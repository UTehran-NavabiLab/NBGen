LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

ENTITY c432 IS
    PORT (
        N1 : IN STD_LOGIC;
        N4 : IN STD_LOGIC;
        N8 : IN STD_LOGIC;
        N11 : IN STD_LOGIC;
        N14 : IN STD_LOGIC;
        N17 : IN STD_LOGIC;
        N21 : IN STD_LOGIC;
        N24 : IN STD_LOGIC;
        N27 : IN STD_LOGIC;
        N30 : IN STD_LOGIC;
        N34 : IN STD_LOGIC;
        N37 : IN STD_LOGIC;
        N40 : IN STD_LOGIC;
        N43 : IN STD_LOGIC;
        N47 : IN STD_LOGIC;
        N50 : IN STD_LOGIC;
        N53 : IN STD_LOGIC;
        N56 : IN STD_LOGIC;
        N60 : IN STD_LOGIC;
        N63 : IN STD_LOGIC;
        N66 : IN STD_LOGIC;
        N69 : IN STD_LOGIC;
        N73 : IN STD_LOGIC;
        N76 : IN STD_LOGIC;
        N79 : IN STD_LOGIC;
        N82 : IN STD_LOGIC;
        N86 : IN STD_LOGIC;
        N89 : IN STD_LOGIC;
        N92 : IN STD_LOGIC;
        N95 : IN STD_LOGIC;
        N99 : IN STD_LOGIC;
        N102 : IN STD_LOGIC;
        N105 : IN STD_LOGIC;
        N108 : IN STD_LOGIC;
        N112 : IN STD_LOGIC;
        N115 : IN STD_LOGIC;
        N223 : OUT STD_LOGIC;
        N329 : OUT STD_LOGIC;
        N370 : OUT STD_LOGIC;
        N421 : OUT STD_LOGIC;
        N430 : OUT STD_LOGIC;
        N431 : OUT STD_LOGIC;
        N432 : OUT STD_LOGIC);
END ENTITY c432;

ARCHITECTURE arch OF c432 IS
    SIGNAL _0_ : STD_LOGIC;
    SIGNAL _100_ : STD_LOGIC;
    SIGNAL _101_ : STD_LOGIC;
    SIGNAL _102_ : STD_LOGIC;
    SIGNAL _103_ : STD_LOGIC;
    SIGNAL _104_ : STD_LOGIC;
    SIGNAL _105_ : STD_LOGIC;
    SIGNAL _106_ : STD_LOGIC;
    SIGNAL _107_ : STD_LOGIC;
    SIGNAL _108_ : STD_LOGIC;
    SIGNAL _109_ : STD_LOGIC;
    SIGNAL _10_ : STD_LOGIC;
    SIGNAL _110_ : STD_LOGIC;
    SIGNAL _111_ : STD_LOGIC;
    SIGNAL _112_ : STD_LOGIC;
    SIGNAL _113_ : STD_LOGIC;
    SIGNAL _114_ : STD_LOGIC;
    SIGNAL _115_ : STD_LOGIC;
    SIGNAL _116_ : STD_LOGIC;
    SIGNAL _117_ : STD_LOGIC;
    SIGNAL _118_ : STD_LOGIC;
    SIGNAL _119_ : STD_LOGIC;
    SIGNAL _11_ : STD_LOGIC;
    SIGNAL _120_ : STD_LOGIC;
    SIGNAL _121_ : STD_LOGIC;
    SIGNAL _122_ : STD_LOGIC;
    SIGNAL _123_ : STD_LOGIC;
    SIGNAL _124_ : STD_LOGIC;
    SIGNAL _125_ : STD_LOGIC;
    SIGNAL _126_ : STD_LOGIC;
    SIGNAL _127_ : STD_LOGIC;
    SIGNAL _128_ : STD_LOGIC;
    SIGNAL _129_ : STD_LOGIC;
    SIGNAL _12_ : STD_LOGIC;
    SIGNAL _130_ : STD_LOGIC;
    SIGNAL _131_ : STD_LOGIC;
    SIGNAL _13_ : STD_LOGIC;
    SIGNAL _14_ : STD_LOGIC;
    SIGNAL _15_ : STD_LOGIC;
    SIGNAL _16_ : STD_LOGIC;
    SIGNAL _17_ : STD_LOGIC;
    SIGNAL _18_ : STD_LOGIC;
    SIGNAL _19_ : STD_LOGIC;
    SIGNAL _1_ : STD_LOGIC;
    SIGNAL _20_ : STD_LOGIC;
    SIGNAL _21_ : STD_LOGIC;
    SIGNAL _22_ : STD_LOGIC;
    SIGNAL _23_ : STD_LOGIC;
    SIGNAL _24_ : STD_LOGIC;
    SIGNAL _25_ : STD_LOGIC;
    SIGNAL _26_ : STD_LOGIC;
    SIGNAL _27_ : STD_LOGIC;
    SIGNAL _28_ : STD_LOGIC;
    SIGNAL _29_ : STD_LOGIC;
    SIGNAL _2_ : STD_LOGIC;
    SIGNAL _30_ : STD_LOGIC;
    SIGNAL _31_ : STD_LOGIC;
    SIGNAL _32_ : STD_LOGIC;
    SIGNAL _33_ : STD_LOGIC;
    SIGNAL _34_ : STD_LOGIC;
    SIGNAL _35_ : STD_LOGIC;
    SIGNAL _36_ : STD_LOGIC;
    SIGNAL _37_ : STD_LOGIC;
    SIGNAL _38_ : STD_LOGIC;
    SIGNAL _39_ : STD_LOGIC;
    SIGNAL _3_ : STD_LOGIC;
    SIGNAL _40_ : STD_LOGIC;
    SIGNAL _41_ : STD_LOGIC;
    SIGNAL _42_ : STD_LOGIC;
    SIGNAL _43_ : STD_LOGIC;
    SIGNAL _44_ : STD_LOGIC;
    SIGNAL _45_ : STD_LOGIC;
    SIGNAL _46_ : STD_LOGIC;
    SIGNAL _47_ : STD_LOGIC;
    SIGNAL _48_ : STD_LOGIC;
    SIGNAL _49_ : STD_LOGIC;
    SIGNAL _4_ : STD_LOGIC;
    SIGNAL _50_ : STD_LOGIC;
    SIGNAL _51_ : STD_LOGIC;
    SIGNAL _52_ : STD_LOGIC;
    SIGNAL _53_ : STD_LOGIC;
    SIGNAL _54_ : STD_LOGIC;
    SIGNAL _55_ : STD_LOGIC;
    SIGNAL _56_ : STD_LOGIC;
    SIGNAL _57_ : STD_LOGIC;
    SIGNAL _58_ : STD_LOGIC;
    SIGNAL _59_ : STD_LOGIC;
    SIGNAL _5_ : STD_LOGIC;
    SIGNAL _60_ : STD_LOGIC;
    SIGNAL _61_ : STD_LOGIC;
    SIGNAL _62_ : STD_LOGIC;
    SIGNAL _63_ : STD_LOGIC;
    SIGNAL _64_ : STD_LOGIC;
    SIGNAL _65_ : STD_LOGIC;
    SIGNAL _66_ : STD_LOGIC;
    SIGNAL _67_ : STD_LOGIC;
    SIGNAL _68_ : STD_LOGIC;
    SIGNAL _69_ : STD_LOGIC;
    SIGNAL _6_ : STD_LOGIC;
    SIGNAL _70_ : STD_LOGIC;
    SIGNAL _71_ : STD_LOGIC;
    SIGNAL _72_ : STD_LOGIC;
    SIGNAL _73_ : STD_LOGIC;
    SIGNAL _74_ : STD_LOGIC;
    SIGNAL _75_ : STD_LOGIC;
    SIGNAL _76_ : STD_LOGIC;
    SIGNAL _77_ : STD_LOGIC;
    SIGNAL _78_ : STD_LOGIC;
    SIGNAL _79_ : STD_LOGIC;
    SIGNAL _7_ : STD_LOGIC;
    SIGNAL _80_ : STD_LOGIC;
    SIGNAL _81_ : STD_LOGIC;
    SIGNAL _82_ : STD_LOGIC;
    SIGNAL _83_ : STD_LOGIC;
    SIGNAL _84_ : STD_LOGIC;
    SIGNAL _85_ : STD_LOGIC;
    SIGNAL _86_ : STD_LOGIC;
    SIGNAL _87_ : STD_LOGIC;
    SIGNAL _88_ : STD_LOGIC;
    SIGNAL _89_ : STD_LOGIC;
    SIGNAL _8_ : STD_LOGIC;
    SIGNAL _90_ : STD_LOGIC;
    SIGNAL _91_ : STD_LOGIC;
    SIGNAL _92_ : STD_LOGIC;
    SIGNAL _93_ : STD_LOGIC;
    SIGNAL _94_ : STD_LOGIC;
    SIGNAL _95_ : STD_LOGIC;
    SIGNAL _96_ : STD_LOGIC;
    SIGNAL _97_ : STD_LOGIC;
    SIGNAL _98_ : STD_LOGIC;
    SIGNAL _99_ : STD_LOGIC;
    SIGNAL _9_ : STD_LOGIC;

BEGIN
INV_X1_1: ENTITY WORK.INV_X1
    PORT MAP (
        A => N56,
        ZN => _69_
    );
NOR2_X1_1: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => _69_,
        A2 => N60,
        ZN => _70_
    );
INV_X1_2: ENTITY WORK.INV_X1
    PORT MAP (
        A => N50,
        ZN => _71_
    );
INV_X1_3: ENTITY WORK.INV_X1
    PORT MAP (
        A => N89,
        ZN => _72_
    );
AOI22_X1_1: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => N95,
        A2 => _72_,
        B1 => _71_,
        B2 => N56,
        ZN => _73_
    );
INV_X1_4: ENTITY WORK.INV_X1
    PORT MAP (
        A => N1,
        ZN => _74_
    );
INV_X1_5: ENTITY WORK.INV_X1
    PORT MAP (
        A => N37,
        ZN => _75_
    );
AOI22_X1_2: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => _74_,
        A2 => N4,
        B1 => _75_,
        B2 => N43,
        ZN => _76_
    );
INV_X1_6: ENTITY WORK.INV_X1
    PORT MAP (
        A => N11,
        ZN => _77_
    );
INV_X1_7: ENTITY WORK.INV_X1
    PORT MAP (
        A => N24,
        ZN => _78_
    );
AOI22_X1_3: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => N30,
        A2 => _78_,
        B1 => _77_,
        B2 => N17,
        ZN => _79_
    );
INV_X1_8: ENTITY WORK.INV_X1
    PORT MAP (
        A => N63,
        ZN => _80_
    );
INV_X1_9: ENTITY WORK.INV_X1
    PORT MAP (
        A => N76,
        ZN => _81_
    );
AOI22_X1_4: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => N82,
        A2 => _81_,
        B1 => _80_,
        B2 => N69,
        ZN => _82_
    );
NAND4_X1_1: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => _79_,
        A2 => _82_,
        A3 => _73_,
        A4 => _76_,
        ZN => _83_
    );
INV_X1_10: ENTITY WORK.INV_X1
    PORT MAP (
        A => N102,
        ZN => _84_
    );
AND2_X1_1: ENTITY WORK.AND2_X1
    PORT MAP (
        A1 => _84_,
        A2 => N108,
        ZN => _85_
    );
OAI21_X1_1: ENTITY WORK.OAI21_X1
    PORT MAP (
        A => N50,
        B1 => _83_,
        B2 => _85_,
        ZN => _86_
    );
NAND2_X1_1: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => _86_,
        A2 => _70_,
        ZN => _87_
    );
INV_X1_11: ENTITY WORK.INV_X1
    PORT MAP (
        A => _87_,
        ZN => _88_
    );
NOR2_X1_2: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => _83_,
        A2 => _85_,
        ZN => _89_
    );
OAI21_X1_2: ENTITY WORK.OAI21_X1
    PORT MAP (
        A => N108,
        B1 => _89_,
        B2 => _84_,
        ZN => _90_
    );
NOR2_X1_3: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => _90_,
        A2 => N112,
        ZN => _91_
    );
INV_X1_12: ENTITY WORK.INV_X1
    PORT MAP (
        A => N43,
        ZN => _92_
    );
NOR2_X1_4: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => _92_,
        A2 => N47,
        ZN => _93_
    );
OAI21_X1_3: ENTITY WORK.OAI21_X1
    PORT MAP (
        A => N37,
        B1 => _83_,
        B2 => _85_,
        ZN => _94_
    );
INV_X1_13: ENTITY WORK.INV_X1
    PORT MAP (
        A => N82,
        ZN => _95_
    );
NOR2_X1_5: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => _95_,
        A2 => N86,
        ZN => _96_
    );
OAI21_X1_4: ENTITY WORK.OAI21_X1
    PORT MAP (
        A => N76,
        B1 => _83_,
        B2 => _85_,
        ZN => _97_
    );
AOI22_X1_5: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => _96_,
        A2 => _97_,
        B1 => _94_,
        B2 => _93_,
        ZN => _98_
    );
INV_X1_14: ENTITY WORK.INV_X1
    PORT MAP (
        A => N69,
        ZN => _99_
    );
NOR2_X1_6: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => _99_,
        A2 => N73,
        ZN => _100_
    );
OAI21_X1_5: ENTITY WORK.OAI21_X1
    PORT MAP (
        A => N63,
        B1 => _83_,
        B2 => _85_,
        ZN => _101_
    );
AOI22_X1_6: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => _70_,
        A2 => _86_,
        B1 => _101_,
        B2 => _100_,
        ZN => _102_
    );
INV_X1_15: ENTITY WORK.INV_X1
    PORT MAP (
        A => N4,
        ZN => _103_
    );
NOR2_X1_7: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => _103_,
        A2 => N8,
        ZN => _104_
    );
OAI21_X1_6: ENTITY WORK.OAI21_X1
    PORT MAP (
        A => N1,
        B1 => _83_,
        B2 => _85_,
        ZN => _105_
    );
INV_X1_16: ENTITY WORK.INV_X1
    PORT MAP (
        A => N17,
        ZN => _106_
    );
NOR2_X1_8: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => _106_,
        A2 => N21,
        ZN => _107_
    );
OAI21_X1_7: ENTITY WORK.OAI21_X1
    PORT MAP (
        A => N11,
        B1 => _83_,
        B2 => _85_,
        ZN => _108_
    );
AOI22_X1_7: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => _107_,
        A2 => _108_,
        B1 => _105_,
        B2 => _104_,
        ZN => _109_
    );
INV_X1_17: ENTITY WORK.INV_X1
    PORT MAP (
        A => N95,
        ZN => _110_
    );
NOR2_X1_9: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => _110_,
        A2 => N99,
        ZN => _111_
    );
OAI21_X1_8: ENTITY WORK.OAI21_X1
    PORT MAP (
        A => N89,
        B1 => _83_,
        B2 => _85_,
        ZN => _112_
    );
INV_X1_18: ENTITY WORK.INV_X1
    PORT MAP (
        A => N30,
        ZN => _113_
    );
NOR2_X1_10: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => _113_,
        A2 => N34,
        ZN => _114_
    );
OAI21_X1_9: ENTITY WORK.OAI21_X1
    PORT MAP (
        A => N24,
        B1 => _83_,
        B2 => _85_,
        ZN => _115_
    );
AOI22_X1_8: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => _114_,
        A2 => _115_,
        B1 => _112_,
        B2 => _111_,
        ZN => _116_
    );
NAND4_X1_2: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => _109_,
        A2 => _116_,
        A3 => _98_,
        A4 => _102_,
        ZN => _117_
    );
NOR2_X1_11: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => _117_,
        A2 => _91_,
        ZN => _118_
    );
NAND2_X1_2: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => _86_,
        A2 => N56,
        ZN => _119_
    );
NOR2_X1_12: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => _119_,
        A2 => N66,
        ZN => _120_
    );
OAI21_X1_10: ENTITY WORK.OAI21_X1
    PORT MAP (
        A => _120_,
        B1 => _118_,
        B2 => _88_,
        ZN => _121_
    );
INV_X1_19: ENTITY WORK.INV_X1
    PORT MAP (
        A => N115,
        ZN => _122_
    );
AOI21_X1_1: ENTITY WORK.AOI21_X1
    PORT MAP (
        A => _90_,
        B1 => _117_,
        B2 => N112,
        ZN => _123_
    );
NAND2_X1_3: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => _123_,
        A2 => _122_,
        ZN => _124_
    );
NAND2_X1_4: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => _108_,
        A2 => _107_,
        ZN => _0_
    );
INV_X1_20: ENTITY WORK.INV_X1
    PORT MAP (
        A => _0_,
        ZN => _1_
    );
NAND2_X1_5: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => _108_,
        A2 => N17,
        ZN => _2_
    );
NOR2_X1_13: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => _2_,
        A2 => N27,
        ZN => _3_
    );
OAI21_X1_11: ENTITY WORK.OAI21_X1
    PORT MAP (
        A => _3_,
        B1 => _118_,
        B2 => _1_,
        ZN => _4_
    );
NAND2_X1_6: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => _105_,
        A2 => _104_,
        ZN => _5_
    );
INV_X1_21: ENTITY WORK.INV_X1
    PORT MAP (
        A => _5_,
        ZN => _6_
    );
NAND2_X1_7: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => _105_,
        A2 => N4,
        ZN => _7_
    );
NOR2_X1_14: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => _7_,
        A2 => N14,
        ZN => _8_
    );
OAI21_X1_12: ENTITY WORK.OAI21_X1
    PORT MAP (
        A => _8_,
        B1 => _118_,
        B2 => _6_,
        ZN => _9_
    );
NAND4_X1_3: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => _4_,
        A2 => _9_,
        A3 => _121_,
        A4 => _124_,
        ZN => _10_
    );
INV_X1_22: ENTITY WORK.INV_X1
    PORT MAP (
        A => N92,
        ZN => _11_
    );
NAND2_X1_8: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => _97_,
        A2 => _96_,
        ZN => _12_
    );
INV_X1_23: ENTITY WORK.INV_X1
    PORT MAP (
        A => _12_,
        ZN => _13_
    );
AND2_X1_2: ENTITY WORK.AND2_X1
    PORT MAP (
        A1 => _97_,
        A2 => N82,
        ZN => _14_
    );
OAI211_X1_1: ENTITY WORK.OAI211_X1
    PORT MAP (
        A => _11_,
        B => _14_,
        C1 => _118_,
        C2 => _13_,
        ZN => _15_
    );
NAND2_X1_9: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => _101_,
        A2 => _100_,
        ZN => _16_
    );
OAI21_X1_13: ENTITY WORK.OAI21_X1
    PORT MAP (
        A => _16_,
        B1 => _117_,
        B2 => _91_,
        ZN => _17_
    );
NAND2_X1_10: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => _101_,
        A2 => N69,
        ZN => _18_
    );
NOR2_X1_15: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => _18_,
        A2 => N79,
        ZN => _19_
    );
NAND2_X1_11: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => _112_,
        A2 => _111_,
        ZN => _20_
    );
OAI21_X1_14: ENTITY WORK.OAI21_X1
    PORT MAP (
        A => _20_,
        B1 => _117_,
        B2 => _91_,
        ZN => _21_
    );
NAND2_X1_12: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => _112_,
        A2 => N95,
        ZN => _22_
    );
NOR2_X1_16: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => _22_,
        A2 => N105,
        ZN => _23_
    );
AOI22_X1_9: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => _19_,
        A2 => _17_,
        B1 => _21_,
        B2 => _23_,
        ZN => _24_
    );
NAND2_X1_13: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => _94_,
        A2 => _93_,
        ZN => _25_
    );
OAI21_X1_15: ENTITY WORK.OAI21_X1
    PORT MAP (
        A => _25_,
        B1 => _117_,
        B2 => _91_,
        ZN => _26_
    );
NAND2_X1_14: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => _94_,
        A2 => N43,
        ZN => _27_
    );
NOR2_X1_17: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => _27_,
        A2 => N53,
        ZN => _28_
    );
NAND2_X1_15: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => _115_,
        A2 => _114_,
        ZN => _29_
    );
OAI21_X1_16: ENTITY WORK.OAI21_X1
    PORT MAP (
        A => _29_,
        B1 => _117_,
        B2 => _91_,
        ZN => _30_
    );
NAND2_X1_16: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => _115_,
        A2 => N30,
        ZN => _31_
    );
NOR2_X1_18: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => _31_,
        A2 => N40,
        ZN => _32_
    );
AOI22_X1_10: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => _28_,
        A2 => _26_,
        B1 => _30_,
        B2 => _32_,
        ZN => _33_
    );
NAND3_X1_1: ENTITY WORK.NAND3_X1
    PORT MAP (
        A1 => _24_,
        A2 => _33_,
        A3 => _15_,
        ZN => _34_
    );
OAI21_X1_17: ENTITY WORK.OAI21_X1
    PORT MAP (
        A => N40,
        B1 => _34_,
        B2 => _10_,
        ZN => _35_
    );
INV_X1_24: ENTITY WORK.INV_X1
    PORT MAP (
        A => _118_,
        ZN => _126_
    );
AOI21_X1_2: ENTITY WORK.AOI21_X1
    PORT MAP (
        A => _31_,
        B1 => _126_,
        B2 => N34,
        ZN => _36_
    );
NAND2_X1_17: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => _35_,
        A2 => _36_,
        ZN => _37_
    );
OAI21_X1_18: ENTITY WORK.OAI21_X1
    PORT MAP (
        A => N27,
        B1 => _34_,
        B2 => _10_,
        ZN => _38_
    );
AOI21_X1_3: ENTITY WORK.AOI21_X1
    PORT MAP (
        A => _2_,
        B1 => _126_,
        B2 => N21,
        ZN => _39_
    );
NAND2_X1_18: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => _38_,
        A2 => _39_,
        ZN => _40_
    );
OAI21_X1_19: ENTITY WORK.OAI21_X1
    PORT MAP (
        A => N66,
        B1 => _34_,
        B2 => _10_,
        ZN => _41_
    );
AOI21_X1_4: ENTITY WORK.AOI21_X1
    PORT MAP (
        A => _119_,
        B1 => _126_,
        B2 => N60,
        ZN => _42_
    );
NAND2_X1_19: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => _41_,
        A2 => _42_,
        ZN => _43_
    );
OAI21_X1_20: ENTITY WORK.OAI21_X1
    PORT MAP (
        A => N53,
        B1 => _34_,
        B2 => _10_,
        ZN => _44_
    );
AOI21_X1_5: ENTITY WORK.AOI21_X1
    PORT MAP (
        A => _27_,
        B1 => _126_,
        B2 => N47,
        ZN => _45_
    );
NAND2_X1_20: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => _44_,
        A2 => _45_,
        ZN => _46_
    );
AND4_X1_1: ENTITY WORK.AND4_X1
    PORT MAP (
        A1 => _37_,
        A2 => _43_,
        A3 => _46_,
        A4 => _40_,
        ZN => _47_
    );
OAI21_X1_21: ENTITY WORK.OAI21_X1
    PORT MAP (
        A => N115,
        B1 => _34_,
        B2 => _10_,
        ZN => _48_
    );
NAND2_X1_21: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => _48_,
        A2 => _123_,
        ZN => _49_
    );
AOI21_X1_6: ENTITY WORK.AOI21_X1
    PORT MAP (
        A => _22_,
        B1 => _126_,
        B2 => N99,
        ZN => _50_
    );
OAI21_X1_22: ENTITY WORK.OAI21_X1
    PORT MAP (
        A => N105,
        B1 => _34_,
        B2 => _10_,
        ZN => _51_
    );
NAND2_X1_22: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => _51_,
        A2 => _50_,
        ZN => _52_
    );
OAI21_X1_23: ENTITY WORK.OAI21_X1
    PORT MAP (
        A => N92,
        B1 => _34_,
        B2 => _10_,
        ZN => _53_
    );
NAND2_X1_23: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => _126_,
        A2 => N86,
        ZN => _54_
    );
NAND3_X1_2: ENTITY WORK.NAND3_X1
    PORT MAP (
        A1 => _53_,
        A2 => _14_,
        A3 => _54_,
        ZN => _55_
    );
AOI21_X1_7: ENTITY WORK.AOI21_X1
    PORT MAP (
        A => _18_,
        B1 => _126_,
        B2 => N73,
        ZN => _56_
    );
OAI21_X1_24: ENTITY WORK.OAI21_X1
    PORT MAP (
        A => N79,
        B1 => _34_,
        B2 => _10_,
        ZN => _57_
    );
NAND2_X1_24: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => _57_,
        A2 => _56_,
        ZN => _58_
    );
AND4_X1_2: ENTITY WORK.AND4_X1
    PORT MAP (
        A1 => _49_,
        A2 => _55_,
        A3 => _58_,
        A4 => _52_,
        ZN => _59_
    );
OR2_X1_1: ENTITY WORK.OR2_X1
    PORT MAP (
        A1 => _34_,
        A2 => _10_,
        ZN => _127_
    );
AND2_X1_3: ENTITY WORK.AND2_X1
    PORT MAP (
        A1 => _126_,
        A2 => N8,
        ZN => _60_
    );
AOI211_X1_1: ENTITY WORK.AOI211_X1
    PORT MAP (
        A => _7_,
        B => _60_,
        C1 => _127_,
        C2 => N14,
        ZN => _61_
    );
AOI21_X1_8: ENTITY WORK.AOI21_X1
    PORT MAP (
        A => _61_,
        B1 => _59_,
        B2 => _47_,
        ZN => _128_
    );
INV_X1_25: ENTITY WORK.INV_X1
    PORT MAP (
        A => _47_,
        ZN => _129_
    );
AND2_X1_4: ENTITY WORK.AND2_X1
    PORT MAP (
        A1 => _40_,
        A2 => _37_,
        ZN => _62_
    );
NAND2_X1_25: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => _43_,
        A2 => _46_,
        ZN => _63_
    );
INV_X1_26: ENTITY WORK.INV_X1
    PORT MAP (
        A => _58_,
        ZN => _64_
    );
NAND4_X1_4: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => _64_,
        A2 => _46_,
        A3 => _43_,
        A4 => _37_,
        ZN => _65_
    );
OAI211_X1_2: ENTITY WORK.OAI211_X1
    PORT MAP (
        A => _65_,
        B => _62_,
        C1 => _63_,
        C2 => _55_,
        ZN => _130_
    );
NAND3_X1_3: ENTITY WORK.NAND3_X1
    PORT MAP (
        A1 => _55_,
        A2 => _37_,
        A3 => _46_,
        ZN => _66_
    );
AND2_X1_5: ENTITY WORK.AND2_X1
    PORT MAP (
        A1 => _44_,
        A2 => _45_,
        ZN => _67_
    );
AOI22_X1_11: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => _67_,
        A2 => _37_,
        B1 => _38_,
        B2 => _39_,
        ZN => _68_
    );
OAI211_X1_3: ENTITY WORK.OAI211_X1
    PORT MAP (
        A => _65_,
        B => _68_,
        C1 => _52_,
        C2 => _66_,
        ZN => _131_
    );
INV_X1_27: ENTITY WORK.INV_X1
    PORT MAP (
        A => _89_,
        ZN => _125_
    );
BUF_X1_1: ENTITY WORK.BUF_X1
    PORT MAP (
        A => _125_,
        Z => N223
    );
BUF_X1_2: ENTITY WORK.BUF_X1
    PORT MAP (
        A => _126_,
        Z => N329
    );
BUF_X1_3: ENTITY WORK.BUF_X1
    PORT MAP (
        A => _127_,
        Z => N370
    );
BUF_X1_4: ENTITY WORK.BUF_X1
    PORT MAP (
        A => _128_,
        Z => N421
    );
BUF_X1_5: ENTITY WORK.BUF_X1
    PORT MAP (
        A => _129_,
        Z => N430
    );
BUF_X1_6: ENTITY WORK.BUF_X1
    PORT MAP (
        A => _130_,
        Z => N431
    );
BUF_X1_7: ENTITY WORK.BUF_X1
    PORT MAP (
        A => _131_,
        Z => N432
    );

END ARCHITECTURE arch;
