LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

ENTITY Puneh_Top IS
    PORT (
        clk : IN STD_LOGIC;
        rst : IN STD_LOGIC;
        dataBus : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
        readMEM : OUT STD_LOGIC;
        writeMEM : OUT STD_LOGIC;
        addrBus : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
        dataBus_out : OUT STD_LOGIC_VECTOR (15 DOWNTO 0));
END ENTITY Puneh_Top;

ARCHITECTURE arch OF Puneh_Top IS
    SIGNAL S0 : STD_LOGIC;
    SIGNAL S1 : STD_LOGIC;
    SIGNAL S2 : STD_LOGIC;
    SIGNAL S3 : STD_LOGIC;
    SIGNAL S4 : STD_LOGIC;
    SIGNAL S5 : STD_LOGIC;
    SIGNAL S6 : STD_LOGIC;
    SIGNAL S7 : STD_LOGIC;
    SIGNAL S8 : STD_LOGIC;
    SIGNAL S9 : STD_LOGIC;
    SIGNAL S10 : STD_LOGIC;
    SIGNAL S11 : STD_LOGIC;
    SIGNAL S12 : STD_LOGIC;
    SIGNAL S13 : STD_LOGIC;
    SIGNAL S14 : STD_LOGIC;
    SIGNAL S15 : STD_LOGIC;
    SIGNAL S16 : STD_LOGIC;
    SIGNAL S17 : STD_LOGIC;
    SIGNAL S18 : STD_LOGIC;
    SIGNAL S19 : STD_LOGIC;
    SIGNAL S20 : STD_LOGIC;
    SIGNAL S21 : STD_LOGIC;
    SIGNAL S22 : STD_LOGIC;
    SIGNAL S23 : STD_LOGIC;
    SIGNAL S24 : STD_LOGIC;
    SIGNAL S25 : STD_LOGIC;
    SIGNAL S26 : STD_LOGIC;
    SIGNAL S27 : STD_LOGIC;
    SIGNAL S28 : STD_LOGIC;
    SIGNAL S29 : STD_LOGIC;
    SIGNAL S30 : STD_LOGIC;
    SIGNAL S31 : STD_LOGIC;
    SIGNAL S32 : STD_LOGIC;
    SIGNAL S33 : STD_LOGIC;
    SIGNAL S34 : STD_LOGIC;
    SIGNAL S35 : STD_LOGIC;
    SIGNAL S36 : STD_LOGIC;
    SIGNAL S37 : STD_LOGIC;
    SIGNAL S38 : STD_LOGIC;
    SIGNAL S39 : STD_LOGIC;
    SIGNAL S40 : STD_LOGIC;
    SIGNAL S41 : STD_LOGIC;
    SIGNAL S42 : STD_LOGIC;
    SIGNAL S43 : STD_LOGIC;
    SIGNAL S44 : STD_LOGIC;
    SIGNAL S45 : STD_LOGIC;
    SIGNAL S46 : STD_LOGIC;
    SIGNAL S47 : STD_LOGIC;
    SIGNAL S48 : STD_LOGIC;
    SIGNAL S49 : STD_LOGIC;
    SIGNAL S50 : STD_LOGIC;
    SIGNAL S51 : STD_LOGIC;
    SIGNAL S52 : STD_LOGIC;
    SIGNAL S53 : STD_LOGIC;
    SIGNAL S54 : STD_LOGIC;
    SIGNAL S55 : STD_LOGIC;
    SIGNAL S56 : STD_LOGIC;
    SIGNAL S57 : STD_LOGIC;
    SIGNAL S58 : STD_LOGIC;
    SIGNAL S59 : STD_LOGIC;
    SIGNAL S60 : STD_LOGIC;
    SIGNAL S61 : STD_LOGIC;
    SIGNAL S62 : STD_LOGIC;
    SIGNAL S63 : STD_LOGIC;
    SIGNAL S64 : STD_LOGIC;
    SIGNAL S65 : STD_LOGIC;
    SIGNAL S66 : STD_LOGIC;
    SIGNAL S67 : STD_LOGIC;
    SIGNAL S68 : STD_LOGIC;
    SIGNAL S69 : STD_LOGIC;
    SIGNAL S70 : STD_LOGIC;
    SIGNAL S71 : STD_LOGIC;
    SIGNAL S72 : STD_LOGIC;
    SIGNAL S73 : STD_LOGIC;
    SIGNAL S74 : STD_LOGIC;
    SIGNAL S75 : STD_LOGIC;
    SIGNAL S76 : STD_LOGIC;
    SIGNAL S77 : STD_LOGIC;
    SIGNAL S78 : STD_LOGIC;
    SIGNAL S79 : STD_LOGIC;
    SIGNAL S80 : STD_LOGIC;
    SIGNAL S81 : STD_LOGIC;
    SIGNAL S82 : STD_LOGIC;
    SIGNAL S83 : STD_LOGIC;
    SIGNAL S84 : STD_LOGIC;
    SIGNAL S85 : STD_LOGIC;
    SIGNAL S86 : STD_LOGIC;
    SIGNAL S87 : STD_LOGIC;
    SIGNAL S88 : STD_LOGIC;
    SIGNAL S89 : STD_LOGIC;
    SIGNAL S90 : STD_LOGIC;
    SIGNAL S91 : STD_LOGIC;
    SIGNAL S92 : STD_LOGIC;
    SIGNAL S93 : STD_LOGIC;
    SIGNAL S94 : STD_LOGIC;
    SIGNAL S95 : STD_LOGIC;
    SIGNAL S96 : STD_LOGIC;
    SIGNAL S97 : STD_LOGIC;
    SIGNAL S98 : STD_LOGIC;
    SIGNAL S99 : STD_LOGIC;
    SIGNAL S100 : STD_LOGIC;
    SIGNAL S101 : STD_LOGIC;
    SIGNAL S102 : STD_LOGIC;
    SIGNAL S103 : STD_LOGIC;
    SIGNAL S104 : STD_LOGIC;
    SIGNAL S105 : STD_LOGIC;
    SIGNAL S106 : STD_LOGIC;
    SIGNAL S107 : STD_LOGIC;
    SIGNAL S108 : STD_LOGIC;
    SIGNAL S109 : STD_LOGIC;
    SIGNAL S110 : STD_LOGIC;
    SIGNAL S111 : STD_LOGIC;
    SIGNAL S112 : STD_LOGIC;
    SIGNAL S113 : STD_LOGIC;
    SIGNAL S114 : STD_LOGIC;
    SIGNAL S115 : STD_LOGIC;
    SIGNAL S116 : STD_LOGIC;
    SIGNAL S117 : STD_LOGIC;
    SIGNAL S118 : STD_LOGIC;
    SIGNAL S119 : STD_LOGIC;
    SIGNAL S120 : STD_LOGIC;
    SIGNAL S121 : STD_LOGIC;
    SIGNAL S122 : STD_LOGIC;
    SIGNAL S123 : STD_LOGIC;
    SIGNAL S124 : STD_LOGIC;
    SIGNAL S125 : STD_LOGIC;
    SIGNAL S126 : STD_LOGIC;
    SIGNAL S127 : STD_LOGIC;
    SIGNAL S128 : STD_LOGIC;
    SIGNAL S129 : STD_LOGIC;
    SIGNAL S130 : STD_LOGIC;
    SIGNAL S131 : STD_LOGIC;
    SIGNAL S132 : STD_LOGIC;
    SIGNAL S133 : STD_LOGIC;
    SIGNAL S134 : STD_LOGIC;
    SIGNAL S135 : STD_LOGIC;
    SIGNAL S136 : STD_LOGIC;
    SIGNAL S137 : STD_LOGIC;
    SIGNAL S138 : STD_LOGIC;
    SIGNAL S139 : STD_LOGIC;
    SIGNAL S140 : STD_LOGIC;
    SIGNAL S141 : STD_LOGIC;
    SIGNAL S142 : STD_LOGIC;
    SIGNAL S143 : STD_LOGIC;
    SIGNAL S144 : STD_LOGIC;
    SIGNAL S145 : STD_LOGIC;
    SIGNAL S146 : STD_LOGIC;
    SIGNAL S147 : STD_LOGIC;
    SIGNAL S148 : STD_LOGIC;
    SIGNAL S149 : STD_LOGIC;
    SIGNAL S150 : STD_LOGIC;
    SIGNAL S151 : STD_LOGIC;
    SIGNAL S152 : STD_LOGIC;
    SIGNAL S153 : STD_LOGIC;
    SIGNAL S154 : STD_LOGIC;
    SIGNAL S155 : STD_LOGIC;
    SIGNAL S156 : STD_LOGIC;
    SIGNAL S157 : STD_LOGIC;
    SIGNAL S158 : STD_LOGIC;
    SIGNAL S159 : STD_LOGIC;
    SIGNAL S160 : STD_LOGIC;
    SIGNAL S161 : STD_LOGIC;
    SIGNAL S162 : STD_LOGIC;
    SIGNAL S163 : STD_LOGIC;
    SIGNAL S164 : STD_LOGIC;
    SIGNAL S165 : STD_LOGIC;
    SIGNAL S166 : STD_LOGIC;
    SIGNAL S167 : STD_LOGIC;
    SIGNAL S168 : STD_LOGIC;
    SIGNAL S169 : STD_LOGIC;
    SIGNAL S170 : STD_LOGIC;
    SIGNAL S171 : STD_LOGIC;
    SIGNAL S172 : STD_LOGIC;
    SIGNAL S173 : STD_LOGIC;
    SIGNAL S174 : STD_LOGIC;
    SIGNAL S175 : STD_LOGIC;
    SIGNAL S176 : STD_LOGIC;
    SIGNAL S177 : STD_LOGIC;
    SIGNAL S178 : STD_LOGIC;
    SIGNAL S179 : STD_LOGIC;
    SIGNAL S180 : STD_LOGIC;
    SIGNAL S181 : STD_LOGIC;
    SIGNAL S182 : STD_LOGIC;
    SIGNAL S183 : STD_LOGIC;
    SIGNAL S184 : STD_LOGIC;
    SIGNAL S185 : STD_LOGIC;
    SIGNAL S186 : STD_LOGIC;
    SIGNAL S187 : STD_LOGIC;
    SIGNAL S188 : STD_LOGIC;
    SIGNAL S189 : STD_LOGIC;
    SIGNAL S190 : STD_LOGIC;
    SIGNAL S191 : STD_LOGIC;
    SIGNAL S192 : STD_LOGIC;
    SIGNAL S193 : STD_LOGIC;
    SIGNAL S194 : STD_LOGIC;
    SIGNAL S195 : STD_LOGIC;
    SIGNAL S196 : STD_LOGIC;
    SIGNAL S197 : STD_LOGIC;
    SIGNAL S198 : STD_LOGIC;
    SIGNAL S199 : STD_LOGIC;
    SIGNAL S200 : STD_LOGIC;
    SIGNAL S201 : STD_LOGIC;
    SIGNAL S202 : STD_LOGIC;
    SIGNAL S203 : STD_LOGIC;
    SIGNAL S204 : STD_LOGIC;
    SIGNAL S205 : STD_LOGIC;
    SIGNAL S206 : STD_LOGIC;
    SIGNAL S207 : STD_LOGIC;
    SIGNAL S208 : STD_LOGIC;
    SIGNAL S209 : STD_LOGIC;
    SIGNAL S210 : STD_LOGIC;
    SIGNAL S211 : STD_LOGIC;
    SIGNAL S212 : STD_LOGIC;
    SIGNAL S213 : STD_LOGIC;
    SIGNAL S214 : STD_LOGIC;
    SIGNAL S215 : STD_LOGIC;
    SIGNAL S216 : STD_LOGIC;
    SIGNAL S217 : STD_LOGIC;
    SIGNAL S218 : STD_LOGIC;
    SIGNAL S219 : STD_LOGIC;
    SIGNAL S220 : STD_LOGIC;
    SIGNAL S221 : STD_LOGIC;
    SIGNAL S222 : STD_LOGIC;
    SIGNAL S223 : STD_LOGIC;
    SIGNAL S224 : STD_LOGIC;
    SIGNAL S225 : STD_LOGIC;
    SIGNAL S226 : STD_LOGIC;
    SIGNAL S227 : STD_LOGIC;
    SIGNAL S228 : STD_LOGIC;
    SIGNAL S229 : STD_LOGIC;
    SIGNAL S230 : STD_LOGIC;
    SIGNAL S231 : STD_LOGIC;
    SIGNAL S232 : STD_LOGIC;
    SIGNAL S233 : STD_LOGIC;
    SIGNAL S234 : STD_LOGIC;
    SIGNAL S235 : STD_LOGIC;
    SIGNAL S236 : STD_LOGIC;
    SIGNAL S237 : STD_LOGIC;
    SIGNAL S238 : STD_LOGIC;
    SIGNAL S239 : STD_LOGIC;
    SIGNAL S240 : STD_LOGIC;
    SIGNAL S241 : STD_LOGIC;
    SIGNAL S242 : STD_LOGIC;
    SIGNAL S243 : STD_LOGIC;
    SIGNAL S244 : STD_LOGIC;
    SIGNAL S245 : STD_LOGIC;
    SIGNAL S246 : STD_LOGIC;
    SIGNAL S247 : STD_LOGIC;
    SIGNAL S248 : STD_LOGIC;
    SIGNAL S249 : STD_LOGIC;
    SIGNAL S250 : STD_LOGIC;
    SIGNAL S251 : STD_LOGIC;
    SIGNAL S252 : STD_LOGIC;
    SIGNAL S253 : STD_LOGIC;
    SIGNAL S254 : STD_LOGIC;
    SIGNAL S255 : STD_LOGIC;
    SIGNAL S256 : STD_LOGIC;
    SIGNAL S257 : STD_LOGIC;
    SIGNAL S258 : STD_LOGIC;
    SIGNAL S259 : STD_LOGIC;
    SIGNAL S260 : STD_LOGIC;
    SIGNAL S261 : STD_LOGIC;
    SIGNAL S262 : STD_LOGIC;
    SIGNAL S263 : STD_LOGIC;
    SIGNAL S264 : STD_LOGIC;
    SIGNAL S265 : STD_LOGIC;
    SIGNAL S266 : STD_LOGIC;
    SIGNAL S267 : STD_LOGIC;
    SIGNAL S268 : STD_LOGIC;
    SIGNAL S269 : STD_LOGIC;
    SIGNAL S270 : STD_LOGIC;
    SIGNAL S271 : STD_LOGIC;
    SIGNAL S272 : STD_LOGIC;
    SIGNAL S273 : STD_LOGIC;
    SIGNAL S274 : STD_LOGIC;
    SIGNAL S275 : STD_LOGIC;
    SIGNAL S276 : STD_LOGIC;
    SIGNAL S277 : STD_LOGIC;
    SIGNAL S278 : STD_LOGIC;
    SIGNAL S279 : STD_LOGIC;
    SIGNAL S280 : STD_LOGIC;
    SIGNAL S281 : STD_LOGIC;
    SIGNAL S282 : STD_LOGIC;
    SIGNAL S283 : STD_LOGIC;
    SIGNAL S284 : STD_LOGIC;
    SIGNAL S285 : STD_LOGIC;
    SIGNAL S286 : STD_LOGIC;
    SIGNAL S287 : STD_LOGIC;
    SIGNAL S288 : STD_LOGIC;
    SIGNAL S289 : STD_LOGIC;
    SIGNAL S290 : STD_LOGIC;
    SIGNAL S291 : STD_LOGIC;
    SIGNAL S292 : STD_LOGIC;
    SIGNAL S293 : STD_LOGIC;
    SIGNAL S294 : STD_LOGIC;
    SIGNAL S295 : STD_LOGIC;
    SIGNAL S296 : STD_LOGIC;
    SIGNAL S297 : STD_LOGIC;
    SIGNAL S298 : STD_LOGIC;
    SIGNAL S299 : STD_LOGIC;
    SIGNAL S300 : STD_LOGIC;
    SIGNAL S301 : STD_LOGIC;
    SIGNAL S302 : STD_LOGIC;
    SIGNAL S303 : STD_LOGIC;
    SIGNAL S304 : STD_LOGIC;
    SIGNAL S305 : STD_LOGIC;
    SIGNAL S306 : STD_LOGIC;
    SIGNAL S307 : STD_LOGIC;
    SIGNAL S308 : STD_LOGIC;
    SIGNAL S309 : STD_LOGIC;
    SIGNAL S310 : STD_LOGIC;
    SIGNAL S311 : STD_LOGIC;
    SIGNAL S312 : STD_LOGIC;
    SIGNAL S313 : STD_LOGIC;
    SIGNAL S314 : STD_LOGIC;
    SIGNAL S315 : STD_LOGIC;
    SIGNAL S316 : STD_LOGIC;
    SIGNAL S317 : STD_LOGIC;
    SIGNAL S318 : STD_LOGIC;
    SIGNAL S319 : STD_LOGIC;
    SIGNAL S320 : STD_LOGIC;
    SIGNAL S321 : STD_LOGIC;
    SIGNAL S322 : STD_LOGIC;
    SIGNAL S323 : STD_LOGIC;
    SIGNAL S324 : STD_LOGIC;
    SIGNAL S325 : STD_LOGIC;
    SIGNAL S326 : STD_LOGIC;
    SIGNAL S327 : STD_LOGIC;
    SIGNAL S328 : STD_LOGIC;
    SIGNAL S329 : STD_LOGIC;
    SIGNAL S330 : STD_LOGIC;
    SIGNAL S331 : STD_LOGIC;
    SIGNAL S332 : STD_LOGIC;
    SIGNAL S333 : STD_LOGIC;
    SIGNAL S334 : STD_LOGIC;
    SIGNAL S335 : STD_LOGIC;
    SIGNAL S336 : STD_LOGIC;
    SIGNAL S337 : STD_LOGIC;
    SIGNAL S338 : STD_LOGIC;
    SIGNAL S339 : STD_LOGIC;
    SIGNAL S340 : STD_LOGIC;
    SIGNAL S341 : STD_LOGIC;
    SIGNAL S342 : STD_LOGIC;
    SIGNAL S343 : STD_LOGIC;
    SIGNAL S344 : STD_LOGIC;
    SIGNAL S345 : STD_LOGIC;
    SIGNAL S346 : STD_LOGIC;
    SIGNAL S347 : STD_LOGIC;
    SIGNAL S348 : STD_LOGIC;
    SIGNAL S349 : STD_LOGIC;
    SIGNAL S350 : STD_LOGIC;
    SIGNAL S351 : STD_LOGIC;
    SIGNAL S352 : STD_LOGIC;
    SIGNAL S353 : STD_LOGIC;
    SIGNAL S354 : STD_LOGIC;
    SIGNAL S355 : STD_LOGIC;
    SIGNAL S356 : STD_LOGIC;
    SIGNAL S357 : STD_LOGIC;
    SIGNAL S358 : STD_LOGIC;
    SIGNAL S359 : STD_LOGIC;
    SIGNAL S360 : STD_LOGIC;
    SIGNAL S361 : STD_LOGIC;
    SIGNAL S362 : STD_LOGIC;
    SIGNAL S363 : STD_LOGIC;
    SIGNAL S364 : STD_LOGIC;
    SIGNAL S365 : STD_LOGIC;
    SIGNAL S366 : STD_LOGIC;
    SIGNAL S367 : STD_LOGIC;
    SIGNAL S368 : STD_LOGIC;
    SIGNAL S369 : STD_LOGIC;
    SIGNAL S370 : STD_LOGIC;
    SIGNAL S371 : STD_LOGIC;
    SIGNAL S372 : STD_LOGIC;
    SIGNAL S373 : STD_LOGIC;
    SIGNAL S374 : STD_LOGIC;
    SIGNAL S375 : STD_LOGIC;
    SIGNAL S376 : STD_LOGIC;
    SIGNAL S377 : STD_LOGIC;
    SIGNAL S378 : STD_LOGIC;
    SIGNAL S379 : STD_LOGIC;
    SIGNAL S380 : STD_LOGIC;
    SIGNAL S381 : STD_LOGIC;
    SIGNAL S382 : STD_LOGIC;
    SIGNAL S383 : STD_LOGIC;
    SIGNAL S384 : STD_LOGIC;
    SIGNAL S385 : STD_LOGIC;
    SIGNAL S386 : STD_LOGIC;
    SIGNAL S387 : STD_LOGIC;
    SIGNAL S388 : STD_LOGIC;
    SIGNAL S389 : STD_LOGIC;
    SIGNAL S390 : STD_LOGIC;
    SIGNAL S391 : STD_LOGIC;
    SIGNAL S392 : STD_LOGIC;
    SIGNAL S393 : STD_LOGIC;
    SIGNAL S394 : STD_LOGIC;
    SIGNAL S395 : STD_LOGIC;
    SIGNAL S396 : STD_LOGIC;
    SIGNAL S397 : STD_LOGIC;
    SIGNAL S398 : STD_LOGIC;
    SIGNAL S399 : STD_LOGIC;
    SIGNAL S400 : STD_LOGIC;
    SIGNAL S401 : STD_LOGIC;
    SIGNAL S402 : STD_LOGIC;
    SIGNAL S403 : STD_LOGIC;
    SIGNAL S404 : STD_LOGIC;
    SIGNAL S405 : STD_LOGIC;
    SIGNAL S406 : STD_LOGIC;
    SIGNAL S407 : STD_LOGIC;
    SIGNAL S408 : STD_LOGIC;
    SIGNAL S409 : STD_LOGIC;
    SIGNAL S410 : STD_LOGIC;
    SIGNAL S411 : STD_LOGIC;
    SIGNAL S412 : STD_LOGIC;
    SIGNAL S413 : STD_LOGIC;
    SIGNAL S414 : STD_LOGIC;
    SIGNAL S415 : STD_LOGIC;
    SIGNAL S416 : STD_LOGIC;
    SIGNAL S417 : STD_LOGIC;
    SIGNAL S418 : STD_LOGIC;
    SIGNAL S419 : STD_LOGIC;
    SIGNAL S420 : STD_LOGIC;
    SIGNAL S421 : STD_LOGIC;
    SIGNAL S422 : STD_LOGIC;
    SIGNAL S423 : STD_LOGIC;
    SIGNAL S424 : STD_LOGIC;
    SIGNAL S425 : STD_LOGIC;
    SIGNAL S426 : STD_LOGIC;
    SIGNAL S427 : STD_LOGIC;
    SIGNAL S428 : STD_LOGIC;
    SIGNAL S429 : STD_LOGIC;
    SIGNAL S430 : STD_LOGIC;
    SIGNAL S431 : STD_LOGIC;
    SIGNAL S432 : STD_LOGIC;
    SIGNAL S433 : STD_LOGIC;
    SIGNAL S434 : STD_LOGIC;
    SIGNAL S435 : STD_LOGIC;
    SIGNAL S436 : STD_LOGIC;
    SIGNAL S437 : STD_LOGIC;
    SIGNAL S438 : STD_LOGIC;
    SIGNAL S439 : STD_LOGIC;
    SIGNAL S440 : STD_LOGIC;
    SIGNAL S441 : STD_LOGIC;
    SIGNAL S442 : STD_LOGIC;
    SIGNAL S443 : STD_LOGIC;
    SIGNAL S444 : STD_LOGIC;
    SIGNAL S445 : STD_LOGIC;
    SIGNAL S446 : STD_LOGIC;
    SIGNAL S447 : STD_LOGIC;
    SIGNAL S448 : STD_LOGIC;
    SIGNAL S449 : STD_LOGIC;
    SIGNAL S450 : STD_LOGIC;
    SIGNAL S451 : STD_LOGIC;
    SIGNAL S452 : STD_LOGIC;
    SIGNAL S453 : STD_LOGIC;
    SIGNAL S454 : STD_LOGIC;
    SIGNAL S455 : STD_LOGIC;
    SIGNAL S456 : STD_LOGIC;
    SIGNAL S457 : STD_LOGIC;
    SIGNAL S458 : STD_LOGIC;
    SIGNAL S459 : STD_LOGIC;
    SIGNAL S460 : STD_LOGIC;
    SIGNAL S461 : STD_LOGIC;
    SIGNAL S462 : STD_LOGIC;
    SIGNAL S463 : STD_LOGIC;
    SIGNAL S464 : STD_LOGIC;
    SIGNAL S465 : STD_LOGIC;
    SIGNAL S466 : STD_LOGIC;
    SIGNAL S467 : STD_LOGIC;
    SIGNAL S468 : STD_LOGIC;
    SIGNAL S469 : STD_LOGIC;
    SIGNAL S470 : STD_LOGIC;
    SIGNAL S471 : STD_LOGIC;
    SIGNAL S472 : STD_LOGIC;
    SIGNAL S473 : STD_LOGIC;
    SIGNAL S474 : STD_LOGIC;
    SIGNAL S475 : STD_LOGIC;
    SIGNAL S476 : STD_LOGIC;
    SIGNAL S477 : STD_LOGIC;
    SIGNAL S478 : STD_LOGIC;
    SIGNAL S479 : STD_LOGIC;
    SIGNAL S480 : STD_LOGIC;
    SIGNAL S481 : STD_LOGIC;
    SIGNAL S482 : STD_LOGIC;
    SIGNAL S483 : STD_LOGIC;
    SIGNAL S484 : STD_LOGIC;
    SIGNAL S485 : STD_LOGIC;
    SIGNAL S486 : STD_LOGIC;
    SIGNAL S487 : STD_LOGIC;
    SIGNAL S488 : STD_LOGIC;
    SIGNAL S489 : STD_LOGIC;
    SIGNAL S490 : STD_LOGIC;
    SIGNAL S491 : STD_LOGIC;
    SIGNAL S492 : STD_LOGIC;
    SIGNAL S493 : STD_LOGIC;
    SIGNAL S494 : STD_LOGIC;
    SIGNAL S495 : STD_LOGIC;
    SIGNAL S496 : STD_LOGIC;
    SIGNAL S497 : STD_LOGIC;
    SIGNAL S498 : STD_LOGIC;
    SIGNAL S499 : STD_LOGIC;
    SIGNAL S500 : STD_LOGIC;
    SIGNAL S501 : STD_LOGIC;
    SIGNAL S502 : STD_LOGIC;
    SIGNAL S503 : STD_LOGIC;
    SIGNAL S504 : STD_LOGIC;
    SIGNAL S505 : STD_LOGIC;
    SIGNAL S506 : STD_LOGIC;
    SIGNAL S507 : STD_LOGIC;
    SIGNAL S508 : STD_LOGIC;
    SIGNAL S509 : STD_LOGIC;
    SIGNAL S510 : STD_LOGIC;
    SIGNAL S511 : STD_LOGIC;
    SIGNAL S512 : STD_LOGIC;
    SIGNAL S513 : STD_LOGIC;
    SIGNAL S514 : STD_LOGIC;
    SIGNAL S515 : STD_LOGIC;
    SIGNAL S516 : STD_LOGIC;
    SIGNAL S517 : STD_LOGIC;
    SIGNAL S518 : STD_LOGIC;
    SIGNAL S519 : STD_LOGIC;
    SIGNAL S520 : STD_LOGIC;
    SIGNAL S521 : STD_LOGIC;
    SIGNAL S522 : STD_LOGIC;
    SIGNAL S523 : STD_LOGIC;
    SIGNAL S524 : STD_LOGIC;
    SIGNAL S525 : STD_LOGIC;
    SIGNAL S526 : STD_LOGIC;
    SIGNAL S527 : STD_LOGIC;
    SIGNAL S528 : STD_LOGIC;
    SIGNAL S529 : STD_LOGIC;
    SIGNAL S530 : STD_LOGIC;
    SIGNAL S531 : STD_LOGIC;
    SIGNAL S532 : STD_LOGIC;
    SIGNAL S533 : STD_LOGIC;
    SIGNAL S534 : STD_LOGIC;
    SIGNAL S535 : STD_LOGIC;
    SIGNAL S536 : STD_LOGIC;
    SIGNAL S537 : STD_LOGIC;
    SIGNAL S538 : STD_LOGIC;
    SIGNAL S539 : STD_LOGIC;
    SIGNAL S540 : STD_LOGIC;
    SIGNAL S541 : STD_LOGIC;
    SIGNAL S542 : STD_LOGIC;
    SIGNAL S543 : STD_LOGIC;
    SIGNAL S544 : STD_LOGIC;
    SIGNAL S545 : STD_LOGIC;
    SIGNAL S546 : STD_LOGIC;
    SIGNAL S547 : STD_LOGIC;
    SIGNAL S548 : STD_LOGIC;
    SIGNAL S549 : STD_LOGIC;
    SIGNAL S550 : STD_LOGIC;
    SIGNAL S551 : STD_LOGIC;
    SIGNAL S552 : STD_LOGIC;
    SIGNAL S553 : STD_LOGIC;
    SIGNAL S554 : STD_LOGIC;
    SIGNAL S555 : STD_LOGIC;
    SIGNAL S556 : STD_LOGIC;
    SIGNAL S557 : STD_LOGIC;
    SIGNAL S558 : STD_LOGIC;
    SIGNAL S559 : STD_LOGIC;
    SIGNAL S560 : STD_LOGIC;
    SIGNAL S561 : STD_LOGIC;
    SIGNAL S562 : STD_LOGIC;
    SIGNAL S563 : STD_LOGIC;
    SIGNAL S564 : STD_LOGIC;
    SIGNAL S565 : STD_LOGIC;
    SIGNAL S566 : STD_LOGIC;
    SIGNAL S567 : STD_LOGIC;
    SIGNAL S568 : STD_LOGIC;
    SIGNAL S569 : STD_LOGIC;
    SIGNAL S570 : STD_LOGIC;
    SIGNAL S571 : STD_LOGIC;
    SIGNAL S572 : STD_LOGIC;
    SIGNAL S573 : STD_LOGIC;
    SIGNAL S574 : STD_LOGIC;
    SIGNAL S575 : STD_LOGIC;
    SIGNAL S576 : STD_LOGIC;
    SIGNAL S577 : STD_LOGIC;
    SIGNAL S578 : STD_LOGIC;
    SIGNAL S579 : STD_LOGIC;
    SIGNAL S580 : STD_LOGIC;
    SIGNAL S581 : STD_LOGIC;
    SIGNAL S582 : STD_LOGIC;
    SIGNAL S583 : STD_LOGIC;
    SIGNAL S584 : STD_LOGIC;
    SIGNAL S585 : STD_LOGIC;
    SIGNAL S586 : STD_LOGIC;
    SIGNAL S587 : STD_LOGIC;
    SIGNAL S588 : STD_LOGIC;
    SIGNAL S589 : STD_LOGIC;
    SIGNAL S590 : STD_LOGIC;
    SIGNAL S591 : STD_LOGIC;
    SIGNAL S592 : STD_LOGIC;
    SIGNAL S593 : STD_LOGIC;
    SIGNAL S594 : STD_LOGIC;
    SIGNAL S595 : STD_LOGIC;
    SIGNAL S596 : STD_LOGIC;
    SIGNAL S597 : STD_LOGIC;
    SIGNAL S598 : STD_LOGIC;
    SIGNAL S599 : STD_LOGIC;
    SIGNAL S600 : STD_LOGIC;
    SIGNAL S601 : STD_LOGIC;
    SIGNAL S602 : STD_LOGIC;
    SIGNAL S603 : STD_LOGIC;
    SIGNAL S604 : STD_LOGIC;
    SIGNAL S605 : STD_LOGIC;
    SIGNAL S606 : STD_LOGIC;
    SIGNAL S607 : STD_LOGIC;
    SIGNAL S608 : STD_LOGIC;
    SIGNAL S609 : STD_LOGIC;
    SIGNAL S610 : STD_LOGIC;
    SIGNAL S611 : STD_LOGIC;
    SIGNAL S612 : STD_LOGIC;
    SIGNAL S613 : STD_LOGIC;
    SIGNAL S614 : STD_LOGIC;
    SIGNAL S615 : STD_LOGIC;
    SIGNAL S616 : STD_LOGIC;
    SIGNAL S617 : STD_LOGIC;
    SIGNAL S618 : STD_LOGIC;
    SIGNAL S619 : STD_LOGIC;
    SIGNAL S620 : STD_LOGIC;
    SIGNAL S621 : STD_LOGIC;
    SIGNAL S622 : STD_LOGIC;
    SIGNAL S623 : STD_LOGIC;
    SIGNAL S624 : STD_LOGIC;
    SIGNAL S625 : STD_LOGIC;
    SIGNAL S626 : STD_LOGIC;
    SIGNAL S627 : STD_LOGIC;
    SIGNAL S628 : STD_LOGIC;
    SIGNAL S629 : STD_LOGIC;
    SIGNAL S630 : STD_LOGIC;
    SIGNAL S631 : STD_LOGIC;
    SIGNAL S632 : STD_LOGIC;
    SIGNAL S633 : STD_LOGIC;
    SIGNAL S634 : STD_LOGIC;
    SIGNAL S635 : STD_LOGIC;
    SIGNAL S636 : STD_LOGIC;
    SIGNAL S637 : STD_LOGIC;
    SIGNAL S638 : STD_LOGIC;
    SIGNAL S639 : STD_LOGIC;
    SIGNAL S640 : STD_LOGIC;
    SIGNAL S641 : STD_LOGIC;
    SIGNAL S642 : STD_LOGIC;
    SIGNAL S643 : STD_LOGIC;
    SIGNAL S644 : STD_LOGIC;
    SIGNAL S645 : STD_LOGIC;
    SIGNAL S646 : STD_LOGIC;
    SIGNAL S647 : STD_LOGIC;
    SIGNAL S648 : STD_LOGIC;
    SIGNAL S649 : STD_LOGIC;
    SIGNAL S650 : STD_LOGIC;
    SIGNAL S651 : STD_LOGIC;
    SIGNAL S652 : STD_LOGIC;
    SIGNAL S653 : STD_LOGIC;
    SIGNAL S654 : STD_LOGIC;
    SIGNAL S655 : STD_LOGIC;
    SIGNAL S656 : STD_LOGIC;
    SIGNAL S657 : STD_LOGIC;
    SIGNAL S658 : STD_LOGIC;
    SIGNAL S659 : STD_LOGIC;
    SIGNAL S660 : STD_LOGIC;
    SIGNAL S661 : STD_LOGIC;
    SIGNAL S662 : STD_LOGIC;
    SIGNAL S663 : STD_LOGIC;
    SIGNAL S664 : STD_LOGIC;
    SIGNAL S665 : STD_LOGIC;
    SIGNAL S666 : STD_LOGIC;
    SIGNAL S667 : STD_LOGIC;
    SIGNAL S668 : STD_LOGIC;
    SIGNAL S669 : STD_LOGIC;
    SIGNAL S670 : STD_LOGIC;
    SIGNAL S671 : STD_LOGIC;
    SIGNAL S672 : STD_LOGIC;
    SIGNAL S673 : STD_LOGIC;
    SIGNAL S674 : STD_LOGIC;
    SIGNAL S675 : STD_LOGIC;
    SIGNAL S676 : STD_LOGIC;
    SIGNAL S677 : STD_LOGIC;
    SIGNAL S678 : STD_LOGIC;
    SIGNAL S679 : STD_LOGIC;
    SIGNAL S680 : STD_LOGIC;
    SIGNAL S681 : STD_LOGIC;
    SIGNAL S682 : STD_LOGIC;
    SIGNAL S683 : STD_LOGIC;
    SIGNAL S684 : STD_LOGIC;
    SIGNAL S685 : STD_LOGIC;
    SIGNAL S686 : STD_LOGIC;
    SIGNAL S687 : STD_LOGIC;
    SIGNAL S688 : STD_LOGIC;
    SIGNAL S689 : STD_LOGIC;
    SIGNAL S690 : STD_LOGIC;
    SIGNAL S691 : STD_LOGIC;
    SIGNAL S692 : STD_LOGIC;
    SIGNAL S693 : STD_LOGIC;
    SIGNAL S694 : STD_LOGIC;
    SIGNAL S695 : STD_LOGIC;
    SIGNAL S696 : STD_LOGIC;
    SIGNAL S697 : STD_LOGIC;
    SIGNAL S698 : STD_LOGIC;
    SIGNAL S699 : STD_LOGIC;
    SIGNAL S700 : STD_LOGIC;
    SIGNAL S701 : STD_LOGIC;
    SIGNAL S702 : STD_LOGIC;
    SIGNAL S703 : STD_LOGIC;
    SIGNAL S704 : STD_LOGIC;
    SIGNAL S705 : STD_LOGIC;
    SIGNAL S706 : STD_LOGIC;
    SIGNAL S707 : STD_LOGIC;
    SIGNAL S708 : STD_LOGIC;
    SIGNAL S709 : STD_LOGIC;
    SIGNAL S710 : STD_LOGIC;
    SIGNAL S711 : STD_LOGIC;
    SIGNAL S712 : STD_LOGIC;
    SIGNAL S713 : STD_LOGIC;
    SIGNAL S714 : STD_LOGIC;
    SIGNAL S715 : STD_LOGIC;
    SIGNAL S716 : STD_LOGIC;
    SIGNAL S717 : STD_LOGIC;
    SIGNAL S718 : STD_LOGIC;
    SIGNAL S719 : STD_LOGIC;
    SIGNAL S720 : STD_LOGIC;
    SIGNAL S721 : STD_LOGIC;
    SIGNAL S722 : STD_LOGIC;
    SIGNAL S723 : STD_LOGIC;
    SIGNAL S724 : STD_LOGIC;
    SIGNAL S725 : STD_LOGIC;
    SIGNAL S726 : STD_LOGIC;
    SIGNAL S727 : STD_LOGIC;
    SIGNAL S728 : STD_LOGIC;
    SIGNAL S729 : STD_LOGIC;
    SIGNAL S730 : STD_LOGIC;
    SIGNAL S731 : STD_LOGIC;
    SIGNAL S732 : STD_LOGIC;
    SIGNAL S733 : STD_LOGIC;
    SIGNAL S734 : STD_LOGIC;
    SIGNAL S735 : STD_LOGIC;
    SIGNAL S736 : STD_LOGIC;
    SIGNAL S737 : STD_LOGIC;
    SIGNAL S738 : STD_LOGIC;
    SIGNAL S739 : STD_LOGIC;
    SIGNAL S740 : STD_LOGIC;
    SIGNAL S741 : STD_LOGIC;
    SIGNAL S742 : STD_LOGIC;
    SIGNAL S743 : STD_LOGIC;
    SIGNAL S744 : STD_LOGIC;
    SIGNAL S745 : STD_LOGIC;
    SIGNAL S746 : STD_LOGIC;
    SIGNAL S747 : STD_LOGIC;
    SIGNAL S748 : STD_LOGIC;
    SIGNAL S749 : STD_LOGIC;
    SIGNAL S750 : STD_LOGIC;
    SIGNAL S751 : STD_LOGIC;
    SIGNAL S752 : STD_LOGIC;
    SIGNAL S753 : STD_LOGIC;
    SIGNAL S754 : STD_LOGIC;
    SIGNAL S755 : STD_LOGIC;
    SIGNAL S756 : STD_LOGIC;
    SIGNAL S757 : STD_LOGIC;
    SIGNAL S758 : STD_LOGIC;
    SIGNAL S759 : STD_LOGIC;
    SIGNAL S760 : STD_LOGIC;
    SIGNAL S761 : STD_LOGIC;
    SIGNAL S762 : STD_LOGIC;
    SIGNAL S763 : STD_LOGIC;
    SIGNAL S764 : STD_LOGIC;
    SIGNAL S765 : STD_LOGIC;
    SIGNAL S766 : STD_LOGIC;
    SIGNAL S767 : STD_LOGIC;
    SIGNAL S768 : STD_LOGIC;
    SIGNAL S769 : STD_LOGIC;
    SIGNAL S770 : STD_LOGIC;
    SIGNAL S771 : STD_LOGIC;
    SIGNAL S772 : STD_LOGIC;
    SIGNAL S773 : STD_LOGIC;
    SIGNAL S774 : STD_LOGIC;
    SIGNAL S775 : STD_LOGIC;
    SIGNAL S776 : STD_LOGIC;
    SIGNAL S777 : STD_LOGIC;
    SIGNAL S778 : STD_LOGIC;
    SIGNAL S779 : STD_LOGIC;
    SIGNAL S780 : STD_LOGIC;
    SIGNAL S781 : STD_LOGIC;
    SIGNAL S782 : STD_LOGIC;
    SIGNAL S783 : STD_LOGIC;
    SIGNAL S784 : STD_LOGIC;
    SIGNAL S785 : STD_LOGIC;
    SIGNAL S786 : STD_LOGIC;
    SIGNAL S787 : STD_LOGIC;
    SIGNAL S788 : STD_LOGIC;
    SIGNAL S789 : STD_LOGIC;
    SIGNAL S790 : STD_LOGIC;
    SIGNAL S791 : STD_LOGIC;
    SIGNAL S792 : STD_LOGIC;
    SIGNAL S793 : STD_LOGIC;
    SIGNAL S794 : STD_LOGIC;
    SIGNAL S795 : STD_LOGIC;
    SIGNAL S796 : STD_LOGIC;
    SIGNAL S797 : STD_LOGIC;
    SIGNAL S798 : STD_LOGIC;
    SIGNAL S799 : STD_LOGIC;
    SIGNAL S800 : STD_LOGIC;
    SIGNAL S801 : STD_LOGIC;
    SIGNAL S802 : STD_LOGIC;
    SIGNAL S803 : STD_LOGIC;
    SIGNAL S804 : STD_LOGIC;
    SIGNAL S805 : STD_LOGIC;
    SIGNAL S806 : STD_LOGIC;
    SIGNAL S807 : STD_LOGIC;
    SIGNAL S808 : STD_LOGIC;
    SIGNAL S809 : STD_LOGIC;
    SIGNAL S810 : STD_LOGIC;
    SIGNAL S811 : STD_LOGIC;
    SIGNAL S812 : STD_LOGIC;
    SIGNAL S813 : STD_LOGIC;
    SIGNAL S814 : STD_LOGIC;
    SIGNAL S815 : STD_LOGIC;
    SIGNAL S816 : STD_LOGIC;
    SIGNAL S817 : STD_LOGIC;
    SIGNAL S818 : STD_LOGIC;
    SIGNAL S819 : STD_LOGIC;
    SIGNAL S820 : STD_LOGIC;
    SIGNAL S821 : STD_LOGIC;
    SIGNAL S822 : STD_LOGIC;
    SIGNAL S823 : STD_LOGIC;
    SIGNAL S824 : STD_LOGIC;
    SIGNAL S825 : STD_LOGIC;
    SIGNAL S826 : STD_LOGIC;
    SIGNAL S827 : STD_LOGIC;
    SIGNAL S828 : STD_LOGIC;
    SIGNAL S829 : STD_LOGIC;
    SIGNAL S830 : STD_LOGIC;
    SIGNAL S831 : STD_LOGIC;
    SIGNAL S832 : STD_LOGIC;
    SIGNAL S833 : STD_LOGIC;
    SIGNAL S834 : STD_LOGIC;
    SIGNAL S835 : STD_LOGIC;
    SIGNAL S836 : STD_LOGIC;
    SIGNAL S837 : STD_LOGIC;
    SIGNAL S838 : STD_LOGIC;
    SIGNAL S839 : STD_LOGIC;
    SIGNAL S840 : STD_LOGIC;
    SIGNAL S841 : STD_LOGIC;
    SIGNAL S842 : STD_LOGIC;
    SIGNAL S843 : STD_LOGIC;
    SIGNAL S844 : STD_LOGIC;
    SIGNAL S845 : STD_LOGIC;
    SIGNAL S846 : STD_LOGIC;
    SIGNAL S847 : STD_LOGIC;
    SIGNAL S848 : STD_LOGIC;
    SIGNAL S849 : STD_LOGIC;
    SIGNAL S850 : STD_LOGIC;
    SIGNAL S851 : STD_LOGIC;
    SIGNAL S852 : STD_LOGIC;
    SIGNAL S853 : STD_LOGIC;
    SIGNAL S854 : STD_LOGIC;
    SIGNAL S855 : STD_LOGIC;
    SIGNAL S856 : STD_LOGIC;
    SIGNAL S857 : STD_LOGIC;
    SIGNAL S858 : STD_LOGIC;
    SIGNAL S859 : STD_LOGIC;
    SIGNAL S860 : STD_LOGIC;
    SIGNAL S861 : STD_LOGIC;
    SIGNAL S862 : STD_LOGIC;
    SIGNAL S863 : STD_LOGIC;
    SIGNAL S864 : STD_LOGIC;
    SIGNAL S865 : STD_LOGIC;
    SIGNAL S866 : STD_LOGIC;
    SIGNAL S867 : STD_LOGIC;
    SIGNAL S868 : STD_LOGIC;
    SIGNAL S869 : STD_LOGIC;
    SIGNAL S870 : STD_LOGIC;
    SIGNAL S871 : STD_LOGIC;
    SIGNAL S872 : STD_LOGIC;
    SIGNAL S873 : STD_LOGIC;
    SIGNAL S874 : STD_LOGIC;
    SIGNAL S875 : STD_LOGIC;
    SIGNAL S876 : STD_LOGIC;
    SIGNAL S877 : STD_LOGIC;
    SIGNAL S878 : STD_LOGIC;
    SIGNAL S879 : STD_LOGIC;
    SIGNAL S880 : STD_LOGIC;
    SIGNAL S881 : STD_LOGIC;
    SIGNAL S882 : STD_LOGIC;
    SIGNAL S883 : STD_LOGIC;
    SIGNAL S884 : STD_LOGIC;
    SIGNAL S885 : STD_LOGIC;
    SIGNAL S886 : STD_LOGIC;
    SIGNAL S887 : STD_LOGIC;
    SIGNAL S888 : STD_LOGIC;
    SIGNAL S889 : STD_LOGIC;
    SIGNAL S890 : STD_LOGIC;
    SIGNAL S891 : STD_LOGIC;
    SIGNAL S892 : STD_LOGIC;
    SIGNAL S893 : STD_LOGIC;
    SIGNAL S894 : STD_LOGIC;
    SIGNAL S895 : STD_LOGIC;
    SIGNAL S896 : STD_LOGIC;
    SIGNAL S897 : STD_LOGIC;
    SIGNAL S898 : STD_LOGIC;
    SIGNAL S899 : STD_LOGIC;
    SIGNAL S900 : STD_LOGIC;
    SIGNAL S901 : STD_LOGIC;
    SIGNAL S902 : STD_LOGIC;
    SIGNAL S903 : STD_LOGIC;
    SIGNAL S904 : STD_LOGIC;
    SIGNAL S905 : STD_LOGIC;
    SIGNAL S906 : STD_LOGIC;
    SIGNAL S907 : STD_LOGIC;
    SIGNAL S908 : STD_LOGIC;
    SIGNAL S909 : STD_LOGIC;
    SIGNAL S910 : STD_LOGIC;
    SIGNAL S911 : STD_LOGIC;
    SIGNAL S912 : STD_LOGIC;
    SIGNAL S913 : STD_LOGIC;
    SIGNAL S914 : STD_LOGIC;
    SIGNAL S915 : STD_LOGIC;
    SIGNAL S916 : STD_LOGIC;
    SIGNAL S917 : STD_LOGIC;
    SIGNAL S918 : STD_LOGIC;
    SIGNAL S919 : STD_LOGIC;
    SIGNAL S920 : STD_LOGIC;
    SIGNAL S921 : STD_LOGIC;
    SIGNAL S922 : STD_LOGIC;
    SIGNAL S923 : STD_LOGIC;
    SIGNAL S924 : STD_LOGIC;
    SIGNAL S925 : STD_LOGIC;
    SIGNAL S926 : STD_LOGIC;
    SIGNAL S927 : STD_LOGIC;
    SIGNAL S928 : STD_LOGIC;
    SIGNAL S929 : STD_LOGIC;
    SIGNAL S930 : STD_LOGIC;
    SIGNAL S931 : STD_LOGIC;
    SIGNAL S932 : STD_LOGIC;
    SIGNAL S933 : STD_LOGIC;
    SIGNAL S934 : STD_LOGIC;
    SIGNAL S935 : STD_LOGIC;
    SIGNAL S936 : STD_LOGIC;
    SIGNAL S937 : STD_LOGIC;
    SIGNAL S938 : STD_LOGIC;
    SIGNAL S939 : STD_LOGIC;
    SIGNAL S940 : STD_LOGIC;
    SIGNAL S941 : STD_LOGIC;
    SIGNAL S942 : STD_LOGIC;
    SIGNAL S943 : STD_LOGIC;
    SIGNAL S944 : STD_LOGIC;
    SIGNAL S945 : STD_LOGIC;
    SIGNAL S946 : STD_LOGIC;
    SIGNAL S947 : STD_LOGIC;
    SIGNAL S948 : STD_LOGIC;
    SIGNAL S949 : STD_LOGIC;
    SIGNAL S950 : STD_LOGIC;
    SIGNAL S951 : STD_LOGIC;
    SIGNAL S952 : STD_LOGIC;
    SIGNAL S953 : STD_LOGIC;
    SIGNAL S954 : STD_LOGIC;
    SIGNAL S955 : STD_LOGIC;
    SIGNAL S956 : STD_LOGIC;
    SIGNAL S957 : STD_LOGIC;
    SIGNAL S958 : STD_LOGIC;
    SIGNAL S959 : STD_LOGIC;
    SIGNAL S960 : STD_LOGIC;
    SIGNAL S961 : STD_LOGIC;
    SIGNAL S962 : STD_LOGIC;
    SIGNAL S963 : STD_LOGIC;
    SIGNAL S964 : STD_LOGIC;
    SIGNAL S965 : STD_LOGIC;
    SIGNAL S966 : STD_LOGIC;
    SIGNAL S967 : STD_LOGIC;
    SIGNAL S968 : STD_LOGIC;
    SIGNAL S969 : STD_LOGIC;
    SIGNAL S970 : STD_LOGIC;
    SIGNAL S971 : STD_LOGIC;
    SIGNAL S972 : STD_LOGIC;
    SIGNAL S973 : STD_LOGIC;
    SIGNAL S974 : STD_LOGIC;
    SIGNAL S975 : STD_LOGIC;
    SIGNAL S976 : STD_LOGIC;
    SIGNAL S977 : STD_LOGIC;
    SIGNAL S978 : STD_LOGIC;
    SIGNAL S979 : STD_LOGIC;
    SIGNAL S980 : STD_LOGIC;
    SIGNAL S981 : STD_LOGIC;
    SIGNAL S982 : STD_LOGIC;
    SIGNAL S983 : STD_LOGIC;
    SIGNAL S984 : STD_LOGIC;
    SIGNAL S985 : STD_LOGIC;
    SIGNAL S986 : STD_LOGIC;
    SIGNAL S987 : STD_LOGIC;
    SIGNAL S988 : STD_LOGIC;
    SIGNAL S989 : STD_LOGIC;
    SIGNAL S990 : STD_LOGIC;
    SIGNAL S991 : STD_LOGIC;
    SIGNAL S992 : STD_LOGIC;
    SIGNAL S993 : STD_LOGIC;
    SIGNAL S994 : STD_LOGIC;
    SIGNAL S995 : STD_LOGIC;
    SIGNAL S996 : STD_LOGIC;
    SIGNAL S997 : STD_LOGIC;
    SIGNAL S998 : STD_LOGIC;
    SIGNAL S999 : STD_LOGIC;
    SIGNAL S1000 : STD_LOGIC;
    SIGNAL S1001 : STD_LOGIC;
    SIGNAL S1002 : STD_LOGIC;
    SIGNAL S1003 : STD_LOGIC;
    SIGNAL S1004 : STD_LOGIC;
    SIGNAL S1005 : STD_LOGIC;
    SIGNAL S1006 : STD_LOGIC;
    SIGNAL S1007 : STD_LOGIC;
    SIGNAL S1008 : STD_LOGIC;
    SIGNAL S1009 : STD_LOGIC;
    SIGNAL S1010 : STD_LOGIC;
    SIGNAL S1011 : STD_LOGIC;
    SIGNAL S1012 : STD_LOGIC;
    SIGNAL S1013 : STD_LOGIC;
    SIGNAL S1014 : STD_LOGIC;
    SIGNAL S1015 : STD_LOGIC;
    SIGNAL S1016 : STD_LOGIC;
    SIGNAL S1017 : STD_LOGIC;
    SIGNAL S1018 : STD_LOGIC;
    SIGNAL S1019 : STD_LOGIC;
    SIGNAL S1020 : STD_LOGIC;
    SIGNAL S1021 : STD_LOGIC;
    SIGNAL S1022 : STD_LOGIC;
    SIGNAL S1023 : STD_LOGIC;
    SIGNAL S1024 : STD_LOGIC;
    SIGNAL S1025 : STD_LOGIC;
    SIGNAL S1026 : STD_LOGIC;
    SIGNAL S1027 : STD_LOGIC;
    SIGNAL S1028 : STD_LOGIC;
    SIGNAL S1029 : STD_LOGIC;
    SIGNAL S1030 : STD_LOGIC;
    SIGNAL S1031 : STD_LOGIC;
    SIGNAL S1032 : STD_LOGIC;
    SIGNAL S1033 : STD_LOGIC;
    SIGNAL S1034 : STD_LOGIC;
    SIGNAL S1035 : STD_LOGIC;
    SIGNAL S1036 : STD_LOGIC;
    SIGNAL S1037 : STD_LOGIC;
    SIGNAL S1038 : STD_LOGIC;
    SIGNAL S1039 : STD_LOGIC;
    SIGNAL S1040 : STD_LOGIC;
    SIGNAL S1041 : STD_LOGIC;
    SIGNAL S1042 : STD_LOGIC;
    SIGNAL S1043 : STD_LOGIC;
    SIGNAL S1044 : STD_LOGIC;
    SIGNAL S1045 : STD_LOGIC;
    SIGNAL S1046 : STD_LOGIC;
    SIGNAL S1047 : STD_LOGIC;
    SIGNAL S1048 : STD_LOGIC;
    SIGNAL S1049 : STD_LOGIC;
    SIGNAL S1050 : STD_LOGIC;
    SIGNAL S1051 : STD_LOGIC;
    SIGNAL S1052 : STD_LOGIC;
    SIGNAL S1053 : STD_LOGIC;
    SIGNAL S1054 : STD_LOGIC;
    SIGNAL S1055 : STD_LOGIC;
    SIGNAL S1056 : STD_LOGIC;
    SIGNAL S1057 : STD_LOGIC;
    SIGNAL S1058 : STD_LOGIC;
    SIGNAL S1059 : STD_LOGIC;
    SIGNAL S1060 : STD_LOGIC;
    SIGNAL S1061 : STD_LOGIC;
    SIGNAL S1062 : STD_LOGIC;
    SIGNAL S1063 : STD_LOGIC;
    SIGNAL S1064 : STD_LOGIC;
    SIGNAL S1065 : STD_LOGIC;
    SIGNAL S1066 : STD_LOGIC;
    SIGNAL S1067 : STD_LOGIC;
    SIGNAL S1068 : STD_LOGIC;
    SIGNAL S1069 : STD_LOGIC;
    SIGNAL S1070 : STD_LOGIC;
    SIGNAL S1071 : STD_LOGIC;
    SIGNAL S1072 : STD_LOGIC;
    SIGNAL S1073 : STD_LOGIC;
    SIGNAL S1074 : STD_LOGIC;
    SIGNAL S1075 : STD_LOGIC;
    SIGNAL S1076 : STD_LOGIC;
    SIGNAL S1077 : STD_LOGIC;
    SIGNAL S1078 : STD_LOGIC;
    SIGNAL S1079 : STD_LOGIC;
    SIGNAL S1080 : STD_LOGIC;
    SIGNAL S1081 : STD_LOGIC;
    SIGNAL S1082 : STD_LOGIC;
    SIGNAL S1083 : STD_LOGIC;
    SIGNAL S1084 : STD_LOGIC;
    SIGNAL S1085 : STD_LOGIC;
    SIGNAL S1086 : STD_LOGIC;
    SIGNAL S1087 : STD_LOGIC;
    SIGNAL S1088 : STD_LOGIC;
    SIGNAL S1089 : STD_LOGIC;
    SIGNAL S1090 : STD_LOGIC;
    SIGNAL S1091 : STD_LOGIC;
    SIGNAL S1092 : STD_LOGIC;
    SIGNAL S1093 : STD_LOGIC;
    SIGNAL S1094 : STD_LOGIC;
    SIGNAL S1095 : STD_LOGIC;
    SIGNAL S1096 : STD_LOGIC;
    SIGNAL S1097 : STD_LOGIC;
    SIGNAL S1098 : STD_LOGIC;
    SIGNAL S1099 : STD_LOGIC;
    SIGNAL S1100 : STD_LOGIC;
    SIGNAL S1101 : STD_LOGIC;
    SIGNAL S1102 : STD_LOGIC;
    SIGNAL S1103 : STD_LOGIC;
    SIGNAL S1104 : STD_LOGIC;
    SIGNAL S1105 : STD_LOGIC;
    SIGNAL S1106 : STD_LOGIC;
    SIGNAL S1107 : STD_LOGIC;
    SIGNAL S1108 : STD_LOGIC;
    SIGNAL S1109 : STD_LOGIC;
    SIGNAL S1110 : STD_LOGIC;
    SIGNAL S1111 : STD_LOGIC;
    SIGNAL S1112 : STD_LOGIC;
    SIGNAL S1113 : STD_LOGIC;
    SIGNAL S1114 : STD_LOGIC;
    SIGNAL S1115 : STD_LOGIC;
    SIGNAL S1116 : STD_LOGIC;
    SIGNAL S1117 : STD_LOGIC;
    SIGNAL S1118 : STD_LOGIC;
    SIGNAL S1119 : STD_LOGIC;
    SIGNAL S1120 : STD_LOGIC;
    SIGNAL S1121 : STD_LOGIC;
    SIGNAL S1122 : STD_LOGIC;
    SIGNAL S1123 : STD_LOGIC;
    SIGNAL S1124 : STD_LOGIC;
    SIGNAL S1125 : STD_LOGIC;
    SIGNAL S1126 : STD_LOGIC;
    SIGNAL S1127 : STD_LOGIC;
    SIGNAL S1128 : STD_LOGIC;
    SIGNAL S1129 : STD_LOGIC;
    SIGNAL S1130 : STD_LOGIC;
    SIGNAL S1131 : STD_LOGIC;
    SIGNAL S1132 : STD_LOGIC;
    SIGNAL S1133 : STD_LOGIC;
    SIGNAL S1134 : STD_LOGIC;
    SIGNAL S1135 : STD_LOGIC;
    SIGNAL S1136 : STD_LOGIC;
    SIGNAL S1137 : STD_LOGIC;
    SIGNAL S1138 : STD_LOGIC;
    SIGNAL S1139 : STD_LOGIC;
    SIGNAL S1140 : STD_LOGIC;
    SIGNAL S1141 : STD_LOGIC;
    SIGNAL S1142 : STD_LOGIC;
    SIGNAL S1143 : STD_LOGIC;
    SIGNAL S1144 : STD_LOGIC;
    SIGNAL S1145 : STD_LOGIC;
    SIGNAL S1146 : STD_LOGIC;
    SIGNAL S1147 : STD_LOGIC;
    SIGNAL S1148 : STD_LOGIC;
    SIGNAL S1149 : STD_LOGIC;
    SIGNAL S1150 : STD_LOGIC;
    SIGNAL S1151 : STD_LOGIC;
    SIGNAL S1152 : STD_LOGIC;
    SIGNAL S1153 : STD_LOGIC;
    SIGNAL S1154 : STD_LOGIC;
    SIGNAL S1155 : STD_LOGIC;
    SIGNAL S1156 : STD_LOGIC;
    SIGNAL S1157 : STD_LOGIC;
    SIGNAL S1158 : STD_LOGIC;
    SIGNAL S1159 : STD_LOGIC;
    SIGNAL S1160 : STD_LOGIC;
    SIGNAL S1161 : STD_LOGIC;
    SIGNAL S1162 : STD_LOGIC;
    SIGNAL S1163 : STD_LOGIC;
    SIGNAL S1164 : STD_LOGIC;
    SIGNAL S1165 : STD_LOGIC;
    SIGNAL S1166 : STD_LOGIC;
    SIGNAL S1167 : STD_LOGIC;
    SIGNAL S1168 : STD_LOGIC;
    SIGNAL S1169 : STD_LOGIC;
    SIGNAL S1170 : STD_LOGIC;
    SIGNAL S1171 : STD_LOGIC;
    SIGNAL S1172 : STD_LOGIC;
    SIGNAL S1173 : STD_LOGIC;
    SIGNAL S1174 : STD_LOGIC;
    SIGNAL S1175 : STD_LOGIC;
    SIGNAL S1176 : STD_LOGIC;
    SIGNAL S1177 : STD_LOGIC;
    SIGNAL S1178 : STD_LOGIC;
    SIGNAL S1179 : STD_LOGIC;
    SIGNAL S1180 : STD_LOGIC;
    SIGNAL S1181 : STD_LOGIC;
    SIGNAL S1182 : STD_LOGIC;
    SIGNAL S1183 : STD_LOGIC;
    SIGNAL S1184 : STD_LOGIC;
    SIGNAL S1185 : STD_LOGIC;
    SIGNAL S1186 : STD_LOGIC;
    SIGNAL S1187 : STD_LOGIC;
    SIGNAL S1188 : STD_LOGIC;
    SIGNAL S1189 : STD_LOGIC;
    SIGNAL S1190 : STD_LOGIC;
    SIGNAL S1191 : STD_LOGIC;
    SIGNAL S1192 : STD_LOGIC;
    SIGNAL S1193 : STD_LOGIC;
    SIGNAL S1194 : STD_LOGIC;
    SIGNAL S1195 : STD_LOGIC;
    SIGNAL S1196 : STD_LOGIC;
    SIGNAL S1197 : STD_LOGIC;
    SIGNAL S1198 : STD_LOGIC;
    SIGNAL S1199 : STD_LOGIC;
    SIGNAL S1200 : STD_LOGIC;
    SIGNAL S1201 : STD_LOGIC;
    SIGNAL S1202 : STD_LOGIC;
    SIGNAL S1203 : STD_LOGIC;
    SIGNAL S1204 : STD_LOGIC;
    SIGNAL S1205 : STD_LOGIC;
    SIGNAL S1206 : STD_LOGIC;
    SIGNAL S1207 : STD_LOGIC;
    SIGNAL S1208 : STD_LOGIC;
    SIGNAL S1209 : STD_LOGIC;
    SIGNAL S1210 : STD_LOGIC;
    SIGNAL S1211 : STD_LOGIC;
    SIGNAL S1212 : STD_LOGIC;
    SIGNAL S1213 : STD_LOGIC;
    SIGNAL S1214 : STD_LOGIC;
    SIGNAL S1215 : STD_LOGIC;
    SIGNAL S1216 : STD_LOGIC;
    SIGNAL S1217 : STD_LOGIC;
    SIGNAL S1218 : STD_LOGIC;
    SIGNAL S1219 : STD_LOGIC;
    SIGNAL S1220 : STD_LOGIC;
    SIGNAL S1221 : STD_LOGIC;
    SIGNAL S1222 : STD_LOGIC;
    SIGNAL S1223 : STD_LOGIC;
    SIGNAL S1224 : STD_LOGIC;
    SIGNAL S1225 : STD_LOGIC;
    SIGNAL S1226 : STD_LOGIC;
    SIGNAL S1227 : STD_LOGIC;
    SIGNAL S1228 : STD_LOGIC;
    SIGNAL S1229 : STD_LOGIC;
    SIGNAL S1230 : STD_LOGIC;
    SIGNAL S1231 : STD_LOGIC;
    SIGNAL S1232 : STD_LOGIC;
    SIGNAL S1233 : STD_LOGIC;
    SIGNAL S1234 : STD_LOGIC;
    SIGNAL S1235 : STD_LOGIC;
    SIGNAL S1236 : STD_LOGIC;
    SIGNAL S1237 : STD_LOGIC;
    SIGNAL S1238 : STD_LOGIC;
    SIGNAL S1239 : STD_LOGIC;
    SIGNAL S1240 : STD_LOGIC;
    SIGNAL S1241 : STD_LOGIC;
    SIGNAL S1242 : STD_LOGIC;
    SIGNAL S1243 : STD_LOGIC;
    SIGNAL S1244 : STD_LOGIC;
    SIGNAL S1245 : STD_LOGIC;
    SIGNAL S1246 : STD_LOGIC;
    SIGNAL S1247 : STD_LOGIC;
    SIGNAL S1248 : STD_LOGIC;
    SIGNAL S1249 : STD_LOGIC;
    SIGNAL S1250 : STD_LOGIC;
    SIGNAL S1251 : STD_LOGIC;
    SIGNAL S1252 : STD_LOGIC;
    SIGNAL S1253 : STD_LOGIC;
    SIGNAL S1254 : STD_LOGIC;
    SIGNAL S1255 : STD_LOGIC;
    SIGNAL S1256 : STD_LOGIC;
    SIGNAL S1257 : STD_LOGIC;
    SIGNAL S1258 : STD_LOGIC;
    SIGNAL S1259 : STD_LOGIC;
    SIGNAL S1260 : STD_LOGIC;
    SIGNAL S1261 : STD_LOGIC;
    SIGNAL S1262 : STD_LOGIC;
    SIGNAL S1263 : STD_LOGIC;
    SIGNAL S1264 : STD_LOGIC;
    SIGNAL S1265 : STD_LOGIC;
    SIGNAL S1266 : STD_LOGIC;
    SIGNAL S1267 : STD_LOGIC;
    SIGNAL S1268 : STD_LOGIC;
    SIGNAL S1269 : STD_LOGIC;
    SIGNAL S1270 : STD_LOGIC;
    SIGNAL S1271 : STD_LOGIC;
    SIGNAL S1272 : STD_LOGIC;
    SIGNAL S1273 : STD_LOGIC;
    SIGNAL S1274 : STD_LOGIC;
    SIGNAL S1275 : STD_LOGIC;
    SIGNAL S1276 : STD_LOGIC;
    SIGNAL S1277 : STD_LOGIC;
    SIGNAL S1278 : STD_LOGIC;
    SIGNAL S1279 : STD_LOGIC;
    SIGNAL S1280 : STD_LOGIC;
    SIGNAL S1281 : STD_LOGIC;
    SIGNAL S1282 : STD_LOGIC;
    SIGNAL S1283 : STD_LOGIC;
    SIGNAL S1284 : STD_LOGIC;
    SIGNAL S1285 : STD_LOGIC;
    SIGNAL S1286 : STD_LOGIC;
    SIGNAL S1287 : STD_LOGIC;
    SIGNAL S1288 : STD_LOGIC;
    SIGNAL S1289 : STD_LOGIC;
    SIGNAL S1290 : STD_LOGIC;
    SIGNAL S1291 : STD_LOGIC;
    SIGNAL S1292 : STD_LOGIC;
    SIGNAL S1293 : STD_LOGIC;
    SIGNAL S1294 : STD_LOGIC;
    SIGNAL S1295 : STD_LOGIC;
    SIGNAL S1296 : STD_LOGIC;
    SIGNAL S1297 : STD_LOGIC;
    SIGNAL S1298 : STD_LOGIC;
    SIGNAL S1299 : STD_LOGIC;
    SIGNAL S1300 : STD_LOGIC;
    SIGNAL S1301 : STD_LOGIC;
    SIGNAL S1302 : STD_LOGIC;
    SIGNAL S1303 : STD_LOGIC;
    SIGNAL S1304 : STD_LOGIC;
    SIGNAL S1305 : STD_LOGIC;
    SIGNAL S1306 : STD_LOGIC;
    SIGNAL S1307 : STD_LOGIC;
    SIGNAL S1308 : STD_LOGIC;
    SIGNAL S1309 : STD_LOGIC;
    SIGNAL S1310 : STD_LOGIC;
    SIGNAL S1311 : STD_LOGIC;
    SIGNAL S1312 : STD_LOGIC;
    SIGNAL S1313 : STD_LOGIC;
    SIGNAL S1314 : STD_LOGIC;
    SIGNAL S1315 : STD_LOGIC;
    SIGNAL S1316 : STD_LOGIC;
    SIGNAL S1317 : STD_LOGIC;
    SIGNAL S1318 : STD_LOGIC;
    SIGNAL S1319 : STD_LOGIC;
    SIGNAL S1320 : STD_LOGIC;
    SIGNAL S1321 : STD_LOGIC;
    SIGNAL S1322 : STD_LOGIC;
    SIGNAL S1323 : STD_LOGIC;
    SIGNAL S1324 : STD_LOGIC;
    SIGNAL S1325 : STD_LOGIC;
    SIGNAL S1326 : STD_LOGIC;
    SIGNAL S1327 : STD_LOGIC;
    SIGNAL S1328 : STD_LOGIC;
    SIGNAL S1329 : STD_LOGIC;
    SIGNAL S1330 : STD_LOGIC;
    SIGNAL S1331 : STD_LOGIC;
    SIGNAL S1332 : STD_LOGIC;
    SIGNAL S1333 : STD_LOGIC;
    SIGNAL S1334 : STD_LOGIC;
    SIGNAL S1335 : STD_LOGIC;
    SIGNAL S1336 : STD_LOGIC;
    SIGNAL S1337 : STD_LOGIC;
    SIGNAL S1338 : STD_LOGIC;
    SIGNAL S1339 : STD_LOGIC;
    SIGNAL S1340 : STD_LOGIC;
    SIGNAL S1341 : STD_LOGIC;
    SIGNAL S1342 : STD_LOGIC;
    SIGNAL S1343 : STD_LOGIC;
    SIGNAL S1344 : STD_LOGIC;
    SIGNAL S1345 : STD_LOGIC;
    SIGNAL S1346 : STD_LOGIC;
    SIGNAL S1347 : STD_LOGIC;
    SIGNAL S1348 : STD_LOGIC;
    SIGNAL S1349 : STD_LOGIC;
    SIGNAL S1350 : STD_LOGIC;
    SIGNAL S1351 : STD_LOGIC;
    SIGNAL S1352 : STD_LOGIC;
    SIGNAL S1353 : STD_LOGIC;
    SIGNAL S1354 : STD_LOGIC;
    SIGNAL S1355 : STD_LOGIC;
    SIGNAL S1356 : STD_LOGIC;
    SIGNAL S1357 : STD_LOGIC;
    SIGNAL S1358 : STD_LOGIC;
    SIGNAL S1359 : STD_LOGIC;
    SIGNAL S1360 : STD_LOGIC;
    SIGNAL S1361 : STD_LOGIC;
    SIGNAL S1362 : STD_LOGIC;
    SIGNAL S1363 : STD_LOGIC;
    SIGNAL S1364 : STD_LOGIC;
    SIGNAL S1365 : STD_LOGIC;
    SIGNAL S1366 : STD_LOGIC;
    SIGNAL S1367 : STD_LOGIC;
    SIGNAL S1368 : STD_LOGIC;
    SIGNAL S1369 : STD_LOGIC;
    SIGNAL S1370 : STD_LOGIC;
    SIGNAL S1371 : STD_LOGIC;
    SIGNAL S1372 : STD_LOGIC;
    SIGNAL S1373 : STD_LOGIC;
    SIGNAL S1374 : STD_LOGIC;
    SIGNAL S1375 : STD_LOGIC;
    SIGNAL S1376 : STD_LOGIC;
    SIGNAL S1377 : STD_LOGIC;
    SIGNAL S1378 : STD_LOGIC;
    SIGNAL S1379 : STD_LOGIC;
    SIGNAL S1380 : STD_LOGIC;
    SIGNAL S1381 : STD_LOGIC;
    SIGNAL S1382 : STD_LOGIC;
    SIGNAL S1383 : STD_LOGIC;
    SIGNAL S1384 : STD_LOGIC;
    SIGNAL S1385 : STD_LOGIC;
    SIGNAL S1386 : STD_LOGIC;
    SIGNAL S1387 : STD_LOGIC;
    SIGNAL S1388 : STD_LOGIC;
    SIGNAL S1389 : STD_LOGIC;
    SIGNAL S1390 : STD_LOGIC;
    SIGNAL S1391 : STD_LOGIC;
    SIGNAL S1392 : STD_LOGIC;
    SIGNAL S1393 : STD_LOGIC;
    SIGNAL S1394 : STD_LOGIC;
    SIGNAL S1395 : STD_LOGIC;
    SIGNAL S1396 : STD_LOGIC;
    SIGNAL S1397 : STD_LOGIC;
    SIGNAL S1398 : STD_LOGIC;
    SIGNAL S1399 : STD_LOGIC;
    SIGNAL S1400 : STD_LOGIC;
    SIGNAL S1401 : STD_LOGIC;
    SIGNAL S1402 : STD_LOGIC;
    SIGNAL S1403 : STD_LOGIC;
    SIGNAL S1404 : STD_LOGIC;
    SIGNAL S1405 : STD_LOGIC;
    SIGNAL S1406 : STD_LOGIC;
    SIGNAL S1407 : STD_LOGIC;
    SIGNAL S1408 : STD_LOGIC;
    SIGNAL S1409 : STD_LOGIC;
    SIGNAL S1410 : STD_LOGIC;
    SIGNAL S1411 : STD_LOGIC;
    SIGNAL S1412 : STD_LOGIC;
    SIGNAL S1413 : STD_LOGIC;
    SIGNAL S1414 : STD_LOGIC;
    SIGNAL S1415 : STD_LOGIC;
    SIGNAL S1416 : STD_LOGIC;
    SIGNAL S1417 : STD_LOGIC;
    SIGNAL S1418 : STD_LOGIC;
    SIGNAL S1419 : STD_LOGIC;
    SIGNAL S1420 : STD_LOGIC;
    SIGNAL S1421 : STD_LOGIC;
    SIGNAL S1422 : STD_LOGIC;
    SIGNAL S1423 : STD_LOGIC;
    SIGNAL S1424 : STD_LOGIC;
    SIGNAL S1425 : STD_LOGIC;
    SIGNAL S1426 : STD_LOGIC;
    SIGNAL S1427 : STD_LOGIC;
    SIGNAL S1428 : STD_LOGIC;
    SIGNAL S1429 : STD_LOGIC;
    SIGNAL S1430 : STD_LOGIC;
    SIGNAL S1431 : STD_LOGIC;
    SIGNAL S1432 : STD_LOGIC;
    SIGNAL S1433 : STD_LOGIC;
    SIGNAL S1434 : STD_LOGIC;
    SIGNAL S1435 : STD_LOGIC;
    SIGNAL S1436 : STD_LOGIC;
    SIGNAL S1437 : STD_LOGIC;
    SIGNAL S1438 : STD_LOGIC;
    SIGNAL S1439 : STD_LOGIC;
    SIGNAL S1440 : STD_LOGIC;
    SIGNAL S1441 : STD_LOGIC;
    SIGNAL S1442 : STD_LOGIC;
    SIGNAL S1443 : STD_LOGIC;
    SIGNAL S1444 : STD_LOGIC;
    SIGNAL S1445 : STD_LOGIC;
    SIGNAL S1446 : STD_LOGIC;
    SIGNAL S1447 : STD_LOGIC;
    SIGNAL S1448 : STD_LOGIC;
    SIGNAL S1449 : STD_LOGIC;
    SIGNAL S1450 : STD_LOGIC;
    SIGNAL S1451 : STD_LOGIC;
    SIGNAL S1452 : STD_LOGIC;
    SIGNAL S1453 : STD_LOGIC;
    SIGNAL S1454 : STD_LOGIC;
    SIGNAL S1455 : STD_LOGIC;
    SIGNAL S1456 : STD_LOGIC;
    SIGNAL S1457 : STD_LOGIC;
    SIGNAL S1458 : STD_LOGIC;
    SIGNAL S1459 : STD_LOGIC;
    SIGNAL S1460 : STD_LOGIC;
    SIGNAL S1461 : STD_LOGIC;
    SIGNAL S1462 : STD_LOGIC;
    SIGNAL S1463 : STD_LOGIC;
    SIGNAL S1464 : STD_LOGIC;
    SIGNAL S1465 : STD_LOGIC;
    SIGNAL S1466 : STD_LOGIC;
    SIGNAL S1467 : STD_LOGIC;
    SIGNAL S1468 : STD_LOGIC;
    SIGNAL S1469 : STD_LOGIC;
    SIGNAL S1470 : STD_LOGIC;
    SIGNAL S1471 : STD_LOGIC;
    SIGNAL S1472 : STD_LOGIC;
    SIGNAL S1473 : STD_LOGIC;
    SIGNAL S1474 : STD_LOGIC;
    SIGNAL S1475 : STD_LOGIC;
    SIGNAL S1476 : STD_LOGIC;
    SIGNAL S1477 : STD_LOGIC;
    SIGNAL S1478 : STD_LOGIC;
    SIGNAL S1479 : STD_LOGIC;
    SIGNAL S1480 : STD_LOGIC;
    SIGNAL S1481 : STD_LOGIC;
    SIGNAL S1482 : STD_LOGIC;
    SIGNAL S1483 : STD_LOGIC;
    SIGNAL S1484 : STD_LOGIC;
    SIGNAL S1485 : STD_LOGIC;
    SIGNAL S1486 : STD_LOGIC;
    SIGNAL S1487 : STD_LOGIC;
    SIGNAL S1488 : STD_LOGIC;
    SIGNAL S1489 : STD_LOGIC;
    SIGNAL S1490 : STD_LOGIC;
    SIGNAL S1491 : STD_LOGIC;
    SIGNAL S1492 : STD_LOGIC;
    SIGNAL S1493 : STD_LOGIC;
    SIGNAL S1494 : STD_LOGIC;
    SIGNAL S1495 : STD_LOGIC;
    SIGNAL S1496 : STD_LOGIC;
    SIGNAL S1497 : STD_LOGIC;
    SIGNAL S1498 : STD_LOGIC;
    SIGNAL S1499 : STD_LOGIC;
    SIGNAL S1500 : STD_LOGIC;
    SIGNAL S1501 : STD_LOGIC;
    SIGNAL S1502 : STD_LOGIC;
    SIGNAL S1503 : STD_LOGIC;
    SIGNAL S1504 : STD_LOGIC;
    SIGNAL S1505 : STD_LOGIC;
    SIGNAL S1506 : STD_LOGIC;
    SIGNAL S1507 : STD_LOGIC;
    SIGNAL S1508 : STD_LOGIC;
    SIGNAL S1509 : STD_LOGIC;
    SIGNAL S1510 : STD_LOGIC;
    SIGNAL S1511 : STD_LOGIC;
    SIGNAL S1512 : STD_LOGIC;
    SIGNAL S1513 : STD_LOGIC;
    SIGNAL S1514 : STD_LOGIC;
    SIGNAL S1515 : STD_LOGIC;
    SIGNAL S1516 : STD_LOGIC;
    SIGNAL S1517 : STD_LOGIC;
    SIGNAL S1518 : STD_LOGIC;
    SIGNAL S1519 : STD_LOGIC;
    SIGNAL S1520 : STD_LOGIC;
    SIGNAL S1521 : STD_LOGIC;
    SIGNAL S1522 : STD_LOGIC;
    SIGNAL S1523 : STD_LOGIC;
    SIGNAL S1524 : STD_LOGIC;
    SIGNAL S1525 : STD_LOGIC;
    SIGNAL S1526 : STD_LOGIC;
    SIGNAL S1527 : STD_LOGIC;
    SIGNAL S1528 : STD_LOGIC;
    SIGNAL S1529 : STD_LOGIC;
    SIGNAL S1530 : STD_LOGIC;
    SIGNAL S1531 : STD_LOGIC;
    SIGNAL S1532 : STD_LOGIC;
    SIGNAL S1533 : STD_LOGIC;
    SIGNAL S1534 : STD_LOGIC;
    SIGNAL S1535 : STD_LOGIC;
    SIGNAL S1536 : STD_LOGIC;
    SIGNAL S1537 : STD_LOGIC;
    SIGNAL S1538 : STD_LOGIC;
    SIGNAL S1539 : STD_LOGIC;
    SIGNAL S1540 : STD_LOGIC;
    SIGNAL S1541 : STD_LOGIC;
    SIGNAL S1542 : STD_LOGIC;
    SIGNAL S1543 : STD_LOGIC;
    SIGNAL S1544 : STD_LOGIC;
    SIGNAL S1545 : STD_LOGIC;
    SIGNAL S1546 : STD_LOGIC;
    SIGNAL S1547 : STD_LOGIC;
    SIGNAL S1548 : STD_LOGIC;
    SIGNAL S1549 : STD_LOGIC;
    SIGNAL S1550 : STD_LOGIC;
    SIGNAL S1551 : STD_LOGIC;
    SIGNAL S1552 : STD_LOGIC;
    SIGNAL S1553 : STD_LOGIC;
    SIGNAL S1554 : STD_LOGIC;
    SIGNAL S1555 : STD_LOGIC;
    SIGNAL S1556 : STD_LOGIC;
    SIGNAL S1557 : STD_LOGIC;
    SIGNAL S1558 : STD_LOGIC;
    SIGNAL S1559 : STD_LOGIC;
    SIGNAL S1560 : STD_LOGIC;
    SIGNAL S1561 : STD_LOGIC;
    SIGNAL S1562 : STD_LOGIC;
    SIGNAL S1563 : STD_LOGIC;
    SIGNAL S1564 : STD_LOGIC;
    SIGNAL S1565 : STD_LOGIC;
    SIGNAL S1566 : STD_LOGIC;
    SIGNAL S1567 : STD_LOGIC;
    SIGNAL S1568 : STD_LOGIC;
    SIGNAL S1569 : STD_LOGIC;
    SIGNAL S1570 : STD_LOGIC;
    SIGNAL S1571 : STD_LOGIC;
    SIGNAL S1572 : STD_LOGIC;
    SIGNAL S1573 : STD_LOGIC;
    SIGNAL S1574 : STD_LOGIC;
    SIGNAL S1575 : STD_LOGIC;
    SIGNAL S1576 : STD_LOGIC;
    SIGNAL S1577 : STD_LOGIC;
    SIGNAL S1578 : STD_LOGIC;
    SIGNAL S1579 : STD_LOGIC;
    SIGNAL S1580 : STD_LOGIC;
    SIGNAL S1581 : STD_LOGIC;
    SIGNAL S1582 : STD_LOGIC;
    SIGNAL S1583 : STD_LOGIC;
    SIGNAL S1584 : STD_LOGIC;
    SIGNAL S1585 : STD_LOGIC;
    SIGNAL S1586 : STD_LOGIC;
    SIGNAL S1587 : STD_LOGIC;
    SIGNAL S1588 : STD_LOGIC;
    SIGNAL S1589 : STD_LOGIC;
    SIGNAL S1590 : STD_LOGIC;
    SIGNAL S1591 : STD_LOGIC;
    SIGNAL S1592 : STD_LOGIC;
    SIGNAL S1593 : STD_LOGIC;
    SIGNAL S1594 : STD_LOGIC;
    SIGNAL S1595 : STD_LOGIC;
    SIGNAL S1596 : STD_LOGIC;
    SIGNAL S1597 : STD_LOGIC;
    SIGNAL S1598 : STD_LOGIC;
    SIGNAL S1599 : STD_LOGIC;
    SIGNAL S1600 : STD_LOGIC;
    SIGNAL S1601 : STD_LOGIC;
    SIGNAL S1602 : STD_LOGIC;
    SIGNAL S1603 : STD_LOGIC;
    SIGNAL S1604 : STD_LOGIC;
    SIGNAL S1605 : STD_LOGIC;
    SIGNAL S1606 : STD_LOGIC;
    SIGNAL S1607 : STD_LOGIC;
    SIGNAL S1608 : STD_LOGIC;
    SIGNAL S1609 : STD_LOGIC;
    SIGNAL S1610 : STD_LOGIC;
    SIGNAL S1611 : STD_LOGIC;
    SIGNAL S1612 : STD_LOGIC;
    SIGNAL S1613 : STD_LOGIC;
    SIGNAL S1614 : STD_LOGIC;
    SIGNAL S1615 : STD_LOGIC;
    SIGNAL S1616 : STD_LOGIC;
    SIGNAL S1617 : STD_LOGIC;
    SIGNAL S1618 : STD_LOGIC;
    SIGNAL S1619 : STD_LOGIC;
    SIGNAL S1620 : STD_LOGIC;
    SIGNAL S1621 : STD_LOGIC;
    SIGNAL S1622 : STD_LOGIC;
    SIGNAL S1623 : STD_LOGIC;
    SIGNAL S1624 : STD_LOGIC;
    SIGNAL S1625 : STD_LOGIC;
    SIGNAL S1626 : STD_LOGIC;
    SIGNAL S1627 : STD_LOGIC;
    SIGNAL S1628 : STD_LOGIC;
    SIGNAL S1629 : STD_LOGIC;
    SIGNAL S1630 : STD_LOGIC;
    SIGNAL S1631 : STD_LOGIC;
    SIGNAL S1632 : STD_LOGIC;
    SIGNAL S1633 : STD_LOGIC;
    SIGNAL S1634 : STD_LOGIC;
    SIGNAL S1635 : STD_LOGIC;
    SIGNAL S1636 : STD_LOGIC;
    SIGNAL S1637 : STD_LOGIC;
    SIGNAL S1638 : STD_LOGIC;
    SIGNAL S1639 : STD_LOGIC;
    SIGNAL S1640 : STD_LOGIC;
    SIGNAL S1641 : STD_LOGIC;
    SIGNAL S1642 : STD_LOGIC;
    SIGNAL S1643 : STD_LOGIC;
    SIGNAL S1644 : STD_LOGIC;
    SIGNAL S1645 : STD_LOGIC;
    SIGNAL S1646 : STD_LOGIC;
    SIGNAL S1647 : STD_LOGIC;
    SIGNAL S1648 : STD_LOGIC;
    SIGNAL S1649 : STD_LOGIC;
    SIGNAL S1650 : STD_LOGIC;
    SIGNAL S1651 : STD_LOGIC;
    SIGNAL S1652 : STD_LOGIC;
    SIGNAL S1653 : STD_LOGIC;
    SIGNAL S1654 : STD_LOGIC;
    SIGNAL S1655 : STD_LOGIC;
    SIGNAL S1656 : STD_LOGIC;
    SIGNAL S1657 : STD_LOGIC;
    SIGNAL S1658 : STD_LOGIC;
    SIGNAL S1659 : STD_LOGIC;
    SIGNAL S1660 : STD_LOGIC;
    SIGNAL S1661 : STD_LOGIC;
    SIGNAL S1662 : STD_LOGIC;
    SIGNAL S1663 : STD_LOGIC;
    SIGNAL S1664 : STD_LOGIC;
    SIGNAL S1665 : STD_LOGIC;
    SIGNAL S1666 : STD_LOGIC;
    SIGNAL S1667 : STD_LOGIC;
    SIGNAL S1668 : STD_LOGIC;
    SIGNAL S1669 : STD_LOGIC;
    SIGNAL S1670 : STD_LOGIC;
    SIGNAL S1671 : STD_LOGIC;
    SIGNAL S1672 : STD_LOGIC;
    SIGNAL S1673 : STD_LOGIC;
    SIGNAL S1674 : STD_LOGIC;
    SIGNAL S1675 : STD_LOGIC;
    SIGNAL S1676 : STD_LOGIC;
    SIGNAL S1677 : STD_LOGIC;
    SIGNAL S1678 : STD_LOGIC;
    SIGNAL S1679 : STD_LOGIC;
    SIGNAL S1680 : STD_LOGIC;
    SIGNAL S1681 : STD_LOGIC;
    SIGNAL S1682 : STD_LOGIC;
    SIGNAL S1683 : STD_LOGIC;
    SIGNAL S1684 : STD_LOGIC;
    SIGNAL S1685 : STD_LOGIC;
    SIGNAL S1686 : STD_LOGIC;
    SIGNAL S1687 : STD_LOGIC;
    SIGNAL S1688 : STD_LOGIC;
    SIGNAL S1689 : STD_LOGIC;
    SIGNAL S1690 : STD_LOGIC;
    SIGNAL S1691 : STD_LOGIC;
    SIGNAL S1692 : STD_LOGIC;
    SIGNAL S1693 : STD_LOGIC;
    SIGNAL S1694 : STD_LOGIC;
    SIGNAL S1695 : STD_LOGIC;
    SIGNAL S1696 : STD_LOGIC;
    SIGNAL S1697 : STD_LOGIC;
    SIGNAL S1698 : STD_LOGIC;
    SIGNAL S1699 : STD_LOGIC;
    SIGNAL S1700 : STD_LOGIC;
    SIGNAL S1701 : STD_LOGIC;
    SIGNAL S1702 : STD_LOGIC;
    SIGNAL S1703 : STD_LOGIC;
    SIGNAL S1704 : STD_LOGIC;
    SIGNAL S1705 : STD_LOGIC;
    SIGNAL S1706 : STD_LOGIC;
    SIGNAL S1707 : STD_LOGIC;
    SIGNAL S1708 : STD_LOGIC;
    SIGNAL S1709 : STD_LOGIC;
    SIGNAL S1710 : STD_LOGIC;
    SIGNAL S1711 : STD_LOGIC;
    SIGNAL S1712 : STD_LOGIC;
    SIGNAL S1713 : STD_LOGIC;
    SIGNAL S1714 : STD_LOGIC;
    SIGNAL S1715 : STD_LOGIC;
    SIGNAL S1716 : STD_LOGIC;
    SIGNAL S1717 : STD_LOGIC;
    SIGNAL S1718 : STD_LOGIC;
    SIGNAL S1719 : STD_LOGIC;
    SIGNAL S1720 : STD_LOGIC;
    SIGNAL S1721 : STD_LOGIC;
    SIGNAL S1722 : STD_LOGIC;
    SIGNAL S1723 : STD_LOGIC;
    SIGNAL S1724 : STD_LOGIC;
    SIGNAL S1725 : STD_LOGIC;
    SIGNAL S1726 : STD_LOGIC;
    SIGNAL S1727 : STD_LOGIC;
    SIGNAL S1728 : STD_LOGIC;
    SIGNAL S1729 : STD_LOGIC;
    SIGNAL S1730 : STD_LOGIC;
    SIGNAL S1731 : STD_LOGIC;
    SIGNAL S1732 : STD_LOGIC;
    SIGNAL S1733 : STD_LOGIC;
    SIGNAL S1734 : STD_LOGIC;
    SIGNAL S1735 : STD_LOGIC;
    SIGNAL S1736 : STD_LOGIC;
    SIGNAL S1737 : STD_LOGIC;
    SIGNAL S1738 : STD_LOGIC;
    SIGNAL S1739 : STD_LOGIC;
    SIGNAL S1740 : STD_LOGIC;
    SIGNAL S1741 : STD_LOGIC;
    SIGNAL S1742 : STD_LOGIC;
    SIGNAL S1743 : STD_LOGIC;
    SIGNAL S1744 : STD_LOGIC;
    SIGNAL S1745 : STD_LOGIC;
    SIGNAL S1746 : STD_LOGIC;
    SIGNAL S1747 : STD_LOGIC;
    SIGNAL S1748 : STD_LOGIC;
    SIGNAL S1749 : STD_LOGIC;
    SIGNAL S1750 : STD_LOGIC;
    SIGNAL S1751 : STD_LOGIC;
    SIGNAL S1752 : STD_LOGIC;
    SIGNAL S1753 : STD_LOGIC;
    SIGNAL S1754 : STD_LOGIC;
    SIGNAL S1755 : STD_LOGIC;
    SIGNAL S1756 : STD_LOGIC;
    SIGNAL S1757 : STD_LOGIC;
    SIGNAL S1758 : STD_LOGIC;
    SIGNAL S1759 : STD_LOGIC;
    SIGNAL S1760 : STD_LOGIC;
    SIGNAL S1761 : STD_LOGIC;
    SIGNAL S1762 : STD_LOGIC;
    SIGNAL S1763 : STD_LOGIC;
    SIGNAL S1764 : STD_LOGIC;
    SIGNAL S1765 : STD_LOGIC;
    SIGNAL S1766 : STD_LOGIC;
    SIGNAL S1767 : STD_LOGIC;
    SIGNAL S1768 : STD_LOGIC;
    SIGNAL S1769 : STD_LOGIC;
    SIGNAL S1770 : STD_LOGIC;
    SIGNAL S1771 : STD_LOGIC;
    SIGNAL S1772 : STD_LOGIC;
    SIGNAL S1773 : STD_LOGIC;
    SIGNAL S1774 : STD_LOGIC;
    SIGNAL S1775 : STD_LOGIC;
    SIGNAL S1776 : STD_LOGIC;
    SIGNAL S1777 : STD_LOGIC;
    SIGNAL S1778 : STD_LOGIC;
    SIGNAL S1779 : STD_LOGIC;
    SIGNAL S1780 : STD_LOGIC;
    SIGNAL S1781 : STD_LOGIC;
    SIGNAL S1782 : STD_LOGIC;
    SIGNAL S1783 : STD_LOGIC;
    SIGNAL S1784 : STD_LOGIC;
    SIGNAL S1785 : STD_LOGIC;
    SIGNAL S1786 : STD_LOGIC;
    SIGNAL S1787 : STD_LOGIC;
    SIGNAL S1788 : STD_LOGIC;
    SIGNAL S1789 : STD_LOGIC;
    SIGNAL S1790 : STD_LOGIC;
    SIGNAL S1791 : STD_LOGIC;
    SIGNAL S1792 : STD_LOGIC;
    SIGNAL S1793 : STD_LOGIC;
    SIGNAL S1794 : STD_LOGIC;
    SIGNAL S1795 : STD_LOGIC;
    SIGNAL S1796 : STD_LOGIC;
    SIGNAL S1797 : STD_LOGIC;
    SIGNAL S1798 : STD_LOGIC;
    SIGNAL S1799 : STD_LOGIC;
    SIGNAL S1800 : STD_LOGIC;
    SIGNAL S1801 : STD_LOGIC;
    SIGNAL S1802 : STD_LOGIC;
    SIGNAL S1803 : STD_LOGIC;
    SIGNAL S1804 : STD_LOGIC;
    SIGNAL S1805 : STD_LOGIC;
    SIGNAL S1806 : STD_LOGIC;
    SIGNAL S1807 : STD_LOGIC;
    SIGNAL S1808 : STD_LOGIC;
    SIGNAL S1809 : STD_LOGIC;
    SIGNAL S1810 : STD_LOGIC;
    SIGNAL S1811 : STD_LOGIC;
    SIGNAL S1812 : STD_LOGIC;
    SIGNAL S1813 : STD_LOGIC;
    SIGNAL S1814 : STD_LOGIC;
    SIGNAL S1815 : STD_LOGIC;
    SIGNAL S1816 : STD_LOGIC;
    SIGNAL S1817 : STD_LOGIC;
    SIGNAL S1818 : STD_LOGIC;
    SIGNAL S1819 : STD_LOGIC;
    SIGNAL S1820 : STD_LOGIC;
    SIGNAL S1821 : STD_LOGIC;
    SIGNAL S1822 : STD_LOGIC;
    SIGNAL S1823 : STD_LOGIC;
    SIGNAL S1824 : STD_LOGIC;
    SIGNAL S1825 : STD_LOGIC;
    SIGNAL S1826 : STD_LOGIC;
    SIGNAL S1827 : STD_LOGIC;
    SIGNAL S1828 : STD_LOGIC;
    SIGNAL S1829 : STD_LOGIC;
    SIGNAL S1830 : STD_LOGIC;
    SIGNAL S1831 : STD_LOGIC;
    SIGNAL S1832 : STD_LOGIC;
    SIGNAL S1833 : STD_LOGIC;
    SIGNAL S1834 : STD_LOGIC;
    SIGNAL S1835 : STD_LOGIC;
    SIGNAL S1836 : STD_LOGIC;
    SIGNAL S1837 : STD_LOGIC;
    SIGNAL S1838 : STD_LOGIC;
    SIGNAL S1839 : STD_LOGIC;
    SIGNAL S1840 : STD_LOGIC;
    SIGNAL S1841 : STD_LOGIC;
    SIGNAL S1842 : STD_LOGIC;
    SIGNAL S1843 : STD_LOGIC;
    SIGNAL S1844 : STD_LOGIC;
    SIGNAL S1845 : STD_LOGIC;
    SIGNAL S1846 : STD_LOGIC;
    SIGNAL S1847 : STD_LOGIC;
    SIGNAL S1848 : STD_LOGIC;
    SIGNAL S1849 : STD_LOGIC;
    SIGNAL S1850 : STD_LOGIC;
    SIGNAL S1851 : STD_LOGIC;
    SIGNAL S1852 : STD_LOGIC;
    SIGNAL S1853 : STD_LOGIC;
    SIGNAL S1854 : STD_LOGIC;
    SIGNAL S1855 : STD_LOGIC;
    SIGNAL S1856 : STD_LOGIC;
    SIGNAL S1857 : STD_LOGIC;
    SIGNAL S1858 : STD_LOGIC;
    SIGNAL S1859 : STD_LOGIC;
    SIGNAL S1860 : STD_LOGIC;
    SIGNAL S1861 : STD_LOGIC;
    SIGNAL S1862 : STD_LOGIC;
    SIGNAL S1863 : STD_LOGIC;
    SIGNAL S1864 : STD_LOGIC;
    SIGNAL S1865 : STD_LOGIC;
    SIGNAL S1866 : STD_LOGIC;
    SIGNAL S1867 : STD_LOGIC;
    SIGNAL S1868 : STD_LOGIC;
    SIGNAL S1869 : STD_LOGIC;
    SIGNAL S1870 : STD_LOGIC;
    SIGNAL S1871 : STD_LOGIC;
    SIGNAL S1872 : STD_LOGIC;
    SIGNAL S1873 : STD_LOGIC;
    SIGNAL S1874 : STD_LOGIC;
    SIGNAL S1875 : STD_LOGIC;
    SIGNAL S1876 : STD_LOGIC;
    SIGNAL S1877 : STD_LOGIC;
    SIGNAL S1878 : STD_LOGIC;
    SIGNAL S1879 : STD_LOGIC;
    SIGNAL S1880 : STD_LOGIC;
    SIGNAL S1881 : STD_LOGIC;
    SIGNAL S1882 : STD_LOGIC;
    SIGNAL S1883 : STD_LOGIC;
    SIGNAL S1884 : STD_LOGIC;
    SIGNAL S1885 : STD_LOGIC;
    SIGNAL S1886 : STD_LOGIC;
    SIGNAL S1887 : STD_LOGIC;
    SIGNAL S1888 : STD_LOGIC;
    SIGNAL S1889 : STD_LOGIC;
    SIGNAL S1890 : STD_LOGIC;
    SIGNAL S1891 : STD_LOGIC;
    SIGNAL S1892 : STD_LOGIC;
    SIGNAL S1893 : STD_LOGIC;
    SIGNAL S1894 : STD_LOGIC;
    SIGNAL S1895 : STD_LOGIC;
    SIGNAL S1896 : STD_LOGIC;
    SIGNAL S1897 : STD_LOGIC;
    SIGNAL S1898 : STD_LOGIC;
    SIGNAL S1899 : STD_LOGIC;
    SIGNAL S1900 : STD_LOGIC;
    SIGNAL S1901 : STD_LOGIC;
    SIGNAL S1902 : STD_LOGIC;
    SIGNAL S1903 : STD_LOGIC;
    SIGNAL S1904 : STD_LOGIC;
    SIGNAL S1905 : STD_LOGIC;
    SIGNAL S1906 : STD_LOGIC;
    SIGNAL S1907 : STD_LOGIC;
    SIGNAL S1908 : STD_LOGIC;
    SIGNAL S1909 : STD_LOGIC;
    SIGNAL S1910 : STD_LOGIC;
    SIGNAL S1911 : STD_LOGIC;
    SIGNAL S1912 : STD_LOGIC;
    SIGNAL S1913 : STD_LOGIC;
    SIGNAL S1914 : STD_LOGIC;
    SIGNAL S1915 : STD_LOGIC;
    SIGNAL S1916 : STD_LOGIC;
    SIGNAL S1917 : STD_LOGIC;
    SIGNAL S1918 : STD_LOGIC;
    SIGNAL S1919 : STD_LOGIC;
    SIGNAL S1920 : STD_LOGIC;
    SIGNAL S1921 : STD_LOGIC;
    SIGNAL S1922 : STD_LOGIC;
    SIGNAL S1923 : STD_LOGIC;
    SIGNAL S1924 : STD_LOGIC;
    SIGNAL S1925 : STD_LOGIC;
    SIGNAL S1926 : STD_LOGIC;
    SIGNAL S1927 : STD_LOGIC;
    SIGNAL S1928 : STD_LOGIC;
    SIGNAL S1929 : STD_LOGIC;
    SIGNAL S1930 : STD_LOGIC;
    SIGNAL S1931 : STD_LOGIC;
    SIGNAL S1932 : STD_LOGIC;
    SIGNAL S1933 : STD_LOGIC;
    SIGNAL S1934 : STD_LOGIC;
    SIGNAL S1935 : STD_LOGIC;
    SIGNAL S1936 : STD_LOGIC;
    SIGNAL S1937 : STD_LOGIC;
    SIGNAL S1938 : STD_LOGIC;
    SIGNAL S1939 : STD_LOGIC;
    SIGNAL S1940 : STD_LOGIC;
    SIGNAL S1941 : STD_LOGIC;
    SIGNAL S1942 : STD_LOGIC;
    SIGNAL S1943 : STD_LOGIC;
    SIGNAL S1944 : STD_LOGIC;
    SIGNAL S1945 : STD_LOGIC;
    SIGNAL S1946 : STD_LOGIC;
    SIGNAL S1947 : STD_LOGIC;
    SIGNAL S1948 : STD_LOGIC;
    SIGNAL S1949 : STD_LOGIC;
    SIGNAL S1950 : STD_LOGIC;
    SIGNAL S1951 : STD_LOGIC;
    SIGNAL S1952 : STD_LOGIC;
    SIGNAL S1953 : STD_LOGIC;
    SIGNAL S1954 : STD_LOGIC;
    SIGNAL S1955 : STD_LOGIC;
    SIGNAL S1956 : STD_LOGIC;
    SIGNAL S1957 : STD_LOGIC;
    SIGNAL S1958 : STD_LOGIC;
    SIGNAL S1959 : STD_LOGIC;
    SIGNAL S1960 : STD_LOGIC;
    SIGNAL S1961 : STD_LOGIC;
    SIGNAL S1962 : STD_LOGIC;
    SIGNAL S1963 : STD_LOGIC;
    SIGNAL S1964 : STD_LOGIC;
    SIGNAL S1965 : STD_LOGIC;
    SIGNAL S1966 : STD_LOGIC;
    SIGNAL S1967 : STD_LOGIC;
    SIGNAL S1968 : STD_LOGIC;
    SIGNAL S1969 : STD_LOGIC;
    SIGNAL S1970 : STD_LOGIC;
    SIGNAL S1971 : STD_LOGIC;
    SIGNAL S1972 : STD_LOGIC;
    SIGNAL S1973 : STD_LOGIC;
    SIGNAL S1974 : STD_LOGIC;
    SIGNAL S1975 : STD_LOGIC;
    SIGNAL S1976 : STD_LOGIC;
    SIGNAL S1977 : STD_LOGIC;
    SIGNAL S1978 : STD_LOGIC;
    SIGNAL S1979 : STD_LOGIC;
    SIGNAL S1980 : STD_LOGIC;
    SIGNAL S1981 : STD_LOGIC;
    SIGNAL S1982 : STD_LOGIC;
    SIGNAL S1983 : STD_LOGIC;
    SIGNAL S1984 : STD_LOGIC;
    SIGNAL S1985 : STD_LOGIC;
    SIGNAL S1986 : STD_LOGIC;
    SIGNAL S1987 : STD_LOGIC;
    SIGNAL S1988 : STD_LOGIC;
    SIGNAL S1989 : STD_LOGIC;
    SIGNAL S1990 : STD_LOGIC;
    SIGNAL S1991 : STD_LOGIC;
    SIGNAL S1992 : STD_LOGIC;
    SIGNAL S1993 : STD_LOGIC;
    SIGNAL S1994 : STD_LOGIC;
    SIGNAL S1995 : STD_LOGIC;
    SIGNAL S1996 : STD_LOGIC;
    SIGNAL S1997 : STD_LOGIC;
    SIGNAL S1998 : STD_LOGIC;
    SIGNAL S1999 : STD_LOGIC;
    SIGNAL S2000 : STD_LOGIC;
    SIGNAL S2001 : STD_LOGIC;
    SIGNAL S2002 : STD_LOGIC;
    SIGNAL S2003 : STD_LOGIC;
    SIGNAL S2004 : STD_LOGIC;
    SIGNAL S2005 : STD_LOGIC;
    SIGNAL S2006 : STD_LOGIC;
    SIGNAL S2007 : STD_LOGIC;
    SIGNAL S2008 : STD_LOGIC;
    SIGNAL S2009 : STD_LOGIC;
    SIGNAL S2010 : STD_LOGIC;
    SIGNAL S2011 : STD_LOGIC;
    SIGNAL S2012 : STD_LOGIC;
    SIGNAL S2013 : STD_LOGIC;
    SIGNAL S2014 : STD_LOGIC;
    SIGNAL S2015 : STD_LOGIC;
    SIGNAL S2016 : STD_LOGIC;
    SIGNAL S2017 : STD_LOGIC;
    SIGNAL S2018 : STD_LOGIC;
    SIGNAL S2019 : STD_LOGIC;
    SIGNAL S2020 : STD_LOGIC;
    SIGNAL S2021 : STD_LOGIC;
    SIGNAL S2022 : STD_LOGIC;
    SIGNAL S2023 : STD_LOGIC;
    SIGNAL S2024 : STD_LOGIC;
    SIGNAL S2025 : STD_LOGIC;
    SIGNAL S2026 : STD_LOGIC;
    SIGNAL S2027 : STD_LOGIC;
    SIGNAL S2028 : STD_LOGIC;
    SIGNAL S2029 : STD_LOGIC;
    SIGNAL S2030 : STD_LOGIC;
    SIGNAL S2031 : STD_LOGIC;
    SIGNAL S2032 : STD_LOGIC;
    SIGNAL S2033 : STD_LOGIC;
    SIGNAL S2034 : STD_LOGIC;
    SIGNAL S2035 : STD_LOGIC;
    SIGNAL S2036 : STD_LOGIC;
    SIGNAL S2037 : STD_LOGIC;
    SIGNAL S2038 : STD_LOGIC;
    SIGNAL S2039 : STD_LOGIC;
    SIGNAL S2040 : STD_LOGIC;
    SIGNAL S2041 : STD_LOGIC;
    SIGNAL S2042 : STD_LOGIC;
    SIGNAL S2043 : STD_LOGIC;
    SIGNAL S2044 : STD_LOGIC;
    SIGNAL S2045 : STD_LOGIC;
    SIGNAL S2046 : STD_LOGIC;
    SIGNAL S2047 : STD_LOGIC;
    SIGNAL S2048 : STD_LOGIC;
    SIGNAL S2049 : STD_LOGIC;
    SIGNAL S2050 : STD_LOGIC;
    SIGNAL S2051 : STD_LOGIC;
    SIGNAL S2052 : STD_LOGIC;
    SIGNAL S2053 : STD_LOGIC;
    SIGNAL S2054 : STD_LOGIC;
    SIGNAL S2055 : STD_LOGIC;
    SIGNAL S2056 : STD_LOGIC;
    SIGNAL S2057 : STD_LOGIC;
    SIGNAL S2058 : STD_LOGIC;
    SIGNAL S2059 : STD_LOGIC;
    SIGNAL S2060 : STD_LOGIC;
    SIGNAL S2061 : STD_LOGIC;
    SIGNAL S2062 : STD_LOGIC;
    SIGNAL S2063 : STD_LOGIC;
    SIGNAL S2064 : STD_LOGIC;
    SIGNAL S2065 : STD_LOGIC;
    SIGNAL S2066 : STD_LOGIC;
    SIGNAL S2067 : STD_LOGIC;
    SIGNAL S2068 : STD_LOGIC;
    SIGNAL S2069 : STD_LOGIC;
    SIGNAL S2070 : STD_LOGIC;
    SIGNAL S2071 : STD_LOGIC;
    SIGNAL S2072 : STD_LOGIC;
    SIGNAL S2073 : STD_LOGIC;
    SIGNAL S2074 : STD_LOGIC;
    SIGNAL S2075 : STD_LOGIC;
    SIGNAL S2076 : STD_LOGIC;
    SIGNAL S2077 : STD_LOGIC;
    SIGNAL S2078 : STD_LOGIC;
    SIGNAL S2079 : STD_LOGIC;
    SIGNAL S2080 : STD_LOGIC;
    SIGNAL S2081 : STD_LOGIC;
    SIGNAL S2082 : STD_LOGIC;
    SIGNAL S2083 : STD_LOGIC;
    SIGNAL S2084 : STD_LOGIC;
    SIGNAL S2085 : STD_LOGIC;
    SIGNAL S2086 : STD_LOGIC;
    SIGNAL S2087 : STD_LOGIC;
    SIGNAL S2088 : STD_LOGIC;
    SIGNAL S2089 : STD_LOGIC;
    SIGNAL S2090 : STD_LOGIC;
    SIGNAL S2091 : STD_LOGIC;
    SIGNAL S2092 : STD_LOGIC;
    SIGNAL S2093 : STD_LOGIC;
    SIGNAL S2094 : STD_LOGIC;
    SIGNAL S2095 : STD_LOGIC;
    SIGNAL S2096 : STD_LOGIC;
    SIGNAL S2097 : STD_LOGIC;
    SIGNAL S2098 : STD_LOGIC;
    SIGNAL S2099 : STD_LOGIC;
    SIGNAL S2100 : STD_LOGIC;
    SIGNAL S2101 : STD_LOGIC;
    SIGNAL S2102 : STD_LOGIC;
    SIGNAL S2103 : STD_LOGIC;
    SIGNAL S2104 : STD_LOGIC;
    SIGNAL S2105 : STD_LOGIC;
    SIGNAL S2106 : STD_LOGIC;
    SIGNAL S2107 : STD_LOGIC;
    SIGNAL S2108 : STD_LOGIC;
    SIGNAL S2109 : STD_LOGIC;
    SIGNAL S2110 : STD_LOGIC;
    SIGNAL S2111 : STD_LOGIC;
    SIGNAL S2112 : STD_LOGIC;
    SIGNAL S2113 : STD_LOGIC;
    SIGNAL S2114 : STD_LOGIC;
    SIGNAL S2115 : STD_LOGIC;
    SIGNAL S2116 : STD_LOGIC;
    SIGNAL S2117 : STD_LOGIC;
    SIGNAL S2118 : STD_LOGIC;
    SIGNAL S2119 : STD_LOGIC;
    SIGNAL S2120 : STD_LOGIC;
    SIGNAL S2121 : STD_LOGIC;
    SIGNAL S2122 : STD_LOGIC;
    SIGNAL S2123 : STD_LOGIC;
    SIGNAL S2124 : STD_LOGIC;
    SIGNAL S2125 : STD_LOGIC;
    SIGNAL S2126 : STD_LOGIC;
    SIGNAL S2127 : STD_LOGIC;
    SIGNAL S2128 : STD_LOGIC;
    SIGNAL S2129 : STD_LOGIC;
    SIGNAL S2130 : STD_LOGIC;
    SIGNAL S2131 : STD_LOGIC;
    SIGNAL S2132 : STD_LOGIC;
    SIGNAL S2133 : STD_LOGIC;
    SIGNAL S2134 : STD_LOGIC;
    SIGNAL S2135 : STD_LOGIC;
    SIGNAL S2136 : STD_LOGIC;
    SIGNAL S2137 : STD_LOGIC;
    SIGNAL S2138 : STD_LOGIC;
    SIGNAL S2139 : STD_LOGIC;
    SIGNAL S2140 : STD_LOGIC;
    SIGNAL S2141 : STD_LOGIC;
    SIGNAL S2142 : STD_LOGIC;
    SIGNAL S2143 : STD_LOGIC;
    SIGNAL S2144 : STD_LOGIC;
    SIGNAL S2145 : STD_LOGIC;
    SIGNAL S2146 : STD_LOGIC;
    SIGNAL S2147 : STD_LOGIC;
    SIGNAL S2148 : STD_LOGIC;
    SIGNAL S2149 : STD_LOGIC;
    SIGNAL S2150 : STD_LOGIC;
    SIGNAL S2151 : STD_LOGIC;
    SIGNAL S2152 : STD_LOGIC;
    SIGNAL S2153 : STD_LOGIC;
    SIGNAL S2154 : STD_LOGIC;
    SIGNAL S2155 : STD_LOGIC;
    SIGNAL S2156 : STD_LOGIC;
    SIGNAL S2157 : STD_LOGIC;
    SIGNAL S2158 : STD_LOGIC;
    SIGNAL S2159 : STD_LOGIC;
    SIGNAL S2160 : STD_LOGIC;
    SIGNAL S2161 : STD_LOGIC;
    SIGNAL S2162 : STD_LOGIC;
    SIGNAL S2163 : STD_LOGIC;
    SIGNAL S2164 : STD_LOGIC;
    SIGNAL S2165 : STD_LOGIC;
    SIGNAL S2166 : STD_LOGIC;
    SIGNAL S2167 : STD_LOGIC;
    SIGNAL S2168 : STD_LOGIC;
    SIGNAL S2169 : STD_LOGIC;
    SIGNAL S2170 : STD_LOGIC;
    SIGNAL S2171 : STD_LOGIC;
    SIGNAL S2172 : STD_LOGIC;
    SIGNAL S2173 : STD_LOGIC;
    SIGNAL S2174 : STD_LOGIC;
    SIGNAL S2175 : STD_LOGIC;
    SIGNAL S2176 : STD_LOGIC;
    SIGNAL S2177 : STD_LOGIC;
    SIGNAL S2178 : STD_LOGIC;
    SIGNAL S2179 : STD_LOGIC;
    SIGNAL S2180 : STD_LOGIC;
    SIGNAL S2181 : STD_LOGIC;
    SIGNAL S2182 : STD_LOGIC;
    SIGNAL S2183 : STD_LOGIC;
    SIGNAL S2184 : STD_LOGIC;
    SIGNAL S2185 : STD_LOGIC;
    SIGNAL S2186 : STD_LOGIC;
    SIGNAL S2187 : STD_LOGIC;
    SIGNAL S2188 : STD_LOGIC;
    SIGNAL S2189 : STD_LOGIC;
    SIGNAL S2190 : STD_LOGIC;
    SIGNAL S2191 : STD_LOGIC;
    SIGNAL S2192 : STD_LOGIC;
    SIGNAL S2193 : STD_LOGIC;
    SIGNAL S2194 : STD_LOGIC;
    SIGNAL S2195 : STD_LOGIC;
    SIGNAL S2196 : STD_LOGIC;
    SIGNAL S2197 : STD_LOGIC;
    SIGNAL S2198 : STD_LOGIC;
    SIGNAL S2199 : STD_LOGIC;
    SIGNAL S2200 : STD_LOGIC;
    SIGNAL S2201 : STD_LOGIC;
    SIGNAL S2202 : STD_LOGIC;
    SIGNAL S2203 : STD_LOGIC;
    SIGNAL S2204 : STD_LOGIC;
    SIGNAL S2205 : STD_LOGIC;
    SIGNAL S2206 : STD_LOGIC;
    SIGNAL S2207 : STD_LOGIC;
    SIGNAL S2208 : STD_LOGIC;
    SIGNAL S2209 : STD_LOGIC;
    SIGNAL S2210 : STD_LOGIC;
    SIGNAL S2211 : STD_LOGIC;
    SIGNAL S2212 : STD_LOGIC;
    SIGNAL S2213 : STD_LOGIC;
    SIGNAL S2214 : STD_LOGIC;
    SIGNAL S2215 : STD_LOGIC;
    SIGNAL S2216 : STD_LOGIC;
    SIGNAL S2217 : STD_LOGIC;
    SIGNAL S2218 : STD_LOGIC;
    SIGNAL S2219 : STD_LOGIC;
    SIGNAL S2220 : STD_LOGIC;
    SIGNAL S2221 : STD_LOGIC;
    SIGNAL S2222 : STD_LOGIC;
    SIGNAL S2223 : STD_LOGIC;
    SIGNAL S2224 : STD_LOGIC;
    SIGNAL S2225 : STD_LOGIC;
    SIGNAL S2226 : STD_LOGIC;
    SIGNAL S2227 : STD_LOGIC;
    SIGNAL S2228 : STD_LOGIC;
    SIGNAL S2229 : STD_LOGIC;
    SIGNAL S2230 : STD_LOGIC;
    SIGNAL S2231 : STD_LOGIC;
    SIGNAL S2232 : STD_LOGIC;
    SIGNAL S2233 : STD_LOGIC;
    SIGNAL S2234 : STD_LOGIC;
    SIGNAL S2235 : STD_LOGIC;
    SIGNAL S2236 : STD_LOGIC;
    SIGNAL S2237 : STD_LOGIC;
    SIGNAL S2238 : STD_LOGIC;
    SIGNAL S2239 : STD_LOGIC;
    SIGNAL S2240 : STD_LOGIC;
    SIGNAL S2241 : STD_LOGIC;
    SIGNAL S2242 : STD_LOGIC;
    SIGNAL S2243 : STD_LOGIC;
    SIGNAL S2244 : STD_LOGIC;
    SIGNAL S2245 : STD_LOGIC;
    SIGNAL S2246 : STD_LOGIC;
    SIGNAL S2247 : STD_LOGIC;
    SIGNAL S2248 : STD_LOGIC;
    SIGNAL S2249 : STD_LOGIC;
    SIGNAL S2250 : STD_LOGIC;
    SIGNAL S2251 : STD_LOGIC;
    SIGNAL S2252 : STD_LOGIC;
    SIGNAL S2253 : STD_LOGIC;
    SIGNAL S2254 : STD_LOGIC;
    SIGNAL S2255 : STD_LOGIC;
    SIGNAL S2256 : STD_LOGIC;
    SIGNAL S2257 : STD_LOGIC;
    SIGNAL S2258 : STD_LOGIC;
    SIGNAL S2259 : STD_LOGIC;
    SIGNAL S2260 : STD_LOGIC;
    SIGNAL S2261 : STD_LOGIC;
    SIGNAL S2262 : STD_LOGIC;
    SIGNAL S2263 : STD_LOGIC;
    SIGNAL S2264 : STD_LOGIC;
    SIGNAL S2265 : STD_LOGIC;
    SIGNAL S2266 : STD_LOGIC;
    SIGNAL S2267 : STD_LOGIC;
    SIGNAL S2268 : STD_LOGIC;
    SIGNAL S2269 : STD_LOGIC;
    SIGNAL S2270 : STD_LOGIC;
    SIGNAL S2271 : STD_LOGIC;
    SIGNAL S2272 : STD_LOGIC;
    SIGNAL S2273 : STD_LOGIC;
    SIGNAL S2274 : STD_LOGIC;
    SIGNAL S2275 : STD_LOGIC;
    SIGNAL S2276 : STD_LOGIC;
    SIGNAL S2277 : STD_LOGIC;
    SIGNAL S2278 : STD_LOGIC;
    SIGNAL S2279 : STD_LOGIC;
    SIGNAL S2280 : STD_LOGIC;
    SIGNAL S2281 : STD_LOGIC;
    SIGNAL S2282 : STD_LOGIC;
    SIGNAL S2283 : STD_LOGIC;
    SIGNAL S2284 : STD_LOGIC;
    SIGNAL S2285 : STD_LOGIC;
    SIGNAL S2286 : STD_LOGIC;
    SIGNAL S2287 : STD_LOGIC;
    SIGNAL S2288 : STD_LOGIC;
    SIGNAL S2289 : STD_LOGIC;
    SIGNAL S2290 : STD_LOGIC;
    SIGNAL S2291 : STD_LOGIC;
    SIGNAL S2292 : STD_LOGIC;
    SIGNAL S2293 : STD_LOGIC;
    SIGNAL S2294 : STD_LOGIC;
    SIGNAL S2295 : STD_LOGIC;
    SIGNAL S2296 : STD_LOGIC;
    SIGNAL S2297 : STD_LOGIC;
    SIGNAL S2298 : STD_LOGIC;
    SIGNAL S2299 : STD_LOGIC;
    SIGNAL S2300 : STD_LOGIC;
    SIGNAL S2301 : STD_LOGIC;
    SIGNAL S2302 : STD_LOGIC;
    SIGNAL S2303 : STD_LOGIC;
    SIGNAL S2304 : STD_LOGIC;
    SIGNAL S2305 : STD_LOGIC;
    SIGNAL S2306 : STD_LOGIC;
    SIGNAL S2307 : STD_LOGIC;
    SIGNAL S2308 : STD_LOGIC;
    SIGNAL S2309 : STD_LOGIC;
    SIGNAL S2310 : STD_LOGIC;
    SIGNAL S2311 : STD_LOGIC;
    SIGNAL S2312 : STD_LOGIC;
    SIGNAL S2313 : STD_LOGIC;
    SIGNAL S2314 : STD_LOGIC;
    SIGNAL S2315 : STD_LOGIC;
    SIGNAL S2316 : STD_LOGIC;
    SIGNAL S2317 : STD_LOGIC;
    SIGNAL S2318 : STD_LOGIC;
    SIGNAL S2319 : STD_LOGIC;
    SIGNAL S2320 : STD_LOGIC;
    SIGNAL S2321 : STD_LOGIC;
    SIGNAL S2322 : STD_LOGIC;
    SIGNAL S2323 : STD_LOGIC;
    SIGNAL S2324 : STD_LOGIC;
    SIGNAL S2325 : STD_LOGIC;
    SIGNAL S2326 : STD_LOGIC;
    SIGNAL S2327 : STD_LOGIC;
    SIGNAL S2328 : STD_LOGIC;
    SIGNAL S2329 : STD_LOGIC;
    SIGNAL S2330 : STD_LOGIC;
    SIGNAL S2331 : STD_LOGIC;
    SIGNAL S2332 : STD_LOGIC;
    SIGNAL S2333 : STD_LOGIC;
    SIGNAL S2334 : STD_LOGIC;
    SIGNAL S2335 : STD_LOGIC;
    SIGNAL S2336 : STD_LOGIC;
    SIGNAL S2337 : STD_LOGIC;
    SIGNAL S2338 : STD_LOGIC;
    SIGNAL S2339 : STD_LOGIC;
    SIGNAL S2340 : STD_LOGIC;
    SIGNAL S2341 : STD_LOGIC;
    SIGNAL S2342 : STD_LOGIC;
    SIGNAL S2343 : STD_LOGIC;
    SIGNAL S2344 : STD_LOGIC;
    SIGNAL S2345 : STD_LOGIC;
    SIGNAL S2346 : STD_LOGIC;
    SIGNAL S2347 : STD_LOGIC;
    SIGNAL S2348 : STD_LOGIC;
    SIGNAL S2349 : STD_LOGIC;
    SIGNAL S2350 : STD_LOGIC;
    SIGNAL S2351 : STD_LOGIC;
    SIGNAL S2352 : STD_LOGIC;
    SIGNAL S2353 : STD_LOGIC;
    SIGNAL S2354 : STD_LOGIC;
    SIGNAL S2355 : STD_LOGIC;
    SIGNAL S2356 : STD_LOGIC;
    SIGNAL S2357 : STD_LOGIC;
    SIGNAL S2358 : STD_LOGIC;
    SIGNAL S2359 : STD_LOGIC;
    SIGNAL S2360 : STD_LOGIC;
    SIGNAL S2361 : STD_LOGIC;
    SIGNAL S2362 : STD_LOGIC;
    SIGNAL S2363 : STD_LOGIC;
    SIGNAL S2364 : STD_LOGIC;
    SIGNAL S2365 : STD_LOGIC;
    SIGNAL S2366 : STD_LOGIC;
    SIGNAL S2367 : STD_LOGIC;
    SIGNAL S2368 : STD_LOGIC;
    SIGNAL S2369 : STD_LOGIC;
    SIGNAL S2370 : STD_LOGIC;
    SIGNAL S2371 : STD_LOGIC;
    SIGNAL S2372 : STD_LOGIC;
    SIGNAL S2373 : STD_LOGIC;
    SIGNAL S2374 : STD_LOGIC;
    SIGNAL S2375 : STD_LOGIC;
    SIGNAL S2376 : STD_LOGIC;
    SIGNAL S2377 : STD_LOGIC;
    SIGNAL S2378 : STD_LOGIC;
    SIGNAL S2379 : STD_LOGIC;
    SIGNAL S2380 : STD_LOGIC;
    SIGNAL S2381 : STD_LOGIC;
    SIGNAL S2382 : STD_LOGIC;
    SIGNAL S2383 : STD_LOGIC;
    SIGNAL S2384 : STD_LOGIC;
    SIGNAL S2385 : STD_LOGIC;
    SIGNAL S2386 : STD_LOGIC;
    SIGNAL S2387 : STD_LOGIC;
    SIGNAL S2388 : STD_LOGIC;
    SIGNAL S2389 : STD_LOGIC;
    SIGNAL S2390 : STD_LOGIC;
    SIGNAL S2391 : STD_LOGIC;
    SIGNAL S2392 : STD_LOGIC;
    SIGNAL S2393 : STD_LOGIC;
    SIGNAL S2394 : STD_LOGIC;
    SIGNAL S2395 : STD_LOGIC;
    SIGNAL S2396 : STD_LOGIC;
    SIGNAL S2397 : STD_LOGIC;
    SIGNAL S2398 : STD_LOGIC;
    SIGNAL S2399 : STD_LOGIC;
    SIGNAL S2400 : STD_LOGIC;
    SIGNAL S2401 : STD_LOGIC;
    SIGNAL S2402 : STD_LOGIC;
    SIGNAL S2403 : STD_LOGIC;
    SIGNAL S2404 : STD_LOGIC;
    SIGNAL S2405 : STD_LOGIC;
    SIGNAL S2406 : STD_LOGIC;
    SIGNAL S2407 : STD_LOGIC;
    SIGNAL S2408 : STD_LOGIC;
    SIGNAL S2409 : STD_LOGIC;
    SIGNAL S2410 : STD_LOGIC;
    SIGNAL S2411 : STD_LOGIC;
    SIGNAL S2412 : STD_LOGIC;
    SIGNAL S2413 : STD_LOGIC;
    SIGNAL S2414 : STD_LOGIC;
    SIGNAL S2415 : STD_LOGIC;
    SIGNAL S2416 : STD_LOGIC;
    SIGNAL S2417 : STD_LOGIC;
    SIGNAL S2418 : STD_LOGIC;
    SIGNAL S2419 : STD_LOGIC;
    SIGNAL S2420 : STD_LOGIC;
    SIGNAL S2421 : STD_LOGIC;
    SIGNAL S2422 : STD_LOGIC;
    SIGNAL S2423 : STD_LOGIC;
    SIGNAL S2424 : STD_LOGIC;
    SIGNAL S2425 : STD_LOGIC;
    SIGNAL S2426 : STD_LOGIC;
    SIGNAL S2427 : STD_LOGIC;
    SIGNAL S2428 : STD_LOGIC;
    SIGNAL S2429 : STD_LOGIC;
    SIGNAL S2430 : STD_LOGIC;
    SIGNAL S2431 : STD_LOGIC;
    SIGNAL S2432 : STD_LOGIC;
    SIGNAL S2433 : STD_LOGIC;
    SIGNAL S2434 : STD_LOGIC;
    SIGNAL S2435 : STD_LOGIC;
    SIGNAL S2436 : STD_LOGIC;
    SIGNAL S2437 : STD_LOGIC;
    SIGNAL S2438 : STD_LOGIC;
    SIGNAL S2439 : STD_LOGIC;
    SIGNAL S2440 : STD_LOGIC;
    SIGNAL S2441 : STD_LOGIC;
    SIGNAL S2442 : STD_LOGIC;
    SIGNAL S2443 : STD_LOGIC;
    SIGNAL S2444 : STD_LOGIC;
    SIGNAL S2445 : STD_LOGIC;
    SIGNAL S2446 : STD_LOGIC;
    SIGNAL S2447 : STD_LOGIC;
    SIGNAL S2448 : STD_LOGIC;
    SIGNAL S2449 : STD_LOGIC;
    SIGNAL S2450 : STD_LOGIC;
    SIGNAL S2451 : STD_LOGIC;
    SIGNAL S2452 : STD_LOGIC;
    SIGNAL S2453 : STD_LOGIC;
    SIGNAL S2454 : STD_LOGIC;
    SIGNAL S2455 : STD_LOGIC;
    SIGNAL S2456 : STD_LOGIC;
    SIGNAL S2457 : STD_LOGIC;
    SIGNAL S2458 : STD_LOGIC;
    SIGNAL S2459 : STD_LOGIC;
    SIGNAL S2460 : STD_LOGIC;
    SIGNAL S2461 : STD_LOGIC;
    SIGNAL S2462 : STD_LOGIC;
    SIGNAL S2463 : STD_LOGIC;
    SIGNAL S2464 : STD_LOGIC;
    SIGNAL S2465 : STD_LOGIC;
    SIGNAL S2466 : STD_LOGIC;
    SIGNAL S2467 : STD_LOGIC;
    SIGNAL S2468 : STD_LOGIC;
    SIGNAL S2469 : STD_LOGIC;
    SIGNAL S2470 : STD_LOGIC;
    SIGNAL S2471 : STD_LOGIC;
    SIGNAL S2472 : STD_LOGIC;
    SIGNAL S2473 : STD_LOGIC;
    SIGNAL S2474 : STD_LOGIC;
    SIGNAL S2475 : STD_LOGIC;
    SIGNAL S2476 : STD_LOGIC;
    SIGNAL S2477 : STD_LOGIC;
    SIGNAL S2478 : STD_LOGIC;
    SIGNAL S2479 : STD_LOGIC;
    SIGNAL S2480 : STD_LOGIC;
    SIGNAL S2481 : STD_LOGIC;
    SIGNAL S2482 : STD_LOGIC;
    SIGNAL S2483 : STD_LOGIC;
    SIGNAL S2484 : STD_LOGIC;
    SIGNAL S2485 : STD_LOGIC;
    SIGNAL S2486 : STD_LOGIC;
    SIGNAL S2487 : STD_LOGIC;
    SIGNAL S2488 : STD_LOGIC;
    SIGNAL S2489 : STD_LOGIC;
    SIGNAL S2490 : STD_LOGIC;
    SIGNAL S2491 : STD_LOGIC;
    SIGNAL S2492 : STD_LOGIC;
    SIGNAL S2493 : STD_LOGIC;
    SIGNAL S2494 : STD_LOGIC;
    SIGNAL S2495 : STD_LOGIC;
    SIGNAL S2496 : STD_LOGIC;
    SIGNAL S2497 : STD_LOGIC;
    SIGNAL S2498 : STD_LOGIC;
    SIGNAL S2499 : STD_LOGIC;
    SIGNAL S2500 : STD_LOGIC;
    SIGNAL S2501 : STD_LOGIC;
    SIGNAL S2502 : STD_LOGIC;
    SIGNAL S2503 : STD_LOGIC;
    SIGNAL S2504 : STD_LOGIC;
    SIGNAL S2505 : STD_LOGIC;
    SIGNAL S2506 : STD_LOGIC;
    SIGNAL S2507 : STD_LOGIC;
    SIGNAL S2508 : STD_LOGIC;
    SIGNAL S2509 : STD_LOGIC;
    SIGNAL S2510 : STD_LOGIC;
    SIGNAL S2511 : STD_LOGIC;
    SIGNAL S2512 : STD_LOGIC;
    SIGNAL S2513 : STD_LOGIC;
    SIGNAL S2514 : STD_LOGIC;
    SIGNAL S2515 : STD_LOGIC;
    SIGNAL S2516 : STD_LOGIC;
    SIGNAL S2517 : STD_LOGIC;
    SIGNAL S2518 : STD_LOGIC;
    SIGNAL S2519 : STD_LOGIC;
    SIGNAL S2520 : STD_LOGIC;
    SIGNAL S2521 : STD_LOGIC;
    SIGNAL S2522 : STD_LOGIC;
    SIGNAL S2523 : STD_LOGIC;
    SIGNAL S2524 : STD_LOGIC;
    SIGNAL S2525 : STD_LOGIC;
    SIGNAL S2526 : STD_LOGIC;
    SIGNAL S2527 : STD_LOGIC;
    SIGNAL S2528 : STD_LOGIC;
    SIGNAL S2529 : STD_LOGIC;
    SIGNAL S2530 : STD_LOGIC;
    SIGNAL S2531 : STD_LOGIC;
    SIGNAL S2532 : STD_LOGIC;
    SIGNAL S2533 : STD_LOGIC;
    SIGNAL S2534 : STD_LOGIC;
    SIGNAL S2535 : STD_LOGIC;
    SIGNAL S2536 : STD_LOGIC;
    SIGNAL S2537 : STD_LOGIC;
    SIGNAL S2538 : STD_LOGIC;
    SIGNAL S2539 : STD_LOGIC;
    SIGNAL S2540 : STD_LOGIC;
    SIGNAL S2541 : STD_LOGIC;
    SIGNAL S2542 : STD_LOGIC;
    SIGNAL S2543 : STD_LOGIC;
    SIGNAL S2544 : STD_LOGIC;
    SIGNAL S2545 : STD_LOGIC;
    SIGNAL S2546 : STD_LOGIC;
    SIGNAL S2547 : STD_LOGIC;
    SIGNAL S2548 : STD_LOGIC;
    SIGNAL S2549 : STD_LOGIC;
    SIGNAL S2550 : STD_LOGIC;
    SIGNAL S2551 : STD_LOGIC;
    SIGNAL S2552 : STD_LOGIC;
    SIGNAL S2553 : STD_LOGIC;
    SIGNAL S2554 : STD_LOGIC;
    SIGNAL S2555 : STD_LOGIC;
    SIGNAL S2556 : STD_LOGIC;
    SIGNAL S2557 : STD_LOGIC;
    SIGNAL S2558 : STD_LOGIC;
    SIGNAL S2559 : STD_LOGIC;
    SIGNAL S2560 : STD_LOGIC;
    SIGNAL S2561 : STD_LOGIC;
    SIGNAL S2562 : STD_LOGIC;
    SIGNAL S2563 : STD_LOGIC;
    SIGNAL S2564 : STD_LOGIC;
    SIGNAL S2565 : STD_LOGIC;
    SIGNAL S2566 : STD_LOGIC;
    SIGNAL S2567 : STD_LOGIC;
    SIGNAL S2568 : STD_LOGIC;
    SIGNAL S2569 : STD_LOGIC;
    SIGNAL S2570 : STD_LOGIC;
    SIGNAL S2571 : STD_LOGIC;
    SIGNAL S2572 : STD_LOGIC;
    SIGNAL S2573 : STD_LOGIC;
    SIGNAL S2574 : STD_LOGIC;
    SIGNAL S2575 : STD_LOGIC;
    SIGNAL S2576 : STD_LOGIC;
    SIGNAL S2577 : STD_LOGIC;
    SIGNAL S2578 : STD_LOGIC;
    SIGNAL S2579 : STD_LOGIC;
    SIGNAL S2580 : STD_LOGIC;
    SIGNAL S2581 : STD_LOGIC;
    SIGNAL S2582 : STD_LOGIC;
    SIGNAL S2583 : STD_LOGIC;
    SIGNAL S2584 : STD_LOGIC;
    SIGNAL S2585 : STD_LOGIC;
    SIGNAL S2586 : STD_LOGIC;
    SIGNAL S2587 : STD_LOGIC;
    SIGNAL S2588 : STD_LOGIC;
    SIGNAL S2589 : STD_LOGIC;
    SIGNAL S2590 : STD_LOGIC;
    SIGNAL S2591 : STD_LOGIC;
    SIGNAL S2592 : STD_LOGIC;
    SIGNAL S2593 : STD_LOGIC;
    SIGNAL S2594 : STD_LOGIC;
    SIGNAL S2595 : STD_LOGIC;
    SIGNAL S2596 : STD_LOGIC;
    SIGNAL S2597 : STD_LOGIC;
    SIGNAL S2598 : STD_LOGIC;
    SIGNAL S2599 : STD_LOGIC;
    SIGNAL S2600 : STD_LOGIC;
    SIGNAL S2601 : STD_LOGIC;
    SIGNAL S2602 : STD_LOGIC;
    SIGNAL S2603 : STD_LOGIC;
    SIGNAL S2604 : STD_LOGIC;
    SIGNAL S2605 : STD_LOGIC;
    SIGNAL S2606 : STD_LOGIC;
    SIGNAL S2607 : STD_LOGIC;
    SIGNAL S2608 : STD_LOGIC;
    SIGNAL S2609 : STD_LOGIC;
    SIGNAL S2610 : STD_LOGIC;
    SIGNAL S2611 : STD_LOGIC;
    SIGNAL S2612 : STD_LOGIC;
    SIGNAL S2613 : STD_LOGIC;
    SIGNAL S2614 : STD_LOGIC;
    SIGNAL S2615 : STD_LOGIC;
    SIGNAL S2616 : STD_LOGIC;
    SIGNAL S2617 : STD_LOGIC;
    SIGNAL S2618 : STD_LOGIC;
    SIGNAL S2619 : STD_LOGIC;
    SIGNAL S2620 : STD_LOGIC;
    SIGNAL S2621 : STD_LOGIC;
    SIGNAL S2622 : STD_LOGIC;
    SIGNAL S2623 : STD_LOGIC;
    SIGNAL S2624 : STD_LOGIC;
    SIGNAL S2625 : STD_LOGIC;
    SIGNAL S2626 : STD_LOGIC;
    SIGNAL S2627 : STD_LOGIC;
    SIGNAL S2628 : STD_LOGIC;
    SIGNAL S2629 : STD_LOGIC;
    SIGNAL S2630 : STD_LOGIC;
    SIGNAL S2631 : STD_LOGIC;
    SIGNAL S2632 : STD_LOGIC;
    SIGNAL S2633 : STD_LOGIC;
    SIGNAL S2634 : STD_LOGIC;
    SIGNAL S2635 : STD_LOGIC;
    SIGNAL S2636 : STD_LOGIC;
    SIGNAL S2637 : STD_LOGIC;
    SIGNAL S2638 : STD_LOGIC;
    SIGNAL S2639 : STD_LOGIC;
    SIGNAL S2640 : STD_LOGIC;
    SIGNAL S2641 : STD_LOGIC;
    SIGNAL S2642 : STD_LOGIC;
    SIGNAL S2643 : STD_LOGIC;
    SIGNAL S2644 : STD_LOGIC;
    SIGNAL S2645 : STD_LOGIC;
    SIGNAL S2646 : STD_LOGIC;
    SIGNAL S2647 : STD_LOGIC;
    SIGNAL S2648 : STD_LOGIC;
    SIGNAL S2649 : STD_LOGIC;
    SIGNAL S2650 : STD_LOGIC;
    SIGNAL S2651 : STD_LOGIC;
    SIGNAL S2652 : STD_LOGIC;
    SIGNAL S2653 : STD_LOGIC;
    SIGNAL S2654 : STD_LOGIC;
    SIGNAL S2655 : STD_LOGIC;
    SIGNAL S2656 : STD_LOGIC;
    SIGNAL S2657 : STD_LOGIC;
    SIGNAL S2658 : STD_LOGIC;
    SIGNAL S2659 : STD_LOGIC;
    SIGNAL S2660 : STD_LOGIC;
    SIGNAL S2661 : STD_LOGIC;
    SIGNAL S2662 : STD_LOGIC;
    SIGNAL S2663 : STD_LOGIC;
    SIGNAL S2664 : STD_LOGIC;
    SIGNAL S2665 : STD_LOGIC;
    SIGNAL S2666 : STD_LOGIC;
    SIGNAL S2667 : STD_LOGIC;
    SIGNAL S2668 : STD_LOGIC;
    SIGNAL S2669 : STD_LOGIC;
    SIGNAL S2670 : STD_LOGIC;
    SIGNAL S2671 : STD_LOGIC;
    SIGNAL S2672 : STD_LOGIC;
    SIGNAL S2673 : STD_LOGIC;
    SIGNAL S2674 : STD_LOGIC;
    SIGNAL S2675 : STD_LOGIC;
    SIGNAL S2676 : STD_LOGIC;
    SIGNAL S2677 : STD_LOGIC;
    SIGNAL S2678 : STD_LOGIC;
    SIGNAL S2679 : STD_LOGIC;
    SIGNAL S2680 : STD_LOGIC;
    SIGNAL S2681 : STD_LOGIC;
    SIGNAL S2682 : STD_LOGIC;
    SIGNAL S2683 : STD_LOGIC;
    SIGNAL S2684 : STD_LOGIC;
    SIGNAL S2685 : STD_LOGIC;
    SIGNAL S2686 : STD_LOGIC;
    SIGNAL S2687 : STD_LOGIC;
    SIGNAL S2688 : STD_LOGIC;
    SIGNAL S2689 : STD_LOGIC;
    SIGNAL S2690 : STD_LOGIC;
    SIGNAL S2691 : STD_LOGIC;
    SIGNAL S2692 : STD_LOGIC;
    SIGNAL S2693 : STD_LOGIC;
    SIGNAL S2694 : STD_LOGIC;
    SIGNAL S2695 : STD_LOGIC;
    SIGNAL S2696 : STD_LOGIC;
    SIGNAL S2697 : STD_LOGIC;
    SIGNAL S2698 : STD_LOGIC;
    SIGNAL S2699 : STD_LOGIC;
    SIGNAL S2700 : STD_LOGIC;
    SIGNAL S2701 : STD_LOGIC;
    SIGNAL S2702 : STD_LOGIC;
    SIGNAL S2703 : STD_LOGIC;
    SIGNAL S2704 : STD_LOGIC;
    SIGNAL S2705 : STD_LOGIC;
    SIGNAL S2706 : STD_LOGIC;
    SIGNAL S2707 : STD_LOGIC;
    SIGNAL S2708 : STD_LOGIC;
    SIGNAL S2709 : STD_LOGIC;
    SIGNAL S2710 : STD_LOGIC;
    SIGNAL S2711 : STD_LOGIC;
    SIGNAL S2712 : STD_LOGIC;
    SIGNAL S2713 : STD_LOGIC;
    SIGNAL S2714 : STD_LOGIC;
    SIGNAL S2715 : STD_LOGIC;
    SIGNAL S2716 : STD_LOGIC;
    SIGNAL S2717 : STD_LOGIC;
    SIGNAL S2718 : STD_LOGIC;
    SIGNAL S2719 : STD_LOGIC;
    SIGNAL S2720 : STD_LOGIC;
    SIGNAL S2721 : STD_LOGIC;
    SIGNAL S2722 : STD_LOGIC;
    SIGNAL S2723 : STD_LOGIC;
    SIGNAL S2724 : STD_LOGIC;
    SIGNAL S2725 : STD_LOGIC;
    SIGNAL S2726 : STD_LOGIC;
    SIGNAL S2727 : STD_LOGIC;
    SIGNAL S2728 : STD_LOGIC;
    SIGNAL S2729 : STD_LOGIC;
    SIGNAL S2730 : STD_LOGIC;
    SIGNAL S2731 : STD_LOGIC;
    SIGNAL S2732 : STD_LOGIC;
    SIGNAL S2733 : STD_LOGIC;
    SIGNAL S2734 : STD_LOGIC;
    SIGNAL S2735 : STD_LOGIC;
    SIGNAL S2736 : STD_LOGIC;
    SIGNAL S2737 : STD_LOGIC;
    SIGNAL S2738 : STD_LOGIC;
    SIGNAL S2739 : STD_LOGIC;
    SIGNAL S2740 : STD_LOGIC;
    SIGNAL S2741 : STD_LOGIC;
    SIGNAL S2742 : STD_LOGIC;
    SIGNAL S2743 : STD_LOGIC;
    SIGNAL S2744 : STD_LOGIC;
    SIGNAL S2745 : STD_LOGIC;
    SIGNAL S2746 : STD_LOGIC;
    SIGNAL S2747 : STD_LOGIC;
    SIGNAL S2748 : STD_LOGIC;
    SIGNAL S2749 : STD_LOGIC;
    SIGNAL S2750 : STD_LOGIC;
    SIGNAL S2751 : STD_LOGIC;
    SIGNAL S2752 : STD_LOGIC;
    SIGNAL S2753 : STD_LOGIC;
    SIGNAL S2754 : STD_LOGIC;
    SIGNAL S2755 : STD_LOGIC;
    SIGNAL S2756 : STD_LOGIC;
    SIGNAL S2757 : STD_LOGIC;
    SIGNAL S2758 : STD_LOGIC;
    SIGNAL S2759 : STD_LOGIC;
    SIGNAL S2760 : STD_LOGIC;
    SIGNAL S2761 : STD_LOGIC;
    SIGNAL S2762 : STD_LOGIC;
    SIGNAL S2763 : STD_LOGIC;
    SIGNAL S2764 : STD_LOGIC;
    SIGNAL S2765 : STD_LOGIC;
    SIGNAL S2766 : STD_LOGIC;
    SIGNAL S2767 : STD_LOGIC;
    SIGNAL S2768 : STD_LOGIC;
    SIGNAL S2769 : STD_LOGIC;
    SIGNAL S2770 : STD_LOGIC;
    SIGNAL S2771 : STD_LOGIC;
    SIGNAL S2772 : STD_LOGIC;
    SIGNAL S2773 : STD_LOGIC;
    SIGNAL S2774 : STD_LOGIC;
    SIGNAL S2775 : STD_LOGIC;
    SIGNAL S2776 : STD_LOGIC;
    SIGNAL S2777 : STD_LOGIC;
    SIGNAL S2778 : STD_LOGIC;
    SIGNAL S2779 : STD_LOGIC;
    SIGNAL S2780 : STD_LOGIC;
    SIGNAL S2781 : STD_LOGIC;
    SIGNAL S2782 : STD_LOGIC;
    SIGNAL S2783 : STD_LOGIC;
    SIGNAL S2784 : STD_LOGIC;
    SIGNAL S2785 : STD_LOGIC;
    SIGNAL S2786 : STD_LOGIC;
    SIGNAL S2787 : STD_LOGIC;
    SIGNAL S2788 : STD_LOGIC;
    SIGNAL S2789 : STD_LOGIC;
    SIGNAL S2790 : STD_LOGIC;
    SIGNAL S2791 : STD_LOGIC;
    SIGNAL S2792 : STD_LOGIC;
    SIGNAL S2793 : STD_LOGIC;
    SIGNAL S2794 : STD_LOGIC;
    SIGNAL S2795 : STD_LOGIC;
    SIGNAL S2796 : STD_LOGIC;
    SIGNAL S2797 : STD_LOGIC;
    SIGNAL S2798 : STD_LOGIC;
    SIGNAL S2799 : STD_LOGIC;
    SIGNAL S2800 : STD_LOGIC;
    SIGNAL S2801 : STD_LOGIC;
    SIGNAL S2802 : STD_LOGIC;
    SIGNAL S2803 : STD_LOGIC;
    SIGNAL S2804 : STD_LOGIC;
    SIGNAL S2805 : STD_LOGIC;
    SIGNAL S2806 : STD_LOGIC;
    SIGNAL S2807 : STD_LOGIC;
    SIGNAL S2808 : STD_LOGIC;
    SIGNAL S2809 : STD_LOGIC;
    SIGNAL S2810 : STD_LOGIC;
    SIGNAL S2811 : STD_LOGIC;
    SIGNAL S2812 : STD_LOGIC;
    SIGNAL S2813 : STD_LOGIC;
    SIGNAL S2814 : STD_LOGIC;
    SIGNAL S2815 : STD_LOGIC;
    SIGNAL S2816 : STD_LOGIC;
    SIGNAL S2817 : STD_LOGIC;
    SIGNAL S2818 : STD_LOGIC;
    SIGNAL S2819 : STD_LOGIC;
    SIGNAL S2820 : STD_LOGIC;
    SIGNAL S2821 : STD_LOGIC;
    SIGNAL S2822 : STD_LOGIC;
    SIGNAL S2823 : STD_LOGIC;
    SIGNAL S2824 : STD_LOGIC;
    SIGNAL S2825 : STD_LOGIC;
    SIGNAL S2826 : STD_LOGIC;
    SIGNAL S2827 : STD_LOGIC;
    SIGNAL S2828 : STD_LOGIC;
    SIGNAL S2829 : STD_LOGIC;
    SIGNAL S2830 : STD_LOGIC;
    SIGNAL S2831 : STD_LOGIC;
    SIGNAL S2832 : STD_LOGIC;
    SIGNAL S2833 : STD_LOGIC;
    SIGNAL S2834 : STD_LOGIC;
    SIGNAL S2835 : STD_LOGIC;
    SIGNAL S2836 : STD_LOGIC;
    SIGNAL S2837 : STD_LOGIC;
    SIGNAL S2838 : STD_LOGIC;
    SIGNAL S2839 : STD_LOGIC;
    SIGNAL S2840 : STD_LOGIC;
    SIGNAL S2841 : STD_LOGIC;
    SIGNAL S2842 : STD_LOGIC;
    SIGNAL S2843 : STD_LOGIC;
    SIGNAL S2844 : STD_LOGIC;
    SIGNAL S2845 : STD_LOGIC;
    SIGNAL S2846 : STD_LOGIC;
    SIGNAL S2847 : STD_LOGIC;
    SIGNAL S2848 : STD_LOGIC;
    SIGNAL S2849 : STD_LOGIC;
    SIGNAL S2850 : STD_LOGIC;
    SIGNAL S2851 : STD_LOGIC;
    SIGNAL S2852 : STD_LOGIC;
    SIGNAL S2853 : STD_LOGIC;
    SIGNAL S2854 : STD_LOGIC;
    SIGNAL S2855 : STD_LOGIC;
    SIGNAL S2856 : STD_LOGIC;
    SIGNAL S2857 : STD_LOGIC;
    SIGNAL S2858 : STD_LOGIC;
    SIGNAL S2859 : STD_LOGIC;
    SIGNAL S2860 : STD_LOGIC;
    SIGNAL S2861 : STD_LOGIC;
    SIGNAL S2862 : STD_LOGIC;
    SIGNAL S2863 : STD_LOGIC;
    SIGNAL S2864 : STD_LOGIC;
    SIGNAL S2865 : STD_LOGIC;
    SIGNAL S2866 : STD_LOGIC;
    SIGNAL S2867 : STD_LOGIC;
    SIGNAL S2868 : STD_LOGIC;
    SIGNAL S2869 : STD_LOGIC;
    SIGNAL S2870 : STD_LOGIC;
    SIGNAL S2871 : STD_LOGIC;
    SIGNAL S2872 : STD_LOGIC;
    SIGNAL S2873 : STD_LOGIC;
    SIGNAL S2874 : STD_LOGIC;
    SIGNAL S2875 : STD_LOGIC;
    SIGNAL S2876 : STD_LOGIC;
    SIGNAL S2877 : STD_LOGIC;
    SIGNAL S2878 : STD_LOGIC;
    SIGNAL S2879 : STD_LOGIC;
    SIGNAL S2880 : STD_LOGIC;
    SIGNAL S2881 : STD_LOGIC;
    SIGNAL S2882 : STD_LOGIC;
    SIGNAL S2883 : STD_LOGIC;
    SIGNAL S2884 : STD_LOGIC;
    SIGNAL S2885 : STD_LOGIC;
    SIGNAL S2886 : STD_LOGIC;
    SIGNAL S2887 : STD_LOGIC;
    SIGNAL S2888 : STD_LOGIC;
    SIGNAL S2889 : STD_LOGIC;
    SIGNAL S2890 : STD_LOGIC;
    SIGNAL S2891 : STD_LOGIC;
    SIGNAL S2892 : STD_LOGIC;
    SIGNAL S2893 : STD_LOGIC;
    SIGNAL S2894 : STD_LOGIC;
    SIGNAL S2895 : STD_LOGIC;
    SIGNAL S2896 : STD_LOGIC;
    SIGNAL S2897 : STD_LOGIC;
    SIGNAL S2898 : STD_LOGIC;
    SIGNAL S2899 : STD_LOGIC;
    SIGNAL S2900 : STD_LOGIC;
    SIGNAL S2901 : STD_LOGIC;
    SIGNAL S2902 : STD_LOGIC;
    SIGNAL S2903 : STD_LOGIC;
    SIGNAL S2904 : STD_LOGIC;
    SIGNAL S2905 : STD_LOGIC;
    SIGNAL U1_AC_out_0 : STD_LOGIC;
    SIGNAL U1_AC_out_10 : STD_LOGIC;
    SIGNAL U1_AC_out_11 : STD_LOGIC;
    SIGNAL U1_AC_out_12 : STD_LOGIC;
    SIGNAL U1_AC_out_13 : STD_LOGIC;
    SIGNAL U1_AC_out_14 : STD_LOGIC;
    SIGNAL U1_AC_out_15 : STD_LOGIC;
    SIGNAL U1_AC_out_1 : STD_LOGIC;
    SIGNAL U1_AC_out_2 : STD_LOGIC;
    SIGNAL U1_AC_out_3 : STD_LOGIC;
    SIGNAL U1_AC_out_4 : STD_LOGIC;
    SIGNAL U1_AC_out_5 : STD_LOGIC;
    SIGNAL U1_AC_out_6 : STD_LOGIC;
    SIGNAL U1_AC_out_7 : STD_LOGIC;
    SIGNAL U1_AC_out_8 : STD_LOGIC;
    SIGNAL U1_AC_out_9 : STD_LOGIC;
    SIGNAL U1_ADD : STD_LOGIC;
    SIGNAL U1_AND : STD_LOGIC;
    SIGNAL U1_C : STD_LOGIC;
    SIGNAL U1_C_out1 : STD_LOGIC;
    SIGNAL U1_INC1 : STD_LOGIC;
    SIGNAL U1_INC2 : STD_LOGIC;
    SIGNAL U1_IN_out_0 : STD_LOGIC;
    SIGNAL U1_IN_out_10 : STD_LOGIC;
    SIGNAL U1_IN_out_11 : STD_LOGIC;
    SIGNAL U1_IN_out_12 : STD_LOGIC;
    SIGNAL U1_IN_out_13 : STD_LOGIC;
    SIGNAL U1_IN_out_14 : STD_LOGIC;
    SIGNAL U1_IN_out_15 : STD_LOGIC;
    SIGNAL U1_IN_out_1 : STD_LOGIC;
    SIGNAL U1_IN_out_2 : STD_LOGIC;
    SIGNAL U1_IN_out_3 : STD_LOGIC;
    SIGNAL U1_IN_out_4 : STD_LOGIC;
    SIGNAL U1_IN_out_5 : STD_LOGIC;
    SIGNAL U1_IN_out_6 : STD_LOGIC;
    SIGNAL U1_IN_out_7 : STD_LOGIC;
    SIGNAL U1_IN_out_8 : STD_LOGIC;
    SIGNAL U1_IN_out_9 : STD_LOGIC;
    SIGNAL U1_IR_out_0 : STD_LOGIC;
    SIGNAL U1_IR_out_10 : STD_LOGIC;
    SIGNAL U1_IR_out_11 : STD_LOGIC;
    SIGNAL U1_IR_out_12 : STD_LOGIC;
    SIGNAL U1_IR_out_13 : STD_LOGIC;
    SIGNAL U1_IR_out_14 : STD_LOGIC;
    SIGNAL U1_IR_out_15 : STD_LOGIC;
    SIGNAL U1_IR_out_1 : STD_LOGIC;
    SIGNAL U1_IR_out_2 : STD_LOGIC;
    SIGNAL U1_IR_out_3 : STD_LOGIC;
    SIGNAL U1_IR_out_4 : STD_LOGIC;
    SIGNAL U1_IR_out_5 : STD_LOGIC;
    SIGNAL U1_IR_out_6 : STD_LOGIC;
    SIGNAL U1_IR_out_7 : STD_LOGIC;
    SIGNAL U1_IR_out_8 : STD_LOGIC;
    SIGNAL U1_IR_out_9 : STD_LOGIC;
    SIGNAL U1_LGU_out_15 : STD_LOGIC;
    SIGNAL U1_MUL : STD_LOGIC;
    SIGNAL U1_NOT : STD_LOGIC;
    SIGNAL U1_N_out1 : STD_LOGIC;
    SIGNAL U1_OF_out_0 : STD_LOGIC;
    SIGNAL U1_OF_out_1 : STD_LOGIC;
    SIGNAL U1_OF_out_2 : STD_LOGIC;
    SIGNAL U1_OF_out_3 : STD_LOGIC;
    SIGNAL U1_PC_out_0 : STD_LOGIC;
    SIGNAL U1_PC_out_10 : STD_LOGIC;
    SIGNAL U1_PC_out_11 : STD_LOGIC;
    SIGNAL U1_PC_out_12 : STD_LOGIC;
    SIGNAL U1_PC_out_13 : STD_LOGIC;
    SIGNAL U1_PC_out_14 : STD_LOGIC;
    SIGNAL U1_PC_out_15 : STD_LOGIC;
    SIGNAL U1_PC_out_1 : STD_LOGIC;
    SIGNAL U1_PC_out_2 : STD_LOGIC;
    SIGNAL U1_PC_out_3 : STD_LOGIC;
    SIGNAL U1_PC_out_4 : STD_LOGIC;
    SIGNAL U1_PC_out_5 : STD_LOGIC;
    SIGNAL U1_PC_out_6 : STD_LOGIC;
    SIGNAL U1_PC_out_7 : STD_LOGIC;
    SIGNAL U1_PC_out_8 : STD_LOGIC;
    SIGNAL U1_PC_out_9 : STD_LOGIC;
    SIGNAL U1_SE12bits : STD_LOGIC;
    SIGNAL U1_SE4bits : STD_LOGIC;
    SIGNAL U1_SHF_0 : STD_LOGIC;
    SIGNAL U1_SHF_1 : STD_LOGIC;
    SIGNAL U1_V : STD_LOGIC;
    SIGNAL U1_V_out1 : STD_LOGIC;
    SIGNAL U1_Z : STD_LOGIC;
    SIGNAL U1_Z_out1 : STD_LOGIC;
    SIGNAL U1_addrBus_0 : STD_LOGIC;
    SIGNAL U1_addrBus_10 : STD_LOGIC;
    SIGNAL U1_addrBus_11 : STD_LOGIC;
    SIGNAL U1_addrBus_12 : STD_LOGIC;
    SIGNAL U1_addrBus_13 : STD_LOGIC;
    SIGNAL U1_addrBus_14 : STD_LOGIC;
    SIGNAL U1_addrBus_15 : STD_LOGIC;
    SIGNAL U1_addrBus_1 : STD_LOGIC;
    SIGNAL U1_addrBus_2 : STD_LOGIC;
    SIGNAL U1_addrBus_3 : STD_LOGIC;
    SIGNAL U1_addrBus_4 : STD_LOGIC;
    SIGNAL U1_addrBus_5 : STD_LOGIC;
    SIGNAL U1_addrBus_6 : STD_LOGIC;
    SIGNAL U1_addrBus_7 : STD_LOGIC;
    SIGNAL U1_addrBus_8 : STD_LOGIC;
    SIGNAL U1_addrBus_9 : STD_LOGIC;
    SIGNAL U1_clk : STD_LOGIC;
    SIGNAL U1_conOF : STD_LOGIC;
    SIGNAL U1_dataBus_0 : STD_LOGIC;
    SIGNAL U1_dataBus_10 : STD_LOGIC;
    SIGNAL U1_dataBus_11 : STD_LOGIC;
    SIGNAL U1_dataBus_12 : STD_LOGIC;
    SIGNAL U1_dataBus_13 : STD_LOGIC;
    SIGNAL U1_dataBus_14 : STD_LOGIC;
    SIGNAL U1_dataBus_15 : STD_LOGIC;
    SIGNAL U1_dataBus_1 : STD_LOGIC;
    SIGNAL U1_dataBus_2 : STD_LOGIC;
    SIGNAL U1_dataBus_3 : STD_LOGIC;
    SIGNAL U1_dataBus_4 : STD_LOGIC;
    SIGNAL U1_dataBus_5 : STD_LOGIC;
    SIGNAL U1_dataBus_6 : STD_LOGIC;
    SIGNAL U1_dataBus_7 : STD_LOGIC;
    SIGNAL U1_dataBus_8 : STD_LOGIC;
    SIGNAL U1_dataBus_9 : STD_LOGIC;
    SIGNAL U1_dataBus_out_0 : STD_LOGIC;
    SIGNAL U1_dataBus_out_10 : STD_LOGIC;
    SIGNAL U1_dataBus_out_11 : STD_LOGIC;
    SIGNAL U1_dataBus_out_12 : STD_LOGIC;
    SIGNAL U1_dataBus_out_13 : STD_LOGIC;
    SIGNAL U1_dataBus_out_14 : STD_LOGIC;
    SIGNAL U1_dataBus_out_15 : STD_LOGIC;
    SIGNAL U1_dataBus_out_1 : STD_LOGIC;
    SIGNAL U1_dataBus_out_2 : STD_LOGIC;
    SIGNAL U1_dataBus_out_3 : STD_LOGIC;
    SIGNAL U1_dataBus_out_4 : STD_LOGIC;
    SIGNAL U1_dataBus_out_5 : STD_LOGIC;
    SIGNAL U1_dataBus_out_6 : STD_LOGIC;
    SIGNAL U1_dataBus_out_7 : STD_LOGIC;
    SIGNAL U1_dataBus_out_8 : STD_LOGIC;
    SIGNAL U1_dataBus_out_9 : STD_LOGIC;
    SIGNAL U1_enSKP : STD_LOGIC;
    SIGNAL U1_ldAC : STD_LOGIC;
    SIGNAL U1_ldIN : STD_LOGIC;
    SIGNAL U1_ldIR : STD_LOGIC;
    SIGNAL U1_ldOF : STD_LOGIC;
    SIGNAL U1_ldPC : STD_LOGIC;
    SIGNAL U1_ldSR_0 : STD_LOGIC;
    SIGNAL U1_rst : STD_LOGIC;
    SIGNAL U1_sel1_ARU : STD_LOGIC;
    SIGNAL U1_selAC_MEM : STD_LOGIC;
    SIGNAL U1_selARU_AC : STD_LOGIC;
    SIGNAL U1_selIMM_AC : STD_LOGIC;
    SIGNAL U1_selIMM_LGU : STD_LOGIC;
    SIGNAL U1_selIMM_OF : STD_LOGIC;
    SIGNAL U1_selIMM_PC : STD_LOGIC;
    SIGNAL U1_selINC_IN : STD_LOGIC;
    SIGNAL U1_selINC_PC : STD_LOGIC;
    SIGNAL U1_selIN_MEM : STD_LOGIC;
    SIGNAL U1_selIR_MEM : STD_LOGIC;
    SIGNAL U1_selLGU_AC : STD_LOGIC;
    SIGNAL U1_selMEM_AC : STD_LOGIC;
    SIGNAL U1_selMEM_IN : STD_LOGIC;
    SIGNAL U1_selMEM_LGU : STD_LOGIC;
    SIGNAL U1_selMEM_PC : STD_LOGIC;
    SIGNAL U1_selMO_ARU : STD_LOGIC;
    SIGNAL U1_selPC_MEM : STD_LOGIC;
    SIGNAL U1_selPC_OF : STD_LOGIC;
    SIGNAL U1_selSET_SR : STD_LOGIC;
    SIGNAL U1_seldataBus : STD_LOGIC;
    SIGNAL U1_zeroAC : STD_LOGIC;
    SIGNAL U2_nstate_1 : STD_LOGIC;
    SIGNAL U2_pstate : STD_LOGIC;
    SIGNAL U2_readMEM : STD_LOGIC;

BEGIN
notg_1: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_INC1,
        out1 => S41
    );
nand_n_1: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_INC1,
        in1(1) => S0,
        out1 => S42
    );
nand_n_2: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S41,
        in1(1) => U1_PC_out_1,
        out1 => S43
    );
nand_n_3: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S43,
        in1(1) => S42,
        out1 => S27
    );
nand_n_4: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2,
        in1(1) => U1_INC1,
        out1 => S44
    );
nand_n_5: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1,
        in1(1) => S41,
        out1 => S45
    );
nand_n_6: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S45,
        in1(1) => S44,
        out1 => S28
    );
nand_n_7: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4,
        in1(1) => U1_INC1,
        out1 => S46
    );
nand_n_8: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3,
        in1(1) => S41,
        out1 => S47
    );
nand_n_9: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S47,
        in1(1) => S46,
        out1 => S29
    );
nand_n_10: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6,
        in1(1) => U1_INC1,
        out1 => S48
    );
nand_n_11: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5,
        in1(1) => S41,
        out1 => S49
    );
nand_n_12: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S49,
        in1(1) => S48,
        out1 => S30
    );
nand_n_13: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S8,
        in1(1) => U1_INC1,
        out1 => S50
    );
nand_n_14: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S7,
        in1(1) => S41,
        out1 => S51
    );
nand_n_15: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S51,
        in1(1) => S50,
        out1 => S31
    );
nand_n_16: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S10,
        in1(1) => U1_INC1,
        out1 => S52
    );
nand_n_17: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S9,
        in1(1) => S41,
        out1 => S53
    );
nand_n_18: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S53,
        in1(1) => S52,
        out1 => S32
    );
nand_n_19: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S12,
        in1(1) => U1_INC1,
        out1 => S54
    );
nand_n_20: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S11,
        in1(1) => S41,
        out1 => S55
    );
nand_n_21: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S55,
        in1(1) => S54,
        out1 => S33
    );
nand_n_22: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S14,
        in1(1) => U1_INC1,
        out1 => S56
    );
nand_n_23: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S13,
        in1(1) => S41,
        out1 => S57
    );
nand_n_24: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S57,
        in1(1) => S56,
        out1 => S34
    );
nand_n_25: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S16,
        in1(1) => U1_INC1,
        out1 => S58
    );
nand_n_26: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S15,
        in1(1) => S41,
        out1 => S59
    );
nand_n_27: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S59,
        in1(1) => S58,
        out1 => S35
    );
nand_n_28: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S18,
        in1(1) => U1_INC1,
        out1 => S60
    );
nand_n_29: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S17,
        in1(1) => S41,
        out1 => S61
    );
nand_n_30: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S61,
        in1(1) => S60,
        out1 => S36
    );
nand_n_31: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S20,
        in1(1) => U1_INC1,
        out1 => S62
    );
nand_n_32: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S19,
        in1(1) => S41,
        out1 => S63
    );
nand_n_33: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S63,
        in1(1) => S62,
        out1 => S37
    );
nand_n_34: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S22,
        in1(1) => U1_INC1,
        out1 => S64
    );
nand_n_35: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S21,
        in1(1) => S41,
        out1 => S65
    );
nand_n_36: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S65,
        in1(1) => S64,
        out1 => S38
    );
nand_n_37: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S24,
        in1(1) => U1_INC1,
        out1 => S66
    );
nand_n_38: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S23,
        in1(1) => S41,
        out1 => S67
    );
nand_n_39: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S67,
        in1(1) => S66,
        out1 => S39
    );
nand_n_40: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S26,
        in1(1) => U1_INC1,
        out1 => S68
    );
nand_n_41: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S25,
        in1(1) => S41,
        out1 => S69
    );
nand_n_42: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S69,
        in1(1) => S68,
        out1 => S40
    );
nor_n_1: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S754,
        in1(1) => S1925,
        out1 => S755
    );
nor_n_2: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S755,
        in1(1) => S750,
        out1 => S756
    );
nor_n_3: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S756,
        in1(1) => U1_AC_out_2,
        out1 => S757
    );
nand_n_43: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S745,
        in1(1) => U1_AC_out_2,
        out1 => S758
    );
nand_n_44: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S758,
        in1(1) => S2029,
        out1 => S759
    );
nor_n_4: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S759,
        in1(1) => S757,
        out1 => S760
    );
nor_n_5: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S760,
        in1(1) => S1939,
        out1 => S761
    );
nor_n_6: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S761,
        in1(1) => S2249,
        out1 => S762
    );
nand_n_45: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S762,
        in1(1) => S736,
        out1 => S763
    );
nor_n_7: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2106,
        in1(1) => S1959,
        out1 => S764
    );
nor_n_8: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S764,
        in1(1) => U1_AND,
        out1 => S765
    );
nand_n_46: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S765,
        in1(1) => S763,
        out1 => S766
    );
nand_n_47: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S602,
        in1(1) => U1_AND,
        out1 => S767
    );
nand_n_48: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S767,
        in1(1) => S766,
        out1 => S768
    );
notg_2: ENTITY WORK.notg
    PORT MAP (
        in1 => S768,
        out1 => S769
    );
nand_n_49: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S625,
        in1(1) => U1_AND,
        out1 => S770
    );
nor_n_9: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2061,
        in1(1) => S1959,
        out1 => S771
    );
nor_n_10: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S771,
        in1(1) => U1_AND,
        out1 => S772
    );
nor_n_11: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_SHF_1,
        in1(1) => S1932,
        out1 => S773
    );
nand_n_50: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1940,
        in1(1) => U1_AC_out_2,
        out1 => S774
    );
nand_n_51: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S773,
        in1(1) => S712,
        out1 => S775
    );
notg_3: ENTITY WORK.notg
    PORT MAP (
        in1 => S775,
        out1 => S776
    );
nand_n_52: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S723,
        in1(1) => S718,
        out1 => S777
    );
notg_4: ENTITY WORK.notg
    PORT MAP (
        in1 => S777,
        out1 => S778
    );
nor_n_12: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S778,
        in1(1) => U1_AC_out_1,
        out1 => S779
    );
nand_n_53: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S777,
        in1(1) => S1925,
        out1 => S780
    );
nand_n_54: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S717,
        in1(1) => S714,
        out1 => S781
    );
notg_5: ENTITY WORK.notg
    PORT MAP (
        in1 => S781,
        out1 => S782
    );
nand_n_55: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S781,
        in1(1) => U1_AC_out_1,
        out1 => S783
    );
notg_6: ENTITY WORK.notg
    PORT MAP (
        in1 => S783,
        out1 => S784
    );
nor_n_13: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S784,
        in1(1) => S779,
        out1 => S785
    );
nand_n_56: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S783,
        in1(1) => S780,
        out1 => S786
    );
nor_n_14: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S786,
        in1(1) => S2100,
        out1 => S787
    );
nor_n_15: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S787,
        in1(1) => S776,
        out1 => S788
    );
nand_n_57: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S756,
        in1(1) => U1_AC_out_2,
        out1 => S789
    );
nor_n_16: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S731,
        in1(1) => U1_AC_out_2,
        out1 => S790
    );
nor_n_17: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S790,
        in1(1) => U1_AC_out_3,
        out1 => S791
    );
nand_n_58: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S791,
        in1(1) => S789,
        out1 => S792
    );
nand_n_59: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S792,
        in1(1) => S2029,
        out1 => S793
    );
nand_n_60: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S793,
        in1(1) => S788,
        out1 => S794
    );
nor_n_18: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S745,
        in1(1) => S2111,
        out1 => S795
    );
nor_n_19: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S795,
        in1(1) => S1939,
        out1 => S796
    );
nor_n_20: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S796,
        in1(1) => S2249,
        out1 => S797
    );
nand_n_61: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S797,
        in1(1) => S794,
        out1 => S798
    );
nand_n_62: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S798,
        in1(1) => S772,
        out1 => S799
    );
nand_n_63: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S799,
        in1(1) => S770,
        out1 => S800
    );
nand_n_64: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S636,
        in1(1) => U1_AND,
        out1 => S801
    );
nor_n_21: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2082,
        in1(1) => S1959,
        out1 => S802
    );
nor_n_22: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S802,
        in1(1) => U1_AND,
        out1 => S803
    );
nor_n_23: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S782,
        in1(1) => U1_AC_out_1,
        out1 => S804
    );
nand_n_65: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S781,
        in1(1) => S1925,
        out1 => S805
    );
nand_n_66: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S711,
        in1(1) => U1_AC_out_1,
        out1 => S806
    );
notg_7: ENTITY WORK.notg
    PORT MAP (
        in1 => S806,
        out1 => S807
    );
nor_n_24: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S807,
        in1(1) => S804,
        out1 => S808
    );
nand_n_67: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S806,
        in1(1) => S805,
        out1 => S809
    );
nor_n_25: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S809,
        in1(1) => S774,
        out1 => S810
    );
nand_n_68: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S727,
        in1(1) => S724,
        out1 => S811
    );
nand_n_69: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S811,
        in1(1) => S1925,
        out1 => S812
    );
nand_n_70: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S777,
        in1(1) => U1_AC_out_1,
        out1 => S813
    );
nand_n_71: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S813,
        in1(1) => S812,
        out1 => S814
    );
nor_n_26: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S814,
        in1(1) => S2100,
        out1 => S815
    );
nor_n_27: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S815,
        in1(1) => S810,
        out1 => S816
    );
nor_n_28: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S754,
        in1(1) => U1_AC_out_1,
        out1 => S817
    );
nor_n_29: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S739,
        in1(1) => S1925,
        out1 => S818
    );
nor_n_30: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S818,
        in1(1) => S817,
        out1 => S819
    );
nand_n_72: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S819,
        in1(1) => U1_AC_out_2,
        out1 => S820
    );
nand_n_73: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S729,
        in1(1) => S1925,
        out1 => S821
    );
nand_n_74: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S748,
        in1(1) => U1_AC_out_1,
        out1 => S822
    );
nand_n_75: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S822,
        in1(1) => S821,
        out1 => S823
    );
nor_n_31: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S823,
        in1(1) => U1_AC_out_2,
        out1 => S824
    );
nor_n_32: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S824,
        in1(1) => U1_AC_out_3,
        out1 => S825
    );
nand_n_76: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S825,
        in1(1) => S820,
        out1 => S826
    );
nand_n_77: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S826,
        in1(1) => S2029,
        out1 => S827
    );
nand_n_78: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S827,
        in1(1) => S816,
        out1 => S828
    );
nand_n_79: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S742,
        in1(1) => S1925,
        out1 => S829
    );
nor_n_33: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S829,
        in1(1) => S2111,
        out1 => S830
    );
nor_n_34: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S830,
        in1(1) => S1939,
        out1 => S831
    );
nor_n_35: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S831,
        in1(1) => S2249,
        out1 => S832
    );
nand_n_80: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S832,
        in1(1) => S828,
        out1 => S833
    );
nand_n_81: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S833,
        in1(1) => S803,
        out1 => S834
    );
nand_n_82: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S834,
        in1(1) => S801,
        out1 => S835
    );
nand_n_83: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S523,
        in1(1) => U1_AND,
        out1 => S836
    );
nand_n_84: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S816,
        in1(1) => U1_AC_out_3,
        out1 => S837
    );
nand_n_85: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S753,
        in1(1) => S747,
        out1 => S838
    );
nand_n_86: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S838,
        in1(1) => S1925,
        out1 => S839
    );
nand_n_87: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S746,
        in1(1) => S728,
        out1 => S840
    );
nand_n_88: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S840,
        in1(1) => U1_AC_out_1,
        out1 => S841
    );
nand_n_89: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S841,
        in1(1) => S839,
        out1 => S842
    );
notg_8: ENTITY WORK.notg
    PORT MAP (
        in1 => S842,
        out1 => S843
    );
nor_n_36: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S842,
        in1(1) => S774,
        out1 => S844
    );
nor_n_37: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_SHF_1,
        in1(1) => S1939,
        out1 => S845
    );
nand_n_90: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1940,
        in1(1) => U1_AC_out_3,
        out1 => S846
    );
nor_n_38: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S845,
        in1(1) => S830,
        out1 => S847
    );
nor_n_39: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S751,
        in1(1) => S737,
        out1 => S848
    );
nand_n_91: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S848,
        in1(1) => U1_AC_out_1,
        out1 => S849
    );
nand_n_92: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2175,
        in1(1) => U1_AC_out_0,
        out1 => S850
    );
nand_n_93: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S850,
        in1(1) => S743,
        out1 => S851
    );
nand_n_94: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S851,
        in1(1) => S1925,
        out1 => S852
    );
nand_n_95: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S852,
        in1(1) => S849,
        out1 => S853
    );
nand_n_96: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S853,
        in1(1) => S2099,
        out1 => S854
    );
nand_n_97: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S854,
        in1(1) => S847,
        out1 => S855
    );
nor_n_40: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S855,
        in1(1) => S844,
        out1 => S856
    );
nor_n_41: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S856,
        in1(1) => S2249,
        out1 => S857
    );
nand_n_98: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S857,
        in1(1) => S837,
        out1 => S858
    );
nor_n_42: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2185,
        in1(1) => S1959,
        out1 => S859
    );
nor_n_43: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S859,
        in1(1) => U1_AND,
        out1 => S860
    );
nand_n_99: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S860,
        in1(1) => S858,
        out1 => S861
    );
nand_n_100: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S861,
        in1(1) => S836,
        out1 => S862
    );
nor_n_44: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2222,
        in1(1) => S2211,
        out1 => S863
    );
nand_n_101: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2237,
        in1(1) => S2152,
        out1 => S864
    );
nand_n_102: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2192,
        in1(1) => S2110,
        out1 => S865
    );
nand_n_103: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S865,
        in1(1) => S846,
        out1 => S866
    );
nor_n_45: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2202,
        in1(1) => S2086,
        out1 => S867
    );
nor_n_46: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S867,
        in1(1) => U1_AC_out_1,
        out1 => S868
    );
nand_n_104: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2077,
        in1(1) => S2065,
        out1 => S869
    );
nor_n_47: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S869,
        in1(1) => S1925,
        out1 => S870
    );
nor_n_48: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S870,
        in1(1) => S868,
        out1 => S871
    );
nand_n_105: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S871,
        in1(1) => S773,
        out1 => S872
    );
nand_n_106: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S863,
        in1(1) => U1_AC_out_1,
        out1 => S873
    );
notg_9: ENTITY WORK.notg
    PORT MAP (
        in1 => S873,
        out1 => S874
    );
nor_n_49: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S864,
        in1(1) => U1_AC_out_1,
        out1 => S875
    );
nor_n_50: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S875,
        in1(1) => S874,
        out1 => S876
    );
nor_n_51: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S876,
        in1(1) => S2100,
        out1 => S877
    );
nor_n_52: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S877,
        in1(1) => S866,
        out1 => S878
    );
nand_n_107: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S878,
        in1(1) => S872,
        out1 => S879
    );
nand_n_108: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S773,
        in1(1) => S2097,
        out1 => S880
    );
nand_n_109: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2129,
        in1(1) => S2056,
        out1 => S881
    );
nor_n_53: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S881,
        in1(1) => U1_AC_out_1,
        out1 => S882
    );
nand_n_110: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2120,
        in1(1) => S2109,
        out1 => S883
    );
nor_n_54: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S883,
        in1(1) => S1925,
        out1 => S884
    );
nor_n_55: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S884,
        in1(1) => S882,
        out1 => S885
    );
nand_n_111: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S885,
        in1(1) => S2099,
        out1 => S886
    );
nand_n_112: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S886,
        in1(1) => S880,
        out1 => S887
    );
notg_10: ENTITY WORK.notg
    PORT MAP (
        in1 => S887,
        out1 => S888
    );
nor_n_56: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S887,
        in1(1) => S1939,
        out1 => S889
    );
nor_n_57: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S889,
        in1(1) => S2249,
        out1 => S890
    );
nand_n_113: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S890,
        in1(1) => S879,
        out1 => S891
    );
nor_n_58: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2148,
        in1(1) => S1959,
        out1 => S892
    );
nor_n_59: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S892,
        in1(1) => U1_AND,
        out1 => S893
    );
nand_n_114: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S893,
        in1(1) => S891,
        out1 => S894
    );
nand_n_115: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2613,
        in1(1) => U1_AND,
        out1 => S895
    );
nand_n_116: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S895,
        in1(1) => S894,
        out1 => S896
    );
nand_n_117: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S608,
        in1(1) => U1_AND,
        out1 => S897
    );
nor_n_60: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2116,
        in1(1) => S1959,
        out1 => S898
    );
nor_n_61: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S898,
        in1(1) => U1_AND,
        out1 => S899
    );
nand_n_118: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2067,
        in1(1) => U1_AC_out_1,
        out1 => S900
    );
nor_n_62: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2130,
        in1(1) => U1_AC_out_1,
        out1 => S901
    );
nor_n_63: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2087,
        in1(1) => U1_AC_out_1,
        out1 => S902
    );
nor_n_64: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2212,
        in1(1) => S1925,
        out1 => S903
    );
nor_n_65: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S903,
        in1(1) => S902,
        out1 => S904
    );
nor_n_66: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S901,
        in1(1) => U1_AC_out_2,
        out1 => S905
    );
nand_n_119: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S905,
        in1(1) => S900,
        out1 => S906
    );
nand_n_120: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S904,
        in1(1) => U1_AC_out_2,
        out1 => S907
    );
nand_n_121: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S907,
        in1(1) => S906,
        out1 => S908
    );
nor_n_67: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S908,
        in1(1) => U1_AC_out_3,
        out1 => S909
    );
nor_n_68: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S909,
        in1(1) => S2030,
        out1 => S910
    );
nor_n_69: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S883,
        in1(1) => U1_AC_out_1,
        out1 => S911
    );
nor_n_70: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2095,
        in1(1) => S1925,
        out1 => S912
    );
nor_n_71: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S912,
        in1(1) => S911,
        out1 => S913
    );
nand_n_122: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S913,
        in1(1) => S2099,
        out1 => S914
    );
notg_11: ENTITY WORK.notg
    PORT MAP (
        in1 => S914,
        out1 => S915
    );
nor_n_72: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S915,
        in1(1) => S910,
        out1 => S916
    );
nor_n_73: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2189,
        in1(1) => U1_AC_out_1,
        out1 => S917
    );
nand_n_123: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S917,
        in1(1) => U1_AC_out_2,
        out1 => S918
    );
nor_n_74: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2238,
        in1(1) => U1_AC_out_1,
        out1 => S919
    );
nand_n_124: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2164,
        in1(1) => U1_AC_out_1,
        out1 => S920
    );
notg_12: ENTITY WORK.notg
    PORT MAP (
        in1 => S920,
        out1 => S921
    );
nor_n_75: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S921,
        in1(1) => S919,
        out1 => S922
    );
nand_n_125: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S922,
        in1(1) => S1932,
        out1 => S923
    );
nand_n_126: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S923,
        in1(1) => S918,
        out1 => S924
    );
nand_n_127: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S924,
        in1(1) => S2029,
        out1 => S925
    );
nand_n_128: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S925,
        in1(1) => U1_AC_out_3,
        out1 => S926
    );
nor_n_76: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S916,
        in1(1) => S2249,
        out1 => S927
    );
nand_n_129: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S927,
        in1(1) => S926,
        out1 => S928
    );
nand_n_130: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S928,
        in1(1) => S899,
        out1 => S929
    );
nand_n_131: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S929,
        in1(1) => S897,
        out1 => S930
    );
nand_n_132: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S613,
        in1(1) => U1_AND,
        out1 => S931
    );
nor_n_77: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2125,
        in1(1) => S1959,
        out1 => S932
    );
nor_n_78: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S932,
        in1(1) => U1_AND,
        out1 => S933
    );
nand_n_133: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S808,
        in1(1) => S2099,
        out1 => S934
    );
nand_n_134: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S725,
        in1(1) => U1_AC_out_1,
        out1 => S935
    );
nand_n_135: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S719,
        in1(1) => S1925,
        out1 => S936
    );
nand_n_136: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S936,
        in1(1) => S935,
        out1 => S937
    );
nand_n_137: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S937,
        in1(1) => S1932,
        out1 => S938
    );
nand_n_138: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S823,
        in1(1) => U1_AC_out_2,
        out1 => S939
    );
nand_n_139: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S939,
        in1(1) => S938,
        out1 => S940
    );
nand_n_140: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S940,
        in1(1) => S1939,
        out1 => S941
    );
nand_n_141: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S941,
        in1(1) => S2029,
        out1 => S942
    );
nand_n_142: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S942,
        in1(1) => S934,
        out1 => S943
    );
nor_n_79: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S819,
        in1(1) => U1_AC_out_2,
        out1 => S944
    );
nand_n_143: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S829,
        in1(1) => U1_AC_out_2,
        out1 => S945
    );
nand_n_144: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S945,
        in1(1) => S2029,
        out1 => S946
    );
nor_n_80: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S946,
        in1(1) => S944,
        out1 => S947
    );
nor_n_81: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S947,
        in1(1) => S1939,
        out1 => S948
    );
nor_n_82: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S948,
        in1(1) => S2249,
        out1 => S949
    );
nand_n_145: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S949,
        in1(1) => S943,
        out1 => S950
    );
nand_n_146: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S950,
        in1(1) => S933,
        out1 => S951
    );
nand_n_147: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S951,
        in1(1) => S931,
        out1 => S952
    );
nand_n_148: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2546,
        in1(1) => U1_AND,
        out1 => S953
    );
nand_n_149: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S843,
        in1(1) => S2099,
        out1 => S954
    );
nor_n_83: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S814,
        in1(1) => S774,
        out1 => S955
    );
nor_n_84: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S955,
        in1(1) => S845,
        out1 => S956
    );
nand_n_150: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S956,
        in1(1) => S954,
        out1 => S957
    );
nor_n_85: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S957,
        in1(1) => S947,
        out1 => S958
    );
nand_n_151: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S934,
        in1(1) => U1_AC_out_3,
        out1 => S959
    );
nand_n_152: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S959,
        in1(1) => S2248,
        out1 => S960
    );
nor_n_86: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S960,
        in1(1) => S958,
        out1 => S961
    );
notg_13: ENTITY WORK.notg
    PORT MAP (
        in1 => S961,
        out1 => S962
    );
nor_n_87: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2232,
        in1(1) => S1959,
        out1 => S963
    );
nor_n_88: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S963,
        in1(1) => U1_AND,
        out1 => S964
    );
nand_n_153: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S964,
        in1(1) => S962,
        out1 => S965
    );
nand_n_154: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S965,
        in1(1) => S953,
        out1 => S966
    );
nand_n_155: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S623,
        in1(1) => U1_AND,
        out1 => S967
    );
nor_n_89: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2053,
        in1(1) => S1959,
        out1 => S968
    );
nor_n_90: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S968,
        in1(1) => U1_AND,
        out1 => S969
    );
nand_n_156: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2242,
        in1(1) => U1_AC_out_2,
        out1 => S970
    );
nand_n_157: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S970,
        in1(1) => S1939,
        out1 => S971
    );
nand_n_158: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S971,
        in1(1) => S2029,
        out1 => S972
    );
nor_n_91: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2111,
        in1(1) => S2090,
        out1 => S973
    );
nand_n_159: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S972,
        in1(1) => S888,
        out1 => S974
    );
nor_n_92: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S974,
        in1(1) => S973,
        out1 => S975
    );
nand_n_160: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S865,
        in1(1) => U1_AC_out_3,
        out1 => S976
    );
nor_n_93: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S975,
        in1(1) => S2249,
        out1 => S977
    );
nand_n_161: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S977,
        in1(1) => S976,
        out1 => S978
    );
nand_n_162: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S978,
        in1(1) => S969,
        out1 => S979
    );
nand_n_163: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S979,
        in1(1) => S967,
        out1 => S980
    );
nand_n_164: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S634,
        in1(1) => U1_AND,
        out1 => S981
    );
nor_n_94: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2073,
        in1(1) => S1959,
        out1 => S982
    );
nor_n_95: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S982,
        in1(1) => U1_AND,
        out1 => S983
    );
nand_n_165: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S922,
        in1(1) => U1_AC_out_2,
        out1 => S984
    );
notg_14: ENTITY WORK.notg
    PORT MAP (
        in1 => S984,
        out1 => S985
    );
nor_n_96: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S985,
        in1(1) => U1_AC_out_3,
        out1 => S986
    );
nor_n_97: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S986,
        in1(1) => S2030,
        out1 => S987
    );
nand_n_166: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S904,
        in1(1) => S2110,
        out1 => S988
    );
nor_n_98: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S869,
        in1(1) => U1_AC_out_1,
        out1 => S989
    );
nor_n_99: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S881,
        in1(1) => S1925,
        out1 => S990
    );
nor_n_100: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S990,
        in1(1) => S989,
        out1 => S991
    );
nand_n_167: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S991,
        in1(1) => S2099,
        out1 => S992
    );
nand_n_168: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S913,
        in1(1) => S773,
        out1 => S993
    );
nand_n_169: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S993,
        in1(1) => S992,
        out1 => S994
    );
notg_15: ENTITY WORK.notg
    PORT MAP (
        in1 => S994,
        out1 => S995
    );
nand_n_170: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S995,
        in1(1) => S988,
        out1 => S996
    );
nor_n_101: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S996,
        in1(1) => S987,
        out1 => S997
    );
nand_n_171: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S917,
        in1(1) => S2110,
        out1 => S998
    );
nand_n_172: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S998,
        in1(1) => U1_AC_out_3,
        out1 => S999
    );
nor_n_102: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S997,
        in1(1) => S2249,
        out1 => S1000
    );
nand_n_173: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1000,
        in1(1) => S999,
        out1 => S1001
    );
nand_n_174: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1001,
        in1(1) => S983,
        out1 => S1002
    );
nand_n_175: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1002,
        in1(1) => S981,
        out1 => S1003
    );
notg_16: ENTITY WORK.notg
    PORT MAP (
        in1 => S1003,
        out1 => S1004
    );
nand_n_176: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2294,
        in1(1) => U1_AND,
        out1 => S1005
    );
nor_n_103: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2207,
        in1(1) => S1959,
        out1 => S1006
    );
nor_n_104: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1006,
        in1(1) => U1_AND,
        out1 => S1007
    );
nand_n_177: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S785,
        in1(1) => S773,
        out1 => S1008
    );
nand_n_178: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S840,
        in1(1) => S1925,
        out1 => S1009
    );
nand_n_179: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S811,
        in1(1) => U1_AC_out_1,
        out1 => S1010
    );
nand_n_180: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1010,
        in1(1) => S1009,
        out1 => S1011
    );
nor_n_105: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1011,
        in1(1) => S2100,
        out1 => S1012
    );
nor_n_106: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1012,
        in1(1) => S845,
        out1 => S1013
    );
nand_n_181: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1013,
        in1(1) => S1008,
        out1 => S1014
    );
nor_n_107: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1014,
        in1(1) => S760,
        out1 => S1015
    );
nand_n_182: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S713,
        in1(1) => U1_AC_out_3,
        out1 => S1016
    );
nor_n_108: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1015,
        in1(1) => S2249,
        out1 => S1017
    );
nand_n_183: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1017,
        in1(1) => S1016,
        out1 => S1018
    );
nand_n_184: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1018,
        in1(1) => S1007,
        out1 => S1019
    );
nand_n_185: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1019,
        in1(1) => S1005,
        out1 => S1020
    );
nand_n_186: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S788,
        in1(1) => U1_AC_out_3,
        out1 => S1021
    );
nor_n_109: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1011,
        in1(1) => S774,
        out1 => S1022
    );
nor_n_110: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S845,
        in1(1) => S795,
        out1 => S1023
    );
nand_n_187: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S838,
        in1(1) => U1_AC_out_1,
        out1 => S1024
    );
nor_n_111: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S848,
        in1(1) => U1_AC_out_1,
        out1 => S1025
    );
nor_n_112: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1025,
        in1(1) => S2100,
        out1 => S1026
    );
nand_n_188: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1026,
        in1(1) => S1024,
        out1 => S1027
    );
nand_n_189: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1027,
        in1(1) => S1023,
        out1 => S1028
    );
nor_n_113: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1028,
        in1(1) => S1022,
        out1 => S1029
    );
nor_n_114: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1029,
        in1(1) => S2249,
        out1 => S1030
    );
nand_n_190: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1030,
        in1(1) => S1021,
        out1 => S1031
    );
nor_n_115: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2159,
        in1(1) => S1959,
        out1 => S1032
    );
nor_n_116: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1032,
        in1(1) => U1_AND,
        out1 => S1033
    );
nand_n_191: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1033,
        in1(1) => S1031,
        out1 => S1034
    );
nand_n_192: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S361,
        in1(1) => U1_AND,
        out1 => S1035
    );
nand_n_193: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1035,
        in1(1) => S1034,
        out1 => S1036
    );
nor_n_117: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S863,
        in1(1) => U1_AC_out_1,
        out1 => S1037
    );
nor_n_118: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S867,
        in1(1) => S1925,
        out1 => S1038
    );
nor_n_119: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1038,
        in1(1) => S1037,
        out1 => S1039
    );
nor_n_120: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1039,
        in1(1) => S1932,
        out1 => S1040
    );
nand_n_194: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2177,
        in1(1) => S2163,
        out1 => S1041
    );
nand_n_195: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1041,
        in1(1) => S1925,
        out1 => S1042
    );
nand_n_196: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S864,
        in1(1) => U1_AC_out_1,
        out1 => S1043
    );
nand_n_197: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1043,
        in1(1) => S1042,
        out1 => S1044
    );
nand_n_198: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1044,
        in1(1) => S1932,
        out1 => S1045
    );
nand_n_199: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1045,
        in1(1) => S1940,
        out1 => S1046
    );
nor_n_121: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1046,
        in1(1) => S1040,
        out1 => S1047
    );
nand_n_200: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S998,
        in1(1) => S846,
        out1 => S1048
    );
nor_n_122: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1048,
        in1(1) => S1047,
        out1 => S1049
    );
nand_n_201: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S995,
        in1(1) => U1_AC_out_3,
        out1 => S1050
    );
nand_n_202: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1050,
        in1(1) => S2248,
        out1 => S1051
    );
nor_n_123: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1051,
        in1(1) => S1049,
        out1 => S1052
    );
nor_n_124: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2173,
        in1(1) => S1959,
        out1 => S1053
    );
nor_n_125: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1053,
        in1(1) => S1052,
        out1 => S1054
    );
nor_n_126: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1054,
        in1(1) => U1_AND,
        out1 => S1055
    );
nand_n_203: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2173,
        in1(1) => U1_AND,
        out1 => S1056
    );
nor_n_127: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1056,
        in1(1) => S1925,
        out1 => S1057
    );
nor_n_128: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1057,
        in1(1) => S1055,
        out1 => S1058
    );
nand_n_204: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2418,
        in1(1) => U1_AND,
        out1 => S1059
    );
nand_n_205: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S885,
        in1(1) => S773,
        out1 => S1060
    );
nand_n_206: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S871,
        in1(1) => S2099,
        out1 => S1061
    );
nand_n_207: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1060,
        in1(1) => S846,
        out1 => S1062
    );
nor_n_129: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1062,
        in1(1) => S2246,
        out1 => S1063
    );
nand_n_208: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1063,
        in1(1) => S1061,
        out1 => S1064
    );
nand_n_209: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2101,
        in1(1) => U1_AC_out_3,
        out1 => S1065
    );
notg_17: ENTITY WORK.notg
    PORT MAP (
        in1 => S1065,
        out1 => S1066
    );
nor_n_130: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1066,
        in1(1) => S2249,
        out1 => S1067
    );
nand_n_210: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1067,
        in1(1) => S1064,
        out1 => S1068
    );
nor_n_131: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2198,
        in1(1) => S1959,
        out1 => S1069
    );
nor_n_132: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1069,
        in1(1) => U1_AND,
        out1 => S1070
    );
nand_n_211: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1070,
        in1(1) => S1068,
        out1 => S1071
    );
nand_n_212: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1071,
        in1(1) => S1059,
        out1 => S1072
    );
nand_n_213: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2329,
        in1(1) => U1_AND,
        out1 => S1073
    );
nand_n_214: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1039,
        in1(1) => S2099,
        out1 => S1074
    );
nand_n_215: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S991,
        in1(1) => S773,
        out1 => S1075
    );
nand_n_216: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1075,
        in1(1) => S1074,
        out1 => S1076
    );
nor_n_133: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1076,
        in1(1) => S845,
        out1 => S1077
    );
nand_n_217: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1077,
        in1(1) => S925,
        out1 => S1078
    );
nand_n_218: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S914,
        in1(1) => U1_AC_out_3,
        out1 => S1079
    );
notg_18: ENTITY WORK.notg
    PORT MAP (
        in1 => S1079,
        out1 => S1080
    );
nor_n_134: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1080,
        in1(1) => S2249,
        out1 => S1081
    );
nand_n_219: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1081,
        in1(1) => S1078,
        out1 => S1082
    );
nor_n_135: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2218,
        in1(1) => S1959,
        out1 => S1083
    );
nor_n_136: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1083,
        in1(1) => U1_AND,
        out1 => S1084
    );
nand_n_220: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1084,
        in1(1) => S1082,
        out1 => S1085
    );
nand_n_221: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1085,
        in1(1) => S1073,
        out1 => S1086
    );
nand_n_222: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S862,
        in1(1) => S2253,
        out1 => S1087
    );
notg_19: ENTITY WORK.notg
    PORT MAP (
        in1 => S1087,
        out1 => S1088
    );
nand_n_223: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1088,
        in1(1) => S1036,
        out1 => S1089
    );
nor_n_137: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1089,
        in1(1) => S769,
        out1 => S1090
    );
nand_n_224: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1086,
        in1(1) => S966,
        out1 => S1091
    );
nor_n_138: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1091,
        in1(1) => S1004,
        out1 => S1092
    );
nand_n_225: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1092,
        in1(1) => S980,
        out1 => S1093
    );
nand_n_226: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1072,
        in1(1) => S835,
        out1 => S1094
    );
nand_n_227: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S930,
        in1(1) => S800,
        out1 => S1095
    );
nor_n_139: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1095,
        in1(1) => S1094,
        out1 => S1096
    );
nand_n_228: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1020,
        in1(1) => S952,
        out1 => S1097
    );
nand_n_229: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1058,
        in1(1) => S896,
        out1 => S1098
    );
nor_n_140: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1098,
        in1(1) => S1097,
        out1 => S1099
    );
nand_n_230: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1099,
        in1(1) => S1096,
        out1 => S1100
    );
nor_n_141: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1100,
        in1(1) => S1093,
        out1 => S1101
    );
nand_n_231: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1101,
        in1(1) => S1090,
        out1 => S1102
    );
notg_20: ENTITY WORK.notg
    PORT MAP (
        in1 => S1102,
        out1 => U1_Z
    );
nand_n_232: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1966,
        in1(1) => U1_INC1,
        out1 => S1103
    );
nand_n_233: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_PC_out_0,
        in1(1) => S1965,
        out1 => S1104
    );
nand_n_234: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1104,
        in1(1) => S1103,
        out1 => S1105
    );
nand_n_235: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1105,
        in1(1) => U1_selPC_MEM,
        out1 => S1106
    );
nand_n_236: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1996,
        in1(1) => U1_IN_out_0,
        out1 => S1107
    );
nand_n_237: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1107,
        in1(1) => S1106,
        out1 => S1108
    );
nand_n_238: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1108,
        in1(1) => S1997,
        out1 => S1109
    );
nand_n_239: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selAC_MEM,
        in1(1) => U1_AC_out_0,
        out1 => S1110
    );
nand_n_240: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1110,
        in1(1) => S1109,
        out1 => U1_dataBus_out_0
    );
nand_n_241: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_PC_out_1,
        in1(1) => U1_INC1,
        out1 => S1111
    );
nor_n_142: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_PC_out_1,
        in1(1) => U1_INC1,
        out1 => S1112
    );
nor_n_143: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1112,
        in1(1) => U1_PC_out_0,
        out1 => S1113
    );
nand_n_242: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1113,
        in1(1) => S1111,
        out1 => S1114
    );
nand_n_243: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1114,
        in1(1) => S2254,
        out1 => S1115
    );
nor_n_144: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1115,
        in1(1) => S1996,
        out1 => S1116
    );
nand_n_244: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_IN_out_1,
        in1(1) => S1996,
        out1 => S1117
    );
nor_n_145: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1997,
        in1(1) => U1_AC_out_1,
        out1 => S1118
    );
nand_n_245: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1117,
        in1(1) => S1997,
        out1 => S1119
    );
nor_n_146: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1119,
        in1(1) => S1116,
        out1 => S1120
    );
nor_n_147: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1120,
        in1(1) => S1118,
        out1 => U1_dataBus_out_1
    );
nand_n_246: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1970,
        in1(1) => S27,
        out1 => S1121
    );
nand_n_247: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_PC_out_2,
        in1(1) => S1969,
        out1 => S1122
    );
nand_n_248: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1122,
        in1(1) => S1121,
        out1 => S1123
    );
nand_n_249: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1123,
        in1(1) => U1_selPC_MEM,
        out1 => S1124
    );
nand_n_250: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_IN_out_2,
        in1(1) => S1996,
        out1 => S1125
    );
nand_n_251: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1125,
        in1(1) => S1124,
        out1 => S1126
    );
nand_n_252: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1126,
        in1(1) => S1997,
        out1 => S1127
    );
nand_n_253: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selAC_MEM,
        in1(1) => U1_AC_out_2,
        out1 => S1128
    );
nand_n_254: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1128,
        in1(1) => S1127,
        out1 => U1_dataBus_out_2
    );
nand_n_255: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1972,
        in1(1) => S28,
        out1 => S1129
    );
nand_n_256: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_PC_out_3,
        in1(1) => S1971,
        out1 => S1130
    );
nand_n_257: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1130,
        in1(1) => S1129,
        out1 => S1131
    );
nand_n_258: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1131,
        in1(1) => U1_selPC_MEM,
        out1 => S1132
    );
nand_n_259: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_IN_out_3,
        in1(1) => S1996,
        out1 => S1133
    );
nand_n_260: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1133,
        in1(1) => S1132,
        out1 => S1134
    );
nand_n_261: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1134,
        in1(1) => S1997,
        out1 => S1135
    );
nand_n_262: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selAC_MEM,
        in1(1) => U1_AC_out_3,
        out1 => S1136
    );
nand_n_263: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1136,
        in1(1) => S1135,
        out1 => U1_dataBus_out_3
    );
nand_n_264: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1974,
        in1(1) => S29,
        out1 => S1137
    );
nand_n_265: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_PC_out_4,
        in1(1) => S1973,
        out1 => S1138
    );
nand_n_266: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1138,
        in1(1) => S1137,
        out1 => S1139
    );
nand_n_267: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1139,
        in1(1) => U1_selPC_MEM,
        out1 => S1140
    );
nand_n_268: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_IN_out_4,
        in1(1) => S1996,
        out1 => S1141
    );
nand_n_269: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1141,
        in1(1) => S1140,
        out1 => S1142
    );
nand_n_270: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1142,
        in1(1) => S1997,
        out1 => S1143
    );
nand_n_271: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selAC_MEM,
        in1(1) => U1_AC_out_4,
        out1 => S1144
    );
nand_n_272: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1144,
        in1(1) => S1143,
        out1 => U1_dataBus_out_4
    );
nand_n_273: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1976,
        in1(1) => S30,
        out1 => S1145
    );
nand_n_274: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_PC_out_5,
        in1(1) => S1975,
        out1 => S1146
    );
nand_n_275: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1146,
        in1(1) => S1145,
        out1 => S1147
    );
nand_n_276: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1147,
        in1(1) => U1_selPC_MEM,
        out1 => S1148
    );
nand_n_277: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_IN_out_5,
        in1(1) => S1996,
        out1 => S1149
    );
nand_n_278: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1149,
        in1(1) => S1148,
        out1 => S1150
    );
nand_n_279: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1150,
        in1(1) => S1997,
        out1 => S1151
    );
nand_n_280: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selAC_MEM,
        in1(1) => U1_AC_out_5,
        out1 => S1152
    );
nand_n_281: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1152,
        in1(1) => S1151,
        out1 => U1_dataBus_out_5
    );
nand_n_282: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1978,
        in1(1) => S31,
        out1 => S1153
    );
nand_n_283: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_PC_out_6,
        in1(1) => S1977,
        out1 => S1154
    );
nand_n_284: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1154,
        in1(1) => S1153,
        out1 => S1155
    );
nand_n_285: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1155,
        in1(1) => U1_selPC_MEM,
        out1 => S1156
    );
nand_n_286: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_IN_out_6,
        in1(1) => S1996,
        out1 => S1157
    );
nand_n_287: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1157,
        in1(1) => S1156,
        out1 => S1158
    );
nand_n_288: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1158,
        in1(1) => S1997,
        out1 => S1159
    );
nand_n_289: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selAC_MEM,
        in1(1) => U1_AC_out_6,
        out1 => S1160
    );
nand_n_290: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1160,
        in1(1) => S1159,
        out1 => U1_dataBus_out_6
    );
nand_n_291: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1980,
        in1(1) => S32,
        out1 => S1161
    );
nand_n_292: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_PC_out_7,
        in1(1) => S1979,
        out1 => S1162
    );
nand_n_293: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1162,
        in1(1) => S1161,
        out1 => S1163
    );
nand_n_294: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1163,
        in1(1) => U1_selPC_MEM,
        out1 => S1164
    );
nand_n_295: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_IN_out_7,
        in1(1) => S1996,
        out1 => S1165
    );
nand_n_296: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1165,
        in1(1) => S1164,
        out1 => S1166
    );
nand_n_297: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1166,
        in1(1) => S1997,
        out1 => S1167
    );
nand_n_298: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selAC_MEM,
        in1(1) => U1_AC_out_7,
        out1 => S1168
    );
nand_n_299: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1168,
        in1(1) => S1167,
        out1 => U1_dataBus_out_7
    );
nand_n_300: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1982,
        in1(1) => S33,
        out1 => S1169
    );
nand_n_301: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_PC_out_8,
        in1(1) => S1981,
        out1 => S1170
    );
nand_n_302: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1170,
        in1(1) => S1169,
        out1 => S1171
    );
nand_n_303: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1171,
        in1(1) => U1_selPC_MEM,
        out1 => S1172
    );
nand_n_304: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_IN_out_8,
        in1(1) => S1996,
        out1 => S1173
    );
nand_n_305: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1173,
        in1(1) => S1172,
        out1 => S1174
    );
nand_n_306: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1174,
        in1(1) => S1997,
        out1 => S1175
    );
nand_n_307: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selAC_MEM,
        in1(1) => U1_AC_out_8,
        out1 => S1176
    );
nand_n_308: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1176,
        in1(1) => S1175,
        out1 => U1_dataBus_out_8
    );
nand_n_309: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1984,
        in1(1) => S34,
        out1 => S1177
    );
nand_n_310: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_PC_out_9,
        in1(1) => S1983,
        out1 => S1178
    );
nand_n_311: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1178,
        in1(1) => S1177,
        out1 => S1179
    );
nand_n_312: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1179,
        in1(1) => U1_selPC_MEM,
        out1 => S1180
    );
nand_n_313: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_IN_out_9,
        in1(1) => S1996,
        out1 => S1181
    );
nand_n_314: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1181,
        in1(1) => S1180,
        out1 => S1182
    );
nand_n_315: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1182,
        in1(1) => S1997,
        out1 => S1183
    );
nand_n_316: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selAC_MEM,
        in1(1) => U1_AC_out_9,
        out1 => S1184
    );
nand_n_317: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1184,
        in1(1) => S1183,
        out1 => U1_dataBus_out_9
    );
nand_n_318: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1986,
        in1(1) => S35,
        out1 => S1185
    );
nand_n_319: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_PC_out_10,
        in1(1) => S1985,
        out1 => S1186
    );
nand_n_320: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1186,
        in1(1) => S1185,
        out1 => S1187
    );
nand_n_321: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1187,
        in1(1) => U1_selPC_MEM,
        out1 => S1188
    );
nand_n_322: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_IN_out_10,
        in1(1) => S1996,
        out1 => S1189
    );
nand_n_323: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1189,
        in1(1) => S1188,
        out1 => S1190
    );
nand_n_324: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1190,
        in1(1) => S1997,
        out1 => S1191
    );
nand_n_325: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selAC_MEM,
        in1(1) => U1_AC_out_10,
        out1 => S1192
    );
nand_n_326: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1192,
        in1(1) => S1191,
        out1 => U1_dataBus_out_10
    );
nand_n_327: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1988,
        in1(1) => S36,
        out1 => S1193
    );
nand_n_328: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_PC_out_11,
        in1(1) => S1987,
        out1 => S1194
    );
nand_n_329: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1194,
        in1(1) => S1193,
        out1 => S1195
    );
nand_n_330: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1195,
        in1(1) => U1_selPC_MEM,
        out1 => S1196
    );
nand_n_331: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_IN_out_11,
        in1(1) => S1996,
        out1 => S1197
    );
nand_n_332: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1197,
        in1(1) => S1196,
        out1 => S1198
    );
nand_n_333: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1198,
        in1(1) => S1997,
        out1 => S1199
    );
nand_n_334: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selAC_MEM,
        in1(1) => U1_AC_out_11,
        out1 => S1200
    );
nand_n_335: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1200,
        in1(1) => S1199,
        out1 => U1_dataBus_out_11
    );
nand_n_336: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1989,
        in1(1) => U1_PC_out_12,
        out1 => S1201
    );
nand_n_337: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S37,
        in1(1) => S1961,
        out1 => S1202
    );
nand_n_338: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1202,
        in1(1) => S1201,
        out1 => S1203
    );
nand_n_339: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1203,
        in1(1) => U1_selPC_MEM,
        out1 => S1204
    );
nand_n_340: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_IN_out_12,
        in1(1) => S1996,
        out1 => S1205
    );
nand_n_341: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1205,
        in1(1) => S1204,
        out1 => S1206
    );
nand_n_342: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1206,
        in1(1) => S1997,
        out1 => S1207
    );
nand_n_343: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selAC_MEM,
        in1(1) => U1_AC_out_12,
        out1 => S1208
    );
nand_n_344: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1208,
        in1(1) => S1207,
        out1 => U1_dataBus_out_12
    );
nand_n_345: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1990,
        in1(1) => U1_PC_out_13,
        out1 => S1209
    );
nand_n_346: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S38,
        in1(1) => S1963,
        out1 => S1210
    );
nand_n_347: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1210,
        in1(1) => S1209,
        out1 => S1211
    );
nand_n_348: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1211,
        in1(1) => U1_selPC_MEM,
        out1 => S1212
    );
nand_n_349: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_IN_out_13,
        in1(1) => S1996,
        out1 => S1213
    );
nand_n_350: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1213,
        in1(1) => S1212,
        out1 => S1214
    );
nand_n_351: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1214,
        in1(1) => S1997,
        out1 => S1215
    );
nand_n_352: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selAC_MEM,
        in1(1) => U1_AC_out_13,
        out1 => S1216
    );
nand_n_353: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1216,
        in1(1) => S1215,
        out1 => U1_dataBus_out_13
    );
nand_n_354: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1991,
        in1(1) => U1_PC_out_14,
        out1 => S1217
    );
nand_n_355: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S39,
        in1(1) => S1964,
        out1 => S1218
    );
nand_n_356: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1218,
        in1(1) => S1217,
        out1 => S1219
    );
nand_n_357: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1219,
        in1(1) => U1_selPC_MEM,
        out1 => S1220
    );
nand_n_358: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_IN_out_14,
        in1(1) => S1996,
        out1 => S1221
    );
nand_n_359: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1221,
        in1(1) => S1220,
        out1 => S1222
    );
nand_n_360: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1222,
        in1(1) => S1997,
        out1 => S1223
    );
nand_n_361: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selAC_MEM,
        in1(1) => U1_AC_out_14,
        out1 => S1224
    );
nand_n_362: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1224,
        in1(1) => S1223,
        out1 => U1_dataBus_out_14
    );
nor_n_148: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S40,
        in1(1) => U1_PC_out_15,
        out1 => S1225
    );
nand_n_363: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S40,
        in1(1) => U1_PC_out_15,
        out1 => S1226
    );
notg_21: ENTITY WORK.notg
    PORT MAP (
        in1 => S1226,
        out1 => S1227
    );
nor_n_149: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1227,
        in1(1) => S1225,
        out1 => S1228
    );
nand_n_364: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1228,
        in1(1) => U1_selPC_MEM,
        out1 => S1229
    );
nand_n_365: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_IN_out_15,
        in1(1) => S1996,
        out1 => S1230
    );
nand_n_366: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1230,
        in1(1) => S1229,
        out1 => S1231
    );
nand_n_367: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1231,
        in1(1) => S1997,
        out1 => S1232
    );
nand_n_368: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selAC_MEM,
        in1(1) => U1_AC_out_15,
        out1 => S1233
    );
nand_n_369: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1233,
        in1(1) => S1232,
        out1 => U1_dataBus_out_15
    );
nor_n_150: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2181,
        in1(1) => S1998,
        out1 => S1234
    );
nand_n_370: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1998,
        in1(1) => U1_IN_out_0,
        out1 => S1235
    );
nor_n_151: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1996,
        in1(1) => U1_PC_out_0,
        out1 => S1236
    );
nand_n_371: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1235,
        in1(1) => S1996,
        out1 => S1237
    );
nor_n_152: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1237,
        in1(1) => S1234,
        out1 => S1238
    );
nor_n_153: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1238,
        in1(1) => S1236,
        out1 => U1_addrBus_0
    );
nor_n_154: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2168,
        in1(1) => S1998,
        out1 => S1239
    );
nand_n_372: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1998,
        in1(1) => U1_IN_out_1,
        out1 => S1240
    );
nor_n_155: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1996,
        in1(1) => U1_PC_out_1,
        out1 => S1241
    );
nand_n_373: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1240,
        in1(1) => S1996,
        out1 => S1242
    );
nor_n_156: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1242,
        in1(1) => S1239,
        out1 => S1243
    );
nor_n_157: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1243,
        in1(1) => S1241,
        out1 => U1_addrBus_1
    );
nor_n_158: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2154,
        in1(1) => S1998,
        out1 => S1244
    );
nand_n_374: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1998,
        in1(1) => U1_IN_out_2,
        out1 => S1245
    );
nor_n_159: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1996,
        in1(1) => U1_PC_out_2,
        out1 => S1246
    );
nand_n_375: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1245,
        in1(1) => S1996,
        out1 => S1247
    );
nor_n_160: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1247,
        in1(1) => S1244,
        out1 => S1248
    );
nor_n_161: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1248,
        in1(1) => S1246,
        out1 => U1_addrBus_2
    );
nor_n_162: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2143,
        in1(1) => S1998,
        out1 => S1249
    );
nand_n_376: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1998,
        in1(1) => U1_IN_out_3,
        out1 => S1250
    );
nor_n_163: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1996,
        in1(1) => U1_PC_out_3,
        out1 => S1251
    );
nand_n_377: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1250,
        in1(1) => S1996,
        out1 => S1252
    );
nor_n_164: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1252,
        in1(1) => S1249,
        out1 => S1253
    );
nor_n_165: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1253,
        in1(1) => S1251,
        out1 => U1_addrBus_3
    );
nand_n_378: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2227,
        in1(1) => U1_selIR_MEM,
        out1 => S1254
    );
nand_n_379: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1998,
        in1(1) => U1_IN_out_4,
        out1 => S1255
    );
nand_n_380: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1255,
        in1(1) => S1254,
        out1 => S1256
    );
nand_n_381: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1256,
        in1(1) => S1996,
        out1 => S1257
    );
nand_n_382: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selPC_MEM,
        in1(1) => U1_PC_out_4,
        out1 => S1258
    );
nand_n_383: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1258,
        in1(1) => S1257,
        out1 => U1_addrBus_4
    );
nand_n_384: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2215,
        in1(1) => U1_selIR_MEM,
        out1 => S1259
    );
nand_n_385: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1998,
        in1(1) => U1_IN_out_5,
        out1 => S1260
    );
nand_n_386: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1260,
        in1(1) => S1259,
        out1 => S1261
    );
nand_n_387: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1261,
        in1(1) => S1996,
        out1 => S1262
    );
nand_n_388: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selPC_MEM,
        in1(1) => U1_PC_out_5,
        out1 => S1263
    );
nand_n_389: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1263,
        in1(1) => S1262,
        out1 => U1_addrBus_5
    );
nand_n_390: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2204,
        in1(1) => U1_selIR_MEM,
        out1 => S1264
    );
nand_n_391: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1998,
        in1(1) => U1_IN_out_6,
        out1 => S1265
    );
nand_n_392: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1265,
        in1(1) => S1264,
        out1 => S1266
    );
nand_n_393: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1266,
        in1(1) => S1996,
        out1 => S1267
    );
nand_n_394: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selPC_MEM,
        in1(1) => U1_PC_out_6,
        out1 => S1268
    );
nand_n_395: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1268,
        in1(1) => S1267,
        out1 => U1_addrBus_6
    );
nand_n_396: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2195,
        in1(1) => U1_selIR_MEM,
        out1 => S1269
    );
nand_n_397: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1998,
        in1(1) => U1_IN_out_7,
        out1 => S1270
    );
nand_n_398: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1270,
        in1(1) => S1269,
        out1 => S1271
    );
nand_n_399: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1271,
        in1(1) => S1996,
        out1 => S1272
    );
nand_n_400: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selPC_MEM,
        in1(1) => U1_PC_out_7,
        out1 => S1273
    );
nand_n_401: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1273,
        in1(1) => S1272,
        out1 => U1_addrBus_7
    );
nand_n_402: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2079,
        in1(1) => U1_selIR_MEM,
        out1 => S1274
    );
nand_n_403: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1998,
        in1(1) => U1_IN_out_8,
        out1 => S1275
    );
nand_n_404: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1275,
        in1(1) => S1274,
        out1 => S1276
    );
nand_n_405: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1276,
        in1(1) => S1996,
        out1 => S1277
    );
nand_n_406: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selPC_MEM,
        in1(1) => U1_PC_out_8,
        out1 => S1278
    );
nand_n_407: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1278,
        in1(1) => S1277,
        out1 => U1_addrBus_8
    );
nand_n_408: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2070,
        in1(1) => U1_selIR_MEM,
        out1 => S1279
    );
nand_n_409: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1998,
        in1(1) => U1_IN_out_9,
        out1 => S1280
    );
nand_n_410: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1280,
        in1(1) => S1279,
        out1 => S1281
    );
nand_n_411: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1281,
        in1(1) => S1996,
        out1 => S1282
    );
nand_n_412: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selPC_MEM,
        in1(1) => U1_PC_out_9,
        out1 => S1283
    );
nand_n_413: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1283,
        in1(1) => S1282,
        out1 => U1_addrBus_9
    );
nand_n_414: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2058,
        in1(1) => U1_selIR_MEM,
        out1 => S1284
    );
nand_n_415: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1998,
        in1(1) => U1_IN_out_10,
        out1 => S1285
    );
nand_n_416: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1285,
        in1(1) => S1284,
        out1 => S1286
    );
nand_n_417: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1286,
        in1(1) => S1996,
        out1 => S1287
    );
nand_n_418: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selPC_MEM,
        in1(1) => U1_PC_out_10,
        out1 => S1288
    );
nand_n_419: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1288,
        in1(1) => S1287,
        out1 => U1_addrBus_10
    );
nand_n_420: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2050,
        in1(1) => U1_selIR_MEM,
        out1 => S1289
    );
nand_n_421: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1998,
        in1(1) => U1_IN_out_11,
        out1 => S1290
    );
nand_n_422: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1290,
        in1(1) => S1289,
        out1 => S1291
    );
nand_n_423: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1291,
        in1(1) => S1996,
        out1 => S1292
    );
nand_n_424: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selPC_MEM,
        in1(1) => U1_PC_out_11,
        out1 => S1293
    );
nand_n_425: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1293,
        in1(1) => S1292,
        out1 => U1_addrBus_11
    );
nand_n_426: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2122,
        in1(1) => U1_selIR_MEM,
        out1 => S1294
    );
nand_n_427: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1998,
        in1(1) => U1_IN_out_12,
        out1 => S1295
    );
nand_n_428: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1295,
        in1(1) => S1294,
        out1 => S1296
    );
nand_n_429: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1296,
        in1(1) => S1996,
        out1 => S1297
    );
nand_n_430: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selPC_MEM,
        in1(1) => U1_PC_out_12,
        out1 => S1298
    );
nand_n_431: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1298,
        in1(1) => S1297,
        out1 => U1_addrBus_12
    );
nand_n_432: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2113,
        in1(1) => U1_selIR_MEM,
        out1 => S1299
    );
nand_n_433: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1998,
        in1(1) => U1_IN_out_13,
        out1 => S1300
    );
nand_n_434: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1300,
        in1(1) => S1299,
        out1 => S1301
    );
nand_n_435: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1301,
        in1(1) => S1996,
        out1 => S1302
    );
nand_n_436: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selPC_MEM,
        in1(1) => U1_PC_out_13,
        out1 => S1303
    );
nand_n_437: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1303,
        in1(1) => S1302,
        out1 => U1_addrBus_13
    );
nand_n_438: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2103,
        in1(1) => U1_selIR_MEM,
        out1 => S1304
    );
nand_n_439: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1998,
        in1(1) => U1_IN_out_14,
        out1 => S1305
    );
nand_n_440: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1305,
        in1(1) => S1304,
        out1 => S1306
    );
nand_n_441: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1306,
        in1(1) => S1996,
        out1 => S1307
    );
nand_n_442: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selPC_MEM,
        in1(1) => U1_PC_out_14,
        out1 => S1308
    );
nand_n_443: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1308,
        in1(1) => S1307,
        out1 => U1_addrBus_14
    );
nand_n_444: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2020,
        in1(1) => U1_selIR_MEM,
        out1 => S1309
    );
nand_n_445: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1998,
        in1(1) => U1_IN_out_15,
        out1 => S1310
    );
nand_n_446: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1310,
        in1(1) => S1309,
        out1 => S1311
    );
nand_n_447: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1311,
        in1(1) => S1996,
        out1 => S1312
    );
nand_n_448: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selPC_MEM,
        in1(1) => U1_PC_out_15,
        out1 => S1313
    );
nand_n_449: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1313,
        in1(1) => S1312,
        out1 => U1_addrBus_15
    );
nor_n_166: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_V_out1,
        in1(1) => U1_IR_out_0,
        out1 => S1314
    );
notg_22: ENTITY WORK.notg
    PORT MAP (
        in1 => S1314,
        out1 => S1315
    );
nand_n_450: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_V_out1,
        in1(1) => U1_IR_out_0,
        out1 => S1316
    );
nand_n_451: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1316,
        in1(1) => S1315,
        out1 => S1317
    );
nor_n_167: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_C_out1,
        in1(1) => U1_IR_out_1,
        out1 => S1318
    );
notg_23: ENTITY WORK.notg
    PORT MAP (
        in1 => S1318,
        out1 => S1319
    );
nand_n_452: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_C_out1,
        in1(1) => U1_IR_out_1,
        out1 => S1320
    );
nand_n_453: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1320,
        in1(1) => S1319,
        out1 => S1321
    );
nor_n_168: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1321,
        in1(1) => S1317,
        out1 => S1322
    );
nor_n_169: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_N_out1,
        in1(1) => U1_IR_out_2,
        out1 => S1323
    );
notg_24: ENTITY WORK.notg
    PORT MAP (
        in1 => S1323,
        out1 => S1324
    );
nand_n_454: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_N_out1,
        in1(1) => U1_IR_out_2,
        out1 => S1325
    );
nand_n_455: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1325,
        in1(1) => S1324,
        out1 => S1326
    );
nor_n_170: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_Z_out1,
        in1(1) => U1_IR_out_3,
        out1 => S1327
    );
notg_25: ENTITY WORK.notg
    PORT MAP (
        in1 => S1327,
        out1 => S1328
    );
nand_n_456: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_Z_out1,
        in1(1) => U1_IR_out_3,
        out1 => S1329
    );
nand_n_457: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1329,
        in1(1) => S1328,
        out1 => S1330
    );
nor_n_171: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1330,
        in1(1) => S1326,
        out1 => S1331
    );
nand_n_458: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1331,
        in1(1) => S1322,
        out1 => U1_enSKP
    );
nor_n_172: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2181,
        in1(1) => S1962,
        out1 => S1332
    );
nand_n_459: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1962,
        in1(1) => U1_PC_out_12,
        out1 => S1333
    );
nor_n_173: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_ldOF,
        in1(1) => U1_OF_out_0,
        out1 => S1334
    );
nand_n_460: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1333,
        in1(1) => U1_ldOF,
        out1 => S1335
    );
nor_n_174: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1335,
        in1(1) => S1332,
        out1 => S1336
    );
nor_n_175: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1336,
        in1(1) => S1334,
        out1 => S70
    );
nor_n_176: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2168,
        in1(1) => S1962,
        out1 => S1337
    );
nand_n_461: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_PC_out_13,
        in1(1) => S1962,
        out1 => S1338
    );
nor_n_177: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_ldOF,
        in1(1) => U1_OF_out_1,
        out1 => S1339
    );
nand_n_462: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1338,
        in1(1) => U1_ldOF,
        out1 => S1340
    );
nor_n_178: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1340,
        in1(1) => S1337,
        out1 => S1341
    );
nor_n_179: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1341,
        in1(1) => S1339,
        out1 => S71
    );
nor_n_180: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2154,
        in1(1) => S1962,
        out1 => S1342
    );
nand_n_463: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_PC_out_14,
        in1(1) => S1962,
        out1 => S1343
    );
nor_n_181: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_ldOF,
        in1(1) => U1_OF_out_2,
        out1 => S1344
    );
nand_n_464: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1343,
        in1(1) => U1_ldOF,
        out1 => S1345
    );
nor_n_182: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1345,
        in1(1) => S1342,
        out1 => S1346
    );
nor_n_183: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1346,
        in1(1) => S1344,
        out1 => S72
    );
nor_n_184: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2143,
        in1(1) => S1962,
        out1 => S1347
    );
nand_n_465: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_PC_out_15,
        in1(1) => S1962,
        out1 => S1348
    );
nor_n_185: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_ldOF,
        in1(1) => U1_OF_out_3,
        out1 => S1349
    );
nand_n_466: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1348,
        in1(1) => U1_ldOF,
        out1 => S1350
    );
nor_n_186: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1350,
        in1(1) => S1347,
        out1 => S1351
    );
nor_n_187: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1351,
        in1(1) => S1349,
        out1 => S73
    );
nor_n_188: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_ldAC,
        in1(1) => U1_zeroAC,
        out1 => S1352
    );
nand_n_467: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1352,
        in1(1) => U1_AC_out_0,
        out1 => S1353
    );
nand_n_468: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2180,
        in1(1) => S1999,
        out1 => S1354
    );
nand_n_469: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selMEM_AC,
        in1(1) => U1_dataBus_0,
        out1 => S1355
    );
nand_n_470: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1355,
        in1(1) => S1354,
        out1 => S1356
    );
nand_n_471: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1356,
        in1(1) => S2000,
        out1 => S1357
    );
nor_n_189: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2518,
        in1(1) => U1_AC_out_0,
        out1 => S1358
    );
nor_n_190: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1358,
        in1(1) => S653,
        out1 => S1359
    );
nand_n_472: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1359,
        in1(1) => U1_ADD,
        out1 => S1360
    );
nand_n_473: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S653,
        in1(1) => S597,
        out1 => S1361
    );
nand_n_474: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1361,
        in1(1) => S1360,
        out1 => S1362
    );
nand_n_475: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1362,
        in1(1) => U1_selARU_AC,
        out1 => S1363
    );
nand_n_476: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1363,
        in1(1) => S1357,
        out1 => S1364
    );
nand_n_477: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S862,
        in1(1) => U1_selLGU_AC,
        out1 => S1365
    );
nor_n_191: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1364,
        in1(1) => U1_selLGU_AC,
        out1 => S1366
    );
nor_n_192: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1366,
        in1(1) => S1960,
        out1 => S1367
    );
nand_n_478: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1367,
        in1(1) => S1365,
        out1 => S1368
    );
nand_n_479: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1368,
        in1(1) => S1353,
        out1 => S74
    );
nand_n_480: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1352,
        in1(1) => U1_AC_out_1,
        out1 => S1369
    );
nand_n_481: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1058,
        in1(1) => U1_selLGU_AC,
        out1 => S1370
    );
nor_n_193: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2168,
        in1(1) => U1_selMEM_AC,
        out1 => S1371
    );
nand_n_482: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selMEM_AC,
        in1(1) => U1_dataBus_1,
        out1 => S1372
    );
nand_n_483: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1372,
        in1(1) => S2000,
        out1 => S1373
    );
nor_n_194: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1373,
        in1(1) => S1371,
        out1 => S1374
    );
nor_n_195: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S655,
        in1(1) => S653,
        out1 => S1375
    );
nand_n_484: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S656,
        in1(1) => U1_ADD,
        out1 => S1376
    );
nor_n_196: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1376,
        in1(1) => S1375,
        out1 => S1377
    );
nor_n_197: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2517,
        in1(1) => S1925,
        out1 => S1378
    );
nor_n_198: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1378,
        in1(1) => S500,
        out1 => S1379
    );
nor_n_199: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1379,
        in1(1) => S598,
        out1 => S1380
    );
nand_n_485: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1380,
        in1(1) => S525,
        out1 => S1381
    );
nand_n_486: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1381,
        in1(1) => U1_selARU_AC,
        out1 => S1382
    );
nor_n_200: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1382,
        in1(1) => S1377,
        out1 => S1383
    );
nor_n_201: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1383,
        in1(1) => S1374,
        out1 => S1384
    );
nor_n_202: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1384,
        in1(1) => U1_selLGU_AC,
        out1 => S1385
    );
nor_n_203: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1385,
        in1(1) => S1960,
        out1 => S1386
    );
nand_n_487: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1386,
        in1(1) => S1370,
        out1 => S1387
    );
nand_n_488: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1387,
        in1(1) => S1369,
        out1 => S75
    );
nand_n_489: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1352,
        in1(1) => U1_AC_out_2,
        out1 => S1388
    );
nand_n_490: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1036,
        in1(1) => U1_selLGU_AC,
        out1 => S1389
    );
nor_n_204: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2154,
        in1(1) => U1_selMEM_AC,
        out1 => S1390
    );
nand_n_491: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selMEM_AC,
        in1(1) => U1_dataBus_2,
        out1 => S1391
    );
nand_n_492: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1391,
        in1(1) => S2000,
        out1 => S1392
    );
nor_n_205: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1392,
        in1(1) => S1390,
        out1 => S1393
    );
nand_n_493: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S527,
        in1(1) => S525,
        out1 => S1394
    );
nand_n_494: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1394,
        in1(1) => S597,
        out1 => S1395
    );
nor_n_206: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1395,
        in1(1) => S528,
        out1 => S1396
    );
nor_n_207: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S657,
        in1(1) => S652,
        out1 => S1397
    );
nor_n_208: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1397,
        in1(1) => S1995,
        out1 => S1398
    );
nand_n_495: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1398,
        in1(1) => S658,
        out1 => S1399
    );
nand_n_496: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1399,
        in1(1) => U1_selARU_AC,
        out1 => S1400
    );
nor_n_209: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1400,
        in1(1) => S1396,
        out1 => S1401
    );
nor_n_210: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1401,
        in1(1) => S1393,
        out1 => S1402
    );
nor_n_211: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1402,
        in1(1) => U1_selLGU_AC,
        out1 => S1403
    );
nor_n_212: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1403,
        in1(1) => S1960,
        out1 => S1404
    );
nand_n_497: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1404,
        in1(1) => S1389,
        out1 => S1405
    );
nand_n_498: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1405,
        in1(1) => S1388,
        out1 => S76
    );
nand_n_499: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1352,
        in1(1) => U1_AC_out_3,
        out1 => S1406
    );
nor_n_213: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S531,
        in1(1) => S528,
        out1 => S1407
    );
notg_26: ENTITY WORK.notg
    PORT MAP (
        in1 => S1407,
        out1 => S1408
    );
nand_n_500: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1408,
        in1(1) => U1_MUL,
        out1 => S1409
    );
nor_n_214: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1409,
        in1(1) => S533,
        out1 => S1410
    );
nor_n_215: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1410,
        in1(1) => U1_ADD,
        out1 => S1411
    );
nand_n_501: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S650,
        in1(1) => S2615,
        out1 => S1412
    );
nand_n_502: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1412,
        in1(1) => S659,
        out1 => S1413
    );
nor_n_216: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1412,
        in1(1) => S659,
        out1 => S1414
    );
nor_n_217: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1414,
        in1(1) => S1995,
        out1 => S1415
    );
nand_n_503: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1415,
        in1(1) => S1413,
        out1 => S1416
    );
nand_n_504: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1416,
        in1(1) => U1_selARU_AC,
        out1 => S1417
    );
nor_n_218: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1417,
        in1(1) => S1411,
        out1 => S1418
    );
nand_n_505: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2143,
        in1(1) => S1999,
        out1 => S1419
    );
nor_n_219: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1999,
        in1(1) => U1_dataBus_3,
        out1 => S1420
    );
nor_n_220: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1420,
        in1(1) => U1_selARU_AC,
        out1 => S1421
    );
nand_n_506: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1421,
        in1(1) => S1419,
        out1 => S1422
    );
nand_n_507: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1422,
        in1(1) => S2001,
        out1 => S1423
    );
nor_n_221: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1423,
        in1(1) => S1418,
        out1 => S1424
    );
nand_n_508: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S896,
        in1(1) => U1_selLGU_AC,
        out1 => S1425
    );
nor_n_222: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1424,
        in1(1) => S1960,
        out1 => S1426
    );
nand_n_509: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1426,
        in1(1) => S1425,
        out1 => S1427
    );
nand_n_510: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1427,
        in1(1) => S1406,
        out1 => S77
    );
nand_n_511: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1352,
        in1(1) => U1_AC_out_4,
        out1 => S1428
    );
nor_n_223: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2226,
        in1(1) => U1_selMEM_AC,
        out1 => S1429
    );
nand_n_512: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selMEM_AC,
        in1(1) => U1_dataBus_4,
        out1 => S1430
    );
nand_n_513: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1430,
        in1(1) => S2000,
        out1 => S1431
    );
nor_n_224: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1431,
        in1(1) => S1429,
        out1 => S1432
    );
nor_n_225: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S535,
        in1(1) => S533,
        out1 => S1433
    );
nand_n_514: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S597,
        in1(1) => S536,
        out1 => S1434
    );
nor_n_226: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1434,
        in1(1) => S1433,
        out1 => S1435
    );
nor_n_227: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S661,
        in1(1) => S649,
        out1 => S1436
    );
nor_n_228: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1436,
        in1(1) => S663,
        out1 => S1437
    );
nand_n_515: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1437,
        in1(1) => U1_ADD,
        out1 => S1438
    );
nand_n_516: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1438,
        in1(1) => U1_selARU_AC,
        out1 => S1439
    );
nor_n_229: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1439,
        in1(1) => S1435,
        out1 => S1440
    );
nor_n_230: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1440,
        in1(1) => S1432,
        out1 => S1441
    );
nor_n_231: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1441,
        in1(1) => U1_selLGU_AC,
        out1 => S1442
    );
nand_n_517: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S966,
        in1(1) => U1_selLGU_AC,
        out1 => S1443
    );
nor_n_232: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1442,
        in1(1) => S1960,
        out1 => S1444
    );
nand_n_518: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1444,
        in1(1) => S1443,
        out1 => S1445
    );
nand_n_519: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1445,
        in1(1) => S1428,
        out1 => S78
    );
nand_n_520: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1352,
        in1(1) => U1_AC_out_5,
        out1 => S1446
    );
nand_n_521: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2215,
        in1(1) => S1999,
        out1 => S1447
    );
nand_n_522: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selMEM_AC,
        in1(1) => U1_dataBus_5,
        out1 => S1448
    );
nand_n_523: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1448,
        in1(1) => S1447,
        out1 => S1449
    );
nor_n_233: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1449,
        in1(1) => U1_selARU_AC,
        out1 => S1450
    );
nand_n_524: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S543,
        in1(1) => S538,
        out1 => S1451
    );
nor_n_234: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S598,
        in1(1) => S544,
        out1 => S1452
    );
nand_n_525: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1452,
        in1(1) => S1451,
        out1 => S1453
    );
nor_n_235: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S664,
        in1(1) => S647,
        out1 => S1454
    );
nand_n_526: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S665,
        in1(1) => U1_ADD,
        out1 => S1455
    );
nor_n_236: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1455,
        in1(1) => S1454,
        out1 => S1456
    );
nand_n_527: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1453,
        in1(1) => U1_selARU_AC,
        out1 => S1457
    );
nor_n_237: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1457,
        in1(1) => S1456,
        out1 => S1458
    );
nor_n_238: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1458,
        in1(1) => S1450,
        out1 => S1459
    );
nor_n_239: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1459,
        in1(1) => U1_selLGU_AC,
        out1 => S1460
    );
nand_n_528: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1086,
        in1(1) => U1_selLGU_AC,
        out1 => S1461
    );
nor_n_240: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1460,
        in1(1) => S1960,
        out1 => S1462
    );
nand_n_529: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1462,
        in1(1) => S1461,
        out1 => S1463
    );
nand_n_530: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1463,
        in1(1) => S1446,
        out1 => S79
    );
nand_n_531: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1352,
        in1(1) => U1_AC_out_6,
        out1 => S1464
    );
nand_n_532: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2204,
        in1(1) => S1999,
        out1 => S1465
    );
nand_n_533: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selMEM_AC,
        in1(1) => U1_dataBus_6,
        out1 => S1466
    );
nand_n_534: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1466,
        in1(1) => S1465,
        out1 => S1467
    );
nor_n_241: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1467,
        in1(1) => U1_selARU_AC,
        out1 => S1468
    );
nand_n_535: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S546,
        in1(1) => S456,
        out1 => S1469
    );
nand_n_536: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1469,
        in1(1) => S597,
        out1 => S1470
    );
nor_n_242: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1470,
        in1(1) => S548,
        out1 => S1471
    );
nor_n_243: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S666,
        in1(1) => S645,
        out1 => S1472
    );
nor_n_244: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1472,
        in1(1) => S1995,
        out1 => S1473
    );
nand_n_537: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1473,
        in1(1) => S667,
        out1 => S1474
    );
nand_n_538: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1474,
        in1(1) => U1_selARU_AC,
        out1 => S1475
    );
nor_n_245: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1475,
        in1(1) => S1471,
        out1 => S1476
    );
nor_n_246: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1476,
        in1(1) => S1468,
        out1 => S1477
    );
nor_n_247: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1477,
        in1(1) => U1_selLGU_AC,
        out1 => S1478
    );
nand_n_539: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1020,
        in1(1) => U1_selLGU_AC,
        out1 => S1479
    );
nor_n_248: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1478,
        in1(1) => S1960,
        out1 => S1480
    );
nand_n_540: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1480,
        in1(1) => S1479,
        out1 => S1481
    );
nand_n_541: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1481,
        in1(1) => S1464,
        out1 => S80
    );
nand_n_542: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1352,
        in1(1) => U1_AC_out_7,
        out1 => S1482
    );
nand_n_543: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2195,
        in1(1) => S1999,
        out1 => S1483
    );
nand_n_544: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selMEM_AC,
        in1(1) => U1_dataBus_7,
        out1 => S1484
    );
nand_n_545: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1484,
        in1(1) => S1483,
        out1 => S1485
    );
nor_n_249: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1485,
        in1(1) => U1_selARU_AC,
        out1 => S1486
    );
nand_n_546: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S550,
        in1(1) => S405,
        out1 => S1487
    );
nor_n_250: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S598,
        in1(1) => S552,
        out1 => S1488
    );
nand_n_547: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1488,
        in1(1) => S1487,
        out1 => S1489
    );
notg_27: ENTITY WORK.notg
    PORT MAP (
        in1 => S1489,
        out1 => S1490
    );
nor_n_251: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S643,
        in1(1) => S2419,
        out1 => S1491
    );
nor_n_252: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1491,
        in1(1) => S668,
        out1 => S1492
    );
nand_n_548: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1491,
        in1(1) => S668,
        out1 => S1493
    );
nor_n_253: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1492,
        in1(1) => S1995,
        out1 => S1494
    );
nand_n_549: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1494,
        in1(1) => S1493,
        out1 => S1495
    );
nand_n_550: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1495,
        in1(1) => U1_selARU_AC,
        out1 => S1496
    );
nor_n_254: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1496,
        in1(1) => S1490,
        out1 => S1497
    );
nor_n_255: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1497,
        in1(1) => S1486,
        out1 => S1498
    );
nor_n_256: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1498,
        in1(1) => U1_selLGU_AC,
        out1 => S1499
    );
nand_n_551: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1072,
        in1(1) => U1_selLGU_AC,
        out1 => S1500
    );
nor_n_257: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1499,
        in1(1) => S1960,
        out1 => S1501
    );
nand_n_552: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1501,
        in1(1) => S1500,
        out1 => S1502
    );
nand_n_553: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1502,
        in1(1) => S1482,
        out1 => S81
    );
nand_n_554: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1352,
        in1(1) => U1_AC_out_8,
        out1 => S1503
    );
nand_n_555: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2079,
        in1(1) => S1999,
        out1 => S1504
    );
nand_n_556: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selMEM_AC,
        in1(1) => U1_dataBus_8,
        out1 => S1505
    );
nand_n_557: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1505,
        in1(1) => S1504,
        out1 => S1506
    );
nor_n_258: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1506,
        in1(1) => U1_selARU_AC,
        out1 => S1507
    );
nor_n_259: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S555,
        in1(1) => S342,
        out1 => S1508
    );
nand_n_558: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S597,
        in1(1) => S557,
        out1 => S1509
    );
nor_n_260: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1509,
        in1(1) => S1508,
        out1 => S1510
    );
nor_n_261: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S670,
        in1(1) => S642,
        out1 => S1511
    );
nor_n_262: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1511,
        in1(1) => S1995,
        out1 => S1512
    );
nand_n_559: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1512,
        in1(1) => S671,
        out1 => S1513
    );
nand_n_560: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1513,
        in1(1) => U1_selARU_AC,
        out1 => S1514
    );
nor_n_263: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1514,
        in1(1) => S1510,
        out1 => S1515
    );
nor_n_264: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1515,
        in1(1) => S1507,
        out1 => S1516
    );
nor_n_265: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1516,
        in1(1) => U1_selLGU_AC,
        out1 => S1517
    );
nand_n_561: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S835,
        in1(1) => U1_selLGU_AC,
        out1 => S1518
    );
nor_n_266: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1517,
        in1(1) => S1960,
        out1 => S1519
    );
nand_n_562: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1519,
        in1(1) => S1518,
        out1 => S1520
    );
nand_n_563: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1520,
        in1(1) => S1503,
        out1 => S82
    );
nand_n_564: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1352,
        in1(1) => U1_AC_out_9,
        out1 => S1521
    );
nand_n_565: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2070,
        in1(1) => S1999,
        out1 => S1522
    );
nand_n_566: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selMEM_AC,
        in1(1) => U1_dataBus_9,
        out1 => S1523
    );
nand_n_567: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1523,
        in1(1) => S1522,
        out1 => S1524
    );
nor_n_267: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1524,
        in1(1) => U1_selARU_AC,
        out1 => S1525
    );
nand_n_568: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S558,
        in1(1) => S270,
        out1 => S1526
    );
nand_n_569: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1526,
        in1(1) => S561,
        out1 => S1527
    );
nor_n_268: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1527,
        in1(1) => S598,
        out1 => S1528
    );
nor_n_269: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S635,
        in1(1) => S633,
        out1 => S1529
    );
nor_n_270: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1529,
        in1(1) => S672,
        out1 => S1530
    );
nand_n_570: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1529,
        in1(1) => S672,
        out1 => S1531
    );
nor_n_271: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1530,
        in1(1) => S1995,
        out1 => S1532
    );
nand_n_571: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1532,
        in1(1) => S1531,
        out1 => S1533
    );
nand_n_572: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1533,
        in1(1) => U1_selARU_AC,
        out1 => S1534
    );
nor_n_272: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1534,
        in1(1) => S1528,
        out1 => S1535
    );
nor_n_273: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1535,
        in1(1) => S1525,
        out1 => S1536
    );
nor_n_274: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1536,
        in1(1) => U1_selLGU_AC,
        out1 => S1537
    );
nand_n_573: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1003,
        in1(1) => U1_selLGU_AC,
        out1 => S1538
    );
nor_n_275: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1537,
        in1(1) => S1960,
        out1 => S1539
    );
nand_n_574: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1539,
        in1(1) => S1538,
        out1 => S1540
    );
nand_n_575: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1540,
        in1(1) => S1521,
        out1 => S83
    );
nand_n_576: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1352,
        in1(1) => U1_AC_out_10,
        out1 => S1541
    );
nand_n_577: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2058,
        in1(1) => S1999,
        out1 => S1542
    );
nand_n_578: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selMEM_AC,
        in1(1) => U1_dataBus_10,
        out1 => S1543
    );
nand_n_579: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1543,
        in1(1) => S1542,
        out1 => S1544
    );
nor_n_276: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1544,
        in1(1) => U1_selARU_AC,
        out1 => S1545
    );
nor_n_277: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S563,
        in1(1) => S193,
        out1 => S1546
    );
nor_n_278: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1546,
        in1(1) => S564,
        out1 => S1547
    );
nand_n_580: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1547,
        in1(1) => S597,
        out1 => S1548
    );
notg_28: ENTITY WORK.notg
    PORT MAP (
        in1 => S1548,
        out1 => S1549
    );
nand_n_581: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S675,
        in1(1) => S630,
        out1 => S1550
    );
nor_n_279: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S676,
        in1(1) => S1995,
        out1 => S1551
    );
nand_n_582: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1551,
        in1(1) => S1550,
        out1 => S1552
    );
nand_n_583: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1552,
        in1(1) => U1_selARU_AC,
        out1 => S1553
    );
nor_n_280: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1553,
        in1(1) => S1549,
        out1 => S1554
    );
nor_n_281: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1554,
        in1(1) => S1545,
        out1 => S1555
    );
nor_n_282: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1555,
        in1(1) => U1_selLGU_AC,
        out1 => S1556
    );
nand_n_584: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S800,
        in1(1) => U1_selLGU_AC,
        out1 => S1557
    );
nor_n_283: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1556,
        in1(1) => S1960,
        out1 => S1558
    );
nand_n_585: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1558,
        in1(1) => S1557,
        out1 => S1559
    );
nand_n_586: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1559,
        in1(1) => S1541,
        out1 => S84
    );
nand_n_587: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1352,
        in1(1) => U1_AC_out_11,
        out1 => S1560
    );
nand_n_588: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2050,
        in1(1) => S1999,
        out1 => S1561
    );
nand_n_589: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selMEM_AC,
        in1(1) => U1_dataBus_11,
        out1 => S1562
    );
nand_n_590: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1562,
        in1(1) => S1561,
        out1 => S1563
    );
nor_n_284: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1563,
        in1(1) => U1_selARU_AC,
        out1 => S1564
    );
nor_n_285: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S567,
        in1(1) => S2595,
        out1 => S1565
    );
nand_n_591: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S597,
        in1(1) => S569,
        out1 => S1566
    );
nor_n_286: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1566,
        in1(1) => S1565,
        out1 => S1567
    );
nor_n_287: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S624,
        in1(1) => S622,
        out1 => S1568
    );
nor_n_288: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1568,
        in1(1) => S678,
        out1 => S1569
    );
nand_n_592: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1568,
        in1(1) => S678,
        out1 => S1570
    );
nor_n_289: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1569,
        in1(1) => S1995,
        out1 => S1571
    );
nand_n_593: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1571,
        in1(1) => S1570,
        out1 => S1572
    );
nand_n_594: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1572,
        in1(1) => U1_selARU_AC,
        out1 => S1573
    );
nor_n_290: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1573,
        in1(1) => S1567,
        out1 => S1574
    );
nor_n_291: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1574,
        in1(1) => S1564,
        out1 => S1575
    );
nor_n_292: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1575,
        in1(1) => U1_selLGU_AC,
        out1 => S1576
    );
nand_n_595: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S980,
        in1(1) => U1_selLGU_AC,
        out1 => S1577
    );
nor_n_293: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1576,
        in1(1) => S1960,
        out1 => S1578
    );
nand_n_596: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1578,
        in1(1) => S1577,
        out1 => S1579
    );
nand_n_597: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1579,
        in1(1) => S1560,
        out1 => S85
    );
nand_n_598: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1352,
        in1(1) => U1_AC_out_12,
        out1 => S1580
    );
nand_n_599: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2122,
        in1(1) => S1999,
        out1 => S1581
    );
nand_n_600: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selMEM_AC,
        in1(1) => U1_dataBus_12,
        out1 => S1582
    );
nand_n_601: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1582,
        in1(1) => S1581,
        out1 => S1583
    );
nor_n_294: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1583,
        in1(1) => U1_selARU_AC,
        out1 => S1584
    );
nand_n_602: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S570,
        in1(1) => S2515,
        out1 => S1585
    );
nor_n_295: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S598,
        in1(1) => S572,
        out1 => S1586
    );
nand_n_603: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1586,
        in1(1) => S1585,
        out1 => S1587
    );
nor_n_296: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S680,
        in1(1) => S619,
        out1 => S1588
    );
nand_n_604: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S681,
        in1(1) => U1_ADD,
        out1 => S1589
    );
nor_n_297: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1589,
        in1(1) => S1588,
        out1 => S1590
    );
nand_n_605: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1587,
        in1(1) => U1_selARU_AC,
        out1 => S1591
    );
nor_n_298: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1591,
        in1(1) => S1590,
        out1 => S1592
    );
nor_n_299: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1592,
        in1(1) => S1584,
        out1 => S1593
    );
nor_n_300: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1593,
        in1(1) => U1_selLGU_AC,
        out1 => S1594
    );
nand_n_606: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S952,
        in1(1) => U1_selLGU_AC,
        out1 => S1595
    );
nor_n_301: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1594,
        in1(1) => S1960,
        out1 => S1596
    );
nand_n_607: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1596,
        in1(1) => S1595,
        out1 => S1597
    );
nand_n_608: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1597,
        in1(1) => S1580,
        out1 => S86
    );
nand_n_609: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1352,
        in1(1) => U1_AC_out_13,
        out1 => S1598
    );
nand_n_610: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2113,
        in1(1) => S1999,
        out1 => S1599
    );
nand_n_611: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selMEM_AC,
        in1(1) => U1_dataBus_13,
        out1 => S1600
    );
nand_n_612: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1600,
        in1(1) => S1599,
        out1 => S1601
    );
nor_n_302: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1601,
        in1(1) => U1_selARU_AC,
        out1 => S1602
    );
nor_n_303: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S575,
        in1(1) => S2438,
        out1 => S1603
    );
nand_n_613: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S597,
        in1(1) => S577,
        out1 => S1604
    );
nor_n_304: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1604,
        in1(1) => S1603,
        out1 => S1605
    );
nor_n_305: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S612,
        in1(1) => S611,
        out1 => S1606
    );
nand_n_614: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1606,
        in1(1) => S682,
        out1 => S1607
    );
nor_n_306: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1606,
        in1(1) => S682,
        out1 => S1608
    );
nor_n_307: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1608,
        in1(1) => S1995,
        out1 => S1609
    );
nand_n_615: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1609,
        in1(1) => S1607,
        out1 => S1610
    );
nand_n_616: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1610,
        in1(1) => U1_selARU_AC,
        out1 => S1611
    );
nor_n_308: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1611,
        in1(1) => S1605,
        out1 => S1612
    );
nor_n_309: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1612,
        in1(1) => S1602,
        out1 => S1613
    );
nor_n_310: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1613,
        in1(1) => U1_selLGU_AC,
        out1 => S1614
    );
nand_n_617: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S930,
        in1(1) => U1_selLGU_AC,
        out1 => S1615
    );
nor_n_311: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1614,
        in1(1) => S1960,
        out1 => S1616
    );
nand_n_618: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1616,
        in1(1) => S1615,
        out1 => S1617
    );
nand_n_619: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1617,
        in1(1) => S1598,
        out1 => S87
    );
nand_n_620: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1352,
        in1(1) => U1_AC_out_14,
        out1 => S1618
    );
nand_n_621: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2103,
        in1(1) => S1999,
        out1 => S1619
    );
nand_n_622: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selMEM_AC,
        in1(1) => U1_dataBus_14,
        out1 => S1620
    );
notg_29: ENTITY WORK.notg
    PORT MAP (
        in1 => S1620,
        out1 => S1621
    );
nor_n_312: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1621,
        in1(1) => U1_selARU_AC,
        out1 => S1622
    );
nand_n_623: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1622,
        in1(1) => S1619,
        out1 => S1623
    );
nor_n_313: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S589,
        in1(1) => S579,
        out1 => S1624
    );
nor_n_314: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1624,
        in1(1) => S590,
        out1 => S1625
    );
nand_n_624: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1625,
        in1(1) => S597,
        out1 => S1626
    );
nand_n_625: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S685,
        in1(1) => S607,
        out1 => S1627
    );
nand_n_626: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1627,
        in1(1) => U1_ADD,
        out1 => S1628
    );
nor_n_315: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1628,
        in1(1) => S686,
        out1 => S1629
    );
nor_n_316: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1629,
        in1(1) => S2000,
        out1 => S1630
    );
nand_n_627: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1630,
        in1(1) => S1626,
        out1 => S1631
    );
nand_n_628: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1631,
        in1(1) => S1623,
        out1 => S1632
    );
nand_n_629: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1632,
        in1(1) => S2001,
        out1 => S1633
    );
nand_n_630: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S768,
        in1(1) => U1_selLGU_AC,
        out1 => S1634
    );
nand_n_631: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1634,
        in1(1) => U1_ldAC,
        out1 => S1635
    );
notg_30: ENTITY WORK.notg
    PORT MAP (
        in1 => S1635,
        out1 => S1636
    );
nand_n_632: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1636,
        in1(1) => S1633,
        out1 => S1637
    );
nand_n_633: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1637,
        in1(1) => S1618,
        out1 => S88
    );
nand_n_634: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1352,
        in1(1) => U1_AC_out_15,
        out1 => S1638
    );
nand_n_635: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S701,
        in1(1) => U1_selARU_AC,
        out1 => S1639
    );
nor_n_317: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2020,
        in1(1) => U1_selMEM_AC,
        out1 => S1640
    );
nand_n_636: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selMEM_AC,
        in1(1) => S1793,
        out1 => S1641
    );
nand_n_637: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1641,
        in1(1) => S2000,
        out1 => S1642
    );
nor_n_318: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1642,
        in1(1) => S1640,
        out1 => S1643
    );
nor_n_319: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1643,
        in1(1) => U1_selLGU_AC,
        out1 => S1644
    );
nand_n_638: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1644,
        in1(1) => S1639,
        out1 => S1645
    );
nor_n_320: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_LGU_out_15,
        in1(1) => S2001,
        out1 => S1646
    );
nor_n_321: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1646,
        in1(1) => S1960,
        out1 => S1647
    );
nand_n_639: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1647,
        in1(1) => S1645,
        out1 => S1648
    );
nand_n_640: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1648,
        in1(1) => S1638,
        out1 => S89
    );
nand_n_641: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2002,
        in1(1) => U1_V_out1,
        out1 => S1649
    );
nand_n_642: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S704,
        in1(1) => U1_selSET_SR,
        out1 => S1650
    );
nor_n_322: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_selSET_SR,
        in1(1) => U1_IR_out_0,
        out1 => S1651
    );
nor_n_323: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1651,
        in1(1) => S2002,
        out1 => S1652
    );
nand_n_643: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1652,
        in1(1) => S1650,
        out1 => S1653
    );
nand_n_644: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1653,
        in1(1) => S1649,
        out1 => S90
    );
nand_n_645: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2003,
        in1(1) => U1_C_out1,
        out1 => S1654
    );
nand_n_646: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S707,
        in1(1) => U1_selSET_SR,
        out1 => S1655
    );
nor_n_324: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_selSET_SR,
        in1(1) => U1_IR_out_1,
        out1 => S1656
    );
nor_n_325: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1656,
        in1(1) => S2003,
        out1 => S1657
    );
nand_n_647: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1657,
        in1(1) => S1655,
        out1 => S1658
    );
nand_n_648: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1658,
        in1(1) => S1654,
        out1 => S91
    );
nand_n_649: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2004,
        in1(1) => U1_N_out1,
        out1 => S1659
    );
nand_n_650: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2253,
        in1(1) => U1_selSET_SR,
        out1 => S1660
    );
nor_n_326: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_selSET_SR,
        in1(1) => U1_IR_out_2,
        out1 => S1661
    );
nor_n_327: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1661,
        in1(1) => S2004,
        out1 => S1662
    );
nand_n_651: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1662,
        in1(1) => S1660,
        out1 => S1663
    );
nand_n_652: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1663,
        in1(1) => S1659,
        out1 => S92
    );
nand_n_653: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2005,
        in1(1) => U1_Z_out1,
        out1 => S1664
    );
nand_n_654: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1102,
        in1(1) => U1_selSET_SR,
        out1 => S1665
    );
nor_n_328: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_selSET_SR,
        in1(1) => U1_IR_out_3,
        out1 => S1666
    );
nor_n_329: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1666,
        in1(1) => S2005,
        out1 => S1667
    );
nand_n_655: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1667,
        in1(1) => S1665,
        out1 => S1668
    );
nand_n_656: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1668,
        in1(1) => S1664,
        out1 => S93
    );
nor_n_330: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1992,
        in1(1) => U1_dataBus_0,
        out1 => S1669
    );
nor_n_331: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_selMEM_IN,
        in1(1) => S1958,
        out1 => S1670
    );
notg_31: ENTITY WORK.notg
    PORT MAP (
        in1 => S1670,
        out1 => S1671
    );
nor_n_332: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1670,
        in1(1) => S1669,
        out1 => S1672
    );
nor_n_333: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1672,
        in1(1) => S2006,
        out1 => S1673
    );
nor_n_334: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_ldIN,
        in1(1) => U1_IN_out_0,
        out1 => S1674
    );
nor_n_335: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1674,
        in1(1) => S1673,
        out1 => S94
    );
nor_n_336: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1670,
        in1(1) => U1_dataBus_1,
        out1 => S1675
    );
nor_n_337: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1671,
        in1(1) => S1956,
        out1 => S1676
    );
nand_n_657: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1670,
        in1(1) => U1_dataBus_1,
        out1 => S1677
    );
nor_n_338: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1675,
        in1(1) => S2006,
        out1 => S1678
    );
nand_n_658: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1678,
        in1(1) => S1677,
        out1 => S1679
    );
nand_n_659: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2006,
        in1(1) => U1_IN_out_1,
        out1 => S1680
    );
nand_n_660: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1680,
        in1(1) => S1679,
        out1 => S95
    );
nor_n_339: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1677,
        in1(1) => S1954,
        out1 => S1681
    );
notg_32: ENTITY WORK.notg
    PORT MAP (
        in1 => S1681,
        out1 => S1682
    );
nor_n_340: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1676,
        in1(1) => U1_dataBus_2,
        out1 => S1683
    );
nor_n_341: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1683,
        in1(1) => S1681,
        out1 => S1684
    );
nor_n_342: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1684,
        in1(1) => S2006,
        out1 => S1685
    );
nor_n_343: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_ldIN,
        in1(1) => U1_IN_out_2,
        out1 => S1686
    );
nor_n_344: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1686,
        in1(1) => S1685,
        out1 => S96
    );
nor_n_345: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1681,
        in1(1) => U1_dataBus_3,
        out1 => S1687
    );
nor_n_346: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1682,
        in1(1) => S1953,
        out1 => S1688
    );
nand_n_661: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1681,
        in1(1) => U1_dataBus_3,
        out1 => S1689
    );
nor_n_347: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1688,
        in1(1) => S1687,
        out1 => S1690
    );
nor_n_348: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1690,
        in1(1) => S2006,
        out1 => S1691
    );
nor_n_349: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_ldIN,
        in1(1) => U1_IN_out_3,
        out1 => S1692
    );
nor_n_350: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1692,
        in1(1) => S1691,
        out1 => S97
    );
nor_n_351: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1688,
        in1(1) => U1_dataBus_4,
        out1 => S1693
    );
nor_n_352: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1689,
        in1(1) => S1951,
        out1 => S1694
    );
nor_n_353: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1694,
        in1(1) => S1693,
        out1 => S1695
    );
nor_n_354: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1695,
        in1(1) => S2006,
        out1 => S1696
    );
nor_n_355: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_ldIN,
        in1(1) => U1_IN_out_4,
        out1 => S1697
    );
nor_n_356: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1697,
        in1(1) => S1696,
        out1 => S98
    );
nand_n_662: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_dataBus_4,
        in1(1) => U1_dataBus_5,
        out1 => S1698
    );
nor_n_357: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1698,
        in1(1) => S1689,
        out1 => S1699
    );
notg_33: ENTITY WORK.notg
    PORT MAP (
        in1 => S1699,
        out1 => S1700
    );
nor_n_358: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1694,
        in1(1) => U1_dataBus_5,
        out1 => S1701
    );
nor_n_359: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1701,
        in1(1) => S1699,
        out1 => S1702
    );
nor_n_360: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1702,
        in1(1) => S2006,
        out1 => S1703
    );
nor_n_361: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_ldIN,
        in1(1) => U1_IN_out_5,
        out1 => S1704
    );
nor_n_362: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1704,
        in1(1) => S1703,
        out1 => S99
    );
nor_n_363: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1700,
        in1(1) => S1950,
        out1 => S1705
    );
notg_34: ENTITY WORK.notg
    PORT MAP (
        in1 => S1705,
        out1 => S1706
    );
nor_n_364: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1699,
        in1(1) => U1_dataBus_6,
        out1 => S1707
    );
nor_n_365: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1707,
        in1(1) => S1705,
        out1 => S1708
    );
nor_n_366: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1708,
        in1(1) => S2006,
        out1 => S1709
    );
nor_n_367: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_ldIN,
        in1(1) => U1_IN_out_6,
        out1 => S1710
    );
nor_n_368: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1710,
        in1(1) => S1709,
        out1 => S100
    );
nand_n_663: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2006,
        in1(1) => U1_IN_out_7,
        out1 => S1711
    );
nor_n_369: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1706,
        in1(1) => S1949,
        out1 => S1712
    );
notg_35: ENTITY WORK.notg
    PORT MAP (
        in1 => S1712,
        out1 => S1713
    );
nor_n_370: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1705,
        in1(1) => U1_dataBus_7,
        out1 => S1714
    );
nor_n_371: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1714,
        in1(1) => S1712,
        out1 => S1715
    );
nand_n_664: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1715,
        in1(1) => U1_ldIN,
        out1 => S1716
    );
nand_n_665: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1716,
        in1(1) => S1711,
        out1 => S101
    );
nand_n_666: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2006,
        in1(1) => U1_IN_out_8,
        out1 => S1717
    );
nor_n_372: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1713,
        in1(1) => S1948,
        out1 => S1718
    );
notg_36: ENTITY WORK.notg
    PORT MAP (
        in1 => S1718,
        out1 => S1719
    );
nor_n_373: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1712,
        in1(1) => U1_dataBus_8,
        out1 => S1720
    );
nor_n_374: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1720,
        in1(1) => S1718,
        out1 => S1721
    );
nand_n_667: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1721,
        in1(1) => U1_ldIN,
        out1 => S1722
    );
nand_n_668: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1722,
        in1(1) => S1717,
        out1 => S102
    );
nand_n_669: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2006,
        in1(1) => U1_IN_out_9,
        out1 => S1723
    );
nor_n_375: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1718,
        in1(1) => U1_dataBus_9,
        out1 => S1724
    );
nor_n_376: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1719,
        in1(1) => S1947,
        out1 => S1725
    );
notg_37: ENTITY WORK.notg
    PORT MAP (
        in1 => S1725,
        out1 => S1726
    );
nor_n_377: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1725,
        in1(1) => S1724,
        out1 => S1727
    );
nand_n_670: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1727,
        in1(1) => U1_ldIN,
        out1 => S1728
    );
nand_n_671: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1728,
        in1(1) => S1723,
        out1 => S103
    );
nand_n_672: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2006,
        in1(1) => U1_IN_out_10,
        out1 => S1729
    );
nor_n_378: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1726,
        in1(1) => S1946,
        out1 => S1730
    );
notg_38: ENTITY WORK.notg
    PORT MAP (
        in1 => S1730,
        out1 => S1731
    );
nor_n_379: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1725,
        in1(1) => U1_dataBus_10,
        out1 => S1732
    );
nor_n_380: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1732,
        in1(1) => S1730,
        out1 => S1733
    );
nand_n_673: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1733,
        in1(1) => U1_ldIN,
        out1 => S1734
    );
nand_n_674: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1734,
        in1(1) => S1729,
        out1 => S104
    );
nand_n_675: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2006,
        in1(1) => U1_IN_out_11,
        out1 => S1735
    );
nor_n_381: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1730,
        in1(1) => U1_dataBus_11,
        out1 => S1736
    );
nor_n_382: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1731,
        in1(1) => S1945,
        out1 => S1737
    );
notg_39: ENTITY WORK.notg
    PORT MAP (
        in1 => S1737,
        out1 => S1738
    );
nor_n_383: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1737,
        in1(1) => S1736,
        out1 => S1739
    );
nand_n_676: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1739,
        in1(1) => U1_ldIN,
        out1 => S1740
    );
nand_n_677: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1740,
        in1(1) => S1735,
        out1 => S105
    );
nand_n_678: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2006,
        in1(1) => U1_IN_out_12,
        out1 => S1741
    );
nor_n_384: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1738,
        in1(1) => S1944,
        out1 => S1742
    );
notg_40: ENTITY WORK.notg
    PORT MAP (
        in1 => S1742,
        out1 => S1743
    );
nor_n_385: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1737,
        in1(1) => U1_dataBus_12,
        out1 => S1744
    );
nor_n_386: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1744,
        in1(1) => S1742,
        out1 => S1745
    );
nand_n_679: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1745,
        in1(1) => U1_ldIN,
        out1 => S1746
    );
nand_n_680: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1746,
        in1(1) => S1741,
        out1 => S106
    );
nand_n_681: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2006,
        in1(1) => U1_IN_out_13,
        out1 => S1747
    );
nor_n_387: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1742,
        in1(1) => U1_dataBus_13,
        out1 => S1748
    );
nor_n_388: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1743,
        in1(1) => S1943,
        out1 => S1749
    );
notg_41: ENTITY WORK.notg
    PORT MAP (
        in1 => S1749,
        out1 => S1750
    );
nor_n_389: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1749,
        in1(1) => S1748,
        out1 => S1751
    );
nand_n_682: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1751,
        in1(1) => U1_ldIN,
        out1 => S1752
    );
nand_n_683: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1752,
        in1(1) => S1747,
        out1 => S107
    );
nand_n_684: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2006,
        in1(1) => U1_IN_out_14,
        out1 => S1753
    );
nor_n_390: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1750,
        in1(1) => S1942,
        out1 => S1754
    );
nor_n_391: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1749,
        in1(1) => U1_dataBus_14,
        out1 => S1755
    );
nor_n_392: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1755,
        in1(1) => S1754,
        out1 => S1756
    );
nand_n_685: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1756,
        in1(1) => U1_ldIN,
        out1 => S1757
    );
nand_n_686: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1757,
        in1(1) => S1753,
        out1 => S108
    );
nand_n_687: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2006,
        in1(1) => U1_IN_out_15,
        out1 => S1758
    );
nand_n_688: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1754,
        in1(1) => U1_dataBus_15,
        out1 => S1759
    );
nor_n_393: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1754,
        in1(1) => U1_dataBus_15,
        out1 => S1760
    );
nor_n_394: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1760,
        in1(1) => S2006,
        out1 => S1761
    );
nand_n_689: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1761,
        in1(1) => S1759,
        out1 => S1762
    );
nand_n_690: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1762,
        in1(1) => S1758,
        out1 => S109
    );
nand_n_691: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2180,
        in1(1) => U1_selIMM_PC,
        out1 => S1763
    );
nand_n_692: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1105,
        in1(1) => S1967,
        out1 => S1764
    );
nand_n_693: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selMEM_PC,
        in1(1) => U1_dataBus_0,
        out1 => S1765
    );
nand_n_694: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1765,
        in1(1) => S1764,
        out1 => S1766
    );
nand_n_695: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1766,
        in1(1) => S1968,
        out1 => S1767
    );
nand_n_696: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1767,
        in1(1) => S1763,
        out1 => S1768
    );
nand_n_697: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1768,
        in1(1) => U1_ldPC,
        out1 => S1769
    );
nand_n_698: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2007,
        in1(1) => U1_PC_out_0,
        out1 => S1770
    );
nand_n_699: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1770,
        in1(1) => S1769,
        out1 => S110
    );
nand_n_700: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2168,
        in1(1) => U1_selIMM_PC,
        out1 => S1771
    );
nor_n_395: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1115,
        in1(1) => U1_selMEM_PC,
        out1 => S1772
    );
nand_n_701: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selMEM_PC,
        in1(1) => U1_dataBus_1,
        out1 => S1773
    );
nand_n_702: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1773,
        in1(1) => S1968,
        out1 => S1774
    );
nor_n_396: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1774,
        in1(1) => S1772,
        out1 => S1775
    );
nand_n_703: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2007,
        in1(1) => U1_PC_out_1,
        out1 => S1776
    );
nor_n_397: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1775,
        in1(1) => S2007,
        out1 => S1777
    );
nand_n_704: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1777,
        in1(1) => S1771,
        out1 => S1778
    );
nand_n_705: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1778,
        in1(1) => S1776,
        out1 => S111
    );
nand_n_706: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2153,
        in1(1) => U1_selIMM_PC,
        out1 => S1779
    );
nand_n_707: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1123,
        in1(1) => S1967,
        out1 => S1780
    );
nand_n_708: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selMEM_PC,
        in1(1) => U1_dataBus_2,
        out1 => S1781
    );
nand_n_709: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1781,
        in1(1) => S1780,
        out1 => S1782
    );
nand_n_710: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1782,
        in1(1) => S1968,
        out1 => S1783
    );
nand_n_711: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1783,
        in1(1) => S1779,
        out1 => S1784
    );
nand_n_712: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1784,
        in1(1) => U1_ldPC,
        out1 => S1785
    );
nand_n_713: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2007,
        in1(1) => U1_PC_out_2,
        out1 => S1786
    );
nand_n_714: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1786,
        in1(1) => S1785,
        out1 => S112
    );
nand_n_715: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2142,
        in1(1) => U1_selIMM_PC,
        out1 => S1787
    );
nand_n_716: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1131,
        in1(1) => S1967,
        out1 => S1788
    );
nand_n_717: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selMEM_PC,
        in1(1) => U1_dataBus_3,
        out1 => S1789
    );
nand_n_718: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1789,
        in1(1) => S1788,
        out1 => S1790
    );
nand_n_719: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1790,
        in1(1) => S1968,
        out1 => S1791
    );
nand_n_720: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1791,
        in1(1) => S1787,
        out1 => S1792
    );
nand_n_721: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1792,
        in1(1) => U1_ldPC,
        out1 => S1794
    );
nand_n_722: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2007,
        in1(1) => U1_PC_out_3,
        out1 => S1795
    );
nand_n_723: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1795,
        in1(1) => S1794,
        out1 => S113
    );
nand_n_724: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2227,
        in1(1) => U1_selIMM_PC,
        out1 => S1796
    );
nand_n_725: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selMEM_PC,
        in1(1) => U1_dataBus_4,
        out1 => S1797
    );
nand_n_726: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1139,
        in1(1) => S1967,
        out1 => S1798
    );
nand_n_727: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1798,
        in1(1) => S1797,
        out1 => S1799
    );
nand_n_728: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1799,
        in1(1) => S1968,
        out1 => S1800
    );
nand_n_729: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1800,
        in1(1) => S1796,
        out1 => S1801
    );
nand_n_730: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1801,
        in1(1) => U1_ldPC,
        out1 => S1802
    );
nand_n_731: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2007,
        in1(1) => U1_PC_out_4,
        out1 => S1804
    );
nand_n_732: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1804,
        in1(1) => S1802,
        out1 => S114
    );
nand_n_733: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2215,
        in1(1) => U1_selIMM_PC,
        out1 => S1805
    );
nand_n_734: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selMEM_PC,
        in1(1) => U1_dataBus_5,
        out1 => S1806
    );
nand_n_735: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1147,
        in1(1) => S1967,
        out1 => S1807
    );
nand_n_736: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1807,
        in1(1) => S1806,
        out1 => S1808
    );
nand_n_737: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1808,
        in1(1) => S1968,
        out1 => S1809
    );
nand_n_738: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1809,
        in1(1) => S1805,
        out1 => S1810
    );
nand_n_739: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1810,
        in1(1) => U1_ldPC,
        out1 => S1811
    );
nand_n_740: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2007,
        in1(1) => U1_PC_out_5,
        out1 => S1812
    );
nand_n_741: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1812,
        in1(1) => S1811,
        out1 => S115
    );
nand_n_742: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2204,
        in1(1) => U1_selIMM_PC,
        out1 => S1814
    );
nand_n_743: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selMEM_PC,
        in1(1) => U1_dataBus_6,
        out1 => S1815
    );
nand_n_744: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1155,
        in1(1) => S1967,
        out1 => S1816
    );
nand_n_745: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1816,
        in1(1) => S1815,
        out1 => S1817
    );
nand_n_746: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1817,
        in1(1) => S1968,
        out1 => S1818
    );
nand_n_747: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1818,
        in1(1) => S1814,
        out1 => S1819
    );
nand_n_748: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1819,
        in1(1) => U1_ldPC,
        out1 => S1820
    );
nand_n_749: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2007,
        in1(1) => U1_PC_out_6,
        out1 => S1821
    );
nand_n_750: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1821,
        in1(1) => S1820,
        out1 => S116
    );
nand_n_751: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2195,
        in1(1) => U1_selIMM_PC,
        out1 => S1823
    );
nand_n_752: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selMEM_PC,
        in1(1) => U1_dataBus_7,
        out1 => S1824
    );
nand_n_753: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1163,
        in1(1) => S1967,
        out1 => S1825
    );
nand_n_754: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1825,
        in1(1) => S1824,
        out1 => S1826
    );
nand_n_755: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1826,
        in1(1) => S1968,
        out1 => S1827
    );
nand_n_756: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1827,
        in1(1) => S1823,
        out1 => S1828
    );
nand_n_757: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1828,
        in1(1) => U1_ldPC,
        out1 => S1829
    );
nand_n_758: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2007,
        in1(1) => U1_PC_out_7,
        out1 => S1830
    );
nand_n_759: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1830,
        in1(1) => S1829,
        out1 => S117
    );
nand_n_760: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2079,
        in1(1) => U1_selIMM_PC,
        out1 => S1831
    );
nand_n_761: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selMEM_PC,
        in1(1) => U1_dataBus_8,
        out1 => S1833
    );
nand_n_762: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1171,
        in1(1) => S1967,
        out1 => S1834
    );
nand_n_763: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1834,
        in1(1) => S1833,
        out1 => S1835
    );
nand_n_764: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1835,
        in1(1) => S1968,
        out1 => S1836
    );
nand_n_765: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1836,
        in1(1) => S1831,
        out1 => S1837
    );
nand_n_766: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1837,
        in1(1) => U1_ldPC,
        out1 => S1838
    );
nand_n_767: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2007,
        in1(1) => U1_PC_out_8,
        out1 => S1839
    );
nand_n_768: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1839,
        in1(1) => S1838,
        out1 => S118
    );
nand_n_769: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2070,
        in1(1) => U1_selIMM_PC,
        out1 => S1840
    );
nand_n_770: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selMEM_PC,
        in1(1) => U1_dataBus_9,
        out1 => S1841
    );
nand_n_771: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1179,
        in1(1) => S1967,
        out1 => S1843
    );
nand_n_772: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1843,
        in1(1) => S1841,
        out1 => S1844
    );
nand_n_773: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1844,
        in1(1) => S1968,
        out1 => S1845
    );
nand_n_774: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1845,
        in1(1) => S1840,
        out1 => S1846
    );
nand_n_775: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1846,
        in1(1) => U1_ldPC,
        out1 => S1847
    );
nand_n_776: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2007,
        in1(1) => U1_PC_out_9,
        out1 => S1848
    );
nand_n_777: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1848,
        in1(1) => S1847,
        out1 => S119
    );
nand_n_778: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2058,
        in1(1) => U1_selIMM_PC,
        out1 => S1849
    );
nand_n_779: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selMEM_PC,
        in1(1) => U1_dataBus_10,
        out1 => S1850
    );
nand_n_780: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1187,
        in1(1) => S1967,
        out1 => S1851
    );
nand_n_781: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1851,
        in1(1) => S1850,
        out1 => S1853
    );
nand_n_782: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1853,
        in1(1) => S1968,
        out1 => S1854
    );
nand_n_783: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1854,
        in1(1) => S1849,
        out1 => S1855
    );
nand_n_784: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1855,
        in1(1) => U1_ldPC,
        out1 => S1856
    );
nand_n_785: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2007,
        in1(1) => U1_PC_out_10,
        out1 => S1857
    );
nand_n_786: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1857,
        in1(1) => S1856,
        out1 => S120
    );
nand_n_787: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2050,
        in1(1) => U1_selIMM_PC,
        out1 => S1858
    );
nand_n_788: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selMEM_PC,
        in1(1) => U1_dataBus_11,
        out1 => S1859
    );
nand_n_789: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1195,
        in1(1) => S1967,
        out1 => S1860
    );
nand_n_790: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1860,
        in1(1) => S1859,
        out1 => S1861
    );
nand_n_791: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1861,
        in1(1) => S1968,
        out1 => S1863
    );
nand_n_792: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1863,
        in1(1) => S1858,
        out1 => S1864
    );
nand_n_793: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1864,
        in1(1) => U1_ldPC,
        out1 => S1865
    );
nand_n_794: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2007,
        in1(1) => U1_PC_out_11,
        out1 => S1866
    );
nand_n_795: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1866,
        in1(1) => S1865,
        out1 => S121
    );
nand_n_796: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2122,
        in1(1) => U1_selIMM_PC,
        out1 => S1867
    );
nand_n_797: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selMEM_PC,
        in1(1) => U1_dataBus_12,
        out1 => S1868
    );
nand_n_798: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1203,
        in1(1) => S1967,
        out1 => S1869
    );
nand_n_799: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1869,
        in1(1) => S1868,
        out1 => S1870
    );
nand_n_800: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1870,
        in1(1) => S1968,
        out1 => S1871
    );
nand_n_801: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1871,
        in1(1) => S1867,
        out1 => S1873
    );
nand_n_802: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1873,
        in1(1) => U1_ldPC,
        out1 => S1874
    );
nand_n_803: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2007,
        in1(1) => U1_PC_out_12,
        out1 => S1875
    );
nand_n_804: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1875,
        in1(1) => S1874,
        out1 => S122
    );
nand_n_805: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2113,
        in1(1) => U1_selIMM_PC,
        out1 => S1876
    );
nand_n_806: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selMEM_PC,
        in1(1) => U1_dataBus_13,
        out1 => S1877
    );
nand_n_807: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1211,
        in1(1) => S1967,
        out1 => S1878
    );
nand_n_808: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1878,
        in1(1) => S1877,
        out1 => S1879
    );
nand_n_809: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1879,
        in1(1) => S1968,
        out1 => S1880
    );
nand_n_810: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1880,
        in1(1) => S1876,
        out1 => S1881
    );
nand_n_811: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1881,
        in1(1) => U1_ldPC,
        out1 => S1883
    );
nand_n_812: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2007,
        in1(1) => U1_PC_out_13,
        out1 => S1884
    );
nand_n_813: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1884,
        in1(1) => S1883,
        out1 => S123
    );
nand_n_814: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2103,
        in1(1) => U1_selIMM_PC,
        out1 => S1885
    );
nand_n_815: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selMEM_PC,
        in1(1) => U1_dataBus_14,
        out1 => S1886
    );
nand_n_816: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1219,
        in1(1) => S1967,
        out1 => S1887
    );
nand_n_817: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1887,
        in1(1) => S1886,
        out1 => S1888
    );
nand_n_818: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1888,
        in1(1) => S1968,
        out1 => S1889
    );
nand_n_819: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1889,
        in1(1) => S1885,
        out1 => S1890
    );
nand_n_820: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1890,
        in1(1) => U1_ldPC,
        out1 => S1891
    );
nand_n_821: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2007,
        in1(1) => U1_PC_out_14,
        out1 => S1893
    );
nand_n_822: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1893,
        in1(1) => S1891,
        out1 => S124
    );
nand_n_823: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2020,
        in1(1) => U1_selIMM_PC,
        out1 => S1894
    );
nand_n_824: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_selMEM_PC,
        in1(1) => U1_dataBus_15,
        out1 => S1895
    );
nand_n_825: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1228,
        in1(1) => S1967,
        out1 => S1896
    );
nand_n_826: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1896,
        in1(1) => S1895,
        out1 => S1897
    );
nand_n_827: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1897,
        in1(1) => S1968,
        out1 => S1898
    );
nand_n_828: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1898,
        in1(1) => S1894,
        out1 => S1899
    );
nand_n_829: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1899,
        in1(1) => U1_ldPC,
        out1 => S1900
    );
nand_n_830: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2007,
        in1(1) => U1_PC_out_15,
        out1 => S1901
    );
nand_n_831: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1901,
        in1(1) => S1900,
        out1 => S125
    );
nand_n_832: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_ldIR,
        in1(1) => U1_dataBus_0,
        out1 => S1903
    );
nand_n_833: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2008,
        in1(1) => U1_IR_out_0,
        out1 => S1904
    );
nand_n_834: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1904,
        in1(1) => S1903,
        out1 => S126
    );
nand_n_835: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_ldIR,
        in1(1) => U1_dataBus_1,
        out1 => S1905
    );
nand_n_836: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2008,
        in1(1) => U1_IR_out_1,
        out1 => S1906
    );
nand_n_837: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1906,
        in1(1) => S1905,
        out1 => S127
    );
nand_n_838: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_ldIR,
        in1(1) => U1_dataBus_2,
        out1 => S1907
    );
nand_n_839: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2008,
        in1(1) => U1_IR_out_2,
        out1 => S1908
    );
nand_n_840: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1908,
        in1(1) => S1907,
        out1 => S128
    );
nand_n_841: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_ldIR,
        in1(1) => U1_dataBus_3,
        out1 => S1910
    );
nand_n_842: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2008,
        in1(1) => U1_IR_out_3,
        out1 => S1911
    );
nand_n_843: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1911,
        in1(1) => S1910,
        out1 => S129
    );
nand_n_844: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_ldIR,
        in1(1) => U1_dataBus_4,
        out1 => S1912
    );
nand_n_845: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2008,
        in1(1) => U1_IR_out_4,
        out1 => S1913
    );
nand_n_846: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1913,
        in1(1) => S1912,
        out1 => S130
    );
nand_n_847: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_ldIR,
        in1(1) => U1_dataBus_5,
        out1 => S1914
    );
nand_n_848: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2008,
        in1(1) => U1_IR_out_5,
        out1 => S1915
    );
nand_n_849: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1915,
        in1(1) => S1914,
        out1 => S131
    );
nand_n_850: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_ldIR,
        in1(1) => U1_dataBus_6,
        out1 => S1916
    );
nand_n_851: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2008,
        in1(1) => U1_IR_out_6,
        out1 => S1918
    );
nand_n_852: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1918,
        in1(1) => S1916,
        out1 => S132
    );
nand_n_853: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_ldIR,
        in1(1) => U1_dataBus_7,
        out1 => S1919
    );
nand_n_854: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2008,
        in1(1) => U1_IR_out_7,
        out1 => S1920
    );
nand_n_855: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1920,
        in1(1) => S1919,
        out1 => S133
    );
nand_n_856: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_ldIR,
        in1(1) => U1_dataBus_8,
        out1 => S1921
    );
nand_n_857: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2008,
        in1(1) => U1_IR_out_8,
        out1 => S1922
    );
nand_n_858: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1922,
        in1(1) => S1921,
        out1 => S134
    );
nand_n_859: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_ldIR,
        in1(1) => U1_dataBus_9,
        out1 => S1923
    );
nand_n_860: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2008,
        in1(1) => U1_IR_out_9,
        out1 => S1924
    );
nand_n_861: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1924,
        in1(1) => S1923,
        out1 => S135
    );
nand_n_862: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_ldIR,
        in1(1) => U1_dataBus_10,
        out1 => S1926
    );
nand_n_863: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2008,
        in1(1) => U1_IR_out_10,
        out1 => S1927
    );
nand_n_864: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1927,
        in1(1) => S1926,
        out1 => S136
    );
nand_n_865: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_ldIR,
        in1(1) => U1_dataBus_11,
        out1 => S1928
    );
nand_n_866: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2008,
        in1(1) => U1_IR_out_11,
        out1 => S1929
    );
nand_n_867: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1929,
        in1(1) => S1928,
        out1 => S137
    );
nand_n_868: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_ldIR,
        in1(1) => U1_dataBus_12,
        out1 => S1930
    );
nand_n_869: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_IR_out_12,
        in1(1) => S2008,
        out1 => S1931
    );
nand_n_870: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1931,
        in1(1) => S1930,
        out1 => S138
    );
nand_n_871: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_ldIR,
        in1(1) => U1_dataBus_13,
        out1 => S1933
    );
nand_n_872: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_IR_out_13,
        in1(1) => S2008,
        out1 => S1934
    );
nand_n_873: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1934,
        in1(1) => S1933,
        out1 => S139
    );
nand_n_874: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_ldIR,
        in1(1) => U1_dataBus_14,
        out1 => S1935
    );
nand_n_875: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_IR_out_14,
        in1(1) => S2008,
        out1 => S1936
    );
nand_n_876: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1936,
        in1(1) => S1935,
        out1 => S140
    );
nand_n_877: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_ldIR,
        in1(1) => U1_dataBus_15,
        out1 => S1937
    );
nand_n_878: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_IR_out_15,
        in1(1) => S2008,
        out1 => S1938
    );
nand_n_879: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1938,
        in1(1) => S1937,
        out1 => S141
    );
notg_42: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_dataBus_15,
        out1 => S1793
    );
notg_43: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_conOF,
        out1 => S1803
    );
notg_44: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_IR_out_3,
        out1 => S1813
    );
notg_45: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_SE12bits,
        out1 => S1822
    );
notg_46: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_SE4bits,
        out1 => S1832
    );
notg_47: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_selMEM_LGU,
        out1 => S1842
    );
notg_48: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_AC_out_4,
        out1 => S1852
    );
notg_49: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_AC_out_6,
        out1 => S1862
    );
notg_50: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_AC_out_5,
        out1 => S1872
    );
notg_51: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_AC_out_7,
        out1 => S1882
    );
notg_52: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_AC_out_10,
        out1 => S1892
    );
notg_53: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_AC_out_14,
        out1 => S1902
    );
notg_54: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_AC_out_15,
        out1 => S1909
    );
notg_55: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_AC_out_0,
        out1 => S1917
    );
notg_56: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_AC_out_1,
        out1 => S1925
    );
notg_57: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_AC_out_2,
        out1 => S1932
    );
notg_58: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_AC_out_3,
        out1 => S1939
    );
notg_59: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_SHF_1,
        out1 => S1940
    );
notg_60: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_SHF_0,
        out1 => S1941
    );
notg_61: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_dataBus_14,
        out1 => S1942
    );
notg_62: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_dataBus_13,
        out1 => S1943
    );
notg_63: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_dataBus_12,
        out1 => S1944
    );
notg_64: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_dataBus_11,
        out1 => S1945
    );
notg_65: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_dataBus_10,
        out1 => S1946
    );
notg_66: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_dataBus_9,
        out1 => S1947
    );
notg_67: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_dataBus_8,
        out1 => S1948
    );
notg_68: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_dataBus_7,
        out1 => S1949
    );
notg_69: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_dataBus_6,
        out1 => S1950
    );
notg_70: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_dataBus_4,
        out1 => S1951
    );
notg_71: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_IR_out_4,
        out1 => S1952
    );
notg_72: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_dataBus_3,
        out1 => S1953
    );
notg_73: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_dataBus_2,
        out1 => S1954
    );
notg_74: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_IR_out_2,
        out1 => S1955
    );
notg_75: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_dataBus_1,
        out1 => S1956
    );
notg_76: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_IR_out_0,
        out1 => S1957
    );
notg_77: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_dataBus_0,
        out1 => S1958
    );
notg_78: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_NOT,
        out1 => S1959
    );
notg_79: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_ldAC,
        out1 => S1960
    );
notg_80: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_PC_out_12,
        out1 => S1961
    );
notg_81: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_selIMM_OF,
        out1 => S1962
    );
notg_82: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_PC_out_13,
        out1 => S1963
    );
notg_83: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_PC_out_14,
        out1 => S1964
    );
notg_84: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_INC1,
        out1 => S1965
    );
notg_85: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_PC_out_0,
        out1 => S1966
    );
notg_86: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_selMEM_PC,
        out1 => S1967
    );
notg_87: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_selIMM_PC,
        out1 => S1968
    );
notg_88: ENTITY WORK.notg
    PORT MAP (
        in1 => S27,
        out1 => S1969
    );
notg_89: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_PC_out_2,
        out1 => S1970
    );
notg_90: ENTITY WORK.notg
    PORT MAP (
        in1 => S28,
        out1 => S1971
    );
notg_91: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_PC_out_3,
        out1 => S1972
    );
notg_92: ENTITY WORK.notg
    PORT MAP (
        in1 => S29,
        out1 => S1973
    );
notg_93: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_PC_out_4,
        out1 => S1974
    );
notg_94: ENTITY WORK.notg
    PORT MAP (
        in1 => S30,
        out1 => S1975
    );
notg_95: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_PC_out_5,
        out1 => S1976
    );
notg_96: ENTITY WORK.notg
    PORT MAP (
        in1 => S31,
        out1 => S1977
    );
notg_97: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_PC_out_6,
        out1 => S1978
    );
notg_98: ENTITY WORK.notg
    PORT MAP (
        in1 => S32,
        out1 => S1979
    );
notg_99: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_PC_out_7,
        out1 => S1980
    );
notg_100: ENTITY WORK.notg
    PORT MAP (
        in1 => S33,
        out1 => S1981
    );
notg_101: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_PC_out_8,
        out1 => S1982
    );
notg_102: ENTITY WORK.notg
    PORT MAP (
        in1 => S34,
        out1 => S1983
    );
notg_103: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_PC_out_9,
        out1 => S1984
    );
notg_104: ENTITY WORK.notg
    PORT MAP (
        in1 => S35,
        out1 => S1985
    );
notg_105: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_PC_out_10,
        out1 => S1986
    );
notg_106: ENTITY WORK.notg
    PORT MAP (
        in1 => S36,
        out1 => S1987
    );
notg_107: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_PC_out_11,
        out1 => S1988
    );
notg_108: ENTITY WORK.notg
    PORT MAP (
        in1 => S37,
        out1 => S1989
    );
notg_109: ENTITY WORK.notg
    PORT MAP (
        in1 => S38,
        out1 => S1990
    );
notg_110: ENTITY WORK.notg
    PORT MAP (
        in1 => S39,
        out1 => S1991
    );
notg_111: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_selMEM_IN,
        out1 => S1992
    );
notg_112: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_selMO_ARU,
        out1 => S1993
    );
notg_113: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_MUL,
        out1 => S1994
    );
notg_114: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_ADD,
        out1 => S1995
    );
notg_115: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_selPC_MEM,
        out1 => S1996
    );
notg_116: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_selAC_MEM,
        out1 => S1997
    );
notg_117: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_selIR_MEM,
        out1 => S1998
    );
notg_118: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_selMEM_AC,
        out1 => S1999
    );
notg_119: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_selARU_AC,
        out1 => S2000
    );
notg_120: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_selLGU_AC,
        out1 => S2001
    );
notg_121: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_ldSR_0,
        out1 => S2002
    );
notg_122: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_ldSR_0,
        out1 => S2003
    );
notg_123: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_ldSR_0,
        out1 => S2004
    );
notg_124: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_ldSR_0,
        out1 => S2005
    );
notg_125: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_ldIN,
        out1 => S2006
    );
notg_126: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_ldPC,
        out1 => S2007
    );
notg_127: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_ldIR,
        out1 => S2008
    );
nor_n_398: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1822,
        in1(1) => S1813,
        out1 => S2009
    );
nand_n_880: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_SE12bits,
        in1(1) => U1_IR_out_3,
        out1 => S2010
    );
nor_n_399: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2010,
        in1(1) => U1_SE4bits,
        out1 => S2011
    );
nand_n_881: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2009,
        in1(1) => S1832,
        out1 => S2012
    );
nand_n_882: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_SE4bits,
        in1(1) => U1_IR_out_11,
        out1 => S2013
    );
notg_128: ENTITY WORK.notg
    PORT MAP (
        in1 => S2013,
        out1 => S2014
    );
nor_n_400: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2014,
        in1(1) => S2011,
        out1 => S2015
    );
nor_n_401: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_SE12bits,
        in1(1) => S1803,
        out1 => S2016
    );
nand_n_883: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1822,
        in1(1) => U1_conOF,
        out1 => S2017
    );
nor_n_402: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2017,
        in1(1) => U1_SE4bits,
        out1 => S2018
    );
nand_n_884: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2018,
        in1(1) => U1_OF_out_3,
        out1 => S2019
    );
nand_n_885: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2019,
        in1(1) => S2015,
        out1 => S2020
    );
nor_n_403: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2020,
        in1(1) => U1_selMEM_LGU,
        out1 => S2021
    );
nor_n_404: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1842,
        in1(1) => U1_dataBus_15,
        out1 => S2022
    );
nor_n_405: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2022,
        in1(1) => S2021,
        out1 => S2023
    );
nand_n_886: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2023,
        in1(1) => U1_AC_out_15,
        out1 => S2024
    );
notg_129: ENTITY WORK.notg
    PORT MAP (
        in1 => S2024,
        out1 => S2025
    );
nand_n_887: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2024,
        in1(1) => U1_AND,
        out1 => S2026
    );
nor_n_406: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2023,
        in1(1) => S1959,
        out1 => S2027
    );
nor_n_407: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2027,
        in1(1) => U1_AND,
        out1 => S2028
    );
nor_n_408: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_SHF_0,
        in1(1) => S1940,
        out1 => S2029
    );
nand_n_888: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1941,
        in1(1) => U1_SHF_1,
        out1 => S2030
    );
nand_n_889: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1909,
        in1(1) => S1902,
        out1 => S2031
    );
nor_n_409: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2031,
        in1(1) => U1_AC_out_13,
        out1 => S2032
    );
nor_n_410: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_AC_out_9,
        in1(1) => U1_AC_out_10,
        out1 => S2033
    );
nor_n_411: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_AC_out_11,
        in1(1) => U1_AC_out_12,
        out1 => S2034
    );
nand_n_890: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2034,
        in1(1) => S2033,
        out1 => S2035
    );
notg_130: ENTITY WORK.notg
    PORT MAP (
        in1 => S2035,
        out1 => S2036
    );
nor_n_412: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_AC_out_5,
        in1(1) => U1_AC_out_6,
        out1 => S2037
    );
nor_n_413: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_AC_out_7,
        in1(1) => U1_AC_out_8,
        out1 => S2038
    );
nand_n_891: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2038,
        in1(1) => S2037,
        out1 => S2039
    );
nor_n_414: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2039,
        in1(1) => S2035,
        out1 => S2040
    );
nor_n_415: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_AC_out_7,
        in1(1) => U1_AC_out_6,
        out1 => S2041
    );
nand_n_892: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2041,
        in1(1) => S2036,
        out1 => S2042
    );
nor_n_416: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_AC_out_8,
        in1(1) => U1_AC_out_5,
        out1 => S2043
    );
nand_n_893: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2043,
        in1(1) => S2032,
        out1 => S2044
    );
nor_n_417: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2044,
        in1(1) => S2042,
        out1 => S2045
    );
nand_n_894: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2040,
        in1(1) => S2032,
        out1 => S2046
    );
nor_n_418: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2016,
        in1(1) => U1_SE4bits,
        out1 => S2047
    );
nand_n_895: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2017,
        in1(1) => S1832,
        out1 => S2048
    );
nand_n_896: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2048,
        in1(1) => U1_IR_out_11,
        out1 => S2049
    );
nand_n_897: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2049,
        in1(1) => S2012,
        out1 => S2050
    );
nor_n_419: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2050,
        in1(1) => U1_selMEM_LGU,
        out1 => S2051
    );
nor_n_420: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_dataBus_11,
        in1(1) => S1842,
        out1 => S2052
    );
nor_n_421: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2052,
        in1(1) => S2051,
        out1 => S2053
    );
nand_n_898: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2053,
        in1(1) => S2045,
        out1 => S2054
    );
nor_n_422: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2054,
        in1(1) => U1_AC_out_0,
        out1 => S2055
    );
notg_131: ENTITY WORK.notg
    PORT MAP (
        in1 => S2055,
        out1 => S2056
    );
nand_n_899: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2048,
        in1(1) => U1_IR_out_10,
        out1 => S2057
    );
nand_n_900: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2057,
        in1(1) => S2012,
        out1 => S2058
    );
nor_n_423: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2058,
        in1(1) => U1_selMEM_LGU,
        out1 => S2059
    );
nor_n_424: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_dataBus_10,
        in1(1) => S1842,
        out1 => S2060
    );
nor_n_425: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2060,
        in1(1) => S2059,
        out1 => S2061
    );
notg_132: ENTITY WORK.notg
    PORT MAP (
        in1 => S2061,
        out1 => S2062
    );
nor_n_426: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2062,
        in1(1) => S2046,
        out1 => S2063
    );
nand_n_901: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2061,
        in1(1) => S2045,
        out1 => S2064
    );
nand_n_902: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2063,
        in1(1) => U1_AC_out_0,
        out1 => S2065
    );
notg_133: ENTITY WORK.notg
    PORT MAP (
        in1 => S2065,
        out1 => S2066
    );
nor_n_427: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2066,
        in1(1) => S2055,
        out1 => S2067
    );
nand_n_903: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2067,
        in1(1) => S1925,
        out1 => S2068
    );
nand_n_904: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2048,
        in1(1) => U1_IR_out_9,
        out1 => S2069
    );
nand_n_905: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2069,
        in1(1) => S2012,
        out1 => S2070
    );
nor_n_428: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2070,
        in1(1) => U1_selMEM_LGU,
        out1 => S2071
    );
nor_n_429: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_dataBus_9,
        in1(1) => S1842,
        out1 => S2072
    );
nor_n_430: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2072,
        in1(1) => S2071,
        out1 => S2073
    );
nand_n_906: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2073,
        in1(1) => S2045,
        out1 => S2074
    );
notg_134: ENTITY WORK.notg
    PORT MAP (
        in1 => S2074,
        out1 => S2075
    );
nor_n_431: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2074,
        in1(1) => U1_AC_out_0,
        out1 => S2076
    );
notg_135: ENTITY WORK.notg
    PORT MAP (
        in1 => S2076,
        out1 => S2077
    );
nand_n_907: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2048,
        in1(1) => U1_IR_out_8,
        out1 => S2078
    );
nand_n_908: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2078,
        in1(1) => S2012,
        out1 => S2079
    );
nor_n_432: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2079,
        in1(1) => U1_selMEM_LGU,
        out1 => S2080
    );
nor_n_433: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_dataBus_8,
        in1(1) => S1842,
        out1 => S2081
    );
nor_n_434: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2081,
        in1(1) => S2080,
        out1 => S2082
    );
nand_n_909: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2082,
        in1(1) => S2045,
        out1 => S2083
    );
notg_136: ENTITY WORK.notg
    PORT MAP (
        in1 => S2083,
        out1 => S2084
    );
nor_n_435: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2075,
        in1(1) => U1_AC_out_0,
        out1 => S2085
    );
nor_n_436: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2084,
        in1(1) => S1917,
        out1 => S2086
    );
nor_n_437: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2086,
        in1(1) => S2085,
        out1 => S2087
    );
notg_137: ENTITY WORK.notg
    PORT MAP (
        in1 => S2087,
        out1 => S2088
    );
nand_n_910: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2088,
        in1(1) => U1_AC_out_1,
        out1 => S2089
    );
nand_n_911: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2089,
        in1(1) => S2068,
        out1 => S2090
    );
nor_n_438: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2090,
        in1(1) => S1932,
        out1 => S2091
    );
nor_n_439: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2091,
        in1(1) => U1_AC_out_3,
        out1 => S2092
    );
nor_n_440: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2092,
        in1(1) => S2030,
        out1 => S2093
    );
nand_n_912: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2045,
        in1(1) => S2023,
        out1 => S2094
    );
nor_n_441: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2094,
        in1(1) => U1_AC_out_0,
        out1 => S2095
    );
notg_138: ENTITY WORK.notg
    PORT MAP (
        in1 => S2095,
        out1 => S2096
    );
nor_n_442: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2096,
        in1(1) => U1_AC_out_1,
        out1 => S2097
    );
notg_139: ENTITY WORK.notg
    PORT MAP (
        in1 => S2097,
        out1 => S2098
    );
nor_n_443: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_SHF_1,
        in1(1) => U1_AC_out_2,
        out1 => S2099
    );
nand_n_913: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1940,
        in1(1) => S1932,
        out1 => S2100
    );
nand_n_914: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2099,
        in1(1) => S2097,
        out1 => S2101
    );
nand_n_915: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2018,
        in1(1) => U1_OF_out_2,
        out1 => S2102
    );
nand_n_916: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2102,
        in1(1) => S2015,
        out1 => S2103
    );
nor_n_444: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2103,
        in1(1) => U1_selMEM_LGU,
        out1 => S2104
    );
nor_n_445: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_dataBus_14,
        in1(1) => S1842,
        out1 => S2105
    );
nor_n_446: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2105,
        in1(1) => S2104,
        out1 => S2106
    );
notg_140: ENTITY WORK.notg
    PORT MAP (
        in1 => S2106,
        out1 => S2107
    );
nor_n_447: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2107,
        in1(1) => S2046,
        out1 => S2108
    );
nand_n_917: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2108,
        in1(1) => U1_AC_out_0,
        out1 => S2109
    );
nor_n_448: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2030,
        in1(1) => U1_AC_out_2,
        out1 => S2110
    );
nand_n_918: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2029,
        in1(1) => S1932,
        out1 => S2111
    );
nand_n_919: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2018,
        in1(1) => U1_OF_out_1,
        out1 => S2112
    );
nand_n_920: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2112,
        in1(1) => S2015,
        out1 => S2113
    );
nor_n_449: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2113,
        in1(1) => U1_selMEM_LGU,
        out1 => S2114
    );
nor_n_450: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_dataBus_13,
        in1(1) => S1842,
        out1 => S2115
    );
nor_n_451: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2115,
        in1(1) => S2114,
        out1 => S2116
    );
notg_141: ENTITY WORK.notg
    PORT MAP (
        in1 => S2116,
        out1 => S2117
    );
nor_n_452: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2117,
        in1(1) => S2046,
        out1 => S2118
    );
nand_n_921: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2116,
        in1(1) => S2045,
        out1 => S2119
    );
nand_n_922: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2118,
        in1(1) => S1917,
        out1 => S2120
    );
nand_n_923: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2018,
        in1(1) => U1_OF_out_0,
        out1 => S2121
    );
nand_n_924: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2121,
        in1(1) => S2015,
        out1 => S2122
    );
nor_n_453: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2122,
        in1(1) => U1_selMEM_LGU,
        out1 => S2123
    );
nor_n_454: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_dataBus_12,
        in1(1) => S1842,
        out1 => S2124
    );
nor_n_455: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2124,
        in1(1) => S2123,
        out1 => S2125
    );
notg_142: ENTITY WORK.notg
    PORT MAP (
        in1 => S2125,
        out1 => S2126
    );
nor_n_456: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2126,
        in1(1) => S2046,
        out1 => S2127
    );
nand_n_925: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2125,
        in1(1) => S2045,
        out1 => S2128
    );
nand_n_926: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2127,
        in1(1) => U1_AC_out_0,
        out1 => S2129
    );
nand_n_927: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2129,
        in1(1) => S2120,
        out1 => S2130
    );
nor_n_457: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2109,
        in1(1) => U1_AC_out_1,
        out1 => S2131
    );
nand_n_928: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2130,
        in1(1) => U1_AC_out_1,
        out1 => S2132
    );
nand_n_929: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2132,
        in1(1) => S2098,
        out1 => S2133
    );
nor_n_458: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2133,
        in1(1) => S2131,
        out1 => S2134
    );
nor_n_459: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2134,
        in1(1) => S2111,
        out1 => S2135
    );
nor_n_460: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2135,
        in1(1) => S2093,
        out1 => S2136
    );
nand_n_930: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2136,
        in1(1) => S2101,
        out1 => S2137
    );
nor_n_461: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_SE12bits,
        in1(1) => U1_conOF,
        out1 => S2138
    );
notg_143: ENTITY WORK.notg
    PORT MAP (
        in1 => S2138,
        out1 => S2139
    );
nor_n_462: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2139,
        in1(1) => U1_SE4bits,
        out1 => S2140
    );
nand_n_931: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2138,
        in1(1) => S1832,
        out1 => S2141
    );
nor_n_463: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2140,
        in1(1) => S1813,
        out1 => S2142
    );
nand_n_932: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2141,
        in1(1) => U1_IR_out_3,
        out1 => S2143
    );
nand_n_933: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_dataBus_3,
        in1(1) => U1_selMEM_LGU,
        out1 => S2144
    );
notg_144: ENTITY WORK.notg
    PORT MAP (
        in1 => S2144,
        out1 => S2145
    );
nor_n_464: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2143,
        in1(1) => U1_selMEM_LGU,
        out1 => S2146
    );
notg_145: ENTITY WORK.notg
    PORT MAP (
        in1 => S2146,
        out1 => S2147
    );
nand_n_934: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2147,
        in1(1) => S2144,
        out1 => S2148
    );
nor_n_465: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2146,
        in1(1) => S2145,
        out1 => S2149
    );
nor_n_466: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2149,
        in1(1) => S2046,
        out1 => S2150
    );
nand_n_935: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2148,
        in1(1) => S2045,
        out1 => S2151
    );
nand_n_936: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2151,
        in1(1) => S1917,
        out1 => S2152
    );
nor_n_467: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2140,
        in1(1) => S1955,
        out1 => S2153
    );
nand_n_937: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2141,
        in1(1) => U1_IR_out_2,
        out1 => S2154
    );
nand_n_938: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_dataBus_2,
        in1(1) => U1_selMEM_LGU,
        out1 => S2155
    );
notg_146: ENTITY WORK.notg
    PORT MAP (
        in1 => S2155,
        out1 => S2156
    );
nor_n_468: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2154,
        in1(1) => U1_selMEM_LGU,
        out1 => S2157
    );
notg_147: ENTITY WORK.notg
    PORT MAP (
        in1 => S2157,
        out1 => S2158
    );
nand_n_939: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2158,
        in1(1) => S2155,
        out1 => S2159
    );
nor_n_469: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2157,
        in1(1) => S2156,
        out1 => S2160
    );
nor_n_470: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2160,
        in1(1) => S2046,
        out1 => S2161
    );
nand_n_940: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2159,
        in1(1) => S2045,
        out1 => S2162
    );
nand_n_941: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2162,
        in1(1) => U1_AC_out_0,
        out1 => S2163
    );
nand_n_942: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2163,
        in1(1) => S2152,
        out1 => S2164
    );
notg_148: ENTITY WORK.notg
    PORT MAP (
        in1 => S2164,
        out1 => S2165
    );
nor_n_471: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2165,
        in1(1) => U1_AC_out_1,
        out1 => S2166
    );
nand_n_943: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2164,
        in1(1) => S1925,
        out1 => S2167
    );
nand_n_944: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2141,
        in1(1) => U1_IR_out_1,
        out1 => S2168
    );
nand_n_945: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_dataBus_1,
        in1(1) => U1_selMEM_LGU,
        out1 => S2169
    );
notg_149: ENTITY WORK.notg
    PORT MAP (
        in1 => S2169,
        out1 => S2170
    );
nor_n_472: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2168,
        in1(1) => U1_selMEM_LGU,
        out1 => S2171
    );
notg_150: ENTITY WORK.notg
    PORT MAP (
        in1 => S2171,
        out1 => S2172
    );
nand_n_946: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2172,
        in1(1) => S2169,
        out1 => S2173
    );
nor_n_473: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2171,
        in1(1) => S2170,
        out1 => S2174
    );
nor_n_474: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2174,
        in1(1) => S2046,
        out1 => S2175
    );
notg_151: ENTITY WORK.notg
    PORT MAP (
        in1 => S2175,
        out1 => S2176
    );
nand_n_947: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2176,
        in1(1) => S1917,
        out1 => S2177
    );
nand_n_948: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_dataBus_0,
        in1(1) => U1_selMEM_LGU,
        out1 => S2178
    );
notg_152: ENTITY WORK.notg
    PORT MAP (
        in1 => S2178,
        out1 => S2179
    );
nor_n_475: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2140,
        in1(1) => S1957,
        out1 => S2180
    );
nand_n_949: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2141,
        in1(1) => U1_IR_out_0,
        out1 => S2181
    );
nor_n_476: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2181,
        in1(1) => U1_selMEM_LGU,
        out1 => S2182
    );
notg_153: ENTITY WORK.notg
    PORT MAP (
        in1 => S2182,
        out1 => S2183
    );
nor_n_477: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2182,
        in1(1) => S2179,
        out1 => S2184
    );
nand_n_950: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2183,
        in1(1) => S2178,
        out1 => S2185
    );
nand_n_951: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2185,
        in1(1) => S2045,
        out1 => S2186
    );
notg_154: ENTITY WORK.notg
    PORT MAP (
        in1 => S2186,
        out1 => S2187
    );
nand_n_952: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2186,
        in1(1) => U1_AC_out_0,
        out1 => S2188
    );
nand_n_953: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2188,
        in1(1) => S2177,
        out1 => S2189
    );
nand_n_954: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2189,
        in1(1) => U1_AC_out_1,
        out1 => S2190
    );
notg_155: ENTITY WORK.notg
    PORT MAP (
        in1 => S2190,
        out1 => S2191
    );
nor_n_478: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2191,
        in1(1) => S2166,
        out1 => S2192
    );
nand_n_955: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2190,
        in1(1) => S2167,
        out1 => S2193
    );
nand_n_956: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2048,
        in1(1) => U1_IR_out_7,
        out1 => S2194
    );
nand_n_957: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2194,
        in1(1) => S2012,
        out1 => S2195
    );
nor_n_479: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2195,
        in1(1) => U1_selMEM_LGU,
        out1 => S2196
    );
nor_n_480: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_dataBus_7,
        in1(1) => S1842,
        out1 => S2197
    );
nor_n_481: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2197,
        in1(1) => S2196,
        out1 => S2198
    );
notg_156: ENTITY WORK.notg
    PORT MAP (
        in1 => S2198,
        out1 => S2199
    );
nor_n_482: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2199,
        in1(1) => S2046,
        out1 => S2200
    );
nand_n_958: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2198,
        in1(1) => S2045,
        out1 => S2201
    );
nor_n_483: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2200,
        in1(1) => U1_AC_out_0,
        out1 => S2202
    );
nand_n_959: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2048,
        in1(1) => U1_IR_out_6,
        out1 => S2203
    );
nand_n_960: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2203,
        in1(1) => S2012,
        out1 => S2204
    );
nor_n_484: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2204,
        in1(1) => U1_selMEM_LGU,
        out1 => S2205
    );
nor_n_485: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_dataBus_6,
        in1(1) => S1842,
        out1 => S2206
    );
nor_n_486: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2206,
        in1(1) => S2205,
        out1 => S2207
    );
notg_157: ENTITY WORK.notg
    PORT MAP (
        in1 => S2207,
        out1 => S2208
    );
nor_n_487: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2208,
        in1(1) => S2046,
        out1 => S2209
    );
nand_n_961: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2207,
        in1(1) => S2045,
        out1 => S2210
    );
nor_n_488: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2209,
        in1(1) => S1917,
        out1 => S2211
    );
nor_n_489: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2211,
        in1(1) => S2202,
        out1 => S2212
    );
nor_n_490: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2212,
        in1(1) => U1_AC_out_1,
        out1 => S2213
    );
nand_n_962: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2048,
        in1(1) => U1_IR_out_5,
        out1 => S2214
    );
nand_n_963: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2214,
        in1(1) => S2012,
        out1 => S2215
    );
nor_n_491: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2215,
        in1(1) => U1_selMEM_LGU,
        out1 => S2216
    );
nor_n_492: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_dataBus_5,
        in1(1) => S1842,
        out1 => S2217
    );
nor_n_493: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2217,
        in1(1) => S2216,
        out1 => S2218
    );
notg_158: ENTITY WORK.notg
    PORT MAP (
        in1 => S2218,
        out1 => S2219
    );
nor_n_494: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2219,
        in1(1) => S2046,
        out1 => S2220
    );
nand_n_964: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2218,
        in1(1) => S2045,
        out1 => S2221
    );
nor_n_495: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2220,
        in1(1) => U1_AC_out_0,
        out1 => S2222
    );
notg_159: ENTITY WORK.notg
    PORT MAP (
        in1 => S2222,
        out1 => S2223
    );
nor_n_496: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2047,
        in1(1) => S1952,
        out1 => S2224
    );
nand_n_965: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2048,
        in1(1) => U1_IR_out_4,
        out1 => S2225
    );
nor_n_497: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2224,
        in1(1) => S2011,
        out1 => S2226
    );
nand_n_966: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2225,
        in1(1) => S2012,
        out1 => S2227
    );
nand_n_967: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_dataBus_4,
        in1(1) => U1_selMEM_LGU,
        out1 => S2228
    );
notg_160: ENTITY WORK.notg
    PORT MAP (
        in1 => S2228,
        out1 => S2229
    );
nor_n_498: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2226,
        in1(1) => U1_selMEM_LGU,
        out1 => S2230
    );
nand_n_968: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2227,
        in1(1) => S1842,
        out1 => S2231
    );
nand_n_969: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2231,
        in1(1) => S2228,
        out1 => S2232
    );
nor_n_499: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2230,
        in1(1) => S2229,
        out1 => S2233
    );
nor_n_500: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2233,
        in1(1) => S2046,
        out1 => S2234
    );
nand_n_970: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2232,
        in1(1) => S2045,
        out1 => S2235
    );
nor_n_501: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2234,
        in1(1) => S1917,
        out1 => S2236
    );
nand_n_971: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2235,
        in1(1) => U1_AC_out_0,
        out1 => S2237
    );
nor_n_502: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2236,
        in1(1) => S2222,
        out1 => S2238
    );
nand_n_972: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2237,
        in1(1) => S2223,
        out1 => S2239
    );
nand_n_973: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2239,
        in1(1) => U1_AC_out_1,
        out1 => S2240
    );
notg_161: ENTITY WORK.notg
    PORT MAP (
        in1 => S2240,
        out1 => S2241
    );
nor_n_503: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2241,
        in1(1) => S2213,
        out1 => S2242
    );
nor_n_504: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2242,
        in1(1) => U1_AC_out_2,
        out1 => S2243
    );
nand_n_974: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2193,
        in1(1) => U1_AC_out_2,
        out1 => S2244
    );
nand_n_975: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2244,
        in1(1) => S2029,
        out1 => S2245
    );
nor_n_505: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2245,
        in1(1) => S2243,
        out1 => S2246
    );
nor_n_506: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2246,
        in1(1) => S1939,
        out1 => S2247
    );
nor_n_507: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_NOT,
        in1(1) => U1_AC_out_4,
        out1 => S2248
    );
nand_n_976: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1959,
        in1(1) => S1852,
        out1 => S2249
    );
nor_n_508: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2249,
        in1(1) => S2247,
        out1 => S2250
    );
nand_n_977: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2250,
        in1(1) => S2137,
        out1 => S2251
    );
nand_n_978: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2251,
        in1(1) => S2028,
        out1 => S2252
    );
nand_n_979: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2252,
        in1(1) => S2026,
        out1 => S2253
    );
notg_162: ENTITY WORK.notg
    PORT MAP (
        in1 => S2253,
        out1 => U1_LGU_out_15
    );
nand_n_980: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_PC_out_1,
        in1(1) => U1_PC_out_0,
        out1 => S2254
    );
notg_163: ENTITY WORK.notg
    PORT MAP (
        in1 => S2254,
        out1 => S0
    );
nand_n_981: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_PC_out_2,
        in1(1) => U1_PC_out_1,
        out1 => S2255
    );
notg_164: ENTITY WORK.notg
    PORT MAP (
        in1 => S2255,
        out1 => S1
    );
nor_n_509: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2254,
        in1(1) => S1970,
        out1 => S2
    );
nand_n_982: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1,
        in1(1) => U1_PC_out_3,
        out1 => S2256
    );
notg_165: ENTITY WORK.notg
    PORT MAP (
        in1 => S2256,
        out1 => S3
    );
nor_n_510: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2256,
        in1(1) => S1966,
        out1 => S4
    );
nand_n_983: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3,
        in1(1) => U1_PC_out_4,
        out1 => S2257
    );
notg_166: ENTITY WORK.notg
    PORT MAP (
        in1 => S2257,
        out1 => S5
    );
nor_n_511: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2257,
        in1(1) => S1966,
        out1 => S6
    );
nand_n_984: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5,
        in1(1) => U1_PC_out_5,
        out1 => S2258
    );
notg_167: ENTITY WORK.notg
    PORT MAP (
        in1 => S2258,
        out1 => S7
    );
nor_n_512: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2258,
        in1(1) => S1966,
        out1 => S8
    );
nand_n_985: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S7,
        in1(1) => U1_PC_out_6,
        out1 => S2259
    );
notg_168: ENTITY WORK.notg
    PORT MAP (
        in1 => S2259,
        out1 => S9
    );
nor_n_513: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2259,
        in1(1) => S1966,
        out1 => S10
    );
nand_n_986: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S9,
        in1(1) => U1_PC_out_7,
        out1 => S2260
    );
notg_169: ENTITY WORK.notg
    PORT MAP (
        in1 => S2260,
        out1 => S11
    );
nor_n_514: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2260,
        in1(1) => S1966,
        out1 => S12
    );
nand_n_987: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S11,
        in1(1) => U1_PC_out_8,
        out1 => S2261
    );
notg_170: ENTITY WORK.notg
    PORT MAP (
        in1 => S2261,
        out1 => S13
    );
nor_n_515: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2261,
        in1(1) => S1966,
        out1 => S14
    );
nand_n_988: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S13,
        in1(1) => U1_PC_out_9,
        out1 => S2262
    );
notg_171: ENTITY WORK.notg
    PORT MAP (
        in1 => S2262,
        out1 => S15
    );
nor_n_516: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2262,
        in1(1) => S1966,
        out1 => S16
    );
nand_n_989: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S15,
        in1(1) => U1_PC_out_10,
        out1 => S2263
    );
notg_172: ENTITY WORK.notg
    PORT MAP (
        in1 => S2263,
        out1 => S17
    );
nor_n_517: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2263,
        in1(1) => S1966,
        out1 => S18
    );
nor_n_518: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2263,
        in1(1) => S1988,
        out1 => S19
    );
nand_n_990: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S19,
        in1(1) => U1_PC_out_0,
        out1 => S2264
    );
notg_173: ENTITY WORK.notg
    PORT MAP (
        in1 => S2264,
        out1 => S20
    );
nand_n_991: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S19,
        in1(1) => U1_PC_out_12,
        out1 => S2265
    );
notg_174: ENTITY WORK.notg
    PORT MAP (
        in1 => S2265,
        out1 => S21
    );
nor_n_519: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2264,
        in1(1) => S1961,
        out1 => S22
    );
nand_n_992: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S21,
        in1(1) => U1_PC_out_13,
        out1 => S2266
    );
notg_175: ENTITY WORK.notg
    PORT MAP (
        in1 => S2266,
        out1 => S23
    );
nand_n_993: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S23,
        in1(1) => U1_PC_out_0,
        out1 => S2267
    );
notg_176: ENTITY WORK.notg
    PORT MAP (
        in1 => S2267,
        out1 => S24
    );
nor_n_520: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2266,
        in1(1) => S1964,
        out1 => S25
    );
nor_n_521: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2267,
        in1(1) => S1964,
        out1 => S26
    );
nand_n_994: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2023,
        in1(1) => U1_selMO_ARU,
        out1 => S2268
    );
nand_n_995: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2025,
        in1(1) => U1_selMO_ARU,
        out1 => S2269
    );
notg_177: ENTITY WORK.notg
    PORT MAP (
        in1 => S2269,
        out1 => S2270
    );
nor_n_522: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2219,
        in1(1) => S1993,
        out1 => S2271
    );
nand_n_996: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2218,
        in1(1) => U1_selMO_ARU,
        out1 => S2272
    );
nand_n_997: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2271,
        in1(1) => U1_AC_out_6,
        out1 => S2273
    );
nor_n_523: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2233,
        in1(1) => S1993,
        out1 => S2274
    );
nand_n_998: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2232,
        in1(1) => U1_selMO_ARU,
        out1 => S2275
    );
nand_n_999: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2274,
        in1(1) => U1_AC_out_7,
        out1 => S2276
    );
nor_n_524: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2272,
        in1(1) => S1882,
        out1 => S2277
    );
nand_n_1000: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2271,
        in1(1) => U1_AC_out_7,
        out1 => S2278
    );
nor_n_525: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2275,
        in1(1) => S1862,
        out1 => S2279
    );
nand_n_1001: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2274,
        in1(1) => U1_AC_out_6,
        out1 => S2280
    );
nor_n_526: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2280,
        in1(1) => S2278,
        out1 => S2281
    );
nand_n_1002: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2279,
        in1(1) => S2277,
        out1 => S2282
    );
nor_n_527: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2208,
        in1(1) => S1993,
        out1 => S2283
    );
nand_n_1003: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2207,
        in1(1) => U1_selMO_ARU,
        out1 => S2284
    );
nand_n_1004: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2283,
        in1(1) => U1_AC_out_5,
        out1 => S2285
    );
notg_178: ENTITY WORK.notg
    PORT MAP (
        in1 => S2285,
        out1 => S2286
    );
nand_n_1005: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2276,
        in1(1) => S2273,
        out1 => S2287
    );
nand_n_1006: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2287,
        in1(1) => S2282,
        out1 => S2288
    );
notg_179: ENTITY WORK.notg
    PORT MAP (
        in1 => S2288,
        out1 => S2289
    );
nor_n_528: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2288,
        in1(1) => S2285,
        out1 => S2290
    );
nand_n_1007: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2289,
        in1(1) => S2286,
        out1 => S2291
    );
nor_n_529: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2290,
        in1(1) => S2281,
        out1 => S2292
    );
nand_n_1008: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2291,
        in1(1) => S2282,
        out1 => S2293
    );
nand_n_1009: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2207,
        in1(1) => U1_AC_out_6,
        out1 => S2294
    );
notg_180: ENTITY WORK.notg
    PORT MAP (
        in1 => S2294,
        out1 => S2295
    );
nor_n_530: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2284,
        in1(1) => S1862,
        out1 => S2296
    );
nand_n_1010: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2283,
        in1(1) => U1_AC_out_6,
        out1 => S2297
    );
nand_n_1011: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2283,
        in1(1) => U1_AC_out_7,
        out1 => S2298
    );
nor_n_531: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2294,
        in1(1) => S2278,
        out1 => S2299
    );
notg_181: ENTITY WORK.notg
    PORT MAP (
        in1 => S2299,
        out1 => S2300
    );
nor_n_532: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2296,
        in1(1) => S2277,
        out1 => S2301
    );
nand_n_1012: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2297,
        in1(1) => S2278,
        out1 => S2302
    );
nor_n_533: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2301,
        in1(1) => S2299,
        out1 => S2303
    );
nand_n_1013: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2302,
        in1(1) => S2300,
        out1 => S2304
    );
nor_n_534: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2199,
        in1(1) => S1993,
        out1 => S2305
    );
nand_n_1014: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2198,
        in1(1) => U1_selMO_ARU,
        out1 => S2306
    );
nor_n_535: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2306,
        in1(1) => S1872,
        out1 => S2307
    );
nand_n_1015: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2305,
        in1(1) => U1_AC_out_5,
        out1 => S2308
    );
nor_n_536: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2308,
        in1(1) => S2304,
        out1 => S2309
    );
notg_182: ENTITY WORK.notg
    PORT MAP (
        in1 => S2309,
        out1 => S2310
    );
nor_n_537: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2307,
        in1(1) => S2303,
        out1 => S2311
    );
nand_n_1016: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2308,
        in1(1) => S2304,
        out1 => S2312
    );
nor_n_538: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2311,
        in1(1) => S2309,
        out1 => S2313
    );
nand_n_1017: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2312,
        in1(1) => S2310,
        out1 => S2314
    );
nor_n_539: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2314,
        in1(1) => S2292,
        out1 => S2315
    );
notg_183: ENTITY WORK.notg
    PORT MAP (
        in1 => S2315,
        out1 => S2316
    );
nor_n_540: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2313,
        in1(1) => S2293,
        out1 => S2317
    );
nand_n_1018: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2314,
        in1(1) => S2292,
        out1 => S2318
    );
nor_n_541: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2317,
        in1(1) => S2315,
        out1 => S2319
    );
nand_n_1019: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2318,
        in1(1) => S2316,
        out1 => S2320
    );
nor_n_542: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2149,
        in1(1) => S1993,
        out1 => S2321
    );
nand_n_1020: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2148,
        in1(1) => U1_selMO_ARU,
        out1 => S2322
    );
nor_n_543: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2322,
        in1(1) => S1882,
        out1 => S2323
    );
nand_n_1021: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2321,
        in1(1) => U1_AC_out_7,
        out1 => S2324
    );
nor_n_544: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2322,
        in1(1) => S1862,
        out1 => S2325
    );
nand_n_1022: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2321,
        in1(1) => U1_AC_out_6,
        out1 => S2326
    );
nor_n_545: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2324,
        in1(1) => S2280,
        out1 => S2327
    );
nand_n_1023: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2323,
        in1(1) => S2279,
        out1 => S2328
    );
nand_n_1024: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2218,
        in1(1) => U1_AC_out_5,
        out1 => S2329
    );
nor_n_546: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2272,
        in1(1) => S1872,
        out1 => S2330
    );
nand_n_1025: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2271,
        in1(1) => U1_AC_out_5,
        out1 => S2331
    );
nor_n_547: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2323,
        in1(1) => S2279,
        out1 => S2332
    );
nand_n_1026: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2324,
        in1(1) => S2280,
        out1 => S2333
    );
nor_n_548: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2332,
        in1(1) => S2327,
        out1 => S2334
    );
nand_n_1027: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2333,
        in1(1) => S2328,
        out1 => S2335
    );
nor_n_549: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2335,
        in1(1) => S2331,
        out1 => S2336
    );
nand_n_1028: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2334,
        in1(1) => S2330,
        out1 => S2337
    );
nor_n_550: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2336,
        in1(1) => S2327,
        out1 => S2338
    );
nand_n_1029: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2337,
        in1(1) => S2328,
        out1 => S2339
    );
nand_n_1030: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2288,
        in1(1) => S2285,
        out1 => S2340
    );
notg_184: ENTITY WORK.notg
    PORT MAP (
        in1 => S2340,
        out1 => S2341
    );
nor_n_551: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2341,
        in1(1) => S2290,
        out1 => S2342
    );
nand_n_1031: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2340,
        in1(1) => S2291,
        out1 => S2343
    );
nor_n_552: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2343,
        in1(1) => S2338,
        out1 => S2344
    );
nand_n_1032: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2342,
        in1(1) => S2339,
        out1 => S2345
    );
nor_n_553: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2306,
        in1(1) => S1852,
        out1 => S2346
    );
nand_n_1033: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2305,
        in1(1) => U1_AC_out_4,
        out1 => S2347
    );
nor_n_554: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2342,
        in1(1) => S2339,
        out1 => S2348
    );
nand_n_1034: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2343,
        in1(1) => S2338,
        out1 => S2349
    );
nor_n_555: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2348,
        in1(1) => S2344,
        out1 => S2350
    );
nand_n_1035: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2349,
        in1(1) => S2345,
        out1 => S2351
    );
nor_n_556: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2351,
        in1(1) => S2347,
        out1 => S2352
    );
nand_n_1036: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2350,
        in1(1) => S2346,
        out1 => S2353
    );
nor_n_557: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2352,
        in1(1) => S2344,
        out1 => S2354
    );
nand_n_1037: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2353,
        in1(1) => S2345,
        out1 => S2355
    );
nor_n_558: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2354,
        in1(1) => S2320,
        out1 => S2356
    );
nor_n_559: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2355,
        in1(1) => S2319,
        out1 => S2357
    );
nor_n_560: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2357,
        in1(1) => S2356,
        out1 => S2358
    );
notg_185: ENTITY WORK.notg
    PORT MAP (
        in1 => S2358,
        out1 => S2359
    );
nor_n_561: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2160,
        in1(1) => S1993,
        out1 => S2360
    );
nand_n_1038: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2159,
        in1(1) => U1_selMO_ARU,
        out1 => S2361
    );
nor_n_562: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2361,
        in1(1) => S1882,
        out1 => S2362
    );
nand_n_1039: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2360,
        in1(1) => U1_AC_out_7,
        out1 => S2363
    );
nand_n_1040: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2360,
        in1(1) => U1_AC_out_6,
        out1 => S2364
    );
nor_n_563: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2363,
        in1(1) => S2326,
        out1 => S2365
    );
nand_n_1041: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2362,
        in1(1) => S2325,
        out1 => S2366
    );
nor_n_564: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2275,
        in1(1) => S1872,
        out1 => S2367
    );
nand_n_1042: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2274,
        in1(1) => U1_AC_out_5,
        out1 => S2368
    );
nor_n_565: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2362,
        in1(1) => S2325,
        out1 => S2369
    );
nand_n_1043: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2363,
        in1(1) => S2326,
        out1 => S2370
    );
nor_n_566: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2369,
        in1(1) => S2365,
        out1 => S2371
    );
nand_n_1044: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2370,
        in1(1) => S2366,
        out1 => S2372
    );
nor_n_567: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2372,
        in1(1) => S2368,
        out1 => S2373
    );
nand_n_1045: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2371,
        in1(1) => S2367,
        out1 => S2374
    );
nor_n_568: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2373,
        in1(1) => S2365,
        out1 => S2375
    );
nand_n_1046: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2374,
        in1(1) => S2366,
        out1 => S2376
    );
nor_n_569: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2334,
        in1(1) => S2330,
        out1 => S2377
    );
nand_n_1047: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2335,
        in1(1) => S2331,
        out1 => S2378
    );
nor_n_570: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2377,
        in1(1) => S2336,
        out1 => S2379
    );
nand_n_1048: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2378,
        in1(1) => S2337,
        out1 => S2380
    );
nor_n_571: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2380,
        in1(1) => S2375,
        out1 => S2381
    );
nand_n_1049: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2379,
        in1(1) => S2376,
        out1 => S2382
    );
nor_n_572: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2379,
        in1(1) => S2376,
        out1 => S2383
    );
nand_n_1050: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2380,
        in1(1) => S2375,
        out1 => S2384
    );
nor_n_573: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2383,
        in1(1) => S2381,
        out1 => S2385
    );
nand_n_1051: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2384,
        in1(1) => S2382,
        out1 => S2386
    );
nand_n_1052: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2305,
        in1(1) => U1_AC_out_3,
        out1 => S2387
    );
nand_n_1053: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2283,
        in1(1) => U1_AC_out_4,
        out1 => S2388
    );
nor_n_574: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2284,
        in1(1) => S1939,
        out1 => S2389
    );
nand_n_1054: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2283,
        in1(1) => U1_AC_out_3,
        out1 => S2390
    );
nor_n_575: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2390,
        in1(1) => S2347,
        out1 => S2391
    );
nand_n_1055: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2389,
        in1(1) => S2346,
        out1 => S2392
    );
nand_n_1056: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2388,
        in1(1) => S2387,
        out1 => S2393
    );
notg_186: ENTITY WORK.notg
    PORT MAP (
        in1 => S2393,
        out1 => S2394
    );
nor_n_576: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2394,
        in1(1) => S2391,
        out1 => S2395
    );
nand_n_1057: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2393,
        in1(1) => S2392,
        out1 => S2396
    );
nor_n_577: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2396,
        in1(1) => S2386,
        out1 => S2397
    );
nand_n_1058: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2395,
        in1(1) => S2385,
        out1 => S2398
    );
nor_n_578: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2397,
        in1(1) => S2381,
        out1 => S2399
    );
nand_n_1059: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2398,
        in1(1) => S2382,
        out1 => S2400
    );
nor_n_579: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2350,
        in1(1) => S2346,
        out1 => S2401
    );
nand_n_1060: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2351,
        in1(1) => S2347,
        out1 => S2402
    );
nor_n_580: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2401,
        in1(1) => S2352,
        out1 => S2403
    );
nand_n_1061: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2402,
        in1(1) => S2353,
        out1 => S2404
    );
nor_n_581: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2404,
        in1(1) => S2399,
        out1 => S2405
    );
nand_n_1062: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2403,
        in1(1) => S2400,
        out1 => S2406
    );
nor_n_582: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2403,
        in1(1) => S2400,
        out1 => S2407
    );
nand_n_1063: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2404,
        in1(1) => S2399,
        out1 => S2408
    );
nor_n_583: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2407,
        in1(1) => S2405,
        out1 => S2409
    );
nand_n_1064: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2408,
        in1(1) => S2406,
        out1 => S2410
    );
nor_n_584: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2410,
        in1(1) => S2392,
        out1 => S2411
    );
nand_n_1065: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2409,
        in1(1) => S2391,
        out1 => S2412
    );
nor_n_585: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2411,
        in1(1) => S2405,
        out1 => S2413
    );
nand_n_1066: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2412,
        in1(1) => S2406,
        out1 => S2414
    );
nand_n_1067: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2414,
        in1(1) => S2358,
        out1 => S2415
    );
notg_187: ENTITY WORK.notg
    PORT MAP (
        in1 => S2415,
        out1 => S2416
    );
nor_n_586: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2309,
        in1(1) => S2299,
        out1 => S2417
    );
nand_n_1068: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2198,
        in1(1) => U1_AC_out_7,
        out1 => S2418
    );
nor_n_587: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2306,
        in1(1) => S1882,
        out1 => S2419
    );
nand_n_1069: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2419,
        in1(1) => S2295,
        out1 => S2420
    );
nand_n_1070: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2305,
        in1(1) => U1_AC_out_6,
        out1 => S2421
    );
nand_n_1071: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2421,
        in1(1) => S2298,
        out1 => S2422
    );
nand_n_1072: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2422,
        in1(1) => S2420,
        out1 => S2423
    );
nor_n_588: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2423,
        in1(1) => S2417,
        out1 => S2424
    );
notg_188: ENTITY WORK.notg
    PORT MAP (
        in1 => S2424,
        out1 => S2425
    );
nand_n_1073: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2423,
        in1(1) => S2417,
        out1 => S2426
    );
nand_n_1074: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2426,
        in1(1) => S2425,
        out1 => S2427
    );
nor_n_589: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2356,
        in1(1) => S2315,
        out1 => S2428
    );
nor_n_590: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2428,
        in1(1) => S2427,
        out1 => S2429
    );
notg_189: ENTITY WORK.notg
    PORT MAP (
        in1 => S2429,
        out1 => S2430
    );
nand_n_1075: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2428,
        in1(1) => S2427,
        out1 => S2431
    );
nand_n_1076: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2431,
        in1(1) => S2430,
        out1 => S2432
    );
notg_190: ENTITY WORK.notg
    PORT MAP (
        in1 => S2432,
        out1 => S2433
    );
nand_n_1077: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2433,
        in1(1) => S2416,
        out1 => S2434
    );
notg_191: ENTITY WORK.notg
    PORT MAP (
        in1 => S2434,
        out1 => S2435
    );
nand_n_1078: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2432,
        in1(1) => S2415,
        out1 => S2436
    );
nand_n_1079: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2436,
        in1(1) => S2434,
        out1 => S2437
    );
notg_192: ENTITY WORK.notg
    PORT MAP (
        in1 => S2437,
        out1 => S2438
    );
nand_n_1080: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2413,
        in1(1) => S2359,
        out1 => S2439
    );
nand_n_1081: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2439,
        in1(1) => S2415,
        out1 => S2440
    );
notg_193: ENTITY WORK.notg
    PORT MAP (
        in1 => S2440,
        out1 => S2441
    );
nor_n_591: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2174,
        in1(1) => S1993,
        out1 => S2442
    );
nand_n_1082: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2173,
        in1(1) => U1_selMO_ARU,
        out1 => S2443
    );
nand_n_1083: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2442,
        in1(1) => U1_AC_out_7,
        out1 => S2444
    );
nor_n_592: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2443,
        in1(1) => S1862,
        out1 => S2445
    );
nand_n_1084: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2442,
        in1(1) => U1_AC_out_6,
        out1 => S2446
    );
nor_n_593: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2446,
        in1(1) => S2363,
        out1 => S2447
    );
nand_n_1085: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2445,
        in1(1) => S2362,
        out1 => S2448
    );
nand_n_1086: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2321,
        in1(1) => U1_AC_out_5,
        out1 => S2449
    );
notg_194: ENTITY WORK.notg
    PORT MAP (
        in1 => S2449,
        out1 => S2450
    );
nand_n_1087: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2444,
        in1(1) => S2364,
        out1 => S2451
    );
nand_n_1088: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2451,
        in1(1) => S2448,
        out1 => S2452
    );
notg_195: ENTITY WORK.notg
    PORT MAP (
        in1 => S2452,
        out1 => S2453
    );
nor_n_594: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2452,
        in1(1) => S2449,
        out1 => S2454
    );
nand_n_1089: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2453,
        in1(1) => S2450,
        out1 => S2455
    );
nor_n_595: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2454,
        in1(1) => S2447,
        out1 => S2456
    );
nand_n_1090: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2455,
        in1(1) => S2448,
        out1 => S2457
    );
nor_n_596: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2371,
        in1(1) => S2367,
        out1 => S2458
    );
nand_n_1091: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2372,
        in1(1) => S2368,
        out1 => S2459
    );
nor_n_597: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2458,
        in1(1) => S2373,
        out1 => S2460
    );
nand_n_1092: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2459,
        in1(1) => S2374,
        out1 => S2461
    );
nor_n_598: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2461,
        in1(1) => S2456,
        out1 => S2462
    );
nand_n_1093: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2460,
        in1(1) => S2457,
        out1 => S2463
    );
nor_n_599: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2460,
        in1(1) => S2457,
        out1 => S2464
    );
nand_n_1094: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2461,
        in1(1) => S2456,
        out1 => S2465
    );
nor_n_600: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2464,
        in1(1) => S2462,
        out1 => S2466
    );
nand_n_1095: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2465,
        in1(1) => S2463,
        out1 => S2467
    );
nor_n_601: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2306,
        in1(1) => S1932,
        out1 => S2468
    );
nand_n_1096: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2305,
        in1(1) => U1_AC_out_2,
        out1 => S2469
    );
nor_n_602: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2272,
        in1(1) => S1852,
        out1 => S2470
    );
nand_n_1097: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2271,
        in1(1) => U1_AC_out_4,
        out1 => S2471
    );
nor_n_603: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2272,
        in1(1) => S1939,
        out1 => S2472
    );
nand_n_1098: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2271,
        in1(1) => U1_AC_out_3,
        out1 => S2473
    );
nor_n_604: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2471,
        in1(1) => S2390,
        out1 => S2474
    );
nand_n_1099: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2470,
        in1(1) => S2389,
        out1 => S2475
    );
nor_n_605: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2470,
        in1(1) => S2389,
        out1 => S2476
    );
nand_n_1100: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2471,
        in1(1) => S2390,
        out1 => S2477
    );
nor_n_606: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2476,
        in1(1) => S2474,
        out1 => S2478
    );
nand_n_1101: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2477,
        in1(1) => S2475,
        out1 => S2479
    );
nor_n_607: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2479,
        in1(1) => S2469,
        out1 => S2480
    );
nand_n_1102: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2478,
        in1(1) => S2468,
        out1 => S2481
    );
nor_n_608: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2478,
        in1(1) => S2468,
        out1 => S2482
    );
nand_n_1103: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2479,
        in1(1) => S2469,
        out1 => S2483
    );
nor_n_609: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2482,
        in1(1) => S2480,
        out1 => S2484
    );
nand_n_1104: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2483,
        in1(1) => S2481,
        out1 => S2485
    );
nor_n_610: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2485,
        in1(1) => S2467,
        out1 => S2486
    );
nand_n_1105: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2484,
        in1(1) => S2466,
        out1 => S2487
    );
nor_n_611: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2486,
        in1(1) => S2462,
        out1 => S2488
    );
nand_n_1106: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2487,
        in1(1) => S2463,
        out1 => S2489
    );
nor_n_612: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2395,
        in1(1) => S2385,
        out1 => S2490
    );
nand_n_1107: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2396,
        in1(1) => S2386,
        out1 => S2491
    );
nor_n_613: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2490,
        in1(1) => S2397,
        out1 => S2492
    );
nand_n_1108: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2491,
        in1(1) => S2398,
        out1 => S2493
    );
nor_n_614: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2493,
        in1(1) => S2488,
        out1 => S2494
    );
nand_n_1109: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2492,
        in1(1) => S2489,
        out1 => S2495
    );
nor_n_615: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2480,
        in1(1) => S2474,
        out1 => S2496
    );
nand_n_1110: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2481,
        in1(1) => S2475,
        out1 => S2497
    );
nor_n_616: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2492,
        in1(1) => S2489,
        out1 => S2498
    );
nand_n_1111: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2493,
        in1(1) => S2488,
        out1 => S2499
    );
nor_n_617: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2498,
        in1(1) => S2494,
        out1 => S2500
    );
nand_n_1112: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2499,
        in1(1) => S2495,
        out1 => S2501
    );
nor_n_618: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2501,
        in1(1) => S2496,
        out1 => S2502
    );
nand_n_1113: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2500,
        in1(1) => S2497,
        out1 => S2503
    );
nor_n_619: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2502,
        in1(1) => S2494,
        out1 => S2504
    );
nand_n_1114: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2503,
        in1(1) => S2495,
        out1 => S2505
    );
nor_n_620: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2409,
        in1(1) => S2391,
        out1 => S2506
    );
nand_n_1115: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2410,
        in1(1) => S2392,
        out1 => S2507
    );
nor_n_621: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2506,
        in1(1) => S2411,
        out1 => S2508
    );
nand_n_1116: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2507,
        in1(1) => S2412,
        out1 => S2509
    );
nand_n_1117: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2508,
        in1(1) => S2505,
        out1 => S2510
    );
notg_196: ENTITY WORK.notg
    PORT MAP (
        in1 => S2510,
        out1 => S2511
    );
nand_n_1118: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2511,
        in1(1) => S2441,
        out1 => S2512
    );
notg_197: ENTITY WORK.notg
    PORT MAP (
        in1 => S2512,
        out1 => S2513
    );
nand_n_1119: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2510,
        in1(1) => S2440,
        out1 => S2514
    );
nand_n_1120: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2514,
        in1(1) => S2512,
        out1 => S2515
    );
notg_198: ENTITY WORK.notg
    PORT MAP (
        in1 => S2515,
        out1 => S2516
    );
nor_n_622: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2185,
        in1(1) => S1993,
        out1 => S2517
    );
nand_n_1121: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2184,
        in1(1) => U1_selMO_ARU,
        out1 => S2518
    );
nor_n_623: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2517,
        in1(1) => S1882,
        out1 => S2519
    );
nand_n_1122: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2518,
        in1(1) => U1_AC_out_7,
        out1 => S2520
    );
nand_n_1123: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2518,
        in1(1) => U1_AC_out_6,
        out1 => S2521
    );
nor_n_624: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2521,
        in1(1) => S2444,
        out1 => S2522
    );
nand_n_1124: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2519,
        in1(1) => S2445,
        out1 => S2523
    );
nor_n_625: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2361,
        in1(1) => S1872,
        out1 => S2524
    );
nand_n_1125: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2360,
        in1(1) => U1_AC_out_5,
        out1 => S2525
    );
nand_n_1126: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2520,
        in1(1) => S2446,
        out1 => S2526
    );
notg_199: ENTITY WORK.notg
    PORT MAP (
        in1 => S2526,
        out1 => S2527
    );
nor_n_626: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2527,
        in1(1) => S2522,
        out1 => S2528
    );
nand_n_1127: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2526,
        in1(1) => S2523,
        out1 => S2529
    );
nor_n_627: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2529,
        in1(1) => S2525,
        out1 => S2530
    );
nand_n_1128: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2528,
        in1(1) => S2524,
        out1 => S2531
    );
nor_n_628: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2530,
        in1(1) => S2522,
        out1 => S2532
    );
nand_n_1129: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2531,
        in1(1) => S2523,
        out1 => S2533
    );
nand_n_1130: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2452,
        in1(1) => S2449,
        out1 => S2534
    );
notg_200: ENTITY WORK.notg
    PORT MAP (
        in1 => S2534,
        out1 => S2535
    );
nor_n_629: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2535,
        in1(1) => S2454,
        out1 => S2536
    );
nand_n_1131: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2534,
        in1(1) => S2455,
        out1 => S2537
    );
nor_n_630: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2537,
        in1(1) => S2532,
        out1 => S2538
    );
nand_n_1132: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2536,
        in1(1) => S2533,
        out1 => S2539
    );
nor_n_631: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2536,
        in1(1) => S2533,
        out1 => S2540
    );
nand_n_1133: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2537,
        in1(1) => S2532,
        out1 => S2541
    );
nor_n_632: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2540,
        in1(1) => S2538,
        out1 => S2542
    );
nand_n_1134: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2541,
        in1(1) => S2539,
        out1 => S2543
    );
nor_n_633: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2284,
        in1(1) => S1932,
        out1 => S2544
    );
nand_n_1135: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2283,
        in1(1) => U1_AC_out_2,
        out1 => S2545
    );
nand_n_1136: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2232,
        in1(1) => U1_AC_out_4,
        out1 => S2546
    );
nor_n_634: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2275,
        in1(1) => S1852,
        out1 => S2547
    );
nand_n_1137: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2274,
        in1(1) => U1_AC_out_4,
        out1 => S2548
    );
nand_n_1138: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2274,
        in1(1) => U1_AC_out_3,
        out1 => S2549
    );
nor_n_635: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2548,
        in1(1) => S2473,
        out1 => S2550
    );
nand_n_1139: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2547,
        in1(1) => S2472,
        out1 => S2551
    );
nor_n_636: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2547,
        in1(1) => S2472,
        out1 => S2552
    );
nand_n_1140: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2548,
        in1(1) => S2473,
        out1 => S2553
    );
nor_n_637: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2552,
        in1(1) => S2550,
        out1 => S2554
    );
nand_n_1141: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2553,
        in1(1) => S2551,
        out1 => S2555
    );
nor_n_638: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2555,
        in1(1) => S2545,
        out1 => S2556
    );
nand_n_1142: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2554,
        in1(1) => S2544,
        out1 => S2557
    );
nor_n_639: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2554,
        in1(1) => S2544,
        out1 => S2558
    );
nand_n_1143: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2555,
        in1(1) => S2545,
        out1 => S2559
    );
nor_n_640: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2558,
        in1(1) => S2556,
        out1 => S2560
    );
nand_n_1144: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2559,
        in1(1) => S2557,
        out1 => S2561
    );
nor_n_641: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2561,
        in1(1) => S2543,
        out1 => S2562
    );
nand_n_1145: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2560,
        in1(1) => S2542,
        out1 => S2563
    );
nor_n_642: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2562,
        in1(1) => S2538,
        out1 => S2564
    );
nand_n_1146: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2563,
        in1(1) => S2539,
        out1 => S2565
    );
nor_n_643: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2484,
        in1(1) => S2466,
        out1 => S2566
    );
nand_n_1147: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2485,
        in1(1) => S2467,
        out1 => S2567
    );
nor_n_644: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2566,
        in1(1) => S2486,
        out1 => S2568
    );
nand_n_1148: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2567,
        in1(1) => S2487,
        out1 => S2569
    );
nor_n_645: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2569,
        in1(1) => S2564,
        out1 => S2570
    );
nand_n_1149: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2568,
        in1(1) => S2565,
        out1 => S2571
    );
nor_n_646: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2556,
        in1(1) => S2550,
        out1 => S2572
    );
nand_n_1150: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2557,
        in1(1) => S2551,
        out1 => S2573
    );
nor_n_647: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2568,
        in1(1) => S2565,
        out1 => S2574
    );
nand_n_1151: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2569,
        in1(1) => S2564,
        out1 => S2575
    );
nor_n_648: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2574,
        in1(1) => S2570,
        out1 => S2576
    );
nand_n_1152: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2575,
        in1(1) => S2571,
        out1 => S2577
    );
nor_n_649: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2577,
        in1(1) => S2572,
        out1 => S2578
    );
nand_n_1153: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2576,
        in1(1) => S2573,
        out1 => S2579
    );
nor_n_650: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2578,
        in1(1) => S2570,
        out1 => S2580
    );
nand_n_1154: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2579,
        in1(1) => S2571,
        out1 => S2581
    );
nor_n_651: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2500,
        in1(1) => S2497,
        out1 => S2582
    );
nand_n_1155: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2501,
        in1(1) => S2496,
        out1 => S2583
    );
nor_n_652: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2582,
        in1(1) => S2502,
        out1 => S2584
    );
nand_n_1156: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2583,
        in1(1) => S2503,
        out1 => S2585
    );
nand_n_1157: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2584,
        in1(1) => S2581,
        out1 => S2586
    );
notg_201: ENTITY WORK.notg
    PORT MAP (
        in1 => S2586,
        out1 => S2587
    );
nand_n_1158: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2509,
        in1(1) => S2504,
        out1 => S2588
    );
nand_n_1159: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2588,
        in1(1) => S2510,
        out1 => S2589
    );
notg_202: ENTITY WORK.notg
    PORT MAP (
        in1 => S2589,
        out1 => S2590
    );
nand_n_1160: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2590,
        in1(1) => S2587,
        out1 => S2591
    );
notg_203: ENTITY WORK.notg
    PORT MAP (
        in1 => S2591,
        out1 => S2592
    );
nand_n_1161: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2589,
        in1(1) => S2586,
        out1 => S2593
    );
nand_n_1162: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2593,
        in1(1) => S2591,
        out1 => S2594
    );
notg_204: ENTITY WORK.notg
    PORT MAP (
        in1 => S2594,
        out1 => S2595
    );
nor_n_653: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2528,
        in1(1) => S2524,
        out1 => S2596
    );
nand_n_1163: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2529,
        in1(1) => S2525,
        out1 => S2597
    );
nor_n_654: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2596,
        in1(1) => S2530,
        out1 => S2598
    );
nand_n_1164: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2597,
        in1(1) => S2531,
        out1 => S2599
    );
nand_n_1165: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2442,
        in1(1) => U1_AC_out_5,
        out1 => S2600
    );
nor_n_655: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2517,
        in1(1) => S1872,
        out1 => S2601
    );
nand_n_1166: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2518,
        in1(1) => U1_AC_out_5,
        out1 => S2602
    );
nor_n_656: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2602,
        in1(1) => S2446,
        out1 => S2603
    );
nand_n_1167: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2601,
        in1(1) => S2445,
        out1 => S2604
    );
nor_n_657: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2604,
        in1(1) => S2599,
        out1 => S2605
    );
nand_n_1168: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2603,
        in1(1) => S2598,
        out1 => S2606
    );
nor_n_658: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2603,
        in1(1) => S2598,
        out1 => S2607
    );
nand_n_1169: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2604,
        in1(1) => S2599,
        out1 => S2608
    );
nor_n_659: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2607,
        in1(1) => S2605,
        out1 => S2609
    );
nand_n_1170: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2608,
        in1(1) => S2606,
        out1 => S2610
    );
nor_n_660: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2272,
        in1(1) => S1932,
        out1 => S2611
    );
nand_n_1171: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2271,
        in1(1) => U1_AC_out_2,
        out1 => S2612
    );
nand_n_1172: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2148,
        in1(1) => U1_AC_out_3,
        out1 => S2613
    );
nor_n_661: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2322,
        in1(1) => S1939,
        out1 => S2614
    );
nand_n_1173: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2321,
        in1(1) => U1_AC_out_3,
        out1 => S2615
    );
nor_n_662: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2615,
        in1(1) => S2546,
        out1 => S2616
    );
notg_205: ENTITY WORK.notg
    PORT MAP (
        in1 => S2616,
        out1 => S2617
    );
nand_n_1174: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2321,
        in1(1) => U1_AC_out_4,
        out1 => S2618
    );
nand_n_1175: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2618,
        in1(1) => S2549,
        out1 => S2619
    );
notg_206: ENTITY WORK.notg
    PORT MAP (
        in1 => S2619,
        out1 => S2620
    );
nor_n_663: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2620,
        in1(1) => S2616,
        out1 => S2621
    );
nand_n_1176: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2619,
        in1(1) => S2617,
        out1 => S2622
    );
nor_n_664: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2622,
        in1(1) => S2612,
        out1 => S142
    );
notg_207: ENTITY WORK.notg
    PORT MAP (
        in1 => S142,
        out1 => S143
    );
nor_n_665: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2621,
        in1(1) => S2611,
        out1 => S144
    );
nand_n_1177: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2622,
        in1(1) => S2612,
        out1 => S145
    );
nor_n_666: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S144,
        in1(1) => S142,
        out1 => S146
    );
nand_n_1178: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S145,
        in1(1) => S143,
        out1 => S147
    );
nor_n_667: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S147,
        in1(1) => S2610,
        out1 => S148
    );
nand_n_1179: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S146,
        in1(1) => S2609,
        out1 => S149
    );
nor_n_668: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S148,
        in1(1) => S2605,
        out1 => S150
    );
nand_n_1180: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S149,
        in1(1) => S2606,
        out1 => S151
    );
nor_n_669: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2560,
        in1(1) => S2542,
        out1 => S152
    );
nand_n_1181: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2561,
        in1(1) => S2543,
        out1 => S153
    );
nor_n_670: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S152,
        in1(1) => S2562,
        out1 => S154
    );
nand_n_1182: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S153,
        in1(1) => S2563,
        out1 => S155
    );
nor_n_671: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S155,
        in1(1) => S150,
        out1 => S156
    );
nand_n_1183: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S154,
        in1(1) => S151,
        out1 => S157
    );
nor_n_672: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S154,
        in1(1) => S151,
        out1 => S158
    );
nand_n_1184: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S155,
        in1(1) => S150,
        out1 => S159
    );
nor_n_673: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S158,
        in1(1) => S156,
        out1 => S160
    );
nand_n_1185: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S159,
        in1(1) => S157,
        out1 => S161
    );
nand_n_1186: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2305,
        in1(1) => U1_AC_out_1,
        out1 => S162
    );
notg_208: ENTITY WORK.notg
    PORT MAP (
        in1 => S162,
        out1 => S163
    );
nor_n_674: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S142,
        in1(1) => S2616,
        out1 => S164
    );
notg_209: ENTITY WORK.notg
    PORT MAP (
        in1 => S164,
        out1 => S165
    );
nor_n_675: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S164,
        in1(1) => S162,
        out1 => S166
    );
nand_n_1187: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S165,
        in1(1) => S163,
        out1 => S167
    );
nand_n_1188: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S164,
        in1(1) => S162,
        out1 => S168
    );
notg_210: ENTITY WORK.notg
    PORT MAP (
        in1 => S168,
        out1 => S169
    );
nor_n_676: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S169,
        in1(1) => S166,
        out1 => S170
    );
nand_n_1189: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S168,
        in1(1) => S167,
        out1 => S171
    );
nor_n_677: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S171,
        in1(1) => S161,
        out1 => S172
    );
nand_n_1190: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S170,
        in1(1) => S160,
        out1 => S173
    );
nor_n_678: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S172,
        in1(1) => S156,
        out1 => S174
    );
nand_n_1191: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2577,
        in1(1) => S2572,
        out1 => S175
    );
nand_n_1192: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S175,
        in1(1) => S2579,
        out1 => S176
    );
nor_n_679: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S176,
        in1(1) => S174,
        out1 => S177
    );
notg_211: ENTITY WORK.notg
    PORT MAP (
        in1 => S177,
        out1 => S178
    );
nand_n_1193: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S176,
        in1(1) => S174,
        out1 => S179
    );
nand_n_1194: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S179,
        in1(1) => S178,
        out1 => S180
    );
notg_212: ENTITY WORK.notg
    PORT MAP (
        in1 => S180,
        out1 => S181
    );
nor_n_680: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S180,
        in1(1) => S167,
        out1 => S182
    );
nand_n_1195: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S181,
        in1(1) => S166,
        out1 => S183
    );
nor_n_681: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S182,
        in1(1) => S177,
        out1 => S184
    );
notg_213: ENTITY WORK.notg
    PORT MAP (
        in1 => S184,
        out1 => S185
    );
nand_n_1196: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2585,
        in1(1) => S2580,
        out1 => S186
    );
nand_n_1197: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S186,
        in1(1) => S2586,
        out1 => S187
    );
notg_214: ENTITY WORK.notg
    PORT MAP (
        in1 => S187,
        out1 => S188
    );
nand_n_1198: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S188,
        in1(1) => S185,
        out1 => S189
    );
notg_215: ENTITY WORK.notg
    PORT MAP (
        in1 => S189,
        out1 => S190
    );
nand_n_1199: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S187,
        in1(1) => S184,
        out1 => S191
    );
nand_n_1200: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S191,
        in1(1) => S189,
        out1 => S192
    );
notg_216: ENTITY WORK.notg
    PORT MAP (
        in1 => S192,
        out1 => S193
    );
nor_n_682: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S146,
        in1(1) => S2609,
        out1 => S194
    );
nand_n_1201: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S147,
        in1(1) => S2610,
        out1 => S195
    );
nor_n_683: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S194,
        in1(1) => S148,
        out1 => S196
    );
nand_n_1202: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S195,
        in1(1) => S149,
        out1 => S197
    );
nand_n_1203: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2600,
        in1(1) => S2521,
        out1 => S198
    );
notg_217: ENTITY WORK.notg
    PORT MAP (
        in1 => S198,
        out1 => S199
    );
nor_n_684: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S199,
        in1(1) => S2603,
        out1 => S200
    );
nand_n_1204: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S198,
        in1(1) => S2604,
        out1 => S201
    );
nor_n_685: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2275,
        in1(1) => S1932,
        out1 => S202
    );
nand_n_1205: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2274,
        in1(1) => U1_AC_out_2,
        out1 => S203
    );
nand_n_1206: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2360,
        in1(1) => U1_AC_out_3,
        out1 => S204
    );
nor_n_686: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2361,
        in1(1) => S1852,
        out1 => S205
    );
nand_n_1207: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2360,
        in1(1) => U1_AC_out_4,
        out1 => S206
    );
nor_n_687: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S206,
        in1(1) => S2615,
        out1 => S207
    );
nand_n_1208: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S205,
        in1(1) => S2614,
        out1 => S208
    );
nor_n_688: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S205,
        in1(1) => S2614,
        out1 => S209
    );
nand_n_1209: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S206,
        in1(1) => S2615,
        out1 => S210
    );
nor_n_689: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S209,
        in1(1) => S207,
        out1 => S211
    );
nand_n_1210: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S210,
        in1(1) => S208,
        out1 => S212
    );
nor_n_690: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S212,
        in1(1) => S203,
        out1 => S213
    );
nand_n_1211: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S211,
        in1(1) => S202,
        out1 => S214
    );
nor_n_691: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S211,
        in1(1) => S202,
        out1 => S215
    );
nand_n_1212: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S212,
        in1(1) => S203,
        out1 => S216
    );
nor_n_692: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S215,
        in1(1) => S213,
        out1 => S217
    );
nand_n_1213: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S216,
        in1(1) => S214,
        out1 => S218
    );
nor_n_693: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S218,
        in1(1) => S201,
        out1 => S219
    );
nand_n_1214: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S217,
        in1(1) => S200,
        out1 => S220
    );
nor_n_694: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S220,
        in1(1) => S197,
        out1 => S221
    );
nand_n_1215: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S219,
        in1(1) => S196,
        out1 => S222
    );
nor_n_695: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S219,
        in1(1) => S196,
        out1 => S223
    );
nand_n_1216: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S220,
        in1(1) => S197,
        out1 => S224
    );
nor_n_696: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S223,
        in1(1) => S221,
        out1 => S225
    );
nand_n_1217: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S224,
        in1(1) => S222,
        out1 => S226
    );
nor_n_697: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2306,
        in1(1) => S1917,
        out1 => S227
    );
nand_n_1218: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2305,
        in1(1) => U1_AC_out_0,
        out1 => S228
    );
nor_n_698: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2284,
        in1(1) => S1925,
        out1 => S229
    );
nand_n_1219: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2283,
        in1(1) => U1_AC_out_1,
        out1 => S230
    );
nor_n_699: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S213,
        in1(1) => S207,
        out1 => S231
    );
nand_n_1220: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S214,
        in1(1) => S208,
        out1 => S232
    );
nor_n_700: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S231,
        in1(1) => S230,
        out1 => S233
    );
nand_n_1221: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S232,
        in1(1) => S229,
        out1 => S234
    );
nor_n_701: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S232,
        in1(1) => S229,
        out1 => S235
    );
nand_n_1222: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S231,
        in1(1) => S230,
        out1 => S236
    );
nor_n_702: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S235,
        in1(1) => S233,
        out1 => S237
    );
nand_n_1223: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S236,
        in1(1) => S234,
        out1 => S238
    );
nor_n_703: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S238,
        in1(1) => S228,
        out1 => S239
    );
nand_n_1224: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S237,
        in1(1) => S227,
        out1 => S240
    );
nor_n_704: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S237,
        in1(1) => S227,
        out1 => S241
    );
nand_n_1225: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S238,
        in1(1) => S228,
        out1 => S242
    );
nor_n_705: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S241,
        in1(1) => S239,
        out1 => S243
    );
nand_n_1226: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S242,
        in1(1) => S240,
        out1 => S244
    );
nor_n_706: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S244,
        in1(1) => S226,
        out1 => S245
    );
nand_n_1227: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S243,
        in1(1) => S225,
        out1 => S246
    );
nor_n_707: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S245,
        in1(1) => S221,
        out1 => S247
    );
nand_n_1228: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S246,
        in1(1) => S222,
        out1 => S248
    );
nor_n_708: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S170,
        in1(1) => S160,
        out1 => S249
    );
nand_n_1229: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S171,
        in1(1) => S161,
        out1 => S250
    );
nor_n_709: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S249,
        in1(1) => S172,
        out1 => S251
    );
nand_n_1230: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S250,
        in1(1) => S173,
        out1 => S252
    );
nor_n_710: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S252,
        in1(1) => S247,
        out1 => S253
    );
notg_218: ENTITY WORK.notg
    PORT MAP (
        in1 => S253,
        out1 => S254
    );
nor_n_711: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S239,
        in1(1) => S233,
        out1 => S255
    );
nand_n_1231: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S240,
        in1(1) => S234,
        out1 => S256
    );
nor_n_712: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S251,
        in1(1) => S248,
        out1 => S257
    );
nand_n_1232: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S252,
        in1(1) => S247,
        out1 => S258
    );
nor_n_713: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S257,
        in1(1) => S253,
        out1 => S259
    );
nand_n_1233: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S258,
        in1(1) => S254,
        out1 => S260
    );
nor_n_714: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S260,
        in1(1) => S255,
        out1 => S261
    );
nor_n_715: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S261,
        in1(1) => S253,
        out1 => S262
    );
notg_219: ENTITY WORK.notg
    PORT MAP (
        in1 => S262,
        out1 => S263
    );
nand_n_1234: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S180,
        in1(1) => S167,
        out1 => S264
    );
nand_n_1235: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S264,
        in1(1) => S183,
        out1 => S265
    );
notg_220: ENTITY WORK.notg
    PORT MAP (
        in1 => S265,
        out1 => S266
    );
nand_n_1236: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S266,
        in1(1) => S263,
        out1 => S267
    );
notg_221: ENTITY WORK.notg
    PORT MAP (
        in1 => S267,
        out1 => S268
    );
nand_n_1237: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S265,
        in1(1) => S262,
        out1 => S269
    );
nand_n_1238: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S269,
        in1(1) => S267,
        out1 => S270
    );
notg_222: ENTITY WORK.notg
    PORT MAP (
        in1 => S270,
        out1 => S271
    );
nor_n_716: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S217,
        in1(1) => S200,
        out1 => S272
    );
nand_n_1239: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S218,
        in1(1) => S201,
        out1 => S273
    );
nor_n_717: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S272,
        in1(1) => S219,
        out1 => S274
    );
nand_n_1240: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S273,
        in1(1) => S220,
        out1 => S275
    );
nand_n_1241: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2321,
        in1(1) => U1_AC_out_2,
        out1 => S276
    );
nand_n_1242: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2442,
        in1(1) => U1_AC_out_4,
        out1 => S277
    );
nor_n_718: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2443,
        in1(1) => S1939,
        out1 => S278
    );
nand_n_1243: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2442,
        in1(1) => U1_AC_out_3,
        out1 => S279
    );
nor_n_719: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S279,
        in1(1) => S206,
        out1 => S280
    );
notg_223: ENTITY WORK.notg
    PORT MAP (
        in1 => S280,
        out1 => S281
    );
nand_n_1244: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S277,
        in1(1) => S204,
        out1 => S282
    );
nand_n_1245: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S282,
        in1(1) => S281,
        out1 => S283
    );
nand_n_1246: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S283,
        in1(1) => S276,
        out1 => S284
    );
notg_224: ENTITY WORK.notg
    PORT MAP (
        in1 => S284,
        out1 => S285
    );
nor_n_720: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S283,
        in1(1) => S276,
        out1 => S286
    );
notg_225: ENTITY WORK.notg
    PORT MAP (
        in1 => S286,
        out1 => S287
    );
nor_n_721: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S286,
        in1(1) => S285,
        out1 => S288
    );
nand_n_1247: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S287,
        in1(1) => S284,
        out1 => S289
    );
nor_n_722: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S289,
        in1(1) => S2602,
        out1 => S290
    );
nand_n_1248: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S288,
        in1(1) => S2601,
        out1 => S291
    );
nor_n_723: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S291,
        in1(1) => S275,
        out1 => S292
    );
nand_n_1249: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S290,
        in1(1) => S274,
        out1 => S293
    );
nor_n_724: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S290,
        in1(1) => S274,
        out1 => S294
    );
nand_n_1250: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S291,
        in1(1) => S275,
        out1 => S295
    );
nor_n_725: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S294,
        in1(1) => S292,
        out1 => S296
    );
nand_n_1251: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S295,
        in1(1) => S293,
        out1 => S297
    );
nor_n_726: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2284,
        in1(1) => S1917,
        out1 => S298
    );
nand_n_1252: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2283,
        in1(1) => U1_AC_out_0,
        out1 => S299
    );
nand_n_1253: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2271,
        in1(1) => U1_AC_out_1,
        out1 => S300
    );
notg_226: ENTITY WORK.notg
    PORT MAP (
        in1 => S300,
        out1 => S301
    );
nor_n_727: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S286,
        in1(1) => S280,
        out1 => S302
    );
notg_227: ENTITY WORK.notg
    PORT MAP (
        in1 => S302,
        out1 => S303
    );
nor_n_728: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S302,
        in1(1) => S300,
        out1 => S304
    );
nand_n_1254: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S303,
        in1(1) => S301,
        out1 => S305
    );
nand_n_1255: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S302,
        in1(1) => S300,
        out1 => S306
    );
notg_228: ENTITY WORK.notg
    PORT MAP (
        in1 => S306,
        out1 => S307
    );
nor_n_729: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S307,
        in1(1) => S304,
        out1 => S308
    );
nand_n_1256: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S306,
        in1(1) => S305,
        out1 => S309
    );
nor_n_730: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S309,
        in1(1) => S299,
        out1 => S310
    );
nand_n_1257: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S308,
        in1(1) => S298,
        out1 => S311
    );
nor_n_731: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S308,
        in1(1) => S298,
        out1 => S312
    );
nand_n_1258: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S309,
        in1(1) => S299,
        out1 => S313
    );
nor_n_732: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S312,
        in1(1) => S310,
        out1 => S314
    );
nand_n_1259: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S313,
        in1(1) => S311,
        out1 => S315
    );
nor_n_733: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S315,
        in1(1) => S297,
        out1 => S316
    );
nand_n_1260: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S314,
        in1(1) => S296,
        out1 => S317
    );
nor_n_734: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S316,
        in1(1) => S292,
        out1 => S318
    );
nand_n_1261: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S317,
        in1(1) => S293,
        out1 => S319
    );
nor_n_735: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S243,
        in1(1) => S225,
        out1 => S320
    );
nand_n_1262: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S244,
        in1(1) => S226,
        out1 => S321
    );
nor_n_736: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S320,
        in1(1) => S245,
        out1 => S322
    );
nand_n_1263: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S321,
        in1(1) => S246,
        out1 => S323
    );
nor_n_737: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S323,
        in1(1) => S318,
        out1 => S324
    );
nand_n_1264: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S322,
        in1(1) => S319,
        out1 => S325
    );
nand_n_1265: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S311,
        in1(1) => S305,
        out1 => S326
    );
notg_229: ENTITY WORK.notg
    PORT MAP (
        in1 => S326,
        out1 => S327
    );
nor_n_738: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S322,
        in1(1) => S319,
        out1 => S328
    );
nand_n_1266: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S323,
        in1(1) => S318,
        out1 => S329
    );
nor_n_739: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S328,
        in1(1) => S324,
        out1 => S330
    );
nand_n_1267: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S329,
        in1(1) => S325,
        out1 => S331
    );
nor_n_740: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S331,
        in1(1) => S327,
        out1 => S332
    );
nand_n_1268: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S330,
        in1(1) => S326,
        out1 => S333
    );
nand_n_1269: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S333,
        in1(1) => S325,
        out1 => S334
    );
notg_230: ENTITY WORK.notg
    PORT MAP (
        in1 => S334,
        out1 => S335
    );
nor_n_741: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S259,
        in1(1) => S256,
        out1 => S336
    );
nor_n_742: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S336,
        in1(1) => S261,
        out1 => S337
    );
notg_231: ENTITY WORK.notg
    PORT MAP (
        in1 => S337,
        out1 => S338
    );
nor_n_743: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S338,
        in1(1) => S335,
        out1 => S339
    );
notg_232: ENTITY WORK.notg
    PORT MAP (
        in1 => S339,
        out1 => S340
    );
nor_n_744: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S337,
        in1(1) => S334,
        out1 => S341
    );
nor_n_745: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S341,
        in1(1) => S339,
        out1 => S342
    );
notg_233: ENTITY WORK.notg
    PORT MAP (
        in1 => S342,
        out1 => S343
    );
nor_n_746: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S314,
        in1(1) => S296,
        out1 => S344
    );
nand_n_1270: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S315,
        in1(1) => S297,
        out1 => S345
    );
nor_n_747: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S344,
        in1(1) => S316,
        out1 => S346
    );
nand_n_1271: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S345,
        in1(1) => S317,
        out1 => S347
    );
nor_n_748: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S288,
        in1(1) => S2601,
        out1 => S348
    );
nand_n_1272: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S289,
        in1(1) => S2602,
        out1 => S349
    );
nor_n_749: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S348,
        in1(1) => S290,
        out1 => S350
    );
nand_n_1273: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S349,
        in1(1) => S291,
        out1 => S351
    );
nor_n_750: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2272,
        in1(1) => S1917,
        out1 => S352
    );
nand_n_1274: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2271,
        in1(1) => U1_AC_out_0,
        out1 => S353
    );
nor_n_751: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2275,
        in1(1) => S1925,
        out1 => S354
    );
nand_n_1275: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2274,
        in1(1) => U1_AC_out_1,
        out1 => S355
    );
nor_n_752: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2517,
        in1(1) => S1852,
        out1 => S356
    );
nand_n_1276: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2518,
        in1(1) => U1_AC_out_4,
        out1 => S357
    );
nand_n_1277: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2518,
        in1(1) => U1_AC_out_3,
        out1 => S358
    );
nor_n_753: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S358,
        in1(1) => S277,
        out1 => S359
    );
nand_n_1278: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S356,
        in1(1) => S278,
        out1 => S360
    );
nand_n_1279: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2159,
        in1(1) => U1_AC_out_2,
        out1 => S361
    );
nor_n_754: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2361,
        in1(1) => S1932,
        out1 => S362
    );
nand_n_1280: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2360,
        in1(1) => U1_AC_out_2,
        out1 => S363
    );
nand_n_1281: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S357,
        in1(1) => S279,
        out1 => S364
    );
notg_234: ENTITY WORK.notg
    PORT MAP (
        in1 => S364,
        out1 => S365
    );
nor_n_755: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S365,
        in1(1) => S359,
        out1 => S366
    );
nand_n_1282: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S364,
        in1(1) => S360,
        out1 => S367
    );
nor_n_756: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S367,
        in1(1) => S363,
        out1 => S368
    );
nand_n_1283: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S366,
        in1(1) => S362,
        out1 => S369
    );
nor_n_757: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S368,
        in1(1) => S359,
        out1 => S370
    );
nand_n_1284: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S369,
        in1(1) => S360,
        out1 => S371
    );
nor_n_758: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S370,
        in1(1) => S355,
        out1 => S372
    );
nand_n_1285: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S371,
        in1(1) => S354,
        out1 => S373
    );
nor_n_759: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S371,
        in1(1) => S354,
        out1 => S374
    );
nand_n_1286: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S370,
        in1(1) => S355,
        out1 => S375
    );
nor_n_760: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S374,
        in1(1) => S372,
        out1 => S376
    );
nand_n_1287: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S375,
        in1(1) => S373,
        out1 => S377
    );
nor_n_761: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S377,
        in1(1) => S353,
        out1 => S378
    );
nand_n_1288: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S376,
        in1(1) => S352,
        out1 => S379
    );
nor_n_762: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S376,
        in1(1) => S352,
        out1 => S380
    );
nand_n_1289: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S377,
        in1(1) => S353,
        out1 => S381
    );
nor_n_763: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S380,
        in1(1) => S378,
        out1 => S382
    );
nand_n_1290: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S381,
        in1(1) => S379,
        out1 => S383
    );
nor_n_764: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S383,
        in1(1) => S351,
        out1 => S384
    );
nand_n_1291: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S382,
        in1(1) => S350,
        out1 => S385
    );
nor_n_765: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S385,
        in1(1) => S347,
        out1 => S386
    );
nand_n_1292: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S384,
        in1(1) => S346,
        out1 => S387
    );
nor_n_766: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S378,
        in1(1) => S372,
        out1 => S388
    );
nand_n_1293: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S379,
        in1(1) => S373,
        out1 => S389
    );
nor_n_767: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S384,
        in1(1) => S346,
        out1 => S390
    );
nand_n_1294: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S385,
        in1(1) => S347,
        out1 => S391
    );
nor_n_768: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S390,
        in1(1) => S386,
        out1 => S392
    );
nand_n_1295: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S391,
        in1(1) => S387,
        out1 => S393
    );
nor_n_769: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S393,
        in1(1) => S388,
        out1 => S394
    );
nand_n_1296: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S392,
        in1(1) => S389,
        out1 => S395
    );
nand_n_1297: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S395,
        in1(1) => S387,
        out1 => S396
    );
notg_235: ENTITY WORK.notg
    PORT MAP (
        in1 => S396,
        out1 => S397
    );
nor_n_770: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S330,
        in1(1) => S326,
        out1 => S398
    );
nor_n_771: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S398,
        in1(1) => S332,
        out1 => S399
    );
notg_236: ENTITY WORK.notg
    PORT MAP (
        in1 => S399,
        out1 => S400
    );
nor_n_772: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S400,
        in1(1) => S397,
        out1 => S401
    );
notg_237: ENTITY WORK.notg
    PORT MAP (
        in1 => S401,
        out1 => S402
    );
nor_n_773: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S399,
        in1(1) => S396,
        out1 => S403
    );
nor_n_774: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S403,
        in1(1) => S401,
        out1 => S404
    );
notg_238: ENTITY WORK.notg
    PORT MAP (
        in1 => S404,
        out1 => S405
    );
nor_n_775: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S382,
        in1(1) => S350,
        out1 => S406
    );
nand_n_1298: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S383,
        in1(1) => S351,
        out1 => S407
    );
nor_n_776: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S406,
        in1(1) => S384,
        out1 => S408
    );
nand_n_1299: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S407,
        in1(1) => S385,
        out1 => S409
    );
nor_n_777: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S366,
        in1(1) => S362,
        out1 => S410
    );
nand_n_1300: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S367,
        in1(1) => S363,
        out1 => S411
    );
nor_n_778: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S410,
        in1(1) => S368,
        out1 => S412
    );
nand_n_1301: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S411,
        in1(1) => S369,
        out1 => S413
    );
nor_n_779: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2275,
        in1(1) => S1917,
        out1 => S414
    );
nand_n_1302: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2274,
        in1(1) => U1_AC_out_0,
        out1 => S415
    );
nor_n_780: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2322,
        in1(1) => S1925,
        out1 => S416
    );
nand_n_1303: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2321,
        in1(1) => U1_AC_out_1,
        out1 => S417
    );
nand_n_1304: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2442,
        in1(1) => U1_AC_out_2,
        out1 => S418
    );
nand_n_1305: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2518,
        in1(1) => U1_AC_out_2,
        out1 => S419
    );
notg_239: ENTITY WORK.notg
    PORT MAP (
        in1 => S419,
        out1 => S420
    );
nor_n_781: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S419,
        in1(1) => S279,
        out1 => S421
    );
nand_n_1306: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S420,
        in1(1) => S278,
        out1 => S422
    );
nor_n_782: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S422,
        in1(1) => S417,
        out1 => S423
    );
nand_n_1307: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S421,
        in1(1) => S416,
        out1 => S424
    );
nor_n_783: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S421,
        in1(1) => S416,
        out1 => S425
    );
nand_n_1308: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S422,
        in1(1) => S417,
        out1 => S426
    );
nor_n_784: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S425,
        in1(1) => S423,
        out1 => S427
    );
nand_n_1309: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S426,
        in1(1) => S424,
        out1 => S428
    );
nor_n_785: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S428,
        in1(1) => S415,
        out1 => S429
    );
nand_n_1310: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S427,
        in1(1) => S414,
        out1 => S430
    );
nor_n_786: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S427,
        in1(1) => S414,
        out1 => S431
    );
nand_n_1311: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S428,
        in1(1) => S415,
        out1 => S432
    );
nor_n_787: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S431,
        in1(1) => S429,
        out1 => S433
    );
nand_n_1312: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S432,
        in1(1) => S430,
        out1 => S434
    );
nor_n_788: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S434,
        in1(1) => S413,
        out1 => S435
    );
nand_n_1313: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S433,
        in1(1) => S412,
        out1 => S436
    );
nor_n_789: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S436,
        in1(1) => S409,
        out1 => S437
    );
nand_n_1314: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S435,
        in1(1) => S408,
        out1 => S438
    );
nor_n_790: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S429,
        in1(1) => S423,
        out1 => S439
    );
nand_n_1315: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S430,
        in1(1) => S424,
        out1 => S440
    );
nor_n_791: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S435,
        in1(1) => S408,
        out1 => S441
    );
nand_n_1316: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S436,
        in1(1) => S409,
        out1 => S442
    );
nor_n_792: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S441,
        in1(1) => S437,
        out1 => S443
    );
nand_n_1317: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S442,
        in1(1) => S438,
        out1 => S444
    );
nor_n_793: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S444,
        in1(1) => S439,
        out1 => S445
    );
nand_n_1318: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S443,
        in1(1) => S440,
        out1 => S446
    );
nor_n_794: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S445,
        in1(1) => S437,
        out1 => S447
    );
notg_240: ENTITY WORK.notg
    PORT MAP (
        in1 => S447,
        out1 => S448
    );
nor_n_795: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S392,
        in1(1) => S389,
        out1 => S449
    );
nand_n_1319: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S393,
        in1(1) => S388,
        out1 => S450
    );
nor_n_796: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S449,
        in1(1) => S394,
        out1 => S451
    );
nand_n_1320: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S450,
        in1(1) => S395,
        out1 => S452
    );
nand_n_1321: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S451,
        in1(1) => S448,
        out1 => S453
    );
notg_241: ENTITY WORK.notg
    PORT MAP (
        in1 => S453,
        out1 => S454
    );
nand_n_1322: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S452,
        in1(1) => S447,
        out1 => S455
    );
nand_n_1323: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S455,
        in1(1) => S453,
        out1 => S456
    );
notg_242: ENTITY WORK.notg
    PORT MAP (
        in1 => S456,
        out1 => S457
    );
nor_n_797: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S433,
        in1(1) => S412,
        out1 => S458
    );
nand_n_1324: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S434,
        in1(1) => S413,
        out1 => S459
    );
nor_n_798: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S458,
        in1(1) => S435,
        out1 => S460
    );
nand_n_1325: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S459,
        in1(1) => S436,
        out1 => S461
    );
nand_n_1326: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S418,
        in1(1) => S358,
        out1 => S462
    );
notg_243: ENTITY WORK.notg
    PORT MAP (
        in1 => S462,
        out1 => S463
    );
nor_n_799: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S463,
        in1(1) => S421,
        out1 => S464
    );
nand_n_1327: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S462,
        in1(1) => S422,
        out1 => S465
    );
nand_n_1328: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2321,
        in1(1) => U1_AC_out_0,
        out1 => S466
    );
nand_n_1329: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2360,
        in1(1) => U1_AC_out_1,
        out1 => S467
    );
nor_n_800: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2361,
        in1(1) => S1917,
        out1 => S468
    );
nand_n_1330: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2360,
        in1(1) => U1_AC_out_0,
        out1 => S469
    );
nor_n_801: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S469,
        in1(1) => S417,
        out1 => S470
    );
nand_n_1331: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S468,
        in1(1) => S416,
        out1 => S471
    );
nand_n_1332: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S467,
        in1(1) => S466,
        out1 => S472
    );
notg_244: ENTITY WORK.notg
    PORT MAP (
        in1 => S472,
        out1 => S473
    );
nor_n_802: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S473,
        in1(1) => S470,
        out1 => S474
    );
nand_n_1333: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S472,
        in1(1) => S471,
        out1 => S475
    );
nor_n_803: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S475,
        in1(1) => S465,
        out1 => S476
    );
nand_n_1334: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S474,
        in1(1) => S464,
        out1 => S477
    );
nor_n_804: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S477,
        in1(1) => S461,
        out1 => S478
    );
nand_n_1335: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S476,
        in1(1) => S460,
        out1 => S479
    );
nor_n_805: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S476,
        in1(1) => S460,
        out1 => S480
    );
nand_n_1336: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S477,
        in1(1) => S461,
        out1 => S481
    );
nor_n_806: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S480,
        in1(1) => S478,
        out1 => S482
    );
nand_n_1337: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S481,
        in1(1) => S479,
        out1 => S483
    );
nor_n_807: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S483,
        in1(1) => S471,
        out1 => S484
    );
nand_n_1338: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S482,
        in1(1) => S470,
        out1 => S485
    );
nor_n_808: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S484,
        in1(1) => S478,
        out1 => S486
    );
nand_n_1339: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S485,
        in1(1) => S479,
        out1 => S487
    );
nor_n_809: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S443,
        in1(1) => S440,
        out1 => S488
    );
nand_n_1340: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S444,
        in1(1) => S439,
        out1 => S489
    );
nor_n_810: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S488,
        in1(1) => S445,
        out1 => S490
    );
nand_n_1341: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S489,
        in1(1) => S446,
        out1 => S491
    );
nor_n_811: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S491,
        in1(1) => S486,
        out1 => S492
    );
nand_n_1342: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S490,
        in1(1) => S487,
        out1 => S493
    );
nor_n_812: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S474,
        in1(1) => S464,
        out1 => S494
    );
nand_n_1343: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S475,
        in1(1) => S465,
        out1 => S495
    );
nor_n_813: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S494,
        in1(1) => S476,
        out1 => S496
    );
nand_n_1344: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S495,
        in1(1) => S477,
        out1 => S497
    );
nor_n_814: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2443,
        in1(1) => S1925,
        out1 => S498
    );
nand_n_1345: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2442,
        in1(1) => U1_AC_out_1,
        out1 => S499
    );
nor_n_815: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2443,
        in1(1) => S1917,
        out1 => S500
    );
nor_n_816: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S499,
        in1(1) => S469,
        out1 => S501
    );
nand_n_1346: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S498,
        in1(1) => S468,
        out1 => S502
    );
nand_n_1347: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S499,
        in1(1) => S469,
        out1 => S503
    );
nand_n_1348: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S503,
        in1(1) => S502,
        out1 => S504
    );
notg_245: ENTITY WORK.notg
    PORT MAP (
        in1 => S504,
        out1 => S505
    );
nor_n_817: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S504,
        in1(1) => S419,
        out1 => S506
    );
nand_n_1349: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S505,
        in1(1) => S420,
        out1 => S507
    );
nor_n_818: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S507,
        in1(1) => S497,
        out1 => S508
    );
nand_n_1350: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S506,
        in1(1) => S496,
        out1 => S509
    );
nor_n_819: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S506,
        in1(1) => S496,
        out1 => S510
    );
nor_n_820: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S510,
        in1(1) => S508,
        out1 => S511
    );
notg_246: ENTITY WORK.notg
    PORT MAP (
        in1 => S511,
        out1 => S512
    );
nor_n_821: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S512,
        in1(1) => S502,
        out1 => S513
    );
notg_247: ENTITY WORK.notg
    PORT MAP (
        in1 => S513,
        out1 => S514
    );
nand_n_1351: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S514,
        in1(1) => S509,
        out1 => S515
    );
notg_248: ENTITY WORK.notg
    PORT MAP (
        in1 => S515,
        out1 => S516
    );
nor_n_822: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S482,
        in1(1) => S470,
        out1 => S517
    );
nand_n_1352: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S483,
        in1(1) => S471,
        out1 => S518
    );
nor_n_823: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S517,
        in1(1) => S484,
        out1 => S519
    );
nand_n_1353: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S518,
        in1(1) => S485,
        out1 => S520
    );
nor_n_824: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S520,
        in1(1) => S516,
        out1 => S521
    );
notg_249: ENTITY WORK.notg
    PORT MAP (
        in1 => S521,
        out1 => S522
    );
nand_n_1354: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2185,
        in1(1) => U1_AC_out_0,
        out1 => S523
    );
notg_250: ENTITY WORK.notg
    PORT MAP (
        in1 => S523,
        out1 => S524
    );
nand_n_1355: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S524,
        in1(1) => S498,
        out1 => S525
    );
nand_n_1356: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S504,
        in1(1) => S419,
        out1 => S526
    );
nand_n_1357: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S526,
        in1(1) => S507,
        out1 => S527
    );
nor_n_825: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S527,
        in1(1) => S525,
        out1 => S528
    );
notg_251: ENTITY WORK.notg
    PORT MAP (
        in1 => S528,
        out1 => S529
    );
nor_n_826: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S511,
        in1(1) => S501,
        out1 => S530
    );
nor_n_827: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S530,
        in1(1) => S513,
        out1 => S531
    );
notg_252: ENTITY WORK.notg
    PORT MAP (
        in1 => S531,
        out1 => S532
    );
nor_n_828: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S532,
        in1(1) => S529,
        out1 => S533
    );
nor_n_829: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S519,
        in1(1) => S515,
        out1 => S534
    );
nor_n_830: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S534,
        in1(1) => S521,
        out1 => S535
    );
nand_n_1358: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S535,
        in1(1) => S533,
        out1 => S536
    );
notg_253: ENTITY WORK.notg
    PORT MAP (
        in1 => S536,
        out1 => S537
    );
nor_n_831: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S537,
        in1(1) => S521,
        out1 => S538
    );
nand_n_1359: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S536,
        in1(1) => S522,
        out1 => S539
    );
nor_n_832: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S490,
        in1(1) => S487,
        out1 => S540
    );
nand_n_1360: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S491,
        in1(1) => S486,
        out1 => S541
    );
nor_n_833: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S540,
        in1(1) => S492,
        out1 => S542
    );
nand_n_1361: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S541,
        in1(1) => S493,
        out1 => S543
    );
nor_n_834: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S543,
        in1(1) => S538,
        out1 => S544
    );
nand_n_1362: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S542,
        in1(1) => S539,
        out1 => S545
    );
nor_n_835: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S544,
        in1(1) => S492,
        out1 => S546
    );
nand_n_1363: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S545,
        in1(1) => S493,
        out1 => S547
    );
nor_n_836: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S546,
        in1(1) => S456,
        out1 => S548
    );
nand_n_1364: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S547,
        in1(1) => S457,
        out1 => S549
    );
nor_n_837: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S548,
        in1(1) => S454,
        out1 => S550
    );
nand_n_1365: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S549,
        in1(1) => S453,
        out1 => S551
    );
nor_n_838: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S550,
        in1(1) => S405,
        out1 => S552
    );
nand_n_1366: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S551,
        in1(1) => S404,
        out1 => S553
    );
nor_n_839: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S552,
        in1(1) => S401,
        out1 => S554
    );
nand_n_1367: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S553,
        in1(1) => S402,
        out1 => S555
    );
nor_n_840: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S554,
        in1(1) => S343,
        out1 => S556
    );
nand_n_1368: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S555,
        in1(1) => S342,
        out1 => S557
    );
nor_n_841: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S556,
        in1(1) => S339,
        out1 => S558
    );
nand_n_1369: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S557,
        in1(1) => S340,
        out1 => S559
    );
nor_n_842: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S558,
        in1(1) => S270,
        out1 => S560
    );
nand_n_1370: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S559,
        in1(1) => S271,
        out1 => S561
    );
nor_n_843: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S560,
        in1(1) => S268,
        out1 => S562
    );
nand_n_1371: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S561,
        in1(1) => S267,
        out1 => S563
    );
nor_n_844: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S562,
        in1(1) => S192,
        out1 => S564
    );
nand_n_1372: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S563,
        in1(1) => S193,
        out1 => S565
    );
nor_n_845: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S564,
        in1(1) => S190,
        out1 => S566
    );
nand_n_1373: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S565,
        in1(1) => S189,
        out1 => S567
    );
nor_n_846: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S566,
        in1(1) => S2594,
        out1 => S568
    );
nand_n_1374: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S567,
        in1(1) => S2595,
        out1 => S569
    );
nor_n_847: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S568,
        in1(1) => S2592,
        out1 => S570
    );
nand_n_1375: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S569,
        in1(1) => S2591,
        out1 => S571
    );
nor_n_848: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S570,
        in1(1) => S2515,
        out1 => S572
    );
nand_n_1376: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S571,
        in1(1) => S2516,
        out1 => S573
    );
nor_n_849: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S572,
        in1(1) => S2513,
        out1 => S574
    );
nand_n_1377: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S573,
        in1(1) => S2512,
        out1 => S575
    );
nor_n_850: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S574,
        in1(1) => S2437,
        out1 => S576
    );
nand_n_1378: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S575,
        in1(1) => S2438,
        out1 => S577
    );
nor_n_851: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S576,
        in1(1) => S2435,
        out1 => S578
    );
nand_n_1379: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S577,
        in1(1) => S2434,
        out1 => S579
    );
nand_n_1380: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2419,
        in1(1) => S2294,
        out1 => S580
    );
notg_254: ENTITY WORK.notg
    PORT MAP (
        in1 => S580,
        out1 => S581
    );
nor_n_852: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2429,
        in1(1) => S2424,
        out1 => S582
    );
notg_255: ENTITY WORK.notg
    PORT MAP (
        in1 => S582,
        out1 => S583
    );
nor_n_853: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S583,
        in1(1) => S580,
        out1 => S584
    );
nand_n_1381: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S582,
        in1(1) => S581,
        out1 => S585
    );
nor_n_854: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S582,
        in1(1) => S581,
        out1 => S586
    );
nand_n_1382: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S583,
        in1(1) => S580,
        out1 => S587
    );
nor_n_855: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S586,
        in1(1) => S584,
        out1 => S588
    );
nand_n_1383: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S587,
        in1(1) => S585,
        out1 => S589
    );
nor_n_856: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S588,
        in1(1) => S578,
        out1 => S590
    );
nand_n_1384: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S589,
        in1(1) => S579,
        out1 => S591
    );
nand_n_1385: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S582,
        in1(1) => S2294,
        out1 => S592
    );
nand_n_1386: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S592,
        in1(1) => S2419,
        out1 => S593
    );
notg_256: ENTITY WORK.notg
    PORT MAP (
        in1 => S593,
        out1 => S594
    );
nor_n_857: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S594,
        in1(1) => S590,
        out1 => S595
    );
nand_n_1387: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S593,
        in1(1) => S591,
        out1 => S596
    );
nor_n_858: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_ADD,
        in1(1) => S1994,
        out1 => S597
    );
nand_n_1388: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1995,
        in1(1) => U1_MUL,
        out1 => S598
    );
nor_n_859: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S598,
        in1(1) => S595,
        out1 => S599
    );
nand_n_1389: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S597,
        in1(1) => S596,
        out1 => S600
    );
nand_n_1390: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2106,
        in1(1) => U1_selMO_ARU,
        out1 => S601
    );
nand_n_1391: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2106,
        in1(1) => U1_AC_out_14,
        out1 => S602
    );
notg_257: ENTITY WORK.notg
    PORT MAP (
        in1 => S602,
        out1 => S603
    );
nand_n_1392: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S603,
        in1(1) => U1_selMO_ARU,
        out1 => S604
    );
notg_258: ENTITY WORK.notg
    PORT MAP (
        in1 => S604,
        out1 => S605
    );
nand_n_1393: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S601,
        in1(1) => S1902,
        out1 => S606
    );
nand_n_1394: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S606,
        in1(1) => S604,
        out1 => S607
    );
nand_n_1395: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2116,
        in1(1) => U1_AC_out_13,
        out1 => S608
    );
nand_n_1396: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2116,
        in1(1) => U1_selMO_ARU,
        out1 => S609
    );
notg_259: ENTITY WORK.notg
    PORT MAP (
        in1 => S609,
        out1 => S610
    );
nor_n_860: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S608,
        in1(1) => S1993,
        out1 => S611
    );
nor_n_861: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S610,
        in1(1) => U1_AC_out_13,
        out1 => S612
    );
nand_n_1397: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2125,
        in1(1) => U1_AC_out_12,
        out1 => S613
    );
nand_n_1398: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2125,
        in1(1) => U1_selMO_ARU,
        out1 => S614
    );
notg_260: ENTITY WORK.notg
    PORT MAP (
        in1 => S614,
        out1 => S615
    );
nor_n_862: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S613,
        in1(1) => S1993,
        out1 => S616
    );
nand_n_1399: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S615,
        in1(1) => U1_AC_out_12,
        out1 => S617
    );
nor_n_863: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S615,
        in1(1) => U1_AC_out_12,
        out1 => S618
    );
nor_n_864: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S618,
        in1(1) => S616,
        out1 => S619
    );
nand_n_1400: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2053,
        in1(1) => U1_selMO_ARU,
        out1 => S620
    );
notg_261: ENTITY WORK.notg
    PORT MAP (
        in1 => S620,
        out1 => S621
    );
nor_n_865: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S621,
        in1(1) => U1_AC_out_11,
        out1 => S622
    );
nand_n_1401: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2053,
        in1(1) => U1_AC_out_11,
        out1 => S623
    );
nor_n_866: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S623,
        in1(1) => S1993,
        out1 => S624
    );
nand_n_1402: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2061,
        in1(1) => U1_AC_out_10,
        out1 => S625
    );
notg_262: ENTITY WORK.notg
    PORT MAP (
        in1 => S625,
        out1 => S626
    );
nand_n_1403: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2061,
        in1(1) => U1_selMO_ARU,
        out1 => S627
    );
nand_n_1404: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S626,
        in1(1) => U1_selMO_ARU,
        out1 => S628
    );
nand_n_1405: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S627,
        in1(1) => S1892,
        out1 => S629
    );
nand_n_1406: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S629,
        in1(1) => S628,
        out1 => S630
    );
nand_n_1407: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2073,
        in1(1) => U1_selMO_ARU,
        out1 => S631
    );
notg_263: ENTITY WORK.notg
    PORT MAP (
        in1 => S631,
        out1 => S632
    );
nor_n_867: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S632,
        in1(1) => U1_AC_out_9,
        out1 => S633
    );
nand_n_1408: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2073,
        in1(1) => U1_AC_out_9,
        out1 => S634
    );
nor_n_868: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S634,
        in1(1) => S1993,
        out1 => S635
    );
nand_n_1409: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2082,
        in1(1) => U1_AC_out_8,
        out1 => S636
    );
nand_n_1410: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2082,
        in1(1) => U1_selMO_ARU,
        out1 => S637
    );
notg_264: ENTITY WORK.notg
    PORT MAP (
        in1 => S637,
        out1 => S638
    );
nor_n_869: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S636,
        in1(1) => S1993,
        out1 => S639
    );
nand_n_1411: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S638,
        in1(1) => U1_AC_out_8,
        out1 => S640
    );
nor_n_870: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S638,
        in1(1) => U1_AC_out_8,
        out1 => S641
    );
nor_n_871: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S641,
        in1(1) => S639,
        out1 => S642
    );
nor_n_872: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2305,
        in1(1) => U1_AC_out_7,
        out1 => S643
    );
nor_n_873: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2283,
        in1(1) => U1_AC_out_6,
        out1 => S644
    );
nor_n_874: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S644,
        in1(1) => S2296,
        out1 => S645
    );
nor_n_875: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2271,
        in1(1) => U1_AC_out_5,
        out1 => S646
    );
nor_n_876: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S646,
        in1(1) => S2330,
        out1 => S647
    );
nor_n_877: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2274,
        in1(1) => U1_AC_out_4,
        out1 => S648
    );
nor_n_878: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S648,
        in1(1) => S2547,
        out1 => S649
    );
nand_n_1412: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2322,
        in1(1) => S1939,
        out1 => S650
    );
nor_n_879: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2360,
        in1(1) => U1_AC_out_2,
        out1 => S651
    );
nor_n_880: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S651,
        in1(1) => S362,
        out1 => S652
    );
nor_n_881: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2517,
        in1(1) => S1917,
        out1 => S653
    );
nor_n_882: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2442,
        in1(1) => U1_AC_out_1,
        out1 => S654
    );
nor_n_883: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S654,
        in1(1) => S498,
        out1 => S655
    );
nand_n_1413: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S655,
        in1(1) => S653,
        out1 => S656
    );
nand_n_1414: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S656,
        in1(1) => S499,
        out1 => S657
    );
nand_n_1415: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S657,
        in1(1) => S652,
        out1 => S658
    );
nand_n_1416: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S658,
        in1(1) => S363,
        out1 => S659
    );
nand_n_1417: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S659,
        in1(1) => S650,
        out1 => S660
    );
nand_n_1418: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S660,
        in1(1) => S2615,
        out1 => S661
    );
nand_n_1419: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S661,
        in1(1) => S649,
        out1 => S662
    );
notg_265: ENTITY WORK.notg
    PORT MAP (
        in1 => S662,
        out1 => S663
    );
nand_n_1420: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S662,
        in1(1) => S2548,
        out1 => S664
    );
nand_n_1421: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S664,
        in1(1) => S647,
        out1 => S665
    );
nand_n_1422: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S665,
        in1(1) => S2331,
        out1 => S666
    );
nand_n_1423: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S666,
        in1(1) => S645,
        out1 => S667
    );
nand_n_1424: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S667,
        in1(1) => S2297,
        out1 => S668
    );
nor_n_884: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S668,
        in1(1) => S2419,
        out1 => S669
    );
nor_n_885: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S669,
        in1(1) => S643,
        out1 => S670
    );
nand_n_1425: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S670,
        in1(1) => S642,
        out1 => S671
    );
nand_n_1426: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S671,
        in1(1) => S640,
        out1 => S672
    );
notg_266: ENTITY WORK.notg
    PORT MAP (
        in1 => S672,
        out1 => S673
    );
nor_n_886: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S673,
        in1(1) => S633,
        out1 => S674
    );
nor_n_887: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S674,
        in1(1) => S635,
        out1 => S675
    );
nor_n_888: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S675,
        in1(1) => S630,
        out1 => S676
    );
notg_267: ENTITY WORK.notg
    PORT MAP (
        in1 => S676,
        out1 => S677
    );
nand_n_1427: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S677,
        in1(1) => S628,
        out1 => S678
    );
nor_n_889: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S678,
        in1(1) => S624,
        out1 => S679
    );
nor_n_890: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S679,
        in1(1) => S622,
        out1 => S680
    );
nand_n_1428: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S680,
        in1(1) => S619,
        out1 => S681
    );
nand_n_1429: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S681,
        in1(1) => S617,
        out1 => S682
    );
notg_268: ENTITY WORK.notg
    PORT MAP (
        in1 => S682,
        out1 => S683
    );
nor_n_891: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S683,
        in1(1) => S612,
        out1 => S684
    );
nor_n_892: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S684,
        in1(1) => S611,
        out1 => S685
    );
nor_n_893: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S685,
        in1(1) => S607,
        out1 => S686
    );
notg_269: ENTITY WORK.notg
    PORT MAP (
        in1 => S686,
        out1 => S687
    );
nor_n_894: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S686,
        in1(1) => S605,
        out1 => S688
    );
nand_n_1430: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S687,
        in1(1) => S604,
        out1 => S689
    );
nand_n_1431: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2268,
        in1(1) => S1909,
        out1 => S690
    );
nand_n_1432: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S690,
        in1(1) => S2269,
        out1 => S691
    );
notg_270: ENTITY WORK.notg
    PORT MAP (
        in1 => S691,
        out1 => S692
    );
nor_n_895: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S691,
        in1(1) => S688,
        out1 => S693
    );
nor_n_896: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S692,
        in1(1) => S689,
        out1 => S694
    );
nand_n_1433: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S691,
        in1(1) => S688,
        out1 => S695
    );
nand_n_1434: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S695,
        in1(1) => U1_ADD,
        out1 => S696
    );
nor_n_897: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S694,
        in1(1) => S693,
        out1 => S697
    );
nor_n_898: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S696,
        in1(1) => S693,
        out1 => S698
    );
nand_n_1435: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S697,
        in1(1) => U1_ADD,
        out1 => S699
    );
nor_n_899: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S698,
        in1(1) => S599,
        out1 => S700
    );
nand_n_1436: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S699,
        in1(1) => S600,
        out1 => S701
    );
nor_n_900: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S701,
        in1(1) => S2269,
        out1 => S702
    );
nor_n_901: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S700,
        in1(1) => S690,
        out1 => S703
    );
nor_n_902: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S703,
        in1(1) => S702,
        out1 => S704
    );
notg_271: ENTITY WORK.notg
    PORT MAP (
        in1 => S704,
        out1 => U1_V
    );
nor_n_903: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S689,
        in1(1) => S2270,
        out1 => S705
    );
nor_n_904: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S705,
        in1(1) => S1995,
        out1 => S706
    );
nand_n_1437: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S706,
        in1(1) => S690,
        out1 => S707
    );
notg_272: ENTITY WORK.notg
    PORT MAP (
        in1 => S707,
        out1 => U1_C
    );
nand_n_1438: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2094,
        in1(1) => U1_AC_out_0,
        out1 => S708
    );
nor_n_905: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2108,
        in1(1) => U1_AC_out_0,
        out1 => S709
    );
notg_273: ENTITY WORK.notg
    PORT MAP (
        in1 => S709,
        out1 => S710
    );
nand_n_1439: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S710,
        in1(1) => S708,
        out1 => S711
    );
nor_n_906: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S711,
        in1(1) => U1_AC_out_1,
        out1 => S712
    );
nand_n_1440: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S712,
        in1(1) => S2099,
        out1 => S713
    );
nand_n_1441: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2119,
        in1(1) => U1_AC_out_0,
        out1 => S714
    );
nand_n_1442: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S714,
        in1(1) => S710,
        out1 => S715
    );
nand_n_1443: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S715,
        in1(1) => S1925,
        out1 => S716
    );
nand_n_1444: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2128,
        in1(1) => S1917,
        out1 => S717
    );
nand_n_1445: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2054,
        in1(1) => U1_AC_out_0,
        out1 => S718
    );
nand_n_1446: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S718,
        in1(1) => S717,
        out1 => S719
    );
nand_n_1447: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S719,
        in1(1) => U1_AC_out_1,
        out1 => S720
    );
nand_n_1448: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S720,
        in1(1) => S716,
        out1 => S721
    );
nand_n_1449: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S721,
        in1(1) => S1932,
        out1 => S722
    );
nand_n_1450: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2064,
        in1(1) => S1917,
        out1 => S723
    );
nand_n_1451: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2074,
        in1(1) => U1_AC_out_0,
        out1 => S724
    );
nand_n_1452: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S724,
        in1(1) => S723,
        out1 => S725
    );
nand_n_1453: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S725,
        in1(1) => S1925,
        out1 => S726
    );
nand_n_1454: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2083,
        in1(1) => S1917,
        out1 => S727
    );
nand_n_1455: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2201,
        in1(1) => U1_AC_out_0,
        out1 => S728
    );
nand_n_1456: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S728,
        in1(1) => S727,
        out1 => S729
    );
nand_n_1457: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S729,
        in1(1) => U1_AC_out_1,
        out1 => S730
    );
nand_n_1458: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S730,
        in1(1) => S726,
        out1 => S731
    );
nand_n_1459: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S731,
        in1(1) => U1_AC_out_2,
        out1 => S732
    );
nand_n_1460: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S732,
        in1(1) => S722,
        out1 => S733
    );
nand_n_1461: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S733,
        in1(1) => S1939,
        out1 => S734
    );
nand_n_1462: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S734,
        in1(1) => S2029,
        out1 => S735
    );
nand_n_1463: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S735,
        in1(1) => S713,
        out1 => S736
    );
nor_n_907: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2161,
        in1(1) => U1_AC_out_0,
        out1 => S737
    );
nor_n_908: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2175,
        in1(1) => S1917,
        out1 => S738
    );
nor_n_909: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S738,
        in1(1) => S737,
        out1 => S739
    );
nor_n_910: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S739,
        in1(1) => U1_AC_out_1,
        out1 => S740
    );
notg_274: ENTITY WORK.notg
    PORT MAP (
        in1 => S740,
        out1 => S741
    );
nor_n_911: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2186,
        in1(1) => U1_AC_out_0,
        out1 => S742
    );
nand_n_1464: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2187,
        in1(1) => S1917,
        out1 => S743
    );
nand_n_1465: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S743,
        in1(1) => U1_AC_out_1,
        out1 => S744
    );
nand_n_1466: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S744,
        in1(1) => S741,
        out1 => S745
    );
nand_n_1467: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2210,
        in1(1) => S1917,
        out1 => S746
    );
nand_n_1468: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2221,
        in1(1) => U1_AC_out_0,
        out1 => S747
    );
nand_n_1469: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S747,
        in1(1) => S746,
        out1 => S748
    );
notg_275: ENTITY WORK.notg
    PORT MAP (
        in1 => S748,
        out1 => S749
    );
nor_n_912: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S749,
        in1(1) => U1_AC_out_1,
        out1 => S750
    );
nor_n_913: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2150,
        in1(1) => S1917,
        out1 => S751
    );
nor_n_914: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2234,
        in1(1) => U1_AC_out_0,
        out1 => S752
    );
notg_276: ENTITY WORK.notg
    PORT MAP (
        in1 => S752,
        out1 => S753
    );
nor_n_915: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S752,
        in1(1) => S751,
        out1 => S754
    );
dff_1: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S70,
        NbarT => '0',
        PRE => '0',
        Q => U1_OF_out_0,
        Si => S2834,
        global_reset => '0'
    );
dff_2: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S71,
        NbarT => '0',
        PRE => '0',
        Q => U1_OF_out_1,
        Si => S2835,
        global_reset => '0'
    );
dff_3: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S72,
        NbarT => '0',
        PRE => '0',
        Q => U1_OF_out_2,
        Si => S2836,
        global_reset => '0'
    );
dff_4: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S73,
        NbarT => '0',
        PRE => '0',
        Q => U1_OF_out_3,
        Si => S2837,
        global_reset => '0'
    );
dff_5: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S74,
        NbarT => '0',
        PRE => '0',
        Q => U1_AC_out_0,
        Si => S2838,
        global_reset => '0'
    );
dff_6: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S75,
        NbarT => '0',
        PRE => '0',
        Q => U1_AC_out_1,
        Si => S2839,
        global_reset => '0'
    );
dff_7: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S76,
        NbarT => '0',
        PRE => '0',
        Q => U1_AC_out_2,
        Si => S2840,
        global_reset => '0'
    );
dff_8: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S77,
        NbarT => '0',
        PRE => '0',
        Q => U1_AC_out_3,
        Si => S2841,
        global_reset => '0'
    );
dff_9: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S78,
        NbarT => '0',
        PRE => '0',
        Q => U1_AC_out_4,
        Si => S2842,
        global_reset => '0'
    );
dff_10: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S79,
        NbarT => '0',
        PRE => '0',
        Q => U1_AC_out_5,
        Si => S2843,
        global_reset => '0'
    );
dff_11: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S80,
        NbarT => '0',
        PRE => '0',
        Q => U1_AC_out_6,
        Si => S2844,
        global_reset => '0'
    );
dff_12: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S81,
        NbarT => '0',
        PRE => '0',
        Q => U1_AC_out_7,
        Si => S2845,
        global_reset => '0'
    );
dff_13: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S82,
        NbarT => '0',
        PRE => '0',
        Q => U1_AC_out_8,
        Si => S2846,
        global_reset => '0'
    );
dff_14: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S83,
        NbarT => '0',
        PRE => '0',
        Q => U1_AC_out_9,
        Si => S2847,
        global_reset => '0'
    );
dff_15: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S84,
        NbarT => '0',
        PRE => '0',
        Q => U1_AC_out_10,
        Si => S2848,
        global_reset => '0'
    );
dff_16: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S85,
        NbarT => '0',
        PRE => '0',
        Q => U1_AC_out_11,
        Si => S2849,
        global_reset => '0'
    );
dff_17: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S86,
        NbarT => '0',
        PRE => '0',
        Q => U1_AC_out_12,
        Si => S2850,
        global_reset => '0'
    );
dff_18: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S87,
        NbarT => '0',
        PRE => '0',
        Q => U1_AC_out_13,
        Si => S2851,
        global_reset => '0'
    );
dff_19: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S88,
        NbarT => '0',
        PRE => '0',
        Q => U1_AC_out_14,
        Si => S2852,
        global_reset => '0'
    );
dff_20: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S89,
        NbarT => '0',
        PRE => '0',
        Q => U1_AC_out_15,
        Si => S2853,
        global_reset => '0'
    );
dff_21: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S90,
        NbarT => '0',
        PRE => '0',
        Q => U1_V_out1,
        Si => S2854,
        global_reset => '0'
    );
dff_22: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S91,
        NbarT => '0',
        PRE => '0',
        Q => U1_C_out1,
        Si => S2855,
        global_reset => '0'
    );
dff_23: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S92,
        NbarT => '0',
        PRE => '0',
        Q => U1_N_out1,
        Si => S2856,
        global_reset => '0'
    );
dff_24: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S93,
        NbarT => '0',
        PRE => '0',
        Q => U1_Z_out1,
        Si => S2857,
        global_reset => '0'
    );
dff_25: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S94,
        NbarT => '0',
        PRE => '0',
        Q => U1_IN_out_0,
        Si => S2858,
        global_reset => '0'
    );
dff_26: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S95,
        NbarT => '0',
        PRE => '0',
        Q => U1_IN_out_1,
        Si => S2859,
        global_reset => '0'
    );
dff_27: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S96,
        NbarT => '0',
        PRE => '0',
        Q => U1_IN_out_2,
        Si => S2860,
        global_reset => '0'
    );
dff_28: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S97,
        NbarT => '0',
        PRE => '0',
        Q => U1_IN_out_3,
        Si => S2861,
        global_reset => '0'
    );
dff_29: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S98,
        NbarT => '0',
        PRE => '0',
        Q => U1_IN_out_4,
        Si => S2862,
        global_reset => '0'
    );
dff_30: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S99,
        NbarT => '0',
        PRE => '0',
        Q => U1_IN_out_5,
        Si => S2863,
        global_reset => '0'
    );
dff_31: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S100,
        NbarT => '0',
        PRE => '0',
        Q => U1_IN_out_6,
        Si => S2864,
        global_reset => '0'
    );
dff_32: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S101,
        NbarT => '0',
        PRE => '0',
        Q => U1_IN_out_7,
        Si => S2865,
        global_reset => '0'
    );
dff_33: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S102,
        NbarT => '0',
        PRE => '0',
        Q => U1_IN_out_8,
        Si => S2866,
        global_reset => '0'
    );
dff_34: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S103,
        NbarT => '0',
        PRE => '0',
        Q => U1_IN_out_9,
        Si => S2867,
        global_reset => '0'
    );
dff_35: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S104,
        NbarT => '0',
        PRE => '0',
        Q => U1_IN_out_10,
        Si => S2868,
        global_reset => '0'
    );
dff_36: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S105,
        NbarT => '0',
        PRE => '0',
        Q => U1_IN_out_11,
        Si => S2869,
        global_reset => '0'
    );
dff_37: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S106,
        NbarT => '0',
        PRE => '0',
        Q => U1_IN_out_12,
        Si => S2870,
        global_reset => '0'
    );
dff_38: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S107,
        NbarT => '0',
        PRE => '0',
        Q => U1_IN_out_13,
        Si => S2871,
        global_reset => '0'
    );
dff_39: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S108,
        NbarT => '0',
        PRE => '0',
        Q => U1_IN_out_14,
        Si => S2872,
        global_reset => '0'
    );
dff_40: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S109,
        NbarT => '0',
        PRE => '0',
        Q => U1_IN_out_15,
        Si => S2873,
        global_reset => '0'
    );
dff_41: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S110,
        NbarT => '0',
        PRE => '0',
        Q => U1_PC_out_0,
        Si => S2874,
        global_reset => '0'
    );
dff_42: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S111,
        NbarT => '0',
        PRE => '0',
        Q => U1_PC_out_1,
        Si => S2875,
        global_reset => '0'
    );
dff_43: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S112,
        NbarT => '0',
        PRE => '0',
        Q => U1_PC_out_2,
        Si => S2876,
        global_reset => '0'
    );
dff_44: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S113,
        NbarT => '0',
        PRE => '0',
        Q => U1_PC_out_3,
        Si => S2877,
        global_reset => '0'
    );
dff_45: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S114,
        NbarT => '0',
        PRE => '0',
        Q => U1_PC_out_4,
        Si => S2878,
        global_reset => '0'
    );
dff_46: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S115,
        NbarT => '0',
        PRE => '0',
        Q => U1_PC_out_5,
        Si => S2879,
        global_reset => '0'
    );
dff_47: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S116,
        NbarT => '0',
        PRE => '0',
        Q => U1_PC_out_6,
        Si => S2880,
        global_reset => '0'
    );
dff_48: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S117,
        NbarT => '0',
        PRE => '0',
        Q => U1_PC_out_7,
        Si => S2881,
        global_reset => '0'
    );
dff_49: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S118,
        NbarT => '0',
        PRE => '0',
        Q => U1_PC_out_8,
        Si => S2882,
        global_reset => '0'
    );
dff_50: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S119,
        NbarT => '0',
        PRE => '0',
        Q => U1_PC_out_9,
        Si => S2883,
        global_reset => '0'
    );
dff_51: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S120,
        NbarT => '0',
        PRE => '0',
        Q => U1_PC_out_10,
        Si => S2884,
        global_reset => '0'
    );
dff_52: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S121,
        NbarT => '0',
        PRE => '0',
        Q => U1_PC_out_11,
        Si => S2885,
        global_reset => '0'
    );
dff_53: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S122,
        NbarT => '0',
        PRE => '0',
        Q => U1_PC_out_12,
        Si => S2886,
        global_reset => '0'
    );
dff_54: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S123,
        NbarT => '0',
        PRE => '0',
        Q => U1_PC_out_13,
        Si => S2887,
        global_reset => '0'
    );
dff_55: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S124,
        NbarT => '0',
        PRE => '0',
        Q => U1_PC_out_14,
        Si => S2888,
        global_reset => '0'
    );
dff_56: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S125,
        NbarT => '0',
        PRE => '0',
        Q => U1_PC_out_15,
        Si => S2889,
        global_reset => '0'
    );
dff_57: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S126,
        NbarT => '0',
        PRE => '0',
        Q => U1_IR_out_0,
        Si => S2890,
        global_reset => '0'
    );
dff_58: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S127,
        NbarT => '0',
        PRE => '0',
        Q => U1_IR_out_1,
        Si => S2891,
        global_reset => '0'
    );
dff_59: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S128,
        NbarT => '0',
        PRE => '0',
        Q => U1_IR_out_2,
        Si => S2892,
        global_reset => '0'
    );
dff_60: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S129,
        NbarT => '0',
        PRE => '0',
        Q => U1_IR_out_3,
        Si => S2893,
        global_reset => '0'
    );
dff_61: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S130,
        NbarT => '0',
        PRE => '0',
        Q => U1_IR_out_4,
        Si => S2894,
        global_reset => '0'
    );
dff_62: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S131,
        NbarT => '0',
        PRE => '0',
        Q => U1_IR_out_5,
        Si => S2895,
        global_reset => '0'
    );
dff_63: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S132,
        NbarT => '0',
        PRE => '0',
        Q => U1_IR_out_6,
        Si => S2896,
        global_reset => '0'
    );
dff_64: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S133,
        NbarT => '0',
        PRE => '0',
        Q => U1_IR_out_7,
        Si => S2897,
        global_reset => '0'
    );
dff_65: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S134,
        NbarT => '0',
        PRE => '0',
        Q => U1_IR_out_8,
        Si => S2898,
        global_reset => '0'
    );
dff_66: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S135,
        NbarT => '0',
        PRE => '0',
        Q => U1_IR_out_9,
        Si => S2899,
        global_reset => '0'
    );
dff_67: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S136,
        NbarT => '0',
        PRE => '0',
        Q => U1_IR_out_10,
        Si => S2900,
        global_reset => '0'
    );
dff_68: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S137,
        NbarT => '0',
        PRE => '0',
        Q => U1_IR_out_11,
        Si => S2901,
        global_reset => '0'
    );
dff_69: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S138,
        NbarT => '0',
        PRE => '0',
        Q => U1_IR_out_12,
        Si => S2902,
        global_reset => '0'
    );
dff_70: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S139,
        NbarT => '0',
        PRE => '0',
        Q => U1_IR_out_13,
        Si => S2903,
        global_reset => '0'
    );
dff_71: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S140,
        NbarT => '0',
        PRE => '0',
        Q => U1_IR_out_14,
        Si => S2904,
        global_reset => '0'
    );
dff_72: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => S141,
        NbarT => '0',
        PRE => '0',
        Q => U1_IR_out_15,
        Si => S2905,
        global_reset => '0'
    );
notg_277: ENTITY WORK.notg
    PORT MAP (
        in1 => S2623,
        out1 => S2796
    );
notg_278: ENTITY WORK.notg
    PORT MAP (
        in1 => U2_pstate,
        out1 => S2797
    );
notg_279: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_IR_out_9,
        out1 => S2798
    );
notg_280: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_IR_out_8,
        out1 => S2799
    );
notg_281: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_IR_out_11,
        out1 => S2800
    );
notg_282: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_IR_out_10,
        out1 => S2801
    );
notg_283: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_IR_out_13,
        out1 => S2802
    );
notg_284: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_IR_out_12,
        out1 => S2803
    );
notg_285: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_IR_out_14,
        out1 => S2804
    );
notg_286: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_IR_out_0,
        out1 => S2805
    );
notg_287: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_IR_out_3,
        out1 => S2806
    );
notg_288: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_IR_out_2,
        out1 => S2807
    );
notg_289: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_IR_out_5,
        out1 => S2808
    );
notg_290: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_IR_out_6,
        out1 => S2809
    );
nor_n_916: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U2_pstate,
        in1(1) => S2623,
        out1 => U1_ldIR
    );
notg_291: ENTITY WORK.notg
    PORT MAP (
        in1 => U1_ldIR,
        out1 => S2810
    );
nor_n_917: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2801,
        in1(1) => U1_IR_out_11,
        out1 => S2811
    );
nand_n_1470: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_IR_out_10,
        in1(1) => S2800,
        out1 => S2812
    );
nor_n_918: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_IR_out_8,
        in1(1) => U1_IR_out_9,
        out1 => S2813
    );
notg_292: ENTITY WORK.notg
    PORT MAP (
        in1 => S2813,
        out1 => S2814
    );
nor_n_919: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2814,
        in1(1) => S2812,
        out1 => S2815
    );
nand_n_1471: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2813,
        in1(1) => S2811,
        out1 => S2816
    );
nor_n_920: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2797,
        in1(1) => S2623,
        out1 => S2817
    );
nand_n_1472: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U2_pstate,
        in1(1) => S2796,
        out1 => S2818
    );
nand_n_1473: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_IR_out_14,
        in1(1) => U1_IR_out_15,
        out1 => S2819
    );
notg_293: ENTITY WORK.notg
    PORT MAP (
        in1 => S2819,
        out1 => S2820
    );
nand_n_1474: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_IR_out_12,
        in1(1) => U1_IR_out_13,
        out1 => S2821
    );
notg_294: ENTITY WORK.notg
    PORT MAP (
        in1 => S2821,
        out1 => S2822
    );
nor_n_921: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2821,
        in1(1) => S2819,
        out1 => S2823
    );
nand_n_1475: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2822,
        in1(1) => S2820,
        out1 => S2824
    );
nor_n_922: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2824,
        in1(1) => S2818,
        out1 => S2825
    );
nand_n_1476: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2823,
        in1(1) => S2817,
        out1 => S2826
    );
nor_n_923: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2826,
        in1(1) => S2816,
        out1 => U1_SHF_0
    );
nor_n_924: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_IR_out_10,
        in1(1) => U1_IR_out_11,
        out1 => S2827
    );
notg_295: ENTITY WORK.notg
    PORT MAP (
        in1 => S2827,
        out1 => S2828
    );
nor_n_925: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2828,
        in1(1) => S2798,
        out1 => S2829
    );
nand_n_1477: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2827,
        in1(1) => U1_IR_out_9,
        out1 => S2830
    );
nand_n_1478: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2829,
        in1(1) => U1_IR_out_8,
        out1 => S2831
    );
nor_n_926: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2831,
        in1(1) => S2826,
        out1 => U1_SHF_1
    );
nor_n_927: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_IR_out_12,
        in1(1) => S2802,
        out1 => S2624
    );
nand_n_1479: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2803,
        in1(1) => U1_IR_out_13,
        out1 => S2625
    );
nand_n_1480: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_IR_out_15,
        in1(1) => S2803,
        out1 => S2626
    );
nor_n_928: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2804,
        in1(1) => S2802,
        out1 => S2627
    );
nand_n_1481: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_IR_out_14,
        in1(1) => U1_IR_out_13,
        out1 => S2628
    );
nor_n_929: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2628,
        in1(1) => S2626,
        out1 => S2629
    );
nand_n_1482: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2627,
        in1(1) => S2817,
        out1 => S2630
    );
nand_n_1483: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2629,
        in1(1) => S2817,
        out1 => S2631
    );
nand_n_1484: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2631,
        in1(1) => S2810,
        out1 => U1_selPC_MEM
    );
nor_n_930: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_IR_out_14,
        in1(1) => U1_IR_out_15,
        out1 => S2632
    );
notg_296: ENTITY WORK.notg
    PORT MAP (
        in1 => S2632,
        out1 => S2633
    );
nand_n_1485: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2632,
        in1(1) => U1_IR_out_12,
        out1 => S2634
    );
notg_297: ENTITY WORK.notg
    PORT MAP (
        in1 => S2634,
        out1 => S2635
    );
nor_n_931: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2634,
        in1(1) => S2802,
        out1 => S2636
    );
notg_298: ENTITY WORK.notg
    PORT MAP (
        in1 => S2636,
        out1 => S2637
    );
nor_n_932: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2636,
        in1(1) => S2629,
        out1 => S2638
    );
notg_299: ENTITY WORK.notg
    PORT MAP (
        in1 => S2638,
        out1 => S2639
    );
nor_n_933: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2804,
        in1(1) => U1_IR_out_15,
        out1 => S2640
    );
nor_n_934: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2628,
        in1(1) => U1_IR_out_15,
        out1 => S2641
    );
nand_n_1486: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2640,
        in1(1) => U1_IR_out_13,
        out1 => S2642
    );
nand_n_1487: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2804,
        in1(1) => U1_IR_out_15,
        out1 => S2643
    );
nor_n_935: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2643,
        in1(1) => U1_IR_out_13,
        out1 => S2644
    );
nor_n_936: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2644,
        in1(1) => S2641,
        out1 => S2645
    );
nor_n_937: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2645,
        in1(1) => U1_IR_out_12,
        out1 => S2646
    );
nor_n_938: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2646,
        in1(1) => S2639,
        out1 => S2647
    );
nor_n_939: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2633,
        in1(1) => U1_IR_out_13,
        out1 => S2648
    );
notg_300: ENTITY WORK.notg
    PORT MAP (
        in1 => S2648,
        out1 => S2649
    );
nand_n_1488: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2648,
        in1(1) => S2803,
        out1 => S2650
    );
nor_n_940: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2823,
        in1(1) => S2818,
        out1 => S2651
    );
nand_n_1489: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2651,
        in1(1) => S2650,
        out1 => S2652
    );
nor_n_941: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2819,
        in1(1) => U1_IR_out_13,
        out1 => S2653
    );
notg_301: ENTITY WORK.notg
    PORT MAP (
        in1 => S2653,
        out1 => S2654
    );
nor_n_942: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2819,
        in1(1) => U1_IR_out_12,
        out1 => S2655
    );
nor_n_943: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2654,
        in1(1) => U1_IR_out_12,
        out1 => S2656
    );
nor_n_944: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2656,
        in1(1) => S2652,
        out1 => S2657
    );
nand_n_1490: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2657,
        in1(1) => S2647,
        out1 => S2658
    );
nand_n_1491: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2797,
        in1(1) => S2623,
        out1 => S2659
    );
nor_n_945: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2659,
        in1(1) => S2625,
        out1 => S2660
    );
notg_302: ENTITY WORK.notg
    PORT MAP (
        in1 => S2660,
        out1 => S2661
    );
nor_n_946: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2661,
        in1(1) => U1_IR_out_14,
        out1 => S2662
    );
notg_303: ENTITY WORK.notg
    PORT MAP (
        in1 => S2662,
        out1 => S2663
    );
nor_n_947: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2662,
        in1(1) => U1_ldIR,
        out1 => S2664
    );
nand_n_1492: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2664,
        in1(1) => S2658,
        out1 => U2_readMEM
    );
nand_n_1493: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2642,
        in1(1) => S2817,
        out1 => S2665
    );
nor_n_948: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2640,
        in1(1) => S2624,
        out1 => S2666
    );
notg_304: ENTITY WORK.notg
    PORT MAP (
        in1 => S2666,
        out1 => S2667
    );
nor_n_949: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2666,
        in1(1) => S2665,
        out1 => U2_nstate_1
    );
nor_n_950: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2627,
        in1(1) => U1_IR_out_15,
        out1 => S2668
    );
nor_n_951: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2668,
        in1(1) => S2629,
        out1 => S2669
    );
notg_305: ENTITY WORK.notg
    PORT MAP (
        in1 => S2669,
        out1 => S2670
    );
nand_n_1494: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2653,
        in1(1) => U1_IR_out_12,
        out1 => S2671
    );
nand_n_1495: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2671,
        in1(1) => S2669,
        out1 => S2672
    );
nand_n_1496: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2672,
        in1(1) => S2817,
        out1 => S2673
    );
nor_n_952: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2661,
        in1(1) => S2819,
        out1 => S2674
    );
notg_306: ENTITY WORK.notg
    PORT MAP (
        in1 => S2674,
        out1 => S2675
    );
nand_n_1497: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2827,
        in1(1) => S2813,
        out1 => S2676
    );
nor_n_953: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2829,
        in1(1) => S2815,
        out1 => S2677
    );
nand_n_1498: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2830,
        in1(1) => S2816,
        out1 => S2678
    );
nand_n_1499: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2677,
        in1(1) => S2676,
        out1 => S2679
    );
nor_n_954: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_IR_out_8,
        in1(1) => S2798,
        out1 => S2680
    );
nand_n_1500: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2799,
        in1(1) => U1_IR_out_9,
        out1 => S2681
    );
nor_n_955: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2681,
        in1(1) => S2812,
        out1 => S2682
    );
nand_n_1501: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2680,
        in1(1) => S2811,
        out1 => S2683
    );
nor_n_956: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2682,
        in1(1) => S2679,
        out1 => S2684
    );
nand_n_1502: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2808,
        in1(1) => S2806,
        out1 => S2685
    );
nor_n_957: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_IR_out_7,
        in1(1) => U1_IR_out_4,
        out1 => S2686
    );
nand_n_1503: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2686,
        in1(1) => S2809,
        out1 => S2687
    );
nor_n_958: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_IR_out_6,
        in1(1) => U1_IR_out_4,
        out1 => S2688
    );
nor_n_959: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2685,
        in1(1) => U1_IR_out_7,
        out1 => S2689
    );
nor_n_960: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2687,
        in1(1) => S2685,
        out1 => S2690
    );
nand_n_1504: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2689,
        in1(1) => S2688,
        out1 => S2691
    );
nor_n_961: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2799,
        in1(1) => U1_IR_out_9,
        out1 => S2692
    );
nand_n_1505: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => U1_IR_out_8,
        in1(1) => S2798,
        out1 => S2693
    );
nor_n_962: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2693,
        in1(1) => S2828,
        out1 => S2694
    );
nand_n_1506: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2692,
        in1(1) => S2827,
        out1 => S2695
    );
nor_n_963: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_IR_out_0,
        in1(1) => U1_IR_out_1,
        out1 => S2696
    );
nand_n_1507: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2696,
        in1(1) => U1_IR_out_2,
        out1 => S2697
    );
nor_n_964: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2697,
        in1(1) => S2695,
        out1 => S2698
    );
nand_n_1508: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2698,
        in1(1) => S2690,
        out1 => S2699
    );
nand_n_1509: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2699,
        in1(1) => S2684,
        out1 => S2700
    );
nor_n_965: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2695,
        in1(1) => U1_IR_out_2,
        out1 => S2701
    );
nand_n_1510: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2694,
        in1(1) => S2807,
        out1 => S2702
    );
nor_n_966: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2702,
        in1(1) => S2691,
        out1 => S2703
    );
nand_n_1511: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2701,
        in1(1) => S2690,
        out1 => S2704
    );
nor_n_967: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2704,
        in1(1) => U1_IR_out_1,
        out1 => S2705
    );
nor_n_968: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2691,
        in1(1) => U1_IR_out_2,
        out1 => S2706
    );
nor_n_969: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2695,
        in1(1) => U1_IR_out_1,
        out1 => S2707
    );
nand_n_1512: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2707,
        in1(1) => S2706,
        out1 => S2708
    );
nor_n_970: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2705,
        in1(1) => S2700,
        out1 => S2709
    );
nor_n_971: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2709,
        in1(1) => S2826,
        out1 => S2710
    );
nor_n_972: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2710,
        in1(1) => S2674,
        out1 => S2711
    );
nand_n_1513: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2711,
        in1(1) => S2673,
        out1 => U1_INC1
    );
nand_n_1514: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2640,
        in1(1) => S2802,
        out1 => S2712
    );
nor_n_973: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2712,
        in1(1) => S2659,
        out1 => S2713
    );
notg_307: ENTITY WORK.notg
    PORT MAP (
        in1 => S2713,
        out1 => S2714
    );
nor_n_974: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2637,
        in1(1) => S2818,
        out1 => S2715
    );
nor_n_975: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2715,
        in1(1) => S2713,
        out1 => S2716
    );
nand_n_1515: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2716,
        in1(1) => S2631,
        out1 => U1_seldataBus
    );
nor_n_976: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2714,
        in1(1) => S2803,
        out1 => S2717
    );
nor_n_977: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2652,
        in1(1) => S2646,
        out1 => S2718
    );
nor_n_978: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2718,
        in1(1) => S2717,
        out1 => S2719
    );
notg_308: ENTITY WORK.notg
    PORT MAP (
        in1 => S2719,
        out1 => U1_conOF
    );
nor_n_979: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2719,
        in1(1) => S2656,
        out1 => U1_selIR_MEM
    );
nor_n_980: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2715,
        in1(1) => S2803,
        out1 => S2720
    );
nor_n_981: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2720,
        in1(1) => S2716,
        out1 => U1_selAC_MEM
    );
nor_n_982: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2812,
        in1(1) => U1_enSKP,
        out1 => S2721
    );
nand_n_1516: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2721,
        in1(1) => S2692,
        out1 => S2722
    );
nand_n_1517: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2722,
        in1(1) => S2823,
        out1 => S2723
    );
notg_309: ENTITY WORK.notg
    PORT MAP (
        in1 => S2723,
        out1 => S2724
    );
nand_n_1518: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2724,
        in1(1) => S2709,
        out1 => S2725
    );
nand_n_1519: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2643,
        in1(1) => S2626,
        out1 => S2726
    );
nor_n_983: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2726,
        in1(1) => S2665,
        out1 => S2727
    );
nand_n_1520: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2727,
        in1(1) => S2725,
        out1 => S2728
    );
nand_n_1521: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2728,
        in1(1) => S2675,
        out1 => U1_selINC_PC
    );
nor_n_984: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2670,
        in1(1) => S2653,
        out1 => S2729
    );
nor_n_985: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2729,
        in1(1) => S2818,
        out1 => S2730
    );
nor_n_986: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2722,
        in1(1) => S2826,
        out1 => U1_INC2
    );
nor_n_987: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_INC2,
        in1(1) => S2730,
        out1 => S2731
    );
nand_n_1522: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2731,
        in1(1) => S2711,
        out1 => U1_ldPC
    );
nand_n_1523: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2662,
        in1(1) => U1_IR_out_15,
        out1 => S2732
    );
nor_n_988: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2653,
        in1(1) => S2818,
        out1 => S2733
    );
nand_n_1524: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2733,
        in1(1) => S2649,
        out1 => S2734
    );
notg_310: ENTITY WORK.notg
    PORT MAP (
        in1 => S2734,
        out1 => S2735
    );
nor_n_989: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2734,
        in1(1) => S2635,
        out1 => S2736
    );
nand_n_1525: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2735,
        in1(1) => S2634,
        out1 => S2737
    );
nor_n_990: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2666,
        in1(1) => S2627,
        out1 => S2738
    );
nand_n_1526: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2667,
        in1(1) => S2628,
        out1 => S2739
    );
nor_n_991: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2643,
        in1(1) => S2821,
        out1 => S2740
    );
notg_311: ENTITY WORK.notg
    PORT MAP (
        in1 => S2740,
        out1 => S2741
    );
nor_n_992: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2740,
        in1(1) => S2629,
        out1 => S2742
    );
nand_n_1527: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2742,
        in1(1) => S2739,
        out1 => S2743
    );
nor_n_993: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2743,
        in1(1) => S2737,
        out1 => S2744
    );
nand_n_1528: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2699,
        in1(1) => S2823,
        out1 => S2745
    );
notg_312: ENTITY WORK.notg
    PORT MAP (
        in1 => S2745,
        out1 => S2746
    );
nor_n_994: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2746,
        in1(1) => S2641,
        out1 => S2747
    );
nand_n_1529: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2747,
        in1(1) => S2744,
        out1 => S2748
    );
nand_n_1530: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2748,
        in1(1) => S2732,
        out1 => U1_ADD
    );
nand_n_1531: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2654,
        in1(1) => S2651,
        out1 => S2749
    );
nor_n_995: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2749,
        in1(1) => S2648,
        out1 => S2750
    );
nor_n_996: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2640,
        in1(1) => U1_IR_out_13,
        out1 => S2751
    );
nor_n_997: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2738,
        in1(1) => S2641,
        out1 => S2752
    );
nand_n_1532: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2739,
        in1(1) => S2638,
        out1 => S2753
    );
nand_n_1533: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2752,
        in1(1) => S2638,
        out1 => S2754
    );
nor_n_998: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2753,
        in1(1) => S2641,
        out1 => S2755
    );
nand_n_1534: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2755,
        in1(1) => S2750,
        out1 => S2756
    );
nand_n_1535: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2756,
        in1(1) => S2732,
        out1 => U1_selMO_ARU
    );
nand_n_1536: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2750,
        in1(1) => S2647,
        out1 => S2757
    );
notg_313: ENTITY WORK.notg
    PORT MAP (
        in1 => S2757,
        out1 => S2758
    );
nand_n_1537: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2758,
        in1(1) => S2739,
        out1 => S2759
    );
nand_n_1538: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2759,
        in1(1) => S2732,
        out1 => U1_selMEM_LGU
    );
nor_n_999: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2678,
        in1(1) => S2824,
        out1 => S2760
    );
notg_314: ENTITY WORK.notg
    PORT MAP (
        in1 => S2760,
        out1 => S2761
    );
nand_n_1539: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2703,
        in1(1) => U1_IR_out_1,
        out1 => S2762
    );
notg_315: ENTITY WORK.notg
    PORT MAP (
        in1 => S2762,
        out1 => S2763
    );
nor_n_1000: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2762,
        in1(1) => S2805,
        out1 => S2764
    );
nand_n_1540: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2763,
        in1(1) => U1_IR_out_0,
        out1 => S2765
    );
nor_n_1001: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2764,
        in1(1) => S2761,
        out1 => S2766
    );
nand_n_1541: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2765,
        in1(1) => S2760,
        out1 => S2767
    );
nand_n_1542: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2766,
        in1(1) => S2699,
        out1 => S2768
    );
nand_n_1543: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2733,
        in1(1) => S2638,
        out1 => S2769
    );
nor_n_1002: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2769,
        in1(1) => S2738,
        out1 => S2770
    );
nand_n_1544: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2770,
        in1(1) => S2768,
        out1 => S2771
    );
nand_n_1545: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2771,
        in1(1) => S2663,
        out1 => U1_ldAC
    );
nor_n_1003: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2754,
        in1(1) => S2734,
        out1 => S2772
    );
nand_n_1546: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2772,
        in1(1) => S2745,
        out1 => S2773
    );
nand_n_1547: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2773,
        in1(1) => S2732,
        out1 => U1_selARU_AC
    );
nor_n_1004: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2818,
        in1(1) => S2803,
        out1 => S2774
    );
nand_n_1548: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2817,
        in1(1) => U1_IR_out_12,
        out1 => S2775
    );
nand_n_1549: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2774,
        in1(1) => S2648,
        out1 => S2776
    );
nand_n_1550: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2660,
        in1(1) => S2632,
        out1 => S2777
    );
nand_n_1551: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2777,
        in1(1) => S2776,
        out1 => U1_selMEM_AC
    );
nor_n_1005: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2763,
        in1(1) => S2824,
        out1 => S2778
    );
nand_n_1552: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2729,
        in1(1) => S2817,
        out1 => S2779
    );
nor_n_1006: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2779,
        in1(1) => S2778,
        out1 => U1_ldSR_0
    );
nor_n_1007: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2683,
        in1(1) => S2826,
        out1 => U1_selSET_SR
    );
nor_n_1008: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2739,
        in1(1) => S2659,
        out1 => U1_selIN_MEM
    );
nor_n_1009: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2739,
        in1(1) => S2818,
        out1 => U1_ldIN
    );
nor_n_1010: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2627,
        in1(1) => U1_IR_out_12,
        out1 => S2780
    );
nand_n_1553: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2780,
        in1(1) => S2817,
        out1 => S2781
    );
nor_n_1011: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2781,
        in1(1) => S2751,
        out1 => U1_selMEM_IN
    );
nor_n_1012: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2775,
        in1(1) => S2712,
        out1 => U1_selINC_IN
    );
nand_n_1554: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2655,
        in1(1) => S2817,
        out1 => S2782
    );
nor_n_1013: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2708,
        in1(1) => S2805,
        out1 => S2783
    );
nand_n_1555: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2783,
        in1(1) => S2825,
        out1 => S2784
    );
nand_n_1556: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2784,
        in1(1) => S2782,
        out1 => U1_selIMM_PC
    );
nor_n_1014: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2775,
        in1(1) => S2654,
        out1 => U1_selMEM_PC
    );
nor_n_1015: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2741,
        in1(1) => S2818,
        out1 => U1_MUL
    );
nor_n_1016: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2765,
        in1(1) => S2826,
        out1 => U1_NOT
    );
nor_n_1017: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2642,
        in1(1) => S2818,
        out1 => U1_AND
    );
nor_n_1018: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2699,
        in1(1) => S2826,
        out1 => U1_sel1_ARU
    );
nor_n_1019: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2645,
        in1(1) => S2803,
        out1 => S2785
    );
nor_n_1020: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2785,
        in1(1) => S2743,
        out1 => S2786
    );
nand_n_1557: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2786,
        in1(1) => S2736,
        out1 => S2787
    );
nor_n_1021: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2787,
        in1(1) => S2760,
        out1 => U1_selIMM_LGU
    );
nor_n_1022: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2826,
        in1(1) => U1_IR_out_0,
        out1 => S2788
    );
notg_316: ENTITY WORK.notg
    PORT MAP (
        in1 => S2788,
        out1 => S2789
    );
nor_n_1023: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2789,
        in1(1) => S2762,
        out1 => U1_zeroAC
    );
nand_n_1558: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2767,
        in1(1) => S2626,
        out1 => S2790
    );
nor_n_1024: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2790,
        in1(1) => S2630,
        out1 => U1_selLGU_AC
    );
nor_n_1025: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2650,
        in1(1) => S2818,
        out1 => U1_selIMM_AC
    );
nor_n_1026: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2783,
        in1(1) => S2679,
        out1 => S2791
    );
nor_n_1027: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2791,
        in1(1) => S2826,
        out1 => U1_SE12bits
    );
nor_n_1028: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2749,
        in1(1) => S2635,
        out1 => S2792
    );
nand_n_1559: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2792,
        in1(1) => S2786,
        out1 => S2793
    );
notg_317: ENTITY WORK.notg
    PORT MAP (
        in1 => S2793,
        out1 => U1_SE4bits
    );
nor_n_1029: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2676,
        in1(1) => S2826,
        out1 => U1_selIMM_OF
    );
nand_n_1560: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2696,
        in1(1) => S2825,
        out1 => S2794
    );
nor_n_1030: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2794,
        in1(1) => S2704,
        out1 => U1_selPC_OF
    );
nor_n_1031: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => U1_selPC_OF,
        in1(1) => U1_selIMM_OF,
        out1 => S2795
    );
notg_318: ENTITY WORK.notg
    PORT MAP (
        in1 => S2795,
        out1 => U1_ldOF
    );
dff_73: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => U1_ldIR,
        NbarT => '0',
        PRE => '0',
        Q => U2_pstate,
        Si => S2832,
        global_reset => '0'
    );
dff_74: ENTITY WORK.dff
    PORT MAP (
        C => U1_clk,
        CE => '1',
        CLR => U1_rst,
        D => U2_nstate_1,
        NbarT => '0',
        PRE => '0',
        Q => S2623,
        Si => S2833,
        global_reset => '0'
    );
bufg_1: ENTITY WORK.bufg
    PORT MAP (
        in1 => U1_addrBus_0,
        out1 => addrBus(0)
    );
bufg_2: ENTITY WORK.bufg
    PORT MAP (
        in1 => U1_addrBus_1,
        out1 => addrBus(1)
    );
bufg_3: ENTITY WORK.bufg
    PORT MAP (
        in1 => U1_addrBus_10,
        out1 => addrBus(10)
    );
bufg_4: ENTITY WORK.bufg
    PORT MAP (
        in1 => U1_addrBus_11,
        out1 => addrBus(11)
    );
bufg_5: ENTITY WORK.bufg
    PORT MAP (
        in1 => U1_addrBus_12,
        out1 => addrBus(12)
    );
bufg_6: ENTITY WORK.bufg
    PORT MAP (
        in1 => U1_addrBus_13,
        out1 => addrBus(13)
    );
bufg_7: ENTITY WORK.bufg
    PORT MAP (
        in1 => U1_addrBus_14,
        out1 => addrBus(14)
    );
bufg_8: ENTITY WORK.bufg
    PORT MAP (
        in1 => U1_addrBus_15,
        out1 => addrBus(15)
    );
bufg_9: ENTITY WORK.bufg
    PORT MAP (
        in1 => U1_addrBus_2,
        out1 => addrBus(2)
    );
bufg_10: ENTITY WORK.bufg
    PORT MAP (
        in1 => U1_addrBus_3,
        out1 => addrBus(3)
    );
bufg_11: ENTITY WORK.bufg
    PORT MAP (
        in1 => U1_addrBus_4,
        out1 => addrBus(4)
    );
bufg_12: ENTITY WORK.bufg
    PORT MAP (
        in1 => U1_addrBus_5,
        out1 => addrBus(5)
    );
bufg_13: ENTITY WORK.bufg
    PORT MAP (
        in1 => U1_addrBus_6,
        out1 => addrBus(6)
    );
bufg_14: ENTITY WORK.bufg
    PORT MAP (
        in1 => U1_addrBus_7,
        out1 => addrBus(7)
    );
bufg_15: ENTITY WORK.bufg
    PORT MAP (
        in1 => U1_addrBus_8,
        out1 => addrBus(8)
    );
bufg_16: ENTITY WORK.bufg
    PORT MAP (
        in1 => U1_addrBus_9,
        out1 => addrBus(9)
    );
bufg_17: ENTITY WORK.bufg
    PORT MAP (
        in1 => clk,
        out1 => U1_clk
    );
bufg_18: ENTITY WORK.bufg
    PORT MAP (
        in1 => dataBus(0),
        out1 => U1_dataBus_0
    );
bufg_19: ENTITY WORK.bufg
    PORT MAP (
        in1 => dataBus(1),
        out1 => U1_dataBus_1
    );
bufg_20: ENTITY WORK.bufg
    PORT MAP (
        in1 => dataBus(10),
        out1 => U1_dataBus_10
    );
bufg_21: ENTITY WORK.bufg
    PORT MAP (
        in1 => dataBus(11),
        out1 => U1_dataBus_11
    );
bufg_22: ENTITY WORK.bufg
    PORT MAP (
        in1 => dataBus(12),
        out1 => U1_dataBus_12
    );
bufg_23: ENTITY WORK.bufg
    PORT MAP (
        in1 => dataBus(13),
        out1 => U1_dataBus_13
    );
bufg_24: ENTITY WORK.bufg
    PORT MAP (
        in1 => dataBus(14),
        out1 => U1_dataBus_14
    );
bufg_25: ENTITY WORK.bufg
    PORT MAP (
        in1 => dataBus(15),
        out1 => U1_dataBus_15
    );
bufg_26: ENTITY WORK.bufg
    PORT MAP (
        in1 => dataBus(2),
        out1 => U1_dataBus_2
    );
bufg_27: ENTITY WORK.bufg
    PORT MAP (
        in1 => dataBus(3),
        out1 => U1_dataBus_3
    );
bufg_28: ENTITY WORK.bufg
    PORT MAP (
        in1 => dataBus(4),
        out1 => U1_dataBus_4
    );
bufg_29: ENTITY WORK.bufg
    PORT MAP (
        in1 => dataBus(5),
        out1 => U1_dataBus_5
    );
bufg_30: ENTITY WORK.bufg
    PORT MAP (
        in1 => dataBus(6),
        out1 => U1_dataBus_6
    );
bufg_31: ENTITY WORK.bufg
    PORT MAP (
        in1 => dataBus(7),
        out1 => U1_dataBus_7
    );
bufg_32: ENTITY WORK.bufg
    PORT MAP (
        in1 => dataBus(8),
        out1 => U1_dataBus_8
    );
bufg_33: ENTITY WORK.bufg
    PORT MAP (
        in1 => dataBus(9),
        out1 => U1_dataBus_9
    );
bufg_34: ENTITY WORK.bufg
    PORT MAP (
        in1 => U1_dataBus_out_0,
        out1 => dataBus_out(0)
    );
bufg_35: ENTITY WORK.bufg
    PORT MAP (
        in1 => U1_dataBus_out_1,
        out1 => dataBus_out(1)
    );
bufg_36: ENTITY WORK.bufg
    PORT MAP (
        in1 => U1_dataBus_out_10,
        out1 => dataBus_out(10)
    );
bufg_37: ENTITY WORK.bufg
    PORT MAP (
        in1 => U1_dataBus_out_11,
        out1 => dataBus_out(11)
    );
bufg_38: ENTITY WORK.bufg
    PORT MAP (
        in1 => U1_dataBus_out_12,
        out1 => dataBus_out(12)
    );
bufg_39: ENTITY WORK.bufg
    PORT MAP (
        in1 => U1_dataBus_out_13,
        out1 => dataBus_out(13)
    );
bufg_40: ENTITY WORK.bufg
    PORT MAP (
        in1 => U1_dataBus_out_14,
        out1 => dataBus_out(14)
    );
bufg_41: ENTITY WORK.bufg
    PORT MAP (
        in1 => U1_dataBus_out_15,
        out1 => dataBus_out(15)
    );
bufg_42: ENTITY WORK.bufg
    PORT MAP (
        in1 => U1_dataBus_out_2,
        out1 => dataBus_out(2)
    );
bufg_43: ENTITY WORK.bufg
    PORT MAP (
        in1 => U1_dataBus_out_3,
        out1 => dataBus_out(3)
    );
bufg_44: ENTITY WORK.bufg
    PORT MAP (
        in1 => U1_dataBus_out_4,
        out1 => dataBus_out(4)
    );
bufg_45: ENTITY WORK.bufg
    PORT MAP (
        in1 => U1_dataBus_out_5,
        out1 => dataBus_out(5)
    );
bufg_46: ENTITY WORK.bufg
    PORT MAP (
        in1 => U1_dataBus_out_6,
        out1 => dataBus_out(6)
    );
bufg_47: ENTITY WORK.bufg
    PORT MAP (
        in1 => U1_dataBus_out_7,
        out1 => dataBus_out(7)
    );
bufg_48: ENTITY WORK.bufg
    PORT MAP (
        in1 => U1_dataBus_out_8,
        out1 => dataBus_out(8)
    );
bufg_49: ENTITY WORK.bufg
    PORT MAP (
        in1 => U1_dataBus_out_9,
        out1 => dataBus_out(9)
    );
bufg_50: ENTITY WORK.bufg
    PORT MAP (
        in1 => U2_readMEM,
        out1 => readMEM
    );
bufg_51: ENTITY WORK.bufg
    PORT MAP (
        in1 => rst,
        out1 => U1_rst
    );
bufg_52: ENTITY WORK.bufg
    PORT MAP (
        in1 => U1_seldataBus,
        out1 => writeMEM
    );

END ARCHITECTURE arch;
