module SAYAC_TOP(clk, rst, readyMEM, dataBusIn, readMEM, writeMEM, readIO, writeIO, dataBusOut, addrBus, readInst, PCout);

wire S0;
wire S1;
wire S2;
wire S3;
wire S4;
wire S5;
wire S6;
wire S7;
wire S8;
wire S9;
wire S10;
wire S11;
wire S12;
wire S13;
wire S14;
wire S15;
wire S16;
wire S17;
wire S18;
wire S19;
wire S20;
wire S21;
wire S22;
wire S23;
wire S24;
wire S25;
wire S26;
wire S27;
wire S28;
wire S29;
wire S30;
wire S31;
wire S32;
wire S33;
wire S34;
wire S35;
wire S36;
wire S37;
wire S38;
wire S39;
wire S40;
wire S41;
wire S42;
wire S43;
wire S44;
wire S45;
wire S46;
wire S47;
wire S48;
wire S49;
wire S50;
wire S51;
wire S52;
wire S53;
wire S54;
wire S55;
wire S56;
wire S57;
wire S58;
wire S59;
wire S60;
wire S61;
wire S62;
wire S63;
wire S64;
wire S65;
wire S66;
wire S67;
wire S68;
wire S69;
wire S70;
wire S71;
wire S72;
wire S73;
wire S74;
wire S75;
wire S76;
wire S77;
wire S78;
wire S79;
wire S80;
wire S81;
wire S82;
wire S83;
wire S84;
wire S85;
wire S86;
wire S87;
wire S88;
wire S89;
wire S90;
wire S91;
wire S92;
wire S93;
wire S94;
wire S95;
wire S96;
wire S97;
wire S98;
wire S99;
wire S100;
wire S101;
wire S102;
wire S103;
wire S104;
wire S105;
wire S106;
wire S107;
wire S108;
wire S109;
wire S110;
wire S111;
wire S112;
wire S113;
wire S114;
wire S115;
wire S116;
wire S117;
wire S118;
wire S119;
wire S120;
wire S121;
wire S122;
wire S123;
wire S124;
wire S125;
wire S126;
wire S127;
wire S128;
wire S129;
wire S130;
wire S131;
wire S132;
wire S133;
wire S134;
wire S135;
wire S136;
wire S137;
wire S138;
wire S139;
wire S140;
wire S141;
wire S142;
wire S143;
wire S144;
wire S145;
wire S146;
wire S147;
wire S148;
wire S149;
wire S150;
wire S151;
wire S152;
wire S153;
wire S154;
wire S155;
wire S156;
wire S157;
wire S158;
wire S159;
wire S160;
wire S161;
wire S162;
wire S163;
wire S164;
wire S165;
wire S166;
wire S167;
wire S168;
wire S169;
wire S170;
wire S171;
wire S172;
wire S173;
wire S174;
wire S175;
wire S176;
wire S177;
wire S178;
wire S179;
wire S180;
wire S181;
wire S182;
wire S183;
wire S184;
wire S185;
wire S186;
wire S187;
wire S188;
wire S189;
wire S190;
wire S191;
wire S192;
wire S193;
wire S194;
wire S195;
wire S196;
wire S197;
wire S198;
wire S199;
wire S200;
wire S201;
wire S202;
wire S203;
wire S204;
wire S205;
wire S206;
wire S207;
wire S208;
wire S209;
wire S210;
wire S211;
wire S212;
wire S213;
wire S214;
wire S215;
wire S216;
wire S217;
wire S218;
wire S219;
wire S220;
wire S221;
wire S222;
wire S223;
wire S224;
wire S225;
wire S226;
wire S227;
wire S228;
wire S229;
wire S230;
wire S231;
wire S232;
wire S233;
wire S234;
wire S235;
wire S236;
wire S237;
wire S238;
wire S239;
wire S240;
wire S241;
wire S242;
wire S243;
wire S244;
wire S245;
wire S246;
wire S247;
wire S248;
wire S249;
wire S250;
wire S251;
wire S252;
wire S253;
wire S254;
wire S255;
wire S256;
wire S257;
wire S258;
wire S259;
wire S260;
wire S261;
wire S262;
wire S263;
wire S264;
wire S265;
wire S266;
wire S267;
wire S268;
wire S269;
wire S270;
wire S271;
wire S272;
wire S273;
wire S274;
wire S275;
wire S276;
wire S277;
wire S278;
wire S279;
wire S280;
wire S281;
wire S282;
wire S283;
wire S284;
wire S285;
wire S286;
wire S287;
wire S288;
wire S289;
wire S290;
wire S291;
wire S292;
wire S293;
wire S294;
wire S295;
wire S296;
wire S297;
wire S298;
wire S299;
wire S300;
wire S301;
wire S302;
wire S303;
wire S304;
wire S305;
wire S306;
wire S307;
wire S308;
wire S309;
wire S310;
wire S311;
wire S312;
wire S313;
wire S314;
wire S315;
wire S316;
wire S317;
wire S318;
wire S319;
wire S320;
wire S321;
wire S322;
wire S323;
wire S324;
wire S325;
wire S326;
wire S327;
wire S328;
wire S329;
wire S330;
wire S331;
wire S332;
wire S333;
wire S334;
wire S335;
wire S336;
wire S337;
wire S338;
wire S339;
wire S340;
wire S341;
wire S342;
wire S343;
wire S344;
wire S345;
wire S346;
wire S347;
wire S348;
wire S349;
wire S350;
wire S351;
wire S352;
wire S353;
wire S354;
wire S355;
wire S356;
wire S357;
wire S358;
wire S359;
wire S360;
wire S361;
wire S362;
wire S363;
wire S364;
wire S365;
wire S366;
wire S367;
wire S368;
wire S369;
wire S370;
wire S371;
wire S372;
wire S373;
wire S374;
wire S375;
wire S376;
wire S377;
wire S378;
wire S379;
wire S380;
wire S381;
wire S382;
wire S383;
wire S384;
wire S385;
wire S386;
wire S387;
wire S388;
wire S389;
wire S390;
wire S391;
wire S392;
wire S393;
wire S394;
wire S395;
wire S396;
wire S397;
wire S398;
wire S399;
wire S400;
wire S401;
wire S402;
wire S403;
wire S404;
wire S405;
wire S406;
wire S407;
wire S408;
wire S409;
wire S410;
wire S411;
wire S412;
wire S413;
wire S414;
wire S415;
wire S416;
wire S417;
wire S418;
wire S419;
wire S420;
wire S421;
wire S422;
wire S423;
wire S424;
wire S425;
wire S426;
wire S427;
wire S428;
wire S429;
wire S430;
wire S431;
wire S432;
wire S433;
wire S434;
wire S435;
wire S436;
wire S437;
wire S438;
wire S439;
wire S440;
wire S441;
wire S442;
wire S443;
wire S444;
wire S445;
wire S446;
wire S447;
wire S448;
wire S449;
wire S450;
wire S451;
wire S452;
wire S453;
wire S454;
wire S455;
wire S456;
wire S457;
wire S458;
wire S459;
wire S460;
wire S461;
wire S462;
wire S463;
wire S464;
wire S465;
wire S466;
wire S467;
wire S468;
wire S469;
wire S470;
wire S471;
wire S472;
wire S473;
wire S474;
wire S475;
wire S476;
wire S477;
wire S478;
wire S479;
wire S480;
wire S481;
wire S482;
wire S483;
wire S484;
wire S485;
wire S486;
wire S487;
wire S488;
wire S489;
wire S490;
wire S491;
wire S492;
wire S493;
wire S494;
wire S495;
wire S496;
wire S497;
wire S498;
wire S499;
wire S500;
wire S501;
wire S502;
wire S503;
wire S504;
wire S505;
wire S506;
wire S507;
wire S508;
wire S509;
wire S510;
wire S511;
wire S512;
wire S513;
wire S514;
wire S515;
wire S516;
wire S517;
wire S518;
wire S519;
wire S520;
wire S521;
wire S522;
wire S523;
wire S524;
wire S525;
wire S526;
wire S527;
wire S528;
wire S529;
wire S530;
wire S531;
wire S532;
wire S533;
wire S534;
wire S535;
wire S536;
wire S537;
wire S538;
wire S539;
wire S540;
wire S541;
wire S542;
wire S543;
wire S544;
wire S545;
wire S546;
wire S547;
wire S548;
wire S549;
wire S550;
wire S551;
wire S552;
wire S553;
wire S554;
wire S555;
wire S556;
wire S557;
wire S558;
wire S559;
wire S560;
wire S561;
wire S562;
wire S563;
wire S564;
wire S565;
wire S566;
wire S567;
wire S568;
wire S569;
wire S570;
wire S571;
wire S572;
wire S573;
wire S574;
wire S575;
wire S576;
wire S577;
wire S578;
wire S579;
wire S580;
wire S581;
wire S582;
wire S583;
wire S584;
wire S585;
wire S586;
wire S587;
wire S588;
wire S589;
wire S590;
wire S591;
wire S592;
wire S593;
wire S594;
wire S595;
wire S596;
wire S597;
wire S598;
wire S599;
wire S600;
wire S601;
wire S602;
wire S603;
wire S604;
wire S605;
wire S606;
wire S607;
wire S608;
wire S609;
wire S610;
wire S611;
wire S612;
wire S613;
wire S614;
wire S615;
wire S616;
wire S617;
wire S618;
wire S619;
wire S620;
wire S621;
wire S622;
wire S623;
wire S624;
wire S625;
wire S626;
wire S627;
wire S628;
wire S629;
wire S630;
wire S631;
wire S632;
wire S633;
wire S634;
wire S635;
wire S636;
wire S637;
wire S638;
wire S639;
wire S640;
wire S641;
wire S642;
wire S643;
wire S644;
wire S645;
wire S646;
wire S647;
wire S648;
wire S649;
wire S650;
wire S651;
wire S652;
wire S653;
wire S654;
wire S655;
wire S656;
wire S657;
wire S658;
wire S659;
wire S660;
wire S661;
wire S662;
wire S663;
wire S664;
wire S665;
wire S666;
wire S667;
wire S668;
wire S669;
wire S670;
wire S671;
wire S672;
wire S673;
wire S674;
wire S675;
wire S676;
wire S677;
wire S678;
wire S679;
wire S680;
wire S681;
wire S682;
wire S683;
wire S684;
wire S685;
wire S686;
wire S687;
wire S688;
wire S689;
wire S690;
wire S691;
wire S692;
wire S693;
wire S694;
wire S695;
wire S696;
wire S697;
wire S698;
wire S699;
wire S700;
wire S701;
wire S702;
wire S703;
wire S704;
wire S705;
wire S706;
wire S707;
wire S708;
wire S709;
wire S710;
wire S711;
wire S712;
wire S713;
wire S714;
wire S715;
wire S716;
wire S717;
wire S718;
wire S719;
wire S720;
wire S721;
wire S722;
wire S723;
wire S724;
wire S725;
wire S726;
wire S727;
wire S728;
wire S729;
wire S730;
wire S731;
wire S732;
wire S733;
wire S734;
wire S735;
wire S736;
wire S737;
wire S738;
wire S739;
wire S740;
wire S741;
wire S742;
wire S743;
wire S744;
wire S745;
wire S746;
wire S747;
wire S748;
wire S749;
wire S750;
wire S751;
wire S752;
wire S753;
wire S754;
wire S755;
wire S756;
wire S757;
wire S758;
wire S759;
wire S760;
wire S761;
wire S762;
wire S763;
wire S764;
wire S765;
wire S766;
wire S767;
wire S768;
wire S769;
wire S770;
wire S771;
wire S772;
wire S773;
wire S774;
wire S775;
wire S776;
wire S777;
wire S778;
wire S779;
wire S780;
wire S781;
wire S782;
wire S783;
wire S784;
wire S785;
wire S786;
wire S787;
wire S788;
wire S789;
wire S790;
wire S791;
wire S792;
wire S793;
wire S794;
wire S795;
wire S796;
wire S797;
wire S798;
wire S799;
wire S800;
wire S801;
wire S802;
wire S803;
wire S804;
wire S805;
wire S806;
wire S807;
wire S808;
wire S809;
wire S810;
wire S811;
wire S812;
wire S813;
wire S814;
wire S815;
wire S816;
wire S817;
wire S818;
wire S819;
wire S820;
wire S821;
wire S822;
wire S823;
wire S824;
wire S825;
wire S826;
wire S827;
wire S828;
wire S829;
wire S830;
wire S831;
wire S832;
wire S833;
wire S834;
wire S835;
wire S836;
wire S837;
wire S838;
wire S839;
wire S840;
wire S841;
wire S842;
wire S843;
wire S844;
wire S845;
wire S846;
wire S847;
wire S848;
wire S849;
wire S850;
wire S851;
wire S852;
wire S853;
wire S854;
wire S855;
wire S856;
wire S857;
wire S858;
wire S859;
wire S860;
wire S861;
wire S862;
wire S863;
wire S864;
wire S865;
wire S866;
wire S867;
wire S868;
wire S869;
wire S870;
wire S871;
wire S872;
wire S873;
wire S874;
wire S875;
wire S876;
wire S877;
wire S878;
wire S879;
wire S880;
wire S881;
wire S882;
wire S883;
wire S884;
wire S885;
wire S886;
wire S887;
wire S888;
wire S889;
wire S890;
wire S891;
wire S892;
wire S893;
wire S894;
wire S895;
wire S896;
wire S897;
wire S898;
wire S899;
wire S900;
wire S901;
wire S902;
wire S903;
wire S904;
wire S905;
wire S906;
wire S907;
wire S908;
wire S909;
wire S910;
wire S911;
wire S912;
wire S913;
wire S914;
wire S915;
wire S916;
wire S917;
wire S918;
wire S919;
wire S920;
wire S921;
wire S922;
wire S923;
wire S924;
wire S925;
wire S926;
wire S927;
wire S928;
wire S929;
wire S930;
wire S931;
wire S932;
wire S933;
wire S934;
wire S935;
wire S936;
wire S937;
wire S938;
wire S939;
wire S940;
wire S941;
wire S942;
wire S943;
wire S944;
wire S945;
wire S946;
wire S947;
wire S948;
wire S949;
wire S950;
wire S951;
wire S952;
wire S953;
wire S954;
wire S955;
wire S956;
wire S957;
wire S958;
wire S959;
wire S960;
wire S961;
wire S962;
wire S963;
wire S964;
wire S965;
wire S966;
wire S967;
wire S968;
wire S969;
wire S970;
wire S971;
wire S972;
wire S973;
wire S974;
wire S975;
wire S976;
wire S977;
wire S978;
wire S979;
wire S980;
wire S981;
wire S982;
wire S983;
wire S984;
wire S985;
wire S986;
wire S987;
wire S988;
wire S989;
wire S990;
wire S991;
wire S992;
wire S993;
wire S994;
wire S995;
wire S996;
wire S997;
wire S998;
wire S999;
wire S1000;
wire S1001;
wire S1002;
wire S1003;
wire S1004;
wire S1005;
wire S1006;
wire S1007;
wire S1008;
wire S1009;
wire S1010;
wire S1011;
wire S1012;
wire S1013;
wire S1014;
wire S1015;
wire S1016;
wire S1017;
wire S1018;
wire S1019;
wire S1020;
wire S1021;
wire S1022;
wire S1023;
wire S1024;
wire S1025;
wire S1026;
wire S1027;
wire S1028;
wire S1029;
wire S1030;
wire S1031;
wire S1032;
wire S1033;
wire S1034;
wire S1035;
wire S1036;
wire S1037;
wire S1038;
wire S1039;
wire S1040;
wire S1041;
wire S1042;
wire S1043;
wire S1044;
wire S1045;
wire S1046;
wire S1047;
wire S1048;
wire S1049;
wire S1050;
wire S1051;
wire S1052;
wire S1053;
wire S1054;
wire S1055;
wire S1056;
wire S1057;
wire S1058;
wire S1059;
wire S1060;
wire S1061;
wire S1062;
wire S1063;
wire S1064;
wire S1065;
wire S1066;
wire S1067;
wire S1068;
wire S1069;
wire S1070;
wire S1071;
wire S1072;
wire S1073;
wire S1074;
wire S1075;
wire S1076;
wire S1077;
wire S1078;
wire S1079;
wire S1080;
wire S1081;
wire S1082;
wire S1083;
wire S1084;
wire S1085;
wire S1086;
wire S1087;
wire S1088;
wire S1089;
wire S1090;
wire S1091;
wire S1092;
wire S1093;
wire S1094;
wire S1095;
wire S1096;
wire S1097;
wire S1098;
wire S1099;
wire S1100;
wire S1101;
wire S1102;
wire S1103;
wire S1104;
wire S1105;
wire S1106;
wire S1107;
wire S1108;
wire S1109;
wire S1110;
wire S1111;
wire S1112;
wire S1113;
wire S1114;
wire S1115;
wire S1116;
wire S1117;
wire S1118;
wire S1119;
wire S1120;
wire S1121;
wire S1122;
wire S1123;
wire S1124;
wire S1125;
wire S1126;
wire S1127;
wire S1128;
wire S1129;
wire S1130;
wire S1131;
wire S1132;
wire S1133;
wire S1134;
wire S1135;
wire S1136;
wire S1137;
wire S1138;
wire S1139;
wire S1140;
wire S1141;
wire S1142;
wire S1143;
wire S1144;
wire S1145;
wire S1146;
wire S1147;
wire S1148;
wire S1149;
wire S1150;
wire S1151;
wire S1152;
wire S1153;
wire S1154;
wire S1155;
wire S1156;
wire S1157;
wire S1158;
wire S1159;
wire S1160;
wire S1161;
wire S1162;
wire S1163;
wire S1164;
wire S1165;
wire S1166;
wire S1167;
wire S1168;
wire S1169;
wire S1170;
wire S1171;
wire S1172;
wire S1173;
wire S1174;
wire S1175;
wire S1176;
wire S1177;
wire S1178;
wire S1179;
wire S1180;
wire S1181;
wire S1182;
wire S1183;
wire S1184;
wire S1185;
wire S1186;
wire S1187;
wire S1188;
wire S1189;
wire S1190;
wire S1191;
wire S1192;
wire S1193;
wire S1194;
wire S1195;
wire S1196;
wire S1197;
wire S1198;
wire S1199;
wire S1200;
wire S1201;
wire S1202;
wire S1203;
wire S1204;
wire S1205;
wire S1206;
wire S1207;
wire S1208;
wire S1209;
wire S1210;
wire S1211;
wire S1212;
wire S1213;
wire S1214;
wire S1215;
wire S1216;
wire S1217;
wire S1218;
wire S1219;
wire S1220;
wire S1221;
wire S1222;
wire S1223;
wire S1224;
wire S1225;
wire S1226;
wire S1227;
wire S1228;
wire S1229;
wire S1230;
wire S1231;
wire S1232;
wire S1233;
wire S1234;
wire S1235;
wire S1236;
wire S1237;
wire S1238;
wire S1239;
wire S1240;
wire S1241;
wire S1242;
wire S1243;
wire S1244;
wire S1245;
wire S1246;
wire S1247;
wire S1248;
wire S1249;
wire S1250;
wire S1251;
wire S1252;
wire S1253;
wire S1254;
wire S1255;
wire S1256;
wire S1257;
wire S1258;
wire S1259;
wire S1260;
wire S1261;
wire S1262;
wire S1263;
wire S1264;
wire S1265;
wire S1266;
wire S1267;
wire S1268;
wire S1269;
wire S1270;
wire S1271;
wire S1272;
wire S1273;
wire S1274;
wire S1275;
wire S1276;
wire S1277;
wire S1278;
wire S1279;
wire S1280;
wire S1281;
wire S1282;
wire S1283;
wire S1284;
wire S1285;
wire S1286;
wire S1287;
wire S1288;
wire S1289;
wire S1290;
wire S1291;
wire S1292;
wire S1293;
wire S1294;
wire S1295;
wire S1296;
wire S1297;
wire S1298;
wire S1299;
wire S1300;
wire S1301;
wire S1302;
wire S1303;
wire S1304;
wire S1305;
wire S1306;
wire S1307;
wire S1308;
wire S1309;
wire S1310;
wire S1311;
wire S1312;
wire S1313;
wire S1314;
wire S1315;
wire S1316;
wire S1317;
wire S1318;
wire S1319;
wire S1320;
wire S1321;
wire S1322;
wire S1323;
wire S1324;
wire S1325;
wire S1326;
wire S1327;
wire S1328;
wire S1329;
wire S1330;
wire S1331;
wire S1332;
wire S1333;
wire S1334;
wire S1335;
wire S1336;
wire S1337;
wire S1338;
wire S1339;
wire S1340;
wire S1341;
wire S1342;
wire S1343;
wire S1344;
wire S1345;
wire S1346;
wire S1347;
wire S1348;
wire S1349;
wire S1350;
wire S1351;
wire S1352;
wire S1353;
wire S1354;
wire S1355;
wire S1356;
wire S1357;
wire S1358;
wire S1359;
wire S1360;
wire S1361;
wire S1362;
wire S1363;
wire S1364;
wire S1365;
wire S1366;
wire S1367;
wire S1368;
wire S1369;
wire S1370;
wire S1371;
wire S1372;
wire S1373;
wire S1374;
wire S1375;
wire S1376;
wire S1377;
wire S1378;
wire S1379;
wire S1380;
wire S1381;
wire S1382;
wire S1383;
wire S1384;
wire S1385;
wire S1386;
wire S1387;
wire S1388;
wire S1389;
wire S1390;
wire S1391;
wire S1392;
wire S1393;
wire S1394;
wire S1395;
wire S1396;
wire S1397;
wire S1398;
wire S1399;
wire S1400;
wire S1401;
wire S1402;
wire S1403;
wire S1404;
wire S1405;
wire S1406;
wire S1407;
wire S1408;
wire S1409;
wire S1410;
wire S1411;
wire S1412;
wire S1413;
wire S1414;
wire S1415;
wire S1416;
wire S1417;
wire S1418;
wire S1419;
wire S1420;
wire S1421;
wire S1422;
wire S1423;
wire S1424;
wire S1425;
wire S1426;
wire S1427;
wire S1428;
wire S1429;
wire S1430;
wire S1431;
wire S1432;
wire S1433;
wire S1434;
wire S1435;
wire S1436;
wire S1437;
wire S1438;
wire S1439;
wire S1440;
wire S1441;
wire S1442;
wire S1443;
wire S1444;
wire S1445;
wire S1446;
wire S1447;
wire S1448;
wire S1449;
wire S1450;
wire S1451;
wire S1452;
wire S1453;
wire S1454;
wire S1455;
wire S1456;
wire S1457;
wire S1458;
wire S1459;
wire S1460;
wire S1461;
wire S1462;
wire S1463;
wire S1464;
wire S1465;
wire S1466;
wire S1467;
wire S1468;
wire S1469;
wire S1470;
wire S1471;
wire S1472;
wire S1473;
wire S1474;
wire S1475;
wire S1476;
wire S1477;
wire S1478;
wire S1479;
wire S1480;
wire S1481;
wire S1482;
wire S1483;
wire S1484;
wire S1485;
wire S1486;
wire S1487;
wire S1488;
wire S1489;
wire S1490;
wire S1491;
wire S1492;
wire S1493;
wire S1494;
wire S1495;
wire S1496;
wire S1497;
wire S1498;
wire S1499;
wire S1500;
wire S1501;
wire S1502;
wire S1503;
wire S1504;
wire S1505;
wire S1506;
wire S1507;
wire S1508;
wire S1509;
wire S1510;
wire S1511;
wire S1512;
wire S1513;
wire S1514;
wire S1515;
wire S1516;
wire S1517;
wire S1518;
wire S1519;
wire S1520;
wire S1521;
wire S1522;
wire S1523;
wire S1524;
wire S1525;
wire S1526;
wire S1527;
wire S1528;
wire S1529;
wire S1530;
wire S1531;
wire S1532;
wire S1533;
wire S1534;
wire S1535;
wire S1536;
wire S1537;
wire S1538;
wire S1539;
wire S1540;
wire S1541;
wire S1542;
wire S1543;
wire S1544;
wire S1545;
wire S1546;
wire S1547;
wire S1548;
wire S1549;
wire S1550;
wire S1551;
wire S1552;
wire S1553;
wire S1554;
wire S1555;
wire S1556;
wire S1557;
wire S1558;
wire S1559;
wire S1560;
wire S1561;
wire S1562;
wire S1563;
wire S1564;
wire S1565;
wire S1566;
wire S1567;
wire S1568;
wire S1569;
wire S1570;
wire S1571;
wire S1572;
wire S1573;
wire S1574;
wire S1575;
wire S1576;
wire S1577;
wire S1578;
wire S1579;
wire S1580;
wire S1581;
wire S1582;
wire S1583;
wire S1584;
wire S1585;
wire S1586;
wire S1587;
wire S1588;
wire S1589;
wire S1590;
wire S1591;
wire S1592;
wire S1593;
wire S1594;
wire S1595;
wire S1596;
wire S1597;
wire S1598;
wire S1599;
wire S1600;
wire S1601;
wire S1602;
wire S1603;
wire S1604;
wire S1605;
wire S1606;
wire S1607;
wire S1608;
wire S1609;
wire S1610;
wire S1611;
wire S1612;
wire S1613;
wire S1614;
wire S1615;
wire S1616;
wire S1617;
wire S1618;
wire S1619;
wire S1620;
wire S1621;
wire S1622;
wire S1623;
wire S1624;
wire S1625;
wire S1626;
wire S1627;
wire S1628;
wire S1629;
wire S1630;
wire S1631;
wire S1632;
wire S1633;
wire S1634;
wire S1635;
wire S1636;
wire S1637;
wire S1638;
wire S1639;
wire S1640;
wire S1641;
wire S1642;
wire S1643;
wire S1644;
wire S1645;
wire S1646;
wire S1647;
wire S1648;
wire S1649;
wire S1650;
wire S1651;
wire S1652;
wire S1653;
wire S1654;
wire S1655;
wire S1656;
wire S1657;
wire S1658;
wire S1659;
wire S1660;
wire S1661;
wire S1662;
wire S1663;
wire S1664;
wire S1665;
wire S1666;
wire S1667;
wire S1668;
wire S1669;
wire S1670;
wire S1671;
wire S1672;
wire S1673;
wire S1674;
wire S1675;
wire S1676;
wire S1677;
wire S1678;
wire S1679;
wire S1680;
wire S1681;
wire S1682;
wire S1683;
wire S1684;
wire S1685;
wire S1686;
wire S1687;
wire S1688;
wire S1689;
wire S1690;
wire S1691;
wire S1692;
wire S1693;
wire S1694;
wire S1695;
wire S1696;
wire S1697;
wire S1698;
wire S1699;
wire S1700;
wire S1701;
wire S1702;
wire S1703;
wire S1704;
wire S1705;
wire S1706;
wire S1707;
wire S1708;
wire S1709;
wire S1710;
wire S1711;
wire S1712;
wire S1713;
wire S1714;
wire S1715;
wire S1716;
wire S1717;
wire S1718;
wire S1719;
wire S1720;
wire S1721;
wire S1722;
wire S1723;
wire S1724;
wire S1725;
wire S1726;
wire S1727;
wire S1728;
wire S1729;
wire S1730;
wire S1731;
wire S1732;
wire S1733;
wire S1734;
wire S1735;
wire S1736;
wire S1737;
wire S1738;
wire S1739;
wire S1740;
wire S1741;
wire S1742;
wire S1743;
wire S1744;
wire S1745;
wire S1746;
wire S1747;
wire S1748;
wire S1749;
wire S1750;
wire S1751;
wire S1752;
wire S1753;
wire S1754;
wire S1755;
wire S1756;
wire S1757;
wire S1758;
wire S1759;
wire S1760;
wire S1761;
wire S1762;
wire S1763;
wire S1764;
wire S1765;
wire S1766;
wire S1767;
wire S1768;
wire S1769;
wire S1770;
wire S1771;
wire S1772;
wire S1773;
wire S1774;
wire S1775;
wire S1776;
wire S1777;
wire S1778;
wire S1779;
wire S1780;
wire S1781;
wire S1782;
wire S1783;
wire S1784;
wire S1785;
wire S1786;
wire S1787;
wire S1788;
wire S1789;
wire S1790;
wire S1791;
wire S1792;
wire S1793;
wire S1794;
wire S1795;
wire S1796;
wire S1797;
wire S1798;
wire S1799;
wire S1800;
wire S1801;
wire S1802;
wire S1803;
wire S1804;
wire S1805;
wire S1806;
wire S1807;
wire S1808;
wire S1809;
wire S1810;
wire S1811;
wire S1812;
wire S1813;
wire S1814;
wire S1815;
wire S1816;
wire S1817;
wire S1818;
wire S1819;
wire S1820;
wire S1821;
wire S1822;
wire S1823;
wire S1824;
wire S1825;
wire S1826;
wire S1827;
wire S1828;
wire S1829;
wire S1830;
wire S1831;
wire S1832;
wire S1833;
wire S1834;
wire S1835;
wire S1836;
wire S1837;
wire S1838;
wire S1839;
wire S1840;
wire S1841;
wire S1842;
wire S1843;
wire S1844;
wire S1845;
wire S1846;
wire S1847;
wire S1848;
wire S1849;
wire S1850;
wire S1851;
wire S1852;
wire S1853;
wire S1854;
wire S1855;
wire S1856;
wire S1857;
wire S1858;
wire S1859;
wire S1860;
wire S1861;
wire S1862;
wire S1863;
wire S1864;
wire S1865;
wire S1866;
wire S1867;
wire S1868;
wire S1869;
wire S1870;
wire S1871;
wire S1872;
wire S1873;
wire S1874;
wire S1875;
wire S1876;
wire S1877;
wire S1878;
wire S1879;
wire S1880;
wire S1881;
wire S1882;
wire S1883;
wire S1884;
wire S1885;
wire S1886;
wire S1887;
wire S1888;
wire S1889;
wire S1890;
wire S1891;
wire S1892;
wire S1893;
wire S1894;
wire S1895;
wire S1896;
wire S1897;
wire S1898;
wire S1899;
wire S1900;
wire S1901;
wire S1902;
wire S1903;
wire S1904;
wire S1905;
wire S1906;
wire S1907;
wire S1908;
wire S1909;
wire S1910;
wire S1911;
wire S1912;
wire S1913;
wire S1914;
wire S1915;
wire S1916;
wire S1917;
wire S1918;
wire S1919;
wire S1920;
wire S1921;
wire S1922;
wire S1923;
wire S1924;
wire S1925;
wire S1926;
wire S1927;
wire S1928;
wire S1929;
wire S1930;
wire S1931;
wire S1932;
wire S1933;
wire S1934;
wire S1935;
wire S1936;
wire S1937;
wire S1938;
wire S1939;
wire S1940;
wire S1941;
wire S1942;
wire S1943;
wire S1944;
wire S1945;
wire S1946;
wire S1947;
wire S1948;
wire S1949;
wire S1950;
wire S1951;
wire S1952;
wire S1953;
wire S1954;
wire S1955;
wire S1956;
wire S1957;
wire S1958;
wire S1959;
wire S1960;
wire S1961;
wire S1962;
wire S1963;
wire S1964;
wire S1965;
wire S1966;
wire S1967;
wire S1968;
wire S1969;
wire S1970;
wire S1971;
wire S1972;
wire S1973;
wire S1974;
wire S1975;
wire S1976;
wire S1977;
wire S1978;
wire S1979;
wire S1980;
wire S1981;
wire S1982;
wire S1983;
wire S1984;
wire S1985;
wire S1986;
wire S1987;
wire S1988;
wire S1989;
wire S1990;
wire S1991;
wire S1992;
wire S1993;
wire S1994;
wire S1995;
wire S1996;
wire S1997;
wire S1998;
wire S1999;
wire S2000;
wire S2001;
wire S2002;
wire S2003;
wire S2004;
wire S2005;
wire S2006;
wire S2007;
wire S2008;
wire S2009;
wire S2010;
wire S2011;
wire S2012;
wire S2013;
wire S2014;
wire S2015;
wire S2016;
wire S2017;
wire S2018;
wire S2019;
wire S2020;
wire S2021;
wire S2022;
wire S2023;
wire S2024;
wire S2025;
wire S2026;
wire S2027;
wire S2028;
wire S2029;
wire S2030;
wire S2031;
wire S2032;
wire S2033;
wire S2034;
wire S2035;
wire S2036;
wire S2037;
wire S2038;
wire S2039;
wire S2040;
wire S2041;
wire S2042;
wire S2043;
wire S2044;
wire S2045;
wire S2046;
wire S2047;
wire S2048;
wire S2049;
wire S2050;
wire S2051;
wire S2052;
wire S2053;
wire S2054;
wire S2055;
wire S2056;
wire S2057;
wire S2058;
wire S2059;
wire S2060;
wire S2061;
wire S2062;
wire S2063;
wire S2064;
wire S2065;
wire S2066;
wire S2067;
wire S2068;
wire S2069;
wire S2070;
wire S2071;
wire S2072;
wire S2073;
wire S2074;
wire S2075;
wire S2076;
wire S2077;
wire S2078;
wire S2079;
wire S2080;
wire S2081;
wire S2082;
wire S2083;
wire S2084;
wire S2085;
wire S2086;
wire S2087;
wire S2088;
wire S2089;
wire S2090;
wire S2091;
wire S2092;
wire S2093;
wire S2094;
wire S2095;
wire S2096;
wire S2097;
wire S2098;
wire S2099;
wire S2100;
wire S2101;
wire S2102;
wire S2103;
wire S2104;
wire S2105;
wire S2106;
wire S2107;
wire S2108;
wire S2109;
wire S2110;
wire S2111;
wire S2112;
wire S2113;
wire S2114;
wire S2115;
wire S2116;
wire S2117;
wire S2118;
wire S2119;
wire S2120;
wire S2121;
wire S2122;
wire S2123;
wire S2124;
wire S2125;
wire S2126;
wire S2127;
wire S2128;
wire S2129;
wire S2130;
wire S2131;
wire S2132;
wire S2133;
wire S2134;
wire S2135;
wire S2136;
wire S2137;
wire S2138;
wire S2139;
wire S2140;
wire S2141;
wire S2142;
wire S2143;
wire S2144;
wire S2145;
wire S2146;
wire S2147;
wire S2148;
wire S2149;
wire S2150;
wire S2151;
wire S2152;
wire S2153;
wire S2154;
wire S2155;
wire S2156;
wire S2157;
wire S2158;
wire S2159;
wire S2160;
wire S2161;
wire S2162;
wire S2163;
wire S2164;
wire S2165;
wire S2166;
wire S2167;
wire S2168;
wire S2169;
wire S2170;
wire S2171;
wire S2172;
wire S2173;
wire S2174;
wire S2175;
wire S2176;
wire S2177;
wire S2178;
wire S2179;
wire S2180;
wire S2181;
wire S2182;
wire S2183;
wire S2184;
wire S2185;
wire S2186;
wire S2187;
wire S2188;
wire S2189;
wire S2190;
wire S2191;
wire S2192;
wire S2193;
wire S2194;
wire S2195;
wire S2196;
wire S2197;
wire S2198;
wire S2199;
wire S2200;
wire S2201;
wire S2202;
wire S2203;
wire S2204;
wire S2205;
wire S2206;
wire S2207;
wire S2208;
wire S2209;
wire S2210;
wire S2211;
wire S2212;
wire S2213;
wire S2214;
wire S2215;
wire S2216;
wire S2217;
wire S2218;
wire S2219;
wire S2220;
wire S2221;
wire S2222;
wire S2223;
wire S2224;
wire S2225;
wire S2226;
wire S2227;
wire S2228;
wire S2229;
wire S2230;
wire S2231;
wire S2232;
wire S2233;
wire S2234;
wire S2235;
wire S2236;
wire S2237;
wire S2238;
wire S2239;
wire S2240;
wire S2241;
wire S2242;
wire S2243;
wire S2244;
wire S2245;
wire S2246;
wire S2247;
wire S2248;
wire S2249;
wire S2250;
wire S2251;
wire S2252;
wire S2253;
wire S2254;
wire S2255;
wire S2256;
wire S2257;
wire S2258;
wire S2259;
wire S2260;
wire S2261;
wire S2262;
wire S2263;
wire S2264;
wire S2265;
wire S2266;
wire S2267;
wire S2268;
wire S2269;
wire S2270;
wire S2271;
wire S2272;
wire S2273;
wire S2274;
wire S2275;
wire S2276;
wire S2277;
wire S2278;
wire S2279;
wire S2280;
wire S2281;
wire S2282;
wire S2283;
wire S2284;
wire S2285;
wire S2286;
wire S2287;
wire S2288;
wire S2289;
wire S2290;
wire S2291;
wire S2292;
wire S2293;
wire S2294;
wire S2295;
wire S2296;
wire S2297;
wire S2298;
wire S2299;
wire S2300;
wire S2301;
wire S2302;
wire S2303;
wire S2304;
wire S2305;
wire S2306;
wire S2307;
wire S2308;
wire S2309;
wire S2310;
wire S2311;
wire S2312;
wire S2313;
wire S2314;
wire S2315;
wire S2316;
wire S2317;
wire S2318;
wire S2319;
wire S2320;
wire S2321;
wire S2322;
wire S2323;
wire S2324;
wire S2325;
wire S2326;
wire S2327;
wire S2328;
wire S2329;
wire S2330;
wire S2331;
wire S2332;
wire S2333;
wire S2334;
wire S2335;
wire S2336;
wire S2337;
wire S2338;
wire S2339;
wire S2340;
wire S2341;
wire S2342;
wire S2343;
wire S2344;
wire S2345;
wire S2346;
wire S2347;
wire S2348;
wire S2349;
wire S2350;
wire S2351;
wire S2352;
wire S2353;
wire S2354;
wire S2355;
wire S2356;
wire S2357;
wire S2358;
wire S2359;
wire S2360;
wire S2361;
wire S2362;
wire S2363;
wire S2364;
wire S2365;
wire S2366;
wire S2367;
wire S2368;
wire S2369;
wire S2370;
wire S2371;
wire S2372;
wire S2373;
wire S2374;
wire S2375;
wire S2376;
wire S2377;
wire S2378;
wire S2379;
wire S2380;
wire S2381;
wire S2382;
wire S2383;
wire S2384;
wire S2385;
wire S2386;
wire S2387;
wire S2388;
wire S2389;
wire S2390;
wire S2391;
wire S2392;
wire S2393;
wire S2394;
wire S2395;
wire S2396;
wire S2397;
wire S2398;
wire S2399;
wire S2400;
wire S2401;
wire S2402;
wire S2403;
wire S2404;
wire S2405;
wire S2406;
wire S2407;
wire S2408;
wire S2409;
wire S2410;
wire S2411;
wire S2412;
wire S2413;
wire S2414;
wire S2415;
wire S2416;
wire S2417;
wire S2418;
wire S2419;
wire S2420;
wire S2421;
wire S2422;
wire S2423;
wire S2424;
wire S2425;
wire S2426;
wire S2427;
wire S2428;
wire S2429;
wire S2430;
wire S2431;
wire S2432;
wire S2433;
wire S2434;
wire S2435;
wire S2436;
wire S2437;
wire S2438;
wire S2439;
wire S2440;
wire S2441;
wire S2442;
wire S2443;
wire S2444;
wire S2445;
wire S2446;
wire S2447;
wire S2448;
wire S2449;
wire S2450;
wire S2451;
wire S2452;
wire S2453;
wire S2454;
wire S2455;
wire S2456;
wire S2457;
wire S2458;
wire S2459;
wire S2460;
wire S2461;
wire S2462;
wire S2463;
wire S2464;
wire S2465;
wire S2466;
wire S2467;
wire S2468;
wire S2469;
wire S2470;
wire S2471;
wire S2472;
wire S2473;
wire S2474;
wire S2475;
wire S2476;
wire S2477;
wire S2478;
wire S2479;
wire S2480;
wire S2481;
wire S2482;
wire S2483;
wire S2484;
wire S2485;
wire S2486;
wire S2487;
wire S2488;
wire S2489;
wire S2490;
wire S2491;
wire S2492;
wire S2493;
wire S2494;
wire S2495;
wire S2496;
wire S2497;
wire S2498;
wire S2499;
wire S2500;
wire S2501;
wire S2502;
wire S2503;
wire S2504;
wire S2505;
wire S2506;
wire S2507;
wire S2508;
wire S2509;
wire S2510;
wire S2511;
wire S2512;
wire S2513;
wire S2514;
wire S2515;
wire S2516;
wire S2517;
wire S2518;
wire S2519;
wire S2520;
wire S2521;
wire S2522;
wire S2523;
wire S2524;
wire S2525;
wire S2526;
wire S2527;
wire S2528;
wire S2529;
wire S2530;
wire S2531;
wire S2532;
wire S2533;
wire S2534;
wire S2535;
wire S2536;
wire S2537;
wire S2538;
wire S2539;
wire S2540;
wire S2541;
wire S2542;
wire S2543;
wire S2544;
wire S2545;
wire S2546;
wire S2547;
wire S2548;
wire S2549;
wire S2550;
wire S2551;
wire S2552;
wire S2553;
wire S2554;
wire S2555;
wire S2556;
wire S2557;
wire S2558;
wire S2559;
wire S2560;
wire S2561;
wire S2562;
wire S2563;
wire S2564;
wire S2565;
wire S2566;
wire S2567;
wire S2568;
wire S2569;
wire S2570;
wire S2571;
wire S2572;
wire S2573;
wire S2574;
wire S2575;
wire S2576;
wire S2577;
wire S2578;
wire S2579;
wire S2580;
wire S2581;
wire S2582;
wire S2583;
wire S2584;
wire S2585;
wire S2586;
wire S2587;
wire S2588;
wire S2589;
wire S2590;
wire S2591;
wire S2592;
wire S2593;
wire S2594;
wire S2595;
wire S2596;
wire S2597;
wire S2598;
wire S2599;
wire S2600;
wire S2601;
wire S2602;
wire S2603;
wire S2604;
wire S2605;
wire S2606;
wire S2607;
wire S2608;
wire S2609;
wire S2610;
wire S2611;
wire S2612;
wire S2613;
wire S2614;
wire S2615;
wire S2616;
wire S2617;
wire S2618;
wire S2619;
wire S2620;
wire S2621;
wire S2622;
wire S2623;
wire S2624;
wire S2625;
wire S2626;
wire S2627;
wire S2628;
wire S2629;
wire S2630;
wire S2631;
wire S2632;
wire S2633;
wire S2634;
wire S2635;
wire S2636;
wire S2637;
wire S2638;
wire S2639;
wire S2640;
wire S2641;
wire S2642;
wire S2643;
wire S2644;
wire S2645;
wire S2646;
wire S2647;
wire S2648;
wire S2649;
wire S2650;
wire S2651;
wire S2652;
wire S2653;
wire S2654;
wire S2655;
wire S2656;
wire S2657;
wire S2658;
wire S2659;
wire S2660;
wire S2661;
wire S2662;
wire S2663;
wire S2664;
wire S2665;
wire S2666;
wire S2667;
wire S2668;
wire S2669;
wire S2670;
wire S2671;
wire S2672;
wire S2673;
wire S2674;
wire S2675;
wire S2676;
wire S2677;
wire S2678;
wire S2679;
wire S2680;
wire S2681;
wire S2682;
wire S2683;
wire S2684;
wire S2685;
wire S2686;
wire S2687;
wire S2688;
wire S2689;
wire S2690;
wire S2691;
wire S2692;
wire S2693;
wire S2694;
wire S2695;
wire S2696;
wire S2697;
wire S2698;
wire S2699;
wire S2700;
wire S2701;
wire S2702;
wire S2703;
wire S2704;
wire S2705;
wire S2706;
wire S2707;
wire S2708;
wire S2709;
wire S2710;
wire S2711;
wire S2712;
wire S2713;
wire S2714;
wire S2715;
wire S2716;
wire S2717;
wire S2718;
wire S2719;
wire S2720;
wire S2721;
wire S2722;
wire S2723;
wire S2724;
wire S2725;
wire S2726;
wire S2727;
wire S2728;
wire S2729;
wire S2730;
wire S2731;
wire S2732;
wire S2733;
wire S2734;
wire S2735;
wire S2736;
wire S2737;
wire S2738;
wire S2739;
wire S2740;
wire S2741;
wire S2742;
wire S2743;
wire S2744;
wire S2745;
wire S2746;
wire S2747;
wire S2748;
wire S2749;
wire S2750;
wire S2751;
wire S2752;
wire S2753;
wire S2754;
wire S2755;
wire S2756;
wire S2757;
wire S2758;
wire S2759;
wire S2760;
wire S2761;
wire S2762;
wire S2763;
wire S2764;
wire S2765;
wire S2766;
wire S2767;
wire S2768;
wire S2769;
wire S2770;
wire S2771;
wire S2772;
wire S2773;
wire S2774;
wire S2775;
wire S2776;
wire S2777;
wire S2778;
wire S2779;
wire S2780;
wire S2781;
wire S2782;
wire S2783;
wire S2784;
wire S2785;
wire S2786;
wire S2787;
wire S2788;
wire S2789;
wire S2790;
wire S2791;
wire S2792;
wire S2793;
wire S2794;
wire S2795;
wire S2796;
wire S2797;
wire S2798;
wire S2799;
wire S2800;
wire S2801;
wire S2802;
wire S2803;
wire S2804;
wire S2805;
wire S2806;
wire S2807;
wire S2808;
wire S2809;
wire S2810;
wire S2811;
wire S2812;
wire S2813;
wire S2814;
wire S2815;
wire S2816;
wire S2817;
wire S2818;
wire S2819;
wire S2820;
wire S2821;
wire S2822;
wire S2823;
wire S2824;
wire S2825;
wire S2826;
wire S2827;
wire S2828;
wire S2829;
wire S2830;
wire S2831;
wire S2832;
wire S2833;
wire S2834;
wire S2835;
wire S2836;
wire S2837;
wire S2838;
wire S2839;
wire S2840;
wire S2841;
wire S2842;
wire S2843;
wire S2844;
wire S2845;
wire S2846;
wire S2847;
wire S2848;
wire S2849;
wire S2850;
wire S2851;
wire S2852;
wire S2853;
wire S2854;
wire S2855;
wire S2856;
wire S2857;
wire S2858;
wire S2859;
wire S2860;
wire S2861;
wire S2862;
wire S2863;
wire S2864;
wire S2865;
wire S2866;
wire S2867;
wire S2868;
wire S2869;
wire S2870;
wire S2871;
wire S2872;
wire S2873;
wire S2874;
wire S2875;
wire S2876;
wire S2877;
wire S2878;
wire S2879;
wire S2880;
wire S2881;
wire S2882;
wire S2883;
wire S2884;
wire S2885;
wire S2886;
wire S2887;
wire S2888;
wire S2889;
wire S2890;
wire S2891;
wire S2892;
wire S2893;
wire S2894;
wire S2895;
wire S2896;
wire S2897;
wire S2898;
wire S2899;
wire S2900;
wire S2901;
wire S2902;
wire S2903;
wire S2904;
wire S2905;
wire S2906;
wire S2907;
wire S2908;
wire S2909;
wire S2910;
wire S2911;
wire S2912;
wire S2913;
wire S2914;
wire S2915;
wire S2916;
wire S2917;
wire S2918;
wire S2919;
wire S2920;
wire S2921;
wire S2922;
wire S2923;
wire S2924;
wire S2925;
wire S2926;
wire S2927;
wire S2928;
wire S2929;
wire S2930;
wire S2931;
wire S2932;
wire S2933;
wire S2934;
wire S2935;
wire S2936;
wire S2937;
wire S2938;
wire S2939;
wire S2940;
wire S2941;
wire S2942;
wire S2943;
wire S2944;
wire S2945;
wire S2946;
wire S2947;
wire S2948;
wire S2949;
wire S2950;
wire S2951;
wire S2952;
wire S2953;
wire S2954;
wire S2955;
wire S2956;
wire S2957;
wire S2958;
wire S2959;
wire S2960;
wire S2961;
wire S2962;
wire S2963;
wire S2964;
wire S2965;
wire S2966;
wire S2967;
wire S2968;
wire S2969;
wire S2970;
wire S2971;
wire S2972;
wire S2973;
wire S2974;
wire S2975;
wire S2976;
wire S2977;
wire S2978;
wire S2979;
wire S2980;
wire S2981;
wire S2982;
wire S2983;
wire S2984;
wire S2985;
wire S2986;
wire S2987;
wire S2988;
wire S2989;
wire S2990;
wire S2991;
wire S2992;
wire S2993;
wire S2994;
wire S2995;
wire S2996;
wire S2997;
wire S2998;
wire S2999;
wire S3000;
wire S3001;
wire S3002;
wire S3003;
wire S3004;
wire S3005;
wire S3006;
wire S3007;
wire S3008;
wire S3009;
wire S3010;
wire S3011;
wire S3012;
wire S3013;
wire S3014;
wire S3015;
wire S3016;
wire S3017;
wire S3018;
wire S3019;
wire S3020;
wire S3021;
wire S3022;
wire S3023;
wire S3024;
wire S3025;
wire S3026;
wire S3027;
wire S3028;
wire S3029;
wire S3030;
wire S3031;
wire S3032;
wire S3033;
wire S3034;
wire S3035;
wire S3036;
wire S3037;
wire S3038;
wire S3039;
wire S3040;
wire S3041;
wire S3042;
wire S3043;
wire S3044;
wire S3045;
wire S3046;
wire S3047;
wire S3048;
wire S3049;
wire S3050;
wire S3051;
wire S3052;
wire S3053;
wire S3054;
wire S3055;
wire S3056;
wire S3057;
wire S3058;
wire S3059;
wire S3060;
wire S3061;
wire S3062;
wire S3063;
wire S3064;
wire S3065;
wire S3066;
wire S3067;
wire S3068;
wire S3069;
wire S3070;
wire S3071;
wire S3072;
wire S3073;
wire S3074;
wire S3075;
wire S3076;
wire S3077;
wire S3078;
wire S3079;
wire S3080;
wire S3081;
wire S3082;
wire S3083;
wire S3084;
wire S3085;
wire S3086;
wire S3087;
wire S3088;
wire S3089;
wire S3090;
wire S3091;
wire S3092;
wire S3093;
wire S3094;
wire S3095;
wire S3096;
wire S3097;
wire S3098;
wire S3099;
wire S3100;
wire S3101;
wire S3102;
wire S3103;
wire S3104;
wire S3105;
wire S3106;
wire S3107;
wire S3108;
wire S3109;
wire S3110;
wire S3111;
wire S3112;
wire S3113;
wire S3114;
wire S3115;
wire S3116;
wire S3117;
wire S3118;
wire S3119;
wire S3120;
wire S3121;
wire S3122;
wire S3123;
wire S3124;
wire S3125;
wire S3126;
wire S3127;
wire S3128;
wire S3129;
wire S3130;
wire S3131;
wire S3132;
wire S3133;
wire S3134;
wire S3135;
wire S3136;
wire S3137;
wire S3138;
wire S3139;
wire S3140;
wire S3141;
wire S3142;
wire S3143;
wire S3144;
wire S3145;
wire S3146;
wire S3147;
wire S3148;
wire S3149;
wire S3150;
wire S3151;
wire S3152;
wire S3153;
wire S3154;
wire S3155;
wire S3156;
wire S3157;
wire S3158;
wire S3159;
wire S3160;
wire S3161;
wire S3162;
wire S3163;
wire S3164;
wire S3165;
wire S3166;
wire S3167;
wire S3168;
wire S3169;
wire S3170;
wire S3171;
wire S3172;
wire S3173;
wire S3174;
wire S3175;
wire S3176;
wire S3177;
wire S3178;
wire S3179;
wire S3180;
wire S3181;
wire S3182;
wire S3183;
wire S3184;
wire S3185;
wire S3186;
wire S3187;
wire S3188;
wire S3189;
wire S3190;
wire S3191;
wire S3192;
wire S3193;
wire S3194;
wire S3195;
wire S3196;
wire S3197;
wire S3198;
wire S3199;
wire S3200;
wire S3201;
wire S3202;
wire S3203;
wire S3204;
wire S3205;
wire S3206;
wire S3207;
wire S3208;
wire S3209;
wire S3210;
wire S3211;
wire S3212;
wire S3213;
wire S3214;
wire S3215;
wire S3216;
wire S3217;
wire S3218;
wire S3219;
wire S3220;
wire S3221;
wire S3222;
wire S3223;
wire S3224;
wire S3225;
wire S3226;
wire S3227;
wire S3228;
wire S3229;
wire S3230;
wire S3231;
wire S3232;
wire S3233;
wire S3234;
wire S3235;
wire S3236;
wire S3237;
wire S3238;
wire S3239;
wire S3240;
wire S3241;
wire S3242;
wire S3243;
wire S3244;
wire S3245;
wire S3246;
wire S3247;
wire S3248;
wire S3249;
wire S3250;
wire S3251;
wire S3252;
wire S3253;
wire S3254;
wire S3255;
wire S3256;
wire S3257;
wire S3258;
wire S3259;
wire S3260;
wire S3261;
wire S3262;
wire S3263;
wire S3264;
wire S3265;
wire S3266;
wire S3267;
wire S3268;
wire S3269;
wire S3270;
wire S3271;
wire S3272;
wire S3273;
wire S3274;
wire S3275;
wire S3276;
wire S3277;
wire S3278;
wire S3279;
wire S3280;
wire S3281;
wire S3282;
wire S3283;
wire S3284;
wire S3285;
wire S3286;
wire S3287;
wire S3288;
wire S3289;
wire S3290;
wire S3291;
wire S3292;
wire S3293;
wire S3294;
wire S3295;
wire S3296;
wire S3297;
wire S3298;
wire S3299;
wire S3300;
wire S3301;
wire S3302;
wire S3303;
wire S3304;
wire S3305;
wire S3306;
wire S3307;
wire S3308;
wire S3309;
wire S3310;
wire S3311;
wire S3312;
wire S3313;
wire S3314;
wire S3315;
wire S3316;
wire S3317;
wire S3318;
wire S3319;
wire S3320;
wire S3321;
wire S3322;
wire S3323;
wire S3324;
wire S3325;
wire S3326;
wire S3327;
wire S3328;
wire S3329;
wire S3330;
wire S3331;
wire S3332;
wire S3333;
wire S3334;
wire S3335;
wire S3336;
wire S3337;
wire S3338;
wire S3339;
wire S3340;
wire S3341;
wire S3342;
wire S3343;
wire S3344;
wire S3345;
wire S3346;
wire S3347;
wire S3348;
wire S3349;
wire S3350;
wire S3351;
wire S3352;
wire S3353;
wire S3354;
wire S3355;
wire S3356;
wire S3357;
wire S3358;
wire S3359;
wire S3360;
wire S3361;
wire S3362;
wire S3363;
wire S3364;
wire S3365;
wire S3366;
wire S3367;
wire S3368;
wire S3369;
wire S3370;
wire S3371;
wire S3372;
wire S3373;
wire S3374;
wire S3375;
wire S3376;
wire S3377;
wire S3378;
wire S3379;
wire S3380;
wire S3381;
wire S3382;
wire S3383;
wire S3384;
wire S3385;
wire S3386;
wire S3387;
wire S3388;
wire S3389;
wire S3390;
wire S3391;
wire S3392;
wire S3393;
wire S3394;
wire S3395;
wire S3396;
wire S3397;
wire S3398;
wire S3399;
wire S3400;
wire S3401;
wire S3402;
wire S3403;
wire S3404;
wire S3405;
wire S3406;
wire S3407;
wire S3408;
wire S3409;
wire S3410;
wire S3411;
wire S3412;
wire S3413;
wire S3414;
wire S3415;
wire S3416;
wire S3417;
wire S3418;
wire S3419;
wire S3420;
wire S3421;
wire S3422;
wire S3423;
wire S3424;
wire S3425;
wire S3426;
wire S3427;
wire S3428;
wire S3429;
wire S3430;
wire S3431;
wire S3432;
wire S3433;
wire S3434;
wire S3435;
wire S3436;
wire S3437;
wire S3438;
wire S3439;
wire S3440;
wire S3441;
wire S3442;
wire S3443;
wire S3444;
wire S3445;
wire S3446;
wire S3447;
wire S3448;
wire S3449;
wire S3450;
wire S3451;
wire S3452;
wire S3453;
wire S3454;
wire S3455;
wire S3456;
wire S3457;
wire S3458;
wire S3459;
wire S3460;
wire S3461;
wire S3462;
wire S3463;
wire S3464;
wire S3465;
wire S3466;
wire S3467;
wire S3468;
wire S3469;
wire S3470;
wire S3471;
wire S3472;
wire S3473;
wire S3474;
wire S3475;
wire S3476;
wire S3477;
wire S3478;
wire S3479;
wire S3480;
wire S3481;
wire S3482;
wire S3483;
wire S3484;
wire S3485;
wire S3486;
wire S3487;
wire S3488;
wire S3489;
wire S3490;
wire S3491;
wire S3492;
wire S3493;
wire S3494;
wire S3495;
wire S3496;
wire S3497;
wire S3498;
wire S3499;
wire S3500;
wire S3501;
wire S3502;
wire S3503;
wire S3504;
wire S3505;
wire S3506;
wire S3507;
wire S3508;
wire S3509;
wire S3510;
wire S3511;
wire S3512;
wire S3513;
wire S3514;
wire S3515;
wire S3516;
wire S3517;
wire S3518;
wire S3519;
wire S3520;
wire S3521;
wire S3522;
wire S3523;
wire S3524;
wire S3525;
wire S3526;
wire S3527;
wire S3528;
wire S3529;
wire S3530;
wire S3531;
wire S3532;
wire S3533;
wire S3534;
wire S3535;
wire S3536;
wire S3537;
wire S3538;
wire S3539;
wire S3540;
wire S3541;
wire S3542;
wire S3543;
wire S3544;
wire S3545;
wire S3546;
wire S3547;
wire S3548;
wire S3549;
wire S3550;
wire S3551;
wire S3552;
wire S3553;
wire S3554;
wire S3555;
wire S3556;
wire S3557;
wire S3558;
wire S3559;
wire S3560;
wire S3561;
wire S3562;
wire S3563;
wire S3564;
wire S3565;
wire S3566;
wire S3567;
wire S3568;
wire S3569;
wire S3570;
wire S3571;
wire S3572;
wire S3573;
wire S3574;
wire S3575;
wire S3576;
wire S3577;
wire S3578;
wire S3579;
wire S3580;
wire S3581;
wire S3582;
wire S3583;
wire S3584;
wire S3585;
wire S3586;
wire S3587;
wire S3588;
wire S3589;
wire S3590;
wire S3591;
wire S3592;
wire S3593;
wire S3594;
wire S3595;
wire S3596;
wire S3597;
wire S3598;
wire S3599;
wire S3600;
wire S3601;
wire S3602;
wire S3603;
wire S3604;
wire S3605;
wire S3606;
wire S3607;
wire S3608;
wire S3609;
wire S3610;
wire S3611;
wire S3612;
wire S3613;
wire S3614;
wire S3615;
wire S3616;
wire S3617;
wire S3618;
wire S3619;
wire S3620;
wire S3621;
wire S3622;
wire S3623;
wire S3624;
wire S3625;
wire S3626;
wire S3627;
wire S3628;
wire S3629;
wire S3630;
wire S3631;
wire S3632;
wire S3633;
wire S3634;
wire S3635;
wire S3636;
wire S3637;
wire S3638;
wire S3639;
wire S3640;
wire S3641;
wire S3642;
wire S3643;
wire S3644;
wire S3645;
wire S3646;
wire S3647;
wire S3648;
wire S3649;
wire S3650;
wire S3651;
wire S3652;
wire S3653;
wire S3654;
wire S3655;
wire S3656;
wire S3657;
wire S3658;
wire S3659;
wire S3660;
wire S3661;
wire S3662;
wire S3663;
wire S3664;
wire S3665;
wire S3666;
wire S3667;
wire S3668;
wire S3669;
wire S3670;
wire S3671;
wire S3672;
wire S3673;
wire S3674;
wire S3675;
wire S3676;
wire S3677;
wire S3678;
wire S3679;
wire S3680;
wire S3681;
wire S3682;
wire S3683;
wire S3684;
wire S3685;
wire S3686;
wire S3687;
wire S3688;
wire S3689;
wire S3690;
wire S3691;
wire S3692;
wire S3693;
wire S3694;
wire S3695;
wire S3696;
wire S3697;
wire S3698;
wire S3699;
wire S3700;
wire S3701;
wire S3702;
wire S3703;
wire S3704;
wire S3705;
wire S3706;
wire S3707;
wire S3708;
wire S3709;
wire S3710;
wire S3711;
wire S3712;
wire S3713;
wire S3714;
wire S3715;
wire S3716;
wire S3717;
wire S3718;
wire S3719;
wire S3720;
wire S3721;
wire S3722;
wire S3723;
wire S3724;
wire S3725;
wire S3726;
wire S3727;
wire S3728;
wire S3729;
wire S3730;
wire S3731;
wire S3732;
wire S3733;
wire S3734;
wire S3735;
wire S3736;
wire S3737;
wire S3738;
wire S3739;
wire S3740;
wire S3741;
wire S3742;
wire S3743;
wire S3744;
wire S3745;
wire S3746;
wire S3747;
wire S3748;
wire S3749;
wire S3750;
wire S3751;
wire S3752;
wire S3753;
wire S3754;
wire S3755;
wire S3756;
wire S3757;
wire S3758;
wire S3759;
wire S3760;
wire S3761;
wire S3762;
wire S3763;
wire S3764;
wire S3765;
wire S3766;
wire S3767;
wire S3768;
wire S3769;
wire S3770;
wire S3771;
wire S3772;
wire S3773;
wire S3774;
wire S3775;
wire S3776;
wire S3777;
wire S3778;
wire S3779;
wire S3780;
wire S3781;
wire S3782;
wire S3783;
wire S3784;
wire S3785;
wire S3786;
wire S3787;
wire S3788;
wire S3789;
wire S3790;
wire S3791;
wire S3792;
wire S3793;
wire S3794;
wire S3795;
wire S3796;
wire S3797;
wire S3798;
wire S3799;
wire S3800;
wire S3801;
wire S3802;
wire S3803;
wire S3804;
wire S3805;
wire S3806;
wire S3807;
wire S3808;
wire S3809;
wire S3810;
wire S3811;
wire S3812;
wire S3813;
wire S3814;
wire S3815;
wire S3816;
wire S3817;
wire S3818;
wire S3819;
wire S3820;
wire S3821;
wire S3822;
wire S3823;
wire S3824;
wire S3825;
wire S3826;
wire S3827;
wire S3828;
wire S3829;
wire S3830;
wire S3831;
wire S3832;
wire S3833;
wire S3834;
wire S3835;
wire S3836;
wire S3837;
wire S3838;
wire S3839;
wire S3840;
wire S3841;
wire S3842;
wire S3843;
wire S3844;
wire S3845;
wire S3846;
wire S3847;
wire S3848;
wire S3849;
wire S3850;
wire S3851;
wire S3852;
wire S3853;
wire S3854;
wire S3855;
wire S3856;
wire S3857;
wire S3858;
wire S3859;
wire S3860;
wire S3861;
wire S3862;
wire S3863;
wire S3864;
wire S3865;
wire S3866;
wire S3867;
wire S3868;
wire S3869;
wire S3870;
wire S3871;
wire S3872;
wire S3873;
wire S3874;
wire S3875;
wire S3876;
wire S3877;
wire S3878;
wire S3879;
wire S3880;
wire S3881;
wire S3882;
wire S3883;
wire S3884;
wire S3885;
wire S3886;
wire S3887;
wire S3888;
wire S3889;
wire S3890;
wire S3891;
wire S3892;
wire S3893;
wire S3894;
wire S3895;
wire S3896;
wire S3897;
wire S3898;
wire S3899;
wire S3900;
wire S3901;
wire S3902;
wire S3903;
wire S3904;
wire S3905;
wire S3906;
wire S3907;
wire S3908;
wire S3909;
wire S3910;
wire S3911;
wire S3912;
wire S3913;
wire S3914;
wire S3915;
wire S3916;
wire S3917;
wire S3918;
wire S3919;
wire S3920;
wire S3921;
wire S3922;
wire S3923;
wire S3924;
wire S3925;
wire S3926;
wire S3927;
wire S3928;
wire S3929;
wire S3930;
wire S3931;
wire S3932;
wire S3933;
wire S3934;
wire S3935;
wire S3936;
wire S3937;
wire S3938;
wire S3939;
wire S3940;
wire S3941;
wire S3942;
wire S3943;
wire S3944;
wire S3945;
wire S3946;
wire S3947;
wire S3948;
wire S3949;
wire S3950;
wire S3951;
wire S3952;
wire S3953;
wire S3954;
wire S3955;
wire S3956;
wire S3957;
wire S3958;
wire S3959;
wire S3960;
wire S3961;
wire S3962;
wire S3963;
wire S3964;
wire S3965;
wire S3966;
wire S3967;
wire S3968;
wire S3969;
wire S3970;
wire S3971;
wire S3972;
wire S3973;
wire S3974;
wire S3975;
wire S3976;
wire S3977;
wire S3978;
wire S3979;
wire S3980;
wire S3981;
wire S3982;
wire S3983;
wire S3984;
wire S3985;
wire S3986;
wire S3987;
wire S3988;
wire S3989;
wire S3990;
wire S3991;
wire S3992;
wire S3993;
wire S3994;
wire S3995;
wire S3996;
wire S3997;
wire S3998;
wire S3999;
wire S4000;
wire S4001;
wire S4002;
wire S4003;
wire S4004;
wire S4005;
wire S4006;
wire S4007;
wire S4008;
wire S4009;
wire S4010;
wire S4011;
wire S4012;
wire S4013;
wire S4014;
wire S4015;
wire S4016;
wire S4017;
wire S4018;
wire S4019;
wire S4020;
wire S4021;
wire S4022;
wire S4023;
wire S4024;
wire S4025;
wire S4026;
wire S4027;
wire S4028;
wire S4029;
wire S4030;
wire S4031;
wire S4032;
wire S4033;
wire S4034;
wire S4035;
wire S4036;
wire S4037;
wire S4038;
wire S4039;
wire S4040;
wire S4041;
wire S4042;
wire S4043;
wire S4044;
wire S4045;
wire S4046;
wire S4047;
wire S4048;
wire S4049;
wire S4050;
wire S4051;
wire S4052;
wire S4053;
wire S4054;
wire S4055;
wire S4056;
wire S4057;
wire S4058;
wire S4059;
wire S4060;
wire S4061;
wire S4062;
wire S4063;
wire S4064;
wire S4065;
wire S4066;
wire S4067;
wire S4068;
wire S4069;
wire S4070;
wire S4071;
wire S4072;
wire S4073;
wire S4074;
wire S4075;
wire S4076;
wire S4077;
wire S4078;
wire S4079;
wire S4080;
wire S4081;
wire S4082;
wire S4083;
wire S4084;
wire S4085;
wire S4086;
wire S4087;
wire S4088;
wire S4089;
wire S4090;
wire S4091;
wire S4092;
wire S4093;
wire S4094;
wire S4095;
wire S4096;
wire S4097;
wire S4098;
wire S4099;
wire S4100;
wire S4101;
wire S4102;
wire S4103;
wire S4104;
wire S4105;
wire S4106;
wire S4107;
wire S4108;
wire S4109;
wire S4110;
wire S4111;
wire S4112;
wire S4113;
wire S4114;
wire S4115;
wire S4116;
wire S4117;
wire S4118;
wire S4119;
wire S4120;
wire S4121;
wire S4122;
wire S4123;
wire S4124;
wire S4125;
wire S4126;
wire S4127;
wire S4128;
wire S4129;
wire S4130;
wire S4131;
wire S4132;
wire S4133;
wire S4134;
wire S4135;
wire S4136;
wire S4137;
wire S4138;
wire S4139;
wire S4140;
wire S4141;
wire S4142;
wire S4143;
wire S4144;
wire S4145;
wire S4146;
wire S4147;
wire S4148;
wire S4149;
wire S4150;
wire S4151;
wire S4152;
wire S4153;
wire S4154;
wire S4155;
wire S4156;
wire S4157;
wire S4158;
wire S4159;
wire S4160;
wire S4161;
wire S4162;
wire S4163;
wire S4164;
wire S4165;
wire S4166;
wire S4167;
wire S4168;
wire S4169;
wire S4170;
wire S4171;
wire S4172;
wire S4173;
wire S4174;
wire S4175;
wire S4176;
wire S4177;
wire S4178;
wire S4179;
wire S4180;
wire S4181;
wire S4182;
wire S4183;
wire S4184;
wire S4185;
wire S4186;
wire S4187;
wire S4188;
wire S4189;
wire S4190;
wire S4191;
wire S4192;
wire S4193;
wire S4194;
wire S4195;
wire S4196;
wire S4197;
wire S4198;
wire S4199;
wire S4200;
wire S4201;
wire S4202;
wire S4203;
wire S4204;
wire S4205;
wire S4206;
wire S4207;
wire S4208;
wire S4209;
wire S4210;
wire S4211;
wire S4212;
wire S4213;
wire S4214;
wire S4215;
wire S4216;
wire S4217;
wire S4218;
wire S4219;
wire S4220;
wire S4221;
wire S4222;
wire S4223;
wire S4224;
wire S4225;
wire S4226;
wire S4227;
wire S4228;
wire S4229;
wire S4230;
wire S4231;
wire S4232;
wire S4233;
wire S4234;
wire S4235;
wire S4236;
wire S4237;
wire S4238;
wire S4239;
wire S4240;
wire S4241;
wire S4242;
wire S4243;
wire S4244;
wire S4245;
wire S4246;
wire S4247;
wire S4248;
wire S4249;
wire S4250;
wire S4251;
wire S4252;
wire S4253;
wire S4254;
wire S4255;
wire S4256;
wire S4257;
wire S4258;
wire S4259;
wire S4260;
wire S4261;
wire S4262;
wire S4263;
wire S4264;
wire S4265;
wire S4266;
wire S4267;
wire S4268;
wire S4269;
wire S4270;
wire S4271;
wire S4272;
wire S4273;
wire S4274;
wire S4275;
wire S4276;
wire S4277;
wire S4278;
wire S4279;
wire S4280;
wire S4281;
wire S4282;
wire S4283;
wire S4284;
wire S4285;
wire S4286;
wire S4287;
wire S4288;
wire S4289;
wire S4290;
wire S4291;
wire S4292;
wire S4293;
wire S4294;
wire S4295;
wire S4296;
wire S4297;
wire S4298;
wire S4299;
wire S4300;
wire S4301;
wire S4302;
wire S4303;
wire S4304;
wire S4305;
wire S4306;
wire S4307;
wire S4308;
wire S4309;
wire S4310;
wire S4311;
wire S4312;
wire S4313;
wire S4314;
wire S4315;
wire S4316;
wire S4317;
wire S4318;
wire S4319;
wire S4320;
wire S4321;
wire S4322;
wire S4323;
wire S4324;
wire S4325;
wire S4326;
wire S4327;
wire S4328;
wire S4329;
wire S4330;
wire S4331;
wire S4332;
wire S4333;
wire S4334;
wire S4335;
wire S4336;
wire S4337;
wire S4338;
wire S4339;
wire S4340;
wire S4341;
wire S4342;
wire S4343;
wire S4344;
wire S4345;
wire S4346;
wire S4347;
wire S4348;
wire S4349;
wire S4350;
wire S4351;
wire S4352;
wire S4353;
wire S4354;
wire S4355;
wire S4356;
wire S4357;
wire S4358;
wire S4359;
wire S4360;
wire S4361;
wire S4362;
wire S4363;
wire S4364;
wire S4365;
wire S4366;
wire S4367;
wire S4368;
wire S4369;
wire S4370;
wire S4371;
wire S4372;
wire S4373;
wire S4374;
wire S4375;
wire S4376;
wire S4377;
wire S4378;
wire S4379;
wire S4380;
wire S4381;
wire S4382;
wire S4383;
wire S4384;
wire S4385;
wire S4386;
wire S4387;
wire S4388;
wire S4389;
wire S4390;
wire S4391;
wire S4392;
wire S4393;
wire S4394;
wire S4395;
wire S4396;
wire S4397;
wire S4398;
wire S4399;
wire S4400;
wire S4401;
wire S4402;
wire S4403;
wire S4404;
wire S4405;
wire S4406;
wire S4407;
wire S4408;
wire S4409;
wire S4410;
wire S4411;
wire S4412;
wire S4413;
wire S4414;
wire S4415;
wire S4416;
wire S4417;
wire S4418;
wire S4419;
wire S4420;
wire S4421;
wire S4422;
wire S4423;
wire S4424;
wire S4425;
wire S4426;
wire S4427;
wire S4428;
wire S4429;
wire S4430;
wire S4431;
wire S4432;
wire S4433;
wire S4434;
wire S4435;
wire S4436;
wire S4437;
wire S4438;
wire S4439;
wire S4440;
wire S4441;
wire S4442;
wire S4443;
wire S4444;
wire S4445;
wire S4446;
wire S4447;
wire S4448;
wire S4449;
wire S4450;
wire S4451;
wire S4452;
wire S4453;
wire S4454;
wire S4455;
wire S4456;
wire S4457;
wire S4458;
wire S4459;
wire S4460;
wire S4461;
wire S4462;
wire S4463;
wire S4464;
wire S4465;
wire S4466;
wire S4467;
wire S4468;
wire S4469;
wire S4470;
wire S4471;
wire S4472;
wire S4473;
wire S4474;
wire S4475;
wire S4476;
wire S4477;
wire S4478;
wire S4479;
wire S4480;
wire S4481;
wire S4482;
wire S4483;
wire S4484;
wire S4485;
wire S4486;
wire S4487;
wire S4488;
wire S4489;
wire S4490;
wire S4491;
wire S4492;
wire S4493;
wire S4494;
wire S4495;
wire S4496;
wire S4497;
wire S4498;
wire S4499;
wire S4500;
wire S4501;
wire S4502;
wire S4503;
wire S4504;
wire S4505;
wire S4506;
wire S4507;
wire S4508;
wire S4509;
wire S4510;
wire S4511;
wire S4512;
wire S4513;
wire S4514;
wire S4515;
wire S4516;
wire S4517;
wire S4518;
wire S4519;
wire S4520;
wire S4521;
wire S4522;
wire S4523;
wire S4524;
wire S4525;
wire S4526;
wire S4527;
wire S4528;
wire S4529;
wire S4530;
wire S4531;
wire S4532;
wire S4533;
wire S4534;
wire S4535;
wire S4536;
wire S4537;
wire S4538;
wire S4539;
wire S4540;
wire S4541;
wire S4542;
wire S4543;
wire S4544;
wire S4545;
wire S4546;
wire S4547;
wire S4548;
wire S4549;
wire S4550;
wire S4551;
wire S4552;
wire S4553;
wire S4554;
wire S4555;
wire S4556;
wire S4557;
wire S4558;
wire S4559;
wire S4560;
wire S4561;
wire S4562;
wire S4563;
wire S4564;
wire S4565;
wire S4566;
wire S4567;
wire S4568;
wire S4569;
wire S4570;
wire S4571;
wire S4572;
wire S4573;
wire S4574;
wire S4575;
wire S4576;
wire S4577;
wire S4578;
wire S4579;
wire S4580;
wire S4581;
wire S4582;
wire S4583;
wire S4584;
wire S4585;
wire S4586;
wire S4587;
wire S4588;
wire S4589;
wire S4590;
wire S4591;
wire S4592;
wire S4593;
wire S4594;
wire S4595;
wire S4596;
wire S4597;
wire S4598;
wire S4599;
wire S4600;
wire S4601;
wire S4602;
wire S4603;
wire S4604;
wire S4605;
wire S4606;
wire S4607;
wire S4608;
wire S4609;
wire S4610;
wire S4611;
wire S4612;
wire S4613;
wire S4614;
wire S4615;
wire S4616;
wire S4617;
wire S4618;
wire S4619;
wire S4620;
wire S4621;
wire S4622;
wire S4623;
wire S4624;
wire S4625;
wire S4626;
wire S4627;
wire S4628;
wire S4629;
wire S4630;
wire S4631;
wire S4632;
wire S4633;
wire S4634;
wire S4635;
wire S4636;
wire S4637;
wire S4638;
wire S4639;
wire S4640;
wire S4641;
wire S4642;
wire S4643;
wire S4644;
wire S4645;
wire S4646;
wire S4647;
wire S4648;
wire S4649;
wire S4650;
wire S4651;
wire S4652;
wire S4653;
wire S4654;
wire S4655;
wire S4656;
wire S4657;
wire S4658;
wire S4659;
wire S4660;
wire S4661;
wire S4662;
wire S4663;
wire S4664;
wire S4665;
wire S4666;
wire S4667;
wire S4668;
wire S4669;
wire S4670;
wire S4671;
wire S4672;
wire S4673;
wire S4674;
wire S4675;
wire S4676;
wire S4677;
wire S4678;
wire S4679;
wire S4680;
wire S4681;
wire S4682;
wire S4683;
wire S4684;
wire S4685;
wire S4686;
wire S4687;
wire S4688;
wire S4689;
wire S4690;
wire S4691;
wire S4692;
wire S4693;
wire S4694;
wire S4695;
wire S4696;
wire S4697;
wire S4698;
wire S4699;
wire S4700;
wire S4701;
wire S4702;
wire S4703;
wire S4704;
wire S4705;
wire S4706;
wire S4707;
wire S4708;
wire S4709;
wire S4710;
wire S4711;
wire S4712;
wire S4713;
wire S4714;
wire S4715;
wire S4716;
wire S4717;
wire S4718;
wire S4719;
wire S4720;
wire S4721;
wire S4722;
wire S4723;
wire S4724;
wire S4725;
wire S4726;
wire S4727;
wire S4728;
wire S4729;
wire S4730;
wire S4731;
wire S4732;
wire S4733;
wire S4734;
wire S4735;
wire S4736;
wire S4737;
wire S4738;
wire S4739;
wire S4740;
wire S4741;
wire S4742;
wire S4743;
wire S4744;
wire S4745;
wire S4746;
wire S4747;
wire S4748;
wire S4749;
wire S4750;
wire S4751;
wire S4752;
wire S4753;
wire S4754;
wire S4755;
wire S4756;
wire S4757;
wire S4758;
wire S4759;
wire S4760;
wire S4761;
wire S4762;
wire S4763;
wire S4764;
wire S4765;
wire S4766;
wire S4767;
wire S4768;
wire S4769;
wire S4770;
wire S4771;
wire S4772;
wire S4773;
wire S4774;
wire S4775;
wire S4776;
wire S4777;
wire S4778;
wire S4779;
wire S4780;
wire S4781;
wire S4782;
wire S4783;
wire S4784;
wire S4785;
wire S4786;
wire S4787;
wire S4788;
wire S4789;
wire S4790;
wire S4791;
wire S4792;
wire S4793;
wire S4794;
wire S4795;
wire S4796;
wire S4797;
wire S4798;
wire S4799;
wire S4800;
wire S4801;
wire S4802;
wire S4803;
wire S4804;
wire S4805;
wire S4806;
wire S4807;
wire S4808;
wire S4809;
wire S4810;
wire S4811;
wire S4812;
wire S4813;
wire S4814;
wire S4815;
wire S4816;
wire S4817;
wire S4818;
wire S4819;
wire S4820;
wire S4821;
wire S4822;
wire S4823;
wire S4824;
wire S4825;
wire S4826;
wire S4827;
wire S4828;
wire S4829;
wire S4830;
wire S4831;
wire S4832;
wire S4833;
wire S4834;
wire S4835;
wire S4836;
wire S4837;
wire S4838;
wire S4839;
wire S4840;
wire S4841;
wire S4842;
wire S4843;
wire S4844;
wire S4845;
wire S4846;
wire S4847;
wire S4848;
wire S4849;
wire S4850;
wire S4851;
wire S4852;
wire S4853;
wire S4854;
wire S4855;
wire S4856;
wire S4857;
wire S4858;
wire S4859;
wire S4860;
wire S4861;
wire S4862;
wire S4863;
wire S4864;
wire S4865;
wire S4866;
wire S4867;
wire S4868;
wire S4869;
wire S4870;
wire S4871;
wire S4872;
wire S4873;
wire S4874;
wire S4875;
wire S4876;
wire S4877;
wire S4878;
wire S4879;
wire S4880;
wire S4881;
wire S4882;
wire S4883;
wire S4884;
wire S4885;
wire S4886;
wire S4887;
wire S4888;
wire S4889;
wire S4890;
wire S4891;
wire S4892;
wire S4893;
wire S4894;
wire S4895;
wire S4896;
wire S4897;
wire S4898;
wire S4899;
wire S4900;
wire S4901;
wire S4902;
wire S4903;
wire S4904;
wire S4905;
wire S4906;
wire S4907;
wire S4908;
wire S4909;
wire S4910;
wire S4911;
wire S4912;
wire S4913;
wire S4914;
wire S4915;
wire S4916;
wire S4917;
wire S4918;
wire S4919;
wire S4920;
wire S4921;
wire S4922;
wire S4923;
wire S4924;
wire S4925;
wire S4926;
wire S4927;
wire S4928;
wire S4929;
wire S4930;
wire S4931;
wire S4932;
wire S4933;
wire S4934;
wire S4935;
wire S4936;
wire S4937;
wire S4938;
wire S4939;
wire S4940;
wire S4941;
wire S4942;
wire S4943;
wire S4944;
wire S4945;
wire S4946;
wire S4947;
wire S4948;
wire S4949;
wire S4950;
wire S4951;
wire S4952;
wire S4953;
wire S4954;
wire S4955;
wire S4956;
wire S4957;
wire S4958;
wire S4959;
wire S4960;
wire S4961;
wire S4962;
wire S4963;
wire S4964;
wire S4965;
wire S4966;
wire S4967;
wire S4968;
wire S4969;
wire S4970;
wire S4971;
wire S4972;
wire S4973;
wire S4974;
wire S4975;
wire S4976;
wire S4977;
wire S4978;
wire S4979;
wire S4980;
wire S4981;
wire S4982;
wire S4983;
wire S4984;
wire S4985;
wire S4986;
wire S4987;
wire S4988;
wire S4989;
wire S4990;
wire S4991;
wire S4992;
wire S4993;
wire S4994;
wire S4995;
wire S4996;
wire S4997;
wire S4998;
wire S4999;
wire S5000;
wire S5001;
wire S5002;
wire S5003;
wire S5004;
wire S5005;
wire S5006;
wire S5007;
wire S5008;
wire S5009;
wire S5010;
wire S5011;
wire S5012;
wire S5013;
wire S5014;
wire S5015;
wire S5016;
wire S5017;
wire S5018;
wire S5019;
wire S5020;
wire S5021;
wire S5022;
wire S5023;
wire S5024;
wire S5025;
wire S5026;
wire S5027;
wire S5028;
wire S5029;
wire S5030;
wire S5031;
wire S5032;
wire S5033;
wire S5034;
wire S5035;
wire S5036;
wire S5037;
wire S5038;
wire S5039;
wire S5040;
wire S5041;
wire S5042;
wire S5043;
wire S5044;
wire S5045;
wire S5046;
wire S5047;
wire S5048;
wire S5049;
wire S5050;
wire S5051;
wire S5052;
wire S5053;
wire S5054;
wire S5055;
wire S5056;
wire S5057;
wire S5058;
wire S5059;
wire S5060;
wire S5061;
wire S5062;
wire S5063;
wire S5064;
wire S5065;
wire S5066;
wire S5067;
wire S5068;
wire S5069;
wire S5070;
wire S5071;
wire S5072;
wire S5073;
wire S5074;
wire S5075;
wire S5076;
wire S5077;
wire S5078;
wire S5079;
wire S5080;
wire S5081;
wire S5082;
wire S5083;
wire S5084;
wire S5085;
wire S5086;
wire S5087;
wire S5088;
wire S5089;
wire S5090;
wire S5091;
wire S5092;
wire S5093;
wire S5094;
wire S5095;
wire S5096;
wire S5097;
wire S5098;
wire S5099;
wire S5100;
wire S5101;
wire S5102;
wire S5103;
wire S5104;
wire S5105;
wire S5106;
wire S5107;
wire S5108;
wire S5109;
wire S5110;
wire S5111;
wire S5112;
wire S5113;
wire S5114;
wire S5115;
wire S5116;
wire S5117;
wire S5118;
wire S5119;
wire S5120;
wire S5121;
wire S5122;
wire S5123;
wire S5124;
wire S5125;
wire S5126;
wire S5127;
wire S5128;
wire S5129;
wire S5130;
wire S5131;
wire S5132;
wire S5133;
wire S5134;
wire S5135;
wire S5136;
wire S5137;
wire S5138;
wire S5139;
wire S5140;
wire S5141;
wire S5142;
wire S5143;
wire S5144;
wire S5145;
wire S5146;
wire S5147;
wire S5148;
wire S5149;
wire S5150;
wire S5151;
wire S5152;
wire S5153;
wire S5154;
wire S5155;
wire S5156;
wire S5157;
wire S5158;
wire S5159;
wire S5160;
wire S5161;
wire S5162;
wire S5163;
wire S5164;
wire S5165;
wire S5166;
wire S5167;
wire S5168;
wire S5169;
wire S5170;
wire S5171;
wire S5172;
wire S5173;
wire S5174;
wire S5175;
wire S5176;
wire S5177;
wire S5178;
wire S5179;
wire S5180;
wire S5181;
wire S5182;
wire S5183;
wire S5184;
wire S5185;
wire S5186;
wire S5187;
wire S5188;
wire S5189;
wire S5190;
wire S5191;
wire S5192;
wire S5193;
wire S5194;
wire S5195;
wire S5196;
wire S5197;
wire S5198;
wire S5199;
wire S5200;
wire S5201;
wire S5202;
wire S5203;
wire S5204;
wire S5205;
wire S5206;
wire S5207;
wire S5208;
wire S5209;
wire S5210;
wire S5211;
wire S5212;
wire S5213;
wire S5214;
wire S5215;
wire S5216;
wire S5217;
wire S5218;
wire S5219;
wire S5220;
wire S5221;
wire S5222;
wire S5223;
wire S5224;
wire S5225;
wire S5226;
wire S5227;
wire S5228;
wire S5229;
wire S5230;
wire S5231;
wire S5232;
wire S5233;
wire S5234;
wire S5235;
wire S5236;
wire S5237;
wire S5238;
wire S5239;
wire S5240;
wire S5241;
wire S5242;
wire S5243;
wire S5244;
wire S5245;
wire S5246;
wire S5247;
wire S5248;
wire S5249;
wire S5250;
wire S5251;
wire S5252;
wire S5253;
wire S5254;
wire S5255;
wire S5256;
wire S5257;
wire S5258;
wire S5259;
wire S5260;
wire S5261;
wire S5262;
wire S5263;
wire S5264;
wire S5265;
wire S5266;
wire S5267;
wire S5268;
wire S5269;
wire S5270;
wire S5271;
wire S5272;
wire S5273;
wire S5274;
wire S5275;
wire S5276;
wire S5277;
wire S5278;
wire S5279;
wire S5280;
wire S5281;
wire S5282;
wire S5283;
wire S5284;
wire S5285;
wire S5286;
wire S5287;
wire S5288;
wire S5289;
wire S5290;
wire S5291;
wire S5292;
wire S5293;
wire S5294;
wire S5295;
wire S5296;
wire S5297;
wire S5298;
wire S5299;
wire S5300;
wire S5301;
wire S5302;
wire S5303;
wire S5304;
wire S5305;
wire S5306;
wire S5307;
wire S5308;
wire S5309;
wire S5310;
wire S5311;
wire S5312;
wire S5313;
wire S5314;
wire S5315;
wire S5316;
wire S5317;
wire S5318;
wire S5319;
wire S5320;
wire S5321;
wire S5322;
wire S5323;
wire S5324;
wire S5325;
wire S5326;
wire S5327;
wire S5328;
wire S5329;
wire S5330;
wire S5331;
wire S5332;
wire S5333;
wire S5334;
wire S5335;
wire S5336;
wire S5337;
wire S5338;
wire S5339;
wire S5340;
wire S5341;
wire S5342;
wire S5343;
wire S5344;
wire S5345;
wire S5346;
wire S5347;
wire S5348;
wire S5349;
wire S5350;
wire S5351;
wire S5352;
wire S5353;
wire S5354;
wire S5355;
wire S5356;
wire S5357;
wire S5358;
wire S5359;
wire S5360;
wire S5361;
wire S5362;
wire S5363;
wire S5364;
wire S5365;
wire S5366;
wire S5367;
wire S5368;
wire S5369;
wire S5370;
wire S5371;
wire S5372;
wire S5373;
wire S5374;
wire S5375;
wire S5376;
wire S5377;
wire S5378;
wire S5379;
wire S5380;
wire S5381;
wire S5382;
wire S5383;
wire S5384;
wire S5385;
wire S5386;
wire S5387;
wire S5388;
wire S5389;
wire S5390;
wire S5391;
wire S5392;
wire S5393;
wire S5394;
wire S5395;
wire S5396;
wire S5397;
wire S5398;
wire S5399;
wire S5400;
wire S5401;
wire S5402;
wire S5403;
wire S5404;
wire S5405;
wire S5406;
wire S5407;
wire S5408;
wire S5409;
wire S5410;
wire S5411;
wire S5412;
wire S5413;
wire S5414;
wire S5415;
wire S5416;
wire S5417;
wire S5418;
wire S5419;
wire S5420;
wire S5421;
wire S5422;
wire S5423;
wire S5424;
wire S5425;
wire S5426;
wire S5427;
wire S5428;
wire S5429;
wire S5430;
wire S5431;
wire S5432;
wire S5433;
wire S5434;
wire S5435;
wire S5436;
wire S5437;
wire S5438;
wire S5439;
wire S5440;
wire S5441;
wire S5442;
wire S5443;
wire S5444;
wire S5445;
wire S5446;
wire S5447;
wire S5448;
wire S5449;
wire S5450;
wire S5451;
wire S5452;
wire S5453;
wire S5454;
wire S5455;
wire S5456;
wire S5457;
wire S5458;
wire S5459;
wire S5460;
wire S5461;
wire S5462;
wire S5463;
wire S5464;
wire S5465;
wire S5466;
wire S5467;
wire S5468;
wire S5469;
wire S5470;
wire S5471;
wire S5472;
wire S5473;
wire S5474;
wire S5475;
wire S5476;
wire S5477;
wire S5478;
wire S5479;
wire S5480;
wire S5481;
wire S5482;
wire S5483;
wire S5484;
wire S5485;
wire S5486;
wire S5487;
wire S5488;
wire S5489;
wire S5490;
wire S5491;
wire S5492;
wire S5493;
wire S5494;
wire S5495;
wire S5496;
wire S5497;
wire S5498;
wire S5499;
wire S5500;
wire S5501;
wire S5502;
wire S5503;
wire S5504;
wire S5505;
wire S5506;
wire S5507;
wire S5508;
wire S5509;
wire S5510;
wire S5511;
wire S5512;
wire S5513;
wire S5514;
wire S5515;
wire S5516;
wire S5517;
wire S5518;
wire S5519;
wire S5520;
wire S5521;
wire S5522;
wire S5523;
wire S5524;
wire S5525;
wire S5526;
wire S5527;
wire S5528;
wire S5529;
wire S5530;
wire S5531;
wire S5532;
wire S5533;
wire S5534;
wire S5535;
wire S5536;
wire S5537;
wire S5538;
wire S5539;
wire S5540;
wire S5541;
wire S5542;
wire S5543;
wire S5544;
wire S5545;
wire S5546;
wire S5547;
wire S5548;
wire S5549;
wire S5550;
wire S5551;
wire S5552;
wire S5553;
wire S5554;
wire S5555;
wire S5556;
wire S5557;
wire S5558;
wire S5559;
wire S5560;
wire S5561;
wire S5562;
wire S5563;
wire S5564;
wire S5565;
wire S5566;
wire S5567;
wire S5568;
wire S5569;
wire S5570;
wire S5571;
wire S5572;
wire S5573;
wire S5574;
wire S5575;
wire S5576;
wire S5577;
wire S5578;
wire S5579;
wire S5580;
wire S5581;
wire S5582;
wire S5583;
wire S5584;
wire S5585;
wire S5586;
wire S5587;
wire S5588;
wire S5589;
wire S5590;
wire S5591;
wire S5592;
wire S5593;
wire S5594;
wire S5595;
wire S5596;
wire S5597;
wire S5598;
wire S5599;
wire S5600;
wire S5601;
wire S5602;
wire S5603;
wire S5604;
wire S5605;
wire S5606;
wire S5607;
wire S5608;
wire S5609;
wire S5610;
wire S5611;
wire S5612;
wire S5613;
wire S5614;
wire S5615;
wire S5616;
wire S5617;
wire S5618;
wire S5619;
wire S5620;
wire S5621;
wire S5622;
wire S5623;
wire S5624;
wire S5625;
wire S5626;
wire S5627;
wire S5628;
wire S5629;
wire S5630;
wire S5631;
wire S5632;
wire S5633;
wire S5634;
wire S5635;
wire S5636;
wire S5637;
wire S5638;
wire S5639;
wire S5640;
wire S5641;
wire S5642;
wire S5643;
wire S5644;
wire S5645;
wire S5646;
wire S5647;
wire S5648;
wire S5649;
wire S5650;
wire S5651;
wire S5652;
wire S5653;
wire S5654;
wire S5655;
wire S5656;
wire S5657;
wire S5658;
wire S5659;
wire S5660;
wire S5661;
wire S5662;
wire S5663;
wire S5664;
wire S5665;
wire S5666;
wire S5667;
wire S5668;
wire S5669;
wire S5670;
wire S5671;
wire S5672;
wire S5673;
wire S5674;
wire S5675;
wire S5676;
wire S5677;
wire S5678;
wire S5679;
wire S5680;
wire S5681;
wire S5682;
wire S5683;
wire S5684;
wire S5685;
wire S5686;
wire S5687;
wire S5688;
wire S5689;
wire S5690;
wire S5691;
wire S5692;
wire S5693;
wire S5694;
wire S5695;
wire S5696;
wire S5697;
wire S5698;
wire S5699;
wire S5700;
wire S5701;
wire S5702;
wire S5703;
wire S5704;
wire S5705;
wire S5706;
wire S5707;
wire S5708;
wire S5709;
wire S5710;
wire S5711;
wire S5712;
wire S5713;
wire S5714;
wire S5715;
wire S5716;
wire S5717;
wire S5718;
wire S5719;
wire S5720;
wire S5721;
wire S5722;
wire S5723;
wire S5724;
wire S5725;
wire S5726;
wire S5727;
wire S5728;
wire S5729;
wire S5730;
wire S5731;
wire S5732;
wire S5733;
wire S5734;
wire S5735;
wire S5736;
wire S5737;
wire S5738;
wire S5739;
wire S5740;
wire S5741;
wire S5742;
wire S5743;
wire S5744;
wire S5745;
wire S5746;
wire S5747;
wire S5748;
wire S5749;
wire S5750;
wire S5751;
wire S5752;
wire S5753;
wire S5754;
wire S5755;
wire S5756;
wire S5757;
wire S5758;
wire S5759;
wire S5760;
wire S5761;
wire S5762;
wire S5763;
wire S5764;
wire S5765;
wire S5766;
wire S5767;
wire S5768;
wire S5769;
wire S5770;
wire S5771;
wire S5772;
wire S5773;
wire S5774;
wire S5775;
wire S5776;
wire S5777;
wire S5778;
wire S5779;
wire S5780;
wire S5781;
wire S5782;
wire S5783;
wire S5784;
wire S5785;
wire S5786;
wire S5787;
wire S5788;
wire S5789;
wire S5790;
wire S5791;
wire S5792;
wire S5793;
wire S5794;
wire S5795;
wire S5796;
wire S5797;
wire S5798;
wire S5799;
wire S5800;
wire S5801;
wire S5802;
wire S5803;
wire S5804;
wire S5805;
wire S5806;
wire S5807;
wire S5808;
wire S5809;
wire S5810;
wire S5811;
wire S5812;
wire S5813;
wire S5814;
wire S5815;
wire S5816;
wire S5817;
wire S5818;
wire S5819;
wire S5820;
wire S5821;
wire S5822;
wire S5823;
wire S5824;
wire S5825;
wire S5826;
wire S5827;
wire S5828;
wire S5829;
wire S5830;
wire S5831;
wire S5832;
wire S5833;
wire S5834;
wire S5835;
wire S5836;
wire S5837;
wire S5838;
wire S5839;
wire S5840;
wire S5841;
wire S5842;
wire S5843;
wire S5844;
wire S5845;
wire S5846;
wire S5847;
wire S5848;
wire S5849;
wire S5850;
wire S5851;
wire S5852;
wire S5853;
wire S5854;
wire S5855;
wire S5856;
wire S5857;
wire S5858;
wire S5859;
wire S5860;
wire S5861;
wire S5862;
wire S5863;
wire S5864;
wire S5865;
wire S5866;
wire S5867;
wire S5868;
wire S5869;
wire S5870;
wire S5871;
wire S5872;
wire S5873;
wire S5874;
wire S5875;
wire S5876;
wire S5877;
wire S5878;
wire S5879;
wire S5880;
wire S5881;
wire S5882;
wire S5883;
wire S5884;
wire S5885;
wire S5886;
wire S5887;
wire S5888;
wire S5889;
wire S5890;
wire S5891;
wire S5892;
wire S5893;
wire S5894;
wire S5895;
wire S5896;
wire S5897;
wire S5898;
wire S5899;
wire S5900;
wire S5901;
wire S5902;
wire S5903;
wire S5904;
wire S5905;
wire S5906;
wire S5907;
wire S5908;
wire S5909;
wire S5910;
wire S5911;
wire S5912;
wire S5913;
wire S5914;
wire S5915;
wire S5916;
wire S5917;
wire S5918;
wire S5919;
wire S5920;
wire S5921;
wire S5922;
wire S5923;
wire S5924;
wire S5925;
wire S5926;
wire S5927;
wire S5928;
wire S5929;
wire S5930;
wire S5931;
wire S5932;
wire S5933;
wire S5934;
wire S5935;
wire S5936;
wire S5937;
wire S5938;
wire S5939;
wire S5940;
wire S5941;
wire S5942;
wire S5943;
wire S5944;
wire S5945;
wire S5946;
wire S5947;
wire S5948;
wire S5949;
wire S5950;
wire S5951;
wire S5952;
wire S5953;
wire S5954;
wire S5955;
wire S5956;
wire S5957;
wire S5958;
wire S5959;
wire S5960;
wire S5961;
wire S5962;
wire S5963;
wire S5964;
wire S5965;
wire S5966;
wire S5967;
wire S5968;
wire S5969;
wire S5970;
wire S5971;
wire S5972;
wire S5973;
wire S5974;
wire S5975;
wire S5976;
wire S5977;
wire S5978;
wire S5979;
wire S5980;
wire S5981;
wire S5982;
wire S5983;
wire S5984;
wire S5985;
wire S5986;
wire S5987;
wire S5988;
wire S5989;
wire S5990;
wire S5991;
wire S5992;
wire S5993;
wire S5994;
wire S5995;
wire S5996;
wire S5997;
wire S5998;
wire S5999;
wire S6000;
wire S6001;
wire S6002;
wire S6003;
wire S6004;
wire S6005;
wire S6006;
wire S6007;
wire S6008;
wire S6009;
wire S6010;
wire S6011;
wire S6012;
wire S6013;
wire S6014;
wire S6015;
wire S6016;
wire S6017;
wire S6018;
wire S6019;
wire S6020;
wire S6021;
wire S6022;
wire S6023;
wire S6024;
wire S6025;
wire S6026;
wire S6027;
wire S6028;
wire S6029;
wire S6030;
wire S6031;
wire S6032;
wire S6033;
wire S6034;
wire S6035;
wire S6036;
wire S6037;
wire S6038;
wire S6039;
wire S6040;
wire S6041;
wire S6042;
wire S6043;
wire S6044;
wire S6045;
wire S6046;
wire S6047;
wire S6048;
wire S6049;
wire S6050;
wire S6051;
wire S6052;
wire S6053;
wire S6054;
wire S6055;
wire S6056;
wire S6057;
wire S6058;
wire S6059;
wire S6060;
wire S6061;
wire S6062;
wire S6063;
wire S6064;
wire S6065;
wire S6066;
wire S6067;
wire S6068;
wire S6069;
wire S6070;
wire S6071;
wire S6072;
wire S6073;
wire S6074;
wire S6075;
wire S6076;
wire S6077;
wire S6078;
wire S6079;
wire S6080;
wire S6081;
wire S6082;
wire S6083;
wire S6084;
wire S6085;
wire S6086;
wire S6087;
wire S6088;
wire S6089;
wire S6090;
wire S6091;
wire S6092;
wire S6093;
wire S6094;
wire S6095;
wire S6096;
wire S6097;
wire S6098;
wire S6099;
wire S6100;
wire S6101;
wire S6102;
wire S6103;
wire S6104;
wire S6105;
wire S6106;
wire S6107;
wire S6108;
wire S6109;
wire S6110;
wire S6111;
wire S6112;
wire S6113;
wire S6114;
wire S6115;
wire S6116;
wire S6117;
wire S6118;
wire S6119;
wire S6120;
wire S6121;
wire S6122;
wire S6123;
wire S6124;
wire S6125;
wire S6126;
wire S6127;
wire S6128;
wire S6129;
wire S6130;
wire S6131;
wire S6132;
wire S6133;
wire S6134;
wire S6135;
wire S6136;
wire S6137;
wire S6138;
wire S6139;
wire S6140;
wire S6141;
wire S6142;
wire S6143;
wire S6144;
wire S6145;
wire S6146;
wire S6147;
wire S6148;
wire S6149;
wire S6150;
wire S6151;
wire S6152;
wire S6153;
wire S6154;
wire S6155;
wire S6156;
wire S6157;
wire S6158;
wire S6159;
wire S6160;
wire S6161;
wire S6162;
wire S6163;
wire S6164;
wire S6165;
wire S6166;
wire S6167;
wire S6168;
wire S6169;
wire S6170;
wire S6171;
wire S6172;
wire S6173;
wire S6174;
wire S6175;
wire S6176;
wire S6177;
wire S6178;
wire S6179;
wire S6180;
wire S6181;
wire S6182;
wire S6183;
wire S6184;
wire S6185;
wire S6186;
wire S6187;
wire S6188;
wire S6189;
wire S6190;
wire S6191;
wire S6192;
wire S6193;
wire S6194;
wire S6195;
wire S6196;
wire S6197;
wire S6198;
wire S6199;
wire S6200;
wire S6201;
wire S6202;
wire S6203;
wire S6204;
wire S6205;
wire S6206;
wire S6207;
wire S6208;
wire S6209;
wire S6210;
wire S6211;
wire S6212;
wire S6213;
wire S6214;
wire S6215;
wire S6216;
wire S6217;
wire S6218;
wire S6219;
wire S6220;
wire S6221;
wire S6222;
wire S6223;
wire S6224;
wire S6225;
wire S6226;
wire S6227;
wire S6228;
wire S6229;
wire S6230;
wire S6231;
wire S6232;
wire S6233;
wire S6234;
wire S6235;
wire S6236;
wire S6237;
wire S6238;
wire S6239;
wire S6240;
wire S6241;
wire S6242;
wire S6243;
wire S6244;
wire S6245;
wire S6246;
wire S6247;
wire S6248;
wire S6249;
wire S6250;
wire S6251;
wire S6252;
wire S6253;
wire S6254;
wire S6255;
wire S6256;
wire S6257;
wire S6258;
wire S6259;
wire S6260;
wire S6261;
wire S6262;
wire S6263;
wire S6264;
wire S6265;
wire S6266;
wire S6267;
wire S6268;
wire S6269;
wire S6270;
wire S6271;
wire S6272;
wire S6273;
wire S6274;
wire S6275;
wire S6276;
wire S6277;
wire S6278;
wire S6279;
wire S6280;
wire S6281;
wire S6282;
wire S6283;
wire S6284;
wire S6285;
wire S6286;
wire S6287;
wire S6288;
wire S6289;
wire S6290;
wire S6291;
wire S6292;
wire S6293;
wire S6294;
wire S6295;
wire S6296;
wire S6297;
wire S6298;
wire S6299;
wire S6300;
wire S6301;
wire S6302;
wire S6303;
wire S6304;
wire S6305;
wire S6306;
wire S6307;
wire S6308;
wire S6309;
wire S6310;
wire S6311;
wire S6312;
wire S6313;
wire S6314;
wire S6315;
wire S6316;
wire S6317;
wire S6318;
wire S6319;
wire S6320;
wire S6321;
wire S6322;
wire S6323;
wire S6324;
wire S6325;
wire S6326;
wire S6327;
wire S6328;
wire S6329;
wire S6330;
wire S6331;
wire S6332;
wire S6333;
wire S6334;
wire S6335;
wire S6336;
wire S6337;
wire S6338;
wire S6339;
wire S6340;
wire S6341;
wire S6342;
wire S6343;
wire S6344;
wire S6345;
wire S6346;
wire S6347;
wire S6348;
wire S6349;
wire S6350;
wire S6351;
wire S6352;
wire S6353;
wire S6354;
wire S6355;
wire S6356;
wire S6357;
wire S6358;
wire S6359;
wire S6360;
wire S6361;
wire S6362;
wire S6363;
wire S6364;
wire S6365;
wire S6366;
wire S6367;
wire S6368;
wire S6369;
wire S6370;
wire S6371;
wire S6372;
wire S6373;
wire S6374;
wire S6375;
wire S6376;
wire S6377;
wire S6378;
wire S6379;
wire S6380;
wire S6381;
wire S6382;
wire S6383;
wire S6384;
wire S6385;
wire S6386;
wire S6387;
wire S6388;
wire S6389;
wire S6390;
wire S6391;
wire S6392;
wire S6393;
wire S6394;
wire S6395;
wire S6396;
wire S6397;
wire S6398;
wire S6399;
wire S6400;
wire S6401;
wire S6402;
wire S6403;
wire S6404;
wire S6405;
wire S6406;
wire S6407;
wire S6408;
wire S6409;
wire S6410;
wire S6411;
wire S6412;
wire S6413;
wire S6414;
wire S6415;
wire S6416;
wire S6417;
wire S6418;
wire S6419;
wire S6420;
wire S6421;
wire S6422;
wire S6423;
wire S6424;
wire S6425;
wire S6426;
wire S6427;
wire S6428;
wire S6429;
wire S6430;
wire S6431;
wire S6432;
wire S6433;
wire S6434;
wire S6435;
wire S6436;
wire S6437;
wire S6438;
wire S6439;
wire S6440;
wire S6441;
wire S6442;
wire S6443;
wire S6444;
wire S6445;
wire S6446;
wire S6447;
wire S6448;
wire S6449;
wire S6450;
wire S6451;
wire S6452;
wire S6453;
wire S6454;
wire S6455;
wire S6456;
wire S6457;
wire S6458;
wire S6459;
wire S6460;
wire S6461;
wire S6462;
wire S6463;
wire S6464;
wire S6465;
wire S6466;
wire S6467;
wire S6468;
wire S6469;
wire S6470;
wire S6471;
wire S6472;
wire S6473;
wire S6474;
wire S6475;
wire S6476;
wire S6477;
wire S6478;
wire S6479;
wire S6480;
wire S6481;
wire S6482;
wire S6483;
wire S6484;
wire S6485;
wire S6486;
wire S6487;
wire S6488;
wire S6489;
wire S6490;
wire S6491;
wire S6492;
wire S6493;
wire S6494;
wire S6495;
wire S6496;
wire S6497;
wire S6498;
wire S6499;
wire S6500;
wire S6501;
wire S6502;
wire S6503;
wire S6504;
wire S6505;
wire S6506;
wire S6507;
wire S6508;
wire S6509;
wire S6510;
wire S6511;
wire S6512;
wire S6513;
wire S6514;
wire S6515;
wire S6516;
wire S6517;
wire S6518;
wire S6519;
wire S6520;
wire S6521;
wire S6522;
wire S6523;
wire S6524;
wire S6525;
wire S6526;
wire S6527;
wire S6528;
wire S6529;
wire S6530;
wire S6531;
wire S6532;
wire S6533;
wire S6534;
wire S6535;
wire S6536;
wire S6537;
wire S6538;
wire S6539;
wire S6540;
wire S6541;
wire S6542;
wire S6543;
wire S6544;
wire S6545;
wire S6546;
wire S6547;
wire S6548;
wire S6549;
wire S6550;
wire S6551;
wire S6552;
wire S6553;
wire S6554;
wire S6555;
wire S6556;
wire S6557;
wire S6558;
wire S6559;
wire S6560;
wire S6561;
wire S6562;
wire S6563;
wire S6564;
wire S6565;
wire S6566;
wire S6567;
wire S6568;
wire S6569;
wire S6570;
wire S6571;
wire S6572;
wire S6573;
wire S6574;
wire S6575;
wire S6576;
wire S6577;
wire S6578;
wire S6579;
wire S6580;
wire S6581;
wire S6582;
wire S6583;
wire S6584;
wire S6585;
wire S6586;
wire S6587;
wire S6588;
wire S6589;
wire S6590;
wire S6591;
wire S6592;
wire S6593;
wire S6594;
wire S6595;
wire S6596;
wire S6597;
wire S6598;
wire S6599;
wire S6600;
wire S6601;
wire S6602;
wire S6603;
wire S6604;
wire S6605;
wire S6606;
wire S6607;
wire S6608;
wire S6609;
wire S6610;
wire S6611;
wire S6612;
wire S6613;
wire S6614;
wire S6615;
wire S6616;
wire S6617;
wire S6618;
wire S6619;
wire S6620;
wire S6621;
wire S6622;
wire S6623;
wire S6624;
wire S6625;
wire S6626;
wire S6627;
wire S6628;
wire S6629;
wire S6630;
wire S6631;
wire S6632;
wire S6633;
wire S6634;
wire S6635;
wire S6636;
wire S6637;
wire S6638;
wire S6639;
wire S6640;
wire S6641;
wire S6642;
wire S6643;
wire S6644;
wire S6645;
wire S6646;
wire S6647;
wire S6648;
wire S6649;
wire S6650;
wire S6651;
wire S6652;
wire S6653;
wire S6654;
wire S6655;
wire S6656;
wire S6657;
wire S6658;
wire S6659;
wire S6660;
wire S6661;
wire S6662;
wire S6663;
wire S6664;
wire S6665;
wire S6666;
wire S6667;
wire S6668;
wire S6669;
wire S6670;
wire S6671;
wire S6672;
wire S6673;
wire S6674;
wire S6675;
wire S6676;
wire S6677;
wire S6678;
wire S6679;
wire S6680;
wire S6681;
wire S6682;
wire S6683;
wire S6684;
wire S6685;
wire S6686;
wire S6687;
wire S6688;
wire S6689;
wire S6690;
wire S6691;
wire S6692;
wire S6693;
wire S6694;
wire S6695;
wire S6696;
wire S6697;
wire S6698;
wire S6699;
wire S6700;
wire S6701;
wire S6702;
wire S6703;
wire S6704;
wire S6705;
wire S6706;
wire S6707;
wire S6708;
wire S6709;
wire S6710;
wire S6711;
wire S6712;
wire S6713;
wire S6714;
wire S6715;
wire S6716;
wire S6717;
wire S6718;
wire S6719;
wire S6720;
wire S6721;
wire S6722;
wire S6723;
wire S6724;
wire S6725;
wire S6726;
wire S6727;
wire S6728;
wire S6729;
wire S6730;
wire S6731;
wire S6732;
wire S6733;
wire S6734;
wire S6735;
wire S6736;
wire S6737;
wire S6738;
wire S6739;
wire S6740;
wire S6741;
wire S6742;
wire S6743;
wire S6744;
wire S6745;
wire S6746;
wire S6747;
wire S6748;
wire S6749;
wire S6750;
wire S6751;
wire S6752;
wire S6753;
wire S6754;
wire S6755;
wire S6756;
wire S6757;
wire S6758;
wire S6759;
wire S6760;
wire S6761;
wire S6762;
wire S6763;
wire S6764;
wire S6765;
wire S6766;
wire S6767;
wire S6768;
wire S6769;
wire S6770;
wire S6771;
wire S6772;
wire S6773;
wire S6774;
wire S6775;
wire S6776;
wire S6777;
wire S6778;
wire S6779;
wire S6780;
wire S6781;
wire S6782;
wire S6783;
wire S6784;
wire S6785;
wire S6786;
wire S6787;
wire S6788;
wire S6789;
wire S6790;
wire S6791;
wire S6792;
wire S6793;
wire S6794;
wire S6795;
wire S6796;
wire S6797;
wire S6798;
wire S6799;
wire S6800;
wire S6801;
wire S6802;
wire S6803;
wire S6804;
wire S6805;
wire S6806;
wire S6807;
wire S6808;
wire S6809;
wire S6810;
wire S6811;
wire S6812;
wire S6813;
wire S6814;
wire S6815;
wire S6816;
wire S6817;
wire S6818;
wire S6819;
wire S6820;
wire S6821;
wire S6822;
wire S6823;
wire S6824;
wire S6825;
wire S6826;
wire S6827;
wire S6828;
wire S6829;
wire S6830;
wire S6831;
wire S6832;
wire S6833;
wire S6834;
wire S6835;
wire S6836;
wire S6837;
wire S6838;
wire S6839;
wire S6840;
wire S6841;
wire S6842;
wire S6843;
wire S6844;
wire S6845;
wire S6846;
wire S6847;
wire S6848;
wire S6849;
wire S6850;
wire S6851;
wire S6852;
wire S6853;
wire S6854;
wire S6855;
wire S6856;
wire S6857;
wire S6858;
wire S6859;
wire S6860;
wire S6861;
wire S6862;
wire S6863;
wire S6864;
wire S6865;
wire S6866;
wire S6867;
wire S6868;
wire S6869;
wire S6870;
wire S6871;
wire S6872;
wire S6873;
wire S6874;
wire S6875;
wire S6876;
wire S6877;
wire S6878;
wire S6879;
wire S6880;
wire S6881;
wire S6882;
wire S6883;
wire S6884;
wire S6885;
wire S6886;
wire S6887;
wire S6888;
wire S6889;
wire S6890;
wire S6891;
wire S6892;
wire S6893;
wire S6894;
wire S6895;
wire S6896;
wire S6897;
wire S6898;
wire S6899;
wire S6900;
wire S6901;
wire S6902;
wire S6903;
wire S6904;
wire S6905;
wire S6906;
wire S6907;
wire S6908;
wire S6909;
wire S6910;
wire S6911;
wire S6912;
wire S6913;
wire S6914;
wire S6915;
wire S6916;
wire S6917;
wire S6918;
wire S6919;
wire S6920;
wire S6921;
wire S6922;
wire S6923;
wire S6924;
wire S6925;
wire S6926;
wire S6927;
wire S6928;
wire S6929;
wire S6930;
wire S6931;
wire S6932;
wire S6933;
wire S6934;
wire S6935;
wire S6936;
wire S6937;
wire S6938;
wire S6939;
wire S6940;
wire S6941;
wire S6942;
wire S6943;
wire S6944;
wire S6945;
wire S6946;
wire S6947;
wire S6948;
wire S6949;
wire S6950;
wire S6951;
wire S6952;
wire S6953;
wire S6954;
wire S6955;
wire S6956;
wire S6957;
wire S6958;
wire S6959;
wire S6960;
wire S6961;
wire S6962;
wire S6963;
wire S6964;
wire S6965;
wire S6966;
wire S6967;
wire S6968;
wire S6969;
wire S6970;
wire S6971;
wire S6972;
wire S6973;
wire S6974;
wire S6975;
wire S6976;
wire S6977;
wire S6978;
wire S6979;
wire S6980;
wire S6981;
wire S6982;
wire S6983;
wire S6984;
wire S6985;
wire S6986;
wire S6987;
wire S6988;
wire S6989;
wire S6990;
wire S6991;
wire S6992;
wire S6993;
wire S6994;
wire S6995;
wire S6996;
wire S6997;
wire S6998;
wire S6999;
wire S7000;
wire S7001;
wire S7002;
wire S7003;
wire S7004;
wire S7005;
wire S7006;
wire S7007;
wire S7008;
wire S7009;
wire S7010;
wire S7011;
wire S7012;
wire S7013;
wire S7014;
wire S7015;
wire S7016;
wire S7017;
wire S7018;
wire S7019;
wire S7020;
wire S7021;
wire S7022;
wire S7023;
wire S7024;
wire S7025;
wire S7026;
wire S7027;
wire S7028;
wire S7029;
wire S7030;
wire S7031;
wire S7032;
wire S7033;
wire S7034;
wire S7035;
wire S7036;
wire S7037;
wire S7038;
wire S7039;
wire S7040;
wire S7041;
wire S7042;
wire S7043;
wire S7044;
wire S7045;
wire S7046;
wire S7047;
wire S7048;
wire S7049;
wire S7050;
wire S7051;
wire S7052;
wire S7053;
wire S7054;
wire S7055;
wire S7056;
wire S7057;
wire S7058;
wire S7059;
wire S7060;
wire S7061;
wire S7062;
wire S7063;
wire S7064;
wire S7065;
wire S7066;
wire S7067;
wire S7068;
wire S7069;
wire S7070;
wire S7071;
wire S7072;
wire S7073;
wire S7074;
wire S7075;
wire S7076;
wire S7077;
wire S7078;
wire S7079;
wire S7080;
wire S7081;
wire S7082;
wire S7083;
wire S7084;
wire S7085;
wire S7086;
wire S7087;
wire S7088;
wire S7089;
wire S7090;
wire S7091;
wire S7092;
wire S7093;
wire S7094;
wire S7095;
wire S7096;
wire S7097;
wire S7098;
wire S7099;
wire S7100;
wire S7101;
wire S7102;
wire S7103;
wire S7104;
wire S7105;
wire S7106;
wire S7107;
wire S7108;
wire S7109;
wire S7110;
wire S7111;
wire S7112;
wire S7113;
wire S7114;
wire S7115;
wire S7116;
wire S7117;
wire S7118;
wire S7119;
wire S7120;
wire S7121;
wire S7122;
wire S7123;
wire S7124;
wire S7125;
wire S7126;
wire S7127;
wire S7128;
wire S7129;
wire S7130;
wire S7131;
wire S7132;
wire S7133;
wire S7134;
wire S7135;
wire S7136;
wire S7137;
wire S7138;
wire S7139;
wire S7140;
wire S7141;
wire S7142;
wire S7143;
wire S7144;
wire S7145;
wire S7146;
wire S7147;
wire S7148;
wire S7149;
wire S7150;
wire S7151;
wire S7152;
wire S7153;
wire S7154;
wire S7155;
wire S7156;
wire S7157;
wire S7158;
wire S7159;
wire S7160;
wire S7161;
wire S7162;
wire S7163;
wire S7164;
wire S7165;
wire S7166;
wire S7167;
wire S7168;
wire S7169;
wire S7170;
wire S7171;
wire S7172;
wire S7173;
wire S7174;
wire S7175;
wire S7176;
wire S7177;
wire S7178;
wire S7179;
wire S7180;
wire S7181;
wire S7182;
wire S7183;
wire S7184;
wire S7185;
wire S7186;
wire S7187;
wire S7188;
wire S7189;
wire S7190;
wire S7191;
wire S7192;
wire S7193;
wire S7194;
wire S7195;
wire S7196;
wire S7197;
wire S7198;
wire S7199;
wire S7200;
wire S7201;
wire S7202;
wire S7203;
wire S7204;
wire S7205;
wire S7206;
wire S7207;
wire S7208;
wire S7209;
wire S7210;
wire S7211;
wire S7212;
wire S7213;
wire S7214;
wire S7215;
wire S7216;
wire S7217;
wire S7218;
wire S7219;
wire S7220;
wire S7221;
wire S7222;
wire S7223;
wire S7224;
wire S7225;
wire S7226;
wire S7227;
wire S7228;
wire S7229;
wire S7230;
wire S7231;
wire S7232;
wire S7233;
wire S7234;
wire S7235;
wire S7236;
wire S7237;
wire S7238;
wire S7239;
wire S7240;
wire S7241;
wire S7242;
wire S7243;
wire S7244;
wire S7245;
wire S7246;
wire S7247;
wire S7248;
wire S7249;
wire S7250;
wire S7251;
wire S7252;
wire S7253;
wire S7254;
wire S7255;
wire S7256;
wire S7257;
wire S7258;
wire S7259;
wire S7260;
wire S7261;
wire S7262;
wire S7263;
wire S7264;
wire S7265;
wire S7266;
wire S7267;
wire S7268;
wire S7269;
wire S7270;
wire S7271;
wire S7272;
wire S7273;
wire S7274;
wire S7275;
wire S7276;
wire S7277;
wire S7278;
wire S7279;
wire S7280;
wire S7281;
wire S7282;
wire S7283;
wire S7284;
wire S7285;
wire S7286;
wire S7287;
wire S7288;
wire S7289;
wire S7290;
wire S7291;
wire S7292;
wire S7293;
wire S7294;
wire S7295;
wire S7296;
wire S7297;
wire S7298;
wire S7299;
wire S7300;
wire S7301;
wire S7302;
wire S7303;
wire S7304;
wire S7305;
wire S7306;
wire S7307;
wire S7308;
wire S7309;
wire S7310;
wire S7311;
wire S7312;
wire S7313;
wire S7314;
wire S7315;
wire S7316;
wire S7317;
wire S7318;
wire S7319;
wire S7320;
wire S7321;
wire S7322;
wire S7323;
wire S7324;
wire S7325;
wire S7326;
wire S7327;
wire S7328;
wire S7329;
wire S7330;
wire S7331;
wire S7332;
wire S7333;
wire S7334;
wire S7335;
wire S7336;
wire S7337;
wire S7338;
wire S7339;
wire S7340;
wire S7341;
wire S7342;
wire S7343;
wire S7344;
wire S7345;
wire S7346;
wire S7347;
wire S7348;
wire S7349;
wire S7350;
wire S7351;
wire S7352;
wire S7353;
wire S7354;
wire S7355;
wire S7356;
wire S7357;
wire S7358;
wire S7359;
wire S7360;
wire S7361;
wire S7362;
wire S7363;
wire S7364;
wire S7365;
wire S7366;
wire S7367;
wire S7368;
wire S7369;
wire S7370;
wire S7371;
wire S7372;
wire S7373;
wire S7374;
wire S7375;
wire S7376;
wire S7377;
wire S7378;
wire S7379;
wire S7380;
wire S7381;
wire S7382;
wire S7383;
wire S7384;
wire S7385;
wire S7386;
wire S7387;
wire S7388;
wire S7389;
wire S7390;
wire S7391;
wire S7392;
wire S7393;
wire S7394;
wire S7395;
wire S7396;
wire S7397;
wire S7398;
wire S7399;
wire S7400;
wire S7401;
wire S7402;
wire S7403;
wire S7404;
wire S7405;
wire S7406;
wire S7407;
wire S7408;
wire S7409;
wire S7410;
wire S7411;
wire S7412;
wire S7413;
wire S7414;
wire S7415;
wire S7416;
wire S7417;
wire S7418;
wire S7419;
wire S7420;
wire S7421;
wire S7422;
wire S7423;
wire S7424;
wire S7425;
wire S7426;
wire S7427;
wire S7428;
wire S7429;
wire S7430;
wire S7431;
wire S7432;
wire S7433;
wire S7434;
wire S7435;
wire S7436;
wire S7437;
wire S7438;
wire S7439;
wire S7440;
wire S7441;
wire S7442;
wire S7443;
wire S7444;
wire S7445;
wire S7446;
wire S7447;
wire S7448;
wire S7449;
wire S7450;
wire S7451;
wire S7452;
wire S7453;
wire S7454;
wire S7455;
wire S7456;
wire S7457;
wire S7458;
wire S7459;
wire S7460;
wire S7461;
wire S7462;
wire S7463;
wire S7464;
wire S7465;
wire S7466;
wire S7467;
wire S7468;
wire S7469;
wire S7470;
wire S7471;
wire S7472;
wire S7473;
wire S7474;
wire S7475;
wire S7476;
wire S7477;
wire S7478;
wire S7479;
wire S7480;
wire S7481;
wire S7482;
wire S7483;
wire S7484;
wire S7485;
wire S7486;
wire S7487;
wire S7488;
wire S7489;
wire S7490;
wire S7491;
wire S7492;
wire S7493;
wire S7494;
wire S7495;
wire S7496;
wire S7497;
wire S7498;
wire S7499;
wire S7500;
wire S7501;
wire S7502;
wire S7503;
wire S7504;
wire S7505;
wire S7506;
wire S7507;
wire S7508;
wire S7509;
wire S7510;
wire S7511;
wire S7512;
wire S7513;
wire S7514;
wire S7515;
wire S7516;
wire S7517;
wire S7518;
wire S7519;
wire S7520;
wire S7521;
wire S7522;
wire S7523;
wire S7524;
wire S7525;
wire S7526;
wire S7527;
wire S7528;
wire S7529;
wire S7530;
wire S7531;
wire S7532;
wire S7533;
wire S7534;
wire S7535;
wire S7536;
wire S7537;
wire S7538;
wire S7539;
wire S7540;
wire S7541;
wire S7542;
wire S7543;
wire S7544;
wire S7545;
wire S7546;
wire S7547;
wire S7548;
wire S7549;
wire S7550;
wire S7551;
wire S7552;
wire S7553;
wire S7554;
wire S7555;
wire S7556;
wire S7557;
wire S7558;
wire S7559;
wire S7560;
wire S7561;
wire S7562;
wire S7563;
wire S7564;
wire S7565;
wire S7566;
wire S7567;
wire S7568;
wire S7569;
wire S7570;
wire S7571;
wire S7572;
wire S7573;
wire S7574;
wire S7575;
wire S7576;
wire S7577;
wire S7578;
wire S7579;
wire S7580;
wire S7581;
wire S7582;
wire S7583;
wire S7584;
wire S7585;
wire S7586;
wire S7587;
wire S7588;
wire S7589;
wire S7590;
wire S7591;
wire S7592;
wire S7593;
wire S7594;
wire S7595;
wire S7596;
wire S7597;
wire S7598;
wire S7599;
wire S7600;
wire S7601;
wire S7602;
wire S7603;
wire S7604;
wire S7605;
wire S7606;
wire S7607;
wire S7608;
wire S7609;
wire S7610;
wire S7611;
wire S7612;
wire S7613;
wire S7614;
wire S7615;
wire S7616;
wire S7617;
wire S7618;
wire S7619;
wire S7620;
wire S7621;
wire S7622;
wire S7623;
wire S7624;
wire S7625;
wire S7626;
wire S7627;
wire S7628;
wire S7629;
wire S7630;
wire S7631;
wire S7632;
wire S7633;
wire S7634;
wire S7635;
wire S7636;
wire S7637;
wire S7638;
wire S7639;
wire S7640;
wire S7641;
wire S7642;
wire S7643;
wire S7644;
wire S7645;
wire S7646;
wire S7647;
wire S7648;
wire S7649;
wire S7650;
wire S7651;
wire S7652;
wire S7653;
wire S7654;
wire S7655;
wire S7656;
wire S7657;
wire S7658;
wire S7659;
wire S7660;
wire S7661;
wire S7662;
wire S7663;
wire S7664;
wire S7665;
wire S7666;
wire S7667;
wire S7668;
wire S7669;
wire S7670;
wire S7671;
wire S7672;
wire S7673;
wire S7674;
wire S7675;
wire S7676;
wire S7677;
wire S7678;
wire S7679;
wire S7680;
wire S7681;
wire S7682;
wire S7683;
wire S7684;
wire S7685;
wire S7686;
wire S7687;
wire S7688;
wire S7689;
wire S7690;
wire S7691;
wire S7692;
wire S7693;
wire S7694;
wire S7695;
wire S7696;
wire S7697;
wire S7698;
wire S7699;
wire S7700;
wire S7701;
wire S7702;
wire S7703;
wire S7704;
wire S7705;
wire S7706;
wire S7707;
wire S7708;
wire S7709;
wire S7710;
wire S7711;
wire S7712;
wire S7713;
wire S7714;
wire S7715;
wire S7716;
wire S7717;
wire S7718;
wire S7719;
wire S7720;
wire S7721;
wire S7722;
wire S7723;
wire S7724;
wire S7725;
wire S7726;
wire S7727;
wire S7728;
wire S7729;
wire S7730;
wire S7731;
wire S7732;
wire S7733;
wire S7734;
wire S7735;
wire S7736;
wire S7737;
wire S7738;
wire S7739;
wire S7740;
wire S7741;
wire S7742;
wire S7743;
wire S7744;
wire S7745;
wire S7746;
wire S7747;
wire S7748;
wire S7749;
wire S7750;
wire S7751;
wire S7752;
wire S7753;
wire S7754;
wire S7755;
wire S7756;
wire S7757;
wire S7758;
wire S7759;
wire S7760;
wire S7761;
wire S7762;
wire S7763;
wire S7764;
wire S7765;
wire S7766;
wire S7767;
wire S7768;
wire S7769;
wire S7770;
wire S7771;
wire S7772;
wire S7773;
wire S7774;
wire S7775;
wire S7776;
wire S7777;
wire S7778;
wire S7779;
wire S7780;
wire S7781;
wire S7782;
wire S7783;
wire S7784;
wire S7785;
wire S7786;
wire S7787;
wire S7788;
wire S7789;
wire S7790;
wire S7791;
wire S7792;
wire S7793;
wire S7794;
wire S7795;
wire S7796;
wire S7797;
wire S7798;
wire S7799;
wire S7800;
wire S7801;
wire S7802;
wire S7803;
wire S7804;
wire S7805;
wire S7806;
wire S7807;
wire S7808;
wire S7809;
wire S7810;
wire S7811;
wire S7812;
wire S7813;
wire S7814;
wire S7815;
wire S7816;
wire S7817;
wire S7818;
wire S7819;
wire S7820;
wire S7821;
wire S7822;
wire S7823;
wire S7824;
wire S7825;
wire S7826;
wire S7827;
wire S7828;
wire S7829;
wire S7830;
wire S7831;
wire S7832;
wire S7833;
wire S7834;
wire S7835;
wire S7836;
wire S7837;
wire S7838;
wire S7839;
wire S7840;
wire S7841;
wire S7842;
wire S7843;
wire S7844;
wire S7845;
wire S7846;
wire S7847;
wire S7848;
wire S7849;
wire S7850;
wire S7851;
wire S7852;
wire S7853;
wire S7854;
wire S7855;
wire S7856;
wire S7857;
wire S7858;
wire S7859;
wire S7860;
wire S7861;
wire S7862;
wire S7863;
wire S7864;
wire S7865;
wire S7866;
wire S7867;
wire S7868;
wire S7869;
wire S7870;
wire S7871;
wire S7872;
wire S7873;
wire S7874;
wire S7875;
wire S7876;
wire S7877;
wire S7878;
wire S7879;
wire S7880;
wire S7881;
wire S7882;
wire S7883;
wire S7884;
wire S7885;
wire S7886;
wire S7887;
wire S7888;
wire S7889;
wire S7890;
wire S7891;
wire S7892;
wire S7893;
wire S7894;
wire S7895;
wire S7896;
wire S7897;
wire S7898;
wire S7899;
wire S7900;
wire S7901;
wire S7902;
wire S7903;
wire S7904;
wire S7905;
wire S7906;
wire S7907;
wire S7908;
wire S7909;
wire S7910;
wire S7911;
wire S7912;
wire S7913;
wire S7914;
wire S7915;
wire S7916;
wire S7917;
wire S7918;
wire S7919;
wire S7920;
wire S7921;
wire S7922;
wire S7923;
wire S7924;
wire S7925;
wire S7926;
wire S7927;
wire S7928;
wire S7929;
wire S7930;
wire S7931;
wire S7932;
wire S7933;
wire S7934;
wire S7935;
wire S7936;
wire S7937;
wire S7938;
wire S7939;
wire S7940;
wire S7941;
wire S7942;
wire S7943;
wire S7944;
wire S7945;
wire S7946;
wire S7947;
wire S7948;
wire S7949;
wire S7950;
wire S7951;
wire S7952;
wire S7953;
wire S7954;
wire S7955;
wire S7956;
wire S7957;
wire S7958;
wire S7959;
wire S7960;
wire S7961;
wire S7962;
wire S7963;
wire S7964;
wire S7965;
wire S7966;
wire S7967;
wire S7968;
wire S7969;
wire S7970;
wire S7971;
wire S7972;
wire S7973;
wire S7974;
wire S7975;
wire S7976;
wire S7977;
wire S7978;
wire S7979;
wire S7980;
wire S7981;
wire S7982;
wire S7983;
wire S7984;
wire S7985;
wire S7986;
wire S7987;
wire S7988;
wire S7989;
wire S7990;
wire S7991;
wire S7992;
wire S7993;
wire S7994;
wire S7995;
wire S7996;
wire S7997;
wire S7998;
wire S7999;
wire S8000;
wire S8001;
wire S8002;
wire S8003;
wire S8004;
wire S8005;
wire S8006;
wire S8007;
wire S8008;
wire S8009;
wire S8010;
wire S8011;
wire S8012;
wire S8013;
wire S8014;
wire S8015;
wire S8016;
wire S8017;
wire S8018;
wire S8019;
wire S8020;
wire S8021;
wire S8022;
wire S8023;
wire S8024;
wire S8025;
wire S8026;
wire S8027;
wire S8028;
wire S8029;
wire S8030;
wire S8031;
wire S8032;
wire S8033;
wire S8034;
wire S8035;
wire S8036;
wire S8037;
wire S8038;
wire S8039;
wire S8040;
wire S8041;
wire S8042;
wire S8043;
wire S8044;
wire S8045;
wire S8046;
wire S8047;
wire S8048;
wire S8049;
wire S8050;
wire S8051;
wire S8052;
wire S8053;
wire S8054;
wire S8055;
wire S8056;
wire S8057;
wire S8058;
wire S8059;
wire S8060;
wire S8061;
wire S8062;
wire S8063;
wire S8064;
wire S8065;
wire S8066;
wire S8067;
wire S8068;
wire S8069;
wire S8070;
wire S8071;
wire S8072;
wire S8073;
wire S8074;
wire S8075;
wire S8076;
wire S8077;
wire S8078;
wire S8079;
wire S8080;
wire S8081;
wire S8082;
wire S8083;
wire S8084;
wire S8085;
wire S8086;
wire S8087;
wire S8088;
wire S8089;
wire S8090;
wire S8091;
wire S8092;
wire S8093;
wire S8094;
wire S8095;
wire S8096;
wire S8097;
wire S8098;
wire S8099;
wire S8100;
wire S8101;
wire S8102;
wire S8103;
wire S8104;
wire S8105;
wire S8106;
wire S8107;
wire S8108;
wire S8109;
wire S8110;
wire S8111;
wire S8112;
wire S8113;
wire S8114;
wire S8115;
wire S8116;
wire S8117;
wire S8118;
wire S8119;
wire S8120;
wire S8121;
wire S8122;
wire S8123;
wire S8124;
wire S8125;
wire S8126;
wire S8127;
wire S8128;
wire S8129;
wire S8130;
wire S8131;
wire S8132;
wire S8133;
wire S8134;
wire S8135;
wire S8136;
wire S8137;
wire S8138;
wire S8139;
wire S8140;
wire S8141;
wire S8142;
wire S8143;
wire S8144;
wire S8145;
wire S8146;
wire S8147;
wire S8148;
wire S8149;
wire S8150;
wire S8151;
wire S8152;
wire S8153;
wire S8154;
wire S8155;
wire S8156;
wire S8157;
wire S8158;
wire S8159;
wire S8160;
wire S8161;
wire S8162;
wire S8163;
wire S8164;
wire S8165;
wire S8166;
wire S8167;
wire S8168;
wire S8169;
wire S8170;
wire S8171;
wire S8172;
wire S8173;
wire S8174;
wire S8175;
wire S8176;
wire S8177;
wire S8178;
wire S8179;
wire S8180;
wire S8181;
wire S8182;
wire S8183;
wire S8184;
wire S8185;
wire S8186;
wire S8187;
wire S8188;
wire S8189;
wire S8190;
wire S8191;
wire S8192;
wire S8193;
wire S8194;
wire S8195;
wire S8196;
wire S8197;
wire S8198;
wire S8199;
wire S8200;
wire S8201;
wire S8202;
wire S8203;
wire S8204;
wire S8205;
wire S8206;
wire S8207;
wire S8208;
wire S8209;
wire S8210;
wire S8211;
wire S8212;
wire S8213;
wire S8214;
wire S8215;
wire S8216;
wire S8217;
wire S8218;
wire S8219;
wire S8220;
wire S8221;
wire S8222;
wire S8223;
wire S8224;
wire S8225;
wire S8226;
wire S8227;
wire S8228;
wire S8229;
wire S8230;
wire S8231;
wire S8232;
wire S8233;
wire S8234;
wire S8235;
wire S8236;
wire S8237;
wire S8238;
wire S8239;
wire S8240;
wire S8241;
wire S8242;
wire S8243;
wire S8244;
wire S8245;
wire S8246;
wire S8247;
wire S8248;
wire S8249;
wire S8250;
wire S8251;
wire S8252;
wire S8253;
wire S8254;
wire S8255;
wire S8256;
wire S8257;
wire S8258;
wire S8259;
wire S8260;
wire S8261;
wire S8262;
wire S8263;
wire S8264;
wire S8265;
wire S8266;
wire S8267;
wire S8268;
wire S8269;
wire S8270;
wire S8271;
wire S8272;
wire S8273;
wire S8274;
wire S8275;
wire S8276;
wire S8277;
wire S8278;
wire S8279;
wire S8280;
wire S8281;
wire S8282;
wire S8283;
wire S8284;
wire S8285;
wire S8286;
wire S8287;
wire S8288;
wire S8289;
wire S8290;
wire S8291;
wire S8292;
wire S8293;
wire S8294;
wire S8295;
wire S8296;
wire S8297;
wire S8298;
wire S8299;
wire S8300;
wire S8301;
wire S8302;
wire S8303;
wire S8304;
wire S8305;
wire S8306;
wire S8307;
wire S8308;
wire S8309;
wire S8310;
wire S8311;
wire S8312;
wire S8313;
wire S8314;
wire S8315;
wire S8316;
wire S8317;
wire S8318;
wire S8319;
wire S8320;
wire S8321;
wire S8322;
wire S8323;
wire S8324;
wire S8325;
wire S8326;
wire S8327;
wire S8328;
wire S8329;
wire S8330;
wire S8331;
wire S8332;
wire S8333;
wire S8334;
wire S8335;
wire S8336;
wire S8337;
wire S8338;
wire S8339;
wire S8340;
wire S8341;
wire S8342;
wire S8343;
wire S8344;
wire S8345;
wire S8346;
wire S8347;
wire S8348;
wire S8349;
wire S8350;
wire S8351;
wire S8352;
wire S8353;
wire S8354;
wire S8355;
wire S8356;
wire S8357;
wire S8358;
wire S8359;
wire S8360;
wire S8361;
wire S8362;
wire S8363;
wire S8364;
wire S8365;
wire S8366;
wire S8367;
wire S8368;
wire S8369;
wire S8370;
wire S8371;
wire S8372;
wire S8373;
wire S8374;
wire S8375;
wire S8376;
wire S8377;
wire S8378;
wire S8379;
wire S8380;
wire S8381;
wire S8382;
wire S8383;
wire S8384;
wire S8385;
wire S8386;
wire S8387;
wire S8388;
wire S8389;
wire S8390;
wire S8391;
wire S8392;
wire S8393;
wire S8394;
wire S8395;
wire S8396;
wire S8397;
wire S8398;
wire S8399;
wire S8400;
wire S8401;
wire S8402;
wire S8403;
wire S8404;
wire S8405;
wire S8406;
wire S8407;
wire S8408;
wire S8409;
wire S8410;
wire S8411;
wire S8412;
wire S8413;
wire S8414;
wire S8415;
wire S8416;
wire S8417;
wire S8418;
wire S8419;
wire S8420;
wire S8421;
wire S8422;
wire S8423;
wire S8424;
wire S8425;
wire S8426;
wire S8427;
wire S8428;
wire S8429;
wire S8430;
wire S8431;
wire S8432;
wire S8433;
wire S8434;
wire S8435;
wire S8436;
wire S8437;
wire S8438;
wire S8439;
wire S8440;
wire S8441;
wire S8442;
wire S8443;
wire S8444;
wire S8445;
wire S8446;
wire S8447;
wire S8448;
wire S8449;
wire S8450;
wire S8451;
wire S8452;
wire S8453;
wire S8454;
wire S8455;
wire S8456;
wire S8457;
wire S8458;
wire S8459;
wire S8460;
wire S8461;
wire S8462;
wire S8463;
wire S8464;
wire S8465;
wire S8466;
wire S8467;
wire S8468;
wire S8469;
wire S8470;
wire S8471;
wire S8472;
wire S8473;
wire S8474;
wire S8475;
wire S8476;
wire S8477;
wire S8478;
wire S8479;
wire S8480;
wire S8481;
wire S8482;
wire S8483;
wire S8484;
wire S8485;
wire S8486;
wire S8487;
wire S8488;
wire S8489;
wire S8490;
wire S8491;
wire S8492;
wire S8493;
wire S8494;
wire S8495;
wire S8496;
wire S8497;
wire S8498;
wire S8499;
wire S8500;
wire S8501;
wire S8502;
wire S8503;
wire S8504;
wire S8505;
wire S8506;
wire S8507;
wire S8508;
wire S8509;
wire S8510;
wire S8511;
wire S8512;
wire S8513;
wire S8514;
wire S8515;
wire S8516;
wire S8517;
wire S8518;
wire S8519;
wire S8520;
wire S8521;
wire S8522;
wire S8523;
wire S8524;
wire S8525;
wire S8526;
wire S8527;
wire S8528;
wire S8529;
wire S8530;
wire S8531;
wire S8532;
wire S8533;
wire S8534;
wire S8535;
wire S8536;
wire S8537;
wire S8538;
wire S8539;
wire S8540;
wire S8541;
wire S8542;
wire S8543;
wire S8544;
wire S8545;
wire S8546;
wire S8547;
wire S8548;
wire S8549;
wire S8550;
wire S8551;
wire S8552;
wire S8553;
wire S8554;
wire S8555;
wire S8556;
wire S8557;
wire S8558;
wire S8559;
wire S8560;
wire S8561;
wire S8562;
wire S8563;
wire S8564;
wire S8565;
wire S8566;
wire S8567;
wire S8568;
wire S8569;
wire S8570;
wire S8571;
wire S8572;
wire S8573;
wire S8574;
wire S8575;
wire S8576;
wire S8577;
wire S8578;
wire S8579;
wire S8580;
wire S8581;
wire S8582;
wire S8583;
wire S8584;
wire S8585;
wire S8586;
wire S8587;
wire S8588;
wire S8589;
wire S8590;
wire S8591;
wire controller_1115_S_0;
wire controller_1405_Y_0;
wire controller_1405_Y_1;
wire controller_216_B_0;
wire controller_389_B_0;
wire controller_389_B_2;
wire controller_clk;
wire controller_fib_0;
wire controller_fib_1;
wire controller_fib_2;
wire controller_fib_3;
wire controller_fib_4;
wire controller_opcode_2;
wire controller_opcode_3;
wire controller_opcode_4;
wire controller_opcode_5;
wire controller_opcode_6;
wire controller_opcode_7;
wire controller_outflag_0;
wire controller_outflag_1;
wire controller_outflag_2;
wire controller_outflag_3;
wire controller_outflag_6;
wire controller_outflag_7;
wire controller_pstate_0;
wire controller_pstate_1;
wire controller_readio;
wire controller_readmem;
wire controller_readymem;
wire controller_rst;
wire controller_writeio;
wire controller_writemem;
wire datapath_addrbus_0;
wire datapath_addrbus_10;
wire datapath_addrbus_11;
wire datapath_addrbus_12;
wire datapath_addrbus_13;
wire datapath_addrbus_14;
wire datapath_addrbus_15;
wire datapath_addrbus_1;
wire datapath_addrbus_2;
wire datapath_addrbus_3;
wire datapath_addrbus_4;
wire datapath_addrbus_5;
wire datapath_addrbus_6;
wire datapath_addrbus_7;
wire datapath_addrbus_8;
wire datapath_addrbus_9;
wire datapath_addsubunit_in1_0;
wire datapath_addsubunit_in1_10;
wire datapath_addsubunit_in1_11;
wire datapath_addsubunit_in1_12;
wire datapath_addsubunit_in1_13;
wire datapath_addsubunit_in1_14;
wire datapath_addsubunit_in1_15;
wire datapath_addsubunit_in1_1;
wire datapath_addsubunit_in1_2;
wire datapath_addsubunit_in1_3;
wire datapath_addsubunit_in1_4;
wire datapath_addsubunit_in1_5;
wire datapath_addsubunit_in1_6;
wire datapath_addsubunit_in1_7;
wire datapath_addsubunit_in1_8;
wire datapath_addsubunit_in1_9;
wire datapath_adr_outreg_0;
wire datapath_adr_outreg_10;
wire datapath_adr_outreg_11;
wire datapath_adr_outreg_12;
wire datapath_adr_outreg_13;
wire datapath_adr_outreg_14;
wire datapath_adr_outreg_15;
wire datapath_adr_outreg_1;
wire datapath_adr_outreg_2;
wire datapath_adr_outreg_3;
wire datapath_adr_outreg_4;
wire datapath_adr_outreg_5;
wire datapath_adr_outreg_6;
wire datapath_adr_outreg_7;
wire datapath_adr_outreg_8;
wire datapath_adr_outreg_9;
wire datapath_databusin_0;
wire datapath_databusin_10;
wire datapath_databusin_11;
wire datapath_databusin_12;
wire datapath_databusin_13;
wire datapath_databusin_14;
wire datapath_databusin_15;
wire datapath_databusin_1;
wire datapath_databusin_2;
wire datapath_databusin_3;
wire datapath_databusin_4;
wire datapath_databusin_5;
wire datapath_databusin_6;
wire datapath_databusin_7;
wire datapath_databusin_8;
wire datapath_databusin_9;
wire datapath_indatatrf_0;
wire datapath_indatatrf_10;
wire datapath_indatatrf_11;
wire datapath_indatatrf_12;
wire datapath_indatatrf_13;
wire datapath_indatatrf_14;
wire datapath_indatatrf_15;
wire datapath_indatatrf_1;
wire datapath_indatatrf_2;
wire datapath_indatatrf_3;
wire datapath_indatatrf_4;
wire datapath_indatatrf_5;
wire datapath_indatatrf_6;
wire datapath_indatatrf_7;
wire datapath_indatatrf_8;
wire datapath_indatatrf_9;
wire datapath_instruction_0;
wire datapath_instruction_1;
wire datapath_instruction_2;
wire datapath_instruction_3;
wire datapath_multdivunit_outmdu1_0;
wire datapath_multdivunit_outmdu1_10;
wire datapath_multdivunit_outmdu1_11;
wire datapath_multdivunit_outmdu1_12;
wire datapath_multdivunit_outmdu1_13;
wire datapath_multdivunit_outmdu1_14;
wire datapath_multdivunit_outmdu1_15;
wire datapath_multdivunit_outmdu1_1;
wire datapath_multdivunit_outmdu1_2;
wire datapath_multdivunit_outmdu1_3;
wire datapath_multdivunit_outmdu1_4;
wire datapath_multdivunit_outmdu1_5;
wire datapath_multdivunit_outmdu1_6;
wire datapath_multdivunit_outmdu1_7;
wire datapath_multdivunit_outmdu1_8;
wire datapath_multdivunit_outmdu1_9;
wire datapath_multdivunit_outmdu2_0;
wire datapath_multdivunit_outmdu2_10;
wire datapath_multdivunit_outmdu2_11;
wire datapath_multdivunit_outmdu2_12;
wire datapath_multdivunit_outmdu2_13;
wire datapath_multdivunit_outmdu2_14;
wire datapath_multdivunit_outmdu2_15;
wire datapath_multdivunit_outmdu2_1;
wire datapath_multdivunit_outmdu2_2;
wire datapath_multdivunit_outmdu2_3;
wire datapath_multdivunit_outmdu2_4;
wire datapath_multdivunit_outmdu2_5;
wire datapath_multdivunit_outmdu2_6;
wire datapath_multdivunit_outmdu2_7;
wire datapath_multdivunit_outmdu2_8;
wire datapath_multdivunit_outmdu2_9;
wire datapath_muxmem_in2_0;
wire datapath_muxmem_in2_10;
wire datapath_muxmem_in2_11;
wire datapath_muxmem_in2_12;
wire datapath_muxmem_in2_13;
wire datapath_muxmem_in2_14;
wire datapath_muxmem_in2_15;
wire datapath_muxmem_in2_1;
wire datapath_muxmem_in2_2;
wire datapath_muxmem_in2_3;
wire datapath_muxmem_in2_4;
wire datapath_muxmem_in2_5;
wire datapath_muxmem_in2_6;
wire datapath_muxmem_in2_7;
wire datapath_muxmem_in2_8;
wire datapath_muxmem_in2_9;
wire datapath_shiftunit_2135_A;
wire datapath_shiftunit_2153_A;
wire datapath_shiftunit_2171_A;
wire datapath_shiftunit_2189_A;
wire datapath_shiftunit_2207_A;
wire datapath_shiftunit_2225_A;
wire datapath_shiftunit_2243_A;
wire datapath_shiftunit_2261_A;
wire datapath_shiftunit_2279_A;
wire datapath_shiftunit_2297_A;
wire datapath_shiftunit_2315_A;
wire datapath_shiftunit_2333_A;
wire datapath_shiftunit_2351_A;
wire datapath_shiftunit_2369_A;
wire datapath_shiftunit_2387_A;
wire datapath_shiftunit_2405_A;
wire datapath_shiftunit_2439_A;
wire datapath_shiftunit_2457_A;
wire datapath_shiftunit_2475_A;
wire datapath_shiftunit_2493_A;
wire datapath_shiftunit_2511_A;
wire datapath_shiftunit_2529_A;
wire datapath_shiftunit_2547_A;
wire datapath_shiftunit_2565_A;
wire datapath_shiftunit_2583_A;
wire datapath_shiftunit_2601_A;
wire datapath_shiftunit_2619_A;
wire datapath_shiftunit_2637_A;
wire datapath_shiftunit_2655_A;
wire datapath_shiftunit_2673_A;
wire datapath_shiftunit_2691_A;
wire datapath_shiftunit_2708_A;
wire datapath_theregisterfile_memtrf_0;
wire datapath_theregisterfile_memtrf_100;
wire datapath_theregisterfile_memtrf_101;
wire datapath_theregisterfile_memtrf_102;
wire datapath_theregisterfile_memtrf_103;
wire datapath_theregisterfile_memtrf_104;
wire datapath_theregisterfile_memtrf_105;
wire datapath_theregisterfile_memtrf_106;
wire datapath_theregisterfile_memtrf_107;
wire datapath_theregisterfile_memtrf_108;
wire datapath_theregisterfile_memtrf_109;
wire datapath_theregisterfile_memtrf_10;
wire datapath_theregisterfile_memtrf_110;
wire datapath_theregisterfile_memtrf_111;
wire datapath_theregisterfile_memtrf_112;
wire datapath_theregisterfile_memtrf_113;
wire datapath_theregisterfile_memtrf_114;
wire datapath_theregisterfile_memtrf_115;
wire datapath_theregisterfile_memtrf_116;
wire datapath_theregisterfile_memtrf_117;
wire datapath_theregisterfile_memtrf_118;
wire datapath_theregisterfile_memtrf_119;
wire datapath_theregisterfile_memtrf_11;
wire datapath_theregisterfile_memtrf_120;
wire datapath_theregisterfile_memtrf_121;
wire datapath_theregisterfile_memtrf_122;
wire datapath_theregisterfile_memtrf_123;
wire datapath_theregisterfile_memtrf_124;
wire datapath_theregisterfile_memtrf_125;
wire datapath_theregisterfile_memtrf_126;
wire datapath_theregisterfile_memtrf_127;
wire datapath_theregisterfile_memtrf_128;
wire datapath_theregisterfile_memtrf_129;
wire datapath_theregisterfile_memtrf_12;
wire datapath_theregisterfile_memtrf_130;
wire datapath_theregisterfile_memtrf_131;
wire datapath_theregisterfile_memtrf_132;
wire datapath_theregisterfile_memtrf_133;
wire datapath_theregisterfile_memtrf_134;
wire datapath_theregisterfile_memtrf_135;
wire datapath_theregisterfile_memtrf_136;
wire datapath_theregisterfile_memtrf_137;
wire datapath_theregisterfile_memtrf_138;
wire datapath_theregisterfile_memtrf_139;
wire datapath_theregisterfile_memtrf_13;
wire datapath_theregisterfile_memtrf_140;
wire datapath_theregisterfile_memtrf_141;
wire datapath_theregisterfile_memtrf_142;
wire datapath_theregisterfile_memtrf_143;
wire datapath_theregisterfile_memtrf_144;
wire datapath_theregisterfile_memtrf_145;
wire datapath_theregisterfile_memtrf_146;
wire datapath_theregisterfile_memtrf_147;
wire datapath_theregisterfile_memtrf_148;
wire datapath_theregisterfile_memtrf_149;
wire datapath_theregisterfile_memtrf_14;
wire datapath_theregisterfile_memtrf_150;
wire datapath_theregisterfile_memtrf_151;
wire datapath_theregisterfile_memtrf_152;
wire datapath_theregisterfile_memtrf_153;
wire datapath_theregisterfile_memtrf_154;
wire datapath_theregisterfile_memtrf_155;
wire datapath_theregisterfile_memtrf_156;
wire datapath_theregisterfile_memtrf_157;
wire datapath_theregisterfile_memtrf_158;
wire datapath_theregisterfile_memtrf_159;
wire datapath_theregisterfile_memtrf_15;
wire datapath_theregisterfile_memtrf_160;
wire datapath_theregisterfile_memtrf_161;
wire datapath_theregisterfile_memtrf_162;
wire datapath_theregisterfile_memtrf_163;
wire datapath_theregisterfile_memtrf_164;
wire datapath_theregisterfile_memtrf_165;
wire datapath_theregisterfile_memtrf_166;
wire datapath_theregisterfile_memtrf_167;
wire datapath_theregisterfile_memtrf_168;
wire datapath_theregisterfile_memtrf_169;
wire datapath_theregisterfile_memtrf_16;
wire datapath_theregisterfile_memtrf_170;
wire datapath_theregisterfile_memtrf_171;
wire datapath_theregisterfile_memtrf_172;
wire datapath_theregisterfile_memtrf_173;
wire datapath_theregisterfile_memtrf_174;
wire datapath_theregisterfile_memtrf_175;
wire datapath_theregisterfile_memtrf_176;
wire datapath_theregisterfile_memtrf_177;
wire datapath_theregisterfile_memtrf_178;
wire datapath_theregisterfile_memtrf_179;
wire datapath_theregisterfile_memtrf_17;
wire datapath_theregisterfile_memtrf_180;
wire datapath_theregisterfile_memtrf_181;
wire datapath_theregisterfile_memtrf_182;
wire datapath_theregisterfile_memtrf_183;
wire datapath_theregisterfile_memtrf_184;
wire datapath_theregisterfile_memtrf_185;
wire datapath_theregisterfile_memtrf_186;
wire datapath_theregisterfile_memtrf_187;
wire datapath_theregisterfile_memtrf_188;
wire datapath_theregisterfile_memtrf_189;
wire datapath_theregisterfile_memtrf_18;
wire datapath_theregisterfile_memtrf_190;
wire datapath_theregisterfile_memtrf_191;
wire datapath_theregisterfile_memtrf_192;
wire datapath_theregisterfile_memtrf_193;
wire datapath_theregisterfile_memtrf_194;
wire datapath_theregisterfile_memtrf_195;
wire datapath_theregisterfile_memtrf_196;
wire datapath_theregisterfile_memtrf_197;
wire datapath_theregisterfile_memtrf_198;
wire datapath_theregisterfile_memtrf_199;
wire datapath_theregisterfile_memtrf_19;
wire datapath_theregisterfile_memtrf_1;
wire datapath_theregisterfile_memtrf_200;
wire datapath_theregisterfile_memtrf_201;
wire datapath_theregisterfile_memtrf_202;
wire datapath_theregisterfile_memtrf_203;
wire datapath_theregisterfile_memtrf_204;
wire datapath_theregisterfile_memtrf_205;
wire datapath_theregisterfile_memtrf_206;
wire datapath_theregisterfile_memtrf_207;
wire datapath_theregisterfile_memtrf_208;
wire datapath_theregisterfile_memtrf_209;
wire datapath_theregisterfile_memtrf_20;
wire datapath_theregisterfile_memtrf_210;
wire datapath_theregisterfile_memtrf_211;
wire datapath_theregisterfile_memtrf_212;
wire datapath_theregisterfile_memtrf_213;
wire datapath_theregisterfile_memtrf_214;
wire datapath_theregisterfile_memtrf_215;
wire datapath_theregisterfile_memtrf_216;
wire datapath_theregisterfile_memtrf_217;
wire datapath_theregisterfile_memtrf_218;
wire datapath_theregisterfile_memtrf_219;
wire datapath_theregisterfile_memtrf_21;
wire datapath_theregisterfile_memtrf_220;
wire datapath_theregisterfile_memtrf_221;
wire datapath_theregisterfile_memtrf_222;
wire datapath_theregisterfile_memtrf_223;
wire datapath_theregisterfile_memtrf_224;
wire datapath_theregisterfile_memtrf_225;
wire datapath_theregisterfile_memtrf_226;
wire datapath_theregisterfile_memtrf_227;
wire datapath_theregisterfile_memtrf_228;
wire datapath_theregisterfile_memtrf_229;
wire datapath_theregisterfile_memtrf_22;
wire datapath_theregisterfile_memtrf_230;
wire datapath_theregisterfile_memtrf_231;
wire datapath_theregisterfile_memtrf_232;
wire datapath_theregisterfile_memtrf_233;
wire datapath_theregisterfile_memtrf_234;
wire datapath_theregisterfile_memtrf_235;
wire datapath_theregisterfile_memtrf_236;
wire datapath_theregisterfile_memtrf_237;
wire datapath_theregisterfile_memtrf_238;
wire datapath_theregisterfile_memtrf_239;
wire datapath_theregisterfile_memtrf_23;
wire datapath_theregisterfile_memtrf_240;
wire datapath_theregisterfile_memtrf_241;
wire datapath_theregisterfile_memtrf_242;
wire datapath_theregisterfile_memtrf_243;
wire datapath_theregisterfile_memtrf_244;
wire datapath_theregisterfile_memtrf_245;
wire datapath_theregisterfile_memtrf_246;
wire datapath_theregisterfile_memtrf_247;
wire datapath_theregisterfile_memtrf_248;
wire datapath_theregisterfile_memtrf_249;
wire datapath_theregisterfile_memtrf_24;
wire datapath_theregisterfile_memtrf_250;
wire datapath_theregisterfile_memtrf_251;
wire datapath_theregisterfile_memtrf_252;
wire datapath_theregisterfile_memtrf_253;
wire datapath_theregisterfile_memtrf_254;
wire datapath_theregisterfile_memtrf_255;
wire datapath_theregisterfile_memtrf_25;
wire datapath_theregisterfile_memtrf_26;
wire datapath_theregisterfile_memtrf_27;
wire datapath_theregisterfile_memtrf_28;
wire datapath_theregisterfile_memtrf_29;
wire datapath_theregisterfile_memtrf_2;
wire datapath_theregisterfile_memtrf_30;
wire datapath_theregisterfile_memtrf_31;
wire datapath_theregisterfile_memtrf_32;
wire datapath_theregisterfile_memtrf_33;
wire datapath_theregisterfile_memtrf_34;
wire datapath_theregisterfile_memtrf_35;
wire datapath_theregisterfile_memtrf_36;
wire datapath_theregisterfile_memtrf_37;
wire datapath_theregisterfile_memtrf_38;
wire datapath_theregisterfile_memtrf_39;
wire datapath_theregisterfile_memtrf_3;
wire datapath_theregisterfile_memtrf_40;
wire datapath_theregisterfile_memtrf_41;
wire datapath_theregisterfile_memtrf_42;
wire datapath_theregisterfile_memtrf_43;
wire datapath_theregisterfile_memtrf_44;
wire datapath_theregisterfile_memtrf_45;
wire datapath_theregisterfile_memtrf_46;
wire datapath_theregisterfile_memtrf_47;
wire datapath_theregisterfile_memtrf_48;
wire datapath_theregisterfile_memtrf_49;
wire datapath_theregisterfile_memtrf_4;
wire datapath_theregisterfile_memtrf_50;
wire datapath_theregisterfile_memtrf_51;
wire datapath_theregisterfile_memtrf_52;
wire datapath_theregisterfile_memtrf_53;
wire datapath_theregisterfile_memtrf_54;
wire datapath_theregisterfile_memtrf_55;
wire datapath_theregisterfile_memtrf_56;
wire datapath_theregisterfile_memtrf_57;
wire datapath_theregisterfile_memtrf_58;
wire datapath_theregisterfile_memtrf_59;
wire datapath_theregisterfile_memtrf_5;
wire datapath_theregisterfile_memtrf_60;
wire datapath_theregisterfile_memtrf_61;
wire datapath_theregisterfile_memtrf_62;
wire datapath_theregisterfile_memtrf_63;
wire datapath_theregisterfile_memtrf_64;
wire datapath_theregisterfile_memtrf_65;
wire datapath_theregisterfile_memtrf_66;
wire datapath_theregisterfile_memtrf_67;
wire datapath_theregisterfile_memtrf_68;
wire datapath_theregisterfile_memtrf_69;
wire datapath_theregisterfile_memtrf_6;
wire datapath_theregisterfile_memtrf_70;
wire datapath_theregisterfile_memtrf_71;
wire datapath_theregisterfile_memtrf_72;
wire datapath_theregisterfile_memtrf_73;
wire datapath_theregisterfile_memtrf_74;
wire datapath_theregisterfile_memtrf_75;
wire datapath_theregisterfile_memtrf_76;
wire datapath_theregisterfile_memtrf_77;
wire datapath_theregisterfile_memtrf_78;
wire datapath_theregisterfile_memtrf_79;
wire datapath_theregisterfile_memtrf_7;
wire datapath_theregisterfile_memtrf_80;
wire datapath_theregisterfile_memtrf_81;
wire datapath_theregisterfile_memtrf_82;
wire datapath_theregisterfile_memtrf_83;
wire datapath_theregisterfile_memtrf_84;
wire datapath_theregisterfile_memtrf_85;
wire datapath_theregisterfile_memtrf_86;
wire datapath_theregisterfile_memtrf_87;
wire datapath_theregisterfile_memtrf_88;
wire datapath_theregisterfile_memtrf_89;
wire datapath_theregisterfile_memtrf_8;
wire datapath_theregisterfile_memtrf_90;
wire datapath_theregisterfile_memtrf_91;
wire datapath_theregisterfile_memtrf_92;
wire datapath_theregisterfile_memtrf_93;
wire datapath_theregisterfile_memtrf_94;
wire datapath_theregisterfile_memtrf_95;
wire datapath_theregisterfile_memtrf_96;
wire datapath_theregisterfile_memtrf_97;
wire datapath_theregisterfile_memtrf_98;
wire datapath_theregisterfile_memtrf_99;
wire datapath_theregisterfile_memtrf_9;
input clk;
input rst;
input readyMEM;
input [15:0] dataBusIn;output readMEM;
output writeMEM;
output readIO;
output writeIO;
output [15:0] dataBusOut;output [15:0] addrBus;output readInst;
output [15:0] PCout;
NOT #() 
NOT_1_ (
  .A({ datapath_multdivunit_outmdu2_15 }),
  .Y({ S7476 })
);
NOT #() 
NOT_2_ (
  .A({ controller_opcode_7 }),
  .Y({ S7487 })
);
NOT #() 
NOT_3_ (
  .A({ datapath_theregisterfile_memtrf_78 }),
  .Y({ S7498 })
);
NOT #() 
NOT_4_ (
  .A({ datapath_theregisterfile_memtrf_62 }),
  .Y({ S7509 })
);
NOT #() 
NOT_5_ (
  .A({ datapath_theregisterfile_memtrf_96 }),
  .Y({ S7520 })
);
NOT #() 
NOT_6_ (
  .A({ datapath_theregisterfile_memtrf_97 }),
  .Y({ S7531 })
);
NOT #() 
NOT_7_ (
  .A({ datapath_theregisterfile_memtrf_14 }),
  .Y({ S7542 })
);
NOT #() 
NOT_8_ (
  .A({ datapath_theregisterfile_memtrf_157 }),
  .Y({ S7553 })
);
NOT #() 
NOT_9_ (
  .A({ datapath_theregisterfile_memtrf_158 }),
  .Y({ S7564 })
);
NOT #() 
NOT_10_ (
  .A({ datapath_theregisterfile_memtrf_175 }),
  .Y({ S7574 })
);
NOT #() 
NOT_11_ (
  .A({ datapath_theregisterfile_memtrf_179 }),
  .Y({ S7585 })
);
NOT #() 
NOT_12_ (
  .A({ datapath_theregisterfile_memtrf_180 }),
  .Y({ S7596 })
);
NOT #() 
NOT_13_ (
  .A({ datapath_theregisterfile_memtrf_184 }),
  .Y({ S7607 })
);
NOT #() 
NOT_14_ (
  .A({ datapath_theregisterfile_memtrf_185 }),
  .Y({ S7618 })
);
NOT #() 
NOT_15_ (
  .A({ datapath_theregisterfile_memtrf_186 }),
  .Y({ S7629 })
);
NOT #() 
NOT_16_ (
  .A({ datapath_theregisterfile_memtrf_187 }),
  .Y({ S7640 })
);
NOT #() 
NOT_17_ (
  .A({ datapath_theregisterfile_memtrf_188 }),
  .Y({ S7651 })
);
NOT #() 
NOT_18_ (
  .A({ datapath_theregisterfile_memtrf_191 }),
  .Y({ S7662 })
);
NOT #() 
NOT_19_ (
  .A({ datapath_theregisterfile_memtrf_192 }),
  .Y({ S7673 })
);
NOT #() 
NOT_20_ (
  .A({ datapath_theregisterfile_memtrf_193 }),
  .Y({ S7684 })
);
NOT #() 
NOT_21_ (
  .A({ datapath_theregisterfile_memtrf_195 }),
  .Y({ S7695 })
);
NOT #() 
NOT_22_ (
  .A({ datapath_theregisterfile_memtrf_197 }),
  .Y({ S7706 })
);
NOT #() 
NOT_23_ (
  .A({ datapath_theregisterfile_memtrf_198 }),
  .Y({ S7717 })
);
NOT #() 
NOT_24_ (
  .A({ datapath_theregisterfile_memtrf_199 }),
  .Y({ S7728 })
);
NOT #() 
NOT_25_ (
  .A({ datapath_theregisterfile_memtrf_200 }),
  .Y({ S7739 })
);
NOT #() 
NOT_26_ (
  .A({ datapath_theregisterfile_memtrf_204 }),
  .Y({ S7750 })
);
NOT #() 
NOT_27_ (
  .A({ datapath_theregisterfile_memtrf_205 }),
  .Y({ S7761 })
);
NOT #() 
NOT_28_ (
  .A({ datapath_theregisterfile_memtrf_206 }),
  .Y({ S7772 })
);
NOT #() 
NOT_29_ (
  .A({ datapath_theregisterfile_memtrf_224 }),
  .Y({ S7783 })
);
NOT #() 
NOT_30_ (
  .A({ datapath_theregisterfile_memtrf_225 }),
  .Y({ S7794 })
);
NOT #() 
NOT_31_ (
  .A({ datapath_theregisterfile_memtrf_226 }),
  .Y({ S7805 })
);
NOT #() 
NOT_32_ (
  .A({ datapath_theregisterfile_memtrf_228 }),
  .Y({ S7816 })
);
NOT #() 
NOT_33_ (
  .A({ datapath_theregisterfile_memtrf_229 }),
  .Y({ S7822 })
);
NOT #() 
NOT_34_ (
  .A({ datapath_theregisterfile_memtrf_230 }),
  .Y({ S7823 })
);
NOT #() 
NOT_35_ (
  .A({ controller_outflag_0 }),
  .Y({ S7830 })
);
NOT #() 
NOT_36_ (
  .A({ controller_outflag_1 }),
  .Y({ S7838 })
);
NOT #() 
NOT_37_ (
  .A({ controller_outflag_2 }),
  .Y({ S7846 })
);
NOT #() 
NOT_38_ (
  .A({ controller_outflag_3 }),
  .Y({ S7853 })
);
NOT #() 
NOT_39_ (
  .A({ controller_389_B_0 }),
  .Y({ S7861 })
);
NOT #() 
NOT_40_ (
  .A({ controller_389_B_2 }),
  .Y({ S7869 })
);
NOT #() 
NOT_41_ (
  .A({ controller_outflag_6 }),
  .Y({ S7876 })
);
NOT #() 
NOT_42_ (
  .A({ datapath_muxmem_in2_0 }),
  .Y({ S7884 })
);
NOT #() 
NOT_43_ (
  .A({ datapath_muxmem_in2_1 }),
  .Y({ S7892 })
);
NOT #() 
NOT_44_ (
  .A({ datapath_muxmem_in2_2 }),
  .Y({ S7897 })
);
NOT #() 
NOT_45_ (
  .A({ datapath_muxmem_in2_3 }),
  .Y({ S7905 })
);
NOT #() 
NOT_46_ (
  .A({ datapath_muxmem_in2_4 }),
  .Y({ S7913 })
);
NOT #() 
NOT_47_ (
  .A({ datapath_muxmem_in2_5 }),
  .Y({ S7920 })
);
NOT #() 
NOT_48_ (
  .A({ datapath_muxmem_in2_6 }),
  .Y({ S7928 })
);
NOT #() 
NOT_49_ (
  .A({ datapath_muxmem_in2_7 }),
  .Y({ S7936 })
);
NOT #() 
NOT_50_ (
  .A({ datapath_muxmem_in2_8 }),
  .Y({ S7946 })
);
NOT #() 
NOT_51_ (
  .A({ datapath_muxmem_in2_9 }),
  .Y({ S7957 })
);
NOT #() 
NOT_52_ (
  .A({ datapath_muxmem_in2_10 }),
  .Y({ S7968 })
);
NOT #() 
NOT_53_ (
  .A({ datapath_muxmem_in2_11 }),
  .Y({ S7978 })
);
NOT #() 
NOT_54_ (
  .A({ datapath_muxmem_in2_12 }),
  .Y({ S7989 })
);
NOT #() 
NOT_55_ (
  .A({ datapath_muxmem_in2_13 }),
  .Y({ S8000 })
);
NOT #() 
NOT_56_ (
  .A({ datapath_multdivunit_outmdu1_2 }),
  .Y({ S8011 })
);
NOT #() 
NOT_57_ (
  .A({ datapath_multdivunit_outmdu1_6 }),
  .Y({ S8022 })
);
NOT #() 
NOT_58_ (
  .A({ datapath_multdivunit_outmdu2_0 }),
  .Y({ S8033 })
);
NOT #() 
NOT_59_ (
  .A({ datapath_multdivunit_outmdu2_1 }),
  .Y({ S8044 })
);
NOT #() 
NOT_60_ (
  .A({ datapath_multdivunit_outmdu2_2 }),
  .Y({ S8054 })
);
NOT #() 
NOT_61_ (
  .A({ datapath_multdivunit_outmdu2_3 }),
  .Y({ S8065 })
);
NOT #() 
NOT_62_ (
  .A({ datapath_multdivunit_outmdu2_4 }),
  .Y({ S8076 })
);
NOT #() 
NOT_63_ (
  .A({ datapath_multdivunit_outmdu2_5 }),
  .Y({ S8087 })
);
NOT #() 
NOT_64_ (
  .A({ datapath_multdivunit_outmdu2_6 }),
  .Y({ S8097 })
);
NOT #() 
NOT_65_ (
  .A({ datapath_multdivunit_outmdu2_7 }),
  .Y({ S8108 })
);
NOT #() 
NOT_66_ (
  .A({ datapath_multdivunit_outmdu2_8 }),
  .Y({ S8119 })
);
NOT #() 
NOT_67_ (
  .A({ datapath_multdivunit_outmdu2_9 }),
  .Y({ S8129 })
);
NOT #() 
NOT_68_ (
  .A({ datapath_multdivunit_outmdu2_10 }),
  .Y({ S8140 })
);
NOT #() 
NOT_69_ (
  .A({ datapath_multdivunit_outmdu2_11 }),
  .Y({ S8151 })
);
NOT #() 
NOT_70_ (
  .A({ datapath_multdivunit_outmdu2_12 }),
  .Y({ S8161 })
);
NOT #() 
NOT_71_ (
  .A({ datapath_multdivunit_outmdu2_13 }),
  .Y({ S8172 })
);
NOT #() 
NOT_72_ (
  .A({ datapath_multdivunit_outmdu2_14 }),
  .Y({ S8183 })
);
NOT #() 
NOT_73_ (
  .A({ datapath_instruction_2 }),
  .Y({ S8193 })
);
NOT #() 
NOT_74_ (
  .A({ datapath_instruction_3 }),
  .Y({ S8204 })
);
NOT #() 
NOT_75_ (
  .A({ controller_fib_0 }),
  .Y({ S8215 })
);
NOT #() 
NOT_76_ (
  .A({ controller_fib_1 }),
  .Y({ S8225 })
);
NOT #() 
NOT_77_ (
  .A({ datapath_databusin_5 }),
  .Y({ S8236 })
);
NOT #() 
NOT_78_ (
  .A({ controller_fib_2 }),
  .Y({ S8246 })
);
NOT #() 
NOT_79_ (
  .A({ datapath_databusin_6 }),
  .Y({ S8257 })
);
NOT #() 
NOT_80_ (
  .A({ controller_fib_4 }),
  .Y({ S8267 })
);
NOT #() 
NOT_81_ (
  .A({ controller_216_B_0 }),
  .Y({ S8278 })
);
NOT #() 
NOT_82_ (
  .A({ datapath_databusin_9 }),
  .Y({ S8288 })
);
NOT #() 
NOT_83_ (
  .A({ controller_opcode_2 }),
  .Y({ S8299 })
);
NOT #() 
NOT_84_ (
  .A({ controller_opcode_3 }),
  .Y({ S8309 })
);
NOT #() 
NOT_85_ (
  .A({ controller_opcode_4 }),
  .Y({ S8319 })
);
NOT #() 
NOT_86_ (
  .A({ controller_opcode_5 }),
  .Y({ S8329 })
);
NOT #() 
NOT_87_ (
  .A({ controller_opcode_6 }),
  .Y({ S8339 })
);
NOT #() 
NOT_88_ (
  .A({ controller_outflag_7 }),
  .Y({ S8349 })
);
NOT #() 
NOT_89_ (
  .A({ controller_pstate_1 }),
  .Y({ S8356 })
);
NOT #() 
NOT_90_ (
  .A({ controller_pstate_0 }),
  .Y({ S8365 })
);
NOR #() 
NOR_1_ (
  .A({ controller_pstate_1 }),
  .B({ S8365 }),
  .Y({ S8375 })
);
NAND #() 
NAND_1_ (
  .A({ S8356 }),
  .B({ controller_pstate_0 }),
  .Y({ S8385 })
);
NOR #() 
NOR_2_ (
  .A({ S7487 }),
  .B({ S8339 }),
  .Y({ S8395 })
);
NAND #() 
NAND_2_ (
  .A({ controller_opcode_7 }),
  .B({ controller_opcode_6 }),
  .Y({ S8405 })
);
NOR #() 
NOR_3_ (
  .A({ controller_opcode_4 }),
  .B({ controller_opcode_5 }),
  .Y({ S8416 })
);
NAND #() 
NAND_3_ (
  .A({ S8319 }),
  .B({ S8329 }),
  .Y({ S8426 })
);
NOR #() 
NOR_4_ (
  .A({ S8405 }),
  .B({ S8416 }),
  .Y({ S8436 })
);
NOT #() 
NOT_91_ (
  .A({ S8436 }),
  .Y({ S8447 })
);
NOR #() 
NOR_5_ (
  .A({ S8319 }),
  .B({ S8329 }),
  .Y({ S8457 })
);
NAND #() 
NAND_4_ (
  .A({ controller_opcode_4 }),
  .B({ controller_opcode_5 }),
  .Y({ S8468 })
);
NOR #() 
NOR_6_ (
  .A({ controller_opcode_7 }),
  .B({ controller_opcode_6 }),
  .Y({ S8478 })
);
NAND #() 
NAND_5_ (
  .A({ S7487 }),
  .B({ S8339 }),
  .Y({ S8489 })
);
NAND #() 
NAND_6_ (
  .A({ S8468 }),
  .B({ S8478 }),
  .Y({ S8499 })
);
NAND #() 
NAND_7_ (
  .A({ S8447 }),
  .B({ S8499 }),
  .Y({ S8510 })
);
NOT #() 
NOT_92_ (
  .A({ S8510 }),
  .Y({ S8520 })
);
NOR #() 
NOR_7_ (
  .A({ controller_opcode_5 }),
  .B({ S8489 }),
  .Y({ S8531 })
);
NOR #() 
NOR_8_ (
  .A({ controller_opcode_2 }),
  .B({ S8309 }),
  .Y({ S8541 })
);
NAND #() 
NAND_8_ (
  .A({ S8299 }),
  .B({ controller_opcode_3 }),
  .Y({ S8542 })
);
NOR #() 
NOR_9_ (
  .A({ S8405 }),
  .B({ S8468 }),
  .Y({ S8543 })
);
NAND #() 
NAND_9_ (
  .A({ S8395 }),
  .B({ S8457 }),
  .Y({ S8544 })
);
NAND #() 
NAND_10_ (
  .A({ S8541 }),
  .B({ S8543 }),
  .Y({ S8545 })
);
NOT #() 
NOT_93_ (
  .A({ S8545 }),
  .Y({ S8546 })
);
NAND #() 
NAND_11_ (
  .A({ S8510 }),
  .B({ S8545 }),
  .Y({ S8547 })
);
NOR #() 
NOR_10_ (
  .A({ S8531 }),
  .B({ S8547 }),
  .Y({ S8548 })
);
NOT #() 
NOT_94_ (
  .A({ S8548 }),
  .Y({ S8549 })
);
NOR #() 
NOR_11_ (
  .A({ S8299 }),
  .B({ controller_opcode_3 }),
  .Y({ S8550 })
);
NAND #() 
NAND_12_ (
  .A({ controller_opcode_2 }),
  .B({ S8309 }),
  .Y({ S8551 })
);
NAND #() 
NAND_13_ (
  .A({ controller_fib_1 }),
  .B({ controller_fib_2 }),
  .Y({ S8552 })
);
NOR #() 
NOR_12_ (
  .A({ S8551 }),
  .B({ S8552 }),
  .Y({ S8553 })
);
NAND #() 
NAND_14_ (
  .A({ S8542 }),
  .B({ S8543 }),
  .Y({ S8554 })
);
NOR #() 
NOR_13_ (
  .A({ S8553 }),
  .B({ S8554 }),
  .Y({ S8555 })
);
NOR #() 
NOR_14_ (
  .A({ controller_opcode_4 }),
  .B({ S8329 }),
  .Y({ S8556 })
);
NAND #() 
NAND_15_ (
  .A({ S8319 }),
  .B({ controller_opcode_5 }),
  .Y({ S8557 })
);
NOR #() 
NOR_15_ (
  .A({ S8489 }),
  .B({ S8557 }),
  .Y({ S8558 })
);
NAND #() 
NAND_16_ (
  .A({ S8478 }),
  .B({ S8556 }),
  .Y({ S8559 })
);
NAND #() 
NAND_17_ (
  .A({ controller_opcode_3 }),
  .B({ S8558 }),
  .Y({ S8560 })
);
NAND #() 
NAND_18_ (
  .A({ S8548 }),
  .B({ S8560 }),
  .Y({ S8561 })
);
NOR #() 
NOR_16_ (
  .A({ S8555 }),
  .B({ S8561 }),
  .Y({ S8562 })
);
NOR #() 
NOR_17_ (
  .A({ S8385 }),
  .B({ S8562 }),
  .Y({ S8563 })
);
NOR #() 
NOR_18_ (
  .A({ S8416 }),
  .B({ S8457 }),
  .Y({ S8564 })
);
NAND #() 
NAND_19_ (
  .A({ S8426 }),
  .B({ S8468 }),
  .Y({ S8565 })
);
NAND #() 
NAND_20_ (
  .A({ controller_pstate_1 }),
  .B({ S8436 }),
  .Y({ S8566 })
);
NOT #() 
NOT_95_ (
  .A({ S8566 }),
  .Y({ S8567 })
);
NOR #() 
NOR_19_ (
  .A({ S8457 }),
  .B({ S8566 }),
  .Y({ S8568 })
);
NAND #() 
NAND_21_ (
  .A({ S8468 }),
  .B({ S8567 }),
  .Y({ S8569 })
);
NOR #() 
NOR_20_ (
  .A({ S8365 }),
  .B({ S8569 }),
  .Y({ S8570 })
);
NAND #() 
NAND_22_ (
  .A({ controller_pstate_0 }),
  .B({ S8568 }),
  .Y({ S8571 })
);
NOR #() 
NOR_21_ (
  .A({ controller_216_B_0 }),
  .B({ controller_readymem }),
  .Y({ S8572 })
);
NOT #() 
NOT_96_ (
  .A({ S8572 }),
  .Y({ S8573 })
);
NOR #() 
NOR_22_ (
  .A({ controller_opcode_3 }),
  .B({ S8356 }),
  .Y({ S8574 })
);
NAND #() 
NAND_23_ (
  .A({ S8365 }),
  .B({ S8574 }),
  .Y({ S8575 })
);
NOR #() 
NOR_23_ (
  .A({ S8559 }),
  .B({ S8575 }),
  .Y({ S8576 })
);
NOT #() 
NOT_97_ (
  .A({ S8576 }),
  .Y({ S8577 })
);
NAND #() 
NAND_24_ (
  .A({ S8573 }),
  .B({ S8576 }),
  .Y({ S8578 })
);
NAND #() 
NAND_25_ (
  .A({ S8571 }),
  .B({ S8578 }),
  .Y({ S8579 })
);
NOR #() 
NOR_24_ (
  .A({ S8563 }),
  .B({ S8579 }),
  .Y({ S8580 })
);
NAND #() 
NAND_26_ (
  .A({ datapath_muxmem_in2_15 }),
  .B({ S8580 }),
  .Y({ S8581 })
);
NAND #() 
NAND_27_ (
  .A({ controller_216_B_0 }),
  .B({ S8543 }),
  .Y({ S8582 })
);
NAND #() 
NAND_28_ (
  .A({ controller_fib_0 }),
  .B({ controller_fib_2 }),
  .Y({ S8583 })
);
NOR #() 
NOR_25_ (
  .A({ controller_fib_1 }),
  .B({ S8583 }),
  .Y({ S8584 })
);
NAND #() 
NAND_29_ (
  .A({ S7861 }),
  .B({ S8584 }),
  .Y({ S8585 })
);
NOR #() 
NOR_26_ (
  .A({ S8225 }),
  .B({ controller_fib_2 }),
  .Y({ S8586 })
);
NOR #() 
NOR_27_ (
  .A({ controller_389_B_0 }),
  .B({ controller_389_B_2 }),
  .Y({ S8587 })
);
NOR #() 
NOR_28_ (
  .A({ controller_389_B_2 }),
  .B({ controller_fib_0 }),
  .Y({ S8588 })
);
NOT #() 
NOT_98_ (
  .A({ S8588 }),
  .Y({ S8589 })
);
NAND #() 
NAND_30_ (
  .A({ S8586 }),
  .B({ S8589 }),
  .Y({ S8590 })
);
NOR #() 
NOR_29_ (
  .A({ S8587 }),
  .B({ S8590 }),
  .Y({ S8591 })
);
NOR #() 
NOR_30_ (
  .A({ S8215 }),
  .B({ controller_fib_2 }),
  .Y({ S344 })
);
NAND #() 
NAND_31_ (
  .A({ controller_fib_0 }),
  .B({ S8246 }),
  .Y({ S345 })
);
NOR #() 
NOR_31_ (
  .A({ controller_fib_1 }),
  .B({ S345 }),
  .Y({ S346 })
);
NOR #() 
NOR_32_ (
  .A({ controller_fib_0 }),
  .B({ controller_fib_1 }),
  .Y({ S347 })
);
NAND #() 
NAND_32_ (
  .A({ controller_fib_2 }),
  .B({ S347 }),
  .Y({ S348 })
);
NOT #() 
NOT_99_ (
  .A({ S348 }),
  .Y({ S349 })
);
NOR #() 
NOR_33_ (
  .A({ S346 }),
  .B({ S349 }),
  .Y({ S350 })
);
NOR #() 
NOR_34_ (
  .A({ controller_389_B_2 }),
  .B({ S350 }),
  .Y({ S351 })
);
NOR #() 
NOR_35_ (
  .A({ controller_389_B_0 }),
  .B({ S351 }),
  .Y({ S352 })
);
NAND #() 
NAND_33_ (
  .A({ S8246 }),
  .B({ S347 }),
  .Y({ S353 })
);
NOR #() 
NOR_36_ (
  .A({ S7861 }),
  .B({ S347 }),
  .Y({ S354 })
);
NOR #() 
NOR_37_ (
  .A({ S352 }),
  .B({ S354 }),
  .Y({ S355 })
);
NOR #() 
NOR_38_ (
  .A({ S8591 }),
  .B({ S355 }),
  .Y({ S356 })
);
NAND #() 
NAND_34_ (
  .A({ S8585 }),
  .B({ S356 }),
  .Y({ S357 })
);
NAND #() 
NAND_35_ (
  .A({ S8550 }),
  .B({ S357 }),
  .Y({ S358 })
);
NOT #() 
NOT_100_ (
  .A({ S358 }),
  .Y({ S359 })
);
NOR #() 
NOR_39_ (
  .A({ S8551 }),
  .B({ S8582 }),
  .Y({ S360 })
);
NOT #() 
NOT_101_ (
  .A({ S360 }),
  .Y({ S361 })
);
NAND #() 
NAND_36_ (
  .A({ S357 }),
  .B({ S360 }),
  .Y({ S362 })
);
NAND #() 
NAND_37_ (
  .A({ S8560 }),
  .B({ S362 }),
  .Y({ S363 })
);
NAND #() 
NAND_38_ (
  .A({ S8375 }),
  .B({ S363 }),
  .Y({ S364 })
);
NOT #() 
NOT_102_ (
  .A({ S364 }),
  .Y({ S365 })
);
NAND #() 
NAND_39_ (
  .A({ controller_opcode_2 }),
  .B({ controller_opcode_3 }),
  .Y({ S366 })
);
NOT #() 
NOT_103_ (
  .A({ S366 }),
  .Y({ S367 })
);
NOR #() 
NOR_40_ (
  .A({ S8385 }),
  .B({ S8559 }),
  .Y({ S368 })
);
NAND #() 
NAND_40_ (
  .A({ S8375 }),
  .B({ S8558 }),
  .Y({ S369 })
);
NOR #() 
NOR_41_ (
  .A({ S366 }),
  .B({ S369 }),
  .Y({ S370 })
);
NOT #() 
NOT_104_ (
  .A({ S370 }),
  .Y({ S371 })
);
NAND #() 
NAND_41_ (
  .A({ controller_216_B_0 }),
  .B({ S370 }),
  .Y({ S372 })
);
NOR #() 
NOR_42_ (
  .A({ S8541 }),
  .B({ S8550 }),
  .Y({ S373 })
);
NAND #() 
NAND_42_ (
  .A({ controller_216_B_0 }),
  .B({ S373 }),
  .Y({ S374 })
);
NAND #() 
NAND_43_ (
  .A({ S358 }),
  .B({ S374 }),
  .Y({ S375 })
);
NOR #() 
NOR_43_ (
  .A({ S8385 }),
  .B({ S8405 }),
  .Y({ S376 })
);
NAND #() 
NAND_44_ (
  .A({ S8375 }),
  .B({ S8395 }),
  .Y({ S377 })
);
NAND #() 
NAND_45_ (
  .A({ controller_opcode_4 }),
  .B({ S8375 }),
  .Y({ S378 })
);
NOR #() 
NOR_44_ (
  .A({ S8385 }),
  .B({ S8544 }),
  .Y({ S379 })
);
NAND #() 
NAND_46_ (
  .A({ S8375 }),
  .B({ S8543 }),
  .Y({ S380 })
);
NAND #() 
NAND_47_ (
  .A({ S375 }),
  .B({ S379 }),
  .Y({ S381 })
);
NOR #() 
NOR_45_ (
  .A({ controller_opcode_7 }),
  .B({ S8339 }),
  .Y({ S382 })
);
NAND #() 
NAND_48_ (
  .A({ S7487 }),
  .B({ controller_opcode_6 }),
  .Y({ S383 })
);
NOR #() 
NOR_46_ (
  .A({ S8557 }),
  .B({ S383 }),
  .Y({ S384 })
);
NOR #() 
NOR_47_ (
  .A({ S8546 }),
  .B({ S384 }),
  .Y({ S385 })
);
NOR #() 
NOR_48_ (
  .A({ S8551 }),
  .B({ S8559 }),
  .Y({ S386 })
);
NAND #() 
NAND_49_ (
  .A({ controller_opcode_7 }),
  .B({ S8339 }),
  .Y({ S387 })
);
NOR #() 
NOR_49_ (
  .A({ S8319 }),
  .B({ S387 }),
  .Y({ S388 })
);
NOR #() 
NOR_50_ (
  .A({ S8468 }),
  .B({ S387 }),
  .Y({ S389 })
);
NOT #() 
NOT_105_ (
  .A({ S389 }),
  .Y({ S390 })
);
NAND #() 
NAND_50_ (
  .A({ controller_opcode_6 }),
  .B({ S8416 }),
  .Y({ S391 })
);
NAND #() 
NAND_51_ (
  .A({ S390 }),
  .B({ S391 }),
  .Y({ S392 })
);
NOR #() 
NOR_51_ (
  .A({ S386 }),
  .B({ S392 }),
  .Y({ S393 })
);
NAND #() 
NAND_52_ (
  .A({ S385 }),
  .B({ S393 }),
  .Y({ S394 })
);
NAND #() 
NAND_53_ (
  .A({ S8375 }),
  .B({ S394 }),
  .Y({ S395 })
);
NAND #() 
NAND_54_ (
  .A({ S381 }),
  .B({ S395 }),
  .Y({ S396 })
);
NAND #() 
NAND_55_ (
  .A({ datapath_instruction_2 }),
  .B({ S396 }),
  .Y({ S397 })
);
NOT #() 
NOT_106_ (
  .A({ S397 }),
  .Y({ S398 })
);
NOR #() 
NOR_52_ (
  .A({ controller_opcode_2 }),
  .B({ S8559 }),
  .Y({ S399 })
);
NOR #() 
NOR_53_ (
  .A({ controller_216_B_0 }),
  .B({ S8544 }),
  .Y({ S400 })
);
NAND #() 
NAND_56_ (
  .A({ S8278 }),
  .B({ S8543 }),
  .Y({ S401 })
);
NAND #() 
NAND_57_ (
  .A({ S373 }),
  .B({ S400 }),
  .Y({ S402 })
);
NAND #() 
NAND_58_ (
  .A({ controller_opcode_2 }),
  .B({ S8576 }),
  .Y({ S403 })
);
NOR #() 
NOR_54_ (
  .A({ controller_opcode_7 }),
  .B({ S8468 }),
  .Y({ S404 })
);
NOT #() 
NOT_107_ (
  .A({ S404 }),
  .Y({ S405 })
);
NAND #() 
NAND_59_ (
  .A({ controller_opcode_7 }),
  .B({ S8468 }),
  .Y({ S406 })
);
NOT #() 
NOT_108_ (
  .A({ S406 }),
  .Y({ S407 })
);
NOR #() 
NOR_55_ (
  .A({ S404 }),
  .B({ S407 }),
  .Y({ S408 })
);
NOR #() 
NOR_56_ (
  .A({ S8405 }),
  .B({ S8426 }),
  .Y({ S409 })
);
NAND #() 
NAND_60_ (
  .A({ S8395 }),
  .B({ S8416 }),
  .Y({ S410 })
);
NAND #() 
NAND_61_ (
  .A({ S8375 }),
  .B({ S410 }),
  .Y({ S411 })
);
NAND #() 
NAND_62_ (
  .A({ S391 }),
  .B({ S407 }),
  .Y({ S412 })
);
NAND #() 
NAND_63_ (
  .A({ S405 }),
  .B({ S412 }),
  .Y({ S413 })
);
NOR #() 
NOR_57_ (
  .A({ S408 }),
  .B({ S411 }),
  .Y({ S414 })
);
NAND #() 
NAND_64_ (
  .A({ S8375 }),
  .B({ S413 }),
  .Y({ S415 })
);
NOR #() 
NOR_58_ (
  .A({ S399 }),
  .B({ S413 }),
  .Y({ S416 })
);
NAND #() 
NAND_65_ (
  .A({ S402 }),
  .B({ S416 }),
  .Y({ S417 })
);
NAND #() 
NAND_66_ (
  .A({ S8375 }),
  .B({ S417 }),
  .Y({ S418 })
);
NAND #() 
NAND_67_ (
  .A({ S403 }),
  .B({ S418 }),
  .Y({ S419 })
);
NAND #() 
NAND_68_ (
  .A({ controller_fib_2 }),
  .B({ S419 }),
  .Y({ S420 })
);
NOT #() 
NOT_109_ (
  .A({ S420 }),
  .Y({ S421 })
);
NOR #() 
NOR_59_ (
  .A({ S398 }),
  .B({ S421 }),
  .Y({ S422 })
);
NAND #() 
NAND_69_ (
  .A({ S397 }),
  .B({ S420 }),
  .Y({ S423 })
);
NAND #() 
NAND_70_ (
  .A({ datapath_instruction_3 }),
  .B({ S396 }),
  .Y({ S424 })
);
NOT #() 
NOT_110_ (
  .A({ S424 }),
  .Y({ S425 })
);
NAND #() 
NAND_71_ (
  .A({ controller_fib_3 }),
  .B({ S419 }),
  .Y({ S426 })
);
NOT #() 
NOT_111_ (
  .A({ S426 }),
  .Y({ S427 })
);
NOR #() 
NOR_60_ (
  .A({ S425 }),
  .B({ S427 }),
  .Y({ S428 })
);
NOR #() 
NOR_61_ (
  .A({ S422 }),
  .B({ S428 }),
  .Y({ S429 })
);
NOT #() 
NOT_112_ (
  .A({ S429 }),
  .Y({ S430 })
);
NAND #() 
NAND_72_ (
  .A({ datapath_instruction_0 }),
  .B({ S396 }),
  .Y({ S431 })
);
NOT #() 
NOT_113_ (
  .A({ S431 }),
  .Y({ S432 })
);
NAND #() 
NAND_73_ (
  .A({ controller_fib_0 }),
  .B({ S419 }),
  .Y({ S433 })
);
NOT #() 
NOT_114_ (
  .A({ S433 }),
  .Y({ S434 })
);
NOR #() 
NOR_62_ (
  .A({ S432 }),
  .B({ S434 }),
  .Y({ S435 })
);
NAND #() 
NAND_74_ (
  .A({ S431 }),
  .B({ S433 }),
  .Y({ S436 })
);
NAND #() 
NAND_75_ (
  .A({ datapath_instruction_1 }),
  .B({ S396 }),
  .Y({ S437 })
);
NOT #() 
NOT_115_ (
  .A({ S437 }),
  .Y({ S438 })
);
NAND #() 
NAND_76_ (
  .A({ controller_fib_1 }),
  .B({ S419 }),
  .Y({ S439 })
);
NOT #() 
NOT_116_ (
  .A({ S439 }),
  .Y({ S440 })
);
NOR #() 
NOR_63_ (
  .A({ S438 }),
  .B({ S440 }),
  .Y({ S441 })
);
NAND #() 
NAND_77_ (
  .A({ S437 }),
  .B({ S439 }),
  .Y({ S442 })
);
NOR #() 
NOR_64_ (
  .A({ S435 }),
  .B({ S441 }),
  .Y({ S443 })
);
NAND #() 
NAND_78_ (
  .A({ S429 }),
  .B({ S442 }),
  .Y({ S444 })
);
NOR #() 
NOR_65_ (
  .A({ S435 }),
  .B({ S444 }),
  .Y({ S445 })
);
NAND #() 
NAND_79_ (
  .A({ S429 }),
  .B({ S443 }),
  .Y({ S446 })
);
NAND #() 
NAND_80_ (
  .A({ datapath_theregisterfile_memtrf_238 }),
  .B({ S436 }),
  .Y({ S447 })
);
NAND #() 
NAND_81_ (
  .A({ datapath_theregisterfile_memtrf_254 }),
  .B({ S435 }),
  .Y({ S448 })
);
NAND #() 
NAND_82_ (
  .A({ S447 }),
  .B({ S448 }),
  .Y({ S449 })
);
NAND #() 
NAND_83_ (
  .A({ S422 }),
  .B({ S449 }),
  .Y({ S450 })
);
NAND #() 
NAND_84_ (
  .A({ datapath_theregisterfile_memtrf_174 }),
  .B({ S436 }),
  .Y({ S451 })
);
NAND #() 
NAND_85_ (
  .A({ datapath_theregisterfile_memtrf_190 }),
  .B({ S435 }),
  .Y({ S452 })
);
NAND #() 
NAND_86_ (
  .A({ S451 }),
  .B({ S452 }),
  .Y({ S453 })
);
NAND #() 
NAND_87_ (
  .A({ S423 }),
  .B({ S453 }),
  .Y({ S454 })
);
NAND #() 
NAND_88_ (
  .A({ S450 }),
  .B({ S454 }),
  .Y({ S455 })
);
NOR #() 
NOR_66_ (
  .A({ datapath_theregisterfile_memtrf_222 }),
  .B({ S423 }),
  .Y({ S456 })
);
NAND #() 
NAND_89_ (
  .A({ S7564 }),
  .B({ S423 }),
  .Y({ S457 })
);
NAND #() 
NAND_90_ (
  .A({ S435 }),
  .B({ S457 }),
  .Y({ S458 })
);
NOR #() 
NOR_67_ (
  .A({ S456 }),
  .B({ S458 }),
  .Y({ S459 })
);
NOR #() 
NOR_68_ (
  .A({ datapath_theregisterfile_memtrf_142 }),
  .B({ S422 }),
  .Y({ S460 })
);
NAND #() 
NAND_91_ (
  .A({ S7772 }),
  .B({ S422 }),
  .Y({ S461 })
);
NAND #() 
NAND_92_ (
  .A({ S436 }),
  .B({ S461 }),
  .Y({ S462 })
);
NOR #() 
NOR_69_ (
  .A({ S460 }),
  .B({ S462 }),
  .Y({ S463 })
);
NOR #() 
NOR_70_ (
  .A({ S459 }),
  .B({ S463 }),
  .Y({ S464 })
);
NAND #() 
NAND_93_ (
  .A({ S442 }),
  .B({ S464 }),
  .Y({ S465 })
);
NOR #() 
NOR_71_ (
  .A({ S442 }),
  .B({ S455 }),
  .Y({ S466 })
);
NAND #() 
NAND_94_ (
  .A({ S428 }),
  .B({ S465 }),
  .Y({ S467 })
);
NOR #() 
NOR_72_ (
  .A({ S466 }),
  .B({ S467 }),
  .Y({ S468 })
);
NAND #() 
NAND_95_ (
  .A({ datapath_theregisterfile_memtrf_62 }),
  .B({ S435 }),
  .Y({ S469 })
);
NAND #() 
NAND_96_ (
  .A({ datapath_theregisterfile_memtrf_46 }),
  .B({ S436 }),
  .Y({ S470 })
);
NAND #() 
NAND_97_ (
  .A({ S469 }),
  .B({ S470 }),
  .Y({ S471 })
);
NAND #() 
NAND_98_ (
  .A({ S441 }),
  .B({ S471 }),
  .Y({ S472 })
);
NAND #() 
NAND_99_ (
  .A({ datapath_theregisterfile_memtrf_30 }),
  .B({ S435 }),
  .Y({ S473 })
);
NAND #() 
NAND_100_ (
  .A({ datapath_theregisterfile_memtrf_14 }),
  .B({ S436 }),
  .Y({ S474 })
);
NAND #() 
NAND_101_ (
  .A({ S473 }),
  .B({ S474 }),
  .Y({ S475 })
);
NAND #() 
NAND_102_ (
  .A({ S442 }),
  .B({ S475 }),
  .Y({ S476 })
);
NAND #() 
NAND_103_ (
  .A({ S472 }),
  .B({ S476 }),
  .Y({ S477 })
);
NAND #() 
NAND_104_ (
  .A({ S429 }),
  .B({ S477 }),
  .Y({ S478 })
);
NOR #() 
NOR_73_ (
  .A({ S423 }),
  .B({ S428 }),
  .Y({ S479 })
);
NAND #() 
NAND_105_ (
  .A({ datapath_theregisterfile_memtrf_126 }),
  .B({ S435 }),
  .Y({ S480 })
);
NAND #() 
NAND_106_ (
  .A({ datapath_theregisterfile_memtrf_110 }),
  .B({ S436 }),
  .Y({ S481 })
);
NAND #() 
NAND_107_ (
  .A({ S480 }),
  .B({ S481 }),
  .Y({ S482 })
);
NAND #() 
NAND_108_ (
  .A({ S441 }),
  .B({ S482 }),
  .Y({ S483 })
);
NAND #() 
NAND_109_ (
  .A({ datapath_theregisterfile_memtrf_94 }),
  .B({ S435 }),
  .Y({ S484 })
);
NAND #() 
NAND_110_ (
  .A({ datapath_theregisterfile_memtrf_78 }),
  .B({ S436 }),
  .Y({ S485 })
);
NAND #() 
NAND_111_ (
  .A({ S484 }),
  .B({ S485 }),
  .Y({ S486 })
);
NAND #() 
NAND_112_ (
  .A({ S442 }),
  .B({ S486 }),
  .Y({ S487 })
);
NAND #() 
NAND_113_ (
  .A({ S483 }),
  .B({ S487 }),
  .Y({ S488 })
);
NAND #() 
NAND_114_ (
  .A({ S479 }),
  .B({ S488 }),
  .Y({ S489 })
);
NAND #() 
NAND_115_ (
  .A({ S478 }),
  .B({ S489 }),
  .Y({ S490 })
);
NOR #() 
NOR_74_ (
  .A({ S468 }),
  .B({ S490 }),
  .Y({ S491 })
);
NOR #() 
NOR_75_ (
  .A({ S445 }),
  .B({ S491 }),
  .Y({ datapath_addsubunit_in1_14 })
);
NOT #() 
NOT_117_ (
  .A({ datapath_addsubunit_in1_14 }),
  .Y({ S492 })
);
NAND #() 
NAND_116_ (
  .A({ S366 }),
  .B({ S368 }),
  .Y({ S493 })
);
NOR #() 
NOR_76_ (
  .A({ S356 }),
  .B({ S361 }),
  .Y({ S494 })
);
NAND #() 
NAND_117_ (
  .A({ S8375 }),
  .B({ S494 }),
  .Y({ S495 })
);
NAND #() 
NAND_118_ (
  .A({ S493 }),
  .B({ S495 }),
  .Y({ S496 })
);
NAND #() 
NAND_119_ (
  .A({ datapath_addsubunit_in1_14 }),
  .B({ S496 }),
  .Y({ S497 })
);
NAND #() 
NAND_120_ (
  .A({ S372 }),
  .B({ S497 }),
  .Y({ S498 })
);
NAND #() 
NAND_121_ (
  .A({ datapath_muxmem_in2_14 }),
  .B({ S498 }),
  .Y({ S499 })
);
NOT #() 
NOT_118_ (
  .A({ S499 }),
  .Y({ S500 })
);
NOR #() 
NOR_77_ (
  .A({ datapath_muxmem_in2_14 }),
  .B({ S498 }),
  .Y({ S501 })
);
NOR #() 
NOR_78_ (
  .A({ S500 }),
  .B({ S501 }),
  .Y({ S502 })
);
NAND #() 
NAND_122_ (
  .A({ datapath_theregisterfile_memtrf_237 }),
  .B({ S436 }),
  .Y({ S503 })
);
NAND #() 
NAND_123_ (
  .A({ datapath_theregisterfile_memtrf_253 }),
  .B({ S435 }),
  .Y({ S504 })
);
NAND #() 
NAND_124_ (
  .A({ S503 }),
  .B({ S504 }),
  .Y({ S505 })
);
NAND #() 
NAND_125_ (
  .A({ S422 }),
  .B({ S505 }),
  .Y({ S506 })
);
NAND #() 
NAND_126_ (
  .A({ datapath_theregisterfile_memtrf_173 }),
  .B({ S436 }),
  .Y({ S507 })
);
NAND #() 
NAND_127_ (
  .A({ datapath_theregisterfile_memtrf_189 }),
  .B({ S435 }),
  .Y({ S508 })
);
NAND #() 
NAND_128_ (
  .A({ S507 }),
  .B({ S508 }),
  .Y({ S509 })
);
NAND #() 
NAND_129_ (
  .A({ S423 }),
  .B({ S509 }),
  .Y({ S510 })
);
NAND #() 
NAND_130_ (
  .A({ S506 }),
  .B({ S510 }),
  .Y({ S511 })
);
NOR #() 
NOR_79_ (
  .A({ datapath_theregisterfile_memtrf_221 }),
  .B({ S423 }),
  .Y({ S512 })
);
NAND #() 
NAND_131_ (
  .A({ S7553 }),
  .B({ S423 }),
  .Y({ S513 })
);
NAND #() 
NAND_132_ (
  .A({ S435 }),
  .B({ S513 }),
  .Y({ S514 })
);
NOR #() 
NOR_80_ (
  .A({ S512 }),
  .B({ S514 }),
  .Y({ S515 })
);
NOR #() 
NOR_81_ (
  .A({ datapath_theregisterfile_memtrf_141 }),
  .B({ S422 }),
  .Y({ S516 })
);
NAND #() 
NAND_133_ (
  .A({ S7761 }),
  .B({ S422 }),
  .Y({ S517 })
);
NAND #() 
NAND_134_ (
  .A({ S436 }),
  .B({ S517 }),
  .Y({ S518 })
);
NOR #() 
NOR_82_ (
  .A({ S516 }),
  .B({ S518 }),
  .Y({ S519 })
);
NOR #() 
NOR_83_ (
  .A({ S515 }),
  .B({ S519 }),
  .Y({ S520 })
);
NAND #() 
NAND_135_ (
  .A({ S442 }),
  .B({ S520 }),
  .Y({ S521 })
);
NOR #() 
NOR_84_ (
  .A({ S442 }),
  .B({ S511 }),
  .Y({ S522 })
);
NAND #() 
NAND_136_ (
  .A({ S428 }),
  .B({ S521 }),
  .Y({ S523 })
);
NOR #() 
NOR_85_ (
  .A({ S522 }),
  .B({ S523 }),
  .Y({ S524 })
);
NAND #() 
NAND_137_ (
  .A({ datapath_theregisterfile_memtrf_61 }),
  .B({ S435 }),
  .Y({ S525 })
);
NAND #() 
NAND_138_ (
  .A({ datapath_theregisterfile_memtrf_45 }),
  .B({ S436 }),
  .Y({ S526 })
);
NAND #() 
NAND_139_ (
  .A({ S525 }),
  .B({ S526 }),
  .Y({ S527 })
);
NAND #() 
NAND_140_ (
  .A({ S441 }),
  .B({ S527 }),
  .Y({ S528 })
);
NAND #() 
NAND_141_ (
  .A({ datapath_theregisterfile_memtrf_29 }),
  .B({ S435 }),
  .Y({ S529 })
);
NAND #() 
NAND_142_ (
  .A({ datapath_theregisterfile_memtrf_13 }),
  .B({ S436 }),
  .Y({ S530 })
);
NAND #() 
NAND_143_ (
  .A({ S529 }),
  .B({ S530 }),
  .Y({ S531 })
);
NAND #() 
NAND_144_ (
  .A({ S442 }),
  .B({ S531 }),
  .Y({ S532 })
);
NAND #() 
NAND_145_ (
  .A({ S528 }),
  .B({ S532 }),
  .Y({ S533 })
);
NAND #() 
NAND_146_ (
  .A({ S429 }),
  .B({ S533 }),
  .Y({ S534 })
);
NAND #() 
NAND_147_ (
  .A({ datapath_theregisterfile_memtrf_125 }),
  .B({ S435 }),
  .Y({ S535 })
);
NAND #() 
NAND_148_ (
  .A({ datapath_theregisterfile_memtrf_109 }),
  .B({ S436 }),
  .Y({ S536 })
);
NAND #() 
NAND_149_ (
  .A({ S535 }),
  .B({ S536 }),
  .Y({ S537 })
);
NAND #() 
NAND_150_ (
  .A({ S441 }),
  .B({ S537 }),
  .Y({ S538 })
);
NAND #() 
NAND_151_ (
  .A({ datapath_theregisterfile_memtrf_93 }),
  .B({ S435 }),
  .Y({ S539 })
);
NAND #() 
NAND_152_ (
  .A({ datapath_theregisterfile_memtrf_77 }),
  .B({ S436 }),
  .Y({ S540 })
);
NAND #() 
NAND_153_ (
  .A({ S539 }),
  .B({ S540 }),
  .Y({ S541 })
);
NAND #() 
NAND_154_ (
  .A({ S442 }),
  .B({ S541 }),
  .Y({ S542 })
);
NAND #() 
NAND_155_ (
  .A({ S538 }),
  .B({ S542 }),
  .Y({ S543 })
);
NAND #() 
NAND_156_ (
  .A({ S479 }),
  .B({ S543 }),
  .Y({ S544 })
);
NOT #() 
NOT_119_ (
  .A({ S544 }),
  .Y({ S545 })
);
NOR #() 
NOR_86_ (
  .A({ S524 }),
  .B({ S545 }),
  .Y({ S546 })
);
NAND #() 
NAND_157_ (
  .A({ S534 }),
  .B({ S546 }),
  .Y({ S547 })
);
NAND #() 
NAND_158_ (
  .A({ S446 }),
  .B({ S547 }),
  .Y({ S548 })
);
NOT #() 
NOT_120_ (
  .A({ S548 }),
  .Y({ datapath_addsubunit_in1_13 })
);
NAND #() 
NAND_159_ (
  .A({ S496 }),
  .B({ datapath_addsubunit_in1_13 }),
  .Y({ S549 })
);
NAND #() 
NAND_160_ (
  .A({ S372 }),
  .B({ S549 }),
  .Y({ S550 })
);
NOT #() 
NOT_121_ (
  .A({ S550 }),
  .Y({ S551 })
);
NOR #() 
NOR_87_ (
  .A({ datapath_muxmem_in2_13 }),
  .B({ S550 }),
  .Y({ S552 })
);
NOR #() 
NOR_88_ (
  .A({ S8000 }),
  .B({ S551 }),
  .Y({ S553 })
);
NOR #() 
NOR_89_ (
  .A({ datapath_theregisterfile_memtrf_172 }),
  .B({ S422 }),
  .Y({ S554 })
);
NOR #() 
NOR_90_ (
  .A({ datapath_theregisterfile_memtrf_236 }),
  .B({ S423 }),
  .Y({ S555 })
);
NOR #() 
NOR_91_ (
  .A({ S554 }),
  .B({ S555 }),
  .Y({ S556 })
);
NAND #() 
NAND_161_ (
  .A({ S436 }),
  .B({ S556 }),
  .Y({ S557 })
);
NOR #() 
NOR_92_ (
  .A({ datapath_theregisterfile_memtrf_252 }),
  .B({ S423 }),
  .Y({ S558 })
);
NAND #() 
NAND_162_ (
  .A({ S7651 }),
  .B({ S423 }),
  .Y({ S559 })
);
NAND #() 
NAND_163_ (
  .A({ S435 }),
  .B({ S559 }),
  .Y({ S560 })
);
NOR #() 
NOR_93_ (
  .A({ S558 }),
  .B({ S560 }),
  .Y({ S561 })
);
NAND #() 
NAND_164_ (
  .A({ datapath_theregisterfile_memtrf_204 }),
  .B({ S436 }),
  .Y({ S562 })
);
NAND #() 
NAND_165_ (
  .A({ datapath_theregisterfile_memtrf_220 }),
  .B({ S435 }),
  .Y({ S563 })
);
NAND #() 
NAND_166_ (
  .A({ S562 }),
  .B({ S563 }),
  .Y({ S564 })
);
NAND #() 
NAND_167_ (
  .A({ S422 }),
  .B({ S564 }),
  .Y({ S565 })
);
NAND #() 
NAND_168_ (
  .A({ datapath_theregisterfile_memtrf_140 }),
  .B({ S436 }),
  .Y({ S566 })
);
NAND #() 
NAND_169_ (
  .A({ datapath_theregisterfile_memtrf_156 }),
  .B({ S435 }),
  .Y({ S567 })
);
NAND #() 
NAND_170_ (
  .A({ S566 }),
  .B({ S567 }),
  .Y({ S568 })
);
NAND #() 
NAND_171_ (
  .A({ S423 }),
  .B({ S568 }),
  .Y({ S569 })
);
NAND #() 
NAND_172_ (
  .A({ S565 }),
  .B({ S569 }),
  .Y({ S570 })
);
NOR #() 
NOR_94_ (
  .A({ S441 }),
  .B({ S570 }),
  .Y({ S571 })
);
NOR #() 
NOR_95_ (
  .A({ S442 }),
  .B({ S561 }),
  .Y({ S572 })
);
NAND #() 
NAND_173_ (
  .A({ S557 }),
  .B({ S572 }),
  .Y({ S573 })
);
NAND #() 
NAND_174_ (
  .A({ S428 }),
  .B({ S573 }),
  .Y({ S574 })
);
NOR #() 
NOR_96_ (
  .A({ S571 }),
  .B({ S574 }),
  .Y({ S575 })
);
NAND #() 
NAND_175_ (
  .A({ datapath_theregisterfile_memtrf_124 }),
  .B({ S435 }),
  .Y({ S576 })
);
NAND #() 
NAND_176_ (
  .A({ datapath_theregisterfile_memtrf_108 }),
  .B({ S436 }),
  .Y({ S577 })
);
NAND #() 
NAND_177_ (
  .A({ S576 }),
  .B({ S577 }),
  .Y({ S578 })
);
NAND #() 
NAND_178_ (
  .A({ S441 }),
  .B({ S578 }),
  .Y({ S579 })
);
NAND #() 
NAND_179_ (
  .A({ datapath_theregisterfile_memtrf_92 }),
  .B({ S435 }),
  .Y({ S580 })
);
NAND #() 
NAND_180_ (
  .A({ datapath_theregisterfile_memtrf_76 }),
  .B({ S436 }),
  .Y({ S581 })
);
NAND #() 
NAND_181_ (
  .A({ S580 }),
  .B({ S581 }),
  .Y({ S582 })
);
NAND #() 
NAND_182_ (
  .A({ S442 }),
  .B({ S582 }),
  .Y({ S583 })
);
NAND #() 
NAND_183_ (
  .A({ S579 }),
  .B({ S583 }),
  .Y({ S584 })
);
NAND #() 
NAND_184_ (
  .A({ S479 }),
  .B({ S584 }),
  .Y({ S585 })
);
NAND #() 
NAND_185_ (
  .A({ datapath_theregisterfile_memtrf_60 }),
  .B({ S435 }),
  .Y({ S586 })
);
NAND #() 
NAND_186_ (
  .A({ datapath_theregisterfile_memtrf_44 }),
  .B({ S436 }),
  .Y({ S587 })
);
NAND #() 
NAND_187_ (
  .A({ S586 }),
  .B({ S587 }),
  .Y({ S588 })
);
NAND #() 
NAND_188_ (
  .A({ S441 }),
  .B({ S588 }),
  .Y({ S589 })
);
NAND #() 
NAND_189_ (
  .A({ datapath_theregisterfile_memtrf_28 }),
  .B({ S435 }),
  .Y({ S590 })
);
NAND #() 
NAND_190_ (
  .A({ datapath_theregisterfile_memtrf_12 }),
  .B({ S436 }),
  .Y({ S591 })
);
NAND #() 
NAND_191_ (
  .A({ S590 }),
  .B({ S591 }),
  .Y({ S592 })
);
NAND #() 
NAND_192_ (
  .A({ S442 }),
  .B({ S592 }),
  .Y({ S593 })
);
NAND #() 
NAND_193_ (
  .A({ S589 }),
  .B({ S593 }),
  .Y({ S594 })
);
NAND #() 
NAND_194_ (
  .A({ S429 }),
  .B({ S594 }),
  .Y({ S595 })
);
NOT #() 
NOT_122_ (
  .A({ S595 }),
  .Y({ S596 })
);
NOR #() 
NOR_97_ (
  .A({ S575 }),
  .B({ S596 }),
  .Y({ S597 })
);
NAND #() 
NAND_195_ (
  .A({ S585 }),
  .B({ S597 }),
  .Y({ S598 })
);
NAND #() 
NAND_196_ (
  .A({ S446 }),
  .B({ S598 }),
  .Y({ S599 })
);
NOT #() 
NOT_123_ (
  .A({ S599 }),
  .Y({ datapath_addsubunit_in1_12 })
);
NAND #() 
NAND_197_ (
  .A({ S496 }),
  .B({ datapath_addsubunit_in1_12 }),
  .Y({ S600 })
);
NAND #() 
NAND_198_ (
  .A({ S372 }),
  .B({ S600 }),
  .Y({ S601 })
);
NAND #() 
NAND_199_ (
  .A({ datapath_muxmem_in2_12 }),
  .B({ S601 }),
  .Y({ S602 })
);
NOT #() 
NOT_124_ (
  .A({ S602 }),
  .Y({ S603 })
);
NOR #() 
NOR_98_ (
  .A({ datapath_muxmem_in2_12 }),
  .B({ S601 }),
  .Y({ S604 })
);
NOR #() 
NOR_99_ (
  .A({ S603 }),
  .B({ S604 }),
  .Y({ S605 })
);
NOR #() 
NOR_100_ (
  .A({ datapath_theregisterfile_memtrf_171 }),
  .B({ S422 }),
  .Y({ S606 })
);
NOR #() 
NOR_101_ (
  .A({ datapath_theregisterfile_memtrf_235 }),
  .B({ S423 }),
  .Y({ S607 })
);
NOR #() 
NOR_102_ (
  .A({ S606 }),
  .B({ S607 }),
  .Y({ S608 })
);
NAND #() 
NAND_200_ (
  .A({ S436 }),
  .B({ S608 }),
  .Y({ S609 })
);
NOR #() 
NOR_103_ (
  .A({ datapath_theregisterfile_memtrf_251 }),
  .B({ S423 }),
  .Y({ S610 })
);
NAND #() 
NAND_201_ (
  .A({ S7640 }),
  .B({ S423 }),
  .Y({ S611 })
);
NAND #() 
NAND_202_ (
  .A({ S435 }),
  .B({ S611 }),
  .Y({ S612 })
);
NOR #() 
NOR_104_ (
  .A({ S610 }),
  .B({ S612 }),
  .Y({ S613 })
);
NAND #() 
NAND_203_ (
  .A({ datapath_theregisterfile_memtrf_203 }),
  .B({ S436 }),
  .Y({ S614 })
);
NAND #() 
NAND_204_ (
  .A({ datapath_theregisterfile_memtrf_219 }),
  .B({ S435 }),
  .Y({ S615 })
);
NAND #() 
NAND_205_ (
  .A({ S614 }),
  .B({ S615 }),
  .Y({ S616 })
);
NAND #() 
NAND_206_ (
  .A({ S422 }),
  .B({ S616 }),
  .Y({ S617 })
);
NAND #() 
NAND_207_ (
  .A({ datapath_theregisterfile_memtrf_139 }),
  .B({ S436 }),
  .Y({ S618 })
);
NAND #() 
NAND_208_ (
  .A({ datapath_theregisterfile_memtrf_155 }),
  .B({ S435 }),
  .Y({ S619 })
);
NAND #() 
NAND_209_ (
  .A({ S618 }),
  .B({ S619 }),
  .Y({ S620 })
);
NAND #() 
NAND_210_ (
  .A({ S423 }),
  .B({ S620 }),
  .Y({ S621 })
);
NAND #() 
NAND_211_ (
  .A({ S617 }),
  .B({ S621 }),
  .Y({ S622 })
);
NOR #() 
NOR_105_ (
  .A({ S441 }),
  .B({ S622 }),
  .Y({ S623 })
);
NOR #() 
NOR_106_ (
  .A({ S442 }),
  .B({ S613 }),
  .Y({ S624 })
);
NAND #() 
NAND_212_ (
  .A({ S609 }),
  .B({ S624 }),
  .Y({ S625 })
);
NAND #() 
NAND_213_ (
  .A({ S428 }),
  .B({ S625 }),
  .Y({ S626 })
);
NOR #() 
NOR_107_ (
  .A({ S623 }),
  .B({ S626 }),
  .Y({ S627 })
);
NAND #() 
NAND_214_ (
  .A({ datapath_theregisterfile_memtrf_59 }),
  .B({ S435 }),
  .Y({ S628 })
);
NAND #() 
NAND_215_ (
  .A({ datapath_theregisterfile_memtrf_43 }),
  .B({ S436 }),
  .Y({ S629 })
);
NAND #() 
NAND_216_ (
  .A({ S628 }),
  .B({ S629 }),
  .Y({ S630 })
);
NAND #() 
NAND_217_ (
  .A({ S441 }),
  .B({ S630 }),
  .Y({ S631 })
);
NAND #() 
NAND_218_ (
  .A({ datapath_theregisterfile_memtrf_27 }),
  .B({ S435 }),
  .Y({ S632 })
);
NAND #() 
NAND_219_ (
  .A({ datapath_theregisterfile_memtrf_11 }),
  .B({ S436 }),
  .Y({ S633 })
);
NAND #() 
NAND_220_ (
  .A({ S632 }),
  .B({ S633 }),
  .Y({ S634 })
);
NAND #() 
NAND_221_ (
  .A({ S442 }),
  .B({ S634 }),
  .Y({ S635 })
);
NAND #() 
NAND_222_ (
  .A({ S631 }),
  .B({ S635 }),
  .Y({ S636 })
);
NAND #() 
NAND_223_ (
  .A({ S429 }),
  .B({ S636 }),
  .Y({ S637 })
);
NAND #() 
NAND_224_ (
  .A({ datapath_theregisterfile_memtrf_123 }),
  .B({ S435 }),
  .Y({ S638 })
);
NAND #() 
NAND_225_ (
  .A({ datapath_theregisterfile_memtrf_107 }),
  .B({ S436 }),
  .Y({ S639 })
);
NAND #() 
NAND_226_ (
  .A({ S638 }),
  .B({ S639 }),
  .Y({ S640 })
);
NAND #() 
NAND_227_ (
  .A({ S441 }),
  .B({ S640 }),
  .Y({ S641 })
);
NAND #() 
NAND_228_ (
  .A({ datapath_theregisterfile_memtrf_91 }),
  .B({ S435 }),
  .Y({ S642 })
);
NAND #() 
NAND_229_ (
  .A({ datapath_theregisterfile_memtrf_75 }),
  .B({ S436 }),
  .Y({ S643 })
);
NAND #() 
NAND_230_ (
  .A({ S642 }),
  .B({ S643 }),
  .Y({ S644 })
);
NAND #() 
NAND_231_ (
  .A({ S442 }),
  .B({ S644 }),
  .Y({ S645 })
);
NAND #() 
NAND_232_ (
  .A({ S641 }),
  .B({ S645 }),
  .Y({ S646 })
);
NAND #() 
NAND_233_ (
  .A({ S479 }),
  .B({ S646 }),
  .Y({ S647 })
);
NOT #() 
NOT_125_ (
  .A({ S647 }),
  .Y({ S648 })
);
NOR #() 
NOR_108_ (
  .A({ S627 }),
  .B({ S648 }),
  .Y({ S649 })
);
NAND #() 
NAND_234_ (
  .A({ S637 }),
  .B({ S649 }),
  .Y({ S650 })
);
NAND #() 
NAND_235_ (
  .A({ S446 }),
  .B({ S650 }),
  .Y({ S651 })
);
NOT #() 
NOT_126_ (
  .A({ S651 }),
  .Y({ datapath_addsubunit_in1_11 })
);
NAND #() 
NAND_236_ (
  .A({ S496 }),
  .B({ datapath_addsubunit_in1_11 }),
  .Y({ S652 })
);
NAND #() 
NAND_237_ (
  .A({ S372 }),
  .B({ S652 }),
  .Y({ S653 })
);
NOT #() 
NOT_127_ (
  .A({ S653 }),
  .Y({ S654 })
);
NOR #() 
NOR_109_ (
  .A({ S7978 }),
  .B({ S654 }),
  .Y({ S655 })
);
NOR #() 
NOR_110_ (
  .A({ datapath_muxmem_in2_11 }),
  .B({ S653 }),
  .Y({ S656 })
);
NOR #() 
NOR_111_ (
  .A({ datapath_theregisterfile_memtrf_170 }),
  .B({ S422 }),
  .Y({ S657 })
);
NOR #() 
NOR_112_ (
  .A({ datapath_theregisterfile_memtrf_234 }),
  .B({ S423 }),
  .Y({ S658 })
);
NOR #() 
NOR_113_ (
  .A({ S657 }),
  .B({ S658 }),
  .Y({ S659 })
);
NAND #() 
NAND_238_ (
  .A({ S436 }),
  .B({ S659 }),
  .Y({ S660 })
);
NOR #() 
NOR_114_ (
  .A({ datapath_theregisterfile_memtrf_250 }),
  .B({ S423 }),
  .Y({ S661 })
);
NAND #() 
NAND_239_ (
  .A({ S7629 }),
  .B({ S423 }),
  .Y({ S662 })
);
NAND #() 
NAND_240_ (
  .A({ S435 }),
  .B({ S662 }),
  .Y({ S663 })
);
NOR #() 
NOR_115_ (
  .A({ S661 }),
  .B({ S663 }),
  .Y({ S664 })
);
NAND #() 
NAND_241_ (
  .A({ datapath_theregisterfile_memtrf_202 }),
  .B({ S436 }),
  .Y({ S665 })
);
NAND #() 
NAND_242_ (
  .A({ datapath_theregisterfile_memtrf_218 }),
  .B({ S435 }),
  .Y({ S666 })
);
NAND #() 
NAND_243_ (
  .A({ S665 }),
  .B({ S666 }),
  .Y({ S667 })
);
NAND #() 
NAND_244_ (
  .A({ S422 }),
  .B({ S667 }),
  .Y({ S668 })
);
NAND #() 
NAND_245_ (
  .A({ datapath_theregisterfile_memtrf_138 }),
  .B({ S436 }),
  .Y({ S669 })
);
NAND #() 
NAND_246_ (
  .A({ datapath_theregisterfile_memtrf_154 }),
  .B({ S435 }),
  .Y({ S670 })
);
NAND #() 
NAND_247_ (
  .A({ S669 }),
  .B({ S670 }),
  .Y({ S671 })
);
NAND #() 
NAND_248_ (
  .A({ S423 }),
  .B({ S671 }),
  .Y({ S672 })
);
NAND #() 
NAND_249_ (
  .A({ S668 }),
  .B({ S672 }),
  .Y({ S673 })
);
NOR #() 
NOR_116_ (
  .A({ S441 }),
  .B({ S673 }),
  .Y({ S674 })
);
NOR #() 
NOR_117_ (
  .A({ S442 }),
  .B({ S664 }),
  .Y({ S675 })
);
NAND #() 
NAND_250_ (
  .A({ S660 }),
  .B({ S675 }),
  .Y({ S676 })
);
NAND #() 
NAND_251_ (
  .A({ S428 }),
  .B({ S676 }),
  .Y({ S677 })
);
NOR #() 
NOR_118_ (
  .A({ S674 }),
  .B({ S677 }),
  .Y({ S678 })
);
NAND #() 
NAND_252_ (
  .A({ datapath_theregisterfile_memtrf_122 }),
  .B({ S435 }),
  .Y({ S679 })
);
NAND #() 
NAND_253_ (
  .A({ datapath_theregisterfile_memtrf_106 }),
  .B({ S436 }),
  .Y({ S680 })
);
NAND #() 
NAND_254_ (
  .A({ S679 }),
  .B({ S680 }),
  .Y({ S681 })
);
NAND #() 
NAND_255_ (
  .A({ S441 }),
  .B({ S681 }),
  .Y({ S682 })
);
NAND #() 
NAND_256_ (
  .A({ datapath_theregisterfile_memtrf_90 }),
  .B({ S435 }),
  .Y({ S683 })
);
NAND #() 
NAND_257_ (
  .A({ datapath_theregisterfile_memtrf_74 }),
  .B({ S436 }),
  .Y({ S684 })
);
NAND #() 
NAND_258_ (
  .A({ S683 }),
  .B({ S684 }),
  .Y({ S685 })
);
NAND #() 
NAND_259_ (
  .A({ S442 }),
  .B({ S685 }),
  .Y({ S686 })
);
NAND #() 
NAND_260_ (
  .A({ S682 }),
  .B({ S686 }),
  .Y({ S687 })
);
NAND #() 
NAND_261_ (
  .A({ S479 }),
  .B({ S687 }),
  .Y({ S688 })
);
NAND #() 
NAND_262_ (
  .A({ datapath_theregisterfile_memtrf_58 }),
  .B({ S435 }),
  .Y({ S689 })
);
NAND #() 
NAND_263_ (
  .A({ datapath_theregisterfile_memtrf_42 }),
  .B({ S436 }),
  .Y({ S690 })
);
NAND #() 
NAND_264_ (
  .A({ S689 }),
  .B({ S690 }),
  .Y({ S691 })
);
NAND #() 
NAND_265_ (
  .A({ S441 }),
  .B({ S691 }),
  .Y({ S692 })
);
NAND #() 
NAND_266_ (
  .A({ datapath_theregisterfile_memtrf_26 }),
  .B({ S435 }),
  .Y({ S693 })
);
NAND #() 
NAND_267_ (
  .A({ datapath_theregisterfile_memtrf_10 }),
  .B({ S436 }),
  .Y({ S694 })
);
NAND #() 
NAND_268_ (
  .A({ S693 }),
  .B({ S694 }),
  .Y({ S695 })
);
NAND #() 
NAND_269_ (
  .A({ S442 }),
  .B({ S695 }),
  .Y({ S696 })
);
NAND #() 
NAND_270_ (
  .A({ S692 }),
  .B({ S696 }),
  .Y({ S697 })
);
NAND #() 
NAND_271_ (
  .A({ S429 }),
  .B({ S697 }),
  .Y({ S698 })
);
NOT #() 
NOT_128_ (
  .A({ S698 }),
  .Y({ S699 })
);
NOR #() 
NOR_119_ (
  .A({ S678 }),
  .B({ S699 }),
  .Y({ S700 })
);
NAND #() 
NAND_272_ (
  .A({ S688 }),
  .B({ S700 }),
  .Y({ S701 })
);
NAND #() 
NAND_273_ (
  .A({ S446 }),
  .B({ S701 }),
  .Y({ S702 })
);
NOT #() 
NOT_129_ (
  .A({ S702 }),
  .Y({ datapath_addsubunit_in1_10 })
);
NAND #() 
NAND_274_ (
  .A({ S496 }),
  .B({ datapath_addsubunit_in1_10 }),
  .Y({ S703 })
);
NAND #() 
NAND_275_ (
  .A({ S372 }),
  .B({ S703 }),
  .Y({ S704 })
);
NAND #() 
NAND_276_ (
  .A({ datapath_muxmem_in2_10 }),
  .B({ S704 }),
  .Y({ S705 })
);
NOT #() 
NOT_130_ (
  .A({ S705 }),
  .Y({ S706 })
);
NOR #() 
NOR_120_ (
  .A({ datapath_muxmem_in2_10 }),
  .B({ S704 }),
  .Y({ S707 })
);
NOR #() 
NOR_121_ (
  .A({ S706 }),
  .B({ S707 }),
  .Y({ S708 })
);
NOR #() 
NOR_122_ (
  .A({ datapath_theregisterfile_memtrf_169 }),
  .B({ S422 }),
  .Y({ S709 })
);
NOR #() 
NOR_123_ (
  .A({ datapath_theregisterfile_memtrf_233 }),
  .B({ S423 }),
  .Y({ S710 })
);
NOR #() 
NOR_124_ (
  .A({ S709 }),
  .B({ S710 }),
  .Y({ S711 })
);
NAND #() 
NAND_277_ (
  .A({ S436 }),
  .B({ S711 }),
  .Y({ S712 })
);
NOR #() 
NOR_125_ (
  .A({ datapath_theregisterfile_memtrf_249 }),
  .B({ S423 }),
  .Y({ S713 })
);
NAND #() 
NAND_278_ (
  .A({ S7618 }),
  .B({ S423 }),
  .Y({ S714 })
);
NAND #() 
NAND_279_ (
  .A({ S435 }),
  .B({ S714 }),
  .Y({ S715 })
);
NOR #() 
NOR_126_ (
  .A({ S713 }),
  .B({ S715 }),
  .Y({ S716 })
);
NAND #() 
NAND_280_ (
  .A({ datapath_theregisterfile_memtrf_201 }),
  .B({ S436 }),
  .Y({ S717 })
);
NAND #() 
NAND_281_ (
  .A({ datapath_theregisterfile_memtrf_217 }),
  .B({ S435 }),
  .Y({ S718 })
);
NAND #() 
NAND_282_ (
  .A({ S717 }),
  .B({ S718 }),
  .Y({ S719 })
);
NAND #() 
NAND_283_ (
  .A({ S422 }),
  .B({ S719 }),
  .Y({ S720 })
);
NAND #() 
NAND_284_ (
  .A({ datapath_theregisterfile_memtrf_137 }),
  .B({ S436 }),
  .Y({ S721 })
);
NAND #() 
NAND_285_ (
  .A({ datapath_theregisterfile_memtrf_153 }),
  .B({ S435 }),
  .Y({ S722 })
);
NAND #() 
NAND_286_ (
  .A({ S721 }),
  .B({ S722 }),
  .Y({ S723 })
);
NAND #() 
NAND_287_ (
  .A({ S423 }),
  .B({ S723 }),
  .Y({ S724 })
);
NAND #() 
NAND_288_ (
  .A({ S720 }),
  .B({ S724 }),
  .Y({ S725 })
);
NOR #() 
NOR_127_ (
  .A({ S441 }),
  .B({ S725 }),
  .Y({ S726 })
);
NOR #() 
NOR_128_ (
  .A({ S442 }),
  .B({ S716 }),
  .Y({ S727 })
);
NAND #() 
NAND_289_ (
  .A({ S712 }),
  .B({ S727 }),
  .Y({ S728 })
);
NAND #() 
NAND_290_ (
  .A({ S428 }),
  .B({ S728 }),
  .Y({ S729 })
);
NOR #() 
NOR_129_ (
  .A({ S726 }),
  .B({ S729 }),
  .Y({ S730 })
);
NAND #() 
NAND_291_ (
  .A({ datapath_theregisterfile_memtrf_121 }),
  .B({ S435 }),
  .Y({ S731 })
);
NAND #() 
NAND_292_ (
  .A({ datapath_theregisterfile_memtrf_105 }),
  .B({ S436 }),
  .Y({ S732 })
);
NAND #() 
NAND_293_ (
  .A({ S731 }),
  .B({ S732 }),
  .Y({ S733 })
);
NAND #() 
NAND_294_ (
  .A({ S441 }),
  .B({ S733 }),
  .Y({ S734 })
);
NAND #() 
NAND_295_ (
  .A({ datapath_theregisterfile_memtrf_89 }),
  .B({ S435 }),
  .Y({ S735 })
);
NAND #() 
NAND_296_ (
  .A({ datapath_theregisterfile_memtrf_73 }),
  .B({ S436 }),
  .Y({ S736 })
);
NAND #() 
NAND_297_ (
  .A({ S735 }),
  .B({ S736 }),
  .Y({ S737 })
);
NAND #() 
NAND_298_ (
  .A({ S442 }),
  .B({ S737 }),
  .Y({ S738 })
);
NAND #() 
NAND_299_ (
  .A({ S734 }),
  .B({ S738 }),
  .Y({ S739 })
);
NAND #() 
NAND_300_ (
  .A({ S479 }),
  .B({ S739 }),
  .Y({ S740 })
);
NAND #() 
NAND_301_ (
  .A({ datapath_theregisterfile_memtrf_57 }),
  .B({ S435 }),
  .Y({ S741 })
);
NAND #() 
NAND_302_ (
  .A({ datapath_theregisterfile_memtrf_41 }),
  .B({ S436 }),
  .Y({ S742 })
);
NAND #() 
NAND_303_ (
  .A({ S741 }),
  .B({ S742 }),
  .Y({ S743 })
);
NAND #() 
NAND_304_ (
  .A({ S441 }),
  .B({ S743 }),
  .Y({ S744 })
);
NAND #() 
NAND_305_ (
  .A({ datapath_theregisterfile_memtrf_25 }),
  .B({ S435 }),
  .Y({ S745 })
);
NAND #() 
NAND_306_ (
  .A({ datapath_theregisterfile_memtrf_9 }),
  .B({ S436 }),
  .Y({ S746 })
);
NAND #() 
NAND_307_ (
  .A({ S745 }),
  .B({ S746 }),
  .Y({ S747 })
);
NAND #() 
NAND_308_ (
  .A({ S442 }),
  .B({ S747 }),
  .Y({ S748 })
);
NAND #() 
NAND_309_ (
  .A({ S744 }),
  .B({ S748 }),
  .Y({ S749 })
);
NAND #() 
NAND_310_ (
  .A({ S429 }),
  .B({ S749 }),
  .Y({ S750 })
);
NOT #() 
NOT_131_ (
  .A({ S750 }),
  .Y({ S751 })
);
NOR #() 
NOR_130_ (
  .A({ S730 }),
  .B({ S751 }),
  .Y({ S752 })
);
NAND #() 
NAND_311_ (
  .A({ S740 }),
  .B({ S752 }),
  .Y({ S753 })
);
NAND #() 
NAND_312_ (
  .A({ S446 }),
  .B({ S753 }),
  .Y({ S754 })
);
NOT #() 
NOT_132_ (
  .A({ S754 }),
  .Y({ datapath_addsubunit_in1_9 })
);
NAND #() 
NAND_313_ (
  .A({ S496 }),
  .B({ datapath_addsubunit_in1_9 }),
  .Y({ S755 })
);
NAND #() 
NAND_314_ (
  .A({ S372 }),
  .B({ S755 }),
  .Y({ S756 })
);
NOT #() 
NOT_133_ (
  .A({ S756 }),
  .Y({ S757 })
);
NOR #() 
NOR_131_ (
  .A({ S7957 }),
  .B({ S757 }),
  .Y({ S758 })
);
NOR #() 
NOR_132_ (
  .A({ datapath_muxmem_in2_9 }),
  .B({ S756 }),
  .Y({ S759 })
);
NOR #() 
NOR_133_ (
  .A({ datapath_theregisterfile_memtrf_168 }),
  .B({ S422 }),
  .Y({ S760 })
);
NOR #() 
NOR_134_ (
  .A({ datapath_theregisterfile_memtrf_232 }),
  .B({ S423 }),
  .Y({ S761 })
);
NOR #() 
NOR_135_ (
  .A({ S760 }),
  .B({ S761 }),
  .Y({ S762 })
);
NAND #() 
NAND_315_ (
  .A({ S436 }),
  .B({ S762 }),
  .Y({ S763 })
);
NOR #() 
NOR_136_ (
  .A({ datapath_theregisterfile_memtrf_248 }),
  .B({ S423 }),
  .Y({ S764 })
);
NAND #() 
NAND_316_ (
  .A({ S7607 }),
  .B({ S423 }),
  .Y({ S765 })
);
NAND #() 
NAND_317_ (
  .A({ S435 }),
  .B({ S765 }),
  .Y({ S766 })
);
NOR #() 
NOR_137_ (
  .A({ S764 }),
  .B({ S766 }),
  .Y({ S767 })
);
NAND #() 
NAND_318_ (
  .A({ datapath_theregisterfile_memtrf_200 }),
  .B({ S436 }),
  .Y({ S768 })
);
NAND #() 
NAND_319_ (
  .A({ datapath_theregisterfile_memtrf_216 }),
  .B({ S435 }),
  .Y({ S769 })
);
NAND #() 
NAND_320_ (
  .A({ S768 }),
  .B({ S769 }),
  .Y({ S770 })
);
NAND #() 
NAND_321_ (
  .A({ S422 }),
  .B({ S770 }),
  .Y({ S771 })
);
NAND #() 
NAND_322_ (
  .A({ datapath_theregisterfile_memtrf_136 }),
  .B({ S436 }),
  .Y({ S772 })
);
NAND #() 
NAND_323_ (
  .A({ datapath_theregisterfile_memtrf_152 }),
  .B({ S435 }),
  .Y({ S773 })
);
NAND #() 
NAND_324_ (
  .A({ S772 }),
  .B({ S773 }),
  .Y({ S774 })
);
NAND #() 
NAND_325_ (
  .A({ S423 }),
  .B({ S774 }),
  .Y({ S775 })
);
NAND #() 
NAND_326_ (
  .A({ S771 }),
  .B({ S775 }),
  .Y({ S776 })
);
NOR #() 
NOR_138_ (
  .A({ S441 }),
  .B({ S776 }),
  .Y({ S777 })
);
NOR #() 
NOR_139_ (
  .A({ S442 }),
  .B({ S767 }),
  .Y({ S778 })
);
NAND #() 
NAND_327_ (
  .A({ S763 }),
  .B({ S778 }),
  .Y({ S779 })
);
NAND #() 
NAND_328_ (
  .A({ S428 }),
  .B({ S779 }),
  .Y({ S780 })
);
NOR #() 
NOR_140_ (
  .A({ S777 }),
  .B({ S780 }),
  .Y({ S781 })
);
NAND #() 
NAND_329_ (
  .A({ datapath_theregisterfile_memtrf_120 }),
  .B({ S435 }),
  .Y({ S782 })
);
NAND #() 
NAND_330_ (
  .A({ datapath_theregisterfile_memtrf_104 }),
  .B({ S436 }),
  .Y({ S783 })
);
NAND #() 
NAND_331_ (
  .A({ S782 }),
  .B({ S783 }),
  .Y({ S784 })
);
NAND #() 
NAND_332_ (
  .A({ S441 }),
  .B({ S784 }),
  .Y({ S785 })
);
NAND #() 
NAND_333_ (
  .A({ datapath_theregisterfile_memtrf_88 }),
  .B({ S435 }),
  .Y({ S786 })
);
NAND #() 
NAND_334_ (
  .A({ datapath_theregisterfile_memtrf_72 }),
  .B({ S436 }),
  .Y({ S787 })
);
NAND #() 
NAND_335_ (
  .A({ S786 }),
  .B({ S787 }),
  .Y({ S788 })
);
NAND #() 
NAND_336_ (
  .A({ S442 }),
  .B({ S788 }),
  .Y({ S789 })
);
NAND #() 
NAND_337_ (
  .A({ S785 }),
  .B({ S789 }),
  .Y({ S790 })
);
NAND #() 
NAND_338_ (
  .A({ S479 }),
  .B({ S790 }),
  .Y({ S791 })
);
NAND #() 
NAND_339_ (
  .A({ datapath_theregisterfile_memtrf_56 }),
  .B({ S435 }),
  .Y({ S792 })
);
NAND #() 
NAND_340_ (
  .A({ datapath_theregisterfile_memtrf_40 }),
  .B({ S436 }),
  .Y({ S793 })
);
NAND #() 
NAND_341_ (
  .A({ S792 }),
  .B({ S793 }),
  .Y({ S794 })
);
NAND #() 
NAND_342_ (
  .A({ S441 }),
  .B({ S794 }),
  .Y({ S795 })
);
NAND #() 
NAND_343_ (
  .A({ datapath_theregisterfile_memtrf_24 }),
  .B({ S435 }),
  .Y({ S796 })
);
NAND #() 
NAND_344_ (
  .A({ datapath_theregisterfile_memtrf_8 }),
  .B({ S436 }),
  .Y({ S797 })
);
NAND #() 
NAND_345_ (
  .A({ S796 }),
  .B({ S797 }),
  .Y({ S798 })
);
NAND #() 
NAND_346_ (
  .A({ S442 }),
  .B({ S798 }),
  .Y({ S799 })
);
NAND #() 
NAND_347_ (
  .A({ S795 }),
  .B({ S799 }),
  .Y({ S800 })
);
NAND #() 
NAND_348_ (
  .A({ S429 }),
  .B({ S800 }),
  .Y({ S801 })
);
NOT #() 
NOT_134_ (
  .A({ S801 }),
  .Y({ S802 })
);
NOR #() 
NOR_141_ (
  .A({ S781 }),
  .B({ S802 }),
  .Y({ S803 })
);
NAND #() 
NAND_349_ (
  .A({ S791 }),
  .B({ S803 }),
  .Y({ S804 })
);
NAND #() 
NAND_350_ (
  .A({ S446 }),
  .B({ S804 }),
  .Y({ S805 })
);
NOT #() 
NOT_135_ (
  .A({ S805 }),
  .Y({ datapath_addsubunit_in1_8 })
);
NAND #() 
NAND_351_ (
  .A({ S496 }),
  .B({ datapath_addsubunit_in1_8 }),
  .Y({ S806 })
);
NAND #() 
NAND_352_ (
  .A({ S372 }),
  .B({ S806 }),
  .Y({ S807 })
);
NAND #() 
NAND_353_ (
  .A({ datapath_muxmem_in2_8 }),
  .B({ S807 }),
  .Y({ S808 })
);
NOT #() 
NOT_136_ (
  .A({ S808 }),
  .Y({ S809 })
);
NOR #() 
NOR_142_ (
  .A({ datapath_muxmem_in2_8 }),
  .B({ S807 }),
  .Y({ S810 })
);
NOR #() 
NOR_143_ (
  .A({ S809 }),
  .B({ S810 }),
  .Y({ S811 })
);
NAND #() 
NAND_354_ (
  .A({ S8349 }),
  .B({ S445 }),
  .Y({ S812 })
);
NAND #() 
NAND_355_ (
  .A({ datapath_theregisterfile_memtrf_183 }),
  .B({ S423 }),
  .Y({ S813 })
);
NAND #() 
NAND_356_ (
  .A({ datapath_theregisterfile_memtrf_247 }),
  .B({ S422 }),
  .Y({ S814 })
);
NAND #() 
NAND_357_ (
  .A({ S813 }),
  .B({ S814 }),
  .Y({ S815 })
);
NAND #() 
NAND_358_ (
  .A({ S435 }),
  .B({ S815 }),
  .Y({ S816 })
);
NOR #() 
NOR_144_ (
  .A({ datapath_theregisterfile_memtrf_167 }),
  .B({ S422 }),
  .Y({ S817 })
);
NOR #() 
NOR_145_ (
  .A({ datapath_theregisterfile_memtrf_231 }),
  .B({ S423 }),
  .Y({ S818 })
);
NOR #() 
NOR_146_ (
  .A({ S817 }),
  .B({ S818 }),
  .Y({ S819 })
);
NAND #() 
NAND_359_ (
  .A({ S436 }),
  .B({ S819 }),
  .Y({ S820 })
);
NAND #() 
NAND_360_ (
  .A({ S816 }),
  .B({ S820 }),
  .Y({ S821 })
);
NAND #() 
NAND_361_ (
  .A({ datapath_theregisterfile_memtrf_215 }),
  .B({ S422 }),
  .Y({ S822 })
);
NAND #() 
NAND_362_ (
  .A({ datapath_theregisterfile_memtrf_151 }),
  .B({ S423 }),
  .Y({ S823 })
);
NAND #() 
NAND_363_ (
  .A({ S822 }),
  .B({ S823 }),
  .Y({ S824 })
);
NAND #() 
NAND_364_ (
  .A({ S435 }),
  .B({ S824 }),
  .Y({ S825 })
);
NOR #() 
NOR_147_ (
  .A({ datapath_theregisterfile_memtrf_135 }),
  .B({ S422 }),
  .Y({ S826 })
);
NAND #() 
NAND_365_ (
  .A({ S7728 }),
  .B({ S422 }),
  .Y({ S827 })
);
NAND #() 
NAND_366_ (
  .A({ S436 }),
  .B({ S827 }),
  .Y({ S828 })
);
NOR #() 
NOR_148_ (
  .A({ S826 }),
  .B({ S828 }),
  .Y({ S829 })
);
NOR #() 
NOR_149_ (
  .A({ S442 }),
  .B({ S821 }),
  .Y({ S830 })
);
NOR #() 
NOR_150_ (
  .A({ S441 }),
  .B({ S829 }),
  .Y({ S831 })
);
NAND #() 
NAND_367_ (
  .A({ S825 }),
  .B({ S831 }),
  .Y({ S832 })
);
NAND #() 
NAND_368_ (
  .A({ S428 }),
  .B({ S832 }),
  .Y({ S833 })
);
NOR #() 
NOR_151_ (
  .A({ S830 }),
  .B({ S833 }),
  .Y({ S834 })
);
NAND #() 
NAND_369_ (
  .A({ datapath_theregisterfile_memtrf_55 }),
  .B({ S435 }),
  .Y({ S835 })
);
NAND #() 
NAND_370_ (
  .A({ datapath_theregisterfile_memtrf_39 }),
  .B({ S436 }),
  .Y({ S836 })
);
NAND #() 
NAND_371_ (
  .A({ S835 }),
  .B({ S836 }),
  .Y({ S837 })
);
NAND #() 
NAND_372_ (
  .A({ S441 }),
  .B({ S837 }),
  .Y({ S838 })
);
NAND #() 
NAND_373_ (
  .A({ datapath_theregisterfile_memtrf_7 }),
  .B({ S436 }),
  .Y({ S839 })
);
NAND #() 
NAND_374_ (
  .A({ datapath_theregisterfile_memtrf_23 }),
  .B({ S435 }),
  .Y({ S840 })
);
NAND #() 
NAND_375_ (
  .A({ S839 }),
  .B({ S840 }),
  .Y({ S841 })
);
NAND #() 
NAND_376_ (
  .A({ S442 }),
  .B({ S841 }),
  .Y({ S842 })
);
NAND #() 
NAND_377_ (
  .A({ S838 }),
  .B({ S842 }),
  .Y({ S843 })
);
NAND #() 
NAND_378_ (
  .A({ S429 }),
  .B({ S843 }),
  .Y({ S844 })
);
NAND #() 
NAND_379_ (
  .A({ datapath_theregisterfile_memtrf_119 }),
  .B({ S435 }),
  .Y({ S845 })
);
NAND #() 
NAND_380_ (
  .A({ datapath_theregisterfile_memtrf_103 }),
  .B({ S436 }),
  .Y({ S846 })
);
NAND #() 
NAND_381_ (
  .A({ S845 }),
  .B({ S846 }),
  .Y({ S847 })
);
NAND #() 
NAND_382_ (
  .A({ S441 }),
  .B({ S847 }),
  .Y({ S848 })
);
NAND #() 
NAND_383_ (
  .A({ datapath_theregisterfile_memtrf_87 }),
  .B({ S435 }),
  .Y({ S849 })
);
NAND #() 
NAND_384_ (
  .A({ datapath_theregisterfile_memtrf_71 }),
  .B({ S436 }),
  .Y({ S850 })
);
NAND #() 
NAND_385_ (
  .A({ S849 }),
  .B({ S850 }),
  .Y({ S851 })
);
NAND #() 
NAND_386_ (
  .A({ S442 }),
  .B({ S851 }),
  .Y({ S852 })
);
NAND #() 
NAND_387_ (
  .A({ S848 }),
  .B({ S852 }),
  .Y({ S853 })
);
NAND #() 
NAND_388_ (
  .A({ S479 }),
  .B({ S853 }),
  .Y({ S854 })
);
NAND #() 
NAND_389_ (
  .A({ S844 }),
  .B({ S854 }),
  .Y({ S855 })
);
NOR #() 
NOR_152_ (
  .A({ S834 }),
  .B({ S855 }),
  .Y({ S856 })
);
NAND #() 
NAND_390_ (
  .A({ S446 }),
  .B({ S856 }),
  .Y({ S857 })
);
NAND #() 
NAND_391_ (
  .A({ S812 }),
  .B({ S857 }),
  .Y({ S858 })
);
NOT #() 
NOT_137_ (
  .A({ S858 }),
  .Y({ datapath_addsubunit_in1_7 })
);
NAND #() 
NAND_392_ (
  .A({ S496 }),
  .B({ datapath_addsubunit_in1_7 }),
  .Y({ S859 })
);
NAND #() 
NAND_393_ (
  .A({ S372 }),
  .B({ S859 }),
  .Y({ S860 })
);
NOT #() 
NOT_138_ (
  .A({ S860 }),
  .Y({ S861 })
);
NOR #() 
NOR_153_ (
  .A({ S7936 }),
  .B({ S861 }),
  .Y({ S862 })
);
NOR #() 
NOR_154_ (
  .A({ datapath_muxmem_in2_7 }),
  .B({ S860 }),
  .Y({ S863 })
);
NAND #() 
NAND_394_ (
  .A({ S7876 }),
  .B({ S445 }),
  .Y({ S864 })
);
NAND #() 
NAND_395_ (
  .A({ datapath_theregisterfile_memtrf_182 }),
  .B({ S423 }),
  .Y({ S865 })
);
NAND #() 
NAND_396_ (
  .A({ datapath_theregisterfile_memtrf_246 }),
  .B({ S422 }),
  .Y({ S866 })
);
NAND #() 
NAND_397_ (
  .A({ S865 }),
  .B({ S866 }),
  .Y({ S867 })
);
NAND #() 
NAND_398_ (
  .A({ S435 }),
  .B({ S867 }),
  .Y({ S868 })
);
NOR #() 
NOR_155_ (
  .A({ datapath_theregisterfile_memtrf_166 }),
  .B({ S422 }),
  .Y({ S869 })
);
NOR #() 
NOR_156_ (
  .A({ datapath_theregisterfile_memtrf_230 }),
  .B({ S423 }),
  .Y({ S870 })
);
NOR #() 
NOR_157_ (
  .A({ S869 }),
  .B({ S870 }),
  .Y({ S871 })
);
NAND #() 
NAND_399_ (
  .A({ S436 }),
  .B({ S871 }),
  .Y({ S872 })
);
NAND #() 
NAND_400_ (
  .A({ S868 }),
  .B({ S872 }),
  .Y({ S873 })
);
NAND #() 
NAND_401_ (
  .A({ datapath_theregisterfile_memtrf_214 }),
  .B({ S422 }),
  .Y({ S874 })
);
NAND #() 
NAND_402_ (
  .A({ datapath_theregisterfile_memtrf_150 }),
  .B({ S423 }),
  .Y({ S875 })
);
NAND #() 
NAND_403_ (
  .A({ S874 }),
  .B({ S875 }),
  .Y({ S876 })
);
NAND #() 
NAND_404_ (
  .A({ S435 }),
  .B({ S876 }),
  .Y({ S877 })
);
NOR #() 
NOR_158_ (
  .A({ datapath_theregisterfile_memtrf_134 }),
  .B({ S422 }),
  .Y({ S878 })
);
NAND #() 
NAND_405_ (
  .A({ S7717 }),
  .B({ S422 }),
  .Y({ S879 })
);
NAND #() 
NAND_406_ (
  .A({ S436 }),
  .B({ S879 }),
  .Y({ S880 })
);
NOR #() 
NOR_159_ (
  .A({ S878 }),
  .B({ S880 }),
  .Y({ S881 })
);
NOR #() 
NOR_160_ (
  .A({ S442 }),
  .B({ S873 }),
  .Y({ S882 })
);
NOR #() 
NOR_161_ (
  .A({ S441 }),
  .B({ S881 }),
  .Y({ S883 })
);
NAND #() 
NAND_407_ (
  .A({ S877 }),
  .B({ S883 }),
  .Y({ S884 })
);
NAND #() 
NAND_408_ (
  .A({ S428 }),
  .B({ S884 }),
  .Y({ S885 })
);
NOR #() 
NOR_162_ (
  .A({ S882 }),
  .B({ S885 }),
  .Y({ S886 })
);
NAND #() 
NAND_409_ (
  .A({ datapath_theregisterfile_memtrf_54 }),
  .B({ S435 }),
  .Y({ S887 })
);
NAND #() 
NAND_410_ (
  .A({ datapath_theregisterfile_memtrf_38 }),
  .B({ S436 }),
  .Y({ S888 })
);
NAND #() 
NAND_411_ (
  .A({ S887 }),
  .B({ S888 }),
  .Y({ S889 })
);
NAND #() 
NAND_412_ (
  .A({ S441 }),
  .B({ S889 }),
  .Y({ S890 })
);
NAND #() 
NAND_413_ (
  .A({ datapath_theregisterfile_memtrf_6 }),
  .B({ S436 }),
  .Y({ S891 })
);
NAND #() 
NAND_414_ (
  .A({ datapath_theregisterfile_memtrf_22 }),
  .B({ S435 }),
  .Y({ S892 })
);
NAND #() 
NAND_415_ (
  .A({ S891 }),
  .B({ S892 }),
  .Y({ S893 })
);
NAND #() 
NAND_416_ (
  .A({ S442 }),
  .B({ S893 }),
  .Y({ S894 })
);
NAND #() 
NAND_417_ (
  .A({ S890 }),
  .B({ S894 }),
  .Y({ S895 })
);
NAND #() 
NAND_418_ (
  .A({ S429 }),
  .B({ S895 }),
  .Y({ S896 })
);
NAND #() 
NAND_419_ (
  .A({ datapath_theregisterfile_memtrf_118 }),
  .B({ S435 }),
  .Y({ S897 })
);
NAND #() 
NAND_420_ (
  .A({ datapath_theregisterfile_memtrf_102 }),
  .B({ S436 }),
  .Y({ S898 })
);
NAND #() 
NAND_421_ (
  .A({ S897 }),
  .B({ S898 }),
  .Y({ S899 })
);
NAND #() 
NAND_422_ (
  .A({ S441 }),
  .B({ S899 }),
  .Y({ S900 })
);
NAND #() 
NAND_423_ (
  .A({ datapath_theregisterfile_memtrf_86 }),
  .B({ S435 }),
  .Y({ S901 })
);
NAND #() 
NAND_424_ (
  .A({ datapath_theregisterfile_memtrf_70 }),
  .B({ S436 }),
  .Y({ S902 })
);
NAND #() 
NAND_425_ (
  .A({ S901 }),
  .B({ S902 }),
  .Y({ S903 })
);
NAND #() 
NAND_426_ (
  .A({ S442 }),
  .B({ S903 }),
  .Y({ S904 })
);
NAND #() 
NAND_427_ (
  .A({ S900 }),
  .B({ S904 }),
  .Y({ S905 })
);
NAND #() 
NAND_428_ (
  .A({ S479 }),
  .B({ S905 }),
  .Y({ S906 })
);
NAND #() 
NAND_429_ (
  .A({ S446 }),
  .B({ S906 }),
  .Y({ S907 })
);
NOR #() 
NOR_163_ (
  .A({ S886 }),
  .B({ S907 }),
  .Y({ S908 })
);
NAND #() 
NAND_430_ (
  .A({ S896 }),
  .B({ S908 }),
  .Y({ S909 })
);
NAND #() 
NAND_431_ (
  .A({ S864 }),
  .B({ S909 }),
  .Y({ S910 })
);
NOT #() 
NOT_139_ (
  .A({ S910 }),
  .Y({ datapath_addsubunit_in1_6 })
);
NAND #() 
NAND_432_ (
  .A({ S496 }),
  .B({ datapath_addsubunit_in1_6 }),
  .Y({ S911 })
);
NAND #() 
NAND_433_ (
  .A({ S372 }),
  .B({ S911 }),
  .Y({ S912 })
);
NAND #() 
NAND_434_ (
  .A({ datapath_muxmem_in2_6 }),
  .B({ S912 }),
  .Y({ S913 })
);
NOT #() 
NOT_140_ (
  .A({ S913 }),
  .Y({ S914 })
);
NOR #() 
NOR_164_ (
  .A({ datapath_muxmem_in2_6 }),
  .B({ S912 }),
  .Y({ S915 })
);
NOR #() 
NOR_165_ (
  .A({ S914 }),
  .B({ S915 }),
  .Y({ S916 })
);
NAND #() 
NAND_435_ (
  .A({ S7869 }),
  .B({ S445 }),
  .Y({ S917 })
);
NAND #() 
NAND_436_ (
  .A({ datapath_theregisterfile_memtrf_181 }),
  .B({ S423 }),
  .Y({ S918 })
);
NAND #() 
NAND_437_ (
  .A({ datapath_theregisterfile_memtrf_245 }),
  .B({ S422 }),
  .Y({ S919 })
);
NAND #() 
NAND_438_ (
  .A({ S918 }),
  .B({ S919 }),
  .Y({ S920 })
);
NAND #() 
NAND_439_ (
  .A({ S435 }),
  .B({ S920 }),
  .Y({ S921 })
);
NOR #() 
NOR_166_ (
  .A({ datapath_theregisterfile_memtrf_165 }),
  .B({ S422 }),
  .Y({ S922 })
);
NOR #() 
NOR_167_ (
  .A({ datapath_theregisterfile_memtrf_229 }),
  .B({ S423 }),
  .Y({ S923 })
);
NOR #() 
NOR_168_ (
  .A({ S922 }),
  .B({ S923 }),
  .Y({ S924 })
);
NAND #() 
NAND_440_ (
  .A({ S436 }),
  .B({ S924 }),
  .Y({ S925 })
);
NAND #() 
NAND_441_ (
  .A({ S921 }),
  .B({ S925 }),
  .Y({ S926 })
);
NAND #() 
NAND_442_ (
  .A({ datapath_theregisterfile_memtrf_213 }),
  .B({ S422 }),
  .Y({ S927 })
);
NAND #() 
NAND_443_ (
  .A({ datapath_theregisterfile_memtrf_149 }),
  .B({ S423 }),
  .Y({ S928 })
);
NAND #() 
NAND_444_ (
  .A({ S927 }),
  .B({ S928 }),
  .Y({ S929 })
);
NAND #() 
NAND_445_ (
  .A({ S435 }),
  .B({ S929 }),
  .Y({ S930 })
);
NOR #() 
NOR_169_ (
  .A({ datapath_theregisterfile_memtrf_133 }),
  .B({ S422 }),
  .Y({ S931 })
);
NAND #() 
NAND_446_ (
  .A({ S7706 }),
  .B({ S422 }),
  .Y({ S932 })
);
NAND #() 
NAND_447_ (
  .A({ S436 }),
  .B({ S932 }),
  .Y({ S933 })
);
NOR #() 
NOR_170_ (
  .A({ S931 }),
  .B({ S933 }),
  .Y({ S934 })
);
NOR #() 
NOR_171_ (
  .A({ S442 }),
  .B({ S926 }),
  .Y({ S935 })
);
NOR #() 
NOR_172_ (
  .A({ S441 }),
  .B({ S934 }),
  .Y({ S936 })
);
NAND #() 
NAND_448_ (
  .A({ S930 }),
  .B({ S936 }),
  .Y({ S937 })
);
NAND #() 
NAND_449_ (
  .A({ S428 }),
  .B({ S937 }),
  .Y({ S938 })
);
NOR #() 
NOR_173_ (
  .A({ S935 }),
  .B({ S938 }),
  .Y({ S939 })
);
NAND #() 
NAND_450_ (
  .A({ datapath_theregisterfile_memtrf_53 }),
  .B({ S435 }),
  .Y({ S940 })
);
NAND #() 
NAND_451_ (
  .A({ datapath_theregisterfile_memtrf_37 }),
  .B({ S436 }),
  .Y({ S941 })
);
NAND #() 
NAND_452_ (
  .A({ S940 }),
  .B({ S941 }),
  .Y({ S942 })
);
NAND #() 
NAND_453_ (
  .A({ S441 }),
  .B({ S942 }),
  .Y({ S943 })
);
NAND #() 
NAND_454_ (
  .A({ datapath_theregisterfile_memtrf_5 }),
  .B({ S436 }),
  .Y({ S944 })
);
NAND #() 
NAND_455_ (
  .A({ datapath_theregisterfile_memtrf_21 }),
  .B({ S435 }),
  .Y({ S945 })
);
NAND #() 
NAND_456_ (
  .A({ S944 }),
  .B({ S945 }),
  .Y({ S946 })
);
NAND #() 
NAND_457_ (
  .A({ S442 }),
  .B({ S946 }),
  .Y({ S947 })
);
NAND #() 
NAND_458_ (
  .A({ S943 }),
  .B({ S947 }),
  .Y({ S948 })
);
NAND #() 
NAND_459_ (
  .A({ S429 }),
  .B({ S948 }),
  .Y({ S949 })
);
NAND #() 
NAND_460_ (
  .A({ datapath_theregisterfile_memtrf_117 }),
  .B({ S435 }),
  .Y({ S950 })
);
NAND #() 
NAND_461_ (
  .A({ datapath_theregisterfile_memtrf_101 }),
  .B({ S436 }),
  .Y({ S951 })
);
NAND #() 
NAND_462_ (
  .A({ S950 }),
  .B({ S951 }),
  .Y({ S952 })
);
NAND #() 
NAND_463_ (
  .A({ S441 }),
  .B({ S952 }),
  .Y({ S953 })
);
NAND #() 
NAND_464_ (
  .A({ datapath_theregisterfile_memtrf_85 }),
  .B({ S435 }),
  .Y({ S954 })
);
NAND #() 
NAND_465_ (
  .A({ datapath_theregisterfile_memtrf_69 }),
  .B({ S436 }),
  .Y({ S955 })
);
NAND #() 
NAND_466_ (
  .A({ S954 }),
  .B({ S955 }),
  .Y({ S956 })
);
NAND #() 
NAND_467_ (
  .A({ S442 }),
  .B({ S956 }),
  .Y({ S957 })
);
NAND #() 
NAND_468_ (
  .A({ S953 }),
  .B({ S957 }),
  .Y({ S958 })
);
NAND #() 
NAND_469_ (
  .A({ S479 }),
  .B({ S958 }),
  .Y({ S959 })
);
NAND #() 
NAND_470_ (
  .A({ S949 }),
  .B({ S959 }),
  .Y({ S960 })
);
NOR #() 
NOR_174_ (
  .A({ S939 }),
  .B({ S960 }),
  .Y({ S961 })
);
NAND #() 
NAND_471_ (
  .A({ S446 }),
  .B({ S961 }),
  .Y({ S962 })
);
NAND #() 
NAND_472_ (
  .A({ S917 }),
  .B({ S962 }),
  .Y({ S963 })
);
NOT #() 
NOT_141_ (
  .A({ S963 }),
  .Y({ datapath_addsubunit_in1_5 })
);
NAND #() 
NAND_473_ (
  .A({ S496 }),
  .B({ datapath_addsubunit_in1_5 }),
  .Y({ S964 })
);
NAND #() 
NAND_474_ (
  .A({ S372 }),
  .B({ S964 }),
  .Y({ S965 })
);
NOT #() 
NOT_142_ (
  .A({ S965 }),
  .Y({ S966 })
);
NOR #() 
NOR_175_ (
  .A({ S7920 }),
  .B({ S966 }),
  .Y({ S967 })
);
NOR #() 
NOR_176_ (
  .A({ datapath_muxmem_in2_5 }),
  .B({ S965 }),
  .Y({ S968 })
);
NAND #() 
NAND_475_ (
  .A({ controller_fib_4 }),
  .B({ S370 }),
  .Y({ S969 })
);
NAND #() 
NAND_476_ (
  .A({ S7861 }),
  .B({ S445 }),
  .Y({ S970 })
);
NOR #() 
NOR_177_ (
  .A({ datapath_theregisterfile_memtrf_164 }),
  .B({ S422 }),
  .Y({ S971 })
);
NOR #() 
NOR_178_ (
  .A({ datapath_theregisterfile_memtrf_228 }),
  .B({ S423 }),
  .Y({ S972 })
);
NOR #() 
NOR_179_ (
  .A({ S971 }),
  .B({ S972 }),
  .Y({ S973 })
);
NAND #() 
NAND_477_ (
  .A({ S436 }),
  .B({ S973 }),
  .Y({ S974 })
);
NOR #() 
NOR_180_ (
  .A({ datapath_theregisterfile_memtrf_244 }),
  .B({ S423 }),
  .Y({ S975 })
);
NAND #() 
NAND_478_ (
  .A({ S7596 }),
  .B({ S423 }),
  .Y({ S976 })
);
NAND #() 
NAND_479_ (
  .A({ S435 }),
  .B({ S976 }),
  .Y({ S977 })
);
NOR #() 
NOR_181_ (
  .A({ S975 }),
  .B({ S977 }),
  .Y({ S978 })
);
NAND #() 
NAND_480_ (
  .A({ datapath_theregisterfile_memtrf_196 }),
  .B({ S436 }),
  .Y({ S979 })
);
NAND #() 
NAND_481_ (
  .A({ datapath_theregisterfile_memtrf_212 }),
  .B({ S435 }),
  .Y({ S980 })
);
NAND #() 
NAND_482_ (
  .A({ S979 }),
  .B({ S980 }),
  .Y({ S981 })
);
NAND #() 
NAND_483_ (
  .A({ S422 }),
  .B({ S981 }),
  .Y({ S982 })
);
NAND #() 
NAND_484_ (
  .A({ datapath_theregisterfile_memtrf_132 }),
  .B({ S436 }),
  .Y({ S983 })
);
NAND #() 
NAND_485_ (
  .A({ datapath_theregisterfile_memtrf_148 }),
  .B({ S435 }),
  .Y({ S984 })
);
NAND #() 
NAND_486_ (
  .A({ S983 }),
  .B({ S984 }),
  .Y({ S985 })
);
NAND #() 
NAND_487_ (
  .A({ S423 }),
  .B({ S985 }),
  .Y({ S986 })
);
NAND #() 
NAND_488_ (
  .A({ S982 }),
  .B({ S986 }),
  .Y({ S987 })
);
NOR #() 
NOR_182_ (
  .A({ S441 }),
  .B({ S987 }),
  .Y({ S988 })
);
NOR #() 
NOR_183_ (
  .A({ S442 }),
  .B({ S978 }),
  .Y({ S989 })
);
NAND #() 
NAND_489_ (
  .A({ S974 }),
  .B({ S989 }),
  .Y({ S990 })
);
NAND #() 
NAND_490_ (
  .A({ S428 }),
  .B({ S990 }),
  .Y({ S991 })
);
NOR #() 
NOR_184_ (
  .A({ S988 }),
  .B({ S991 }),
  .Y({ S992 })
);
NAND #() 
NAND_491_ (
  .A({ datapath_theregisterfile_memtrf_116 }),
  .B({ S435 }),
  .Y({ S993 })
);
NAND #() 
NAND_492_ (
  .A({ datapath_theregisterfile_memtrf_100 }),
  .B({ S436 }),
  .Y({ S994 })
);
NAND #() 
NAND_493_ (
  .A({ S993 }),
  .B({ S994 }),
  .Y({ S995 })
);
NAND #() 
NAND_494_ (
  .A({ S441 }),
  .B({ S995 }),
  .Y({ S996 })
);
NAND #() 
NAND_495_ (
  .A({ datapath_theregisterfile_memtrf_84 }),
  .B({ S435 }),
  .Y({ S997 })
);
NAND #() 
NAND_496_ (
  .A({ datapath_theregisterfile_memtrf_68 }),
  .B({ S436 }),
  .Y({ S998 })
);
NAND #() 
NAND_497_ (
  .A({ S997 }),
  .B({ S998 }),
  .Y({ S999 })
);
NAND #() 
NAND_498_ (
  .A({ S442 }),
  .B({ S999 }),
  .Y({ S1000 })
);
NAND #() 
NAND_499_ (
  .A({ S996 }),
  .B({ S1000 }),
  .Y({ S1001 })
);
NAND #() 
NAND_500_ (
  .A({ S479 }),
  .B({ S1001 }),
  .Y({ S1002 })
);
NOR #() 
NOR_185_ (
  .A({ S436 }),
  .B({ S442 }),
  .Y({ S1003 })
);
NAND #() 
NAND_501_ (
  .A({ datapath_theregisterfile_memtrf_52 }),
  .B({ S1003 }),
  .Y({ S1004 })
);
NOR #() 
NOR_186_ (
  .A({ datapath_theregisterfile_memtrf_20 }),
  .B({ S436 }),
  .Y({ S1005 })
);
NOR #() 
NOR_187_ (
  .A({ S441 }),
  .B({ S1005 }),
  .Y({ S1006 })
);
NAND #() 
NAND_502_ (
  .A({ datapath_theregisterfile_memtrf_36 }),
  .B({ S436 }),
  .Y({ S1007 })
);
NAND #() 
NAND_503_ (
  .A({ S1004 }),
  .B({ S1007 }),
  .Y({ S1008 })
);
NOR #() 
NOR_188_ (
  .A({ S1006 }),
  .B({ S1008 }),
  .Y({ S1009 })
);
NOR #() 
NOR_189_ (
  .A({ S430 }),
  .B({ S1009 }),
  .Y({ S1010 })
);
NOR #() 
NOR_190_ (
  .A({ S992 }),
  .B({ S1010 }),
  .Y({ S1011 })
);
NAND #() 
NAND_504_ (
  .A({ S1002 }),
  .B({ S1011 }),
  .Y({ S1012 })
);
NAND #() 
NAND_505_ (
  .A({ S970 }),
  .B({ S1012 }),
  .Y({ S1013 })
);
NOT #() 
NOT_143_ (
  .A({ S1013 }),
  .Y({ datapath_addsubunit_in1_4 })
);
NAND #() 
NAND_506_ (
  .A({ S496 }),
  .B({ datapath_addsubunit_in1_4 }),
  .Y({ S1014 })
);
NAND #() 
NAND_507_ (
  .A({ S969 }),
  .B({ S1014 }),
  .Y({ S1015 })
);
NAND #() 
NAND_508_ (
  .A({ datapath_muxmem_in2_4 }),
  .B({ S1015 }),
  .Y({ S1016 })
);
NOT #() 
NOT_144_ (
  .A({ S1016 }),
  .Y({ S1017 })
);
NOR #() 
NOR_191_ (
  .A({ datapath_muxmem_in2_4 }),
  .B({ S1015 }),
  .Y({ S1018 })
);
NOR #() 
NOR_192_ (
  .A({ S1017 }),
  .B({ S1018 }),
  .Y({ S1019 })
);
NAND #() 
NAND_509_ (
  .A({ controller_fib_3 }),
  .B({ S370 }),
  .Y({ S1020 })
);
NAND #() 
NAND_510_ (
  .A({ S7853 }),
  .B({ S445 }),
  .Y({ S1021 })
);
NOR #() 
NOR_193_ (
  .A({ datapath_theregisterfile_memtrf_163 }),
  .B({ S422 }),
  .Y({ S1022 })
);
NOR #() 
NOR_194_ (
  .A({ datapath_theregisterfile_memtrf_227 }),
  .B({ S423 }),
  .Y({ S1023 })
);
NOR #() 
NOR_195_ (
  .A({ S1022 }),
  .B({ S1023 }),
  .Y({ S1024 })
);
NAND #() 
NAND_511_ (
  .A({ S436 }),
  .B({ S1024 }),
  .Y({ S1025 })
);
NOR #() 
NOR_196_ (
  .A({ datapath_theregisterfile_memtrf_243 }),
  .B({ S423 }),
  .Y({ S1026 })
);
NAND #() 
NAND_512_ (
  .A({ S7585 }),
  .B({ S423 }),
  .Y({ S1027 })
);
NAND #() 
NAND_513_ (
  .A({ S435 }),
  .B({ S1027 }),
  .Y({ S1028 })
);
NOR #() 
NOR_197_ (
  .A({ S1026 }),
  .B({ S1028 }),
  .Y({ S1029 })
);
NAND #() 
NAND_514_ (
  .A({ datapath_theregisterfile_memtrf_195 }),
  .B({ S436 }),
  .Y({ S1030 })
);
NAND #() 
NAND_515_ (
  .A({ datapath_theregisterfile_memtrf_211 }),
  .B({ S435 }),
  .Y({ S1031 })
);
NAND #() 
NAND_516_ (
  .A({ S1030 }),
  .B({ S1031 }),
  .Y({ S1032 })
);
NAND #() 
NAND_517_ (
  .A({ S422 }),
  .B({ S1032 }),
  .Y({ S1033 })
);
NAND #() 
NAND_518_ (
  .A({ datapath_theregisterfile_memtrf_131 }),
  .B({ S436 }),
  .Y({ S1034 })
);
NAND #() 
NAND_519_ (
  .A({ datapath_theregisterfile_memtrf_147 }),
  .B({ S435 }),
  .Y({ S1035 })
);
NAND #() 
NAND_520_ (
  .A({ S1034 }),
  .B({ S1035 }),
  .Y({ S1036 })
);
NAND #() 
NAND_521_ (
  .A({ S423 }),
  .B({ S1036 }),
  .Y({ S1037 })
);
NAND #() 
NAND_522_ (
  .A({ S1033 }),
  .B({ S1037 }),
  .Y({ S1038 })
);
NOR #() 
NOR_198_ (
  .A({ S441 }),
  .B({ S1038 }),
  .Y({ S1039 })
);
NOR #() 
NOR_199_ (
  .A({ S442 }),
  .B({ S1029 }),
  .Y({ S1040 })
);
NAND #() 
NAND_523_ (
  .A({ S1025 }),
  .B({ S1040 }),
  .Y({ S1041 })
);
NAND #() 
NAND_524_ (
  .A({ S428 }),
  .B({ S1041 }),
  .Y({ S1042 })
);
NOR #() 
NOR_200_ (
  .A({ S1039 }),
  .B({ S1042 }),
  .Y({ S1043 })
);
NAND #() 
NAND_525_ (
  .A({ datapath_theregisterfile_memtrf_83 }),
  .B({ S442 }),
  .Y({ S1044 })
);
NAND #() 
NAND_526_ (
  .A({ datapath_theregisterfile_memtrf_115 }),
  .B({ S441 }),
  .Y({ S1045 })
);
NAND #() 
NAND_527_ (
  .A({ S1044 }),
  .B({ S1045 }),
  .Y({ S1046 })
);
NAND #() 
NAND_528_ (
  .A({ S435 }),
  .B({ S1046 }),
  .Y({ S1047 })
);
NAND #() 
NAND_529_ (
  .A({ datapath_theregisterfile_memtrf_99 }),
  .B({ S441 }),
  .Y({ S1048 })
);
NAND #() 
NAND_530_ (
  .A({ datapath_theregisterfile_memtrf_67 }),
  .B({ S442 }),
  .Y({ S1049 })
);
NAND #() 
NAND_531_ (
  .A({ S1048 }),
  .B({ S1049 }),
  .Y({ S1050 })
);
NAND #() 
NAND_532_ (
  .A({ S436 }),
  .B({ S1050 }),
  .Y({ S1051 })
);
NAND #() 
NAND_533_ (
  .A({ S1047 }),
  .B({ S1051 }),
  .Y({ S1052 })
);
NAND #() 
NAND_534_ (
  .A({ S479 }),
  .B({ S1052 }),
  .Y({ S1053 })
);
NAND #() 
NAND_535_ (
  .A({ datapath_theregisterfile_memtrf_51 }),
  .B({ S1003 }),
  .Y({ S1054 })
);
NAND #() 
NAND_536_ (
  .A({ datapath_theregisterfile_memtrf_35 }),
  .B({ S436 }),
  .Y({ S1055 })
);
NOT #() 
NOT_145_ (
  .A({ S1055 }),
  .Y({ S1056 })
);
NOR #() 
NOR_201_ (
  .A({ datapath_theregisterfile_memtrf_19 }),
  .B({ S436 }),
  .Y({ S1057 })
);
NOR #() 
NOR_202_ (
  .A({ S441 }),
  .B({ S1057 }),
  .Y({ S1058 })
);
NOR #() 
NOR_203_ (
  .A({ S1056 }),
  .B({ S1058 }),
  .Y({ S1059 })
);
NAND #() 
NAND_537_ (
  .A({ S1054 }),
  .B({ S1059 }),
  .Y({ S1060 })
);
NAND #() 
NAND_538_ (
  .A({ S429 }),
  .B({ S1060 }),
  .Y({ S1061 })
);
NOT #() 
NOT_146_ (
  .A({ S1061 }),
  .Y({ S1062 })
);
NOR #() 
NOR_204_ (
  .A({ S1043 }),
  .B({ S1062 }),
  .Y({ S1063 })
);
NAND #() 
NAND_539_ (
  .A({ S1053 }),
  .B({ S1063 }),
  .Y({ S1064 })
);
NAND #() 
NAND_540_ (
  .A({ S1021 }),
  .B({ S1064 }),
  .Y({ S1065 })
);
NOT #() 
NOT_147_ (
  .A({ S1065 }),
  .Y({ datapath_addsubunit_in1_3 })
);
NAND #() 
NAND_541_ (
  .A({ S496 }),
  .B({ datapath_addsubunit_in1_3 }),
  .Y({ S1066 })
);
NAND #() 
NAND_542_ (
  .A({ S1020 }),
  .B({ S1066 }),
  .Y({ S1067 })
);
NAND #() 
NAND_543_ (
  .A({ datapath_muxmem_in2_3 }),
  .B({ S1067 }),
  .Y({ S1068 })
);
NOT #() 
NOT_148_ (
  .A({ S1068 }),
  .Y({ S1069 })
);
NOR #() 
NOR_205_ (
  .A({ datapath_muxmem_in2_3 }),
  .B({ S1067 }),
  .Y({ S1070 })
);
NAND #() 
NAND_544_ (
  .A({ controller_fib_2 }),
  .B({ S370 }),
  .Y({ S1071 })
);
NAND #() 
NAND_545_ (
  .A({ S7846 }),
  .B({ S445 }),
  .Y({ S1072 })
);
NAND #() 
NAND_546_ (
  .A({ datapath_theregisterfile_memtrf_178 }),
  .B({ S423 }),
  .Y({ S1073 })
);
NAND #() 
NAND_547_ (
  .A({ datapath_theregisterfile_memtrf_242 }),
  .B({ S422 }),
  .Y({ S1074 })
);
NAND #() 
NAND_548_ (
  .A({ S1073 }),
  .B({ S1074 }),
  .Y({ S1075 })
);
NAND #() 
NAND_549_ (
  .A({ S435 }),
  .B({ S1075 }),
  .Y({ S1076 })
);
NOR #() 
NOR_206_ (
  .A({ datapath_theregisterfile_memtrf_162 }),
  .B({ S422 }),
  .Y({ S1077 })
);
NOR #() 
NOR_207_ (
  .A({ datapath_theregisterfile_memtrf_226 }),
  .B({ S423 }),
  .Y({ S1078 })
);
NOR #() 
NOR_208_ (
  .A({ S1077 }),
  .B({ S1078 }),
  .Y({ S1079 })
);
NAND #() 
NAND_550_ (
  .A({ S436 }),
  .B({ S1079 }),
  .Y({ S1080 })
);
NAND #() 
NAND_551_ (
  .A({ S1076 }),
  .B({ S1080 }),
  .Y({ S1081 })
);
NAND #() 
NAND_552_ (
  .A({ S441 }),
  .B({ S1081 }),
  .Y({ S1082 })
);
NAND #() 
NAND_553_ (
  .A({ datapath_theregisterfile_memtrf_210 }),
  .B({ S422 }),
  .Y({ S1083 })
);
NAND #() 
NAND_554_ (
  .A({ datapath_theregisterfile_memtrf_146 }),
  .B({ S423 }),
  .Y({ S1084 })
);
NAND #() 
NAND_555_ (
  .A({ S1083 }),
  .B({ S1084 }),
  .Y({ S1085 })
);
NAND #() 
NAND_556_ (
  .A({ S435 }),
  .B({ S1085 }),
  .Y({ S1086 })
);
NOR #() 
NOR_209_ (
  .A({ datapath_theregisterfile_memtrf_130 }),
  .B({ S422 }),
  .Y({ S1087 })
);
NOR #() 
NOR_210_ (
  .A({ datapath_theregisterfile_memtrf_194 }),
  .B({ S423 }),
  .Y({ S1088 })
);
NOR #() 
NOR_211_ (
  .A({ S1087 }),
  .B({ S1088 }),
  .Y({ S1089 })
);
NAND #() 
NAND_557_ (
  .A({ S436 }),
  .B({ S1089 }),
  .Y({ S1090 })
);
NAND #() 
NAND_558_ (
  .A({ S1086 }),
  .B({ S1090 }),
  .Y({ S1091 })
);
NAND #() 
NAND_559_ (
  .A({ S442 }),
  .B({ S1091 }),
  .Y({ S1092 })
);
NAND #() 
NAND_560_ (
  .A({ S1082 }),
  .B({ S1092 }),
  .Y({ S1093 })
);
NAND #() 
NAND_561_ (
  .A({ S428 }),
  .B({ S1093 }),
  .Y({ S1094 })
);
NAND #() 
NAND_562_ (
  .A({ datapath_theregisterfile_memtrf_114 }),
  .B({ S435 }),
  .Y({ S1095 })
);
NAND #() 
NAND_563_ (
  .A({ datapath_theregisterfile_memtrf_98 }),
  .B({ S436 }),
  .Y({ S1096 })
);
NAND #() 
NAND_564_ (
  .A({ S1095 }),
  .B({ S1096 }),
  .Y({ S1097 })
);
NAND #() 
NAND_565_ (
  .A({ S441 }),
  .B({ S1097 }),
  .Y({ S1098 })
);
NAND #() 
NAND_566_ (
  .A({ datapath_theregisterfile_memtrf_82 }),
  .B({ S435 }),
  .Y({ S1099 })
);
NAND #() 
NAND_567_ (
  .A({ datapath_theregisterfile_memtrf_66 }),
  .B({ S436 }),
  .Y({ S1100 })
);
NAND #() 
NAND_568_ (
  .A({ S1099 }),
  .B({ S1100 }),
  .Y({ S1101 })
);
NAND #() 
NAND_569_ (
  .A({ S442 }),
  .B({ S1101 }),
  .Y({ S1102 })
);
NAND #() 
NAND_570_ (
  .A({ S1098 }),
  .B({ S1102 }),
  .Y({ S1103 })
);
NAND #() 
NAND_571_ (
  .A({ S479 }),
  .B({ S1103 }),
  .Y({ S1104 })
);
NOT #() 
NOT_149_ (
  .A({ S1104 }),
  .Y({ S1105 })
);
NOR #() 
NOR_212_ (
  .A({ datapath_theregisterfile_memtrf_18 }),
  .B({ S441 }),
  .Y({ S1106 })
);
NOR #() 
NOR_213_ (
  .A({ datapath_theregisterfile_memtrf_50 }),
  .B({ S442 }),
  .Y({ S1107 })
);
NOR #() 
NOR_214_ (
  .A({ S1106 }),
  .B({ S1107 }),
  .Y({ S1108 })
);
NOR #() 
NOR_215_ (
  .A({ S436 }),
  .B({ S1108 }),
  .Y({ S1109 })
);
NOR #() 
NOR_216_ (
  .A({ datapath_theregisterfile_memtrf_34 }),
  .B({ S442 }),
  .Y({ S1110 })
);
NAND #() 
NAND_572_ (
  .A({ S436 }),
  .B({ S1110 }),
  .Y({ S1111 })
);
NAND #() 
NAND_573_ (
  .A({ S429 }),
  .B({ S1111 }),
  .Y({ S1112 })
);
NOR #() 
NOR_217_ (
  .A({ S1109 }),
  .B({ S1112 }),
  .Y({ S1113 })
);
NOR #() 
NOR_218_ (
  .A({ S1105 }),
  .B({ S1113 }),
  .Y({ S1114 })
);
NAND #() 
NAND_574_ (
  .A({ S1094 }),
  .B({ S1114 }),
  .Y({ S1115 })
);
NAND #() 
NAND_575_ (
  .A({ S1072 }),
  .B({ S1115 }),
  .Y({ S1116 })
);
NOT #() 
NOT_150_ (
  .A({ S1116 }),
  .Y({ datapath_addsubunit_in1_2 })
);
NAND #() 
NAND_576_ (
  .A({ S496 }),
  .B({ datapath_addsubunit_in1_2 }),
  .Y({ S1117 })
);
NAND #() 
NAND_577_ (
  .A({ S1071 }),
  .B({ S1117 }),
  .Y({ S1118 })
);
NAND #() 
NAND_578_ (
  .A({ datapath_muxmem_in2_2 }),
  .B({ S1118 }),
  .Y({ S1119 })
);
NOT #() 
NOT_151_ (
  .A({ S1119 }),
  .Y({ S1120 })
);
NAND #() 
NAND_579_ (
  .A({ controller_fib_1 }),
  .B({ S370 }),
  .Y({ S1121 })
);
NAND #() 
NAND_580_ (
  .A({ S7838 }),
  .B({ S445 }),
  .Y({ S1122 })
);
NAND #() 
NAND_581_ (
  .A({ datapath_theregisterfile_memtrf_177 }),
  .B({ S423 }),
  .Y({ S1123 })
);
NAND #() 
NAND_582_ (
  .A({ datapath_theregisterfile_memtrf_241 }),
  .B({ S422 }),
  .Y({ S1124 })
);
NAND #() 
NAND_583_ (
  .A({ S1123 }),
  .B({ S1124 }),
  .Y({ S1125 })
);
NAND #() 
NAND_584_ (
  .A({ S435 }),
  .B({ S1125 }),
  .Y({ S1126 })
);
NOR #() 
NOR_219_ (
  .A({ datapath_theregisterfile_memtrf_161 }),
  .B({ S422 }),
  .Y({ S1127 })
);
NOR #() 
NOR_220_ (
  .A({ datapath_theregisterfile_memtrf_225 }),
  .B({ S423 }),
  .Y({ S1128 })
);
NOR #() 
NOR_221_ (
  .A({ S1127 }),
  .B({ S1128 }),
  .Y({ S1129 })
);
NAND #() 
NAND_585_ (
  .A({ S436 }),
  .B({ S1129 }),
  .Y({ S1130 })
);
NAND #() 
NAND_586_ (
  .A({ S1126 }),
  .B({ S1130 }),
  .Y({ S1131 })
);
NAND #() 
NAND_587_ (
  .A({ datapath_theregisterfile_memtrf_209 }),
  .B({ S422 }),
  .Y({ S1132 })
);
NAND #() 
NAND_588_ (
  .A({ datapath_theregisterfile_memtrf_145 }),
  .B({ S423 }),
  .Y({ S1133 })
);
NAND #() 
NAND_589_ (
  .A({ S1132 }),
  .B({ S1133 }),
  .Y({ S1134 })
);
NAND #() 
NAND_590_ (
  .A({ S435 }),
  .B({ S1134 }),
  .Y({ S1135 })
);
NOR #() 
NOR_222_ (
  .A({ datapath_theregisterfile_memtrf_129 }),
  .B({ S422 }),
  .Y({ S1136 })
);
NAND #() 
NAND_591_ (
  .A({ S7684 }),
  .B({ S422 }),
  .Y({ S1137 })
);
NAND #() 
NAND_592_ (
  .A({ S436 }),
  .B({ S1137 }),
  .Y({ S1138 })
);
NOR #() 
NOR_223_ (
  .A({ S1136 }),
  .B({ S1138 }),
  .Y({ S1139 })
);
NOR #() 
NOR_224_ (
  .A({ S442 }),
  .B({ S1131 }),
  .Y({ S1140 })
);
NOR #() 
NOR_225_ (
  .A({ S441 }),
  .B({ S1139 }),
  .Y({ S1141 })
);
NAND #() 
NAND_593_ (
  .A({ S1135 }),
  .B({ S1141 }),
  .Y({ S1142 })
);
NAND #() 
NAND_594_ (
  .A({ S428 }),
  .B({ S1142 }),
  .Y({ S1143 })
);
NOR #() 
NOR_226_ (
  .A({ S1140 }),
  .B({ S1143 }),
  .Y({ S1144 })
);
NAND #() 
NAND_595_ (
  .A({ datapath_theregisterfile_memtrf_17 }),
  .B({ S442 }),
  .Y({ S1145 })
);
NAND #() 
NAND_596_ (
  .A({ datapath_theregisterfile_memtrf_49 }),
  .B({ S441 }),
  .Y({ S1146 })
);
NAND #() 
NAND_597_ (
  .A({ S1145 }),
  .B({ S1146 }),
  .Y({ S1147 })
);
NAND #() 
NAND_598_ (
  .A({ S435 }),
  .B({ S1147 }),
  .Y({ S1148 })
);
NAND #() 
NAND_599_ (
  .A({ datapath_theregisterfile_memtrf_1 }),
  .B({ S442 }),
  .Y({ S1149 })
);
NAND #() 
NAND_600_ (
  .A({ datapath_theregisterfile_memtrf_33 }),
  .B({ S441 }),
  .Y({ S1150 })
);
NAND #() 
NAND_601_ (
  .A({ S1149 }),
  .B({ S1150 }),
  .Y({ S1151 })
);
NAND #() 
NAND_602_ (
  .A({ S436 }),
  .B({ S1151 }),
  .Y({ S1152 })
);
NAND #() 
NAND_603_ (
  .A({ S1148 }),
  .B({ S1152 }),
  .Y({ S1153 })
);
NAND #() 
NAND_604_ (
  .A({ S429 }),
  .B({ S1153 }),
  .Y({ S1154 })
);
NAND #() 
NAND_605_ (
  .A({ S7531 }),
  .B({ S436 }),
  .Y({ S1155 })
);
NOR #() 
NOR_227_ (
  .A({ datapath_theregisterfile_memtrf_113 }),
  .B({ S436 }),
  .Y({ S1156 })
);
NOR #() 
NOR_228_ (
  .A({ S442 }),
  .B({ S1156 }),
  .Y({ S1157 })
);
NAND #() 
NAND_606_ (
  .A({ S1155 }),
  .B({ S1157 }),
  .Y({ S1158 })
);
NOR #() 
NOR_229_ (
  .A({ datapath_theregisterfile_memtrf_65 }),
  .B({ S435 }),
  .Y({ S1159 })
);
NOR #() 
NOR_230_ (
  .A({ datapath_theregisterfile_memtrf_81 }),
  .B({ S436 }),
  .Y({ S1160 })
);
NOR #() 
NOR_231_ (
  .A({ S1159 }),
  .B({ S1160 }),
  .Y({ S1161 })
);
NAND #() 
NAND_607_ (
  .A({ S442 }),
  .B({ S1161 }),
  .Y({ S1162 })
);
NAND #() 
NAND_608_ (
  .A({ S1158 }),
  .B({ S1162 }),
  .Y({ S1163 })
);
NAND #() 
NAND_609_ (
  .A({ S479 }),
  .B({ S1163 }),
  .Y({ S1164 })
);
NAND #() 
NAND_610_ (
  .A({ S1154 }),
  .B({ S1164 }),
  .Y({ S1165 })
);
NOR #() 
NOR_232_ (
  .A({ S1144 }),
  .B({ S1165 }),
  .Y({ S1166 })
);
NAND #() 
NAND_611_ (
  .A({ S446 }),
  .B({ S1166 }),
  .Y({ S1167 })
);
NAND #() 
NAND_612_ (
  .A({ S1122 }),
  .B({ S1167 }),
  .Y({ S1168 })
);
NOT #() 
NOT_152_ (
  .A({ S1168 }),
  .Y({ datapath_addsubunit_in1_1 })
);
NAND #() 
NAND_613_ (
  .A({ S496 }),
  .B({ datapath_addsubunit_in1_1 }),
  .Y({ S1169 })
);
NAND #() 
NAND_614_ (
  .A({ S1121 }),
  .B({ S1169 }),
  .Y({ S1170 })
);
NAND #() 
NAND_615_ (
  .A({ datapath_muxmem_in2_1 }),
  .B({ S1170 }),
  .Y({ S1171 })
);
NOT #() 
NOT_153_ (
  .A({ S1171 }),
  .Y({ S1172 })
);
NAND #() 
NAND_616_ (
  .A({ controller_fib_0 }),
  .B({ S370 }),
  .Y({ S1173 })
);
NAND #() 
NAND_617_ (
  .A({ S7830 }),
  .B({ S445 }),
  .Y({ S1174 })
);
NAND #() 
NAND_618_ (
  .A({ datapath_theregisterfile_memtrf_176 }),
  .B({ S423 }),
  .Y({ S1175 })
);
NAND #() 
NAND_619_ (
  .A({ datapath_theregisterfile_memtrf_240 }),
  .B({ S422 }),
  .Y({ S1176 })
);
NAND #() 
NAND_620_ (
  .A({ S1175 }),
  .B({ S1176 }),
  .Y({ S1177 })
);
NAND #() 
NAND_621_ (
  .A({ S435 }),
  .B({ S1177 }),
  .Y({ S1178 })
);
NOR #() 
NOR_233_ (
  .A({ datapath_theregisterfile_memtrf_160 }),
  .B({ S422 }),
  .Y({ S1179 })
);
NOR #() 
NOR_234_ (
  .A({ datapath_theregisterfile_memtrf_224 }),
  .B({ S423 }),
  .Y({ S1180 })
);
NOR #() 
NOR_235_ (
  .A({ S1179 }),
  .B({ S1180 }),
  .Y({ S1181 })
);
NAND #() 
NAND_622_ (
  .A({ S436 }),
  .B({ S1181 }),
  .Y({ S1182 })
);
NAND #() 
NAND_623_ (
  .A({ S1178 }),
  .B({ S1182 }),
  .Y({ S1183 })
);
NAND #() 
NAND_624_ (
  .A({ datapath_theregisterfile_memtrf_208 }),
  .B({ S422 }),
  .Y({ S1184 })
);
NAND #() 
NAND_625_ (
  .A({ datapath_theregisterfile_memtrf_144 }),
  .B({ S423 }),
  .Y({ S1185 })
);
NAND #() 
NAND_626_ (
  .A({ S1184 }),
  .B({ S1185 }),
  .Y({ S1186 })
);
NAND #() 
NAND_627_ (
  .A({ S435 }),
  .B({ S1186 }),
  .Y({ S1187 })
);
NOR #() 
NOR_236_ (
  .A({ datapath_theregisterfile_memtrf_128 }),
  .B({ S422 }),
  .Y({ S1188 })
);
NAND #() 
NAND_628_ (
  .A({ S7673 }),
  .B({ S422 }),
  .Y({ S1189 })
);
NAND #() 
NAND_629_ (
  .A({ S436 }),
  .B({ S1189 }),
  .Y({ S1190 })
);
NOR #() 
NOR_237_ (
  .A({ S1188 }),
  .B({ S1190 }),
  .Y({ S1191 })
);
NOR #() 
NOR_238_ (
  .A({ S442 }),
  .B({ S1183 }),
  .Y({ S1192 })
);
NOR #() 
NOR_239_ (
  .A({ S441 }),
  .B({ S1191 }),
  .Y({ S1193 })
);
NAND #() 
NAND_630_ (
  .A({ S1187 }),
  .B({ S1193 }),
  .Y({ S1194 })
);
NAND #() 
NAND_631_ (
  .A({ S428 }),
  .B({ S1194 }),
  .Y({ S1195 })
);
NOR #() 
NOR_240_ (
  .A({ S1192 }),
  .B({ S1195 }),
  .Y({ S1196 })
);
NAND #() 
NAND_632_ (
  .A({ datapath_theregisterfile_memtrf_16 }),
  .B({ S442 }),
  .Y({ S1197 })
);
NAND #() 
NAND_633_ (
  .A({ datapath_theregisterfile_memtrf_48 }),
  .B({ S441 }),
  .Y({ S1198 })
);
NAND #() 
NAND_634_ (
  .A({ S1197 }),
  .B({ S1198 }),
  .Y({ S1199 })
);
NAND #() 
NAND_635_ (
  .A({ S435 }),
  .B({ S1199 }),
  .Y({ S1200 })
);
NAND #() 
NAND_636_ (
  .A({ datapath_theregisterfile_memtrf_0 }),
  .B({ S442 }),
  .Y({ S1201 })
);
NAND #() 
NAND_637_ (
  .A({ datapath_theregisterfile_memtrf_32 }),
  .B({ S441 }),
  .Y({ S1202 })
);
NAND #() 
NAND_638_ (
  .A({ S1201 }),
  .B({ S1202 }),
  .Y({ S1203 })
);
NAND #() 
NAND_639_ (
  .A({ S436 }),
  .B({ S1203 }),
  .Y({ S1204 })
);
NAND #() 
NAND_640_ (
  .A({ S1200 }),
  .B({ S1204 }),
  .Y({ S1205 })
);
NAND #() 
NAND_641_ (
  .A({ S429 }),
  .B({ S1205 }),
  .Y({ S1206 })
);
NAND #() 
NAND_642_ (
  .A({ S7520 }),
  .B({ S436 }),
  .Y({ S1207 })
);
NOR #() 
NOR_241_ (
  .A({ datapath_theregisterfile_memtrf_112 }),
  .B({ S436 }),
  .Y({ S1208 })
);
NOR #() 
NOR_242_ (
  .A({ S442 }),
  .B({ S1208 }),
  .Y({ S1209 })
);
NAND #() 
NAND_643_ (
  .A({ S1207 }),
  .B({ S1209 }),
  .Y({ S1210 })
);
NOR #() 
NOR_243_ (
  .A({ datapath_theregisterfile_memtrf_64 }),
  .B({ S435 }),
  .Y({ S1211 })
);
NOR #() 
NOR_244_ (
  .A({ datapath_theregisterfile_memtrf_80 }),
  .B({ S436 }),
  .Y({ S1212 })
);
NOR #() 
NOR_245_ (
  .A({ S1211 }),
  .B({ S1212 }),
  .Y({ S1213 })
);
NAND #() 
NAND_644_ (
  .A({ S442 }),
  .B({ S1213 }),
  .Y({ S1214 })
);
NAND #() 
NAND_645_ (
  .A({ S1210 }),
  .B({ S1214 }),
  .Y({ S1215 })
);
NAND #() 
NAND_646_ (
  .A({ S479 }),
  .B({ S1215 }),
  .Y({ S1216 })
);
NAND #() 
NAND_647_ (
  .A({ S1206 }),
  .B({ S1216 }),
  .Y({ S1217 })
);
NOR #() 
NOR_246_ (
  .A({ S1196 }),
  .B({ S1217 }),
  .Y({ S1218 })
);
NAND #() 
NAND_648_ (
  .A({ S446 }),
  .B({ S1218 }),
  .Y({ S1219 })
);
NAND #() 
NAND_649_ (
  .A({ S1174 }),
  .B({ S1219 }),
  .Y({ S1220 })
);
NOT #() 
NOT_154_ (
  .A({ S1220 }),
  .Y({ datapath_addsubunit_in1_0 })
);
NAND #() 
NAND_650_ (
  .A({ S496 }),
  .B({ datapath_addsubunit_in1_0 }),
  .Y({ S1221 })
);
NAND #() 
NAND_651_ (
  .A({ S1173 }),
  .B({ S1221 }),
  .Y({ S1222 })
);
NAND #() 
NAND_652_ (
  .A({ datapath_muxmem_in2_0 }),
  .B({ S1222 }),
  .Y({ S1223 })
);
NOT #() 
NOT_155_ (
  .A({ S1223 }),
  .Y({ S1224 })
);
NOR #() 
NOR_247_ (
  .A({ datapath_muxmem_in2_1 }),
  .B({ S1170 }),
  .Y({ S1225 })
);
NOR #() 
NOR_248_ (
  .A({ S1172 }),
  .B({ S1225 }),
  .Y({ S1226 })
);
NAND #() 
NAND_653_ (
  .A({ S1224 }),
  .B({ S1226 }),
  .Y({ S1227 })
);
NOT #() 
NOT_156_ (
  .A({ S1227 }),
  .Y({ S1228 })
);
NAND #() 
NAND_654_ (
  .A({ S1171 }),
  .B({ S1227 }),
  .Y({ S1229 })
);
NOR #() 
NOR_249_ (
  .A({ datapath_muxmem_in2_2 }),
  .B({ S1118 }),
  .Y({ S1230 })
);
NOR #() 
NOR_250_ (
  .A({ S1120 }),
  .B({ S1230 }),
  .Y({ S1231 })
);
NAND #() 
NAND_655_ (
  .A({ S1229 }),
  .B({ S1231 }),
  .Y({ S1232 })
);
NAND #() 
NAND_656_ (
  .A({ S1119 }),
  .B({ S1232 }),
  .Y({ S1233 })
);
NOR #() 
NOR_251_ (
  .A({ S1069 }),
  .B({ S1233 }),
  .Y({ S1234 })
);
NOR #() 
NOR_252_ (
  .A({ S1070 }),
  .B({ S1234 }),
  .Y({ S1235 })
);
NAND #() 
NAND_657_ (
  .A({ S1019 }),
  .B({ S1235 }),
  .Y({ S1236 })
);
NAND #() 
NAND_658_ (
  .A({ S1016 }),
  .B({ S1236 }),
  .Y({ S1237 })
);
NOR #() 
NOR_253_ (
  .A({ S967 }),
  .B({ S1237 }),
  .Y({ S1238 })
);
NOR #() 
NOR_254_ (
  .A({ S968 }),
  .B({ S1238 }),
  .Y({ S1239 })
);
NAND #() 
NAND_659_ (
  .A({ S916 }),
  .B({ S1239 }),
  .Y({ S1240 })
);
NAND #() 
NAND_660_ (
  .A({ S913 }),
  .B({ S1240 }),
  .Y({ S1241 })
);
NOR #() 
NOR_255_ (
  .A({ S862 }),
  .B({ S1241 }),
  .Y({ S1242 })
);
NOR #() 
NOR_256_ (
  .A({ S863 }),
  .B({ S1242 }),
  .Y({ S1243 })
);
NAND #() 
NAND_661_ (
  .A({ S811 }),
  .B({ S1243 }),
  .Y({ S1244 })
);
NAND #() 
NAND_662_ (
  .A({ S808 }),
  .B({ S1244 }),
  .Y({ S1245 })
);
NOR #() 
NOR_257_ (
  .A({ S758 }),
  .B({ S1245 }),
  .Y({ S1246 })
);
NOR #() 
NOR_258_ (
  .A({ S759 }),
  .B({ S1246 }),
  .Y({ S1247 })
);
NAND #() 
NAND_663_ (
  .A({ S708 }),
  .B({ S1247 }),
  .Y({ S1248 })
);
NAND #() 
NAND_664_ (
  .A({ S705 }),
  .B({ S1248 }),
  .Y({ S1249 })
);
NOR #() 
NOR_259_ (
  .A({ S655 }),
  .B({ S1249 }),
  .Y({ S1250 })
);
NOR #() 
NOR_260_ (
  .A({ S656 }),
  .B({ S1250 }),
  .Y({ S1251 })
);
NAND #() 
NAND_665_ (
  .A({ S605 }),
  .B({ S1251 }),
  .Y({ S1252 })
);
NAND #() 
NAND_666_ (
  .A({ S602 }),
  .B({ S1252 }),
  .Y({ S1253 })
);
NOR #() 
NOR_261_ (
  .A({ S553 }),
  .B({ S1253 }),
  .Y({ S1254 })
);
NOR #() 
NOR_262_ (
  .A({ S552 }),
  .B({ S1254 }),
  .Y({ S1255 })
);
NAND #() 
NAND_667_ (
  .A({ S502 }),
  .B({ S1255 }),
  .Y({ S1256 })
);
NAND #() 
NAND_668_ (
  .A({ S499 }),
  .B({ S1256 }),
  .Y({ S1257 })
);
NOT #() 
NOT_157_ (
  .A({ S1257 }),
  .Y({ S1258 })
);
NAND #() 
NAND_669_ (
  .A({ S7574 }),
  .B({ S423 }),
  .Y({ S1259 })
);
NOR #() 
NOR_263_ (
  .A({ datapath_theregisterfile_memtrf_239 }),
  .B({ S423 }),
  .Y({ S1260 })
);
NOR #() 
NOR_264_ (
  .A({ S435 }),
  .B({ S1260 }),
  .Y({ S1261 })
);
NAND #() 
NAND_670_ (
  .A({ S1259 }),
  .B({ S1261 }),
  .Y({ S1262 })
);
NOR #() 
NOR_265_ (
  .A({ datapath_theregisterfile_memtrf_255 }),
  .B({ S423 }),
  .Y({ S1263 })
);
NAND #() 
NAND_671_ (
  .A({ S7662 }),
  .B({ S423 }),
  .Y({ S1264 })
);
NAND #() 
NAND_672_ (
  .A({ S435 }),
  .B({ S1264 }),
  .Y({ S1265 })
);
NOR #() 
NOR_266_ (
  .A({ S1263 }),
  .B({ S1265 }),
  .Y({ S1266 })
);
NAND #() 
NAND_673_ (
  .A({ datapath_theregisterfile_memtrf_207 }),
  .B({ S436 }),
  .Y({ S1267 })
);
NAND #() 
NAND_674_ (
  .A({ datapath_theregisterfile_memtrf_223 }),
  .B({ S435 }),
  .Y({ S1268 })
);
NAND #() 
NAND_675_ (
  .A({ S1267 }),
  .B({ S1268 }),
  .Y({ S1269 })
);
NAND #() 
NAND_676_ (
  .A({ S422 }),
  .B({ S1269 }),
  .Y({ S1270 })
);
NAND #() 
NAND_677_ (
  .A({ datapath_theregisterfile_memtrf_143 }),
  .B({ S436 }),
  .Y({ S1271 })
);
NAND #() 
NAND_678_ (
  .A({ datapath_theregisterfile_memtrf_159 }),
  .B({ S435 }),
  .Y({ S1272 })
);
NAND #() 
NAND_679_ (
  .A({ S1271 }),
  .B({ S1272 }),
  .Y({ S1273 })
);
NAND #() 
NAND_680_ (
  .A({ S423 }),
  .B({ S1273 }),
  .Y({ S1274 })
);
NAND #() 
NAND_681_ (
  .A({ S1270 }),
  .B({ S1274 }),
  .Y({ S1275 })
);
NOR #() 
NOR_267_ (
  .A({ S441 }),
  .B({ S1275 }),
  .Y({ S1276 })
);
NOR #() 
NOR_268_ (
  .A({ S442 }),
  .B({ S1266 }),
  .Y({ S1277 })
);
NAND #() 
NAND_682_ (
  .A({ S1262 }),
  .B({ S1277 }),
  .Y({ S1278 })
);
NAND #() 
NAND_683_ (
  .A({ S428 }),
  .B({ S1278 }),
  .Y({ S1279 })
);
NOR #() 
NOR_269_ (
  .A({ S1276 }),
  .B({ S1279 }),
  .Y({ S1280 })
);
NAND #() 
NAND_684_ (
  .A({ datapath_theregisterfile_memtrf_127 }),
  .B({ S435 }),
  .Y({ S1281 })
);
NAND #() 
NAND_685_ (
  .A({ datapath_theregisterfile_memtrf_111 }),
  .B({ S436 }),
  .Y({ S1282 })
);
NAND #() 
NAND_686_ (
  .A({ S1281 }),
  .B({ S1282 }),
  .Y({ S1283 })
);
NAND #() 
NAND_687_ (
  .A({ S441 }),
  .B({ S1283 }),
  .Y({ S1284 })
);
NAND #() 
NAND_688_ (
  .A({ datapath_theregisterfile_memtrf_95 }),
  .B({ S435 }),
  .Y({ S1285 })
);
NAND #() 
NAND_689_ (
  .A({ datapath_theregisterfile_memtrf_79 }),
  .B({ S436 }),
  .Y({ S1286 })
);
NAND #() 
NAND_690_ (
  .A({ S1285 }),
  .B({ S1286 }),
  .Y({ S1287 })
);
NAND #() 
NAND_691_ (
  .A({ S442 }),
  .B({ S1287 }),
  .Y({ S1288 })
);
NAND #() 
NAND_692_ (
  .A({ S1284 }),
  .B({ S1288 }),
  .Y({ S1289 })
);
NAND #() 
NAND_693_ (
  .A({ S479 }),
  .B({ S1289 }),
  .Y({ S1290 })
);
NAND #() 
NAND_694_ (
  .A({ datapath_theregisterfile_memtrf_63 }),
  .B({ S435 }),
  .Y({ S1291 })
);
NAND #() 
NAND_695_ (
  .A({ datapath_theregisterfile_memtrf_47 }),
  .B({ S436 }),
  .Y({ S1292 })
);
NAND #() 
NAND_696_ (
  .A({ S1291 }),
  .B({ S1292 }),
  .Y({ S1293 })
);
NAND #() 
NAND_697_ (
  .A({ S441 }),
  .B({ S1293 }),
  .Y({ S1294 })
);
NAND #() 
NAND_698_ (
  .A({ datapath_theregisterfile_memtrf_31 }),
  .B({ S435 }),
  .Y({ S1295 })
);
NAND #() 
NAND_699_ (
  .A({ datapath_theregisterfile_memtrf_15 }),
  .B({ S436 }),
  .Y({ S1296 })
);
NAND #() 
NAND_700_ (
  .A({ S1295 }),
  .B({ S1296 }),
  .Y({ S1297 })
);
NAND #() 
NAND_701_ (
  .A({ S442 }),
  .B({ S1297 }),
  .Y({ S1298 })
);
NAND #() 
NAND_702_ (
  .A({ S1294 }),
  .B({ S1298 }),
  .Y({ S1299 })
);
NAND #() 
NAND_703_ (
  .A({ S429 }),
  .B({ S1299 }),
  .Y({ S1300 })
);
NOT #() 
NOT_158_ (
  .A({ S1300 }),
  .Y({ S1301 })
);
NOR #() 
NOR_270_ (
  .A({ S1280 }),
  .B({ S1301 }),
  .Y({ S1302 })
);
NAND #() 
NAND_704_ (
  .A({ S1290 }),
  .B({ S1302 }),
  .Y({ S1303 })
);
NAND #() 
NAND_705_ (
  .A({ S446 }),
  .B({ S1303 }),
  .Y({ S1304 })
);
NOT #() 
NOT_159_ (
  .A({ S1304 }),
  .Y({ datapath_addsubunit_in1_15 })
);
NAND #() 
NAND_706_ (
  .A({ S496 }),
  .B({ datapath_addsubunit_in1_15 }),
  .Y({ S1305 })
);
NAND #() 
NAND_707_ (
  .A({ S372 }),
  .B({ S1305 }),
  .Y({ S1306 })
);
NAND #() 
NAND_708_ (
  .A({ datapath_muxmem_in2_15 }),
  .B({ S1306 }),
  .Y({ S1307 })
);
NOT #() 
NOT_160_ (
  .A({ S1307 }),
  .Y({ S1308 })
);
NOR #() 
NOR_271_ (
  .A({ datapath_muxmem_in2_15 }),
  .B({ S1306 }),
  .Y({ S1309 })
);
NOT #() 
NOT_161_ (
  .A({ S1309 }),
  .Y({ S1310 })
);
NOR #() 
NOR_272_ (
  .A({ S1308 }),
  .B({ S1309 }),
  .Y({ S1311 })
);
NAND #() 
NAND_709_ (
  .A({ S1307 }),
  .B({ S1310 }),
  .Y({ S1312 })
);
NAND #() 
NAND_710_ (
  .A({ S1258 }),
  .B({ S1311 }),
  .Y({ S1313 })
);
NAND #() 
NAND_711_ (
  .A({ S1257 }),
  .B({ S1312 }),
  .Y({ S1314 })
);
NAND #() 
NAND_712_ (
  .A({ S1313 }),
  .B({ S1314 }),
  .Y({ S1315 })
);
NAND #() 
NAND_713_ (
  .A({ S365 }),
  .B({ S1315 }),
  .Y({ S1316 })
);
NOR #() 
NOR_273_ (
  .A({ controller_389_B_0 }),
  .B({ S348 }),
  .Y({ S1317 })
);
NOR #() 
NOR_274_ (
  .A({ S346 }),
  .B({ S1317 }),
  .Y({ S1318 })
);
NOR #() 
NOR_275_ (
  .A({ S8587 }),
  .B({ S1318 }),
  .Y({ S1319 })
);
NAND #() 
NAND_714_ (
  .A({ S8587 }),
  .B({ S344 }),
  .Y({ S1320 })
);
NOR #() 
NOR_276_ (
  .A({ S8225 }),
  .B({ S1320 }),
  .Y({ S1321 })
);
NAND #() 
NAND_715_ (
  .A({ S8586 }),
  .B({ S8588 }),
  .Y({ S1322 })
);
NOR #() 
NOR_277_ (
  .A({ controller_389_B_0 }),
  .B({ S353 }),
  .Y({ S1323 })
);
NAND #() 
NAND_716_ (
  .A({ controller_389_B_0 }),
  .B({ S8584 }),
  .Y({ S1324 })
);
NOR #() 
NOR_278_ (
  .A({ S1321 }),
  .B({ S1323 }),
  .Y({ S1325 })
);
NAND #() 
NAND_717_ (
  .A({ S1322 }),
  .B({ S1324 }),
  .Y({ S1326 })
);
NOR #() 
NOR_279_ (
  .A({ S8551 }),
  .B({ S1326 }),
  .Y({ S1327 })
);
NAND #() 
NAND_718_ (
  .A({ S1325 }),
  .B({ S1327 }),
  .Y({ S1328 })
);
NOR #() 
NOR_280_ (
  .A({ S1319 }),
  .B({ S1328 }),
  .Y({ S1329 })
);
NOR #() 
NOR_281_ (
  .A({ S8554 }),
  .B({ S1329 }),
  .Y({ S1330 })
);
NOR #() 
NOR_282_ (
  .A({ S8549 }),
  .B({ S1330 }),
  .Y({ S1331 })
);
NOR #() 
NOR_283_ (
  .A({ S8385 }),
  .B({ S1331 }),
  .Y({ S1332 })
);
NAND #() 
NAND_719_ (
  .A({ S8571 }),
  .B({ S8577 }),
  .Y({ S1333 })
);
NOR #() 
NOR_284_ (
  .A({ S1332 }),
  .B({ S1333 }),
  .Y({ S1334 })
);
NOR #() 
NOR_285_ (
  .A({ S7884 }),
  .B({ S7892 }),
  .Y({ S1335 })
);
NAND #() 
NAND_720_ (
  .A({ datapath_muxmem_in2_0 }),
  .B({ datapath_muxmem_in2_1 }),
  .Y({ S1336 })
);
NOR #() 
NOR_286_ (
  .A({ S7897 }),
  .B({ S1336 }),
  .Y({ S1337 })
);
NAND #() 
NAND_721_ (
  .A({ datapath_muxmem_in2_2 }),
  .B({ S1335 }),
  .Y({ S1338 })
);
NOR #() 
NOR_287_ (
  .A({ S7905 }),
  .B({ S1338 }),
  .Y({ S1339 })
);
NAND #() 
NAND_722_ (
  .A({ datapath_muxmem_in2_3 }),
  .B({ S1337 }),
  .Y({ S1340 })
);
NAND #() 
NAND_723_ (
  .A({ datapath_muxmem_in2_4 }),
  .B({ S1339 }),
  .Y({ S1341 })
);
NOT #() 
NOT_162_ (
  .A({ S1341 }),
  .Y({ S1342 })
);
NOR #() 
NOR_288_ (
  .A({ S7920 }),
  .B({ S1341 }),
  .Y({ S1343 })
);
NAND #() 
NAND_724_ (
  .A({ datapath_muxmem_in2_5 }),
  .B({ S1342 }),
  .Y({ S1344 })
);
NOR #() 
NOR_289_ (
  .A({ S7928 }),
  .B({ S1344 }),
  .Y({ S1345 })
);
NAND #() 
NAND_725_ (
  .A({ datapath_muxmem_in2_6 }),
  .B({ S1343 }),
  .Y({ S1346 })
);
NAND #() 
NAND_726_ (
  .A({ datapath_muxmem_in2_7 }),
  .B({ S1345 }),
  .Y({ S1347 })
);
NOT #() 
NOT_163_ (
  .A({ S1347 }),
  .Y({ S1348 })
);
NOR #() 
NOR_290_ (
  .A({ S7946 }),
  .B({ S1347 }),
  .Y({ S1349 })
);
NAND #() 
NAND_727_ (
  .A({ datapath_muxmem_in2_8 }),
  .B({ S1348 }),
  .Y({ S1350 })
);
NOR #() 
NOR_291_ (
  .A({ S7957 }),
  .B({ S1350 }),
  .Y({ S1351 })
);
NAND #() 
NAND_728_ (
  .A({ datapath_muxmem_in2_9 }),
  .B({ S1349 }),
  .Y({ S1352 })
);
NOR #() 
NOR_292_ (
  .A({ S7968 }),
  .B({ S1352 }),
  .Y({ S1353 })
);
NAND #() 
NAND_729_ (
  .A({ datapath_muxmem_in2_10 }),
  .B({ S1351 }),
  .Y({ S1354 })
);
NOR #() 
NOR_293_ (
  .A({ S7978 }),
  .B({ S1354 }),
  .Y({ S1355 })
);
NAND #() 
NAND_730_ (
  .A({ datapath_muxmem_in2_11 }),
  .B({ S1353 }),
  .Y({ S1356 })
);
NOR #() 
NOR_294_ (
  .A({ S7989 }),
  .B({ S1356 }),
  .Y({ S1357 })
);
NAND #() 
NAND_731_ (
  .A({ datapath_muxmem_in2_12 }),
  .B({ S1355 }),
  .Y({ S1358 })
);
NOR #() 
NOR_295_ (
  .A({ S8000 }),
  .B({ S1358 }),
  .Y({ S1359 })
);
NAND #() 
NAND_732_ (
  .A({ datapath_muxmem_in2_14 }),
  .B({ S1359 }),
  .Y({ S1360 })
);
NAND #() 
NAND_733_ (
  .A({ datapath_muxmem_in2_15 }),
  .B({ S1360 }),
  .Y({ S1361 })
);
NOR #() 
NOR_296_ (
  .A({ datapath_muxmem_in2_15 }),
  .B({ S1360 }),
  .Y({ S1362 })
);
NOT #() 
NOT_164_ (
  .A({ S1362 }),
  .Y({ S1363 })
);
NAND #() 
NAND_734_ (
  .A({ S1361 }),
  .B({ S1363 }),
  .Y({ S1364 })
);
NOT #() 
NOT_165_ (
  .A({ S1364 }),
  .Y({ S1365 })
);
NOR #() 
NOR_297_ (
  .A({ S1334 }),
  .B({ S1365 }),
  .Y({ S1366 })
);
NAND #() 
NAND_735_ (
  .A({ controller_216_B_0 }),
  .B({ S8585 }),
  .Y({ S1367 })
);
NAND #() 
NAND_736_ (
  .A({ S379 }),
  .B({ S1367 }),
  .Y({ S1368 })
);
NOT #() 
NOT_166_ (
  .A({ S1368 }),
  .Y({ S1369 })
);
NOR #() 
NOR_298_ (
  .A({ S358 }),
  .B({ S1368 }),
  .Y({ S1370 })
);
NAND #() 
NAND_737_ (
  .A({ S359 }),
  .B({ S1369 }),
  .Y({ S1371 })
);
NOR #() 
NOR_299_ (
  .A({ S1366 }),
  .B({ S1370 }),
  .Y({ S1372 })
);
NAND #() 
NAND_738_ (
  .A({ S1316 }),
  .B({ S1372 }),
  .Y({ S1373 })
);
NOR #() 
NOR_300_ (
  .A({ datapath_addsubunit_in1_15 }),
  .B({ S1371 }),
  .Y({ S1374 })
);
NOR #() 
NOR_301_ (
  .A({ S8580 }),
  .B({ S1374 }),
  .Y({ S1375 })
);
NAND #() 
NAND_739_ (
  .A({ S1373 }),
  .B({ S1375 }),
  .Y({ S1376 })
);
NAND #() 
NAND_740_ (
  .A({ S8581 }),
  .B({ S1376 }),
  .Y({ S0 })
);
NOR #() 
NOR_302_ (
  .A({ controller_pstate_0 }),
  .B({ S8569 }),
  .Y({ S1377 })
);
NAND #() 
NAND_741_ (
  .A({ S8365 }),
  .B({ S8568 }),
  .Y({ S1378 })
);
NOR #() 
NOR_303_ (
  .A({ S7476 }),
  .B({ S1377 }),
  .Y({ S1 })
);
NAND #() 
NAND_742_ (
  .A({ S8356 }),
  .B({ S8365 }),
  .Y({ S1379 })
);
NOT #() 
NOT_167_ (
  .A({ S1379 }),
  .Y({ controller_1115_S_0 })
);
NAND #() 
NAND_743_ (
  .A({ datapath_databusin_15 }),
  .B({ controller_1115_S_0 }),
  .Y({ S1380 })
);
NAND #() 
NAND_744_ (
  .A({ controller_opcode_7 }),
  .B({ S1379 }),
  .Y({ S1381 })
);
NAND #() 
NAND_745_ (
  .A({ S1380 }),
  .B({ S1381 }),
  .Y({ S2 })
);
NOR #() 
NOR_304_ (
  .A({ controller_opcode_3 }),
  .B({ S369 }),
  .Y({ S1382 })
);
NAND #() 
NAND_746_ (
  .A({ S8309 }),
  .B({ S368 }),
  .Y({ S1383 })
);
NAND #() 
NAND_747_ (
  .A({ datapath_adr_outreg_15 }),
  .B({ S1383 }),
  .Y({ S1384 })
);
NAND #() 
NAND_748_ (
  .A({ S1306 }),
  .B({ S1382 }),
  .Y({ S1385 })
);
NAND #() 
NAND_749_ (
  .A({ S1384 }),
  .B({ S1385 }),
  .Y({ S3 })
);
NOR #() 
NOR_305_ (
  .A({ S8385 }),
  .B({ S383 }),
  .Y({ S1386 })
);
NAND #() 
NAND_750_ (
  .A({ S8375 }),
  .B({ S382 }),
  .Y({ S1387 })
);
NOR #() 
NOR_306_ (
  .A({ S8557 }),
  .B({ S1387 }),
  .Y({ S1388 })
);
NAND #() 
NAND_751_ (
  .A({ S8375 }),
  .B({ S384 }),
  .Y({ S1389 })
);
NOR #() 
NOR_307_ (
  .A({ S1220 }),
  .B({ S1389 }),
  .Y({ S1390 })
);
NOR #() 
NOR_308_ (
  .A({ S8319 }),
  .B({ controller_opcode_5 }),
  .Y({ S1391 })
);
NOT #() 
NOT_168_ (
  .A({ S1391 }),
  .Y({ S1392 })
);
NAND #() 
NAND_752_ (
  .A({ S382 }),
  .B({ S1391 }),
  .Y({ S1393 })
);
NAND #() 
NAND_753_ (
  .A({ S410 }),
  .B({ S1393 }),
  .Y({ S1394 })
);
NOR #() 
NOR_309_ (
  .A({ S389 }),
  .B({ S1394 }),
  .Y({ S1395 })
);
NOR #() 
NOR_310_ (
  .A({ S8385 }),
  .B({ S1395 }),
  .Y({ S1396 })
);
NOT #() 
NOT_169_ (
  .A({ S1396 }),
  .Y({ S1397 })
);
NAND #() 
NAND_754_ (
  .A({ S8375 }),
  .B({ S8416 }),
  .Y({ S1398 })
);
NAND #() 
NAND_755_ (
  .A({ S8416 }),
  .B({ S1386 }),
  .Y({ S1399 })
);
NOT #() 
NOT_170_ (
  .A({ S1399 }),
  .Y({ S1400 })
);
NAND #() 
NAND_756_ (
  .A({ S1397 }),
  .B({ S1399 }),
  .Y({ S1401 })
);
NOR #() 
NOR_311_ (
  .A({ controller_opcode_2 }),
  .B({ controller_opcode_3 }),
  .Y({ S1402 })
);
NAND #() 
NAND_757_ (
  .A({ S8299 }),
  .B({ S8309 }),
  .Y({ S1403 })
);
NOR #() 
NOR_312_ (
  .A({ S380 }),
  .B({ S1403 }),
  .Y({ S1404 })
);
NAND #() 
NAND_758_ (
  .A({ S379 }),
  .B({ S1402 }),
  .Y({ S1405 })
);
NOR #() 
NOR_313_ (
  .A({ S8278 }),
  .B({ S1405 }),
  .Y({ S1406 })
);
NOT #() 
NOT_171_ (
  .A({ S1406 }),
  .Y({ S1407 })
);
NOR #() 
NOR_314_ (
  .A({ S1401 }),
  .B({ S1406 }),
  .Y({ S1408 })
);
NAND #() 
NAND_759_ (
  .A({ S371 }),
  .B({ S1408 }),
  .Y({ S1409 })
);
NAND #() 
NAND_760_ (
  .A({ controller_fib_0 }),
  .B({ S1409 }),
  .Y({ S1410 })
);
NOT #() 
NOT_172_ (
  .A({ S1410 }),
  .Y({ S1411 })
);
NOR #() 
NOR_315_ (
  .A({ S1390 }),
  .B({ S1411 }),
  .Y({ S1412 })
);
NOT #() 
NOT_173_ (
  .A({ S1412 }),
  .Y({ S1413 })
);
NAND #() 
NAND_761_ (
  .A({ S8375 }),
  .B({ S392 }),
  .Y({ S1414 })
);
NOT #() 
NOT_174_ (
  .A({ S1414 }),
  .Y({ S1415 })
);
NOR #() 
NOR_316_ (
  .A({ S1406 }),
  .B({ S1415 }),
  .Y({ S1416 })
);
NAND #() 
NAND_762_ (
  .A({ S1407 }),
  .B({ S1414 }),
  .Y({ S1417 })
);
NAND #() 
NAND_763_ (
  .A({ S1413 }),
  .B({ S1417 }),
  .Y({ S1418 })
);
NOR #() 
NOR_317_ (
  .A({ S401 }),
  .B({ S1403 }),
  .Y({ S1419 })
);
NAND #() 
NAND_764_ (
  .A({ S400 }),
  .B({ S1402 }),
  .Y({ S1420 })
);
NAND #() 
NAND_765_ (
  .A({ S8457 }),
  .B({ S8478 }),
  .Y({ S1421 })
);
NOR #() 
NOR_318_ (
  .A({ S8557 }),
  .B({ S387 }),
  .Y({ S1422 })
);
NOT #() 
NOT_175_ (
  .A({ S1422 }),
  .Y({ S1423 })
);
NOR #() 
NOR_319_ (
  .A({ S8565 }),
  .B({ S387 }),
  .Y({ S1424 })
);
NAND #() 
NAND_766_ (
  .A({ S1420 }),
  .B({ S1421 }),
  .Y({ S1425 })
);
NOR #() 
NOR_320_ (
  .A({ S1419 }),
  .B({ S1424 }),
  .Y({ S1426 })
);
NOR #() 
NOR_321_ (
  .A({ S1424 }),
  .B({ S1425 }),
  .Y({ S1427 })
);
NAND #() 
NAND_767_ (
  .A({ S1421 }),
  .B({ S1426 }),
  .Y({ S1428 })
);
NOR #() 
NOR_322_ (
  .A({ S8385 }),
  .B({ S1427 }),
  .Y({ S1429 })
);
NAND #() 
NAND_768_ (
  .A({ S8375 }),
  .B({ S1428 }),
  .Y({ S1430 })
);
NOR #() 
NOR_323_ (
  .A({ S8385 }),
  .B({ S1420 }),
  .Y({ S1431 })
);
NAND #() 
NAND_769_ (
  .A({ S8375 }),
  .B({ S1419 }),
  .Y({ S1432 })
);
NOR #() 
NOR_324_ (
  .A({ S8193 }),
  .B({ S1432 }),
  .Y({ S1433 })
);
NAND #() 
NAND_770_ (
  .A({ datapath_instruction_2 }),
  .B({ S1431 }),
  .Y({ S1434 })
);
NOR #() 
NOR_325_ (
  .A({ S8299 }),
  .B({ S415 }),
  .Y({ S1435 })
);
NAND #() 
NAND_771_ (
  .A({ controller_opcode_2 }),
  .B({ S414 }),
  .Y({ S1436 })
);
NOR #() 
NOR_326_ (
  .A({ S1433 }),
  .B({ S1435 }),
  .Y({ S1437 })
);
NAND #() 
NAND_772_ (
  .A({ S1434 }),
  .B({ S1436 }),
  .Y({ S1438 })
);
NAND #() 
NAND_773_ (
  .A({ datapath_instruction_1 }),
  .B({ S1431 }),
  .Y({ S1439 })
);
NOT #() 
NOT_176_ (
  .A({ S1439 }),
  .Y({ S1440 })
);
NAND #() 
NAND_774_ (
  .A({ controller_216_B_0 }),
  .B({ S414 }),
  .Y({ S1441 })
);
NOT #() 
NOT_177_ (
  .A({ S1441 }),
  .Y({ S1442 })
);
NOR #() 
NOR_327_ (
  .A({ S1440 }),
  .B({ S1442 }),
  .Y({ S1443 })
);
NAND #() 
NAND_775_ (
  .A({ S1439 }),
  .B({ S1441 }),
  .Y({ S1444 })
);
NAND #() 
NAND_776_ (
  .A({ datapath_instruction_3 }),
  .B({ S1431 }),
  .Y({ S1445 })
);
NOT #() 
NOT_178_ (
  .A({ S1445 }),
  .Y({ S1446 })
);
NAND #() 
NAND_777_ (
  .A({ controller_opcode_3 }),
  .B({ S414 }),
  .Y({ S1447 })
);
NOT #() 
NOT_179_ (
  .A({ S1447 }),
  .Y({ S1448 })
);
NOR #() 
NOR_328_ (
  .A({ S1446 }),
  .B({ S1448 }),
  .Y({ S1449 })
);
NAND #() 
NAND_778_ (
  .A({ S1445 }),
  .B({ S1447 }),
  .Y({ S1450 })
);
NOR #() 
NOR_329_ (
  .A({ S1443 }),
  .B({ S1449 }),
  .Y({ S1451 })
);
NAND #() 
NAND_779_ (
  .A({ S1444 }),
  .B({ S1450 }),
  .Y({ S1452 })
);
NAND #() 
NAND_780_ (
  .A({ datapath_instruction_0 }),
  .B({ S1431 }),
  .Y({ S1453 })
);
NOT #() 
NOT_180_ (
  .A({ S1453 }),
  .Y({ S1454 })
);
NAND #() 
NAND_781_ (
  .A({ controller_fib_4 }),
  .B({ S414 }),
  .Y({ S1455 })
);
NOT #() 
NOT_181_ (
  .A({ S1455 }),
  .Y({ S1456 })
);
NOR #() 
NOR_330_ (
  .A({ S1454 }),
  .B({ S1456 }),
  .Y({ S1457 })
);
NAND #() 
NAND_782_ (
  .A({ S1453 }),
  .B({ S1455 }),
  .Y({ S1458 })
);
NOR #() 
NOR_331_ (
  .A({ S1452 }),
  .B({ S1457 }),
  .Y({ S1459 })
);
NAND #() 
NAND_783_ (
  .A({ S1451 }),
  .B({ S1458 }),
  .Y({ S1460 })
);
NOR #() 
NOR_332_ (
  .A({ S1437 }),
  .B({ S1460 }),
  .Y({ S1461 })
);
NAND #() 
NAND_784_ (
  .A({ S1438 }),
  .B({ S1459 }),
  .Y({ S1462 })
);
NOR #() 
NOR_333_ (
  .A({ controller_outflag_0 }),
  .B({ S1462 }),
  .Y({ S1463 })
);
NOT #() 
NOT_182_ (
  .A({ S1463 }),
  .Y({ S1464 })
);
NAND #() 
NAND_785_ (
  .A({ datapath_theregisterfile_memtrf_240 }),
  .B({ S1437 }),
  .Y({ S1465 })
);
NAND #() 
NAND_786_ (
  .A({ datapath_theregisterfile_memtrf_176 }),
  .B({ S1438 }),
  .Y({ S1466 })
);
NAND #() 
NAND_787_ (
  .A({ S1465 }),
  .B({ S1466 }),
  .Y({ S1467 })
);
NAND #() 
NAND_788_ (
  .A({ S1457 }),
  .B({ S1467 }),
  .Y({ S1468 })
);
NAND #() 
NAND_789_ (
  .A({ S7783 }),
  .B({ S1437 }),
  .Y({ S1469 })
);
NOR #() 
NOR_334_ (
  .A({ datapath_theregisterfile_memtrf_160 }),
  .B({ S1437 }),
  .Y({ S1470 })
);
NAND #() 
NAND_790_ (
  .A({ S1458 }),
  .B({ S1469 }),
  .Y({ S1471 })
);
NOR #() 
NOR_335_ (
  .A({ S1470 }),
  .B({ S1471 }),
  .Y({ S1472 })
);
NAND #() 
NAND_791_ (
  .A({ datapath_theregisterfile_memtrf_208 }),
  .B({ S1437 }),
  .Y({ S1473 })
);
NAND #() 
NAND_792_ (
  .A({ datapath_theregisterfile_memtrf_144 }),
  .B({ S1438 }),
  .Y({ S1474 })
);
NAND #() 
NAND_793_ (
  .A({ S1473 }),
  .B({ S1474 }),
  .Y({ S1475 })
);
NAND #() 
NAND_794_ (
  .A({ S1457 }),
  .B({ S1475 }),
  .Y({ S1476 })
);
NOR #() 
NOR_336_ (
  .A({ datapath_theregisterfile_memtrf_128 }),
  .B({ S1437 }),
  .Y({ S1477 })
);
NOR #() 
NOR_337_ (
  .A({ datapath_theregisterfile_memtrf_192 }),
  .B({ S1438 }),
  .Y({ S1478 })
);
NOR #() 
NOR_338_ (
  .A({ S1477 }),
  .B({ S1478 }),
  .Y({ S1479 })
);
NAND #() 
NAND_795_ (
  .A({ S1458 }),
  .B({ S1479 }),
  .Y({ S1480 })
);
NAND #() 
NAND_796_ (
  .A({ S1476 }),
  .B({ S1480 }),
  .Y({ S1481 })
);
NOR #() 
NOR_339_ (
  .A({ S1443 }),
  .B({ S1481 }),
  .Y({ S1482 })
);
NOR #() 
NOR_340_ (
  .A({ S1444 }),
  .B({ S1472 }),
  .Y({ S1483 })
);
NAND #() 
NAND_797_ (
  .A({ S1468 }),
  .B({ S1483 }),
  .Y({ S1484 })
);
NAND #() 
NAND_798_ (
  .A({ S1449 }),
  .B({ S1484 }),
  .Y({ S1485 })
);
NOR #() 
NOR_341_ (
  .A({ S1482 }),
  .B({ S1485 }),
  .Y({ S1486 })
);
NOR #() 
NOR_342_ (
  .A({ S1444 }),
  .B({ S1449 }),
  .Y({ S1487 })
);
NAND #() 
NAND_799_ (
  .A({ datapath_theregisterfile_memtrf_48 }),
  .B({ S1438 }),
  .Y({ S1488 })
);
NAND #() 
NAND_800_ (
  .A({ datapath_theregisterfile_memtrf_112 }),
  .B({ S1437 }),
  .Y({ S1489 })
);
NAND #() 
NAND_801_ (
  .A({ S1488 }),
  .B({ S1489 }),
  .Y({ S1490 })
);
NAND #() 
NAND_802_ (
  .A({ S1457 }),
  .B({ S1490 }),
  .Y({ S1491 })
);
NAND #() 
NAND_803_ (
  .A({ datapath_theregisterfile_memtrf_96 }),
  .B({ S1437 }),
  .Y({ S1492 })
);
NAND #() 
NAND_804_ (
  .A({ datapath_theregisterfile_memtrf_32 }),
  .B({ S1438 }),
  .Y({ S1493 })
);
NAND #() 
NAND_805_ (
  .A({ S1492 }),
  .B({ S1493 }),
  .Y({ S1494 })
);
NAND #() 
NAND_806_ (
  .A({ S1458 }),
  .B({ S1494 }),
  .Y({ S1495 })
);
NAND #() 
NAND_807_ (
  .A({ S1491 }),
  .B({ S1495 }),
  .Y({ S1496 })
);
NAND #() 
NAND_808_ (
  .A({ S1487 }),
  .B({ S1496 }),
  .Y({ S1497 })
);
NOR #() 
NOR_343_ (
  .A({ S1438 }),
  .B({ S1458 }),
  .Y({ S1498 })
);
NAND #() 
NAND_809_ (
  .A({ datapath_theregisterfile_memtrf_80 }),
  .B({ S1498 }),
  .Y({ S1499 })
);
NAND #() 
NAND_810_ (
  .A({ datapath_theregisterfile_memtrf_16 }),
  .B({ S1438 }),
  .Y({ S1500 })
);
NAND #() 
NAND_811_ (
  .A({ S1499 }),
  .B({ S1500 }),
  .Y({ S1501 })
);
NOT #() 
NOT_183_ (
  .A({ S1501 }),
  .Y({ S1502 })
);
NOR #() 
NOR_344_ (
  .A({ S1452 }),
  .B({ S1502 }),
  .Y({ S1503 })
);
NAND #() 
NAND_812_ (
  .A({ S1451 }),
  .B({ S1501 }),
  .Y({ S1504 })
);
NOR #() 
NOR_345_ (
  .A({ datapath_theregisterfile_memtrf_64 }),
  .B({ S1438 }),
  .Y({ S1505 })
);
NOT #() 
NOT_184_ (
  .A({ S1505 }),
  .Y({ S1506 })
);
NOR #() 
NOR_346_ (
  .A({ S1460 }),
  .B({ S1505 }),
  .Y({ S1507 })
);
NAND #() 
NAND_813_ (
  .A({ S1459 }),
  .B({ S1506 }),
  .Y({ S1508 })
);
NOR #() 
NOR_347_ (
  .A({ S1503 }),
  .B({ S1507 }),
  .Y({ S1509 })
);
NAND #() 
NAND_814_ (
  .A({ S1504 }),
  .B({ S1508 }),
  .Y({ S1510 })
);
NAND #() 
NAND_815_ (
  .A({ S1497 }),
  .B({ S1509 }),
  .Y({ S1511 })
);
NOR #() 
NOR_348_ (
  .A({ S1486 }),
  .B({ S1510 }),
  .Y({ S1512 })
);
NOR #() 
NOR_349_ (
  .A({ S1486 }),
  .B({ S1511 }),
  .Y({ S1513 })
);
NAND #() 
NAND_816_ (
  .A({ S1497 }),
  .B({ S1512 }),
  .Y({ S1514 })
);
NOR #() 
NOR_350_ (
  .A({ S1463 }),
  .B({ S1513 }),
  .Y({ S1515 })
);
NAND #() 
NAND_817_ (
  .A({ S1464 }),
  .B({ S1514 }),
  .Y({ S1516 })
);
NAND #() 
NAND_818_ (
  .A({ S1429 }),
  .B({ S1515 }),
  .Y({ S1517 })
);
NAND #() 
NAND_819_ (
  .A({ S1418 }),
  .B({ S1517 }),
  .Y({ S1518 })
);
NOT #() 
NOT_185_ (
  .A({ S1518 }),
  .Y({ S1519 })
);
NOR #() 
NOR_351_ (
  .A({ datapath_addsubunit_in1_0 }),
  .B({ S1519 }),
  .Y({ S1520 })
);
NOR #() 
NOR_352_ (
  .A({ S1220 }),
  .B({ S1518 }),
  .Y({ S1521 })
);
NOR #() 
NOR_353_ (
  .A({ S1520 }),
  .B({ S1521 }),
  .Y({ S1522 })
);
NOR #() 
NOR_354_ (
  .A({ S409 }),
  .B({ S1422 }),
  .Y({ S1523 })
);
NAND #() 
NAND_820_ (
  .A({ S410 }),
  .B({ S1423 }),
  .Y({ S1524 })
);
NOR #() 
NOR_355_ (
  .A({ S8385 }),
  .B({ S1523 }),
  .Y({ S1525 })
);
NAND #() 
NAND_821_ (
  .A({ S8375 }),
  .B({ S1524 }),
  .Y({ S1526 })
);
NOR #() 
NOR_356_ (
  .A({ S378 }),
  .B({ S387 }),
  .Y({ S1527 })
);
NAND #() 
NAND_822_ (
  .A({ S8375 }),
  .B({ S388 }),
  .Y({ S1528 })
);
NOR #() 
NOR_357_ (
  .A({ S1525 }),
  .B({ S1527 }),
  .Y({ S1529 })
);
NOR #() 
NOR_358_ (
  .A({ S1522 }),
  .B({ S1529 }),
  .Y({ S1530 })
);
NAND #() 
NAND_823_ (
  .A({ datapath_addsubunit_in1_0 }),
  .B({ S1518 }),
  .Y({ S1531 })
);
NOR #() 
NOR_359_ (
  .A({ S8385 }),
  .B({ S1421 }),
  .Y({ S1532 })
);
NOR #() 
NOR_360_ (
  .A({ S1400 }),
  .B({ S1532 }),
  .Y({ S1533 })
);
NOT #() 
NOT_186_ (
  .A({ S1533 }),
  .Y({ S1534 })
);
NOR #() 
NOR_361_ (
  .A({ S1531 }),
  .B({ S1533 }),
  .Y({ S1535 })
);
NOT #() 
NOT_187_ (
  .A({ S1535 }),
  .Y({ S1536 })
);
NAND #() 
NAND_824_ (
  .A({ controller_opcode_3 }),
  .B({ S379 }),
  .Y({ S1537 })
);
NOR #() 
NOR_362_ (
  .A({ S366 }),
  .B({ S380 }),
  .Y({ S1538 })
);
NAND #() 
NAND_825_ (
  .A({ S367 }),
  .B({ S379 }),
  .Y({ S1539 })
);
NOR #() 
NOR_363_ (
  .A({ S8267 }),
  .B({ S1539 }),
  .Y({ S1540 })
);
NAND #() 
NAND_826_ (
  .A({ S1220 }),
  .B({ S1540 }),
  .Y({ S1541 })
);
NOT #() 
NOT_188_ (
  .A({ S1541 }),
  .Y({ S1542 })
);
NOR #() 
NOR_364_ (
  .A({ S1220 }),
  .B({ S1540 }),
  .Y({ S1543 })
);
NOR #() 
NOR_365_ (
  .A({ S1539 }),
  .B({ S1543 }),
  .Y({ S1544 })
);
NAND #() 
NAND_827_ (
  .A({ S1541 }),
  .B({ S1544 }),
  .Y({ S1545 })
);
NOR #() 
NOR_366_ (
  .A({ S8565 }),
  .B({ S1387 }),
  .Y({ S1546 })
);
NAND #() 
NAND_828_ (
  .A({ S8564 }),
  .B({ S1386 }),
  .Y({ S1547 })
);
NOR #() 
NOR_367_ (
  .A({ S1412 }),
  .B({ S1547 }),
  .Y({ S1548 })
);
NOR #() 
NOR_368_ (
  .A({ controller_389_B_0 }),
  .B({ S1462 }),
  .Y({ S1549 })
);
NOT #() 
NOT_189_ (
  .A({ S1549 }),
  .Y({ S1550 })
);
NAND #() 
NAND_829_ (
  .A({ datapath_theregisterfile_memtrf_244 }),
  .B({ S1437 }),
  .Y({ S1551 })
);
NAND #() 
NAND_830_ (
  .A({ datapath_theregisterfile_memtrf_180 }),
  .B({ S1438 }),
  .Y({ S1552 })
);
NAND #() 
NAND_831_ (
  .A({ S1551 }),
  .B({ S1552 }),
  .Y({ S1553 })
);
NAND #() 
NAND_832_ (
  .A({ S1457 }),
  .B({ S1553 }),
  .Y({ S1554 })
);
NAND #() 
NAND_833_ (
  .A({ S7816 }),
  .B({ S1437 }),
  .Y({ S1555 })
);
NOR #() 
NOR_369_ (
  .A({ datapath_theregisterfile_memtrf_164 }),
  .B({ S1437 }),
  .Y({ S1556 })
);
NAND #() 
NAND_834_ (
  .A({ S1458 }),
  .B({ S1555 }),
  .Y({ S1557 })
);
NOR #() 
NOR_370_ (
  .A({ S1556 }),
  .B({ S1557 }),
  .Y({ S1558 })
);
NAND #() 
NAND_835_ (
  .A({ datapath_theregisterfile_memtrf_148 }),
  .B({ S1438 }),
  .Y({ S1559 })
);
NAND #() 
NAND_836_ (
  .A({ datapath_theregisterfile_memtrf_212 }),
  .B({ S1437 }),
  .Y({ S1560 })
);
NAND #() 
NAND_837_ (
  .A({ S1559 }),
  .B({ S1560 }),
  .Y({ S1561 })
);
NAND #() 
NAND_838_ (
  .A({ S1457 }),
  .B({ S1561 }),
  .Y({ S1562 })
);
NOR #() 
NOR_371_ (
  .A({ datapath_theregisterfile_memtrf_132 }),
  .B({ S1437 }),
  .Y({ S1563 })
);
NOR #() 
NOR_372_ (
  .A({ datapath_theregisterfile_memtrf_196 }),
  .B({ S1438 }),
  .Y({ S1564 })
);
NOR #() 
NOR_373_ (
  .A({ S1563 }),
  .B({ S1564 }),
  .Y({ S1565 })
);
NAND #() 
NAND_839_ (
  .A({ S1458 }),
  .B({ S1565 }),
  .Y({ S1566 })
);
NAND #() 
NAND_840_ (
  .A({ S1562 }),
  .B({ S1566 }),
  .Y({ S1567 })
);
NOR #() 
NOR_374_ (
  .A({ S1443 }),
  .B({ S1567 }),
  .Y({ S1568 })
);
NOR #() 
NOR_375_ (
  .A({ S1444 }),
  .B({ S1558 }),
  .Y({ S1569 })
);
NAND #() 
NAND_841_ (
  .A({ S1554 }),
  .B({ S1569 }),
  .Y({ S1570 })
);
NAND #() 
NAND_842_ (
  .A({ S1449 }),
  .B({ S1570 }),
  .Y({ S1571 })
);
NOR #() 
NOR_376_ (
  .A({ S1568 }),
  .B({ S1571 }),
  .Y({ S1572 })
);
NAND #() 
NAND_843_ (
  .A({ datapath_theregisterfile_memtrf_100 }),
  .B({ S1458 }),
  .Y({ S1573 })
);
NAND #() 
NAND_844_ (
  .A({ datapath_theregisterfile_memtrf_116 }),
  .B({ S1457 }),
  .Y({ S1574 })
);
NAND #() 
NAND_845_ (
  .A({ S1573 }),
  .B({ S1574 }),
  .Y({ S1575 })
);
NAND #() 
NAND_846_ (
  .A({ S1437 }),
  .B({ S1575 }),
  .Y({ S1576 })
);
NAND #() 
NAND_847_ (
  .A({ datapath_theregisterfile_memtrf_36 }),
  .B({ S1458 }),
  .Y({ S1577 })
);
NAND #() 
NAND_848_ (
  .A({ datapath_theregisterfile_memtrf_52 }),
  .B({ S1457 }),
  .Y({ S1578 })
);
NAND #() 
NAND_849_ (
  .A({ S1577 }),
  .B({ S1578 }),
  .Y({ S1579 })
);
NAND #() 
NAND_850_ (
  .A({ S1438 }),
  .B({ S1579 }),
  .Y({ S1580 })
);
NAND #() 
NAND_851_ (
  .A({ S1576 }),
  .B({ S1580 }),
  .Y({ S1581 })
);
NAND #() 
NAND_852_ (
  .A({ S1487 }),
  .B({ S1581 }),
  .Y({ S1582 })
);
NAND #() 
NAND_853_ (
  .A({ datapath_theregisterfile_memtrf_84 }),
  .B({ S1498 }),
  .Y({ S1583 })
);
NOR #() 
NOR_377_ (
  .A({ datapath_theregisterfile_memtrf_68 }),
  .B({ S1438 }),
  .Y({ S1584 })
);
NOT #() 
NOT_190_ (
  .A({ S1584 }),
  .Y({ S1585 })
);
NAND #() 
NAND_854_ (
  .A({ datapath_theregisterfile_memtrf_20 }),
  .B({ S1438 }),
  .Y({ S1586 })
);
NAND #() 
NAND_855_ (
  .A({ S1457 }),
  .B({ S1586 }),
  .Y({ S1587 })
);
NAND #() 
NAND_856_ (
  .A({ S1585 }),
  .B({ S1587 }),
  .Y({ S1588 })
);
NAND #() 
NAND_857_ (
  .A({ S1583 }),
  .B({ S1588 }),
  .Y({ S1589 })
);
NOT #() 
NOT_191_ (
  .A({ S1589 }),
  .Y({ S1590 })
);
NOR #() 
NOR_378_ (
  .A({ S1452 }),
  .B({ S1590 }),
  .Y({ S1591 })
);
NAND #() 
NAND_858_ (
  .A({ S1451 }),
  .B({ S1589 }),
  .Y({ S1592 })
);
NAND #() 
NAND_859_ (
  .A({ S1582 }),
  .B({ S1592 }),
  .Y({ S1593 })
);
NOR #() 
NOR_379_ (
  .A({ S1572 }),
  .B({ S1591 }),
  .Y({ S1594 })
);
NOR #() 
NOR_380_ (
  .A({ S1572 }),
  .B({ S1593 }),
  .Y({ S1595 })
);
NAND #() 
NAND_860_ (
  .A({ S1582 }),
  .B({ S1594 }),
  .Y({ S1596 })
);
NOR #() 
NOR_381_ (
  .A({ S1549 }),
  .B({ S1595 }),
  .Y({ S1597 })
);
NAND #() 
NAND_861_ (
  .A({ S1550 }),
  .B({ S1596 }),
  .Y({ S1598 })
);
NOR #() 
NOR_382_ (
  .A({ S8468 }),
  .B({ S1387 }),
  .Y({ S1599 })
);
NAND #() 
NAND_862_ (
  .A({ S8457 }),
  .B({ S1386 }),
  .Y({ S1600 })
);
NOR #() 
NOR_383_ (
  .A({ S8426 }),
  .B({ S387 }),
  .Y({ S1601 })
);
NOR #() 
NOR_384_ (
  .A({ S387 }),
  .B({ S1398 }),
  .Y({ S1602 })
);
NAND #() 
NAND_863_ (
  .A({ S8375 }),
  .B({ S1601 }),
  .Y({ S1603 })
);
NOR #() 
NOR_385_ (
  .A({ S1599 }),
  .B({ S1602 }),
  .Y({ S1604 })
);
NAND #() 
NAND_864_ (
  .A({ S1600 }),
  .B({ S1603 }),
  .Y({ S1605 })
);
NAND #() 
NAND_865_ (
  .A({ S1597 }),
  .B({ S1605 }),
  .Y({ S1606 })
);
NOR #() 
NOR_386_ (
  .A({ S8385 }),
  .B({ S8545 }),
  .Y({ S1607 })
);
NAND #() 
NAND_866_ (
  .A({ controller_fib_4 }),
  .B({ S1607 }),
  .Y({ S1608 })
);
NAND #() 
NAND_867_ (
  .A({ S1606 }),
  .B({ S1608 }),
  .Y({ S1609 })
);
NAND #() 
NAND_868_ (
  .A({ controller_216_B_0 }),
  .B({ S1607 }),
  .Y({ S1610 })
);
NAND #() 
NAND_869_ (
  .A({ S1603 }),
  .B({ S1610 }),
  .Y({ S1611 })
);
NOT #() 
NOT_192_ (
  .A({ S1611 }),
  .Y({ S1612 })
);
NOR #() 
NOR_387_ (
  .A({ S1605 }),
  .B({ S1607 }),
  .Y({ S1613 })
);
NOR #() 
NOR_388_ (
  .A({ S1609 }),
  .B({ S1613 }),
  .Y({ S1614 })
);
NAND #() 
NAND_870_ (
  .A({ datapath_shiftunit_2135_A }),
  .B({ S1614 }),
  .Y({ S1615 })
);
NAND #() 
NAND_871_ (
  .A({ datapath_shiftunit_2439_A }),
  .B({ S1609 }),
  .Y({ S1616 })
);
NAND #() 
NAND_872_ (
  .A({ datapath_multdivunit_outmdu2_0 }),
  .B({ S8570 }),
  .Y({ S1617 })
);
NOR #() 
NOR_389_ (
  .A({ controller_216_B_0 }),
  .B({ controller_opcode_2 }),
  .Y({ S1618 })
);
NOT #() 
NOT_193_ (
  .A({ S1618 }),
  .Y({ S1619 })
);
NOR #() 
NOR_390_ (
  .A({ S8309 }),
  .B({ S1618 }),
  .Y({ S1620 })
);
NAND #() 
NAND_873_ (
  .A({ controller_opcode_3 }),
  .B({ S1619 }),
  .Y({ S1621 })
);
NOR #() 
NOR_391_ (
  .A({ S369 }),
  .B({ S1621 }),
  .Y({ S1622 })
);
NAND #() 
NAND_874_ (
  .A({ S368 }),
  .B({ S1620 }),
  .Y({ S1623 })
);
NAND #() 
NAND_875_ (
  .A({ S7884 }),
  .B({ S1622 }),
  .Y({ S1624 })
);
NAND #() 
NAND_876_ (
  .A({ S1617 }),
  .B({ S1624 }),
  .Y({ S1625 })
);
NAND #() 
NAND_877_ (
  .A({ datapath_multdivunit_outmdu1_0 }),
  .B({ S1377 }),
  .Y({ S1626 })
);
NOR #() 
NOR_392_ (
  .A({ controller_opcode_2 }),
  .B({ S8577 }),
  .Y({ S1627 })
);
NAND #() 
NAND_878_ (
  .A({ S8299 }),
  .B({ S8576 }),
  .Y({ S1628 })
);
NAND #() 
NAND_879_ (
  .A({ datapath_databusin_0 }),
  .B({ S1627 }),
  .Y({ S1629 })
);
NAND #() 
NAND_880_ (
  .A({ S1626 }),
  .B({ S1629 }),
  .Y({ S1630 })
);
NOR #() 
NOR_393_ (
  .A({ S1625 }),
  .B({ S1630 }),
  .Y({ S1631 })
);
NAND #() 
NAND_881_ (
  .A({ S1616 }),
  .B({ S1631 }),
  .Y({ S1632 })
);
NOT #() 
NOT_194_ (
  .A({ S1632 }),
  .Y({ S1633 })
);
NAND #() 
NAND_882_ (
  .A({ S1615 }),
  .B({ S1633 }),
  .Y({ S1634 })
);
NOR #() 
NOR_394_ (
  .A({ S1548 }),
  .B({ S1634 }),
  .Y({ S1635 })
);
NAND #() 
NAND_883_ (
  .A({ S1536 }),
  .B({ S1635 }),
  .Y({ S1636 })
);
NOR #() 
NOR_395_ (
  .A({ S1530 }),
  .B({ S1636 }),
  .Y({ S1637 })
);
NAND #() 
NAND_884_ (
  .A({ S1545 }),
  .B({ S1637 }),
  .Y({ datapath_indatatrf_0 })
);
NAND #() 
NAND_885_ (
  .A({ S8375 }),
  .B({ S8520 }),
  .Y({ S1638 })
);
NAND #() 
NAND_886_ (
  .A({ S1537 }),
  .B({ S1638 }),
  .Y({ S1639 })
);
NOR #() 
NOR_396_ (
  .A({ S1622 }),
  .B({ S1639 }),
  .Y({ S1640 })
);
NOR #() 
NOR_397_ (
  .A({ S1377 }),
  .B({ S1627 }),
  .Y({ S1641 })
);
NAND #() 
NAND_887_ (
  .A({ S1640 }),
  .B({ S1641 }),
  .Y({ S1642 })
);
NOT #() 
NOT_195_ (
  .A({ S1642 }),
  .Y({ S1643 })
);
NAND #() 
NAND_888_ (
  .A({ datapath_instruction_0 }),
  .B({ datapath_instruction_1 }),
  .Y({ S1644 })
);
NOT #() 
NOT_196_ (
  .A({ S1644 }),
  .Y({ S1645 })
);
NAND #() 
NAND_889_ (
  .A({ datapath_instruction_2 }),
  .B({ S1645 }),
  .Y({ S1646 })
);
NAND #() 
NAND_890_ (
  .A({ S8570 }),
  .B({ S1646 }),
  .Y({ S1647 })
);
NOT #() 
NOT_197_ (
  .A({ S1647 }),
  .Y({ S1648 })
);
NOR #() 
NOR_398_ (
  .A({ S1642 }),
  .B({ S1648 }),
  .Y({ S1649 })
);
NAND #() 
NAND_891_ (
  .A({ S1643 }),
  .B({ S1647 }),
  .Y({ S1650 })
);
NOR #() 
NOR_399_ (
  .A({ S8571 }),
  .B({ S1644 }),
  .Y({ S1651 })
);
NOR #() 
NOR_400_ (
  .A({ datapath_instruction_2 }),
  .B({ S1651 }),
  .Y({ S1652 })
);
NOT #() 
NOT_198_ (
  .A({ S1652 }),
  .Y({ S1653 })
);
NOR #() 
NOR_401_ (
  .A({ S1649 }),
  .B({ S1652 }),
  .Y({ S1654 })
);
NAND #() 
NAND_892_ (
  .A({ S1650 }),
  .B({ S1653 }),
  .Y({ S1655 })
);
NOR #() 
NOR_402_ (
  .A({ S8571 }),
  .B({ S1646 }),
  .Y({ S1656 })
);
NOR #() 
NOR_403_ (
  .A({ datapath_instruction_3 }),
  .B({ S1656 }),
  .Y({ S1657 })
);
NOT #() 
NOT_199_ (
  .A({ S1657 }),
  .Y({ S1658 })
);
NOR #() 
NOR_404_ (
  .A({ S8204 }),
  .B({ S1650 }),
  .Y({ S1659 })
);
NAND #() 
NAND_893_ (
  .A({ datapath_instruction_3 }),
  .B({ S1649 }),
  .Y({ S1660 })
);
NOR #() 
NOR_405_ (
  .A({ S1657 }),
  .B({ S1659 }),
  .Y({ S1661 })
);
NAND #() 
NAND_894_ (
  .A({ S1658 }),
  .B({ S1660 }),
  .Y({ S1662 })
);
NOR #() 
NOR_406_ (
  .A({ S1654 }),
  .B({ S1662 }),
  .Y({ S1663 })
);
NAND #() 
NAND_895_ (
  .A({ S1655 }),
  .B({ S1661 }),
  .Y({ S1664 })
);
NOR #() 
NOR_407_ (
  .A({ datapath_instruction_0 }),
  .B({ datapath_instruction_1 }),
  .Y({ S1665 })
);
NOT #() 
NOT_200_ (
  .A({ S1665 }),
  .Y({ S1666 })
);
NAND #() 
NAND_896_ (
  .A({ datapath_instruction_1 }),
  .B({ S1642 }),
  .Y({ S1667 })
);
NAND #() 
NAND_897_ (
  .A({ S8570 }),
  .B({ S1644 }),
  .Y({ S1668 })
);
NAND #() 
NAND_898_ (
  .A({ S1667 }),
  .B({ S1668 }),
  .Y({ S1669 })
);
NOT #() 
NOT_201_ (
  .A({ S1669 }),
  .Y({ S1670 })
);
NOR #() 
NOR_408_ (
  .A({ S1665 }),
  .B({ S1670 }),
  .Y({ S1671 })
);
NAND #() 
NAND_899_ (
  .A({ S1666 }),
  .B({ S1669 }),
  .Y({ S1672 })
);
NOR #() 
NOR_409_ (
  .A({ S1664 }),
  .B({ S1672 }),
  .Y({ S1673 })
);
NAND #() 
NAND_900_ (
  .A({ S1663 }),
  .B({ S1671 }),
  .Y({ S1674 })
);
NOR #() 
NOR_410_ (
  .A({ S8572 }),
  .B({ S1628 }),
  .Y({ S1675 })
);
NOR #() 
NOR_411_ (
  .A({ S8568 }),
  .B({ S1675 }),
  .Y({ S1676 })
);
NAND #() 
NAND_901_ (
  .A({ S8569 }),
  .B({ S1640 }),
  .Y({ S1677 })
);
NOR #() 
NOR_412_ (
  .A({ S1675 }),
  .B({ S1677 }),
  .Y({ S1678 })
);
NAND #() 
NAND_902_ (
  .A({ S1640 }),
  .B({ S1676 }),
  .Y({ S1679 })
);
NAND #() 
NAND_903_ (
  .A({ datapath_instruction_0 }),
  .B({ S1642 }),
  .Y({ S1680 })
);
NOT #() 
NOT_202_ (
  .A({ S1680 }),
  .Y({ S1681 })
);
NOR #() 
NOR_413_ (
  .A({ datapath_instruction_0 }),
  .B({ S8571 }),
  .Y({ S1682 })
);
NOT #() 
NOT_203_ (
  .A({ S1682 }),
  .Y({ S1683 })
);
NOR #() 
NOR_414_ (
  .A({ S1681 }),
  .B({ S1682 }),
  .Y({ S1684 })
);
NAND #() 
NAND_904_ (
  .A({ S1680 }),
  .B({ S1683 }),
  .Y({ S1685 })
);
NOR #() 
NOR_415_ (
  .A({ S1678 }),
  .B({ S1684 }),
  .Y({ S1686 })
);
NAND #() 
NAND_905_ (
  .A({ S1679 }),
  .B({ S1685 }),
  .Y({ S1687 })
);
NOR #() 
NOR_416_ (
  .A({ S1674 }),
  .B({ S1687 }),
  .Y({ S1688 })
);
NAND #() 
NAND_906_ (
  .A({ S1673 }),
  .B({ S1686 }),
  .Y({ S1689 })
);
NAND #() 
NAND_907_ (
  .A({ datapath_indatatrf_0 }),
  .B({ S1688 }),
  .Y({ S1690 })
);
NAND #() 
NAND_908_ (
  .A({ datapath_theregisterfile_memtrf_64 }),
  .B({ S1689 }),
  .Y({ S1691 })
);
NAND #() 
NAND_909_ (
  .A({ S1690 }),
  .B({ S1691 }),
  .Y({ S4 })
);
NOR #() 
NOR_417_ (
  .A({ S1168 }),
  .B({ S1389 }),
  .Y({ S1692 })
);
NAND #() 
NAND_910_ (
  .A({ controller_fib_1 }),
  .B({ S1409 }),
  .Y({ S1693 })
);
NOT #() 
NOT_204_ (
  .A({ S1693 }),
  .Y({ S1694 })
);
NOR #() 
NOR_418_ (
  .A({ S1692 }),
  .B({ S1694 }),
  .Y({ S1695 })
);
NOR #() 
NOR_419_ (
  .A({ S1416 }),
  .B({ S1695 }),
  .Y({ S1696 })
);
NOR #() 
NOR_420_ (
  .A({ controller_outflag_1 }),
  .B({ S1462 }),
  .Y({ S1697 })
);
NOT #() 
NOT_205_ (
  .A({ S1697 }),
  .Y({ S1698 })
);
NAND #() 
NAND_911_ (
  .A({ datapath_theregisterfile_memtrf_241 }),
  .B({ S1437 }),
  .Y({ S1699 })
);
NAND #() 
NAND_912_ (
  .A({ datapath_theregisterfile_memtrf_177 }),
  .B({ S1438 }),
  .Y({ S1700 })
);
NAND #() 
NAND_913_ (
  .A({ S1699 }),
  .B({ S1700 }),
  .Y({ S1701 })
);
NAND #() 
NAND_914_ (
  .A({ S1457 }),
  .B({ S1701 }),
  .Y({ S1702 })
);
NAND #() 
NAND_915_ (
  .A({ S7794 }),
  .B({ S1437 }),
  .Y({ S1703 })
);
NOR #() 
NOR_421_ (
  .A({ datapath_theregisterfile_memtrf_161 }),
  .B({ S1437 }),
  .Y({ S1704 })
);
NAND #() 
NAND_916_ (
  .A({ S1458 }),
  .B({ S1703 }),
  .Y({ S1705 })
);
NOR #() 
NOR_422_ (
  .A({ S1704 }),
  .B({ S1705 }),
  .Y({ S1706 })
);
NAND #() 
NAND_917_ (
  .A({ datapath_theregisterfile_memtrf_145 }),
  .B({ S1438 }),
  .Y({ S1707 })
);
NAND #() 
NAND_918_ (
  .A({ datapath_theregisterfile_memtrf_209 }),
  .B({ S1437 }),
  .Y({ S1708 })
);
NAND #() 
NAND_919_ (
  .A({ S1707 }),
  .B({ S1708 }),
  .Y({ S1709 })
);
NAND #() 
NAND_920_ (
  .A({ S1457 }),
  .B({ S1709 }),
  .Y({ S1710 })
);
NOR #() 
NOR_423_ (
  .A({ datapath_theregisterfile_memtrf_129 }),
  .B({ S1437 }),
  .Y({ S1711 })
);
NOR #() 
NOR_424_ (
  .A({ datapath_theregisterfile_memtrf_193 }),
  .B({ S1438 }),
  .Y({ S1712 })
);
NOR #() 
NOR_425_ (
  .A({ S1711 }),
  .B({ S1712 }),
  .Y({ S1713 })
);
NAND #() 
NAND_921_ (
  .A({ S1458 }),
  .B({ S1713 }),
  .Y({ S1714 })
);
NAND #() 
NAND_922_ (
  .A({ S1710 }),
  .B({ S1714 }),
  .Y({ S1715 })
);
NOR #() 
NOR_426_ (
  .A({ S1443 }),
  .B({ S1715 }),
  .Y({ S1716 })
);
NOR #() 
NOR_427_ (
  .A({ S1444 }),
  .B({ S1706 }),
  .Y({ S1717 })
);
NAND #() 
NAND_923_ (
  .A({ S1702 }),
  .B({ S1717 }),
  .Y({ S1718 })
);
NAND #() 
NAND_924_ (
  .A({ S1449 }),
  .B({ S1718 }),
  .Y({ S1719 })
);
NOR #() 
NOR_428_ (
  .A({ S1716 }),
  .B({ S1719 }),
  .Y({ S1720 })
);
NAND #() 
NAND_925_ (
  .A({ datapath_theregisterfile_memtrf_97 }),
  .B({ S1458 }),
  .Y({ S1721 })
);
NAND #() 
NAND_926_ (
  .A({ datapath_theregisterfile_memtrf_113 }),
  .B({ S1457 }),
  .Y({ S1722 })
);
NAND #() 
NAND_927_ (
  .A({ S1721 }),
  .B({ S1722 }),
  .Y({ S1723 })
);
NAND #() 
NAND_928_ (
  .A({ S1437 }),
  .B({ S1723 }),
  .Y({ S1724 })
);
NAND #() 
NAND_929_ (
  .A({ datapath_theregisterfile_memtrf_33 }),
  .B({ S1458 }),
  .Y({ S1725 })
);
NAND #() 
NAND_930_ (
  .A({ datapath_theregisterfile_memtrf_49 }),
  .B({ S1457 }),
  .Y({ S1726 })
);
NAND #() 
NAND_931_ (
  .A({ S1725 }),
  .B({ S1726 }),
  .Y({ S1727 })
);
NAND #() 
NAND_932_ (
  .A({ S1438 }),
  .B({ S1727 }),
  .Y({ S1728 })
);
NAND #() 
NAND_933_ (
  .A({ S1724 }),
  .B({ S1728 }),
  .Y({ S1729 })
);
NAND #() 
NAND_934_ (
  .A({ S1487 }),
  .B({ S1729 }),
  .Y({ S1730 })
);
NAND #() 
NAND_935_ (
  .A({ datapath_theregisterfile_memtrf_81 }),
  .B({ S1498 }),
  .Y({ S1731 })
);
NOR #() 
NOR_429_ (
  .A({ datapath_theregisterfile_memtrf_65 }),
  .B({ S1438 }),
  .Y({ S1732 })
);
NOT #() 
NOT_206_ (
  .A({ S1732 }),
  .Y({ S1733 })
);
NAND #() 
NAND_936_ (
  .A({ datapath_theregisterfile_memtrf_17 }),
  .B({ S1438 }),
  .Y({ S1734 })
);
NAND #() 
NAND_937_ (
  .A({ S1457 }),
  .B({ S1734 }),
  .Y({ S1735 })
);
NAND #() 
NAND_938_ (
  .A({ S1733 }),
  .B({ S1735 }),
  .Y({ S1736 })
);
NAND #() 
NAND_939_ (
  .A({ S1731 }),
  .B({ S1736 }),
  .Y({ S1737 })
);
NOT #() 
NOT_207_ (
  .A({ S1737 }),
  .Y({ S1738 })
);
NOR #() 
NOR_430_ (
  .A({ S1452 }),
  .B({ S1738 }),
  .Y({ S1739 })
);
NAND #() 
NAND_940_ (
  .A({ S1451 }),
  .B({ S1737 }),
  .Y({ S1740 })
);
NAND #() 
NAND_941_ (
  .A({ S1730 }),
  .B({ S1740 }),
  .Y({ S1741 })
);
NOR #() 
NOR_431_ (
  .A({ S1720 }),
  .B({ S1739 }),
  .Y({ S1742 })
);
NOR #() 
NOR_432_ (
  .A({ S1720 }),
  .B({ S1741 }),
  .Y({ S1743 })
);
NAND #() 
NAND_942_ (
  .A({ S1730 }),
  .B({ S1742 }),
  .Y({ S1744 })
);
NOR #() 
NOR_433_ (
  .A({ S1697 }),
  .B({ S1743 }),
  .Y({ S1745 })
);
NAND #() 
NAND_943_ (
  .A({ S1698 }),
  .B({ S1744 }),
  .Y({ S1746 })
);
NOR #() 
NOR_434_ (
  .A({ S1430 }),
  .B({ S1746 }),
  .Y({ S1747 })
);
NOR #() 
NOR_435_ (
  .A({ S1696 }),
  .B({ S1747 }),
  .Y({ S1748 })
);
NOT #() 
NOT_208_ (
  .A({ S1748 }),
  .Y({ S1749 })
);
NOR #() 
NOR_436_ (
  .A({ S1168 }),
  .B({ S1749 }),
  .Y({ S1750 })
);
NAND #() 
NAND_944_ (
  .A({ datapath_addsubunit_in1_1 }),
  .B({ S1748 }),
  .Y({ S1751 })
);
NAND #() 
NAND_945_ (
  .A({ S1168 }),
  .B({ S1749 }),
  .Y({ S1752 })
);
NOT #() 
NOT_209_ (
  .A({ S1752 }),
  .Y({ S1753 })
);
NOR #() 
NOR_437_ (
  .A({ S1750 }),
  .B({ S1753 }),
  .Y({ S1754 })
);
NOT #() 
NOT_210_ (
  .A({ S1754 }),
  .Y({ S1755 })
);
NAND #() 
NAND_946_ (
  .A({ S1520 }),
  .B({ S1755 }),
  .Y({ S1756 })
);
NOR #() 
NOR_438_ (
  .A({ S1520 }),
  .B({ S1755 }),
  .Y({ S1757 })
);
NOR #() 
NOR_439_ (
  .A({ S1526 }),
  .B({ S1757 }),
  .Y({ S1758 })
);
NAND #() 
NAND_947_ (
  .A({ S1756 }),
  .B({ S1758 }),
  .Y({ S1759 })
);
NOR #() 
NOR_440_ (
  .A({ S1531 }),
  .B({ S1754 }),
  .Y({ S1760 })
);
NOT #() 
NOT_211_ (
  .A({ S1760 }),
  .Y({ S1761 })
);
NAND #() 
NAND_948_ (
  .A({ S1531 }),
  .B({ S1754 }),
  .Y({ S1762 })
);
NAND #() 
NAND_949_ (
  .A({ S1527 }),
  .B({ S1762 }),
  .Y({ S1763 })
);
NOR #() 
NOR_441_ (
  .A({ S1760 }),
  .B({ S1763 }),
  .Y({ S1764 })
);
NOR #() 
NOR_442_ (
  .A({ datapath_addsubunit_in1_1 }),
  .B({ S1541 }),
  .Y({ S1765 })
);
NOT #() 
NOT_212_ (
  .A({ S1765 }),
  .Y({ S1766 })
);
NOR #() 
NOR_443_ (
  .A({ datapath_addsubunit_in1_1 }),
  .B({ S1539 }),
  .Y({ S1767 })
);
NOR #() 
NOR_444_ (
  .A({ S1542 }),
  .B({ S1767 }),
  .Y({ S1768 })
);
NOR #() 
NOR_445_ (
  .A({ S1765 }),
  .B({ S1768 }),
  .Y({ S1769 })
);
NOR #() 
NOR_446_ (
  .A({ S1547 }),
  .B({ S1695 }),
  .Y({ S1770 })
);
NAND #() 
NAND_950_ (
  .A({ datapath_shiftunit_2153_A }),
  .B({ S1614 }),
  .Y({ S1771 })
);
NOR #() 
NOR_447_ (
  .A({ datapath_muxmem_in2_0 }),
  .B({ datapath_muxmem_in2_1 }),
  .Y({ S1772 })
);
NOR #() 
NOR_448_ (
  .A({ S1335 }),
  .B({ S1772 }),
  .Y({ S1773 })
);
NOT #() 
NOT_213_ (
  .A({ S1773 }),
  .Y({ S1774 })
);
NAND #() 
NAND_951_ (
  .A({ S1622 }),
  .B({ S1773 }),
  .Y({ S1775 })
);
NAND #() 
NAND_952_ (
  .A({ datapath_multdivunit_outmdu2_1 }),
  .B({ S8570 }),
  .Y({ S1776 })
);
NAND #() 
NAND_953_ (
  .A({ S1775 }),
  .B({ S1776 }),
  .Y({ S1777 })
);
NAND #() 
NAND_954_ (
  .A({ datapath_multdivunit_outmdu1_1 }),
  .B({ S1377 }),
  .Y({ S1778 })
);
NAND #() 
NAND_955_ (
  .A({ datapath_databusin_1 }),
  .B({ S1627 }),
  .Y({ S1779 })
);
NAND #() 
NAND_956_ (
  .A({ S1778 }),
  .B({ S1779 }),
  .Y({ S1780 })
);
NOR #() 
NOR_449_ (
  .A({ S1777 }),
  .B({ S1780 }),
  .Y({ S1781 })
);
NAND #() 
NAND_957_ (
  .A({ datapath_shiftunit_2457_A }),
  .B({ S1609 }),
  .Y({ S1782 })
);
NAND #() 
NAND_958_ (
  .A({ S1771 }),
  .B({ S1781 }),
  .Y({ S1783 })
);
NOR #() 
NOR_450_ (
  .A({ S1770 }),
  .B({ S1783 }),
  .Y({ S1784 })
);
NAND #() 
NAND_959_ (
  .A({ S1782 }),
  .B({ S1784 }),
  .Y({ S1785 })
);
NOR #() 
NOR_451_ (
  .A({ S1769 }),
  .B({ S1785 }),
  .Y({ S1786 })
);
NOR #() 
NOR_452_ (
  .A({ S1168 }),
  .B({ S1748 }),
  .Y({ S1787 })
);
NOT #() 
NOT_214_ (
  .A({ S1787 }),
  .Y({ S1788 })
);
NAND #() 
NAND_960_ (
  .A({ S1534 }),
  .B({ S1787 }),
  .Y({ S1789 })
);
NAND #() 
NAND_961_ (
  .A({ S1786 }),
  .B({ S1789 }),
  .Y({ S1790 })
);
NOR #() 
NOR_453_ (
  .A({ S1764 }),
  .B({ S1790 }),
  .Y({ S1791 })
);
NAND #() 
NAND_962_ (
  .A({ S1759 }),
  .B({ S1791 }),
  .Y({ datapath_indatatrf_1 })
);
NAND #() 
NAND_963_ (
  .A({ datapath_indatatrf_1 }),
  .B({ S1688 }),
  .Y({ S1792 })
);
NAND #() 
NAND_964_ (
  .A({ datapath_theregisterfile_memtrf_65 }),
  .B({ S1689 }),
  .Y({ S1793 })
);
NAND #() 
NAND_965_ (
  .A({ S1792 }),
  .B({ S1793 }),
  .Y({ S5 })
);
NOR #() 
NOR_454_ (
  .A({ S1116 }),
  .B({ S1389 }),
  .Y({ S1794 })
);
NAND #() 
NAND_966_ (
  .A({ controller_fib_2 }),
  .B({ S1409 }),
  .Y({ S1795 })
);
NOT #() 
NOT_215_ (
  .A({ S1795 }),
  .Y({ S1796 })
);
NOR #() 
NOR_455_ (
  .A({ S1794 }),
  .B({ S1796 }),
  .Y({ S1797 })
);
NOT #() 
NOT_216_ (
  .A({ S1797 }),
  .Y({ S1798 })
);
NAND #() 
NAND_967_ (
  .A({ S1417 }),
  .B({ S1798 }),
  .Y({ S1799 })
);
NOR #() 
NOR_456_ (
  .A({ controller_outflag_2 }),
  .B({ S1462 }),
  .Y({ S1800 })
);
NOT #() 
NOT_217_ (
  .A({ S1800 }),
  .Y({ S1801 })
);
NAND #() 
NAND_968_ (
  .A({ datapath_theregisterfile_memtrf_242 }),
  .B({ S1437 }),
  .Y({ S1802 })
);
NAND #() 
NAND_969_ (
  .A({ datapath_theregisterfile_memtrf_178 }),
  .B({ S1438 }),
  .Y({ S1803 })
);
NAND #() 
NAND_970_ (
  .A({ S1802 }),
  .B({ S1803 }),
  .Y({ S1804 })
);
NAND #() 
NAND_971_ (
  .A({ S1457 }),
  .B({ S1804 }),
  .Y({ S1805 })
);
NAND #() 
NAND_972_ (
  .A({ S7805 }),
  .B({ S1437 }),
  .Y({ S1806 })
);
NOR #() 
NOR_457_ (
  .A({ datapath_theregisterfile_memtrf_162 }),
  .B({ S1437 }),
  .Y({ S1807 })
);
NAND #() 
NAND_973_ (
  .A({ S1458 }),
  .B({ S1806 }),
  .Y({ S1808 })
);
NOR #() 
NOR_458_ (
  .A({ S1807 }),
  .B({ S1808 }),
  .Y({ S1809 })
);
NAND #() 
NAND_974_ (
  .A({ datapath_theregisterfile_memtrf_146 }),
  .B({ S1438 }),
  .Y({ S1810 })
);
NAND #() 
NAND_975_ (
  .A({ datapath_theregisterfile_memtrf_210 }),
  .B({ S1437 }),
  .Y({ S1811 })
);
NAND #() 
NAND_976_ (
  .A({ S1810 }),
  .B({ S1811 }),
  .Y({ S1812 })
);
NAND #() 
NAND_977_ (
  .A({ S1457 }),
  .B({ S1812 }),
  .Y({ S1813 })
);
NOR #() 
NOR_459_ (
  .A({ datapath_theregisterfile_memtrf_130 }),
  .B({ S1437 }),
  .Y({ S1814 })
);
NOR #() 
NOR_460_ (
  .A({ datapath_theregisterfile_memtrf_194 }),
  .B({ S1438 }),
  .Y({ S1815 })
);
NOR #() 
NOR_461_ (
  .A({ S1814 }),
  .B({ S1815 }),
  .Y({ S1816 })
);
NAND #() 
NAND_978_ (
  .A({ S1458 }),
  .B({ S1816 }),
  .Y({ S1817 })
);
NAND #() 
NAND_979_ (
  .A({ S1813 }),
  .B({ S1817 }),
  .Y({ S1818 })
);
NOR #() 
NOR_462_ (
  .A({ S1443 }),
  .B({ S1818 }),
  .Y({ S1819 })
);
NOR #() 
NOR_463_ (
  .A({ S1444 }),
  .B({ S1809 }),
  .Y({ S1820 })
);
NAND #() 
NAND_980_ (
  .A({ S1805 }),
  .B({ S1820 }),
  .Y({ S1821 })
);
NAND #() 
NAND_981_ (
  .A({ S1449 }),
  .B({ S1821 }),
  .Y({ S1822 })
);
NOR #() 
NOR_464_ (
  .A({ S1819 }),
  .B({ S1822 }),
  .Y({ S1823 })
);
NAND #() 
NAND_982_ (
  .A({ datapath_theregisterfile_memtrf_98 }),
  .B({ S1458 }),
  .Y({ S1824 })
);
NAND #() 
NAND_983_ (
  .A({ datapath_theregisterfile_memtrf_114 }),
  .B({ S1457 }),
  .Y({ S1825 })
);
NAND #() 
NAND_984_ (
  .A({ S1824 }),
  .B({ S1825 }),
  .Y({ S1826 })
);
NAND #() 
NAND_985_ (
  .A({ S1437 }),
  .B({ S1826 }),
  .Y({ S1827 })
);
NAND #() 
NAND_986_ (
  .A({ datapath_theregisterfile_memtrf_34 }),
  .B({ S1458 }),
  .Y({ S1828 })
);
NAND #() 
NAND_987_ (
  .A({ datapath_theregisterfile_memtrf_50 }),
  .B({ S1457 }),
  .Y({ S1829 })
);
NAND #() 
NAND_988_ (
  .A({ S1828 }),
  .B({ S1829 }),
  .Y({ S1830 })
);
NAND #() 
NAND_989_ (
  .A({ S1438 }),
  .B({ S1830 }),
  .Y({ S1831 })
);
NAND #() 
NAND_990_ (
  .A({ S1827 }),
  .B({ S1831 }),
  .Y({ S1832 })
);
NAND #() 
NAND_991_ (
  .A({ S1487 }),
  .B({ S1832 }),
  .Y({ S1833 })
);
NAND #() 
NAND_992_ (
  .A({ datapath_theregisterfile_memtrf_82 }),
  .B({ S1498 }),
  .Y({ S1834 })
);
NOR #() 
NOR_465_ (
  .A({ datapath_theregisterfile_memtrf_66 }),
  .B({ S1438 }),
  .Y({ S1835 })
);
NOT #() 
NOT_218_ (
  .A({ S1835 }),
  .Y({ S1836 })
);
NAND #() 
NAND_993_ (
  .A({ datapath_theregisterfile_memtrf_18 }),
  .B({ S1438 }),
  .Y({ S1837 })
);
NAND #() 
NAND_994_ (
  .A({ S1457 }),
  .B({ S1837 }),
  .Y({ S1838 })
);
NAND #() 
NAND_995_ (
  .A({ S1836 }),
  .B({ S1838 }),
  .Y({ S1839 })
);
NAND #() 
NAND_996_ (
  .A({ S1834 }),
  .B({ S1839 }),
  .Y({ S1840 })
);
NOT #() 
NOT_219_ (
  .A({ S1840 }),
  .Y({ S1841 })
);
NOR #() 
NOR_466_ (
  .A({ S1452 }),
  .B({ S1841 }),
  .Y({ S1842 })
);
NAND #() 
NAND_997_ (
  .A({ S1451 }),
  .B({ S1840 }),
  .Y({ S1843 })
);
NAND #() 
NAND_998_ (
  .A({ S1833 }),
  .B({ S1843 }),
  .Y({ S1844 })
);
NOR #() 
NOR_467_ (
  .A({ S1823 }),
  .B({ S1842 }),
  .Y({ S1845 })
);
NOR #() 
NOR_468_ (
  .A({ S1823 }),
  .B({ S1844 }),
  .Y({ S1846 })
);
NAND #() 
NAND_999_ (
  .A({ S1833 }),
  .B({ S1845 }),
  .Y({ S1847 })
);
NOR #() 
NOR_469_ (
  .A({ S1800 }),
  .B({ S1846 }),
  .Y({ S1848 })
);
NAND #() 
NAND_1000_ (
  .A({ S1801 }),
  .B({ S1847 }),
  .Y({ S1849 })
);
NAND #() 
NAND_1001_ (
  .A({ S1429 }),
  .B({ S1848 }),
  .Y({ S1850 })
);
NAND #() 
NAND_1002_ (
  .A({ S1799 }),
  .B({ S1850 }),
  .Y({ S1851 })
);
NOT #() 
NOT_220_ (
  .A({ S1851 }),
  .Y({ S1852 })
);
NOR #() 
NOR_470_ (
  .A({ datapath_addsubunit_in1_2 }),
  .B({ S1852 }),
  .Y({ S1853 })
);
NOT #() 
NOT_221_ (
  .A({ S1853 }),
  .Y({ S1854 })
);
NOR #() 
NOR_471_ (
  .A({ S1116 }),
  .B({ S1851 }),
  .Y({ S1855 })
);
NOT #() 
NOT_222_ (
  .A({ S1855 }),
  .Y({ S1856 })
);
NAND #() 
NAND_1003_ (
  .A({ S1854 }),
  .B({ S1856 }),
  .Y({ S1857 })
);
NOR #() 
NOR_472_ (
  .A({ S1750 }),
  .B({ S1757 }),
  .Y({ S1858 })
);
NOR #() 
NOR_473_ (
  .A({ S1857 }),
  .B({ S1858 }),
  .Y({ S1859 })
);
NAND #() 
NAND_1004_ (
  .A({ S1857 }),
  .B({ S1858 }),
  .Y({ S1860 })
);
NOT #() 
NOT_223_ (
  .A({ S1860 }),
  .Y({ S1861 })
);
NOR #() 
NOR_474_ (
  .A({ S1859 }),
  .B({ S1861 }),
  .Y({ S1862 })
);
NAND #() 
NAND_1005_ (
  .A({ S1525 }),
  .B({ S1862 }),
  .Y({ S1863 })
);
NAND #() 
NAND_1006_ (
  .A({ S1761 }),
  .B({ S1788 }),
  .Y({ S1864 })
);
NOR #() 
NOR_475_ (
  .A({ S1857 }),
  .B({ S1864 }),
  .Y({ S1865 })
);
NAND #() 
NAND_1007_ (
  .A({ S1857 }),
  .B({ S1864 }),
  .Y({ S1866 })
);
NAND #() 
NAND_1008_ (
  .A({ S1527 }),
  .B({ S1866 }),
  .Y({ S1867 })
);
NOR #() 
NOR_476_ (
  .A({ S1865 }),
  .B({ S1867 }),
  .Y({ S1868 })
);
NAND #() 
NAND_1009_ (
  .A({ datapath_addsubunit_in1_2 }),
  .B({ S1851 }),
  .Y({ S1869 })
);
NOR #() 
NOR_477_ (
  .A({ S1533 }),
  .B({ S1869 }),
  .Y({ S1870 })
);
NOR #() 
NOR_478_ (
  .A({ S1547 }),
  .B({ S1797 }),
  .Y({ S1871 })
);
NAND #() 
NAND_1010_ (
  .A({ datapath_shiftunit_2171_A }),
  .B({ S1614 }),
  .Y({ S1872 })
);
NAND #() 
NAND_1011_ (
  .A({ datapath_shiftunit_2475_A }),
  .B({ S1609 }),
  .Y({ S1873 })
);
NAND #() 
NAND_1012_ (
  .A({ S7897 }),
  .B({ S1336 }),
  .Y({ S1874 })
);
NAND #() 
NAND_1013_ (
  .A({ S1338 }),
  .B({ S1874 }),
  .Y({ S1875 })
);
NOR #() 
NOR_479_ (
  .A({ S1623 }),
  .B({ S1875 }),
  .Y({ S1876 })
);
NOR #() 
NOR_480_ (
  .A({ S8054 }),
  .B({ S8571 }),
  .Y({ S1877 })
);
NOR #() 
NOR_481_ (
  .A({ S8011 }),
  .B({ S1378 }),
  .Y({ S1878 })
);
NAND #() 
NAND_1014_ (
  .A({ datapath_databusin_2 }),
  .B({ S1627 }),
  .Y({ S1879 })
);
NOR #() 
NOR_482_ (
  .A({ S1876 }),
  .B({ S1878 }),
  .Y({ S1880 })
);
NAND #() 
NAND_1015_ (
  .A({ S1879 }),
  .B({ S1880 }),
  .Y({ S1881 })
);
NOR #() 
NOR_483_ (
  .A({ S1877 }),
  .B({ S1881 }),
  .Y({ S1882 })
);
NAND #() 
NAND_1016_ (
  .A({ S1873 }),
  .B({ S1882 }),
  .Y({ S1883 })
);
NOR #() 
NOR_484_ (
  .A({ S1871 }),
  .B({ S1883 }),
  .Y({ S1884 })
);
NAND #() 
NAND_1017_ (
  .A({ S1872 }),
  .B({ S1884 }),
  .Y({ S1885 })
);
NOR #() 
NOR_485_ (
  .A({ S1116 }),
  .B({ S1765 }),
  .Y({ S1886 })
);
NOR #() 
NOR_486_ (
  .A({ datapath_addsubunit_in1_2 }),
  .B({ S1766 }),
  .Y({ S1887 })
);
NOR #() 
NOR_487_ (
  .A({ S1886 }),
  .B({ S1887 }),
  .Y({ S1888 })
);
NAND #() 
NAND_1018_ (
  .A({ S1538 }),
  .B({ S1888 }),
  .Y({ S1889 })
);
NOR #() 
NOR_488_ (
  .A({ S1870 }),
  .B({ S1885 }),
  .Y({ S1890 })
);
NAND #() 
NAND_1019_ (
  .A({ S1889 }),
  .B({ S1890 }),
  .Y({ S1891 })
);
NOR #() 
NOR_489_ (
  .A({ S1868 }),
  .B({ S1891 }),
  .Y({ S1892 })
);
NAND #() 
NAND_1020_ (
  .A({ S1863 }),
  .B({ S1892 }),
  .Y({ datapath_indatatrf_2 })
);
NAND #() 
NAND_1021_ (
  .A({ datapath_indatatrf_2 }),
  .B({ S1688 }),
  .Y({ S1893 })
);
NAND #() 
NAND_1022_ (
  .A({ datapath_theregisterfile_memtrf_66 }),
  .B({ S1689 }),
  .Y({ S1894 })
);
NAND #() 
NAND_1023_ (
  .A({ S1893 }),
  .B({ S1894 }),
  .Y({ S6 })
);
NAND #() 
NAND_1024_ (
  .A({ datapath_addsubunit_in1_3 }),
  .B({ S1388 }),
  .Y({ S1895 })
);
NAND #() 
NAND_1025_ (
  .A({ controller_fib_3 }),
  .B({ S1409 }),
  .Y({ S1896 })
);
NAND #() 
NAND_1026_ (
  .A({ S1895 }),
  .B({ S1896 }),
  .Y({ S1897 })
);
NOT #() 
NOT_224_ (
  .A({ S1897 }),
  .Y({ S1898 })
);
NAND #() 
NAND_1027_ (
  .A({ S1417 }),
  .B({ S1897 }),
  .Y({ S1899 })
);
NOR #() 
NOR_490_ (
  .A({ controller_outflag_3 }),
  .B({ S1462 }),
  .Y({ S1900 })
);
NOT #() 
NOT_225_ (
  .A({ S1900 }),
  .Y({ S1901 })
);
NAND #() 
NAND_1028_ (
  .A({ datapath_theregisterfile_memtrf_243 }),
  .B({ S1437 }),
  .Y({ S1902 })
);
NAND #() 
NAND_1029_ (
  .A({ datapath_theregisterfile_memtrf_179 }),
  .B({ S1438 }),
  .Y({ S1903 })
);
NAND #() 
NAND_1030_ (
  .A({ S1902 }),
  .B({ S1903 }),
  .Y({ S1904 })
);
NAND #() 
NAND_1031_ (
  .A({ S1457 }),
  .B({ S1904 }),
  .Y({ S1905 })
);
NAND #() 
NAND_1032_ (
  .A({ datapath_theregisterfile_memtrf_163 }),
  .B({ S1438 }),
  .Y({ S1906 })
);
NAND #() 
NAND_1033_ (
  .A({ datapath_theregisterfile_memtrf_227 }),
  .B({ S1437 }),
  .Y({ S1907 })
);
NAND #() 
NAND_1034_ (
  .A({ S1906 }),
  .B({ S1907 }),
  .Y({ S1908 })
);
NAND #() 
NAND_1035_ (
  .A({ S1458 }),
  .B({ S1908 }),
  .Y({ S1909 })
);
NAND #() 
NAND_1036_ (
  .A({ S1905 }),
  .B({ S1909 }),
  .Y({ S1910 })
);
NAND #() 
NAND_1037_ (
  .A({ datapath_theregisterfile_memtrf_147 }),
  .B({ S1438 }),
  .Y({ S1911 })
);
NAND #() 
NAND_1038_ (
  .A({ datapath_theregisterfile_memtrf_211 }),
  .B({ S1437 }),
  .Y({ S1912 })
);
NAND #() 
NAND_1039_ (
  .A({ S1911 }),
  .B({ S1912 }),
  .Y({ S1913 })
);
NAND #() 
NAND_1040_ (
  .A({ S1457 }),
  .B({ S1913 }),
  .Y({ S1914 })
);
NOR #() 
NOR_491_ (
  .A({ datapath_theregisterfile_memtrf_131 }),
  .B({ S1437 }),
  .Y({ S1915 })
);
NAND #() 
NAND_1041_ (
  .A({ S7695 }),
  .B({ S1437 }),
  .Y({ S1916 })
);
NAND #() 
NAND_1042_ (
  .A({ S1458 }),
  .B({ S1916 }),
  .Y({ S1917 })
);
NOR #() 
NOR_492_ (
  .A({ S1915 }),
  .B({ S1917 }),
  .Y({ S1918 })
);
NOR #() 
NOR_493_ (
  .A({ S1444 }),
  .B({ S1910 }),
  .Y({ S1919 })
);
NOR #() 
NOR_494_ (
  .A({ S1443 }),
  .B({ S1918 }),
  .Y({ S1920 })
);
NAND #() 
NAND_1043_ (
  .A({ S1914 }),
  .B({ S1920 }),
  .Y({ S1921 })
);
NAND #() 
NAND_1044_ (
  .A({ S1449 }),
  .B({ S1921 }),
  .Y({ S1922 })
);
NOR #() 
NOR_495_ (
  .A({ S1919 }),
  .B({ S1922 }),
  .Y({ S1923 })
);
NAND #() 
NAND_1045_ (
  .A({ datapath_theregisterfile_memtrf_67 }),
  .B({ S1459 }),
  .Y({ S1924 })
);
NOT #() 
NOT_226_ (
  .A({ S1924 }),
  .Y({ S1925 })
);
NOR #() 
NOR_496_ (
  .A({ S1452 }),
  .B({ S1458 }),
  .Y({ S1926 })
);
NAND #() 
NAND_1046_ (
  .A({ datapath_theregisterfile_memtrf_19 }),
  .B({ S1438 }),
  .Y({ S1927 })
);
NAND #() 
NAND_1047_ (
  .A({ datapath_theregisterfile_memtrf_83 }),
  .B({ S1437 }),
  .Y({ S1928 })
);
NAND #() 
NAND_1048_ (
  .A({ S1927 }),
  .B({ S1928 }),
  .Y({ S1929 })
);
NAND #() 
NAND_1049_ (
  .A({ S1926 }),
  .B({ S1929 }),
  .Y({ S1930 })
);
NAND #() 
NAND_1050_ (
  .A({ S1462 }),
  .B({ S1930 }),
  .Y({ S1931 })
);
NOR #() 
NOR_497_ (
  .A({ S1925 }),
  .B({ S1931 }),
  .Y({ S1932 })
);
NAND #() 
NAND_1051_ (
  .A({ datapath_theregisterfile_memtrf_115 }),
  .B({ S1437 }),
  .Y({ S1933 })
);
NAND #() 
NAND_1052_ (
  .A({ datapath_theregisterfile_memtrf_51 }),
  .B({ S1438 }),
  .Y({ S1934 })
);
NAND #() 
NAND_1053_ (
  .A({ S1933 }),
  .B({ S1934 }),
  .Y({ S1935 })
);
NAND #() 
NAND_1054_ (
  .A({ S1457 }),
  .B({ S1935 }),
  .Y({ S1936 })
);
NAND #() 
NAND_1055_ (
  .A({ datapath_theregisterfile_memtrf_99 }),
  .B({ S1437 }),
  .Y({ S1937 })
);
NAND #() 
NAND_1056_ (
  .A({ datapath_theregisterfile_memtrf_35 }),
  .B({ S1438 }),
  .Y({ S1938 })
);
NAND #() 
NAND_1057_ (
  .A({ S1937 }),
  .B({ S1938 }),
  .Y({ S1939 })
);
NOT #() 
NOT_227_ (
  .A({ S1939 }),
  .Y({ S1940 })
);
NAND #() 
NAND_1058_ (
  .A({ S1458 }),
  .B({ S1939 }),
  .Y({ S1941 })
);
NAND #() 
NAND_1059_ (
  .A({ S1936 }),
  .B({ S1941 }),
  .Y({ S1942 })
);
NOR #() 
NOR_498_ (
  .A({ S1458 }),
  .B({ S1935 }),
  .Y({ S1943 })
);
NAND #() 
NAND_1060_ (
  .A({ S1458 }),
  .B({ S1940 }),
  .Y({ S1944 })
);
NAND #() 
NAND_1061_ (
  .A({ S1487 }),
  .B({ S1944 }),
  .Y({ S1945 })
);
NOR #() 
NOR_499_ (
  .A({ S1943 }),
  .B({ S1945 }),
  .Y({ S1946 })
);
NAND #() 
NAND_1062_ (
  .A({ S1487 }),
  .B({ S1942 }),
  .Y({ S1947 })
);
NAND #() 
NAND_1063_ (
  .A({ S1932 }),
  .B({ S1947 }),
  .Y({ S1948 })
);
NOR #() 
NOR_500_ (
  .A({ S1923 }),
  .B({ S1946 }),
  .Y({ S1949 })
);
NOR #() 
NOR_501_ (
  .A({ S1923 }),
  .B({ S1948 }),
  .Y({ S1950 })
);
NAND #() 
NAND_1064_ (
  .A({ S1932 }),
  .B({ S1949 }),
  .Y({ S1951 })
);
NOR #() 
NOR_502_ (
  .A({ S1900 }),
  .B({ S1950 }),
  .Y({ S1952 })
);
NAND #() 
NAND_1065_ (
  .A({ S1901 }),
  .B({ S1951 }),
  .Y({ S1953 })
);
NAND #() 
NAND_1066_ (
  .A({ S1429 }),
  .B({ S1952 }),
  .Y({ S1954 })
);
NAND #() 
NAND_1067_ (
  .A({ S1899 }),
  .B({ S1954 }),
  .Y({ S1955 })
);
NOT #() 
NOT_228_ (
  .A({ S1955 }),
  .Y({ S1956 })
);
NOR #() 
NOR_503_ (
  .A({ S1065 }),
  .B({ S1955 }),
  .Y({ S1957 })
);
NOR #() 
NOR_504_ (
  .A({ datapath_addsubunit_in1_3 }),
  .B({ S1956 }),
  .Y({ S1958 })
);
NOR #() 
NOR_505_ (
  .A({ S1065 }),
  .B({ S1956 }),
  .Y({ S1959 })
);
NOT #() 
NOT_229_ (
  .A({ S1959 }),
  .Y({ S1960 })
);
NOR #() 
NOR_506_ (
  .A({ datapath_addsubunit_in1_3 }),
  .B({ S1955 }),
  .Y({ S1961 })
);
NOR #() 
NOR_507_ (
  .A({ S1959 }),
  .B({ S1961 }),
  .Y({ S1962 })
);
NAND #() 
NAND_1068_ (
  .A({ S1866 }),
  .B({ S1869 }),
  .Y({ S1963 })
);
NOR #() 
NOR_508_ (
  .A({ S1962 }),
  .B({ S1963 }),
  .Y({ S1964 })
);
NAND #() 
NAND_1069_ (
  .A({ S1962 }),
  .B({ S1963 }),
  .Y({ S1965 })
);
NOR #() 
NOR_509_ (
  .A({ S1528 }),
  .B({ S1964 }),
  .Y({ S1966 })
);
NAND #() 
NAND_1070_ (
  .A({ S1965 }),
  .B({ S1966 }),
  .Y({ S1967 })
);
NOR #() 
NOR_510_ (
  .A({ S1855 }),
  .B({ S1859 }),
  .Y({ S1968 })
);
NOR #() 
NOR_511_ (
  .A({ S1962 }),
  .B({ S1968 }),
  .Y({ S1969 })
);
NAND #() 
NAND_1071_ (
  .A({ S1962 }),
  .B({ S1968 }),
  .Y({ S1970 })
);
NAND #() 
NAND_1072_ (
  .A({ S1525 }),
  .B({ S1970 }),
  .Y({ S1971 })
);
NOR #() 
NOR_512_ (
  .A({ S1969 }),
  .B({ S1971 }),
  .Y({ S1972 })
);
NOR #() 
NOR_513_ (
  .A({ S1533 }),
  .B({ S1960 }),
  .Y({ S1973 })
);
NAND #() 
NAND_1073_ (
  .A({ datapath_shiftunit_2189_A }),
  .B({ S1614 }),
  .Y({ S1974 })
);
NAND #() 
NAND_1074_ (
  .A({ datapath_shiftunit_2493_A }),
  .B({ S1609 }),
  .Y({ S1975 })
);
NOR #() 
NOR_514_ (
  .A({ datapath_muxmem_in2_3 }),
  .B({ S1337 }),
  .Y({ S1976 })
);
NOR #() 
NOR_515_ (
  .A({ S1339 }),
  .B({ S1976 }),
  .Y({ S1977 })
);
NOT #() 
NOT_230_ (
  .A({ S1977 }),
  .Y({ S1978 })
);
NAND #() 
NAND_1075_ (
  .A({ S1622 }),
  .B({ S1977 }),
  .Y({ S1979 })
);
NAND #() 
NAND_1076_ (
  .A({ datapath_multdivunit_outmdu2_3 }),
  .B({ S8570 }),
  .Y({ S1980 })
);
NAND #() 
NAND_1077_ (
  .A({ S1979 }),
  .B({ S1980 }),
  .Y({ S1981 })
);
NAND #() 
NAND_1078_ (
  .A({ datapath_multdivunit_outmdu1_3 }),
  .B({ S1377 }),
  .Y({ S1982 })
);
NAND #() 
NAND_1079_ (
  .A({ datapath_databusin_3 }),
  .B({ S1627 }),
  .Y({ S1983 })
);
NAND #() 
NAND_1080_ (
  .A({ S1982 }),
  .B({ S1983 }),
  .Y({ S1984 })
);
NOR #() 
NOR_516_ (
  .A({ S1981 }),
  .B({ S1984 }),
  .Y({ S1985 })
);
NAND #() 
NAND_1081_ (
  .A({ S1975 }),
  .B({ S1985 }),
  .Y({ S1986 })
);
NOR #() 
NOR_517_ (
  .A({ S1547 }),
  .B({ S1898 }),
  .Y({ S1987 })
);
NOR #() 
NOR_518_ (
  .A({ S1986 }),
  .B({ S1987 }),
  .Y({ S1988 })
);
NAND #() 
NAND_1082_ (
  .A({ S1974 }),
  .B({ S1988 }),
  .Y({ S1989 })
);
NOR #() 
NOR_519_ (
  .A({ S1973 }),
  .B({ S1989 }),
  .Y({ S1990 })
);
NOR #() 
NOR_520_ (
  .A({ S1065 }),
  .B({ S1887 }),
  .Y({ S1991 })
);
NAND #() 
NAND_1083_ (
  .A({ S1065 }),
  .B({ S1887 }),
  .Y({ S1992 })
);
NOR #() 
NOR_521_ (
  .A({ S1539 }),
  .B({ S1991 }),
  .Y({ S1993 })
);
NAND #() 
NAND_1084_ (
  .A({ S1992 }),
  .B({ S1993 }),
  .Y({ S1994 })
);
NAND #() 
NAND_1085_ (
  .A({ S1990 }),
  .B({ S1994 }),
  .Y({ S1995 })
);
NOR #() 
NOR_522_ (
  .A({ S1972 }),
  .B({ S1995 }),
  .Y({ S1996 })
);
NAND #() 
NAND_1086_ (
  .A({ S1967 }),
  .B({ S1996 }),
  .Y({ datapath_indatatrf_3 })
);
NAND #() 
NAND_1087_ (
  .A({ datapath_indatatrf_3 }),
  .B({ S1688 }),
  .Y({ S1997 })
);
NAND #() 
NAND_1088_ (
  .A({ datapath_theregisterfile_memtrf_67 }),
  .B({ S1689 }),
  .Y({ S1998 })
);
NAND #() 
NAND_1089_ (
  .A({ S1997 }),
  .B({ S1998 }),
  .Y({ S7 })
);
NAND #() 
NAND_1090_ (
  .A({ datapath_addsubunit_in1_4 }),
  .B({ S1388 }),
  .Y({ S1999 })
);
NAND #() 
NAND_1091_ (
  .A({ controller_fib_4 }),
  .B({ S1409 }),
  .Y({ S2000 })
);
NAND #() 
NAND_1092_ (
  .A({ S1999 }),
  .B({ S2000 }),
  .Y({ S2001 })
);
NOT #() 
NOT_231_ (
  .A({ S2001 }),
  .Y({ S2002 })
);
NAND #() 
NAND_1093_ (
  .A({ S1417 }),
  .B({ S2001 }),
  .Y({ S2003 })
);
NAND #() 
NAND_1094_ (
  .A({ S1429 }),
  .B({ S1597 }),
  .Y({ S2004 })
);
NAND #() 
NAND_1095_ (
  .A({ S2003 }),
  .B({ S2004 }),
  .Y({ S2005 })
);
NOT #() 
NOT_232_ (
  .A({ S2005 }),
  .Y({ S2006 })
);
NOR #() 
NOR_523_ (
  .A({ S1013 }),
  .B({ S2005 }),
  .Y({ S2007 })
);
NOT #() 
NOT_233_ (
  .A({ S2007 }),
  .Y({ S2008 })
);
NOR #() 
NOR_524_ (
  .A({ datapath_addsubunit_in1_4 }),
  .B({ S2006 }),
  .Y({ S2009 })
);
NOT #() 
NOT_234_ (
  .A({ S2009 }),
  .Y({ S2010 })
);
NAND #() 
NAND_1096_ (
  .A({ S2008 }),
  .B({ S2010 }),
  .Y({ S2011 })
);
NOR #() 
NOR_525_ (
  .A({ S1957 }),
  .B({ S1969 }),
  .Y({ S2012 })
);
NAND #() 
NAND_1097_ (
  .A({ S2011 }),
  .B({ S2012 }),
  .Y({ S2013 })
);
NOR #() 
NOR_526_ (
  .A({ S2011 }),
  .B({ S2012 }),
  .Y({ S2014 })
);
NAND #() 
NAND_1098_ (
  .A({ S1525 }),
  .B({ S2013 }),
  .Y({ S2015 })
);
NOR #() 
NOR_527_ (
  .A({ S2014 }),
  .B({ S2015 }),
  .Y({ S2016 })
);
NOR #() 
NOR_528_ (
  .A({ S1959 }),
  .B({ S1963 }),
  .Y({ S2017 })
);
NOR #() 
NOR_529_ (
  .A({ S1961 }),
  .B({ S2017 }),
  .Y({ S2018 })
);
NAND #() 
NAND_1099_ (
  .A({ S2011 }),
  .B({ S2018 }),
  .Y({ S2019 })
);
NOR #() 
NOR_530_ (
  .A({ S2011 }),
  .B({ S2018 }),
  .Y({ S2020 })
);
NOR #() 
NOR_531_ (
  .A({ S1528 }),
  .B({ S2020 }),
  .Y({ S2021 })
);
NAND #() 
NAND_1100_ (
  .A({ S2019 }),
  .B({ S2021 }),
  .Y({ S2022 })
);
NAND #() 
NAND_1101_ (
  .A({ datapath_addsubunit_in1_4 }),
  .B({ S2005 }),
  .Y({ S2023 })
);
NOR #() 
NOR_532_ (
  .A({ S1533 }),
  .B({ S2023 }),
  .Y({ S2024 })
);
NOR #() 
NOR_533_ (
  .A({ S1547 }),
  .B({ S2002 }),
  .Y({ S2025 })
);
NAND #() 
NAND_1102_ (
  .A({ datapath_shiftunit_2207_A }),
  .B({ S1614 }),
  .Y({ S2026 })
);
NAND #() 
NAND_1103_ (
  .A({ datapath_shiftunit_2511_A }),
  .B({ S1609 }),
  .Y({ S2027 })
);
NAND #() 
NAND_1104_ (
  .A({ S7913 }),
  .B({ S1340 }),
  .Y({ S2028 })
);
NAND #() 
NAND_1105_ (
  .A({ S1341 }),
  .B({ S2028 }),
  .Y({ S2029 })
);
NOR #() 
NOR_534_ (
  .A({ S1623 }),
  .B({ S2029 }),
  .Y({ S2030 })
);
NAND #() 
NAND_1106_ (
  .A({ datapath_databusin_4 }),
  .B({ S1627 }),
  .Y({ S2031 })
);
NAND #() 
NAND_1107_ (
  .A({ datapath_multdivunit_outmdu2_4 }),
  .B({ S8570 }),
  .Y({ S2032 })
);
NAND #() 
NAND_1108_ (
  .A({ datapath_multdivunit_outmdu1_4 }),
  .B({ S1377 }),
  .Y({ S2033 })
);
NAND #() 
NAND_1109_ (
  .A({ S2032 }),
  .B({ S2033 }),
  .Y({ S2034 })
);
NAND #() 
NAND_1110_ (
  .A({ S2026 }),
  .B({ S2027 }),
  .Y({ S2035 })
);
NOR #() 
NOR_535_ (
  .A({ S2025 }),
  .B({ S2035 }),
  .Y({ S2036 })
);
NOR #() 
NOR_536_ (
  .A({ S2030 }),
  .B({ S2034 }),
  .Y({ S2037 })
);
NAND #() 
NAND_1111_ (
  .A({ S2036 }),
  .B({ S2037 }),
  .Y({ S2038 })
);
NOT #() 
NOT_235_ (
  .A({ S2038 }),
  .Y({ S2039 })
);
NAND #() 
NAND_1112_ (
  .A({ S2031 }),
  .B({ S2039 }),
  .Y({ S2040 })
);
NOR #() 
NOR_537_ (
  .A({ S2024 }),
  .B({ S2040 }),
  .Y({ S2041 })
);
NAND #() 
NAND_1113_ (
  .A({ datapath_addsubunit_in1_4 }),
  .B({ S1992 }),
  .Y({ S2042 })
);
NOR #() 
NOR_538_ (
  .A({ datapath_addsubunit_in1_4 }),
  .B({ S1992 }),
  .Y({ S2043 })
);
NOR #() 
NOR_539_ (
  .A({ S1539 }),
  .B({ S2043 }),
  .Y({ S2044 })
);
NAND #() 
NAND_1114_ (
  .A({ S2042 }),
  .B({ S2044 }),
  .Y({ S2045 })
);
NAND #() 
NAND_1115_ (
  .A({ S2041 }),
  .B({ S2045 }),
  .Y({ S2046 })
);
NOR #() 
NOR_540_ (
  .A({ S2016 }),
  .B({ S2046 }),
  .Y({ S2047 })
);
NAND #() 
NAND_1116_ (
  .A({ S2022 }),
  .B({ S2047 }),
  .Y({ datapath_indatatrf_4 })
);
NAND #() 
NAND_1117_ (
  .A({ datapath_indatatrf_4 }),
  .B({ S1688 }),
  .Y({ S2048 })
);
NAND #() 
NAND_1118_ (
  .A({ datapath_theregisterfile_memtrf_68 }),
  .B({ S1689 }),
  .Y({ S2049 })
);
NAND #() 
NAND_1119_ (
  .A({ S2048 }),
  .B({ S2049 }),
  .Y({ S8 })
);
NOR #() 
NOR_541_ (
  .A({ S963 }),
  .B({ S1389 }),
  .Y({ S2050 })
);
NAND #() 
NAND_1120_ (
  .A({ controller_216_B_0 }),
  .B({ S1401 }),
  .Y({ S2051 })
);
NAND #() 
NAND_1121_ (
  .A({ controller_fib_4 }),
  .B({ S1406 }),
  .Y({ S2052 })
);
NAND #() 
NAND_1122_ (
  .A({ S372 }),
  .B({ S2052 }),
  .Y({ S2053 })
);
NOT #() 
NOT_236_ (
  .A({ S2053 }),
  .Y({ S2054 })
);
NOR #() 
NOR_542_ (
  .A({ S2050 }),
  .B({ S2053 }),
  .Y({ S2055 })
);
NAND #() 
NAND_1123_ (
  .A({ S2051 }),
  .B({ S2055 }),
  .Y({ S2056 })
);
NAND #() 
NAND_1124_ (
  .A({ S1417 }),
  .B({ S2056 }),
  .Y({ S2057 })
);
NOR #() 
NOR_543_ (
  .A({ controller_389_B_2 }),
  .B({ S1462 }),
  .Y({ S2058 })
);
NOT #() 
NOT_237_ (
  .A({ S2058 }),
  .Y({ S2059 })
);
NAND #() 
NAND_1125_ (
  .A({ datapath_theregisterfile_memtrf_245 }),
  .B({ S1437 }),
  .Y({ S2060 })
);
NAND #() 
NAND_1126_ (
  .A({ datapath_theregisterfile_memtrf_181 }),
  .B({ S1438 }),
  .Y({ S2061 })
);
NAND #() 
NAND_1127_ (
  .A({ S2060 }),
  .B({ S2061 }),
  .Y({ S2062 })
);
NAND #() 
NAND_1128_ (
  .A({ S1457 }),
  .B({ S2062 }),
  .Y({ S2063 })
);
NAND #() 
NAND_1129_ (
  .A({ S7822 }),
  .B({ S1437 }),
  .Y({ S2064 })
);
NOR #() 
NOR_544_ (
  .A({ datapath_theregisterfile_memtrf_165 }),
  .B({ S1437 }),
  .Y({ S2065 })
);
NAND #() 
NAND_1130_ (
  .A({ S1458 }),
  .B({ S2064 }),
  .Y({ S2066 })
);
NOR #() 
NOR_545_ (
  .A({ S2065 }),
  .B({ S2066 }),
  .Y({ S2067 })
);
NAND #() 
NAND_1131_ (
  .A({ datapath_theregisterfile_memtrf_149 }),
  .B({ S1438 }),
  .Y({ S2068 })
);
NAND #() 
NAND_1132_ (
  .A({ datapath_theregisterfile_memtrf_213 }),
  .B({ S1437 }),
  .Y({ S2069 })
);
NAND #() 
NAND_1133_ (
  .A({ S2068 }),
  .B({ S2069 }),
  .Y({ S2070 })
);
NAND #() 
NAND_1134_ (
  .A({ S1457 }),
  .B({ S2070 }),
  .Y({ S2071 })
);
NOR #() 
NOR_546_ (
  .A({ datapath_theregisterfile_memtrf_133 }),
  .B({ S1437 }),
  .Y({ S2072 })
);
NOR #() 
NOR_547_ (
  .A({ datapath_theregisterfile_memtrf_197 }),
  .B({ S1438 }),
  .Y({ S2073 })
);
NOR #() 
NOR_548_ (
  .A({ S2072 }),
  .B({ S2073 }),
  .Y({ S2074 })
);
NAND #() 
NAND_1135_ (
  .A({ S1458 }),
  .B({ S2074 }),
  .Y({ S2075 })
);
NAND #() 
NAND_1136_ (
  .A({ S2071 }),
  .B({ S2075 }),
  .Y({ S2076 })
);
NOR #() 
NOR_549_ (
  .A({ S1443 }),
  .B({ S2076 }),
  .Y({ S2077 })
);
NOR #() 
NOR_550_ (
  .A({ S1444 }),
  .B({ S2067 }),
  .Y({ S2078 })
);
NAND #() 
NAND_1137_ (
  .A({ S2063 }),
  .B({ S2078 }),
  .Y({ S2079 })
);
NAND #() 
NAND_1138_ (
  .A({ S1449 }),
  .B({ S2079 }),
  .Y({ S2080 })
);
NOR #() 
NOR_551_ (
  .A({ S2077 }),
  .B({ S2080 }),
  .Y({ S2081 })
);
NAND #() 
NAND_1139_ (
  .A({ datapath_theregisterfile_memtrf_101 }),
  .B({ S1458 }),
  .Y({ S2082 })
);
NAND #() 
NAND_1140_ (
  .A({ datapath_theregisterfile_memtrf_117 }),
  .B({ S1457 }),
  .Y({ S2083 })
);
NAND #() 
NAND_1141_ (
  .A({ S2082 }),
  .B({ S2083 }),
  .Y({ S2084 })
);
NAND #() 
NAND_1142_ (
  .A({ S1437 }),
  .B({ S2084 }),
  .Y({ S2085 })
);
NAND #() 
NAND_1143_ (
  .A({ datapath_theregisterfile_memtrf_37 }),
  .B({ S1458 }),
  .Y({ S2086 })
);
NAND #() 
NAND_1144_ (
  .A({ datapath_theregisterfile_memtrf_53 }),
  .B({ S1457 }),
  .Y({ S2087 })
);
NAND #() 
NAND_1145_ (
  .A({ S2086 }),
  .B({ S2087 }),
  .Y({ S2088 })
);
NAND #() 
NAND_1146_ (
  .A({ S1438 }),
  .B({ S2088 }),
  .Y({ S2089 })
);
NAND #() 
NAND_1147_ (
  .A({ S2085 }),
  .B({ S2089 }),
  .Y({ S2090 })
);
NAND #() 
NAND_1148_ (
  .A({ S1487 }),
  .B({ S2090 }),
  .Y({ S2091 })
);
NAND #() 
NAND_1149_ (
  .A({ datapath_theregisterfile_memtrf_85 }),
  .B({ S1498 }),
  .Y({ S2092 })
);
NOR #() 
NOR_552_ (
  .A({ datapath_theregisterfile_memtrf_69 }),
  .B({ S1438 }),
  .Y({ S2093 })
);
NOT #() 
NOT_238_ (
  .A({ S2093 }),
  .Y({ S2094 })
);
NAND #() 
NAND_1150_ (
  .A({ datapath_theregisterfile_memtrf_21 }),
  .B({ S1438 }),
  .Y({ S2095 })
);
NAND #() 
NAND_1151_ (
  .A({ S1457 }),
  .B({ S2095 }),
  .Y({ S2096 })
);
NAND #() 
NAND_1152_ (
  .A({ S2094 }),
  .B({ S2096 }),
  .Y({ S2097 })
);
NAND #() 
NAND_1153_ (
  .A({ S2092 }),
  .B({ S2097 }),
  .Y({ S2098 })
);
NOT #() 
NOT_239_ (
  .A({ S2098 }),
  .Y({ S2099 })
);
NOR #() 
NOR_553_ (
  .A({ S1452 }),
  .B({ S2099 }),
  .Y({ S2100 })
);
NAND #() 
NAND_1154_ (
  .A({ S1451 }),
  .B({ S2098 }),
  .Y({ S2101 })
);
NAND #() 
NAND_1155_ (
  .A({ S2091 }),
  .B({ S2101 }),
  .Y({ S2102 })
);
NOR #() 
NOR_554_ (
  .A({ S2081 }),
  .B({ S2100 }),
  .Y({ S2103 })
);
NOR #() 
NOR_555_ (
  .A({ S2081 }),
  .B({ S2102 }),
  .Y({ S2104 })
);
NAND #() 
NAND_1156_ (
  .A({ S2091 }),
  .B({ S2103 }),
  .Y({ S2105 })
);
NOR #() 
NOR_556_ (
  .A({ S2058 }),
  .B({ S2104 }),
  .Y({ S2106 })
);
NAND #() 
NAND_1157_ (
  .A({ S2059 }),
  .B({ S2105 }),
  .Y({ S2107 })
);
NAND #() 
NAND_1158_ (
  .A({ S1429 }),
  .B({ S2106 }),
  .Y({ S2108 })
);
NAND #() 
NAND_1159_ (
  .A({ S2057 }),
  .B({ S2108 }),
  .Y({ S2109 })
);
NOR #() 
NOR_557_ (
  .A({ S963 }),
  .B({ S2109 }),
  .Y({ S2110 })
);
NOT #() 
NOT_240_ (
  .A({ S2110 }),
  .Y({ S2111 })
);
NAND #() 
NAND_1160_ (
  .A({ S963 }),
  .B({ S2109 }),
  .Y({ S2112 })
);
NAND #() 
NAND_1161_ (
  .A({ S2111 }),
  .B({ S2112 }),
  .Y({ S2113 })
);
NOR #() 
NOR_558_ (
  .A({ S2007 }),
  .B({ S2014 }),
  .Y({ S2114 })
);
NAND #() 
NAND_1162_ (
  .A({ S2113 }),
  .B({ S2114 }),
  .Y({ S2115 })
);
NOR #() 
NOR_559_ (
  .A({ S2113 }),
  .B({ S2114 }),
  .Y({ S2116 })
);
NAND #() 
NAND_1163_ (
  .A({ S1525 }),
  .B({ S2115 }),
  .Y({ S2117 })
);
NOR #() 
NOR_560_ (
  .A({ S2116 }),
  .B({ S2117 }),
  .Y({ S2118 })
);
NAND #() 
NAND_1164_ (
  .A({ S2019 }),
  .B({ S2023 }),
  .Y({ S2119 })
);
NAND #() 
NAND_1165_ (
  .A({ S2113 }),
  .B({ S2119 }),
  .Y({ S2120 })
);
NOR #() 
NOR_561_ (
  .A({ S2113 }),
  .B({ S2119 }),
  .Y({ S2121 })
);
NOR #() 
NOR_562_ (
  .A({ S1528 }),
  .B({ S2121 }),
  .Y({ S2122 })
);
NAND #() 
NAND_1166_ (
  .A({ S2120 }),
  .B({ S2122 }),
  .Y({ S2123 })
);
NOR #() 
NOR_563_ (
  .A({ S963 }),
  .B({ S2043 }),
  .Y({ S2124 })
);
NAND #() 
NAND_1167_ (
  .A({ S963 }),
  .B({ S2043 }),
  .Y({ S2125 })
);
NOT #() 
NOT_241_ (
  .A({ S2125 }),
  .Y({ S2126 })
);
NOR #() 
NOR_564_ (
  .A({ S2124 }),
  .B({ S2126 }),
  .Y({ S2127 })
);
NAND #() 
NAND_1168_ (
  .A({ S1538 }),
  .B({ S2127 }),
  .Y({ S2128 })
);
NAND #() 
NAND_1169_ (
  .A({ datapath_addsubunit_in1_5 }),
  .B({ S2109 }),
  .Y({ S2129 })
);
NOR #() 
NOR_565_ (
  .A({ S1533 }),
  .B({ S2129 }),
  .Y({ S2130 })
);
NAND #() 
NAND_1170_ (
  .A({ S1546 }),
  .B({ S2056 }),
  .Y({ S2131 })
);
NAND #() 
NAND_1171_ (
  .A({ datapath_shiftunit_2225_A }),
  .B({ S1614 }),
  .Y({ S2132 })
);
NOT #() 
NOT_242_ (
  .A({ S2132 }),
  .Y({ S2133 })
);
NAND #() 
NAND_1172_ (
  .A({ datapath_shiftunit_2529_A }),
  .B({ S1609 }),
  .Y({ S2134 })
);
NAND #() 
NAND_1173_ (
  .A({ S7920 }),
  .B({ S1341 }),
  .Y({ S2135 })
);
NAND #() 
NAND_1174_ (
  .A({ S1344 }),
  .B({ S2135 }),
  .Y({ S2136 })
);
NOR #() 
NOR_566_ (
  .A({ S1623 }),
  .B({ S2136 }),
  .Y({ S2137 })
);
NOR #() 
NOR_567_ (
  .A({ S8236 }),
  .B({ S1628 }),
  .Y({ S2138 })
);
NAND #() 
NAND_1175_ (
  .A({ datapath_multdivunit_outmdu1_5 }),
  .B({ S1377 }),
  .Y({ S2139 })
);
NOR #() 
NOR_568_ (
  .A({ S8087 }),
  .B({ S8571 }),
  .Y({ S2140 })
);
NOR #() 
NOR_569_ (
  .A({ S2138 }),
  .B({ S2140 }),
  .Y({ S2141 })
);
NAND #() 
NAND_1176_ (
  .A({ S2139 }),
  .B({ S2141 }),
  .Y({ S2142 })
);
NOR #() 
NOR_570_ (
  .A({ S2137 }),
  .B({ S2142 }),
  .Y({ S2143 })
);
NAND #() 
NAND_1177_ (
  .A({ S2134 }),
  .B({ S2143 }),
  .Y({ S2144 })
);
NOR #() 
NOR_571_ (
  .A({ S2133 }),
  .B({ S2144 }),
  .Y({ S2145 })
);
NAND #() 
NAND_1178_ (
  .A({ S2131 }),
  .B({ S2145 }),
  .Y({ S2146 })
);
NOR #() 
NOR_572_ (
  .A({ S2130 }),
  .B({ S2146 }),
  .Y({ S2147 })
);
NAND #() 
NAND_1179_ (
  .A({ S2128 }),
  .B({ S2147 }),
  .Y({ S2148 })
);
NOR #() 
NOR_573_ (
  .A({ S2118 }),
  .B({ S2148 }),
  .Y({ S2149 })
);
NAND #() 
NAND_1180_ (
  .A({ S2123 }),
  .B({ S2149 }),
  .Y({ datapath_indatatrf_5 })
);
NAND #() 
NAND_1181_ (
  .A({ datapath_indatatrf_5 }),
  .B({ S1688 }),
  .Y({ S2150 })
);
NAND #() 
NAND_1182_ (
  .A({ datapath_theregisterfile_memtrf_69 }),
  .B({ S1689 }),
  .Y({ S2151 })
);
NAND #() 
NAND_1183_ (
  .A({ S2150 }),
  .B({ S2151 }),
  .Y({ S9 })
);
NOR #() 
NOR_574_ (
  .A({ S910 }),
  .B({ S1389 }),
  .Y({ S2152 })
);
NAND #() 
NAND_1184_ (
  .A({ controller_opcode_2 }),
  .B({ S1401 }),
  .Y({ S2153 })
);
NAND #() 
NAND_1185_ (
  .A({ S2054 }),
  .B({ S2153 }),
  .Y({ S2154 })
);
NOR #() 
NOR_575_ (
  .A({ S2152 }),
  .B({ S2154 }),
  .Y({ S2155 })
);
NOR #() 
NOR_576_ (
  .A({ S1416 }),
  .B({ S2155 }),
  .Y({ S2156 })
);
NOR #() 
NOR_577_ (
  .A({ controller_outflag_6 }),
  .B({ S1462 }),
  .Y({ S2157 })
);
NOT #() 
NOT_243_ (
  .A({ S2157 }),
  .Y({ S2158 })
);
NAND #() 
NAND_1186_ (
  .A({ datapath_theregisterfile_memtrf_246 }),
  .B({ S1437 }),
  .Y({ S2159 })
);
NAND #() 
NAND_1187_ (
  .A({ datapath_theregisterfile_memtrf_182 }),
  .B({ S1438 }),
  .Y({ S2160 })
);
NAND #() 
NAND_1188_ (
  .A({ S2159 }),
  .B({ S2160 }),
  .Y({ S2161 })
);
NAND #() 
NAND_1189_ (
  .A({ S1457 }),
  .B({ S2161 }),
  .Y({ S2162 })
);
NAND #() 
NAND_1190_ (
  .A({ S7823 }),
  .B({ S1437 }),
  .Y({ S2163 })
);
NOR #() 
NOR_578_ (
  .A({ datapath_theregisterfile_memtrf_166 }),
  .B({ S1437 }),
  .Y({ S2164 })
);
NAND #() 
NAND_1191_ (
  .A({ S1458 }),
  .B({ S2163 }),
  .Y({ S2165 })
);
NOR #() 
NOR_579_ (
  .A({ S2164 }),
  .B({ S2165 }),
  .Y({ S2166 })
);
NAND #() 
NAND_1192_ (
  .A({ datapath_theregisterfile_memtrf_150 }),
  .B({ S1438 }),
  .Y({ S2167 })
);
NAND #() 
NAND_1193_ (
  .A({ datapath_theregisterfile_memtrf_214 }),
  .B({ S1437 }),
  .Y({ S2168 })
);
NAND #() 
NAND_1194_ (
  .A({ S2167 }),
  .B({ S2168 }),
  .Y({ S2169 })
);
NAND #() 
NAND_1195_ (
  .A({ S1457 }),
  .B({ S2169 }),
  .Y({ S2170 })
);
NOR #() 
NOR_580_ (
  .A({ datapath_theregisterfile_memtrf_134 }),
  .B({ S1437 }),
  .Y({ S2171 })
);
NOR #() 
NOR_581_ (
  .A({ datapath_theregisterfile_memtrf_198 }),
  .B({ S1438 }),
  .Y({ S2172 })
);
NOR #() 
NOR_582_ (
  .A({ S2171 }),
  .B({ S2172 }),
  .Y({ S2173 })
);
NAND #() 
NAND_1196_ (
  .A({ S1458 }),
  .B({ S2173 }),
  .Y({ S2174 })
);
NAND #() 
NAND_1197_ (
  .A({ S2170 }),
  .B({ S2174 }),
  .Y({ S2175 })
);
NOR #() 
NOR_583_ (
  .A({ S1443 }),
  .B({ S2175 }),
  .Y({ S2176 })
);
NOR #() 
NOR_584_ (
  .A({ S1444 }),
  .B({ S2166 }),
  .Y({ S2177 })
);
NAND #() 
NAND_1198_ (
  .A({ S2162 }),
  .B({ S2177 }),
  .Y({ S2178 })
);
NAND #() 
NAND_1199_ (
  .A({ S1449 }),
  .B({ S2178 }),
  .Y({ S2179 })
);
NOR #() 
NOR_585_ (
  .A({ S2176 }),
  .B({ S2179 }),
  .Y({ S2180 })
);
NAND #() 
NAND_1200_ (
  .A({ datapath_theregisterfile_memtrf_102 }),
  .B({ S1458 }),
  .Y({ S2181 })
);
NAND #() 
NAND_1201_ (
  .A({ datapath_theregisterfile_memtrf_118 }),
  .B({ S1457 }),
  .Y({ S2182 })
);
NAND #() 
NAND_1202_ (
  .A({ S2181 }),
  .B({ S2182 }),
  .Y({ S2183 })
);
NAND #() 
NAND_1203_ (
  .A({ S1437 }),
  .B({ S2183 }),
  .Y({ S2184 })
);
NAND #() 
NAND_1204_ (
  .A({ datapath_theregisterfile_memtrf_38 }),
  .B({ S1458 }),
  .Y({ S2185 })
);
NAND #() 
NAND_1205_ (
  .A({ datapath_theregisterfile_memtrf_54 }),
  .B({ S1457 }),
  .Y({ S2186 })
);
NAND #() 
NAND_1206_ (
  .A({ S2185 }),
  .B({ S2186 }),
  .Y({ S2187 })
);
NAND #() 
NAND_1207_ (
  .A({ S1438 }),
  .B({ S2187 }),
  .Y({ S2188 })
);
NAND #() 
NAND_1208_ (
  .A({ S2184 }),
  .B({ S2188 }),
  .Y({ S2189 })
);
NAND #() 
NAND_1209_ (
  .A({ S1487 }),
  .B({ S2189 }),
  .Y({ S2190 })
);
NAND #() 
NAND_1210_ (
  .A({ datapath_theregisterfile_memtrf_86 }),
  .B({ S1498 }),
  .Y({ S2191 })
);
NOR #() 
NOR_586_ (
  .A({ datapath_theregisterfile_memtrf_70 }),
  .B({ S1438 }),
  .Y({ S2192 })
);
NOT #() 
NOT_244_ (
  .A({ S2192 }),
  .Y({ S2193 })
);
NAND #() 
NAND_1211_ (
  .A({ datapath_theregisterfile_memtrf_22 }),
  .B({ S1438 }),
  .Y({ S2194 })
);
NAND #() 
NAND_1212_ (
  .A({ S1457 }),
  .B({ S2194 }),
  .Y({ S2195 })
);
NAND #() 
NAND_1213_ (
  .A({ S2193 }),
  .B({ S2195 }),
  .Y({ S2196 })
);
NAND #() 
NAND_1214_ (
  .A({ S2191 }),
  .B({ S2196 }),
  .Y({ S2197 })
);
NOT #() 
NOT_245_ (
  .A({ S2197 }),
  .Y({ S2198 })
);
NOR #() 
NOR_587_ (
  .A({ S1452 }),
  .B({ S2198 }),
  .Y({ S2199 })
);
NAND #() 
NAND_1215_ (
  .A({ S1451 }),
  .B({ S2197 }),
  .Y({ S2200 })
);
NAND #() 
NAND_1216_ (
  .A({ S2190 }),
  .B({ S2200 }),
  .Y({ S2201 })
);
NOR #() 
NOR_588_ (
  .A({ S2180 }),
  .B({ S2199 }),
  .Y({ S2202 })
);
NOR #() 
NOR_589_ (
  .A({ S2180 }),
  .B({ S2201 }),
  .Y({ S2203 })
);
NAND #() 
NAND_1217_ (
  .A({ S2190 }),
  .B({ S2202 }),
  .Y({ S2204 })
);
NOR #() 
NOR_590_ (
  .A({ S2157 }),
  .B({ S2203 }),
  .Y({ S2205 })
);
NAND #() 
NAND_1218_ (
  .A({ S2158 }),
  .B({ S2204 }),
  .Y({ S2206 })
);
NOR #() 
NOR_591_ (
  .A({ S1430 }),
  .B({ S2206 }),
  .Y({ S2207 })
);
NOR #() 
NOR_592_ (
  .A({ S2156 }),
  .B({ S2207 }),
  .Y({ S2208 })
);
NOT #() 
NOT_246_ (
  .A({ S2208 }),
  .Y({ S2209 })
);
NOR #() 
NOR_593_ (
  .A({ datapath_addsubunit_in1_6 }),
  .B({ S2208 }),
  .Y({ S2210 })
);
NOT #() 
NOT_247_ (
  .A({ S2210 }),
  .Y({ S2211 })
);
NOR #() 
NOR_594_ (
  .A({ S910 }),
  .B({ S2209 }),
  .Y({ S2212 })
);
NOR #() 
NOR_595_ (
  .A({ S2210 }),
  .B({ S2212 }),
  .Y({ S2213 })
);
NAND #() 
NAND_1219_ (
  .A({ S2111 }),
  .B({ S2114 }),
  .Y({ S2214 })
);
NAND #() 
NAND_1220_ (
  .A({ S2112 }),
  .B({ S2214 }),
  .Y({ S2215 })
);
NOT #() 
NOT_248_ (
  .A({ S2215 }),
  .Y({ S2216 })
);
NOR #() 
NOR_596_ (
  .A({ S2213 }),
  .B({ S2216 }),
  .Y({ S2217 })
);
NAND #() 
NAND_1221_ (
  .A({ S2213 }),
  .B({ S2216 }),
  .Y({ S2218 })
);
NOT #() 
NOT_249_ (
  .A({ S2218 }),
  .Y({ S2219 })
);
NAND #() 
NAND_1222_ (
  .A({ S1525 }),
  .B({ S2218 }),
  .Y({ S2220 })
);
NOR #() 
NOR_597_ (
  .A({ S2217 }),
  .B({ S2220 }),
  .Y({ S2221 })
);
NAND #() 
NAND_1223_ (
  .A({ S2120 }),
  .B({ S2129 }),
  .Y({ S2222 })
);
NOT #() 
NOT_250_ (
  .A({ S2222 }),
  .Y({ S2223 })
);
NAND #() 
NAND_1224_ (
  .A({ S2213 }),
  .B({ S2223 }),
  .Y({ S2224 })
);
NOR #() 
NOR_598_ (
  .A({ S2213 }),
  .B({ S2223 }),
  .Y({ S2225 })
);
NOR #() 
NOR_599_ (
  .A({ S1528 }),
  .B({ S2225 }),
  .Y({ S2226 })
);
NAND #() 
NAND_1225_ (
  .A({ S2224 }),
  .B({ S2226 }),
  .Y({ S2227 })
);
NOR #() 
NOR_600_ (
  .A({ S910 }),
  .B({ S2208 }),
  .Y({ S2228 })
);
NOT #() 
NOT_251_ (
  .A({ S2228 }),
  .Y({ S2229 })
);
NOR #() 
NOR_601_ (
  .A({ S1533 }),
  .B({ S2229 }),
  .Y({ S2230 })
);
NOR #() 
NOR_602_ (
  .A({ S1547 }),
  .B({ S2155 }),
  .Y({ S2231 })
);
NAND #() 
NAND_1226_ (
  .A({ datapath_shiftunit_2243_A }),
  .B({ S1614 }),
  .Y({ S2232 })
);
NAND #() 
NAND_1227_ (
  .A({ datapath_shiftunit_2547_A }),
  .B({ S1609 }),
  .Y({ S2233 })
);
NAND #() 
NAND_1228_ (
  .A({ S7928 }),
  .B({ S1344 }),
  .Y({ S2234 })
);
NAND #() 
NAND_1229_ (
  .A({ S1346 }),
  .B({ S2234 }),
  .Y({ S2235 })
);
NOR #() 
NOR_603_ (
  .A({ S1623 }),
  .B({ S2235 }),
  .Y({ S2236 })
);
NAND #() 
NAND_1230_ (
  .A({ datapath_multdivunit_outmdu2_6 }),
  .B({ S8570 }),
  .Y({ S2237 })
);
NOR #() 
NOR_604_ (
  .A({ S8022 }),
  .B({ S1378 }),
  .Y({ S2238 })
);
NOR #() 
NOR_605_ (
  .A({ S8257 }),
  .B({ S1628 }),
  .Y({ S2239 })
);
NOR #() 
NOR_606_ (
  .A({ S2238 }),
  .B({ S2239 }),
  .Y({ S2240 })
);
NAND #() 
NAND_1231_ (
  .A({ S2237 }),
  .B({ S2240 }),
  .Y({ S2241 })
);
NOR #() 
NOR_607_ (
  .A({ S2236 }),
  .B({ S2241 }),
  .Y({ S2242 })
);
NAND #() 
NAND_1232_ (
  .A({ S2232 }),
  .B({ S2233 }),
  .Y({ S2243 })
);
NOR #() 
NOR_608_ (
  .A({ S2231 }),
  .B({ S2243 }),
  .Y({ S2244 })
);
NAND #() 
NAND_1233_ (
  .A({ S2242 }),
  .B({ S2244 }),
  .Y({ S2245 })
);
NOR #() 
NOR_609_ (
  .A({ S2230 }),
  .B({ S2245 }),
  .Y({ S2246 })
);
NAND #() 
NAND_1234_ (
  .A({ datapath_addsubunit_in1_6 }),
  .B({ S2125 }),
  .Y({ S2247 })
);
NOR #() 
NOR_610_ (
  .A({ datapath_addsubunit_in1_6 }),
  .B({ S2125 }),
  .Y({ S2248 })
);
NOR #() 
NOR_611_ (
  .A({ S1539 }),
  .B({ S2248 }),
  .Y({ S2249 })
);
NAND #() 
NAND_1235_ (
  .A({ S2247 }),
  .B({ S2249 }),
  .Y({ S2250 })
);
NAND #() 
NAND_1236_ (
  .A({ S2246 }),
  .B({ S2250 }),
  .Y({ S2251 })
);
NOR #() 
NOR_612_ (
  .A({ S2221 }),
  .B({ S2251 }),
  .Y({ S2252 })
);
NAND #() 
NAND_1237_ (
  .A({ S2227 }),
  .B({ S2252 }),
  .Y({ datapath_indatatrf_6 })
);
NAND #() 
NAND_1238_ (
  .A({ datapath_indatatrf_6 }),
  .B({ S1688 }),
  .Y({ S2253 })
);
NAND #() 
NAND_1239_ (
  .A({ datapath_theregisterfile_memtrf_70 }),
  .B({ S1689 }),
  .Y({ S2254 })
);
NAND #() 
NAND_1240_ (
  .A({ S2253 }),
  .B({ S2254 }),
  .Y({ S10 })
);
NOR #() 
NOR_613_ (
  .A({ S858 }),
  .B({ S1389 }),
  .Y({ S2255 })
);
NAND #() 
NAND_1241_ (
  .A({ controller_opcode_3 }),
  .B({ S1401 }),
  .Y({ S2256 })
);
NOR #() 
NOR_614_ (
  .A({ S2053 }),
  .B({ S2255 }),
  .Y({ S2257 })
);
NAND #() 
NAND_1242_ (
  .A({ S2256 }),
  .B({ S2257 }),
  .Y({ S2258 })
);
NAND #() 
NAND_1243_ (
  .A({ S1417 }),
  .B({ S2258 }),
  .Y({ S2259 })
);
NOR #() 
NOR_615_ (
  .A({ controller_outflag_7 }),
  .B({ S1462 }),
  .Y({ S2260 })
);
NOT #() 
NOT_252_ (
  .A({ S2260 }),
  .Y({ S2261 })
);
NAND #() 
NAND_1244_ (
  .A({ datapath_theregisterfile_memtrf_247 }),
  .B({ S1437 }),
  .Y({ S2262 })
);
NAND #() 
NAND_1245_ (
  .A({ datapath_theregisterfile_memtrf_183 }),
  .B({ S1438 }),
  .Y({ S2263 })
);
NAND #() 
NAND_1246_ (
  .A({ S2262 }),
  .B({ S2263 }),
  .Y({ S2264 })
);
NAND #() 
NAND_1247_ (
  .A({ S1457 }),
  .B({ S2264 }),
  .Y({ S2265 })
);
NAND #() 
NAND_1248_ (
  .A({ datapath_theregisterfile_memtrf_167 }),
  .B({ S1438 }),
  .Y({ S2266 })
);
NAND #() 
NAND_1249_ (
  .A({ datapath_theregisterfile_memtrf_231 }),
  .B({ S1437 }),
  .Y({ S2267 })
);
NAND #() 
NAND_1250_ (
  .A({ S2266 }),
  .B({ S2267 }),
  .Y({ S2268 })
);
NAND #() 
NAND_1251_ (
  .A({ S1458 }),
  .B({ S2268 }),
  .Y({ S2269 })
);
NAND #() 
NAND_1252_ (
  .A({ S2265 }),
  .B({ S2269 }),
  .Y({ S2270 })
);
NAND #() 
NAND_1253_ (
  .A({ datapath_theregisterfile_memtrf_151 }),
  .B({ S1438 }),
  .Y({ S2271 })
);
NAND #() 
NAND_1254_ (
  .A({ datapath_theregisterfile_memtrf_215 }),
  .B({ S1437 }),
  .Y({ S2272 })
);
NAND #() 
NAND_1255_ (
  .A({ S2271 }),
  .B({ S2272 }),
  .Y({ S2273 })
);
NAND #() 
NAND_1256_ (
  .A({ S1457 }),
  .B({ S2273 }),
  .Y({ S2274 })
);
NOR #() 
NOR_616_ (
  .A({ datapath_theregisterfile_memtrf_135 }),
  .B({ S1437 }),
  .Y({ S2275 })
);
NAND #() 
NAND_1257_ (
  .A({ S7728 }),
  .B({ S1437 }),
  .Y({ S2276 })
);
NAND #() 
NAND_1258_ (
  .A({ S1458 }),
  .B({ S2276 }),
  .Y({ S2277 })
);
NOR #() 
NOR_617_ (
  .A({ S2275 }),
  .B({ S2277 }),
  .Y({ S2278 })
);
NOR #() 
NOR_618_ (
  .A({ S1444 }),
  .B({ S2270 }),
  .Y({ S2279 })
);
NOR #() 
NOR_619_ (
  .A({ S1443 }),
  .B({ S2278 }),
  .Y({ S2280 })
);
NAND #() 
NAND_1259_ (
  .A({ S2274 }),
  .B({ S2280 }),
  .Y({ S2281 })
);
NAND #() 
NAND_1260_ (
  .A({ S1449 }),
  .B({ S2281 }),
  .Y({ S2282 })
);
NOR #() 
NOR_620_ (
  .A({ S2279 }),
  .B({ S2282 }),
  .Y({ S2283 })
);
NAND #() 
NAND_1261_ (
  .A({ datapath_theregisterfile_memtrf_71 }),
  .B({ S1459 }),
  .Y({ S2284 })
);
NOT #() 
NOT_253_ (
  .A({ S2284 }),
  .Y({ S2285 })
);
NAND #() 
NAND_1262_ (
  .A({ datapath_theregisterfile_memtrf_23 }),
  .B({ S1438 }),
  .Y({ S2286 })
);
NAND #() 
NAND_1263_ (
  .A({ datapath_theregisterfile_memtrf_87 }),
  .B({ S1437 }),
  .Y({ S2287 })
);
NAND #() 
NAND_1264_ (
  .A({ S2286 }),
  .B({ S2287 }),
  .Y({ S2288 })
);
NAND #() 
NAND_1265_ (
  .A({ S1926 }),
  .B({ S2288 }),
  .Y({ S2289 })
);
NAND #() 
NAND_1266_ (
  .A({ S1462 }),
  .B({ S2289 }),
  .Y({ S2290 })
);
NOR #() 
NOR_621_ (
  .A({ S2285 }),
  .B({ S2290 }),
  .Y({ S2291 })
);
NAND #() 
NAND_1267_ (
  .A({ datapath_theregisterfile_memtrf_119 }),
  .B({ S1437 }),
  .Y({ S2292 })
);
NAND #() 
NAND_1268_ (
  .A({ datapath_theregisterfile_memtrf_55 }),
  .B({ S1438 }),
  .Y({ S2293 })
);
NAND #() 
NAND_1269_ (
  .A({ S2292 }),
  .B({ S2293 }),
  .Y({ S2294 })
);
NAND #() 
NAND_1270_ (
  .A({ S1457 }),
  .B({ S2294 }),
  .Y({ S2295 })
);
NAND #() 
NAND_1271_ (
  .A({ datapath_theregisterfile_memtrf_103 }),
  .B({ S1437 }),
  .Y({ S2296 })
);
NAND #() 
NAND_1272_ (
  .A({ datapath_theregisterfile_memtrf_39 }),
  .B({ S1438 }),
  .Y({ S2297 })
);
NAND #() 
NAND_1273_ (
  .A({ S2296 }),
  .B({ S2297 }),
  .Y({ S2298 })
);
NOT #() 
NOT_254_ (
  .A({ S2298 }),
  .Y({ S2299 })
);
NAND #() 
NAND_1274_ (
  .A({ S1458 }),
  .B({ S2298 }),
  .Y({ S2300 })
);
NAND #() 
NAND_1275_ (
  .A({ S2295 }),
  .B({ S2300 }),
  .Y({ S2301 })
);
NOR #() 
NOR_622_ (
  .A({ S1458 }),
  .B({ S2294 }),
  .Y({ S2302 })
);
NAND #() 
NAND_1276_ (
  .A({ S1458 }),
  .B({ S2299 }),
  .Y({ S2303 })
);
NAND #() 
NAND_1277_ (
  .A({ S1487 }),
  .B({ S2303 }),
  .Y({ S2304 })
);
NOR #() 
NOR_623_ (
  .A({ S2302 }),
  .B({ S2304 }),
  .Y({ S2305 })
);
NAND #() 
NAND_1278_ (
  .A({ S1487 }),
  .B({ S2301 }),
  .Y({ S2306 })
);
NAND #() 
NAND_1279_ (
  .A({ S2291 }),
  .B({ S2306 }),
  .Y({ S2307 })
);
NOR #() 
NOR_624_ (
  .A({ S2283 }),
  .B({ S2305 }),
  .Y({ S2308 })
);
NOR #() 
NOR_625_ (
  .A({ S2283 }),
  .B({ S2307 }),
  .Y({ S2309 })
);
NAND #() 
NAND_1280_ (
  .A({ S2291 }),
  .B({ S2308 }),
  .Y({ S2310 })
);
NOR #() 
NOR_626_ (
  .A({ S2260 }),
  .B({ S2309 }),
  .Y({ S2311 })
);
NAND #() 
NAND_1281_ (
  .A({ S2261 }),
  .B({ S2310 }),
  .Y({ S2312 })
);
NAND #() 
NAND_1282_ (
  .A({ S1429 }),
  .B({ S2311 }),
  .Y({ S2313 })
);
NAND #() 
NAND_1283_ (
  .A({ S2259 }),
  .B({ S2313 }),
  .Y({ S2314 })
);
NOT #() 
NOT_255_ (
  .A({ S2314 }),
  .Y({ S2315 })
);
NOR #() 
NOR_627_ (
  .A({ S858 }),
  .B({ S2314 }),
  .Y({ S2316 })
);
NAND #() 
NAND_1284_ (
  .A({ datapath_addsubunit_in1_7 }),
  .B({ S2315 }),
  .Y({ S2317 })
);
NOR #() 
NOR_628_ (
  .A({ datapath_addsubunit_in1_7 }),
  .B({ S2315 }),
  .Y({ S2318 })
);
NAND #() 
NAND_1285_ (
  .A({ S858 }),
  .B({ S2314 }),
  .Y({ S2319 })
);
NAND #() 
NAND_1286_ (
  .A({ datapath_addsubunit_in1_7 }),
  .B({ S2314 }),
  .Y({ S2320 })
);
NOR #() 
NOR_629_ (
  .A({ datapath_addsubunit_in1_7 }),
  .B({ S2314 }),
  .Y({ S2321 })
);
NOR #() 
NOR_630_ (
  .A({ S2316 }),
  .B({ S2318 }),
  .Y({ S2322 })
);
NOR #() 
NOR_631_ (
  .A({ S2225 }),
  .B({ S2228 }),
  .Y({ S2323 })
);
NOR #() 
NOR_632_ (
  .A({ S2212 }),
  .B({ S2219 }),
  .Y({ S2324 })
);
NOR #() 
NOR_633_ (
  .A({ S1533 }),
  .B({ S2320 }),
  .Y({ S2325 })
);
NAND #() 
NAND_1287_ (
  .A({ S1546 }),
  .B({ S2258 }),
  .Y({ S2326 })
);
NAND #() 
NAND_1288_ (
  .A({ datapath_shiftunit_2261_A }),
  .B({ S1614 }),
  .Y({ S2327 })
);
NAND #() 
NAND_1289_ (
  .A({ datapath_shiftunit_2565_A }),
  .B({ S1609 }),
  .Y({ S2328 })
);
NOT #() 
NOT_256_ (
  .A({ S2328 }),
  .Y({ S2329 })
);
NAND #() 
NAND_1290_ (
  .A({ S7936 }),
  .B({ S1346 }),
  .Y({ S2330 })
);
NAND #() 
NAND_1291_ (
  .A({ S1347 }),
  .B({ S2330 }),
  .Y({ S2331 })
);
NOR #() 
NOR_634_ (
  .A({ S1623 }),
  .B({ S2331 }),
  .Y({ S2332 })
);
NAND #() 
NAND_1292_ (
  .A({ datapath_multdivunit_outmdu1_7 }),
  .B({ S1377 }),
  .Y({ S2333 })
);
NAND #() 
NAND_1293_ (
  .A({ datapath_multdivunit_outmdu2_7 }),
  .B({ S8570 }),
  .Y({ S2334 })
);
NAND #() 
NAND_1294_ (
  .A({ datapath_databusin_7 }),
  .B({ S1627 }),
  .Y({ S2335 })
);
NAND #() 
NAND_1295_ (
  .A({ S2333 }),
  .B({ S2335 }),
  .Y({ S2336 })
);
NOR #() 
NOR_635_ (
  .A({ S2332 }),
  .B({ S2336 }),
  .Y({ S2337 })
);
NAND #() 
NAND_1296_ (
  .A({ S2334 }),
  .B({ S2337 }),
  .Y({ S2338 })
);
NOR #() 
NOR_636_ (
  .A({ S2329 }),
  .B({ S2338 }),
  .Y({ S2339 })
);
NOR #() 
NOR_637_ (
  .A({ S858 }),
  .B({ S2248 }),
  .Y({ S2340 })
);
NAND #() 
NAND_1297_ (
  .A({ S858 }),
  .B({ S2248 }),
  .Y({ S2341 })
);
NAND #() 
NAND_1298_ (
  .A({ S2326 }),
  .B({ S2339 }),
  .Y({ S2342 })
);
NOR #() 
NOR_638_ (
  .A({ S2325 }),
  .B({ S2342 }),
  .Y({ S2343 })
);
NOR #() 
NOR_639_ (
  .A({ S1539 }),
  .B({ S2340 }),
  .Y({ S2344 })
);
NAND #() 
NAND_1299_ (
  .A({ S2341 }),
  .B({ S2344 }),
  .Y({ S2345 })
);
NAND #() 
NAND_1300_ (
  .A({ S2327 }),
  .B({ S2345 }),
  .Y({ S2346 })
);
NOT #() 
NOT_257_ (
  .A({ S2346 }),
  .Y({ S2347 })
);
NAND #() 
NAND_1301_ (
  .A({ S2343 }),
  .B({ S2347 }),
  .Y({ S2348 })
);
NOR #() 
NOR_640_ (
  .A({ S2322 }),
  .B({ S2324 }),
  .Y({ S2349 })
);
NOT #() 
NOT_258_ (
  .A({ S2349 }),
  .Y({ S2350 })
);
NAND #() 
NAND_1302_ (
  .A({ S2322 }),
  .B({ S2324 }),
  .Y({ S2351 })
);
NAND #() 
NAND_1303_ (
  .A({ S2350 }),
  .B({ S2351 }),
  .Y({ S2352 })
);
NAND #() 
NAND_1304_ (
  .A({ S1525 }),
  .B({ S2352 }),
  .Y({ S2353 })
);
NOR #() 
NOR_641_ (
  .A({ S2322 }),
  .B({ S2323 }),
  .Y({ S2354 })
);
NAND #() 
NAND_1305_ (
  .A({ S2322 }),
  .B({ S2323 }),
  .Y({ S2355 })
);
NAND #() 
NAND_1306_ (
  .A({ S1527 }),
  .B({ S2355 }),
  .Y({ S2356 })
);
NOR #() 
NOR_642_ (
  .A({ S2354 }),
  .B({ S2356 }),
  .Y({ S2357 })
);
NOR #() 
NOR_643_ (
  .A({ S2348 }),
  .B({ S2357 }),
  .Y({ S2358 })
);
NAND #() 
NAND_1307_ (
  .A({ S2353 }),
  .B({ S2358 }),
  .Y({ datapath_indatatrf_7 })
);
NAND #() 
NAND_1308_ (
  .A({ datapath_indatatrf_7 }),
  .B({ S1688 }),
  .Y({ S2359 })
);
NAND #() 
NAND_1309_ (
  .A({ datapath_theregisterfile_memtrf_71 }),
  .B({ S1689 }),
  .Y({ S2360 })
);
NAND #() 
NAND_1310_ (
  .A({ S2359 }),
  .B({ S2360 }),
  .Y({ S11 })
);
NOR #() 
NOR_644_ (
  .A({ controller_fib_0 }),
  .B({ S1396 }),
  .Y({ S2361 })
);
NOR #() 
NOR_645_ (
  .A({ S1388 }),
  .B({ S1396 }),
  .Y({ S2362 })
);
NOR #() 
NOR_646_ (
  .A({ S8309 }),
  .B({ S2362 }),
  .Y({ S2363 })
);
NOR #() 
NOR_647_ (
  .A({ S1388 }),
  .B({ S2363 }),
  .Y({ S2364 })
);
NOR #() 
NOR_648_ (
  .A({ S2361 }),
  .B({ S2364 }),
  .Y({ S2365 })
);
NOR #() 
NOR_649_ (
  .A({ S2053 }),
  .B({ S2365 }),
  .Y({ S2366 })
);
NOT #() 
NOT_259_ (
  .A({ S2366 }),
  .Y({ S2367 })
);
NOR #() 
NOR_650_ (
  .A({ S1416 }),
  .B({ S2366 }),
  .Y({ S2368 })
);
NAND #() 
NAND_1311_ (
  .A({ S1417 }),
  .B({ S2367 }),
  .Y({ S2369 })
);
NAND #() 
NAND_1312_ (
  .A({ datapath_theregisterfile_memtrf_248 }),
  .B({ S1437 }),
  .Y({ S2370 })
);
NAND #() 
NAND_1313_ (
  .A({ datapath_theregisterfile_memtrf_184 }),
  .B({ S1438 }),
  .Y({ S2371 })
);
NAND #() 
NAND_1314_ (
  .A({ S2370 }),
  .B({ S2371 }),
  .Y({ S2372 })
);
NAND #() 
NAND_1315_ (
  .A({ S1457 }),
  .B({ S2372 }),
  .Y({ S2373 })
);
NAND #() 
NAND_1316_ (
  .A({ datapath_theregisterfile_memtrf_168 }),
  .B({ S1438 }),
  .Y({ S2374 })
);
NAND #() 
NAND_1317_ (
  .A({ datapath_theregisterfile_memtrf_232 }),
  .B({ S1437 }),
  .Y({ S2375 })
);
NAND #() 
NAND_1318_ (
  .A({ S2374 }),
  .B({ S2375 }),
  .Y({ S2376 })
);
NAND #() 
NAND_1319_ (
  .A({ S1458 }),
  .B({ S2376 }),
  .Y({ S2377 })
);
NAND #() 
NAND_1320_ (
  .A({ S2373 }),
  .B({ S2377 }),
  .Y({ S2378 })
);
NAND #() 
NAND_1321_ (
  .A({ datapath_theregisterfile_memtrf_152 }),
  .B({ S1438 }),
  .Y({ S2379 })
);
NAND #() 
NAND_1322_ (
  .A({ datapath_theregisterfile_memtrf_216 }),
  .B({ S1437 }),
  .Y({ S2380 })
);
NAND #() 
NAND_1323_ (
  .A({ S2379 }),
  .B({ S2380 }),
  .Y({ S2381 })
);
NAND #() 
NAND_1324_ (
  .A({ S1457 }),
  .B({ S2381 }),
  .Y({ S2382 })
);
NOR #() 
NOR_651_ (
  .A({ datapath_theregisterfile_memtrf_136 }),
  .B({ S1437 }),
  .Y({ S2383 })
);
NAND #() 
NAND_1325_ (
  .A({ S7739 }),
  .B({ S1437 }),
  .Y({ S2384 })
);
NAND #() 
NAND_1326_ (
  .A({ S1458 }),
  .B({ S2384 }),
  .Y({ S2385 })
);
NOR #() 
NOR_652_ (
  .A({ S2383 }),
  .B({ S2385 }),
  .Y({ S2386 })
);
NOR #() 
NOR_653_ (
  .A({ S1444 }),
  .B({ S2378 }),
  .Y({ S2387 })
);
NOR #() 
NOR_654_ (
  .A({ S1443 }),
  .B({ S2386 }),
  .Y({ S2388 })
);
NAND #() 
NAND_1327_ (
  .A({ S2382 }),
  .B({ S2388 }),
  .Y({ S2389 })
);
NAND #() 
NAND_1328_ (
  .A({ S1449 }),
  .B({ S2389 }),
  .Y({ S2390 })
);
NOR #() 
NOR_655_ (
  .A({ S2387 }),
  .B({ S2390 }),
  .Y({ S2391 })
);
NAND #() 
NAND_1329_ (
  .A({ datapath_theregisterfile_memtrf_104 }),
  .B({ S1458 }),
  .Y({ S2392 })
);
NAND #() 
NAND_1330_ (
  .A({ datapath_theregisterfile_memtrf_120 }),
  .B({ S1457 }),
  .Y({ S2393 })
);
NAND #() 
NAND_1331_ (
  .A({ S2392 }),
  .B({ S2393 }),
  .Y({ S2394 })
);
NAND #() 
NAND_1332_ (
  .A({ S1437 }),
  .B({ S2394 }),
  .Y({ S2395 })
);
NAND #() 
NAND_1333_ (
  .A({ datapath_theregisterfile_memtrf_40 }),
  .B({ S1458 }),
  .Y({ S2396 })
);
NAND #() 
NAND_1334_ (
  .A({ datapath_theregisterfile_memtrf_56 }),
  .B({ S1457 }),
  .Y({ S2397 })
);
NAND #() 
NAND_1335_ (
  .A({ S2396 }),
  .B({ S2397 }),
  .Y({ S2398 })
);
NAND #() 
NAND_1336_ (
  .A({ S1438 }),
  .B({ S2398 }),
  .Y({ S2399 })
);
NAND #() 
NAND_1337_ (
  .A({ S2395 }),
  .B({ S2399 }),
  .Y({ S2400 })
);
NAND #() 
NAND_1338_ (
  .A({ S1487 }),
  .B({ S2400 }),
  .Y({ S2401 })
);
NOR #() 
NOR_656_ (
  .A({ datapath_theregisterfile_memtrf_72 }),
  .B({ S1438 }),
  .Y({ S2402 })
);
NOR #() 
NOR_657_ (
  .A({ datapath_theregisterfile_memtrf_8 }),
  .B({ S1437 }),
  .Y({ S2403 })
);
NOR #() 
NOR_658_ (
  .A({ S2402 }),
  .B({ S2403 }),
  .Y({ S2404 })
);
NAND #() 
NAND_1339_ (
  .A({ S1459 }),
  .B({ S2404 }),
  .Y({ S2405 })
);
NAND #() 
NAND_1340_ (
  .A({ datapath_theregisterfile_memtrf_24 }),
  .B({ S1438 }),
  .Y({ S2406 })
);
NAND #() 
NAND_1341_ (
  .A({ datapath_theregisterfile_memtrf_88 }),
  .B({ S1437 }),
  .Y({ S2407 })
);
NAND #() 
NAND_1342_ (
  .A({ S2406 }),
  .B({ S2407 }),
  .Y({ S2408 })
);
NAND #() 
NAND_1343_ (
  .A({ S1926 }),
  .B({ S2408 }),
  .Y({ S2409 })
);
NAND #() 
NAND_1344_ (
  .A({ S2405 }),
  .B({ S2409 }),
  .Y({ S2410 })
);
NOT #() 
NOT_260_ (
  .A({ S2410 }),
  .Y({ S2411 })
);
NAND #() 
NAND_1345_ (
  .A({ S2401 }),
  .B({ S2411 }),
  .Y({ S2412 })
);
NAND #() 
NAND_1346_ (
  .A({ S2401 }),
  .B({ S2409 }),
  .Y({ S2413 })
);
NOR #() 
NOR_659_ (
  .A({ S2391 }),
  .B({ S2413 }),
  .Y({ S2414 })
);
NOR #() 
NOR_660_ (
  .A({ S2391 }),
  .B({ S2412 }),
  .Y({ S2415 })
);
NAND #() 
NAND_1347_ (
  .A({ S2405 }),
  .B({ S2414 }),
  .Y({ S2416 })
);
NOR #() 
NOR_661_ (
  .A({ S1461 }),
  .B({ S2415 }),
  .Y({ S2417 })
);
NAND #() 
NAND_1348_ (
  .A({ S1462 }),
  .B({ S2416 }),
  .Y({ S2418 })
);
NOR #() 
NOR_662_ (
  .A({ S1430 }),
  .B({ S2418 }),
  .Y({ S2419 })
);
NOR #() 
NOR_663_ (
  .A({ S2368 }),
  .B({ S2419 }),
  .Y({ S2420 })
);
NAND #() 
NAND_1349_ (
  .A({ datapath_addsubunit_in1_8 }),
  .B({ S2420 }),
  .Y({ S2421 })
);
NOR #() 
NOR_664_ (
  .A({ datapath_addsubunit_in1_8 }),
  .B({ S2420 }),
  .Y({ S2422 })
);
NOT #() 
NOT_261_ (
  .A({ S2422 }),
  .Y({ S2423 })
);
NAND #() 
NAND_1350_ (
  .A({ S2421 }),
  .B({ S2423 }),
  .Y({ S2424 })
);
NOT #() 
NOT_262_ (
  .A({ S2424 }),
  .Y({ S2425 })
);
NOR #() 
NOR_665_ (
  .A({ S2321 }),
  .B({ S2323 }),
  .Y({ S2426 })
);
NOT #() 
NOT_263_ (
  .A({ S2426 }),
  .Y({ S2427 })
);
NAND #() 
NAND_1351_ (
  .A({ S2320 }),
  .B({ S2427 }),
  .Y({ S2428 })
);
NOT #() 
NOT_264_ (
  .A({ S2428 }),
  .Y({ S2429 })
);
NOR #() 
NOR_666_ (
  .A({ S2424 }),
  .B({ S2428 }),
  .Y({ S2430 })
);
NOR #() 
NOR_667_ (
  .A({ S2425 }),
  .B({ S2429 }),
  .Y({ S2431 })
);
NOR #() 
NOR_668_ (
  .A({ S2430 }),
  .B({ S2431 }),
  .Y({ S2432 })
);
NAND #() 
NAND_1352_ (
  .A({ S1527 }),
  .B({ S2432 }),
  .Y({ S2433 })
);
NOR #() 
NOR_669_ (
  .A({ S2318 }),
  .B({ S2324 }),
  .Y({ S2434 })
);
NAND #() 
NAND_1353_ (
  .A({ S2213 }),
  .B({ S2322 }),
  .Y({ S2435 })
);
NOR #() 
NOR_670_ (
  .A({ S2316 }),
  .B({ S2434 }),
  .Y({ S2436 })
);
NOR #() 
NOR_671_ (
  .A({ S2424 }),
  .B({ S2436 }),
  .Y({ S2437 })
);
NOT #() 
NOT_265_ (
  .A({ S2437 }),
  .Y({ S2438 })
);
NAND #() 
NAND_1354_ (
  .A({ S2424 }),
  .B({ S2436 }),
  .Y({ S2439 })
);
NAND #() 
NAND_1355_ (
  .A({ S1525 }),
  .B({ S2439 }),
  .Y({ S2440 })
);
NOR #() 
NOR_672_ (
  .A({ S2437 }),
  .B({ S2440 }),
  .Y({ S2441 })
);
NOR #() 
NOR_673_ (
  .A({ S805 }),
  .B({ S2420 }),
  .Y({ S2442 })
);
NOT #() 
NOT_266_ (
  .A({ S2442 }),
  .Y({ S2443 })
);
NOR #() 
NOR_674_ (
  .A({ S1533 }),
  .B({ S2443 }),
  .Y({ S2444 })
);
NAND #() 
NAND_1356_ (
  .A({ datapath_shiftunit_2279_A }),
  .B({ S1614 }),
  .Y({ S2445 })
);
NAND #() 
NAND_1357_ (
  .A({ datapath_shiftunit_2583_A }),
  .B({ S1609 }),
  .Y({ S2446 })
);
NOR #() 
NOR_675_ (
  .A({ S1547 }),
  .B({ S2366 }),
  .Y({ S2447 })
);
NAND #() 
NAND_1358_ (
  .A({ S7946 }),
  .B({ S1347 }),
  .Y({ S2448 })
);
NAND #() 
NAND_1359_ (
  .A({ S1350 }),
  .B({ S2448 }),
  .Y({ S2449 })
);
NOR #() 
NOR_676_ (
  .A({ S1623 }),
  .B({ S2449 }),
  .Y({ S2450 })
);
NAND #() 
NAND_1360_ (
  .A({ datapath_databusin_8 }),
  .B({ S1627 }),
  .Y({ S2451 })
);
NAND #() 
NAND_1361_ (
  .A({ datapath_multdivunit_outmdu1_8 }),
  .B({ S1377 }),
  .Y({ S2452 })
);
NAND #() 
NAND_1362_ (
  .A({ datapath_multdivunit_outmdu2_8 }),
  .B({ S8570 }),
  .Y({ S2453 })
);
NAND #() 
NAND_1363_ (
  .A({ S2451 }),
  .B({ S2452 }),
  .Y({ S2454 })
);
NOR #() 
NOR_677_ (
  .A({ S2447 }),
  .B({ S2454 }),
  .Y({ S2455 })
);
NAND #() 
NAND_1364_ (
  .A({ S2453 }),
  .B({ S2455 }),
  .Y({ S2456 })
);
NOR #() 
NOR_678_ (
  .A({ S2450 }),
  .B({ S2456 }),
  .Y({ S2457 })
);
NAND #() 
NAND_1365_ (
  .A({ S2445 }),
  .B({ S2457 }),
  .Y({ S2458 })
);
NOT #() 
NOT_267_ (
  .A({ S2458 }),
  .Y({ S2459 })
);
NAND #() 
NAND_1366_ (
  .A({ S2446 }),
  .B({ S2459 }),
  .Y({ S2460 })
);
NOR #() 
NOR_679_ (
  .A({ S2444 }),
  .B({ S2460 }),
  .Y({ S2461 })
);
NAND #() 
NAND_1367_ (
  .A({ datapath_addsubunit_in1_8 }),
  .B({ S2341 }),
  .Y({ S2462 })
);
NOR #() 
NOR_680_ (
  .A({ datapath_addsubunit_in1_8 }),
  .B({ S2341 }),
  .Y({ S2463 })
);
NOT #() 
NOT_268_ (
  .A({ S2463 }),
  .Y({ S2464 })
);
NOR #() 
NOR_681_ (
  .A({ S1539 }),
  .B({ S2463 }),
  .Y({ S2465 })
);
NAND #() 
NAND_1368_ (
  .A({ S2462 }),
  .B({ S2465 }),
  .Y({ S2466 })
);
NAND #() 
NAND_1369_ (
  .A({ S2461 }),
  .B({ S2466 }),
  .Y({ S2467 })
);
NOR #() 
NOR_682_ (
  .A({ S2441 }),
  .B({ S2467 }),
  .Y({ S2468 })
);
NAND #() 
NAND_1370_ (
  .A({ S2433 }),
  .B({ S2468 }),
  .Y({ datapath_indatatrf_8 })
);
NAND #() 
NAND_1371_ (
  .A({ datapath_indatatrf_8 }),
  .B({ S1688 }),
  .Y({ S2469 })
);
NAND #() 
NAND_1372_ (
  .A({ datapath_theregisterfile_memtrf_72 }),
  .B({ S1689 }),
  .Y({ S2470 })
);
NAND #() 
NAND_1373_ (
  .A({ S2469 }),
  .B({ S2470 }),
  .Y({ S12 })
);
NAND #() 
NAND_1374_ (
  .A({ datapath_theregisterfile_memtrf_249 }),
  .B({ S1437 }),
  .Y({ S2471 })
);
NAND #() 
NAND_1375_ (
  .A({ datapath_theregisterfile_memtrf_185 }),
  .B({ S1438 }),
  .Y({ S2472 })
);
NAND #() 
NAND_1376_ (
  .A({ S2471 }),
  .B({ S2472 }),
  .Y({ S2473 })
);
NAND #() 
NAND_1377_ (
  .A({ S1457 }),
  .B({ S2473 }),
  .Y({ S2474 })
);
NAND #() 
NAND_1378_ (
  .A({ datapath_theregisterfile_memtrf_169 }),
  .B({ S1438 }),
  .Y({ S2475 })
);
NAND #() 
NAND_1379_ (
  .A({ datapath_theregisterfile_memtrf_233 }),
  .B({ S1437 }),
  .Y({ S2476 })
);
NAND #() 
NAND_1380_ (
  .A({ S2475 }),
  .B({ S2476 }),
  .Y({ S2477 })
);
NAND #() 
NAND_1381_ (
  .A({ S1458 }),
  .B({ S2477 }),
  .Y({ S2478 })
);
NAND #() 
NAND_1382_ (
  .A({ S2474 }),
  .B({ S2478 }),
  .Y({ S2479 })
);
NAND #() 
NAND_1383_ (
  .A({ S1443 }),
  .B({ S2479 }),
  .Y({ S2480 })
);
NAND #() 
NAND_1384_ (
  .A({ datapath_theregisterfile_memtrf_153 }),
  .B({ S1438 }),
  .Y({ S2481 })
);
NAND #() 
NAND_1385_ (
  .A({ datapath_theregisterfile_memtrf_217 }),
  .B({ S1437 }),
  .Y({ S2482 })
);
NAND #() 
NAND_1386_ (
  .A({ S2481 }),
  .B({ S2482 }),
  .Y({ S2483 })
);
NAND #() 
NAND_1387_ (
  .A({ S1457 }),
  .B({ S2483 }),
  .Y({ S2484 })
);
NOR #() 
NOR_683_ (
  .A({ datapath_theregisterfile_memtrf_137 }),
  .B({ S1437 }),
  .Y({ S2485 })
);
NOR #() 
NOR_684_ (
  .A({ datapath_theregisterfile_memtrf_201 }),
  .B({ S1438 }),
  .Y({ S2486 })
);
NOR #() 
NOR_685_ (
  .A({ S2485 }),
  .B({ S2486 }),
  .Y({ S2487 })
);
NAND #() 
NAND_1388_ (
  .A({ S1458 }),
  .B({ S2487 }),
  .Y({ S2488 })
);
NAND #() 
NAND_1389_ (
  .A({ S2484 }),
  .B({ S2488 }),
  .Y({ S2489 })
);
NAND #() 
NAND_1390_ (
  .A({ S1444 }),
  .B({ S2489 }),
  .Y({ S2490 })
);
NAND #() 
NAND_1391_ (
  .A({ S2480 }),
  .B({ S2490 }),
  .Y({ S2491 })
);
NAND #() 
NAND_1392_ (
  .A({ S1449 }),
  .B({ S2491 }),
  .Y({ S2492 })
);
NAND #() 
NAND_1393_ (
  .A({ datapath_theregisterfile_memtrf_25 }),
  .B({ S1438 }),
  .Y({ S2493 })
);
NAND #() 
NAND_1394_ (
  .A({ datapath_theregisterfile_memtrf_89 }),
  .B({ S1437 }),
  .Y({ S2494 })
);
NAND #() 
NAND_1395_ (
  .A({ S2493 }),
  .B({ S2494 }),
  .Y({ S2495 })
);
NAND #() 
NAND_1396_ (
  .A({ S1926 }),
  .B({ S2495 }),
  .Y({ S2496 })
);
NAND #() 
NAND_1397_ (
  .A({ datapath_theregisterfile_memtrf_9 }),
  .B({ S1438 }),
  .Y({ S2497 })
);
NAND #() 
NAND_1398_ (
  .A({ datapath_theregisterfile_memtrf_73 }),
  .B({ S1437 }),
  .Y({ S2498 })
);
NAND #() 
NAND_1399_ (
  .A({ S2497 }),
  .B({ S2498 }),
  .Y({ S2499 })
);
NAND #() 
NAND_1400_ (
  .A({ S1459 }),
  .B({ S2499 }),
  .Y({ S2500 })
);
NAND #() 
NAND_1401_ (
  .A({ S2496 }),
  .B({ S2500 }),
  .Y({ S2501 })
);
NAND #() 
NAND_1402_ (
  .A({ datapath_theregisterfile_memtrf_57 }),
  .B({ S1438 }),
  .Y({ S2502 })
);
NAND #() 
NAND_1403_ (
  .A({ datapath_theregisterfile_memtrf_121 }),
  .B({ S1437 }),
  .Y({ S2503 })
);
NAND #() 
NAND_1404_ (
  .A({ S2502 }),
  .B({ S2503 }),
  .Y({ S2504 })
);
NOR #() 
NOR_686_ (
  .A({ S1458 }),
  .B({ S2504 }),
  .Y({ S2505 })
);
NOR #() 
NOR_687_ (
  .A({ datapath_theregisterfile_memtrf_41 }),
  .B({ S1437 }),
  .Y({ S2506 })
);
NOR #() 
NOR_688_ (
  .A({ datapath_theregisterfile_memtrf_105 }),
  .B({ S1438 }),
  .Y({ S2507 })
);
NOR #() 
NOR_689_ (
  .A({ S2506 }),
  .B({ S2507 }),
  .Y({ S2508 })
);
NOR #() 
NOR_690_ (
  .A({ S1457 }),
  .B({ S2508 }),
  .Y({ S2509 })
);
NOR #() 
NOR_691_ (
  .A({ S2505 }),
  .B({ S2509 }),
  .Y({ S2510 })
);
NAND #() 
NAND_1405_ (
  .A({ S1487 }),
  .B({ S2510 }),
  .Y({ S2511 })
);
NOT #() 
NOT_269_ (
  .A({ S2511 }),
  .Y({ S2512 })
);
NOR #() 
NOR_692_ (
  .A({ S2501 }),
  .B({ S2512 }),
  .Y({ S2513 })
);
NAND #() 
NAND_1406_ (
  .A({ S2492 }),
  .B({ S2511 }),
  .Y({ S2514 })
);
NOR #() 
NOR_693_ (
  .A({ S2501 }),
  .B({ S2514 }),
  .Y({ S2515 })
);
NAND #() 
NAND_1407_ (
  .A({ S2492 }),
  .B({ S2513 }),
  .Y({ S2516 })
);
NOR #() 
NOR_694_ (
  .A({ S1461 }),
  .B({ S2515 }),
  .Y({ S2517 })
);
NAND #() 
NAND_1408_ (
  .A({ S1462 }),
  .B({ S2516 }),
  .Y({ S2518 })
);
NOR #() 
NOR_695_ (
  .A({ S1430 }),
  .B({ S2518 }),
  .Y({ S2519 })
);
NAND #() 
NAND_1409_ (
  .A({ S1429 }),
  .B({ S2517 }),
  .Y({ S2520 })
);
NOR #() 
NOR_696_ (
  .A({ S2368 }),
  .B({ S2519 }),
  .Y({ S2521 })
);
NAND #() 
NAND_1410_ (
  .A({ S2369 }),
  .B({ S2520 }),
  .Y({ S2522 })
);
NOR #() 
NOR_697_ (
  .A({ S754 }),
  .B({ S2522 }),
  .Y({ S2523 })
);
NOR #() 
NOR_698_ (
  .A({ datapath_addsubunit_in1_9 }),
  .B({ S2521 }),
  .Y({ S2524 })
);
NOR #() 
NOR_699_ (
  .A({ S2523 }),
  .B({ S2524 }),
  .Y({ S2525 })
);
NOT #() 
NOT_270_ (
  .A({ S2525 }),
  .Y({ S2526 })
);
NAND #() 
NAND_1411_ (
  .A({ S2421 }),
  .B({ S2438 }),
  .Y({ S2527 })
);
NOR #() 
NOR_700_ (
  .A({ S2525 }),
  .B({ S2527 }),
  .Y({ S2528 })
);
NAND #() 
NAND_1412_ (
  .A({ S2525 }),
  .B({ S2527 }),
  .Y({ S2529 })
);
NOR #() 
NOR_701_ (
  .A({ S1526 }),
  .B({ S2528 }),
  .Y({ S2530 })
);
NAND #() 
NAND_1413_ (
  .A({ S2529 }),
  .B({ S2530 }),
  .Y({ S2531 })
);
NAND #() 
NAND_1414_ (
  .A({ S2431 }),
  .B({ S2526 }),
  .Y({ S2532 })
);
NOR #() 
NOR_702_ (
  .A({ S2431 }),
  .B({ S2442 }),
  .Y({ S2533 })
);
NAND #() 
NAND_1415_ (
  .A({ S2525 }),
  .B({ S2533 }),
  .Y({ S2534 })
);
NOR #() 
NOR_703_ (
  .A({ S2443 }),
  .B({ S2525 }),
  .Y({ S2535 })
);
NOR #() 
NOR_704_ (
  .A({ S2525 }),
  .B({ S2533 }),
  .Y({ S2536 })
);
NOR #() 
NOR_705_ (
  .A({ S1528 }),
  .B({ S2536 }),
  .Y({ S2537 })
);
NAND #() 
NAND_1416_ (
  .A({ S2534 }),
  .B({ S2537 }),
  .Y({ S2538 })
);
NAND #() 
NAND_1417_ (
  .A({ datapath_addsubunit_in1_9 }),
  .B({ S2464 }),
  .Y({ S2539 })
);
NAND #() 
NAND_1418_ (
  .A({ S754 }),
  .B({ S2463 }),
  .Y({ S2540 })
);
NOT #() 
NOT_271_ (
  .A({ S2540 }),
  .Y({ S2541 })
);
NAND #() 
NAND_1419_ (
  .A({ datapath_shiftunit_2297_A }),
  .B({ S1614 }),
  .Y({ S2542 })
);
NAND #() 
NAND_1420_ (
  .A({ datapath_shiftunit_2601_A }),
  .B({ S1609 }),
  .Y({ S2543 })
);
NOT #() 
NOT_272_ (
  .A({ S2543 }),
  .Y({ S2544 })
);
NOR #() 
NOR_706_ (
  .A({ controller_fib_1 }),
  .B({ S1396 }),
  .Y({ S2545 })
);
NOR #() 
NOR_707_ (
  .A({ S2364 }),
  .B({ S2545 }),
  .Y({ S2546 })
);
NOR #() 
NOR_708_ (
  .A({ S2053 }),
  .B({ S2546 }),
  .Y({ S2547 })
);
NOR #() 
NOR_709_ (
  .A({ S1547 }),
  .B({ S2547 }),
  .Y({ S2548 })
);
NOT #() 
NOT_273_ (
  .A({ S2548 }),
  .Y({ S2549 })
);
NAND #() 
NAND_1421_ (
  .A({ S7957 }),
  .B({ S1350 }),
  .Y({ S2550 })
);
NAND #() 
NAND_1422_ (
  .A({ S1352 }),
  .B({ S2550 }),
  .Y({ S2551 })
);
NOR #() 
NOR_710_ (
  .A({ S1623 }),
  .B({ S2551 }),
  .Y({ S2552 })
);
NOR #() 
NOR_711_ (
  .A({ S8129 }),
  .B({ S8571 }),
  .Y({ S2553 })
);
NAND #() 
NAND_1423_ (
  .A({ datapath_multdivunit_outmdu1_9 }),
  .B({ S1377 }),
  .Y({ S2554 })
);
NOR #() 
NOR_712_ (
  .A({ S8288 }),
  .B({ S1628 }),
  .Y({ S2555 })
);
NOR #() 
NOR_713_ (
  .A({ S2553 }),
  .B({ S2555 }),
  .Y({ S2556 })
);
NAND #() 
NAND_1424_ (
  .A({ S2549 }),
  .B({ S2556 }),
  .Y({ S2557 })
);
NOR #() 
NOR_714_ (
  .A({ S2552 }),
  .B({ S2557 }),
  .Y({ S2558 })
);
NAND #() 
NAND_1425_ (
  .A({ S2554 }),
  .B({ S2558 }),
  .Y({ S2559 })
);
NOR #() 
NOR_715_ (
  .A({ S2544 }),
  .B({ S2559 }),
  .Y({ S2560 })
);
NAND #() 
NAND_1426_ (
  .A({ S2542 }),
  .B({ S2560 }),
  .Y({ S2561 })
);
NAND #() 
NAND_1427_ (
  .A({ datapath_addsubunit_in1_9 }),
  .B({ S2522 }),
  .Y({ S2562 })
);
NOR #() 
NOR_716_ (
  .A({ S1533 }),
  .B({ S2562 }),
  .Y({ S2563 })
);
NAND #() 
NAND_1428_ (
  .A({ S2539 }),
  .B({ S2540 }),
  .Y({ S2564 })
);
NOR #() 
NOR_717_ (
  .A({ S1539 }),
  .B({ S2564 }),
  .Y({ S2565 })
);
NOR #() 
NOR_718_ (
  .A({ S2563 }),
  .B({ S2565 }),
  .Y({ S2566 })
);
NAND #() 
NAND_1429_ (
  .A({ S2531 }),
  .B({ S2566 }),
  .Y({ S2567 })
);
NOR #() 
NOR_719_ (
  .A({ S2561 }),
  .B({ S2567 }),
  .Y({ S2568 })
);
NAND #() 
NAND_1430_ (
  .A({ S2538 }),
  .B({ S2568 }),
  .Y({ datapath_indatatrf_9 })
);
NAND #() 
NAND_1431_ (
  .A({ datapath_indatatrf_9 }),
  .B({ S1688 }),
  .Y({ S2569 })
);
NAND #() 
NAND_1432_ (
  .A({ datapath_theregisterfile_memtrf_73 }),
  .B({ S1689 }),
  .Y({ S2570 })
);
NAND #() 
NAND_1433_ (
  .A({ S2569 }),
  .B({ S2570 }),
  .Y({ S13 })
);
NAND #() 
NAND_1434_ (
  .A({ datapath_theregisterfile_memtrf_250 }),
  .B({ S1443 }),
  .Y({ S2571 })
);
NAND #() 
NAND_1435_ (
  .A({ datapath_theregisterfile_memtrf_218 }),
  .B({ S1444 }),
  .Y({ S2572 })
);
NAND #() 
NAND_1436_ (
  .A({ S2571 }),
  .B({ S2572 }),
  .Y({ S2573 })
);
NAND #() 
NAND_1437_ (
  .A({ S1437 }),
  .B({ S2573 }),
  .Y({ S2574 })
);
NAND #() 
NAND_1438_ (
  .A({ datapath_theregisterfile_memtrf_186 }),
  .B({ S1443 }),
  .Y({ S2575 })
);
NAND #() 
NAND_1439_ (
  .A({ datapath_theregisterfile_memtrf_154 }),
  .B({ S1444 }),
  .Y({ S2576 })
);
NAND #() 
NAND_1440_ (
  .A({ S2575 }),
  .B({ S2576 }),
  .Y({ S2577 })
);
NAND #() 
NAND_1441_ (
  .A({ S1438 }),
  .B({ S2577 }),
  .Y({ S2578 })
);
NAND #() 
NAND_1442_ (
  .A({ S2574 }),
  .B({ S2578 }),
  .Y({ S2579 })
);
NAND #() 
NAND_1443_ (
  .A({ S1457 }),
  .B({ S2579 }),
  .Y({ S2580 })
);
NAND #() 
NAND_1444_ (
  .A({ datapath_theregisterfile_memtrf_234 }),
  .B({ S1443 }),
  .Y({ S2581 })
);
NAND #() 
NAND_1445_ (
  .A({ datapath_theregisterfile_memtrf_202 }),
  .B({ S1444 }),
  .Y({ S2582 })
);
NAND #() 
NAND_1446_ (
  .A({ S2581 }),
  .B({ S2582 }),
  .Y({ S2583 })
);
NAND #() 
NAND_1447_ (
  .A({ S1437 }),
  .B({ S2583 }),
  .Y({ S2584 })
);
NAND #() 
NAND_1448_ (
  .A({ datapath_theregisterfile_memtrf_170 }),
  .B({ S1443 }),
  .Y({ S2585 })
);
NAND #() 
NAND_1449_ (
  .A({ datapath_theregisterfile_memtrf_138 }),
  .B({ S1444 }),
  .Y({ S2586 })
);
NAND #() 
NAND_1450_ (
  .A({ S2585 }),
  .B({ S2586 }),
  .Y({ S2587 })
);
NAND #() 
NAND_1451_ (
  .A({ S1438 }),
  .B({ S2587 }),
  .Y({ S2588 })
);
NAND #() 
NAND_1452_ (
  .A({ S2584 }),
  .B({ S2588 }),
  .Y({ S2589 })
);
NAND #() 
NAND_1453_ (
  .A({ S1458 }),
  .B({ S2589 }),
  .Y({ S2590 })
);
NAND #() 
NAND_1454_ (
  .A({ S2580 }),
  .B({ S2590 }),
  .Y({ S2591 })
);
NAND #() 
NAND_1455_ (
  .A({ S1449 }),
  .B({ S2591 }),
  .Y({ S2592 })
);
NOR #() 
NOR_720_ (
  .A({ datapath_theregisterfile_memtrf_74 }),
  .B({ S1438 }),
  .Y({ S2593 })
);
NOR #() 
NOR_721_ (
  .A({ datapath_theregisterfile_memtrf_10 }),
  .B({ S1437 }),
  .Y({ S2594 })
);
NOR #() 
NOR_722_ (
  .A({ S2593 }),
  .B({ S2594 }),
  .Y({ S2595 })
);
NAND #() 
NAND_1456_ (
  .A({ S1459 }),
  .B({ S2595 }),
  .Y({ S2596 })
);
NAND #() 
NAND_1457_ (
  .A({ datapath_theregisterfile_memtrf_26 }),
  .B({ S1438 }),
  .Y({ S2597 })
);
NAND #() 
NAND_1458_ (
  .A({ datapath_theregisterfile_memtrf_90 }),
  .B({ S1437 }),
  .Y({ S2598 })
);
NAND #() 
NAND_1459_ (
  .A({ S2597 }),
  .B({ S2598 }),
  .Y({ S2599 })
);
NAND #() 
NAND_1460_ (
  .A({ S1926 }),
  .B({ S2599 }),
  .Y({ S2600 })
);
NAND #() 
NAND_1461_ (
  .A({ S2596 }),
  .B({ S2600 }),
  .Y({ S2601 })
);
NAND #() 
NAND_1462_ (
  .A({ datapath_theregisterfile_memtrf_58 }),
  .B({ S1438 }),
  .Y({ S2602 })
);
NAND #() 
NAND_1463_ (
  .A({ datapath_theregisterfile_memtrf_122 }),
  .B({ S1437 }),
  .Y({ S2603 })
);
NAND #() 
NAND_1464_ (
  .A({ S2602 }),
  .B({ S2603 }),
  .Y({ S2604 })
);
NOR #() 
NOR_723_ (
  .A({ S1458 }),
  .B({ S2604 }),
  .Y({ S2605 })
);
NOR #() 
NOR_724_ (
  .A({ datapath_theregisterfile_memtrf_42 }),
  .B({ S1437 }),
  .Y({ S2606 })
);
NOR #() 
NOR_725_ (
  .A({ datapath_theregisterfile_memtrf_106 }),
  .B({ S1438 }),
  .Y({ S2607 })
);
NOR #() 
NOR_726_ (
  .A({ S2606 }),
  .B({ S2607 }),
  .Y({ S2608 })
);
NOR #() 
NOR_727_ (
  .A({ S1457 }),
  .B({ S2608 }),
  .Y({ S2609 })
);
NOR #() 
NOR_728_ (
  .A({ S2605 }),
  .B({ S2609 }),
  .Y({ S2610 })
);
NAND #() 
NAND_1465_ (
  .A({ S1487 }),
  .B({ S2610 }),
  .Y({ S2611 })
);
NOT #() 
NOT_274_ (
  .A({ S2611 }),
  .Y({ S2612 })
);
NOR #() 
NOR_729_ (
  .A({ S2601 }),
  .B({ S2612 }),
  .Y({ S2613 })
);
NAND #() 
NAND_1466_ (
  .A({ S2592 }),
  .B({ S2611 }),
  .Y({ S2614 })
);
NOR #() 
NOR_730_ (
  .A({ S2601 }),
  .B({ S2614 }),
  .Y({ S2615 })
);
NAND #() 
NAND_1467_ (
  .A({ S2592 }),
  .B({ S2613 }),
  .Y({ S2616 })
);
NOR #() 
NOR_731_ (
  .A({ S1461 }),
  .B({ S2615 }),
  .Y({ S2617 })
);
NAND #() 
NAND_1468_ (
  .A({ S1462 }),
  .B({ S2616 }),
  .Y({ S2618 })
);
NAND #() 
NAND_1469_ (
  .A({ S1429 }),
  .B({ S2617 }),
  .Y({ S2619 })
);
NAND #() 
NAND_1470_ (
  .A({ S2369 }),
  .B({ S2619 }),
  .Y({ S2620 })
);
NOT #() 
NOT_275_ (
  .A({ S2620 }),
  .Y({ S2621 })
);
NAND #() 
NAND_1471_ (
  .A({ S702 }),
  .B({ S2620 }),
  .Y({ S2622 })
);
NOT #() 
NOT_276_ (
  .A({ S2622 }),
  .Y({ S2623 })
);
NAND #() 
NAND_1472_ (
  .A({ datapath_addsubunit_in1_10 }),
  .B({ S2621 }),
  .Y({ S2624 })
);
NOT #() 
NOT_277_ (
  .A({ S2624 }),
  .Y({ S2625 })
);
NOR #() 
NOR_732_ (
  .A({ S2623 }),
  .B({ S2625 }),
  .Y({ S2626 })
);
NOR #() 
NOR_733_ (
  .A({ S2523 }),
  .B({ S2527 }),
  .Y({ S2627 })
);
NOR #() 
NOR_734_ (
  .A({ S2524 }),
  .B({ S2627 }),
  .Y({ S2628 })
);
NOR #() 
NOR_735_ (
  .A({ S2626 }),
  .B({ S2628 }),
  .Y({ S2629 })
);
NAND #() 
NAND_1473_ (
  .A({ S2626 }),
  .B({ S2628 }),
  .Y({ S2630 })
);
NOR #() 
NOR_736_ (
  .A({ S1526 }),
  .B({ S2629 }),
  .Y({ S2631 })
);
NAND #() 
NAND_1474_ (
  .A({ S2630 }),
  .B({ S2631 }),
  .Y({ S2632 })
);
NAND #() 
NAND_1475_ (
  .A({ S2532 }),
  .B({ S2562 }),
  .Y({ S2633 })
);
NOR #() 
NOR_737_ (
  .A({ S2535 }),
  .B({ S2633 }),
  .Y({ S2634 })
);
NOR #() 
NOR_738_ (
  .A({ S2626 }),
  .B({ S2634 }),
  .Y({ S2635 })
);
NAND #() 
NAND_1476_ (
  .A({ S2626 }),
  .B({ S2634 }),
  .Y({ S2636 })
);
NAND #() 
NAND_1477_ (
  .A({ S1527 }),
  .B({ S2636 }),
  .Y({ S2637 })
);
NOR #() 
NOR_739_ (
  .A({ S2635 }),
  .B({ S2637 }),
  .Y({ S2638 })
);
NAND #() 
NAND_1478_ (
  .A({ datapath_addsubunit_in1_10 }),
  .B({ S2620 }),
  .Y({ S2639 })
);
NOT #() 
NOT_278_ (
  .A({ S2639 }),
  .Y({ S2640 })
);
NOR #() 
NOR_740_ (
  .A({ S1533 }),
  .B({ S2639 }),
  .Y({ S2641 })
);
NAND #() 
NAND_1479_ (
  .A({ datapath_shiftunit_2315_A }),
  .B({ S1614 }),
  .Y({ S2642 })
);
NAND #() 
NAND_1480_ (
  .A({ datapath_shiftunit_2619_A }),
  .B({ S1609 }),
  .Y({ S2643 })
);
NOT #() 
NOT_279_ (
  .A({ S2643 }),
  .Y({ S2644 })
);
NAND #() 
NAND_1481_ (
  .A({ S7968 }),
  .B({ S1352 }),
  .Y({ S2645 })
);
NAND #() 
NAND_1482_ (
  .A({ S1354 }),
  .B({ S2645 }),
  .Y({ S2646 })
);
NOR #() 
NOR_741_ (
  .A({ S1623 }),
  .B({ S2646 }),
  .Y({ S2647 })
);
NOR #() 
NOR_742_ (
  .A({ controller_fib_2 }),
  .B({ S1396 }),
  .Y({ S2648 })
);
NOR #() 
NOR_743_ (
  .A({ S2364 }),
  .B({ S2648 }),
  .Y({ S2649 })
);
NOR #() 
NOR_744_ (
  .A({ S2053 }),
  .B({ S2649 }),
  .Y({ S2650 })
);
NOR #() 
NOR_745_ (
  .A({ S1547 }),
  .B({ S2650 }),
  .Y({ S2651 })
);
NAND #() 
NAND_1483_ (
  .A({ datapath_multdivunit_outmdu1_10 }),
  .B({ S1377 }),
  .Y({ S2652 })
);
NAND #() 
NAND_1484_ (
  .A({ datapath_databusin_10 }),
  .B({ S1627 }),
  .Y({ S2653 })
);
NAND #() 
NAND_1485_ (
  .A({ datapath_multdivunit_outmdu2_10 }),
  .B({ S8570 }),
  .Y({ S2654 })
);
NOT #() 
NOT_280_ (
  .A({ S2654 }),
  .Y({ S2655 })
);
NAND #() 
NAND_1486_ (
  .A({ S2652 }),
  .B({ S2653 }),
  .Y({ S2656 })
);
NOR #() 
NOR_746_ (
  .A({ S2651 }),
  .B({ S2656 }),
  .Y({ S2657 })
);
NOR #() 
NOR_747_ (
  .A({ S2647 }),
  .B({ S2655 }),
  .Y({ S2658 })
);
NAND #() 
NAND_1487_ (
  .A({ S2657 }),
  .B({ S2658 }),
  .Y({ S2659 })
);
NOR #() 
NOR_748_ (
  .A({ S2644 }),
  .B({ S2659 }),
  .Y({ S2660 })
);
NAND #() 
NAND_1488_ (
  .A({ S2642 }),
  .B({ S2660 }),
  .Y({ S2661 })
);
NOR #() 
NOR_749_ (
  .A({ S2641 }),
  .B({ S2661 }),
  .Y({ S2662 })
);
NOR #() 
NOR_750_ (
  .A({ S702 }),
  .B({ S2541 }),
  .Y({ S2663 })
);
NAND #() 
NAND_1489_ (
  .A({ S702 }),
  .B({ S2541 }),
  .Y({ S2664 })
);
NOR #() 
NOR_751_ (
  .A({ S1539 }),
  .B({ S2663 }),
  .Y({ S2665 })
);
NAND #() 
NAND_1490_ (
  .A({ S2664 }),
  .B({ S2665 }),
  .Y({ S2666 })
);
NAND #() 
NAND_1491_ (
  .A({ S2662 }),
  .B({ S2666 }),
  .Y({ S2667 })
);
NOR #() 
NOR_752_ (
  .A({ S2638 }),
  .B({ S2667 }),
  .Y({ S2668 })
);
NAND #() 
NAND_1492_ (
  .A({ S2632 }),
  .B({ S2668 }),
  .Y({ datapath_indatatrf_10 })
);
NAND #() 
NAND_1493_ (
  .A({ datapath_indatatrf_10 }),
  .B({ S1688 }),
  .Y({ S2669 })
);
NAND #() 
NAND_1494_ (
  .A({ datapath_theregisterfile_memtrf_74 }),
  .B({ S1689 }),
  .Y({ S2670 })
);
NAND #() 
NAND_1495_ (
  .A({ S2669 }),
  .B({ S2670 }),
  .Y({ S14 })
);
NAND #() 
NAND_1496_ (
  .A({ datapath_theregisterfile_memtrf_251 }),
  .B({ S1437 }),
  .Y({ S2671 })
);
NAND #() 
NAND_1497_ (
  .A({ datapath_theregisterfile_memtrf_187 }),
  .B({ S1438 }),
  .Y({ S2672 })
);
NAND #() 
NAND_1498_ (
  .A({ S2671 }),
  .B({ S2672 }),
  .Y({ S2673 })
);
NAND #() 
NAND_1499_ (
  .A({ S1457 }),
  .B({ S2673 }),
  .Y({ S2674 })
);
NAND #() 
NAND_1500_ (
  .A({ datapath_theregisterfile_memtrf_171 }),
  .B({ S1438 }),
  .Y({ S2675 })
);
NAND #() 
NAND_1501_ (
  .A({ datapath_theregisterfile_memtrf_235 }),
  .B({ S1437 }),
  .Y({ S2676 })
);
NAND #() 
NAND_1502_ (
  .A({ S2675 }),
  .B({ S2676 }),
  .Y({ S2677 })
);
NAND #() 
NAND_1503_ (
  .A({ S1458 }),
  .B({ S2677 }),
  .Y({ S2678 })
);
NAND #() 
NAND_1504_ (
  .A({ S2674 }),
  .B({ S2678 }),
  .Y({ S2679 })
);
NAND #() 
NAND_1505_ (
  .A({ S1443 }),
  .B({ S2679 }),
  .Y({ S2680 })
);
NAND #() 
NAND_1506_ (
  .A({ datapath_theregisterfile_memtrf_155 }),
  .B({ S1438 }),
  .Y({ S2681 })
);
NAND #() 
NAND_1507_ (
  .A({ datapath_theregisterfile_memtrf_219 }),
  .B({ S1437 }),
  .Y({ S2682 })
);
NAND #() 
NAND_1508_ (
  .A({ S2681 }),
  .B({ S2682 }),
  .Y({ S2683 })
);
NAND #() 
NAND_1509_ (
  .A({ S1457 }),
  .B({ S2683 }),
  .Y({ S2684 })
);
NOR #() 
NOR_753_ (
  .A({ datapath_theregisterfile_memtrf_139 }),
  .B({ S1437 }),
  .Y({ S2685 })
);
NOR #() 
NOR_754_ (
  .A({ datapath_theregisterfile_memtrf_203 }),
  .B({ S1438 }),
  .Y({ S2686 })
);
NOR #() 
NOR_755_ (
  .A({ S2685 }),
  .B({ S2686 }),
  .Y({ S2687 })
);
NAND #() 
NAND_1510_ (
  .A({ S1458 }),
  .B({ S2687 }),
  .Y({ S2688 })
);
NAND #() 
NAND_1511_ (
  .A({ S2684 }),
  .B({ S2688 }),
  .Y({ S2689 })
);
NAND #() 
NAND_1512_ (
  .A({ S1444 }),
  .B({ S2689 }),
  .Y({ S2690 })
);
NAND #() 
NAND_1513_ (
  .A({ S2680 }),
  .B({ S2690 }),
  .Y({ S2691 })
);
NAND #() 
NAND_1514_ (
  .A({ S1449 }),
  .B({ S2691 }),
  .Y({ S2692 })
);
NAND #() 
NAND_1515_ (
  .A({ datapath_theregisterfile_memtrf_27 }),
  .B({ S1438 }),
  .Y({ S2693 })
);
NAND #() 
NAND_1516_ (
  .A({ datapath_theregisterfile_memtrf_91 }),
  .B({ S1437 }),
  .Y({ S2694 })
);
NAND #() 
NAND_1517_ (
  .A({ S2693 }),
  .B({ S2694 }),
  .Y({ S2695 })
);
NAND #() 
NAND_1518_ (
  .A({ S1926 }),
  .B({ S2695 }),
  .Y({ S2696 })
);
NAND #() 
NAND_1519_ (
  .A({ datapath_theregisterfile_memtrf_11 }),
  .B({ S1438 }),
  .Y({ S2697 })
);
NAND #() 
NAND_1520_ (
  .A({ datapath_theregisterfile_memtrf_75 }),
  .B({ S1437 }),
  .Y({ S2698 })
);
NAND #() 
NAND_1521_ (
  .A({ S2697 }),
  .B({ S2698 }),
  .Y({ S2699 })
);
NAND #() 
NAND_1522_ (
  .A({ S1459 }),
  .B({ S2699 }),
  .Y({ S2700 })
);
NAND #() 
NAND_1523_ (
  .A({ S2696 }),
  .B({ S2700 }),
  .Y({ S2701 })
);
NAND #() 
NAND_1524_ (
  .A({ datapath_theregisterfile_memtrf_123 }),
  .B({ S1437 }),
  .Y({ S2702 })
);
NAND #() 
NAND_1525_ (
  .A({ datapath_theregisterfile_memtrf_59 }),
  .B({ S1438 }),
  .Y({ S2703 })
);
NAND #() 
NAND_1526_ (
  .A({ S2702 }),
  .B({ S2703 }),
  .Y({ S2704 })
);
NAND #() 
NAND_1527_ (
  .A({ S1457 }),
  .B({ S2704 }),
  .Y({ S2705 })
);
NAND #() 
NAND_1528_ (
  .A({ datapath_theregisterfile_memtrf_107 }),
  .B({ S1437 }),
  .Y({ S2706 })
);
NAND #() 
NAND_1529_ (
  .A({ datapath_theregisterfile_memtrf_43 }),
  .B({ S1438 }),
  .Y({ S2707 })
);
NAND #() 
NAND_1530_ (
  .A({ S2706 }),
  .B({ S2707 }),
  .Y({ S2708 })
);
NAND #() 
NAND_1531_ (
  .A({ S1458 }),
  .B({ S2708 }),
  .Y({ S2709 })
);
NAND #() 
NAND_1532_ (
  .A({ S2705 }),
  .B({ S2709 }),
  .Y({ S2710 })
);
NAND #() 
NAND_1533_ (
  .A({ S1487 }),
  .B({ S2710 }),
  .Y({ S2711 })
);
NOT #() 
NOT_281_ (
  .A({ S2711 }),
  .Y({ S2712 })
);
NOR #() 
NOR_756_ (
  .A({ S2701 }),
  .B({ S2712 }),
  .Y({ S2713 })
);
NAND #() 
NAND_1534_ (
  .A({ S2692 }),
  .B({ S2711 }),
  .Y({ S2714 })
);
NOR #() 
NOR_757_ (
  .A({ S2701 }),
  .B({ S2714 }),
  .Y({ S2715 })
);
NAND #() 
NAND_1535_ (
  .A({ S2692 }),
  .B({ S2713 }),
  .Y({ S2716 })
);
NOR #() 
NOR_758_ (
  .A({ S1461 }),
  .B({ S2715 }),
  .Y({ S2717 })
);
NAND #() 
NAND_1536_ (
  .A({ S1462 }),
  .B({ S2716 }),
  .Y({ S2718 })
);
NAND #() 
NAND_1537_ (
  .A({ S1429 }),
  .B({ S2717 }),
  .Y({ S2719 })
);
NAND #() 
NAND_1538_ (
  .A({ S2369 }),
  .B({ S2719 }),
  .Y({ S2720 })
);
NOT #() 
NOT_282_ (
  .A({ S2720 }),
  .Y({ S2721 })
);
NOR #() 
NOR_759_ (
  .A({ S651 }),
  .B({ S2720 }),
  .Y({ S2722 })
);
NOR #() 
NOR_760_ (
  .A({ datapath_addsubunit_in1_11 }),
  .B({ S2721 }),
  .Y({ S2723 })
);
NOR #() 
NOR_761_ (
  .A({ S2722 }),
  .B({ S2723 }),
  .Y({ S2724 })
);
NOT #() 
NOT_283_ (
  .A({ S2724 }),
  .Y({ S2725 })
);
NAND #() 
NAND_1539_ (
  .A({ S2624 }),
  .B({ S2630 }),
  .Y({ S2726 })
);
NOR #() 
NOR_762_ (
  .A({ S2724 }),
  .B({ S2726 }),
  .Y({ S2727 })
);
NAND #() 
NAND_1540_ (
  .A({ S2724 }),
  .B({ S2726 }),
  .Y({ S2728 })
);
NAND #() 
NAND_1541_ (
  .A({ S1525 }),
  .B({ S2728 }),
  .Y({ S2729 })
);
NOR #() 
NOR_763_ (
  .A({ S2727 }),
  .B({ S2729 }),
  .Y({ S2730 })
);
NOR #() 
NOR_764_ (
  .A({ S2635 }),
  .B({ S2640 }),
  .Y({ S2731 })
);
NAND #() 
NAND_1542_ (
  .A({ S2724 }),
  .B({ S2731 }),
  .Y({ S2732 })
);
NOR #() 
NOR_765_ (
  .A({ S2724 }),
  .B({ S2731 }),
  .Y({ S2733 })
);
NOR #() 
NOR_766_ (
  .A({ S1528 }),
  .B({ S2733 }),
  .Y({ S2734 })
);
NAND #() 
NAND_1543_ (
  .A({ S2732 }),
  .B({ S2734 }),
  .Y({ S2735 })
);
NAND #() 
NAND_1544_ (
  .A({ datapath_addsubunit_in1_11 }),
  .B({ S2664 }),
  .Y({ S2736 })
);
NOR #() 
NOR_767_ (
  .A({ datapath_addsubunit_in1_11 }),
  .B({ S2664 }),
  .Y({ S2737 })
);
NOR #() 
NOR_768_ (
  .A({ S1539 }),
  .B({ S2737 }),
  .Y({ S2738 })
);
NAND #() 
NAND_1545_ (
  .A({ S2736 }),
  .B({ S2738 }),
  .Y({ S2739 })
);
NAND #() 
NAND_1546_ (
  .A({ datapath_addsubunit_in1_11 }),
  .B({ S2720 }),
  .Y({ S2740 })
);
NOR #() 
NOR_769_ (
  .A({ S1533 }),
  .B({ S2740 }),
  .Y({ S2741 })
);
NAND #() 
NAND_1547_ (
  .A({ datapath_shiftunit_2333_A }),
  .B({ S1614 }),
  .Y({ S2742 })
);
NAND #() 
NAND_1548_ (
  .A({ datapath_shiftunit_2637_A }),
  .B({ S1609 }),
  .Y({ S2743 })
);
NOT #() 
NOT_284_ (
  .A({ S2743 }),
  .Y({ S2744 })
);
NOR #() 
NOR_770_ (
  .A({ datapath_muxmem_in2_11 }),
  .B({ S1353 }),
  .Y({ S2745 })
);
NAND #() 
NAND_1549_ (
  .A({ S7978 }),
  .B({ S1354 }),
  .Y({ S2746 })
);
NOR #() 
NOR_771_ (
  .A({ S1355 }),
  .B({ S2745 }),
  .Y({ S2747 })
);
NAND #() 
NAND_1550_ (
  .A({ S1356 }),
  .B({ S2746 }),
  .Y({ S2748 })
);
NAND #() 
NAND_1551_ (
  .A({ S1622 }),
  .B({ S2747 }),
  .Y({ S2749 })
);
NOR #() 
NOR_772_ (
  .A({ controller_fib_3 }),
  .B({ S1396 }),
  .Y({ S2750 })
);
NOR #() 
NOR_773_ (
  .A({ S2364 }),
  .B({ S2750 }),
  .Y({ S2751 })
);
NOR #() 
NOR_774_ (
  .A({ S2053 }),
  .B({ S2751 }),
  .Y({ S2752 })
);
NOR #() 
NOR_775_ (
  .A({ S1547 }),
  .B({ S2752 }),
  .Y({ S2753 })
);
NAND #() 
NAND_1552_ (
  .A({ datapath_databusin_11 }),
  .B({ S1627 }),
  .Y({ S2754 })
);
NAND #() 
NAND_1553_ (
  .A({ datapath_multdivunit_outmdu1_11 }),
  .B({ S1377 }),
  .Y({ S2755 })
);
NAND #() 
NAND_1554_ (
  .A({ datapath_multdivunit_outmdu2_11 }),
  .B({ S8570 }),
  .Y({ S2756 })
);
NAND #() 
NAND_1555_ (
  .A({ S2755 }),
  .B({ S2756 }),
  .Y({ S2757 })
);
NOT #() 
NOT_285_ (
  .A({ S2757 }),
  .Y({ S2758 })
);
NAND #() 
NAND_1556_ (
  .A({ S2754 }),
  .B({ S2758 }),
  .Y({ S2759 })
);
NOR #() 
NOR_776_ (
  .A({ S2753 }),
  .B({ S2759 }),
  .Y({ S2760 })
);
NAND #() 
NAND_1557_ (
  .A({ S2749 }),
  .B({ S2760 }),
  .Y({ S2761 })
);
NOR #() 
NOR_777_ (
  .A({ S2744 }),
  .B({ S2761 }),
  .Y({ S2762 })
);
NAND #() 
NAND_1558_ (
  .A({ S2742 }),
  .B({ S2762 }),
  .Y({ S2763 })
);
NOR #() 
NOR_778_ (
  .A({ S2741 }),
  .B({ S2763 }),
  .Y({ S2764 })
);
NAND #() 
NAND_1559_ (
  .A({ S2739 }),
  .B({ S2764 }),
  .Y({ S2765 })
);
NOR #() 
NOR_779_ (
  .A({ S2730 }),
  .B({ S2765 }),
  .Y({ S2766 })
);
NAND #() 
NAND_1560_ (
  .A({ S2735 }),
  .B({ S2766 }),
  .Y({ datapath_indatatrf_11 })
);
NAND #() 
NAND_1561_ (
  .A({ datapath_indatatrf_11 }),
  .B({ S1688 }),
  .Y({ S2767 })
);
NAND #() 
NAND_1562_ (
  .A({ datapath_theregisterfile_memtrf_75 }),
  .B({ S1689 }),
  .Y({ S2768 })
);
NAND #() 
NAND_1563_ (
  .A({ S2767 }),
  .B({ S2768 }),
  .Y({ S15 })
);
NAND #() 
NAND_1564_ (
  .A({ datapath_theregisterfile_memtrf_252 }),
  .B({ S1437 }),
  .Y({ S2769 })
);
NAND #() 
NAND_1565_ (
  .A({ datapath_theregisterfile_memtrf_188 }),
  .B({ S1438 }),
  .Y({ S2770 })
);
NAND #() 
NAND_1566_ (
  .A({ S2769 }),
  .B({ S2770 }),
  .Y({ S2771 })
);
NAND #() 
NAND_1567_ (
  .A({ S1457 }),
  .B({ S2771 }),
  .Y({ S2772 })
);
NAND #() 
NAND_1568_ (
  .A({ datapath_theregisterfile_memtrf_172 }),
  .B({ S1438 }),
  .Y({ S2773 })
);
NAND #() 
NAND_1569_ (
  .A({ datapath_theregisterfile_memtrf_236 }),
  .B({ S1437 }),
  .Y({ S2774 })
);
NAND #() 
NAND_1570_ (
  .A({ S2773 }),
  .B({ S2774 }),
  .Y({ S2775 })
);
NAND #() 
NAND_1571_ (
  .A({ S1458 }),
  .B({ S2775 }),
  .Y({ S2776 })
);
NAND #() 
NAND_1572_ (
  .A({ S2772 }),
  .B({ S2776 }),
  .Y({ S2777 })
);
NAND #() 
NAND_1573_ (
  .A({ datapath_theregisterfile_memtrf_156 }),
  .B({ S1438 }),
  .Y({ S2778 })
);
NAND #() 
NAND_1574_ (
  .A({ datapath_theregisterfile_memtrf_220 }),
  .B({ S1437 }),
  .Y({ S2779 })
);
NAND #() 
NAND_1575_ (
  .A({ S2778 }),
  .B({ S2779 }),
  .Y({ S2780 })
);
NAND #() 
NAND_1576_ (
  .A({ S1457 }),
  .B({ S2780 }),
  .Y({ S2781 })
);
NOR #() 
NOR_780_ (
  .A({ datapath_theregisterfile_memtrf_140 }),
  .B({ S1437 }),
  .Y({ S2782 })
);
NAND #() 
NAND_1577_ (
  .A({ S7750 }),
  .B({ S1437 }),
  .Y({ S2783 })
);
NAND #() 
NAND_1578_ (
  .A({ S1458 }),
  .B({ S2783 }),
  .Y({ S2784 })
);
NOR #() 
NOR_781_ (
  .A({ S2782 }),
  .B({ S2784 }),
  .Y({ S2785 })
);
NOR #() 
NOR_782_ (
  .A({ S1444 }),
  .B({ S2777 }),
  .Y({ S2786 })
);
NOR #() 
NOR_783_ (
  .A({ S1443 }),
  .B({ S2785 }),
  .Y({ S2787 })
);
NAND #() 
NAND_1579_ (
  .A({ S2781 }),
  .B({ S2787 }),
  .Y({ S2788 })
);
NAND #() 
NAND_1580_ (
  .A({ S1449 }),
  .B({ S2788 }),
  .Y({ S2789 })
);
NOR #() 
NOR_784_ (
  .A({ S2786 }),
  .B({ S2789 }),
  .Y({ S2790 })
);
NAND #() 
NAND_1581_ (
  .A({ datapath_theregisterfile_memtrf_108 }),
  .B({ S1458 }),
  .Y({ S2791 })
);
NAND #() 
NAND_1582_ (
  .A({ datapath_theregisterfile_memtrf_124 }),
  .B({ S1457 }),
  .Y({ S2792 })
);
NAND #() 
NAND_1583_ (
  .A({ S2791 }),
  .B({ S2792 }),
  .Y({ S2793 })
);
NAND #() 
NAND_1584_ (
  .A({ S1437 }),
  .B({ S2793 }),
  .Y({ S2794 })
);
NAND #() 
NAND_1585_ (
  .A({ datapath_theregisterfile_memtrf_44 }),
  .B({ S1458 }),
  .Y({ S2795 })
);
NAND #() 
NAND_1586_ (
  .A({ datapath_theregisterfile_memtrf_60 }),
  .B({ S1457 }),
  .Y({ S2796 })
);
NAND #() 
NAND_1587_ (
  .A({ S2795 }),
  .B({ S2796 }),
  .Y({ S2797 })
);
NAND #() 
NAND_1588_ (
  .A({ S1438 }),
  .B({ S2797 }),
  .Y({ S2798 })
);
NAND #() 
NAND_1589_ (
  .A({ S2794 }),
  .B({ S2798 }),
  .Y({ S2799 })
);
NAND #() 
NAND_1590_ (
  .A({ S1487 }),
  .B({ S2799 }),
  .Y({ S2800 })
);
NOR #() 
NOR_785_ (
  .A({ datapath_theregisterfile_memtrf_76 }),
  .B({ S1438 }),
  .Y({ S2801 })
);
NOR #() 
NOR_786_ (
  .A({ datapath_theregisterfile_memtrf_12 }),
  .B({ S1437 }),
  .Y({ S2802 })
);
NOR #() 
NOR_787_ (
  .A({ S2801 }),
  .B({ S2802 }),
  .Y({ S2803 })
);
NAND #() 
NAND_1591_ (
  .A({ S1459 }),
  .B({ S2803 }),
  .Y({ S2804 })
);
NAND #() 
NAND_1592_ (
  .A({ datapath_theregisterfile_memtrf_28 }),
  .B({ S1438 }),
  .Y({ S2805 })
);
NAND #() 
NAND_1593_ (
  .A({ datapath_theregisterfile_memtrf_92 }),
  .B({ S1437 }),
  .Y({ S2806 })
);
NAND #() 
NAND_1594_ (
  .A({ S2805 }),
  .B({ S2806 }),
  .Y({ S2807 })
);
NAND #() 
NAND_1595_ (
  .A({ S1926 }),
  .B({ S2807 }),
  .Y({ S2808 })
);
NAND #() 
NAND_1596_ (
  .A({ S2804 }),
  .B({ S2808 }),
  .Y({ S2809 })
);
NOT #() 
NOT_286_ (
  .A({ S2809 }),
  .Y({ S2810 })
);
NAND #() 
NAND_1597_ (
  .A({ S2800 }),
  .B({ S2810 }),
  .Y({ S2811 })
);
NAND #() 
NAND_1598_ (
  .A({ S2800 }),
  .B({ S2808 }),
  .Y({ S2812 })
);
NOR #() 
NOR_788_ (
  .A({ S2790 }),
  .B({ S2812 }),
  .Y({ S2813 })
);
NOR #() 
NOR_789_ (
  .A({ S2790 }),
  .B({ S2811 }),
  .Y({ S2814 })
);
NAND #() 
NAND_1599_ (
  .A({ S2804 }),
  .B({ S2813 }),
  .Y({ S2815 })
);
NOR #() 
NOR_790_ (
  .A({ S1461 }),
  .B({ S2814 }),
  .Y({ S2816 })
);
NAND #() 
NAND_1600_ (
  .A({ S1462 }),
  .B({ S2815 }),
  .Y({ S2817 })
);
NAND #() 
NAND_1601_ (
  .A({ S1429 }),
  .B({ S2816 }),
  .Y({ S2818 })
);
NAND #() 
NAND_1602_ (
  .A({ S2369 }),
  .B({ S2818 }),
  .Y({ S2819 })
);
NOT #() 
NOT_287_ (
  .A({ S2819 }),
  .Y({ S2820 })
);
NOR #() 
NOR_791_ (
  .A({ S599 }),
  .B({ S2819 }),
  .Y({ S2821 })
);
NOT #() 
NOT_288_ (
  .A({ S2821 }),
  .Y({ S2822 })
);
NOR #() 
NOR_792_ (
  .A({ datapath_addsubunit_in1_12 }),
  .B({ S2820 }),
  .Y({ S2823 })
);
NOR #() 
NOR_793_ (
  .A({ S2821 }),
  .B({ S2823 }),
  .Y({ S2824 })
);
NOR #() 
NOR_794_ (
  .A({ S2722 }),
  .B({ S2726 }),
  .Y({ S2825 })
);
NOR #() 
NOR_795_ (
  .A({ S2723 }),
  .B({ S2825 }),
  .Y({ S2826 })
);
NOR #() 
NOR_796_ (
  .A({ S2824 }),
  .B({ S2826 }),
  .Y({ S2827 })
);
NAND #() 
NAND_1603_ (
  .A({ S2824 }),
  .B({ S2826 }),
  .Y({ S2828 })
);
NAND #() 
NAND_1604_ (
  .A({ S1525 }),
  .B({ S2828 }),
  .Y({ S2829 })
);
NOR #() 
NOR_797_ (
  .A({ S2827 }),
  .B({ S2829 }),
  .Y({ S2830 })
);
NAND #() 
NAND_1605_ (
  .A({ S2635 }),
  .B({ S2725 }),
  .Y({ S2831 })
);
NOR #() 
NOR_798_ (
  .A({ S2639 }),
  .B({ S2724 }),
  .Y({ S2832 })
);
NAND #() 
NAND_1606_ (
  .A({ S2740 }),
  .B({ S2831 }),
  .Y({ S2833 })
);
NOR #() 
NOR_799_ (
  .A({ S2832 }),
  .B({ S2833 }),
  .Y({ S2834 })
);
NAND #() 
NAND_1607_ (
  .A({ S2824 }),
  .B({ S2834 }),
  .Y({ S2835 })
);
NOR #() 
NOR_800_ (
  .A({ S2824 }),
  .B({ S2834 }),
  .Y({ S2836 })
);
NOR #() 
NOR_801_ (
  .A({ S1528 }),
  .B({ S2836 }),
  .Y({ S2837 })
);
NAND #() 
NAND_1608_ (
  .A({ S2835 }),
  .B({ S2837 }),
  .Y({ S2838 })
);
NAND #() 
NAND_1609_ (
  .A({ datapath_addsubunit_in1_12 }),
  .B({ S2819 }),
  .Y({ S2839 })
);
NOR #() 
NOR_802_ (
  .A({ S1533 }),
  .B({ S2839 }),
  .Y({ S2840 })
);
NAND #() 
NAND_1610_ (
  .A({ datapath_shiftunit_2351_A }),
  .B({ S1614 }),
  .Y({ S2841 })
);
NAND #() 
NAND_1611_ (
  .A({ datapath_shiftunit_2655_A }),
  .B({ S1609 }),
  .Y({ S2842 })
);
NOT #() 
NOT_289_ (
  .A({ S2842 }),
  .Y({ S2843 })
);
NOR #() 
NOR_803_ (
  .A({ datapath_muxmem_in2_12 }),
  .B({ S1355 }),
  .Y({ S2844 })
);
NAND #() 
NAND_1612_ (
  .A({ S7989 }),
  .B({ S1356 }),
  .Y({ S2845 })
);
NOR #() 
NOR_804_ (
  .A({ S1357 }),
  .B({ S2844 }),
  .Y({ S2846 })
);
NAND #() 
NAND_1613_ (
  .A({ S1358 }),
  .B({ S2845 }),
  .Y({ S2847 })
);
NAND #() 
NAND_1614_ (
  .A({ S1622 }),
  .B({ S2846 }),
  .Y({ S2848 })
);
NOR #() 
NOR_805_ (
  .A({ controller_fib_4 }),
  .B({ S1396 }),
  .Y({ S2849 })
);
NOR #() 
NOR_806_ (
  .A({ S2364 }),
  .B({ S2849 }),
  .Y({ S2850 })
);
NOR #() 
NOR_807_ (
  .A({ S2053 }),
  .B({ S2850 }),
  .Y({ S2851 })
);
NOR #() 
NOR_808_ (
  .A({ S1547 }),
  .B({ S2851 }),
  .Y({ S2852 })
);
NAND #() 
NAND_1615_ (
  .A({ datapath_databusin_12 }),
  .B({ S1627 }),
  .Y({ S2853 })
);
NAND #() 
NAND_1616_ (
  .A({ datapath_multdivunit_outmdu1_12 }),
  .B({ S1377 }),
  .Y({ S2854 })
);
NAND #() 
NAND_1617_ (
  .A({ datapath_multdivunit_outmdu2_12 }),
  .B({ S8570 }),
  .Y({ S2855 })
);
NAND #() 
NAND_1618_ (
  .A({ S2854 }),
  .B({ S2855 }),
  .Y({ S2856 })
);
NOT #() 
NOT_290_ (
  .A({ S2856 }),
  .Y({ S2857 })
);
NAND #() 
NAND_1619_ (
  .A({ S2853 }),
  .B({ S2857 }),
  .Y({ S2858 })
);
NOR #() 
NOR_809_ (
  .A({ S2852 }),
  .B({ S2858 }),
  .Y({ S2859 })
);
NAND #() 
NAND_1620_ (
  .A({ S2848 }),
  .B({ S2859 }),
  .Y({ S2860 })
);
NOR #() 
NOR_810_ (
  .A({ S2843 }),
  .B({ S2860 }),
  .Y({ S2861 })
);
NAND #() 
NAND_1621_ (
  .A({ S2841 }),
  .B({ S2861 }),
  .Y({ S2862 })
);
NOR #() 
NOR_811_ (
  .A({ S2840 }),
  .B({ S2862 }),
  .Y({ S2863 })
);
NAND #() 
NAND_1622_ (
  .A({ S599 }),
  .B({ S2737 }),
  .Y({ S2864 })
);
NOR #() 
NOR_812_ (
  .A({ S599 }),
  .B({ S2737 }),
  .Y({ S2865 })
);
NOR #() 
NOR_813_ (
  .A({ S1539 }),
  .B({ S2865 }),
  .Y({ S2866 })
);
NAND #() 
NAND_1623_ (
  .A({ S2864 }),
  .B({ S2866 }),
  .Y({ S2867 })
);
NAND #() 
NAND_1624_ (
  .A({ S2863 }),
  .B({ S2867 }),
  .Y({ S2868 })
);
NOR #() 
NOR_814_ (
  .A({ S2830 }),
  .B({ S2868 }),
  .Y({ S2869 })
);
NAND #() 
NAND_1625_ (
  .A({ S2838 }),
  .B({ S2869 }),
  .Y({ datapath_indatatrf_12 })
);
NAND #() 
NAND_1626_ (
  .A({ datapath_indatatrf_12 }),
  .B({ S1688 }),
  .Y({ S2870 })
);
NAND #() 
NAND_1627_ (
  .A({ datapath_theregisterfile_memtrf_76 }),
  .B({ S1689 }),
  .Y({ S2871 })
);
NAND #() 
NAND_1628_ (
  .A({ S2870 }),
  .B({ S2871 }),
  .Y({ S16 })
);
NAND #() 
NAND_1629_ (
  .A({ datapath_theregisterfile_memtrf_253 }),
  .B({ S1437 }),
  .Y({ S2872 })
);
NAND #() 
NAND_1630_ (
  .A({ datapath_theregisterfile_memtrf_189 }),
  .B({ S1438 }),
  .Y({ S2873 })
);
NAND #() 
NAND_1631_ (
  .A({ S2872 }),
  .B({ S2873 }),
  .Y({ S2874 })
);
NAND #() 
NAND_1632_ (
  .A({ S1457 }),
  .B({ S2874 }),
  .Y({ S2875 })
);
NAND #() 
NAND_1633_ (
  .A({ datapath_theregisterfile_memtrf_173 }),
  .B({ S1438 }),
  .Y({ S2876 })
);
NAND #() 
NAND_1634_ (
  .A({ datapath_theregisterfile_memtrf_237 }),
  .B({ S1437 }),
  .Y({ S2877 })
);
NAND #() 
NAND_1635_ (
  .A({ S2876 }),
  .B({ S2877 }),
  .Y({ S2878 })
);
NAND #() 
NAND_1636_ (
  .A({ S1458 }),
  .B({ S2878 }),
  .Y({ S2879 })
);
NAND #() 
NAND_1637_ (
  .A({ S2875 }),
  .B({ S2879 }),
  .Y({ S2880 })
);
NAND #() 
NAND_1638_ (
  .A({ datapath_theregisterfile_memtrf_157 }),
  .B({ S1438 }),
  .Y({ S2881 })
);
NAND #() 
NAND_1639_ (
  .A({ datapath_theregisterfile_memtrf_221 }),
  .B({ S1437 }),
  .Y({ S2882 })
);
NAND #() 
NAND_1640_ (
  .A({ S2881 }),
  .B({ S2882 }),
  .Y({ S2883 })
);
NAND #() 
NAND_1641_ (
  .A({ S1457 }),
  .B({ S2883 }),
  .Y({ S2884 })
);
NOR #() 
NOR_815_ (
  .A({ datapath_theregisterfile_memtrf_141 }),
  .B({ S1437 }),
  .Y({ S2885 })
);
NAND #() 
NAND_1642_ (
  .A({ S7761 }),
  .B({ S1437 }),
  .Y({ S2886 })
);
NAND #() 
NAND_1643_ (
  .A({ S1458 }),
  .B({ S2886 }),
  .Y({ S2887 })
);
NOR #() 
NOR_816_ (
  .A({ S2885 }),
  .B({ S2887 }),
  .Y({ S2888 })
);
NOR #() 
NOR_817_ (
  .A({ S1444 }),
  .B({ S2880 }),
  .Y({ S2889 })
);
NOR #() 
NOR_818_ (
  .A({ S1443 }),
  .B({ S2888 }),
  .Y({ S2890 })
);
NAND #() 
NAND_1644_ (
  .A({ S2884 }),
  .B({ S2890 }),
  .Y({ S2891 })
);
NAND #() 
NAND_1645_ (
  .A({ S1449 }),
  .B({ S2891 }),
  .Y({ S2892 })
);
NOR #() 
NOR_819_ (
  .A({ S2889 }),
  .B({ S2892 }),
  .Y({ S2893 })
);
NAND #() 
NAND_1646_ (
  .A({ datapath_theregisterfile_memtrf_109 }),
  .B({ S1458 }),
  .Y({ S2894 })
);
NAND #() 
NAND_1647_ (
  .A({ datapath_theregisterfile_memtrf_125 }),
  .B({ S1457 }),
  .Y({ S2895 })
);
NAND #() 
NAND_1648_ (
  .A({ S2894 }),
  .B({ S2895 }),
  .Y({ S2896 })
);
NAND #() 
NAND_1649_ (
  .A({ S1437 }),
  .B({ S2896 }),
  .Y({ S2897 })
);
NAND #() 
NAND_1650_ (
  .A({ datapath_theregisterfile_memtrf_45 }),
  .B({ S1458 }),
  .Y({ S2898 })
);
NAND #() 
NAND_1651_ (
  .A({ datapath_theregisterfile_memtrf_61 }),
  .B({ S1457 }),
  .Y({ S2899 })
);
NAND #() 
NAND_1652_ (
  .A({ S2898 }),
  .B({ S2899 }),
  .Y({ S2900 })
);
NAND #() 
NAND_1653_ (
  .A({ S1438 }),
  .B({ S2900 }),
  .Y({ S2901 })
);
NAND #() 
NAND_1654_ (
  .A({ S2897 }),
  .B({ S2901 }),
  .Y({ S2902 })
);
NAND #() 
NAND_1655_ (
  .A({ S1487 }),
  .B({ S2902 }),
  .Y({ S2903 })
);
NOR #() 
NOR_820_ (
  .A({ datapath_theregisterfile_memtrf_77 }),
  .B({ S1438 }),
  .Y({ S2904 })
);
NOR #() 
NOR_821_ (
  .A({ datapath_theregisterfile_memtrf_13 }),
  .B({ S1437 }),
  .Y({ S2905 })
);
NOR #() 
NOR_822_ (
  .A({ S2904 }),
  .B({ S2905 }),
  .Y({ S2906 })
);
NAND #() 
NAND_1656_ (
  .A({ S1459 }),
  .B({ S2906 }),
  .Y({ S2907 })
);
NAND #() 
NAND_1657_ (
  .A({ datapath_theregisterfile_memtrf_29 }),
  .B({ S1438 }),
  .Y({ S2908 })
);
NAND #() 
NAND_1658_ (
  .A({ datapath_theregisterfile_memtrf_93 }),
  .B({ S1437 }),
  .Y({ S2909 })
);
NAND #() 
NAND_1659_ (
  .A({ S2908 }),
  .B({ S2909 }),
  .Y({ S2910 })
);
NAND #() 
NAND_1660_ (
  .A({ S1926 }),
  .B({ S2910 }),
  .Y({ S2911 })
);
NAND #() 
NAND_1661_ (
  .A({ S2907 }),
  .B({ S2911 }),
  .Y({ S2912 })
);
NOT #() 
NOT_291_ (
  .A({ S2912 }),
  .Y({ S2913 })
);
NAND #() 
NAND_1662_ (
  .A({ S2903 }),
  .B({ S2913 }),
  .Y({ S2914 })
);
NAND #() 
NAND_1663_ (
  .A({ S2903 }),
  .B({ S2911 }),
  .Y({ S2915 })
);
NOR #() 
NOR_823_ (
  .A({ S2893 }),
  .B({ S2915 }),
  .Y({ S2916 })
);
NOR #() 
NOR_824_ (
  .A({ S2893 }),
  .B({ S2914 }),
  .Y({ S2917 })
);
NAND #() 
NAND_1664_ (
  .A({ S2907 }),
  .B({ S2916 }),
  .Y({ S2918 })
);
NOR #() 
NOR_825_ (
  .A({ S1461 }),
  .B({ S2917 }),
  .Y({ S2919 })
);
NAND #() 
NAND_1665_ (
  .A({ S1462 }),
  .B({ S2918 }),
  .Y({ S2920 })
);
NOR #() 
NOR_826_ (
  .A({ S1430 }),
  .B({ S2920 }),
  .Y({ S2921 })
);
NOT #() 
NOT_292_ (
  .A({ S2921 }),
  .Y({ S2922 })
);
NAND #() 
NAND_1666_ (
  .A({ S2369 }),
  .B({ S2922 }),
  .Y({ S2923 })
);
NOT #() 
NOT_293_ (
  .A({ S2923 }),
  .Y({ S2924 })
);
NOR #() 
NOR_827_ (
  .A({ S548 }),
  .B({ S2923 }),
  .Y({ S2925 })
);
NOT #() 
NOT_294_ (
  .A({ S2925 }),
  .Y({ S2926 })
);
NOR #() 
NOR_828_ (
  .A({ datapath_addsubunit_in1_13 }),
  .B({ S2924 }),
  .Y({ S2927 })
);
NOT #() 
NOT_295_ (
  .A({ S2927 }),
  .Y({ S2928 })
);
NAND #() 
NAND_1667_ (
  .A({ S2926 }),
  .B({ S2928 }),
  .Y({ S2929 })
);
NOT #() 
NOT_296_ (
  .A({ S2929 }),
  .Y({ S2930 })
);
NAND #() 
NAND_1668_ (
  .A({ S2822 }),
  .B({ S2828 }),
  .Y({ S2931 })
);
NAND #() 
NAND_1669_ (
  .A({ S2929 }),
  .B({ S2931 }),
  .Y({ S2932 })
);
NOR #() 
NOR_829_ (
  .A({ S2929 }),
  .B({ S2931 }),
  .Y({ S2933 })
);
NOT #() 
NOT_297_ (
  .A({ S2933 }),
  .Y({ S2934 })
);
NAND #() 
NAND_1670_ (
  .A({ S2932 }),
  .B({ S2934 }),
  .Y({ S2935 })
);
NAND #() 
NAND_1671_ (
  .A({ S1525 }),
  .B({ S2935 }),
  .Y({ S2936 })
);
NAND #() 
NAND_1672_ (
  .A({ S2839 }),
  .B({ S2930 }),
  .Y({ S2937 })
);
NOR #() 
NOR_830_ (
  .A({ S2836 }),
  .B({ S2937 }),
  .Y({ S2938 })
);
NAND #() 
NAND_1673_ (
  .A({ S2836 }),
  .B({ S2929 }),
  .Y({ S2939 })
);
NOR #() 
NOR_831_ (
  .A({ S2839 }),
  .B({ S2930 }),
  .Y({ S2940 })
);
NOR #() 
NOR_832_ (
  .A({ S1528 }),
  .B({ S2940 }),
  .Y({ S2941 })
);
NAND #() 
NAND_1674_ (
  .A({ S2939 }),
  .B({ S2941 }),
  .Y({ S2942 })
);
NOR #() 
NOR_833_ (
  .A({ S2938 }),
  .B({ S2942 }),
  .Y({ S2943 })
);
NAND #() 
NAND_1675_ (
  .A({ datapath_addsubunit_in1_13 }),
  .B({ S2864 }),
  .Y({ S2944 })
);
NOR #() 
NOR_834_ (
  .A({ datapath_addsubunit_in1_13 }),
  .B({ S2864 }),
  .Y({ S2945 })
);
NOT #() 
NOT_298_ (
  .A({ S2945 }),
  .Y({ S2946 })
);
NOR #() 
NOR_835_ (
  .A({ S1539 }),
  .B({ S2945 }),
  .Y({ S2947 })
);
NAND #() 
NAND_1676_ (
  .A({ S2944 }),
  .B({ S2947 }),
  .Y({ S2948 })
);
NAND #() 
NAND_1677_ (
  .A({ datapath_addsubunit_in1_13 }),
  .B({ S2923 }),
  .Y({ S2949 })
);
NOR #() 
NOR_836_ (
  .A({ S1533 }),
  .B({ S2949 }),
  .Y({ S2950 })
);
NAND #() 
NAND_1678_ (
  .A({ datapath_shiftunit_2369_A }),
  .B({ S1614 }),
  .Y({ S2951 })
);
NAND #() 
NAND_1679_ (
  .A({ datapath_shiftunit_2673_A }),
  .B({ S1609 }),
  .Y({ S2952 })
);
NOT #() 
NOT_299_ (
  .A({ S2952 }),
  .Y({ S2953 })
);
NOR #() 
NOR_837_ (
  .A({ datapath_muxmem_in2_13 }),
  .B({ S1357 }),
  .Y({ S2954 })
);
NOR #() 
NOR_838_ (
  .A({ S1359 }),
  .B({ S2954 }),
  .Y({ S2955 })
);
NOT #() 
NOT_300_ (
  .A({ S2955 }),
  .Y({ S2956 })
);
NAND #() 
NAND_1680_ (
  .A({ S1622 }),
  .B({ S2955 }),
  .Y({ S2957 })
);
NOR #() 
NOR_839_ (
  .A({ controller_216_B_0 }),
  .B({ S1396 }),
  .Y({ S2958 })
);
NOR #() 
NOR_840_ (
  .A({ S2364 }),
  .B({ S2958 }),
  .Y({ S2959 })
);
NOR #() 
NOR_841_ (
  .A({ S2053 }),
  .B({ S2959 }),
  .Y({ S2960 })
);
NOR #() 
NOR_842_ (
  .A({ S1547 }),
  .B({ S2960 }),
  .Y({ S2961 })
);
NAND #() 
NAND_1681_ (
  .A({ datapath_multdivunit_outmdu1_13 }),
  .B({ S1377 }),
  .Y({ S2962 })
);
NAND #() 
NAND_1682_ (
  .A({ datapath_multdivunit_outmdu2_13 }),
  .B({ S8570 }),
  .Y({ S2963 })
);
NAND #() 
NAND_1683_ (
  .A({ datapath_databusin_13 }),
  .B({ S1627 }),
  .Y({ S2964 })
);
NAND #() 
NAND_1684_ (
  .A({ S2963 }),
  .B({ S2964 }),
  .Y({ S2965 })
);
NOT #() 
NOT_301_ (
  .A({ S2965 }),
  .Y({ S2966 })
);
NAND #() 
NAND_1685_ (
  .A({ S2962 }),
  .B({ S2966 }),
  .Y({ S2967 })
);
NOR #() 
NOR_843_ (
  .A({ S2961 }),
  .B({ S2967 }),
  .Y({ S2968 })
);
NAND #() 
NAND_1686_ (
  .A({ S2957 }),
  .B({ S2968 }),
  .Y({ S2969 })
);
NOR #() 
NOR_844_ (
  .A({ S2953 }),
  .B({ S2969 }),
  .Y({ S2970 })
);
NAND #() 
NAND_1687_ (
  .A({ S2951 }),
  .B({ S2970 }),
  .Y({ S2971 })
);
NOR #() 
NOR_845_ (
  .A({ S2950 }),
  .B({ S2971 }),
  .Y({ S2972 })
);
NAND #() 
NAND_1688_ (
  .A({ S2948 }),
  .B({ S2972 }),
  .Y({ S2973 })
);
NOR #() 
NOR_846_ (
  .A({ S2943 }),
  .B({ S2973 }),
  .Y({ S2974 })
);
NAND #() 
NAND_1689_ (
  .A({ S2936 }),
  .B({ S2974 }),
  .Y({ datapath_indatatrf_13 })
);
NAND #() 
NAND_1690_ (
  .A({ datapath_indatatrf_13 }),
  .B({ S1688 }),
  .Y({ S2975 })
);
NAND #() 
NAND_1691_ (
  .A({ datapath_theregisterfile_memtrf_77 }),
  .B({ S1689 }),
  .Y({ S2976 })
);
NAND #() 
NAND_1692_ (
  .A({ S2975 }),
  .B({ S2976 }),
  .Y({ S17 })
);
NAND #() 
NAND_1693_ (
  .A({ datapath_theregisterfile_memtrf_254 }),
  .B({ S1437 }),
  .Y({ S2977 })
);
NAND #() 
NAND_1694_ (
  .A({ datapath_theregisterfile_memtrf_190 }),
  .B({ S1438 }),
  .Y({ S2978 })
);
NAND #() 
NAND_1695_ (
  .A({ S2977 }),
  .B({ S2978 }),
  .Y({ S2979 })
);
NAND #() 
NAND_1696_ (
  .A({ S1457 }),
  .B({ S2979 }),
  .Y({ S2980 })
);
NAND #() 
NAND_1697_ (
  .A({ datapath_theregisterfile_memtrf_174 }),
  .B({ S1438 }),
  .Y({ S2981 })
);
NAND #() 
NAND_1698_ (
  .A({ datapath_theregisterfile_memtrf_238 }),
  .B({ S1437 }),
  .Y({ S2982 })
);
NAND #() 
NAND_1699_ (
  .A({ S2981 }),
  .B({ S2982 }),
  .Y({ S2983 })
);
NAND #() 
NAND_1700_ (
  .A({ S1458 }),
  .B({ S2983 }),
  .Y({ S2984 })
);
NAND #() 
NAND_1701_ (
  .A({ S2980 }),
  .B({ S2984 }),
  .Y({ S2985 })
);
NAND #() 
NAND_1702_ (
  .A({ S1443 }),
  .B({ S2985 }),
  .Y({ S2986 })
);
NAND #() 
NAND_1703_ (
  .A({ datapath_theregisterfile_memtrf_158 }),
  .B({ S1438 }),
  .Y({ S2987 })
);
NAND #() 
NAND_1704_ (
  .A({ datapath_theregisterfile_memtrf_222 }),
  .B({ S1437 }),
  .Y({ S2988 })
);
NAND #() 
NAND_1705_ (
  .A({ S2987 }),
  .B({ S2988 }),
  .Y({ S2989 })
);
NAND #() 
NAND_1706_ (
  .A({ S1457 }),
  .B({ S2989 }),
  .Y({ S2990 })
);
NOR #() 
NOR_847_ (
  .A({ datapath_theregisterfile_memtrf_142 }),
  .B({ S1437 }),
  .Y({ S2991 })
);
NOR #() 
NOR_848_ (
  .A({ datapath_theregisterfile_memtrf_206 }),
  .B({ S1438 }),
  .Y({ S2992 })
);
NAND #() 
NAND_1707_ (
  .A({ S7772 }),
  .B({ S1437 }),
  .Y({ S2993 })
);
NOR #() 
NOR_849_ (
  .A({ S2991 }),
  .B({ S2992 }),
  .Y({ S2994 })
);
NAND #() 
NAND_1708_ (
  .A({ S1458 }),
  .B({ S2993 }),
  .Y({ S2995 })
);
NOR #() 
NOR_850_ (
  .A({ S2991 }),
  .B({ S2995 }),
  .Y({ S2996 })
);
NAND #() 
NAND_1709_ (
  .A({ S1458 }),
  .B({ S2994 }),
  .Y({ S2997 })
);
NAND #() 
NAND_1710_ (
  .A({ S2990 }),
  .B({ S2997 }),
  .Y({ S2998 })
);
NAND #() 
NAND_1711_ (
  .A({ S1444 }),
  .B({ S2998 }),
  .Y({ S2999 })
);
NAND #() 
NAND_1712_ (
  .A({ S2986 }),
  .B({ S2999 }),
  .Y({ S3000 })
);
NOR #() 
NOR_851_ (
  .A({ S1444 }),
  .B({ S2985 }),
  .Y({ S3001 })
);
NOR #() 
NOR_852_ (
  .A({ S1443 }),
  .B({ S2996 }),
  .Y({ S3002 })
);
NAND #() 
NAND_1713_ (
  .A({ S2990 }),
  .B({ S3002 }),
  .Y({ S3003 })
);
NAND #() 
NAND_1714_ (
  .A({ S1449 }),
  .B({ S3003 }),
  .Y({ S3004 })
);
NOR #() 
NOR_853_ (
  .A({ S3001 }),
  .B({ S3004 }),
  .Y({ S3005 })
);
NAND #() 
NAND_1715_ (
  .A({ S1449 }),
  .B({ S3000 }),
  .Y({ S3006 })
);
NOR #() 
NOR_854_ (
  .A({ datapath_theregisterfile_memtrf_78 }),
  .B({ S1438 }),
  .Y({ S3007 })
);
NAND #() 
NAND_1716_ (
  .A({ S7498 }),
  .B({ S1437 }),
  .Y({ S3008 })
);
NOR #() 
NOR_855_ (
  .A({ datapath_theregisterfile_memtrf_14 }),
  .B({ S1437 }),
  .Y({ S3009 })
);
NAND #() 
NAND_1717_ (
  .A({ S7542 }),
  .B({ S1438 }),
  .Y({ S3010 })
);
NOR #() 
NOR_856_ (
  .A({ S3007 }),
  .B({ S3009 }),
  .Y({ S3011 })
);
NAND #() 
NAND_1718_ (
  .A({ S3008 }),
  .B({ S3010 }),
  .Y({ S3012 })
);
NOR #() 
NOR_857_ (
  .A({ S1460 }),
  .B({ S3012 }),
  .Y({ S3013 })
);
NAND #() 
NAND_1719_ (
  .A({ S1459 }),
  .B({ S3011 }),
  .Y({ S3014 })
);
NAND #() 
NAND_1720_ (
  .A({ datapath_theregisterfile_memtrf_30 }),
  .B({ S1438 }),
  .Y({ S3015 })
);
NAND #() 
NAND_1721_ (
  .A({ datapath_theregisterfile_memtrf_94 }),
  .B({ S1437 }),
  .Y({ S3016 })
);
NAND #() 
NAND_1722_ (
  .A({ S3015 }),
  .B({ S3016 }),
  .Y({ S3017 })
);
NAND #() 
NAND_1723_ (
  .A({ S1926 }),
  .B({ S3017 }),
  .Y({ S3018 })
);
NAND #() 
NAND_1724_ (
  .A({ S3014 }),
  .B({ S3018 }),
  .Y({ S3019 })
);
NOT #() 
NOT_302_ (
  .A({ S3019 }),
  .Y({ S3020 })
);
NAND #() 
NAND_1725_ (
  .A({ S7509 }),
  .B({ S1438 }),
  .Y({ S3021 })
);
NOR #() 
NOR_858_ (
  .A({ datapath_theregisterfile_memtrf_126 }),
  .B({ S1438 }),
  .Y({ S3022 })
);
NOR #() 
NOR_859_ (
  .A({ S1458 }),
  .B({ S3022 }),
  .Y({ S3023 })
);
NAND #() 
NAND_1726_ (
  .A({ S3021 }),
  .B({ S3023 }),
  .Y({ S3024 })
);
NOR #() 
NOR_860_ (
  .A({ datapath_theregisterfile_memtrf_46 }),
  .B({ S1437 }),
  .Y({ S3025 })
);
NOR #() 
NOR_861_ (
  .A({ datapath_theregisterfile_memtrf_110 }),
  .B({ S1438 }),
  .Y({ S3026 })
);
NOR #() 
NOR_862_ (
  .A({ S3025 }),
  .B({ S3026 }),
  .Y({ S3027 })
);
NAND #() 
NAND_1727_ (
  .A({ S1458 }),
  .B({ S3027 }),
  .Y({ S3028 })
);
NAND #() 
NAND_1728_ (
  .A({ S3024 }),
  .B({ S3028 }),
  .Y({ S3029 })
);
NAND #() 
NAND_1729_ (
  .A({ S1487 }),
  .B({ S3029 }),
  .Y({ S3030 })
);
NAND #() 
NAND_1730_ (
  .A({ S3018 }),
  .B({ S3030 }),
  .Y({ S3031 })
);
NOR #() 
NOR_863_ (
  .A({ S3013 }),
  .B({ S3031 }),
  .Y({ S3032 })
);
NAND #() 
NAND_1731_ (
  .A({ S3020 }),
  .B({ S3030 }),
  .Y({ S3033 })
);
NOR #() 
NOR_864_ (
  .A({ S3005 }),
  .B({ S3033 }),
  .Y({ S3034 })
);
NAND #() 
NAND_1732_ (
  .A({ S3006 }),
  .B({ S3032 }),
  .Y({ S3035 })
);
NOR #() 
NOR_865_ (
  .A({ S1461 }),
  .B({ S3034 }),
  .Y({ S3036 })
);
NAND #() 
NAND_1733_ (
  .A({ S1462 }),
  .B({ S3035 }),
  .Y({ S3037 })
);
NAND #() 
NAND_1734_ (
  .A({ S1429 }),
  .B({ S3036 }),
  .Y({ S3038 })
);
NAND #() 
NAND_1735_ (
  .A({ S2369 }),
  .B({ S3038 }),
  .Y({ S3039 })
);
NOT #() 
NOT_303_ (
  .A({ S3039 }),
  .Y({ S3040 })
);
NAND #() 
NAND_1736_ (
  .A({ datapath_addsubunit_in1_14 }),
  .B({ S3040 }),
  .Y({ S3041 })
);
NOT #() 
NOT_304_ (
  .A({ S3041 }),
  .Y({ S3042 })
);
NAND #() 
NAND_1737_ (
  .A({ S492 }),
  .B({ S3039 }),
  .Y({ S3043 })
);
NOT #() 
NOT_305_ (
  .A({ S3043 }),
  .Y({ S3044 })
);
NOR #() 
NOR_866_ (
  .A({ S3042 }),
  .B({ S3044 }),
  .Y({ S3045 })
);
NOT #() 
NOT_306_ (
  .A({ S3045 }),
  .Y({ S3046 })
);
NOR #() 
NOR_867_ (
  .A({ S2925 }),
  .B({ S2931 }),
  .Y({ S3047 })
);
NOR #() 
NOR_868_ (
  .A({ S2927 }),
  .B({ S3047 }),
  .Y({ S3048 })
);
NAND #() 
NAND_1738_ (
  .A({ S3045 }),
  .B({ S3048 }),
  .Y({ S3049 })
);
NOR #() 
NOR_869_ (
  .A({ S3045 }),
  .B({ S3048 }),
  .Y({ S3050 })
);
NOR #() 
NOR_870_ (
  .A({ S1526 }),
  .B({ S3050 }),
  .Y({ S3051 })
);
NAND #() 
NAND_1739_ (
  .A({ S3049 }),
  .B({ S3051 }),
  .Y({ S3052 })
);
NAND #() 
NAND_1740_ (
  .A({ S2939 }),
  .B({ S2949 }),
  .Y({ S3053 })
);
NOR #() 
NOR_871_ (
  .A({ S2940 }),
  .B({ S3053 }),
  .Y({ S3054 })
);
NOR #() 
NOR_872_ (
  .A({ S3045 }),
  .B({ S3054 }),
  .Y({ S3055 })
);
NOT #() 
NOT_307_ (
  .A({ S3055 }),
  .Y({ S3056 })
);
NAND #() 
NAND_1741_ (
  .A({ S3045 }),
  .B({ S3054 }),
  .Y({ S3057 })
);
NAND #() 
NAND_1742_ (
  .A({ S1527 }),
  .B({ S3057 }),
  .Y({ S3058 })
);
NOR #() 
NOR_873_ (
  .A({ S3055 }),
  .B({ S3058 }),
  .Y({ S3059 })
);
NAND #() 
NAND_1743_ (
  .A({ datapath_addsubunit_in1_14 }),
  .B({ S3039 }),
  .Y({ S3060 })
);
NOR #() 
NOR_874_ (
  .A({ S1533 }),
  .B({ S3060 }),
  .Y({ S3061 })
);
NAND #() 
NAND_1744_ (
  .A({ datapath_shiftunit_2387_A }),
  .B({ S1614 }),
  .Y({ S3062 })
);
NAND #() 
NAND_1745_ (
  .A({ datapath_shiftunit_2691_A }),
  .B({ S1609 }),
  .Y({ S3063 })
);
NOR #() 
NOR_875_ (
  .A({ datapath_muxmem_in2_14 }),
  .B({ S1359 }),
  .Y({ S3064 })
);
NOT #() 
NOT_308_ (
  .A({ S3064 }),
  .Y({ S3065 })
);
NAND #() 
NAND_1746_ (
  .A({ S1360 }),
  .B({ S3065 }),
  .Y({ S3066 })
);
NOR #() 
NOR_876_ (
  .A({ S1623 }),
  .B({ S3066 }),
  .Y({ S3067 })
);
NOR #() 
NOR_877_ (
  .A({ controller_opcode_2 }),
  .B({ S1396 }),
  .Y({ S3068 })
);
NOR #() 
NOR_878_ (
  .A({ S2364 }),
  .B({ S3068 }),
  .Y({ S3069 })
);
NOR #() 
NOR_879_ (
  .A({ S2053 }),
  .B({ S3069 }),
  .Y({ S3070 })
);
NOR #() 
NOR_880_ (
  .A({ S1547 }),
  .B({ S3070 }),
  .Y({ S3071 })
);
NAND #() 
NAND_1747_ (
  .A({ datapath_multdivunit_outmdu2_14 }),
  .B({ S8570 }),
  .Y({ S3072 })
);
NAND #() 
NAND_1748_ (
  .A({ datapath_databusin_14 }),
  .B({ S1627 }),
  .Y({ S3073 })
);
NAND #() 
NAND_1749_ (
  .A({ datapath_multdivunit_outmdu1_14 }),
  .B({ S1377 }),
  .Y({ S3074 })
);
NAND #() 
NAND_1750_ (
  .A({ S3072 }),
  .B({ S3073 }),
  .Y({ S3075 })
);
NOR #() 
NOR_881_ (
  .A({ S3071 }),
  .B({ S3075 }),
  .Y({ S3076 })
);
NAND #() 
NAND_1751_ (
  .A({ S3074 }),
  .B({ S3076 }),
  .Y({ S3077 })
);
NOR #() 
NOR_882_ (
  .A({ S3067 }),
  .B({ S3077 }),
  .Y({ S3078 })
);
NAND #() 
NAND_1752_ (
  .A({ S3063 }),
  .B({ S3078 }),
  .Y({ S3079 })
);
NOT #() 
NOT_309_ (
  .A({ S3079 }),
  .Y({ S3080 })
);
NAND #() 
NAND_1753_ (
  .A({ S3062 }),
  .B({ S3080 }),
  .Y({ S3081 })
);
NOR #() 
NOR_883_ (
  .A({ S3061 }),
  .B({ S3081 }),
  .Y({ S3082 })
);
NOR #() 
NOR_884_ (
  .A({ S492 }),
  .B({ S2945 }),
  .Y({ S3083 })
);
NOR #() 
NOR_885_ (
  .A({ datapath_addsubunit_in1_14 }),
  .B({ S2946 }),
  .Y({ S3084 })
);
NOR #() 
NOR_886_ (
  .A({ S3083 }),
  .B({ S3084 }),
  .Y({ S3085 })
);
NAND #() 
NAND_1754_ (
  .A({ S1538 }),
  .B({ S3085 }),
  .Y({ S3086 })
);
NAND #() 
NAND_1755_ (
  .A({ S3082 }),
  .B({ S3086 }),
  .Y({ S3087 })
);
NOR #() 
NOR_887_ (
  .A({ S3059 }),
  .B({ S3087 }),
  .Y({ S3088 })
);
NAND #() 
NAND_1756_ (
  .A({ S3052 }),
  .B({ S3088 }),
  .Y({ datapath_indatatrf_14 })
);
NAND #() 
NAND_1757_ (
  .A({ datapath_indatatrf_14 }),
  .B({ S1688 }),
  .Y({ S3089 })
);
NAND #() 
NAND_1758_ (
  .A({ datapath_theregisterfile_memtrf_78 }),
  .B({ S1689 }),
  .Y({ S3090 })
);
NAND #() 
NAND_1759_ (
  .A({ S3089 }),
  .B({ S3090 }),
  .Y({ S18 })
);
NAND #() 
NAND_1760_ (
  .A({ datapath_theregisterfile_memtrf_159 }),
  .B({ S1438 }),
  .Y({ S3091 })
);
NAND #() 
NAND_1761_ (
  .A({ datapath_theregisterfile_memtrf_223 }),
  .B({ S1437 }),
  .Y({ S3092 })
);
NAND #() 
NAND_1762_ (
  .A({ S3091 }),
  .B({ S3092 }),
  .Y({ S3093 })
);
NAND #() 
NAND_1763_ (
  .A({ S1457 }),
  .B({ S3093 }),
  .Y({ S3094 })
);
NOR #() 
NOR_888_ (
  .A({ datapath_theregisterfile_memtrf_143 }),
  .B({ S1437 }),
  .Y({ S3095 })
);
NOR #() 
NOR_889_ (
  .A({ datapath_theregisterfile_memtrf_207 }),
  .B({ S1438 }),
  .Y({ S3096 })
);
NOR #() 
NOR_890_ (
  .A({ S3095 }),
  .B({ S3096 }),
  .Y({ S3097 })
);
NAND #() 
NAND_1764_ (
  .A({ S1458 }),
  .B({ S3097 }),
  .Y({ S3098 })
);
NAND #() 
NAND_1765_ (
  .A({ S3094 }),
  .B({ S3098 }),
  .Y({ S3099 })
);
NOR #() 
NOR_891_ (
  .A({ S1443 }),
  .B({ S3099 }),
  .Y({ S3100 })
);
NOR #() 
NOR_892_ (
  .A({ datapath_theregisterfile_memtrf_255 }),
  .B({ S1438 }),
  .Y({ S3101 })
);
NAND #() 
NAND_1766_ (
  .A({ S7662 }),
  .B({ S1438 }),
  .Y({ S3102 })
);
NAND #() 
NAND_1767_ (
  .A({ S1457 }),
  .B({ S3102 }),
  .Y({ S3103 })
);
NOR #() 
NOR_893_ (
  .A({ S3101 }),
  .B({ S3103 }),
  .Y({ S3104 })
);
NOR #() 
NOR_894_ (
  .A({ datapath_theregisterfile_memtrf_239 }),
  .B({ S1438 }),
  .Y({ S3105 })
);
NAND #() 
NAND_1768_ (
  .A({ S7574 }),
  .B({ S1438 }),
  .Y({ S3106 })
);
NAND #() 
NAND_1769_ (
  .A({ S1458 }),
  .B({ S3106 }),
  .Y({ S3107 })
);
NOR #() 
NOR_895_ (
  .A({ S3105 }),
  .B({ S3107 }),
  .Y({ S3108 })
);
NOR #() 
NOR_896_ (
  .A({ S3104 }),
  .B({ S3108 }),
  .Y({ S3109 })
);
NAND #() 
NAND_1770_ (
  .A({ S1443 }),
  .B({ S3109 }),
  .Y({ S3110 })
);
NAND #() 
NAND_1771_ (
  .A({ S1449 }),
  .B({ S3110 }),
  .Y({ S3111 })
);
NOR #() 
NOR_897_ (
  .A({ S1450 }),
  .B({ S3100 }),
  .Y({ S3112 })
);
NOR #() 
NOR_898_ (
  .A({ S3100 }),
  .B({ S3111 }),
  .Y({ S3113 })
);
NAND #() 
NAND_1772_ (
  .A({ S3110 }),
  .B({ S3112 }),
  .Y({ S3114 })
);
NAND #() 
NAND_1773_ (
  .A({ datapath_theregisterfile_memtrf_63 }),
  .B({ S1438 }),
  .Y({ S3115 })
);
NAND #() 
NAND_1774_ (
  .A({ datapath_theregisterfile_memtrf_127 }),
  .B({ S1437 }),
  .Y({ S3116 })
);
NAND #() 
NAND_1775_ (
  .A({ S3115 }),
  .B({ S3116 }),
  .Y({ S3117 })
);
NOR #() 
NOR_899_ (
  .A({ S1458 }),
  .B({ S3117 }),
  .Y({ S3118 })
);
NOR #() 
NOR_900_ (
  .A({ datapath_theregisterfile_memtrf_47 }),
  .B({ S1437 }),
  .Y({ S3119 })
);
NOR #() 
NOR_901_ (
  .A({ datapath_theregisterfile_memtrf_111 }),
  .B({ S1438 }),
  .Y({ S3120 })
);
NOR #() 
NOR_902_ (
  .A({ S3119 }),
  .B({ S3120 }),
  .Y({ S3121 })
);
NOR #() 
NOR_903_ (
  .A({ S1457 }),
  .B({ S3121 }),
  .Y({ S3122 })
);
NOR #() 
NOR_904_ (
  .A({ S3118 }),
  .B({ S3122 }),
  .Y({ S3123 })
);
NAND #() 
NAND_1776_ (
  .A({ S1487 }),
  .B({ S3123 }),
  .Y({ S3124 })
);
NAND #() 
NAND_1777_ (
  .A({ datapath_theregisterfile_memtrf_15 }),
  .B({ S1438 }),
  .Y({ S3125 })
);
NAND #() 
NAND_1778_ (
  .A({ datapath_theregisterfile_memtrf_79 }),
  .B({ S1437 }),
  .Y({ S3126 })
);
NAND #() 
NAND_1779_ (
  .A({ S3125 }),
  .B({ S3126 }),
  .Y({ S3127 })
);
NOT #() 
NOT_310_ (
  .A({ S3127 }),
  .Y({ S3128 })
);
NOR #() 
NOR_905_ (
  .A({ S1460 }),
  .B({ S3128 }),
  .Y({ S3129 })
);
NAND #() 
NAND_1780_ (
  .A({ datapath_theregisterfile_memtrf_31 }),
  .B({ S1438 }),
  .Y({ S3130 })
);
NAND #() 
NAND_1781_ (
  .A({ datapath_theregisterfile_memtrf_95 }),
  .B({ S1437 }),
  .Y({ S3131 })
);
NAND #() 
NAND_1782_ (
  .A({ S3130 }),
  .B({ S3131 }),
  .Y({ S3132 })
);
NAND #() 
NAND_1783_ (
  .A({ S1926 }),
  .B({ S3132 }),
  .Y({ S3133 })
);
NOT #() 
NOT_311_ (
  .A({ S3133 }),
  .Y({ S3134 })
);
NOR #() 
NOR_906_ (
  .A({ S3129 }),
  .B({ S3134 }),
  .Y({ S3135 })
);
NAND #() 
NAND_1784_ (
  .A({ S3124 }),
  .B({ S3133 }),
  .Y({ S3136 })
);
NOR #() 
NOR_907_ (
  .A({ S3129 }),
  .B({ S3136 }),
  .Y({ S3137 })
);
NAND #() 
NAND_1785_ (
  .A({ S3124 }),
  .B({ S3135 }),
  .Y({ S3138 })
);
NOR #() 
NOR_908_ (
  .A({ S3113 }),
  .B({ S3138 }),
  .Y({ S3139 })
);
NAND #() 
NAND_1786_ (
  .A({ S3114 }),
  .B({ S3137 }),
  .Y({ S3140 })
);
NOR #() 
NOR_909_ (
  .A({ S1461 }),
  .B({ S3139 }),
  .Y({ S3141 })
);
NAND #() 
NAND_1787_ (
  .A({ S1462 }),
  .B({ S3140 }),
  .Y({ S3142 })
);
NOR #() 
NOR_910_ (
  .A({ S1430 }),
  .B({ S3142 }),
  .Y({ S3143 })
);
NOR #() 
NOR_911_ (
  .A({ S2368 }),
  .B({ S3143 }),
  .Y({ S3144 })
);
NOT #() 
NOT_312_ (
  .A({ S3144 }),
  .Y({ S3145 })
);
NOR #() 
NOR_912_ (
  .A({ datapath_addsubunit_in1_15 }),
  .B({ S3144 }),
  .Y({ S3146 })
);
NOT #() 
NOT_313_ (
  .A({ S3146 }),
  .Y({ S3147 })
);
NOR #() 
NOR_913_ (
  .A({ S1304 }),
  .B({ S3145 }),
  .Y({ S3148 })
);
NOT #() 
NOT_314_ (
  .A({ S3148 }),
  .Y({ S3149 })
);
NAND #() 
NAND_1788_ (
  .A({ S3147 }),
  .B({ S3149 }),
  .Y({ S3150 })
);
NAND #() 
NAND_1789_ (
  .A({ S3041 }),
  .B({ S3049 }),
  .Y({ S3151 })
);
NOR #() 
NOR_914_ (
  .A({ S3150 }),
  .B({ S3151 }),
  .Y({ S3152 })
);
NOT #() 
NOT_315_ (
  .A({ S3152 }),
  .Y({ S3153 })
);
NAND #() 
NAND_1790_ (
  .A({ S3150 }),
  .B({ S3151 }),
  .Y({ S3154 })
);
NAND #() 
NAND_1791_ (
  .A({ S3153 }),
  .B({ S3154 }),
  .Y({ S3155 })
);
NAND #() 
NAND_1792_ (
  .A({ S1525 }),
  .B({ S3155 }),
  .Y({ S3156 })
);
NAND #() 
NAND_1793_ (
  .A({ S3056 }),
  .B({ S3060 }),
  .Y({ S3157 })
);
NAND #() 
NAND_1794_ (
  .A({ S3150 }),
  .B({ S3157 }),
  .Y({ S3158 })
);
NOR #() 
NOR_915_ (
  .A({ S3150 }),
  .B({ S3157 }),
  .Y({ S3159 })
);
NAND #() 
NAND_1795_ (
  .A({ S1527 }),
  .B({ S3158 }),
  .Y({ S3160 })
);
NOR #() 
NOR_916_ (
  .A({ S3159 }),
  .B({ S3160 }),
  .Y({ S3161 })
);
NAND #() 
NAND_1796_ (
  .A({ datapath_shiftunit_2405_A }),
  .B({ S1614 }),
  .Y({ S3162 })
);
NOT #() 
NOT_316_ (
  .A({ S3162 }),
  .Y({ S3163 })
);
NAND #() 
NAND_1797_ (
  .A({ datapath_shiftunit_2708_A }),
  .B({ S1609 }),
  .Y({ S3164 })
);
NAND #() 
NAND_1798_ (
  .A({ S1364 }),
  .B({ S1622 }),
  .Y({ S3165 })
);
NOR #() 
NOR_917_ (
  .A({ S2053 }),
  .B({ S2363 }),
  .Y({ S3166 })
);
NOR #() 
NOR_918_ (
  .A({ S1547 }),
  .B({ S3166 }),
  .Y({ S3167 })
);
NAND #() 
NAND_1799_ (
  .A({ datapath_databusin_15 }),
  .B({ S1627 }),
  .Y({ S3168 })
);
NAND #() 
NAND_1800_ (
  .A({ datapath_multdivunit_outmdu2_15 }),
  .B({ S8570 }),
  .Y({ S3169 })
);
NAND #() 
NAND_1801_ (
  .A({ datapath_multdivunit_outmdu1_15 }),
  .B({ S1377 }),
  .Y({ S3170 })
);
NAND #() 
NAND_1802_ (
  .A({ S3169 }),
  .B({ S3170 }),
  .Y({ S3171 })
);
NOT #() 
NOT_317_ (
  .A({ S3171 }),
  .Y({ S3172 })
);
NAND #() 
NAND_1803_ (
  .A({ S3168 }),
  .B({ S3172 }),
  .Y({ S3173 })
);
NOR #() 
NOR_919_ (
  .A({ S3167 }),
  .B({ S3173 }),
  .Y({ S3174 })
);
NAND #() 
NAND_1804_ (
  .A({ S3165 }),
  .B({ S3174 }),
  .Y({ S3175 })
);
NOR #() 
NOR_920_ (
  .A({ S3163 }),
  .B({ S3175 }),
  .Y({ S3176 })
);
NAND #() 
NAND_1805_ (
  .A({ S3164 }),
  .B({ S3176 }),
  .Y({ S3177 })
);
NAND #() 
NAND_1806_ (
  .A({ S1534 }),
  .B({ S3145 }),
  .Y({ S3178 })
);
NOR #() 
NOR_921_ (
  .A({ S1304 }),
  .B({ S3178 }),
  .Y({ S3179 })
);
NOR #() 
NOR_922_ (
  .A({ S3177 }),
  .B({ S3179 }),
  .Y({ S3180 })
);
NAND #() 
NAND_1807_ (
  .A({ S1304 }),
  .B({ S3084 }),
  .Y({ S3181 })
);
NOR #() 
NOR_923_ (
  .A({ S1304 }),
  .B({ S3084 }),
  .Y({ S3182 })
);
NOR #() 
NOR_924_ (
  .A({ S1539 }),
  .B({ S3182 }),
  .Y({ S3183 })
);
NAND #() 
NAND_1808_ (
  .A({ S3181 }),
  .B({ S3183 }),
  .Y({ S3184 })
);
NAND #() 
NAND_1809_ (
  .A({ S3180 }),
  .B({ S3184 }),
  .Y({ S3185 })
);
NOR #() 
NOR_925_ (
  .A({ S3161 }),
  .B({ S3185 }),
  .Y({ S3186 })
);
NAND #() 
NAND_1810_ (
  .A({ S3156 }),
  .B({ S3186 }),
  .Y({ datapath_indatatrf_15 })
);
NAND #() 
NAND_1811_ (
  .A({ datapath_indatatrf_15 }),
  .B({ S1688 }),
  .Y({ S3187 })
);
NAND #() 
NAND_1812_ (
  .A({ datapath_theregisterfile_memtrf_79 }),
  .B({ S1689 }),
  .Y({ S3188 })
);
NAND #() 
NAND_1813_ (
  .A({ S3187 }),
  .B({ S3188 }),
  .Y({ S19 })
);
NOR #() 
NOR_926_ (
  .A({ S1655 }),
  .B({ S1662 }),
  .Y({ S3189 })
);
NAND #() 
NAND_1814_ (
  .A({ S1654 }),
  .B({ S1661 }),
  .Y({ S3190 })
);
NOR #() 
NOR_927_ (
  .A({ S1671 }),
  .B({ S1687 }),
  .Y({ S3191 })
);
NAND #() 
NAND_1815_ (
  .A({ S1672 }),
  .B({ S1686 }),
  .Y({ S3192 })
);
NOR #() 
NOR_928_ (
  .A({ S3190 }),
  .B({ S3192 }),
  .Y({ S3193 })
);
NAND #() 
NAND_1816_ (
  .A({ S3189 }),
  .B({ S3191 }),
  .Y({ S3194 })
);
NAND #() 
NAND_1817_ (
  .A({ datapath_indatatrf_0 }),
  .B({ S3193 }),
  .Y({ S3195 })
);
NAND #() 
NAND_1818_ (
  .A({ datapath_theregisterfile_memtrf_32 }),
  .B({ S3194 }),
  .Y({ S3196 })
);
NAND #() 
NAND_1819_ (
  .A({ S3195 }),
  .B({ S3196 }),
  .Y({ S20 })
);
NAND #() 
NAND_1820_ (
  .A({ datapath_indatatrf_1 }),
  .B({ S3193 }),
  .Y({ S3197 })
);
NAND #() 
NAND_1821_ (
  .A({ datapath_theregisterfile_memtrf_33 }),
  .B({ S3194 }),
  .Y({ S3198 })
);
NAND #() 
NAND_1822_ (
  .A({ S3197 }),
  .B({ S3198 }),
  .Y({ S21 })
);
NAND #() 
NAND_1823_ (
  .A({ datapath_indatatrf_2 }),
  .B({ S3193 }),
  .Y({ S3199 })
);
NAND #() 
NAND_1824_ (
  .A({ datapath_theregisterfile_memtrf_34 }),
  .B({ S3194 }),
  .Y({ S3200 })
);
NAND #() 
NAND_1825_ (
  .A({ S3199 }),
  .B({ S3200 }),
  .Y({ S22 })
);
NAND #() 
NAND_1826_ (
  .A({ datapath_indatatrf_3 }),
  .B({ S3193 }),
  .Y({ S3201 })
);
NAND #() 
NAND_1827_ (
  .A({ datapath_theregisterfile_memtrf_35 }),
  .B({ S3194 }),
  .Y({ S3202 })
);
NAND #() 
NAND_1828_ (
  .A({ S3201 }),
  .B({ S3202 }),
  .Y({ S23 })
);
NAND #() 
NAND_1829_ (
  .A({ datapath_indatatrf_4 }),
  .B({ S3193 }),
  .Y({ S3203 })
);
NAND #() 
NAND_1830_ (
  .A({ datapath_theregisterfile_memtrf_36 }),
  .B({ S3194 }),
  .Y({ S3204 })
);
NAND #() 
NAND_1831_ (
  .A({ S3203 }),
  .B({ S3204 }),
  .Y({ S24 })
);
NAND #() 
NAND_1832_ (
  .A({ datapath_indatatrf_5 }),
  .B({ S3193 }),
  .Y({ S3205 })
);
NAND #() 
NAND_1833_ (
  .A({ datapath_theregisterfile_memtrf_37 }),
  .B({ S3194 }),
  .Y({ S3206 })
);
NAND #() 
NAND_1834_ (
  .A({ S3205 }),
  .B({ S3206 }),
  .Y({ S25 })
);
NAND #() 
NAND_1835_ (
  .A({ datapath_indatatrf_6 }),
  .B({ S3193 }),
  .Y({ S3207 })
);
NAND #() 
NAND_1836_ (
  .A({ datapath_theregisterfile_memtrf_38 }),
  .B({ S3194 }),
  .Y({ S3208 })
);
NAND #() 
NAND_1837_ (
  .A({ S3207 }),
  .B({ S3208 }),
  .Y({ S26 })
);
NAND #() 
NAND_1838_ (
  .A({ datapath_indatatrf_7 }),
  .B({ S3193 }),
  .Y({ S3209 })
);
NAND #() 
NAND_1839_ (
  .A({ datapath_theregisterfile_memtrf_39 }),
  .B({ S3194 }),
  .Y({ S3210 })
);
NAND #() 
NAND_1840_ (
  .A({ S3209 }),
  .B({ S3210 }),
  .Y({ S27 })
);
NAND #() 
NAND_1841_ (
  .A({ datapath_indatatrf_8 }),
  .B({ S3193 }),
  .Y({ S3211 })
);
NAND #() 
NAND_1842_ (
  .A({ datapath_theregisterfile_memtrf_40 }),
  .B({ S3194 }),
  .Y({ S3212 })
);
NAND #() 
NAND_1843_ (
  .A({ S3211 }),
  .B({ S3212 }),
  .Y({ S28 })
);
NAND #() 
NAND_1844_ (
  .A({ datapath_indatatrf_9 }),
  .B({ S3193 }),
  .Y({ S3213 })
);
NAND #() 
NAND_1845_ (
  .A({ datapath_theregisterfile_memtrf_41 }),
  .B({ S3194 }),
  .Y({ S3214 })
);
NAND #() 
NAND_1846_ (
  .A({ S3213 }),
  .B({ S3214 }),
  .Y({ S29 })
);
NAND #() 
NAND_1847_ (
  .A({ datapath_indatatrf_10 }),
  .B({ S3193 }),
  .Y({ S3215 })
);
NAND #() 
NAND_1848_ (
  .A({ datapath_theregisterfile_memtrf_42 }),
  .B({ S3194 }),
  .Y({ S3216 })
);
NAND #() 
NAND_1849_ (
  .A({ S3215 }),
  .B({ S3216 }),
  .Y({ S30 })
);
NAND #() 
NAND_1850_ (
  .A({ datapath_indatatrf_11 }),
  .B({ S3193 }),
  .Y({ S3217 })
);
NAND #() 
NAND_1851_ (
  .A({ datapath_theregisterfile_memtrf_43 }),
  .B({ S3194 }),
  .Y({ S3218 })
);
NAND #() 
NAND_1852_ (
  .A({ S3217 }),
  .B({ S3218 }),
  .Y({ S31 })
);
NAND #() 
NAND_1853_ (
  .A({ datapath_indatatrf_12 }),
  .B({ S3193 }),
  .Y({ S3219 })
);
NAND #() 
NAND_1854_ (
  .A({ datapath_theregisterfile_memtrf_44 }),
  .B({ S3194 }),
  .Y({ S3220 })
);
NAND #() 
NAND_1855_ (
  .A({ S3219 }),
  .B({ S3220 }),
  .Y({ S32 })
);
NAND #() 
NAND_1856_ (
  .A({ datapath_indatatrf_13 }),
  .B({ S3193 }),
  .Y({ S3221 })
);
NAND #() 
NAND_1857_ (
  .A({ datapath_theregisterfile_memtrf_45 }),
  .B({ S3194 }),
  .Y({ S3222 })
);
NAND #() 
NAND_1858_ (
  .A({ S3221 }),
  .B({ S3222 }),
  .Y({ S33 })
);
NAND #() 
NAND_1859_ (
  .A({ datapath_indatatrf_14 }),
  .B({ S3193 }),
  .Y({ S3223 })
);
NAND #() 
NAND_1860_ (
  .A({ datapath_theregisterfile_memtrf_46 }),
  .B({ S3194 }),
  .Y({ S3224 })
);
NAND #() 
NAND_1861_ (
  .A({ S3223 }),
  .B({ S3224 }),
  .Y({ S34 })
);
NAND #() 
NAND_1862_ (
  .A({ datapath_indatatrf_15 }),
  .B({ S3193 }),
  .Y({ S3225 })
);
NAND #() 
NAND_1863_ (
  .A({ datapath_theregisterfile_memtrf_47 }),
  .B({ S3194 }),
  .Y({ S3226 })
);
NAND #() 
NAND_1864_ (
  .A({ S3225 }),
  .B({ S3226 }),
  .Y({ S35 })
);
NOR #() 
NOR_929_ (
  .A({ S1678 }),
  .B({ S1685 }),
  .Y({ S3227 })
);
NAND #() 
NAND_1865_ (
  .A({ S1679 }),
  .B({ S1684 }),
  .Y({ S3228 })
);
NOR #() 
NOR_930_ (
  .A({ S1671 }),
  .B({ S3228 }),
  .Y({ S3229 })
);
NAND #() 
NAND_1866_ (
  .A({ S1672 }),
  .B({ S3227 }),
  .Y({ S3230 })
);
NOR #() 
NOR_931_ (
  .A({ S3190 }),
  .B({ S3230 }),
  .Y({ S3231 })
);
NAND #() 
NAND_1867_ (
  .A({ S3189 }),
  .B({ S3229 }),
  .Y({ S3232 })
);
NAND #() 
NAND_1868_ (
  .A({ datapath_indatatrf_0 }),
  .B({ S3231 }),
  .Y({ S3233 })
);
NAND #() 
NAND_1869_ (
  .A({ datapath_theregisterfile_memtrf_48 }),
  .B({ S3232 }),
  .Y({ S3234 })
);
NAND #() 
NAND_1870_ (
  .A({ S3233 }),
  .B({ S3234 }),
  .Y({ S36 })
);
NAND #() 
NAND_1871_ (
  .A({ datapath_indatatrf_1 }),
  .B({ S3231 }),
  .Y({ S3235 })
);
NAND #() 
NAND_1872_ (
  .A({ datapath_theregisterfile_memtrf_49 }),
  .B({ S3232 }),
  .Y({ S3236 })
);
NAND #() 
NAND_1873_ (
  .A({ S3235 }),
  .B({ S3236 }),
  .Y({ S37 })
);
NAND #() 
NAND_1874_ (
  .A({ datapath_indatatrf_2 }),
  .B({ S3231 }),
  .Y({ S3237 })
);
NAND #() 
NAND_1875_ (
  .A({ datapath_theregisterfile_memtrf_50 }),
  .B({ S3232 }),
  .Y({ S3238 })
);
NAND #() 
NAND_1876_ (
  .A({ S3237 }),
  .B({ S3238 }),
  .Y({ S38 })
);
NAND #() 
NAND_1877_ (
  .A({ datapath_indatatrf_3 }),
  .B({ S3231 }),
  .Y({ S3239 })
);
NAND #() 
NAND_1878_ (
  .A({ datapath_theregisterfile_memtrf_51 }),
  .B({ S3232 }),
  .Y({ S3240 })
);
NAND #() 
NAND_1879_ (
  .A({ S3239 }),
  .B({ S3240 }),
  .Y({ S39 })
);
NAND #() 
NAND_1880_ (
  .A({ datapath_indatatrf_4 }),
  .B({ S3231 }),
  .Y({ S3241 })
);
NAND #() 
NAND_1881_ (
  .A({ datapath_theregisterfile_memtrf_52 }),
  .B({ S3232 }),
  .Y({ S3242 })
);
NAND #() 
NAND_1882_ (
  .A({ S3241 }),
  .B({ S3242 }),
  .Y({ S40 })
);
NAND #() 
NAND_1883_ (
  .A({ datapath_indatatrf_5 }),
  .B({ S3231 }),
  .Y({ S3243 })
);
NAND #() 
NAND_1884_ (
  .A({ datapath_theregisterfile_memtrf_53 }),
  .B({ S3232 }),
  .Y({ S3244 })
);
NAND #() 
NAND_1885_ (
  .A({ S3243 }),
  .B({ S3244 }),
  .Y({ S41 })
);
NAND #() 
NAND_1886_ (
  .A({ datapath_indatatrf_6 }),
  .B({ S3231 }),
  .Y({ S3245 })
);
NAND #() 
NAND_1887_ (
  .A({ datapath_theregisterfile_memtrf_54 }),
  .B({ S3232 }),
  .Y({ S3246 })
);
NAND #() 
NAND_1888_ (
  .A({ S3245 }),
  .B({ S3246 }),
  .Y({ S42 })
);
NAND #() 
NAND_1889_ (
  .A({ datapath_indatatrf_7 }),
  .B({ S3231 }),
  .Y({ S3247 })
);
NAND #() 
NAND_1890_ (
  .A({ datapath_theregisterfile_memtrf_55 }),
  .B({ S3232 }),
  .Y({ S3248 })
);
NAND #() 
NAND_1891_ (
  .A({ S3247 }),
  .B({ S3248 }),
  .Y({ S43 })
);
NAND #() 
NAND_1892_ (
  .A({ datapath_indatatrf_8 }),
  .B({ S3231 }),
  .Y({ S3249 })
);
NAND #() 
NAND_1893_ (
  .A({ datapath_theregisterfile_memtrf_56 }),
  .B({ S3232 }),
  .Y({ S3250 })
);
NAND #() 
NAND_1894_ (
  .A({ S3249 }),
  .B({ S3250 }),
  .Y({ S44 })
);
NAND #() 
NAND_1895_ (
  .A({ datapath_indatatrf_9 }),
  .B({ S3231 }),
  .Y({ S3251 })
);
NAND #() 
NAND_1896_ (
  .A({ datapath_theregisterfile_memtrf_57 }),
  .B({ S3232 }),
  .Y({ S3252 })
);
NAND #() 
NAND_1897_ (
  .A({ S3251 }),
  .B({ S3252 }),
  .Y({ S45 })
);
NAND #() 
NAND_1898_ (
  .A({ datapath_indatatrf_10 }),
  .B({ S3231 }),
  .Y({ S3253 })
);
NAND #() 
NAND_1899_ (
  .A({ datapath_theregisterfile_memtrf_58 }),
  .B({ S3232 }),
  .Y({ S3254 })
);
NAND #() 
NAND_1900_ (
  .A({ S3253 }),
  .B({ S3254 }),
  .Y({ S46 })
);
NAND #() 
NAND_1901_ (
  .A({ datapath_indatatrf_11 }),
  .B({ S3231 }),
  .Y({ S3255 })
);
NAND #() 
NAND_1902_ (
  .A({ datapath_theregisterfile_memtrf_59 }),
  .B({ S3232 }),
  .Y({ S3256 })
);
NAND #() 
NAND_1903_ (
  .A({ S3255 }),
  .B({ S3256 }),
  .Y({ S47 })
);
NAND #() 
NAND_1904_ (
  .A({ datapath_indatatrf_12 }),
  .B({ S3231 }),
  .Y({ S3257 })
);
NAND #() 
NAND_1905_ (
  .A({ datapath_theregisterfile_memtrf_60 }),
  .B({ S3232 }),
  .Y({ S3258 })
);
NAND #() 
NAND_1906_ (
  .A({ S3257 }),
  .B({ S3258 }),
  .Y({ S48 })
);
NAND #() 
NAND_1907_ (
  .A({ datapath_indatatrf_13 }),
  .B({ S3231 }),
  .Y({ S3259 })
);
NAND #() 
NAND_1908_ (
  .A({ datapath_theregisterfile_memtrf_61 }),
  .B({ S3232 }),
  .Y({ S3260 })
);
NAND #() 
NAND_1909_ (
  .A({ S3259 }),
  .B({ S3260 }),
  .Y({ S49 })
);
NAND #() 
NAND_1910_ (
  .A({ datapath_indatatrf_14 }),
  .B({ S3231 }),
  .Y({ S3261 })
);
NAND #() 
NAND_1911_ (
  .A({ datapath_theregisterfile_memtrf_62 }),
  .B({ S3232 }),
  .Y({ S3262 })
);
NAND #() 
NAND_1912_ (
  .A({ S3261 }),
  .B({ S3262 }),
  .Y({ S50 })
);
NAND #() 
NAND_1913_ (
  .A({ datapath_indatatrf_15 }),
  .B({ S3231 }),
  .Y({ S3263 })
);
NAND #() 
NAND_1914_ (
  .A({ datapath_theregisterfile_memtrf_63 }),
  .B({ S3232 }),
  .Y({ S3264 })
);
NAND #() 
NAND_1915_ (
  .A({ S3263 }),
  .B({ S3264 }),
  .Y({ S51 })
);
NOR #() 
NOR_932_ (
  .A({ S1655 }),
  .B({ S1661 }),
  .Y({ S3265 })
);
NAND #() 
NAND_1916_ (
  .A({ S1654 }),
  .B({ S1662 }),
  .Y({ S3266 })
);
NOR #() 
NOR_933_ (
  .A({ S1672 }),
  .B({ S3266 }),
  .Y({ S3267 })
);
NAND #() 
NAND_1917_ (
  .A({ S1671 }),
  .B({ S3265 }),
  .Y({ S3268 })
);
NOR #() 
NOR_934_ (
  .A({ S1687 }),
  .B({ S3268 }),
  .Y({ S3269 })
);
NAND #() 
NAND_1918_ (
  .A({ S1686 }),
  .B({ S3267 }),
  .Y({ S3270 })
);
NAND #() 
NAND_1919_ (
  .A({ datapath_indatatrf_0 }),
  .B({ S3269 }),
  .Y({ S3271 })
);
NAND #() 
NAND_1920_ (
  .A({ datapath_theregisterfile_memtrf_128 }),
  .B({ S3270 }),
  .Y({ S3272 })
);
NAND #() 
NAND_1921_ (
  .A({ S3271 }),
  .B({ S3272 }),
  .Y({ S52 })
);
NAND #() 
NAND_1922_ (
  .A({ datapath_indatatrf_1 }),
  .B({ S3269 }),
  .Y({ S3273 })
);
NAND #() 
NAND_1923_ (
  .A({ datapath_theregisterfile_memtrf_129 }),
  .B({ S3270 }),
  .Y({ S3274 })
);
NAND #() 
NAND_1924_ (
  .A({ S3273 }),
  .B({ S3274 }),
  .Y({ S53 })
);
NAND #() 
NAND_1925_ (
  .A({ datapath_indatatrf_2 }),
  .B({ S3269 }),
  .Y({ S3275 })
);
NAND #() 
NAND_1926_ (
  .A({ datapath_theregisterfile_memtrf_130 }),
  .B({ S3270 }),
  .Y({ S3276 })
);
NAND #() 
NAND_1927_ (
  .A({ S3275 }),
  .B({ S3276 }),
  .Y({ S54 })
);
NAND #() 
NAND_1928_ (
  .A({ datapath_indatatrf_3 }),
  .B({ S3269 }),
  .Y({ S3277 })
);
NAND #() 
NAND_1929_ (
  .A({ datapath_theregisterfile_memtrf_131 }),
  .B({ S3270 }),
  .Y({ S3278 })
);
NAND #() 
NAND_1930_ (
  .A({ S3277 }),
  .B({ S3278 }),
  .Y({ S55 })
);
NAND #() 
NAND_1931_ (
  .A({ datapath_indatatrf_4 }),
  .B({ S3269 }),
  .Y({ S3279 })
);
NAND #() 
NAND_1932_ (
  .A({ datapath_theregisterfile_memtrf_132 }),
  .B({ S3270 }),
  .Y({ S3280 })
);
NAND #() 
NAND_1933_ (
  .A({ S3279 }),
  .B({ S3280 }),
  .Y({ S56 })
);
NAND #() 
NAND_1934_ (
  .A({ datapath_indatatrf_5 }),
  .B({ S3269 }),
  .Y({ S3281 })
);
NAND #() 
NAND_1935_ (
  .A({ datapath_theregisterfile_memtrf_133 }),
  .B({ S3270 }),
  .Y({ S3282 })
);
NAND #() 
NAND_1936_ (
  .A({ S3281 }),
  .B({ S3282 }),
  .Y({ S57 })
);
NAND #() 
NAND_1937_ (
  .A({ datapath_indatatrf_6 }),
  .B({ S3269 }),
  .Y({ S3283 })
);
NAND #() 
NAND_1938_ (
  .A({ datapath_theregisterfile_memtrf_134 }),
  .B({ S3270 }),
  .Y({ S3284 })
);
NAND #() 
NAND_1939_ (
  .A({ S3283 }),
  .B({ S3284 }),
  .Y({ S58 })
);
NAND #() 
NAND_1940_ (
  .A({ datapath_indatatrf_7 }),
  .B({ S3269 }),
  .Y({ S3285 })
);
NAND #() 
NAND_1941_ (
  .A({ datapath_theregisterfile_memtrf_135 }),
  .B({ S3270 }),
  .Y({ S3286 })
);
NAND #() 
NAND_1942_ (
  .A({ S3285 }),
  .B({ S3286 }),
  .Y({ S59 })
);
NAND #() 
NAND_1943_ (
  .A({ datapath_indatatrf_8 }),
  .B({ S3269 }),
  .Y({ S3287 })
);
NAND #() 
NAND_1944_ (
  .A({ datapath_theregisterfile_memtrf_136 }),
  .B({ S3270 }),
  .Y({ S3288 })
);
NAND #() 
NAND_1945_ (
  .A({ S3287 }),
  .B({ S3288 }),
  .Y({ S60 })
);
NAND #() 
NAND_1946_ (
  .A({ datapath_indatatrf_9 }),
  .B({ S3269 }),
  .Y({ S3289 })
);
NAND #() 
NAND_1947_ (
  .A({ datapath_theregisterfile_memtrf_137 }),
  .B({ S3270 }),
  .Y({ S3290 })
);
NAND #() 
NAND_1948_ (
  .A({ S3289 }),
  .B({ S3290 }),
  .Y({ S61 })
);
NAND #() 
NAND_1949_ (
  .A({ datapath_indatatrf_10 }),
  .B({ S3269 }),
  .Y({ S3291 })
);
NAND #() 
NAND_1950_ (
  .A({ datapath_theregisterfile_memtrf_138 }),
  .B({ S3270 }),
  .Y({ S3292 })
);
NAND #() 
NAND_1951_ (
  .A({ S3291 }),
  .B({ S3292 }),
  .Y({ S62 })
);
NAND #() 
NAND_1952_ (
  .A({ datapath_indatatrf_11 }),
  .B({ S3269 }),
  .Y({ S3293 })
);
NAND #() 
NAND_1953_ (
  .A({ datapath_theregisterfile_memtrf_139 }),
  .B({ S3270 }),
  .Y({ S3294 })
);
NAND #() 
NAND_1954_ (
  .A({ S3293 }),
  .B({ S3294 }),
  .Y({ S63 })
);
NAND #() 
NAND_1955_ (
  .A({ datapath_indatatrf_12 }),
  .B({ S3269 }),
  .Y({ S3295 })
);
NAND #() 
NAND_1956_ (
  .A({ datapath_theregisterfile_memtrf_140 }),
  .B({ S3270 }),
  .Y({ S3296 })
);
NAND #() 
NAND_1957_ (
  .A({ S3295 }),
  .B({ S3296 }),
  .Y({ S64 })
);
NAND #() 
NAND_1958_ (
  .A({ datapath_indatatrf_13 }),
  .B({ S3269 }),
  .Y({ S3297 })
);
NAND #() 
NAND_1959_ (
  .A({ datapath_theregisterfile_memtrf_141 }),
  .B({ S3270 }),
  .Y({ S3298 })
);
NAND #() 
NAND_1960_ (
  .A({ S3297 }),
  .B({ S3298 }),
  .Y({ S65 })
);
NAND #() 
NAND_1961_ (
  .A({ datapath_indatatrf_14 }),
  .B({ S3269 }),
  .Y({ S3299 })
);
NAND #() 
NAND_1962_ (
  .A({ datapath_theregisterfile_memtrf_142 }),
  .B({ S3270 }),
  .Y({ S3300 })
);
NAND #() 
NAND_1963_ (
  .A({ S3299 }),
  .B({ S3300 }),
  .Y({ S66 })
);
NAND #() 
NAND_1964_ (
  .A({ datapath_indatatrf_15 }),
  .B({ S3269 }),
  .Y({ S3301 })
);
NAND #() 
NAND_1965_ (
  .A({ datapath_theregisterfile_memtrf_143 }),
  .B({ S3270 }),
  .Y({ S3302 })
);
NAND #() 
NAND_1966_ (
  .A({ S3301 }),
  .B({ S3302 }),
  .Y({ S67 })
);
NOR #() 
NOR_935_ (
  .A({ S1672 }),
  .B({ S3190 }),
  .Y({ S3303 })
);
NAND #() 
NAND_1967_ (
  .A({ S1671 }),
  .B({ S3189 }),
  .Y({ S3304 })
);
NOR #() 
NOR_936_ (
  .A({ S3228 }),
  .B({ S3304 }),
  .Y({ S3305 })
);
NAND #() 
NAND_1968_ (
  .A({ S3227 }),
  .B({ S3303 }),
  .Y({ S3306 })
);
NAND #() 
NAND_1969_ (
  .A({ datapath_indatatrf_0 }),
  .B({ S3305 }),
  .Y({ S3307 })
);
NAND #() 
NAND_1970_ (
  .A({ datapath_theregisterfile_memtrf_16 }),
  .B({ S3306 }),
  .Y({ S3308 })
);
NAND #() 
NAND_1971_ (
  .A({ S3307 }),
  .B({ S3308 }),
  .Y({ S68 })
);
NAND #() 
NAND_1972_ (
  .A({ datapath_indatatrf_1 }),
  .B({ S3305 }),
  .Y({ S3309 })
);
NAND #() 
NAND_1973_ (
  .A({ datapath_theregisterfile_memtrf_17 }),
  .B({ S3306 }),
  .Y({ S3310 })
);
NAND #() 
NAND_1974_ (
  .A({ S3309 }),
  .B({ S3310 }),
  .Y({ S69 })
);
NAND #() 
NAND_1975_ (
  .A({ datapath_indatatrf_2 }),
  .B({ S3305 }),
  .Y({ S3311 })
);
NAND #() 
NAND_1976_ (
  .A({ datapath_theregisterfile_memtrf_18 }),
  .B({ S3306 }),
  .Y({ S3312 })
);
NAND #() 
NAND_1977_ (
  .A({ S3311 }),
  .B({ S3312 }),
  .Y({ S70 })
);
NAND #() 
NAND_1978_ (
  .A({ datapath_indatatrf_3 }),
  .B({ S3305 }),
  .Y({ S3313 })
);
NAND #() 
NAND_1979_ (
  .A({ datapath_theregisterfile_memtrf_19 }),
  .B({ S3306 }),
  .Y({ S3314 })
);
NAND #() 
NAND_1980_ (
  .A({ S3313 }),
  .B({ S3314 }),
  .Y({ S71 })
);
NAND #() 
NAND_1981_ (
  .A({ datapath_indatatrf_4 }),
  .B({ S3305 }),
  .Y({ S3315 })
);
NAND #() 
NAND_1982_ (
  .A({ datapath_theregisterfile_memtrf_20 }),
  .B({ S3306 }),
  .Y({ S3316 })
);
NAND #() 
NAND_1983_ (
  .A({ S3315 }),
  .B({ S3316 }),
  .Y({ S72 })
);
NAND #() 
NAND_1984_ (
  .A({ datapath_indatatrf_5 }),
  .B({ S3305 }),
  .Y({ S3317 })
);
NAND #() 
NAND_1985_ (
  .A({ datapath_theregisterfile_memtrf_21 }),
  .B({ S3306 }),
  .Y({ S3318 })
);
NAND #() 
NAND_1986_ (
  .A({ S3317 }),
  .B({ S3318 }),
  .Y({ S73 })
);
NAND #() 
NAND_1987_ (
  .A({ datapath_indatatrf_6 }),
  .B({ S3305 }),
  .Y({ S3319 })
);
NAND #() 
NAND_1988_ (
  .A({ datapath_theregisterfile_memtrf_22 }),
  .B({ S3306 }),
  .Y({ S3320 })
);
NAND #() 
NAND_1989_ (
  .A({ S3319 }),
  .B({ S3320 }),
  .Y({ S74 })
);
NAND #() 
NAND_1990_ (
  .A({ datapath_indatatrf_7 }),
  .B({ S3305 }),
  .Y({ S3321 })
);
NAND #() 
NAND_1991_ (
  .A({ datapath_theregisterfile_memtrf_23 }),
  .B({ S3306 }),
  .Y({ S3322 })
);
NAND #() 
NAND_1992_ (
  .A({ S3321 }),
  .B({ S3322 }),
  .Y({ S75 })
);
NAND #() 
NAND_1993_ (
  .A({ datapath_indatatrf_8 }),
  .B({ S3305 }),
  .Y({ S3323 })
);
NAND #() 
NAND_1994_ (
  .A({ datapath_theregisterfile_memtrf_24 }),
  .B({ S3306 }),
  .Y({ S3324 })
);
NAND #() 
NAND_1995_ (
  .A({ S3323 }),
  .B({ S3324 }),
  .Y({ S76 })
);
NAND #() 
NAND_1996_ (
  .A({ datapath_indatatrf_9 }),
  .B({ S3305 }),
  .Y({ S3325 })
);
NAND #() 
NAND_1997_ (
  .A({ datapath_theregisterfile_memtrf_25 }),
  .B({ S3306 }),
  .Y({ S3326 })
);
NAND #() 
NAND_1998_ (
  .A({ S3325 }),
  .B({ S3326 }),
  .Y({ S77 })
);
NAND #() 
NAND_1999_ (
  .A({ datapath_indatatrf_10 }),
  .B({ S3305 }),
  .Y({ S3327 })
);
NAND #() 
NAND_2000_ (
  .A({ datapath_theregisterfile_memtrf_26 }),
  .B({ S3306 }),
  .Y({ S3328 })
);
NAND #() 
NAND_2001_ (
  .A({ S3327 }),
  .B({ S3328 }),
  .Y({ S78 })
);
NAND #() 
NAND_2002_ (
  .A({ datapath_indatatrf_11 }),
  .B({ S3305 }),
  .Y({ S3329 })
);
NAND #() 
NAND_2003_ (
  .A({ datapath_theregisterfile_memtrf_27 }),
  .B({ S3306 }),
  .Y({ S3330 })
);
NAND #() 
NAND_2004_ (
  .A({ S3329 }),
  .B({ S3330 }),
  .Y({ S79 })
);
NAND #() 
NAND_2005_ (
  .A({ datapath_indatatrf_12 }),
  .B({ S3305 }),
  .Y({ S3331 })
);
NAND #() 
NAND_2006_ (
  .A({ datapath_theregisterfile_memtrf_28 }),
  .B({ S3306 }),
  .Y({ S3332 })
);
NAND #() 
NAND_2007_ (
  .A({ S3331 }),
  .B({ S3332 }),
  .Y({ S80 })
);
NAND #() 
NAND_2008_ (
  .A({ datapath_indatatrf_13 }),
  .B({ S3305 }),
  .Y({ S3333 })
);
NAND #() 
NAND_2009_ (
  .A({ datapath_theregisterfile_memtrf_29 }),
  .B({ S3306 }),
  .Y({ S3334 })
);
NAND #() 
NAND_2010_ (
  .A({ S3333 }),
  .B({ S3334 }),
  .Y({ S81 })
);
NAND #() 
NAND_2011_ (
  .A({ datapath_indatatrf_14 }),
  .B({ S3305 }),
  .Y({ S3335 })
);
NAND #() 
NAND_2012_ (
  .A({ datapath_theregisterfile_memtrf_30 }),
  .B({ S3306 }),
  .Y({ S3336 })
);
NAND #() 
NAND_2013_ (
  .A({ S3335 }),
  .B({ S3336 }),
  .Y({ S82 })
);
NAND #() 
NAND_2014_ (
  .A({ datapath_indatatrf_15 }),
  .B({ S3305 }),
  .Y({ S3337 })
);
NAND #() 
NAND_2015_ (
  .A({ datapath_theregisterfile_memtrf_31 }),
  .B({ S3306 }),
  .Y({ S3338 })
);
NAND #() 
NAND_2016_ (
  .A({ S3337 }),
  .B({ S3338 }),
  .Y({ S83 })
);
NOR #() 
NOR_937_ (
  .A({ S1674 }),
  .B({ S3228 }),
  .Y({ S3339 })
);
NAND #() 
NAND_2017_ (
  .A({ S1673 }),
  .B({ S3227 }),
  .Y({ S3340 })
);
NAND #() 
NAND_2018_ (
  .A({ datapath_indatatrf_0 }),
  .B({ S3339 }),
  .Y({ S3341 })
);
NAND #() 
NAND_2019_ (
  .A({ datapath_theregisterfile_memtrf_80 }),
  .B({ S3340 }),
  .Y({ S3342 })
);
NAND #() 
NAND_2020_ (
  .A({ S3341 }),
  .B({ S3342 }),
  .Y({ S84 })
);
NAND #() 
NAND_2021_ (
  .A({ datapath_indatatrf_1 }),
  .B({ S3339 }),
  .Y({ S3343 })
);
NAND #() 
NAND_2022_ (
  .A({ datapath_theregisterfile_memtrf_81 }),
  .B({ S3340 }),
  .Y({ S3344 })
);
NAND #() 
NAND_2023_ (
  .A({ S3343 }),
  .B({ S3344 }),
  .Y({ S85 })
);
NAND #() 
NAND_2024_ (
  .A({ datapath_indatatrf_2 }),
  .B({ S3339 }),
  .Y({ S3345 })
);
NAND #() 
NAND_2025_ (
  .A({ datapath_theregisterfile_memtrf_82 }),
  .B({ S3340 }),
  .Y({ S3346 })
);
NAND #() 
NAND_2026_ (
  .A({ S3345 }),
  .B({ S3346 }),
  .Y({ S86 })
);
NAND #() 
NAND_2027_ (
  .A({ datapath_indatatrf_3 }),
  .B({ S3339 }),
  .Y({ S3347 })
);
NAND #() 
NAND_2028_ (
  .A({ datapath_theregisterfile_memtrf_83 }),
  .B({ S3340 }),
  .Y({ S3348 })
);
NAND #() 
NAND_2029_ (
  .A({ S3347 }),
  .B({ S3348 }),
  .Y({ S87 })
);
NAND #() 
NAND_2030_ (
  .A({ datapath_indatatrf_4 }),
  .B({ S3339 }),
  .Y({ S3349 })
);
NAND #() 
NAND_2031_ (
  .A({ datapath_theregisterfile_memtrf_84 }),
  .B({ S3340 }),
  .Y({ S3350 })
);
NAND #() 
NAND_2032_ (
  .A({ S3349 }),
  .B({ S3350 }),
  .Y({ S88 })
);
NAND #() 
NAND_2033_ (
  .A({ datapath_indatatrf_5 }),
  .B({ S3339 }),
  .Y({ S3351 })
);
NAND #() 
NAND_2034_ (
  .A({ datapath_theregisterfile_memtrf_85 }),
  .B({ S3340 }),
  .Y({ S3352 })
);
NAND #() 
NAND_2035_ (
  .A({ S3351 }),
  .B({ S3352 }),
  .Y({ S89 })
);
NAND #() 
NAND_2036_ (
  .A({ datapath_indatatrf_6 }),
  .B({ S3339 }),
  .Y({ S3353 })
);
NAND #() 
NAND_2037_ (
  .A({ datapath_theregisterfile_memtrf_86 }),
  .B({ S3340 }),
  .Y({ S3354 })
);
NAND #() 
NAND_2038_ (
  .A({ S3353 }),
  .B({ S3354 }),
  .Y({ S90 })
);
NAND #() 
NAND_2039_ (
  .A({ datapath_indatatrf_7 }),
  .B({ S3339 }),
  .Y({ S3355 })
);
NAND #() 
NAND_2040_ (
  .A({ datapath_theregisterfile_memtrf_87 }),
  .B({ S3340 }),
  .Y({ S3356 })
);
NAND #() 
NAND_2041_ (
  .A({ S3355 }),
  .B({ S3356 }),
  .Y({ S91 })
);
NAND #() 
NAND_2042_ (
  .A({ datapath_indatatrf_8 }),
  .B({ S3339 }),
  .Y({ S3357 })
);
NAND #() 
NAND_2043_ (
  .A({ datapath_theregisterfile_memtrf_88 }),
  .B({ S3340 }),
  .Y({ S3358 })
);
NAND #() 
NAND_2044_ (
  .A({ S3357 }),
  .B({ S3358 }),
  .Y({ S92 })
);
NAND #() 
NAND_2045_ (
  .A({ datapath_indatatrf_9 }),
  .B({ S3339 }),
  .Y({ S3359 })
);
NAND #() 
NAND_2046_ (
  .A({ datapath_theregisterfile_memtrf_89 }),
  .B({ S3340 }),
  .Y({ S3360 })
);
NAND #() 
NAND_2047_ (
  .A({ S3359 }),
  .B({ S3360 }),
  .Y({ S93 })
);
NAND #() 
NAND_2048_ (
  .A({ datapath_indatatrf_10 }),
  .B({ S3339 }),
  .Y({ S3361 })
);
NAND #() 
NAND_2049_ (
  .A({ datapath_theregisterfile_memtrf_90 }),
  .B({ S3340 }),
  .Y({ S3362 })
);
NAND #() 
NAND_2050_ (
  .A({ S3361 }),
  .B({ S3362 }),
  .Y({ S94 })
);
NAND #() 
NAND_2051_ (
  .A({ datapath_indatatrf_11 }),
  .B({ S3339 }),
  .Y({ S3363 })
);
NAND #() 
NAND_2052_ (
  .A({ datapath_theregisterfile_memtrf_91 }),
  .B({ S3340 }),
  .Y({ S3364 })
);
NAND #() 
NAND_2053_ (
  .A({ S3363 }),
  .B({ S3364 }),
  .Y({ S95 })
);
NAND #() 
NAND_2054_ (
  .A({ datapath_indatatrf_12 }),
  .B({ S3339 }),
  .Y({ S3365 })
);
NAND #() 
NAND_2055_ (
  .A({ datapath_theregisterfile_memtrf_92 }),
  .B({ S3340 }),
  .Y({ S3366 })
);
NAND #() 
NAND_2056_ (
  .A({ S3365 }),
  .B({ S3366 }),
  .Y({ S96 })
);
NAND #() 
NAND_2057_ (
  .A({ datapath_indatatrf_13 }),
  .B({ S3339 }),
  .Y({ S3367 })
);
NAND #() 
NAND_2058_ (
  .A({ datapath_theregisterfile_memtrf_93 }),
  .B({ S3340 }),
  .Y({ S3368 })
);
NAND #() 
NAND_2059_ (
  .A({ S3367 }),
  .B({ S3368 }),
  .Y({ S97 })
);
NAND #() 
NAND_2060_ (
  .A({ datapath_indatatrf_14 }),
  .B({ S3339 }),
  .Y({ S3369 })
);
NAND #() 
NAND_2061_ (
  .A({ datapath_theregisterfile_memtrf_94 }),
  .B({ S3340 }),
  .Y({ S3370 })
);
NAND #() 
NAND_2062_ (
  .A({ S3369 }),
  .B({ S3370 }),
  .Y({ S98 })
);
NAND #() 
NAND_2063_ (
  .A({ datapath_indatatrf_15 }),
  .B({ S3339 }),
  .Y({ S3371 })
);
NAND #() 
NAND_2064_ (
  .A({ datapath_theregisterfile_memtrf_95 }),
  .B({ S3340 }),
  .Y({ S3372 })
);
NAND #() 
NAND_2065_ (
  .A({ S3371 }),
  .B({ S3372 }),
  .Y({ S99 })
);
NOR #() 
NOR_938_ (
  .A({ S1664 }),
  .B({ S3192 }),
  .Y({ S3373 })
);
NAND #() 
NAND_2066_ (
  .A({ S1663 }),
  .B({ S3191 }),
  .Y({ S3374 })
);
NAND #() 
NAND_2067_ (
  .A({ datapath_indatatrf_0 }),
  .B({ S3373 }),
  .Y({ S3375 })
);
NAND #() 
NAND_2068_ (
  .A({ datapath_theregisterfile_memtrf_96 }),
  .B({ S3374 }),
  .Y({ S3376 })
);
NAND #() 
NAND_2069_ (
  .A({ S3375 }),
  .B({ S3376 }),
  .Y({ S100 })
);
NAND #() 
NAND_2070_ (
  .A({ datapath_indatatrf_1 }),
  .B({ S3373 }),
  .Y({ S3377 })
);
NAND #() 
NAND_2071_ (
  .A({ datapath_theregisterfile_memtrf_97 }),
  .B({ S3374 }),
  .Y({ S3378 })
);
NAND #() 
NAND_2072_ (
  .A({ S3377 }),
  .B({ S3378 }),
  .Y({ S101 })
);
NAND #() 
NAND_2073_ (
  .A({ datapath_indatatrf_2 }),
  .B({ S3373 }),
  .Y({ S3379 })
);
NAND #() 
NAND_2074_ (
  .A({ datapath_theregisterfile_memtrf_98 }),
  .B({ S3374 }),
  .Y({ S3380 })
);
NAND #() 
NAND_2075_ (
  .A({ S3379 }),
  .B({ S3380 }),
  .Y({ S102 })
);
NAND #() 
NAND_2076_ (
  .A({ datapath_indatatrf_3 }),
  .B({ S3373 }),
  .Y({ S3381 })
);
NAND #() 
NAND_2077_ (
  .A({ datapath_theregisterfile_memtrf_99 }),
  .B({ S3374 }),
  .Y({ S3382 })
);
NAND #() 
NAND_2078_ (
  .A({ S3381 }),
  .B({ S3382 }),
  .Y({ S103 })
);
NAND #() 
NAND_2079_ (
  .A({ datapath_indatatrf_4 }),
  .B({ S3373 }),
  .Y({ S3383 })
);
NAND #() 
NAND_2080_ (
  .A({ datapath_theregisterfile_memtrf_100 }),
  .B({ S3374 }),
  .Y({ S3384 })
);
NAND #() 
NAND_2081_ (
  .A({ S3383 }),
  .B({ S3384 }),
  .Y({ S104 })
);
NAND #() 
NAND_2082_ (
  .A({ datapath_indatatrf_5 }),
  .B({ S3373 }),
  .Y({ S3385 })
);
NAND #() 
NAND_2083_ (
  .A({ datapath_theregisterfile_memtrf_101 }),
  .B({ S3374 }),
  .Y({ S3386 })
);
NAND #() 
NAND_2084_ (
  .A({ S3385 }),
  .B({ S3386 }),
  .Y({ S105 })
);
NAND #() 
NAND_2085_ (
  .A({ datapath_indatatrf_6 }),
  .B({ S3373 }),
  .Y({ S3387 })
);
NAND #() 
NAND_2086_ (
  .A({ datapath_theregisterfile_memtrf_102 }),
  .B({ S3374 }),
  .Y({ S3388 })
);
NAND #() 
NAND_2087_ (
  .A({ S3387 }),
  .B({ S3388 }),
  .Y({ S106 })
);
NAND #() 
NAND_2088_ (
  .A({ datapath_indatatrf_7 }),
  .B({ S3373 }),
  .Y({ S3389 })
);
NAND #() 
NAND_2089_ (
  .A({ datapath_theregisterfile_memtrf_103 }),
  .B({ S3374 }),
  .Y({ S3390 })
);
NAND #() 
NAND_2090_ (
  .A({ S3389 }),
  .B({ S3390 }),
  .Y({ S107 })
);
NAND #() 
NAND_2091_ (
  .A({ datapath_indatatrf_8 }),
  .B({ S3373 }),
  .Y({ S3391 })
);
NAND #() 
NAND_2092_ (
  .A({ datapath_theregisterfile_memtrf_104 }),
  .B({ S3374 }),
  .Y({ S3392 })
);
NAND #() 
NAND_2093_ (
  .A({ S3391 }),
  .B({ S3392 }),
  .Y({ S108 })
);
NAND #() 
NAND_2094_ (
  .A({ datapath_indatatrf_9 }),
  .B({ S3373 }),
  .Y({ S3393 })
);
NAND #() 
NAND_2095_ (
  .A({ datapath_theregisterfile_memtrf_105 }),
  .B({ S3374 }),
  .Y({ S3394 })
);
NAND #() 
NAND_2096_ (
  .A({ S3393 }),
  .B({ S3394 }),
  .Y({ S109 })
);
NAND #() 
NAND_2097_ (
  .A({ datapath_indatatrf_10 }),
  .B({ S3373 }),
  .Y({ S3395 })
);
NAND #() 
NAND_2098_ (
  .A({ datapath_theregisterfile_memtrf_106 }),
  .B({ S3374 }),
  .Y({ S3396 })
);
NAND #() 
NAND_2099_ (
  .A({ S3395 }),
  .B({ S3396 }),
  .Y({ S110 })
);
NAND #() 
NAND_2100_ (
  .A({ datapath_indatatrf_11 }),
  .B({ S3373 }),
  .Y({ S3397 })
);
NAND #() 
NAND_2101_ (
  .A({ datapath_theregisterfile_memtrf_107 }),
  .B({ S3374 }),
  .Y({ S3398 })
);
NAND #() 
NAND_2102_ (
  .A({ S3397 }),
  .B({ S3398 }),
  .Y({ S111 })
);
NAND #() 
NAND_2103_ (
  .A({ datapath_indatatrf_12 }),
  .B({ S3373 }),
  .Y({ S3399 })
);
NAND #() 
NAND_2104_ (
  .A({ datapath_theregisterfile_memtrf_108 }),
  .B({ S3374 }),
  .Y({ S3400 })
);
NAND #() 
NAND_2105_ (
  .A({ S3399 }),
  .B({ S3400 }),
  .Y({ S112 })
);
NAND #() 
NAND_2106_ (
  .A({ datapath_indatatrf_13 }),
  .B({ S3373 }),
  .Y({ S3401 })
);
NAND #() 
NAND_2107_ (
  .A({ datapath_theregisterfile_memtrf_109 }),
  .B({ S3374 }),
  .Y({ S3402 })
);
NAND #() 
NAND_2108_ (
  .A({ S3401 }),
  .B({ S3402 }),
  .Y({ S113 })
);
NAND #() 
NAND_2109_ (
  .A({ datapath_indatatrf_14 }),
  .B({ S3373 }),
  .Y({ S3403 })
);
NAND #() 
NAND_2110_ (
  .A({ datapath_theregisterfile_memtrf_110 }),
  .B({ S3374 }),
  .Y({ S3404 })
);
NAND #() 
NAND_2111_ (
  .A({ S3403 }),
  .B({ S3404 }),
  .Y({ S114 })
);
NAND #() 
NAND_2112_ (
  .A({ datapath_indatatrf_15 }),
  .B({ S3373 }),
  .Y({ S3405 })
);
NAND #() 
NAND_2113_ (
  .A({ datapath_theregisterfile_memtrf_111 }),
  .B({ S3374 }),
  .Y({ S3406 })
);
NAND #() 
NAND_2114_ (
  .A({ S3405 }),
  .B({ S3406 }),
  .Y({ S115 })
);
NOR #() 
NOR_939_ (
  .A({ S1664 }),
  .B({ S3230 }),
  .Y({ S3407 })
);
NAND #() 
NAND_2115_ (
  .A({ S1663 }),
  .B({ S3229 }),
  .Y({ S3408 })
);
NAND #() 
NAND_2116_ (
  .A({ datapath_indatatrf_0 }),
  .B({ S3407 }),
  .Y({ S3409 })
);
NAND #() 
NAND_2117_ (
  .A({ datapath_theregisterfile_memtrf_112 }),
  .B({ S3408 }),
  .Y({ S3410 })
);
NAND #() 
NAND_2118_ (
  .A({ S3409 }),
  .B({ S3410 }),
  .Y({ S116 })
);
NAND #() 
NAND_2119_ (
  .A({ datapath_indatatrf_1 }),
  .B({ S3407 }),
  .Y({ S3411 })
);
NAND #() 
NAND_2120_ (
  .A({ datapath_theregisterfile_memtrf_113 }),
  .B({ S3408 }),
  .Y({ S3412 })
);
NAND #() 
NAND_2121_ (
  .A({ S3411 }),
  .B({ S3412 }),
  .Y({ S117 })
);
NAND #() 
NAND_2122_ (
  .A({ datapath_indatatrf_2 }),
  .B({ S3407 }),
  .Y({ S3413 })
);
NAND #() 
NAND_2123_ (
  .A({ datapath_theregisterfile_memtrf_114 }),
  .B({ S3408 }),
  .Y({ S3414 })
);
NAND #() 
NAND_2124_ (
  .A({ S3413 }),
  .B({ S3414 }),
  .Y({ S118 })
);
NAND #() 
NAND_2125_ (
  .A({ datapath_indatatrf_3 }),
  .B({ S3407 }),
  .Y({ S3415 })
);
NAND #() 
NAND_2126_ (
  .A({ datapath_theregisterfile_memtrf_115 }),
  .B({ S3408 }),
  .Y({ S3416 })
);
NAND #() 
NAND_2127_ (
  .A({ S3415 }),
  .B({ S3416 }),
  .Y({ S119 })
);
NAND #() 
NAND_2128_ (
  .A({ datapath_indatatrf_4 }),
  .B({ S3407 }),
  .Y({ S3417 })
);
NAND #() 
NAND_2129_ (
  .A({ datapath_theregisterfile_memtrf_116 }),
  .B({ S3408 }),
  .Y({ S3418 })
);
NAND #() 
NAND_2130_ (
  .A({ S3417 }),
  .B({ S3418 }),
  .Y({ S120 })
);
NAND #() 
NAND_2131_ (
  .A({ datapath_indatatrf_5 }),
  .B({ S3407 }),
  .Y({ S3419 })
);
NAND #() 
NAND_2132_ (
  .A({ datapath_theregisterfile_memtrf_117 }),
  .B({ S3408 }),
  .Y({ S3420 })
);
NAND #() 
NAND_2133_ (
  .A({ S3419 }),
  .B({ S3420 }),
  .Y({ S121 })
);
NAND #() 
NAND_2134_ (
  .A({ datapath_indatatrf_6 }),
  .B({ S3407 }),
  .Y({ S3421 })
);
NAND #() 
NAND_2135_ (
  .A({ datapath_theregisterfile_memtrf_118 }),
  .B({ S3408 }),
  .Y({ S3422 })
);
NAND #() 
NAND_2136_ (
  .A({ S3421 }),
  .B({ S3422 }),
  .Y({ S122 })
);
NAND #() 
NAND_2137_ (
  .A({ datapath_indatatrf_7 }),
  .B({ S3407 }),
  .Y({ S3423 })
);
NAND #() 
NAND_2138_ (
  .A({ datapath_theregisterfile_memtrf_119 }),
  .B({ S3408 }),
  .Y({ S3424 })
);
NAND #() 
NAND_2139_ (
  .A({ S3423 }),
  .B({ S3424 }),
  .Y({ S123 })
);
NAND #() 
NAND_2140_ (
  .A({ datapath_indatatrf_8 }),
  .B({ S3407 }),
  .Y({ S3425 })
);
NAND #() 
NAND_2141_ (
  .A({ datapath_theregisterfile_memtrf_120 }),
  .B({ S3408 }),
  .Y({ S3426 })
);
NAND #() 
NAND_2142_ (
  .A({ S3425 }),
  .B({ S3426 }),
  .Y({ S124 })
);
NAND #() 
NAND_2143_ (
  .A({ datapath_indatatrf_9 }),
  .B({ S3407 }),
  .Y({ S3427 })
);
NAND #() 
NAND_2144_ (
  .A({ datapath_theregisterfile_memtrf_121 }),
  .B({ S3408 }),
  .Y({ S3428 })
);
NAND #() 
NAND_2145_ (
  .A({ S3427 }),
  .B({ S3428 }),
  .Y({ S125 })
);
NAND #() 
NAND_2146_ (
  .A({ datapath_indatatrf_10 }),
  .B({ S3407 }),
  .Y({ S3429 })
);
NAND #() 
NAND_2147_ (
  .A({ datapath_theregisterfile_memtrf_122 }),
  .B({ S3408 }),
  .Y({ S3430 })
);
NAND #() 
NAND_2148_ (
  .A({ S3429 }),
  .B({ S3430 }),
  .Y({ S126 })
);
NAND #() 
NAND_2149_ (
  .A({ datapath_indatatrf_11 }),
  .B({ S3407 }),
  .Y({ S3431 })
);
NAND #() 
NAND_2150_ (
  .A({ datapath_theregisterfile_memtrf_123 }),
  .B({ S3408 }),
  .Y({ S3432 })
);
NAND #() 
NAND_2151_ (
  .A({ S3431 }),
  .B({ S3432 }),
  .Y({ S127 })
);
NAND #() 
NAND_2152_ (
  .A({ datapath_indatatrf_12 }),
  .B({ S3407 }),
  .Y({ S3433 })
);
NAND #() 
NAND_2153_ (
  .A({ datapath_theregisterfile_memtrf_124 }),
  .B({ S3408 }),
  .Y({ S3434 })
);
NAND #() 
NAND_2154_ (
  .A({ S3433 }),
  .B({ S3434 }),
  .Y({ S128 })
);
NAND #() 
NAND_2155_ (
  .A({ datapath_indatatrf_13 }),
  .B({ S3407 }),
  .Y({ S3435 })
);
NAND #() 
NAND_2156_ (
  .A({ datapath_theregisterfile_memtrf_125 }),
  .B({ S3408 }),
  .Y({ S3436 })
);
NAND #() 
NAND_2157_ (
  .A({ S3435 }),
  .B({ S3436 }),
  .Y({ S129 })
);
NAND #() 
NAND_2158_ (
  .A({ datapath_indatatrf_14 }),
  .B({ S3407 }),
  .Y({ S3437 })
);
NAND #() 
NAND_2159_ (
  .A({ datapath_theregisterfile_memtrf_126 }),
  .B({ S3408 }),
  .Y({ S3438 })
);
NAND #() 
NAND_2160_ (
  .A({ S3437 }),
  .B({ S3438 }),
  .Y({ S130 })
);
NAND #() 
NAND_2161_ (
  .A({ datapath_indatatrf_15 }),
  .B({ S3407 }),
  .Y({ S3439 })
);
NAND #() 
NAND_2162_ (
  .A({ datapath_theregisterfile_memtrf_127 }),
  .B({ S3408 }),
  .Y({ S3440 })
);
NAND #() 
NAND_2163_ (
  .A({ S3439 }),
  .B({ S3440 }),
  .Y({ S131 })
);
NOR #() 
NOR_940_ (
  .A({ S1687 }),
  .B({ S3304 }),
  .Y({ S3441 })
);
NAND #() 
NAND_2164_ (
  .A({ S1686 }),
  .B({ S3303 }),
  .Y({ S3442 })
);
NAND #() 
NAND_2165_ (
  .A({ datapath_indatatrf_0 }),
  .B({ S3441 }),
  .Y({ S3443 })
);
NAND #() 
NAND_2166_ (
  .A({ datapath_theregisterfile_memtrf_0 }),
  .B({ S3442 }),
  .Y({ S3444 })
);
NAND #() 
NAND_2167_ (
  .A({ S3443 }),
  .B({ S3444 }),
  .Y({ S132 })
);
NAND #() 
NAND_2168_ (
  .A({ datapath_indatatrf_1 }),
  .B({ S3441 }),
  .Y({ S3445 })
);
NAND #() 
NAND_2169_ (
  .A({ datapath_theregisterfile_memtrf_1 }),
  .B({ S3442 }),
  .Y({ S3446 })
);
NAND #() 
NAND_2170_ (
  .A({ S3445 }),
  .B({ S3446 }),
  .Y({ S133 })
);
NAND #() 
NAND_2171_ (
  .A({ datapath_indatatrf_2 }),
  .B({ S3441 }),
  .Y({ S3447 })
);
NAND #() 
NAND_2172_ (
  .A({ datapath_theregisterfile_memtrf_2 }),
  .B({ S3442 }),
  .Y({ S3448 })
);
NAND #() 
NAND_2173_ (
  .A({ S3447 }),
  .B({ S3448 }),
  .Y({ S134 })
);
NAND #() 
NAND_2174_ (
  .A({ datapath_indatatrf_3 }),
  .B({ S3441 }),
  .Y({ S3449 })
);
NAND #() 
NAND_2175_ (
  .A({ datapath_theregisterfile_memtrf_3 }),
  .B({ S3442 }),
  .Y({ S3450 })
);
NAND #() 
NAND_2176_ (
  .A({ S3449 }),
  .B({ S3450 }),
  .Y({ S135 })
);
NAND #() 
NAND_2177_ (
  .A({ datapath_indatatrf_4 }),
  .B({ S3441 }),
  .Y({ S3451 })
);
NAND #() 
NAND_2178_ (
  .A({ datapath_theregisterfile_memtrf_4 }),
  .B({ S3442 }),
  .Y({ S3452 })
);
NAND #() 
NAND_2179_ (
  .A({ S3451 }),
  .B({ S3452 }),
  .Y({ S136 })
);
NAND #() 
NAND_2180_ (
  .A({ datapath_indatatrf_5 }),
  .B({ S3441 }),
  .Y({ S3453 })
);
NAND #() 
NAND_2181_ (
  .A({ datapath_theregisterfile_memtrf_5 }),
  .B({ S3442 }),
  .Y({ S3454 })
);
NAND #() 
NAND_2182_ (
  .A({ S3453 }),
  .B({ S3454 }),
  .Y({ S137 })
);
NAND #() 
NAND_2183_ (
  .A({ datapath_indatatrf_6 }),
  .B({ S3441 }),
  .Y({ S3455 })
);
NAND #() 
NAND_2184_ (
  .A({ datapath_theregisterfile_memtrf_6 }),
  .B({ S3442 }),
  .Y({ S3456 })
);
NAND #() 
NAND_2185_ (
  .A({ S3455 }),
  .B({ S3456 }),
  .Y({ S138 })
);
NAND #() 
NAND_2186_ (
  .A({ datapath_indatatrf_7 }),
  .B({ S3441 }),
  .Y({ S3457 })
);
NAND #() 
NAND_2187_ (
  .A({ datapath_theregisterfile_memtrf_7 }),
  .B({ S3442 }),
  .Y({ S3458 })
);
NAND #() 
NAND_2188_ (
  .A({ S3457 }),
  .B({ S3458 }),
  .Y({ S139 })
);
NAND #() 
NAND_2189_ (
  .A({ datapath_indatatrf_8 }),
  .B({ S3441 }),
  .Y({ S3459 })
);
NAND #() 
NAND_2190_ (
  .A({ datapath_theregisterfile_memtrf_8 }),
  .B({ S3442 }),
  .Y({ S3460 })
);
NAND #() 
NAND_2191_ (
  .A({ S3459 }),
  .B({ S3460 }),
  .Y({ S140 })
);
NAND #() 
NAND_2192_ (
  .A({ datapath_indatatrf_9 }),
  .B({ S3441 }),
  .Y({ S3461 })
);
NAND #() 
NAND_2193_ (
  .A({ datapath_theregisterfile_memtrf_9 }),
  .B({ S3442 }),
  .Y({ S3462 })
);
NAND #() 
NAND_2194_ (
  .A({ S3461 }),
  .B({ S3462 }),
  .Y({ S141 })
);
NAND #() 
NAND_2195_ (
  .A({ datapath_indatatrf_10 }),
  .B({ S3441 }),
  .Y({ S3463 })
);
NAND #() 
NAND_2196_ (
  .A({ datapath_theregisterfile_memtrf_10 }),
  .B({ S3442 }),
  .Y({ S3464 })
);
NAND #() 
NAND_2197_ (
  .A({ S3463 }),
  .B({ S3464 }),
  .Y({ S142 })
);
NAND #() 
NAND_2198_ (
  .A({ datapath_indatatrf_11 }),
  .B({ S3441 }),
  .Y({ S3465 })
);
NAND #() 
NAND_2199_ (
  .A({ datapath_theregisterfile_memtrf_11 }),
  .B({ S3442 }),
  .Y({ S3466 })
);
NAND #() 
NAND_2200_ (
  .A({ S3465 }),
  .B({ S3466 }),
  .Y({ S143 })
);
NAND #() 
NAND_2201_ (
  .A({ datapath_indatatrf_12 }),
  .B({ S3441 }),
  .Y({ S3467 })
);
NAND #() 
NAND_2202_ (
  .A({ datapath_theregisterfile_memtrf_12 }),
  .B({ S3442 }),
  .Y({ S3468 })
);
NAND #() 
NAND_2203_ (
  .A({ S3467 }),
  .B({ S3468 }),
  .Y({ S144 })
);
NAND #() 
NAND_2204_ (
  .A({ datapath_indatatrf_13 }),
  .B({ S3441 }),
  .Y({ S3469 })
);
NAND #() 
NAND_2205_ (
  .A({ datapath_theregisterfile_memtrf_13 }),
  .B({ S3442 }),
  .Y({ S3470 })
);
NAND #() 
NAND_2206_ (
  .A({ S3469 }),
  .B({ S3470 }),
  .Y({ S145 })
);
NAND #() 
NAND_2207_ (
  .A({ datapath_indatatrf_14 }),
  .B({ S3441 }),
  .Y({ S3471 })
);
NAND #() 
NAND_2208_ (
  .A({ datapath_theregisterfile_memtrf_14 }),
  .B({ S3442 }),
  .Y({ S3472 })
);
NAND #() 
NAND_2209_ (
  .A({ S3471 }),
  .B({ S3472 }),
  .Y({ S146 })
);
NAND #() 
NAND_2210_ (
  .A({ datapath_indatatrf_15 }),
  .B({ S3441 }),
  .Y({ S3473 })
);
NAND #() 
NAND_2211_ (
  .A({ datapath_theregisterfile_memtrf_15 }),
  .B({ S3442 }),
  .Y({ S3474 })
);
NAND #() 
NAND_2212_ (
  .A({ S3473 }),
  .B({ S3474 }),
  .Y({ S147 })
);
NOR #() 
NOR_941_ (
  .A({ S3228 }),
  .B({ S3268 }),
  .Y({ S3475 })
);
NAND #() 
NAND_2213_ (
  .A({ S3227 }),
  .B({ S3267 }),
  .Y({ S3476 })
);
NAND #() 
NAND_2214_ (
  .A({ datapath_indatatrf_0 }),
  .B({ S3475 }),
  .Y({ S3477 })
);
NAND #() 
NAND_2215_ (
  .A({ datapath_theregisterfile_memtrf_144 }),
  .B({ S3476 }),
  .Y({ S3478 })
);
NAND #() 
NAND_2216_ (
  .A({ S3477 }),
  .B({ S3478 }),
  .Y({ S148 })
);
NAND #() 
NAND_2217_ (
  .A({ datapath_indatatrf_1 }),
  .B({ S3475 }),
  .Y({ S3479 })
);
NAND #() 
NAND_2218_ (
  .A({ datapath_theregisterfile_memtrf_145 }),
  .B({ S3476 }),
  .Y({ S3480 })
);
NAND #() 
NAND_2219_ (
  .A({ S3479 }),
  .B({ S3480 }),
  .Y({ S149 })
);
NAND #() 
NAND_2220_ (
  .A({ datapath_indatatrf_2 }),
  .B({ S3475 }),
  .Y({ S3481 })
);
NAND #() 
NAND_2221_ (
  .A({ datapath_theregisterfile_memtrf_146 }),
  .B({ S3476 }),
  .Y({ S3482 })
);
NAND #() 
NAND_2222_ (
  .A({ S3481 }),
  .B({ S3482 }),
  .Y({ S150 })
);
NAND #() 
NAND_2223_ (
  .A({ datapath_indatatrf_3 }),
  .B({ S3475 }),
  .Y({ S3483 })
);
NAND #() 
NAND_2224_ (
  .A({ datapath_theregisterfile_memtrf_147 }),
  .B({ S3476 }),
  .Y({ S3484 })
);
NAND #() 
NAND_2225_ (
  .A({ S3483 }),
  .B({ S3484 }),
  .Y({ S151 })
);
NAND #() 
NAND_2226_ (
  .A({ datapath_indatatrf_4 }),
  .B({ S3475 }),
  .Y({ S3485 })
);
NAND #() 
NAND_2227_ (
  .A({ datapath_theregisterfile_memtrf_148 }),
  .B({ S3476 }),
  .Y({ S3486 })
);
NAND #() 
NAND_2228_ (
  .A({ S3485 }),
  .B({ S3486 }),
  .Y({ S152 })
);
NAND #() 
NAND_2229_ (
  .A({ datapath_indatatrf_5 }),
  .B({ S3475 }),
  .Y({ S3487 })
);
NAND #() 
NAND_2230_ (
  .A({ datapath_theregisterfile_memtrf_149 }),
  .B({ S3476 }),
  .Y({ S3488 })
);
NAND #() 
NAND_2231_ (
  .A({ S3487 }),
  .B({ S3488 }),
  .Y({ S153 })
);
NAND #() 
NAND_2232_ (
  .A({ datapath_indatatrf_6 }),
  .B({ S3475 }),
  .Y({ S3489 })
);
NAND #() 
NAND_2233_ (
  .A({ datapath_theregisterfile_memtrf_150 }),
  .B({ S3476 }),
  .Y({ S3490 })
);
NAND #() 
NAND_2234_ (
  .A({ S3489 }),
  .B({ S3490 }),
  .Y({ S154 })
);
NAND #() 
NAND_2235_ (
  .A({ datapath_indatatrf_7 }),
  .B({ S3475 }),
  .Y({ S3491 })
);
NAND #() 
NAND_2236_ (
  .A({ datapath_theregisterfile_memtrf_151 }),
  .B({ S3476 }),
  .Y({ S3492 })
);
NAND #() 
NAND_2237_ (
  .A({ S3491 }),
  .B({ S3492 }),
  .Y({ S155 })
);
NAND #() 
NAND_2238_ (
  .A({ datapath_indatatrf_8 }),
  .B({ S3475 }),
  .Y({ S3493 })
);
NAND #() 
NAND_2239_ (
  .A({ datapath_theregisterfile_memtrf_152 }),
  .B({ S3476 }),
  .Y({ S3494 })
);
NAND #() 
NAND_2240_ (
  .A({ S3493 }),
  .B({ S3494 }),
  .Y({ S156 })
);
NAND #() 
NAND_2241_ (
  .A({ datapath_indatatrf_9 }),
  .B({ S3475 }),
  .Y({ S3495 })
);
NAND #() 
NAND_2242_ (
  .A({ datapath_theregisterfile_memtrf_153 }),
  .B({ S3476 }),
  .Y({ S3496 })
);
NAND #() 
NAND_2243_ (
  .A({ S3495 }),
  .B({ S3496 }),
  .Y({ S157 })
);
NAND #() 
NAND_2244_ (
  .A({ datapath_indatatrf_10 }),
  .B({ S3475 }),
  .Y({ S3497 })
);
NAND #() 
NAND_2245_ (
  .A({ datapath_theregisterfile_memtrf_154 }),
  .B({ S3476 }),
  .Y({ S3498 })
);
NAND #() 
NAND_2246_ (
  .A({ S3497 }),
  .B({ S3498 }),
  .Y({ S158 })
);
NAND #() 
NAND_2247_ (
  .A({ datapath_indatatrf_11 }),
  .B({ S3475 }),
  .Y({ S3499 })
);
NAND #() 
NAND_2248_ (
  .A({ datapath_theregisterfile_memtrf_155 }),
  .B({ S3476 }),
  .Y({ S3500 })
);
NAND #() 
NAND_2249_ (
  .A({ S3499 }),
  .B({ S3500 }),
  .Y({ S159 })
);
NAND #() 
NAND_2250_ (
  .A({ datapath_indatatrf_12 }),
  .B({ S3475 }),
  .Y({ S3501 })
);
NAND #() 
NAND_2251_ (
  .A({ datapath_theregisterfile_memtrf_156 }),
  .B({ S3476 }),
  .Y({ S3502 })
);
NAND #() 
NAND_2252_ (
  .A({ S3501 }),
  .B({ S3502 }),
  .Y({ S160 })
);
NAND #() 
NAND_2253_ (
  .A({ datapath_indatatrf_13 }),
  .B({ S3475 }),
  .Y({ S3503 })
);
NAND #() 
NAND_2254_ (
  .A({ datapath_theregisterfile_memtrf_157 }),
  .B({ S3476 }),
  .Y({ S3504 })
);
NAND #() 
NAND_2255_ (
  .A({ S3503 }),
  .B({ S3504 }),
  .Y({ S161 })
);
NAND #() 
NAND_2256_ (
  .A({ datapath_indatatrf_14 }),
  .B({ S3475 }),
  .Y({ S3505 })
);
NAND #() 
NAND_2257_ (
  .A({ datapath_theregisterfile_memtrf_158 }),
  .B({ S3476 }),
  .Y({ S3506 })
);
NAND #() 
NAND_2258_ (
  .A({ S3505 }),
  .B({ S3506 }),
  .Y({ S162 })
);
NAND #() 
NAND_2259_ (
  .A({ datapath_indatatrf_15 }),
  .B({ S3475 }),
  .Y({ S3507 })
);
NAND #() 
NAND_2260_ (
  .A({ datapath_theregisterfile_memtrf_159 }),
  .B({ S3476 }),
  .Y({ S3508 })
);
NAND #() 
NAND_2261_ (
  .A({ S3507 }),
  .B({ S3508 }),
  .Y({ S163 })
);
NOR #() 
NOR_942_ (
  .A({ S3192 }),
  .B({ S3266 }),
  .Y({ S3509 })
);
NAND #() 
NAND_2262_ (
  .A({ S3191 }),
  .B({ S3265 }),
  .Y({ S3510 })
);
NAND #() 
NAND_2263_ (
  .A({ datapath_indatatrf_0 }),
  .B({ S3509 }),
  .Y({ S3511 })
);
NAND #() 
NAND_2264_ (
  .A({ datapath_theregisterfile_memtrf_160 }),
  .B({ S3510 }),
  .Y({ S3512 })
);
NAND #() 
NAND_2265_ (
  .A({ S3511 }),
  .B({ S3512 }),
  .Y({ S164 })
);
NAND #() 
NAND_2266_ (
  .A({ datapath_indatatrf_1 }),
  .B({ S3509 }),
  .Y({ S3513 })
);
NAND #() 
NAND_2267_ (
  .A({ datapath_theregisterfile_memtrf_161 }),
  .B({ S3510 }),
  .Y({ S3514 })
);
NAND #() 
NAND_2268_ (
  .A({ S3513 }),
  .B({ S3514 }),
  .Y({ S165 })
);
NAND #() 
NAND_2269_ (
  .A({ datapath_indatatrf_2 }),
  .B({ S3509 }),
  .Y({ S3515 })
);
NAND #() 
NAND_2270_ (
  .A({ datapath_theregisterfile_memtrf_162 }),
  .B({ S3510 }),
  .Y({ S3516 })
);
NAND #() 
NAND_2271_ (
  .A({ S3515 }),
  .B({ S3516 }),
  .Y({ S166 })
);
NAND #() 
NAND_2272_ (
  .A({ datapath_indatatrf_3 }),
  .B({ S3509 }),
  .Y({ S3517 })
);
NAND #() 
NAND_2273_ (
  .A({ datapath_theregisterfile_memtrf_163 }),
  .B({ S3510 }),
  .Y({ S3518 })
);
NAND #() 
NAND_2274_ (
  .A({ S3517 }),
  .B({ S3518 }),
  .Y({ S167 })
);
NAND #() 
NAND_2275_ (
  .A({ datapath_indatatrf_4 }),
  .B({ S3509 }),
  .Y({ S3519 })
);
NAND #() 
NAND_2276_ (
  .A({ datapath_theregisterfile_memtrf_164 }),
  .B({ S3510 }),
  .Y({ S3520 })
);
NAND #() 
NAND_2277_ (
  .A({ S3519 }),
  .B({ S3520 }),
  .Y({ S168 })
);
NAND #() 
NAND_2278_ (
  .A({ datapath_indatatrf_5 }),
  .B({ S3509 }),
  .Y({ S3521 })
);
NAND #() 
NAND_2279_ (
  .A({ datapath_theregisterfile_memtrf_165 }),
  .B({ S3510 }),
  .Y({ S3522 })
);
NAND #() 
NAND_2280_ (
  .A({ S3521 }),
  .B({ S3522 }),
  .Y({ S169 })
);
NAND #() 
NAND_2281_ (
  .A({ datapath_indatatrf_6 }),
  .B({ S3509 }),
  .Y({ S3523 })
);
NAND #() 
NAND_2282_ (
  .A({ datapath_theregisterfile_memtrf_166 }),
  .B({ S3510 }),
  .Y({ S3524 })
);
NAND #() 
NAND_2283_ (
  .A({ S3523 }),
  .B({ S3524 }),
  .Y({ S170 })
);
NAND #() 
NAND_2284_ (
  .A({ datapath_indatatrf_7 }),
  .B({ S3509 }),
  .Y({ S3525 })
);
NAND #() 
NAND_2285_ (
  .A({ datapath_theregisterfile_memtrf_167 }),
  .B({ S3510 }),
  .Y({ S3526 })
);
NAND #() 
NAND_2286_ (
  .A({ S3525 }),
  .B({ S3526 }),
  .Y({ S171 })
);
NAND #() 
NAND_2287_ (
  .A({ datapath_indatatrf_8 }),
  .B({ S3509 }),
  .Y({ S3527 })
);
NAND #() 
NAND_2288_ (
  .A({ datapath_theregisterfile_memtrf_168 }),
  .B({ S3510 }),
  .Y({ S3528 })
);
NAND #() 
NAND_2289_ (
  .A({ S3527 }),
  .B({ S3528 }),
  .Y({ S172 })
);
NAND #() 
NAND_2290_ (
  .A({ datapath_indatatrf_9 }),
  .B({ S3509 }),
  .Y({ S3529 })
);
NAND #() 
NAND_2291_ (
  .A({ datapath_theregisterfile_memtrf_169 }),
  .B({ S3510 }),
  .Y({ S3530 })
);
NAND #() 
NAND_2292_ (
  .A({ S3529 }),
  .B({ S3530 }),
  .Y({ S173 })
);
NAND #() 
NAND_2293_ (
  .A({ datapath_indatatrf_10 }),
  .B({ S3509 }),
  .Y({ S3531 })
);
NAND #() 
NAND_2294_ (
  .A({ datapath_theregisterfile_memtrf_170 }),
  .B({ S3510 }),
  .Y({ S3532 })
);
NAND #() 
NAND_2295_ (
  .A({ S3531 }),
  .B({ S3532 }),
  .Y({ S174 })
);
NAND #() 
NAND_2296_ (
  .A({ datapath_indatatrf_11 }),
  .B({ S3509 }),
  .Y({ S3533 })
);
NAND #() 
NAND_2297_ (
  .A({ datapath_theregisterfile_memtrf_171 }),
  .B({ S3510 }),
  .Y({ S3534 })
);
NAND #() 
NAND_2298_ (
  .A({ S3533 }),
  .B({ S3534 }),
  .Y({ S175 })
);
NAND #() 
NAND_2299_ (
  .A({ datapath_indatatrf_12 }),
  .B({ S3509 }),
  .Y({ S3535 })
);
NAND #() 
NAND_2300_ (
  .A({ datapath_theregisterfile_memtrf_172 }),
  .B({ S3510 }),
  .Y({ S3536 })
);
NAND #() 
NAND_2301_ (
  .A({ S3535 }),
  .B({ S3536 }),
  .Y({ S176 })
);
NAND #() 
NAND_2302_ (
  .A({ datapath_indatatrf_13 }),
  .B({ S3509 }),
  .Y({ S3537 })
);
NAND #() 
NAND_2303_ (
  .A({ datapath_theregisterfile_memtrf_173 }),
  .B({ S3510 }),
  .Y({ S3538 })
);
NAND #() 
NAND_2304_ (
  .A({ S3537 }),
  .B({ S3538 }),
  .Y({ S177 })
);
NAND #() 
NAND_2305_ (
  .A({ datapath_indatatrf_14 }),
  .B({ S3509 }),
  .Y({ S3539 })
);
NAND #() 
NAND_2306_ (
  .A({ datapath_theregisterfile_memtrf_174 }),
  .B({ S3510 }),
  .Y({ S3540 })
);
NAND #() 
NAND_2307_ (
  .A({ S3539 }),
  .B({ S3540 }),
  .Y({ S178 })
);
NAND #() 
NAND_2308_ (
  .A({ datapath_indatatrf_15 }),
  .B({ S3509 }),
  .Y({ S3541 })
);
NAND #() 
NAND_2309_ (
  .A({ datapath_theregisterfile_memtrf_175 }),
  .B({ S3510 }),
  .Y({ S3542 })
);
NAND #() 
NAND_2310_ (
  .A({ S3541 }),
  .B({ S3542 }),
  .Y({ S179 })
);
NOR #() 
NOR_943_ (
  .A({ S3230 }),
  .B({ S3266 }),
  .Y({ S3543 })
);
NAND #() 
NAND_2311_ (
  .A({ S3229 }),
  .B({ S3265 }),
  .Y({ S3544 })
);
NAND #() 
NAND_2312_ (
  .A({ datapath_indatatrf_0 }),
  .B({ S3543 }),
  .Y({ S3545 })
);
NAND #() 
NAND_2313_ (
  .A({ datapath_theregisterfile_memtrf_176 }),
  .B({ S3544 }),
  .Y({ S3546 })
);
NAND #() 
NAND_2314_ (
  .A({ S3545 }),
  .B({ S3546 }),
  .Y({ S180 })
);
NAND #() 
NAND_2315_ (
  .A({ datapath_indatatrf_1 }),
  .B({ S3543 }),
  .Y({ S3547 })
);
NAND #() 
NAND_2316_ (
  .A({ datapath_theregisterfile_memtrf_177 }),
  .B({ S3544 }),
  .Y({ S3548 })
);
NAND #() 
NAND_2317_ (
  .A({ S3547 }),
  .B({ S3548 }),
  .Y({ S181 })
);
NAND #() 
NAND_2318_ (
  .A({ datapath_indatatrf_2 }),
  .B({ S3543 }),
  .Y({ S3549 })
);
NAND #() 
NAND_2319_ (
  .A({ datapath_theregisterfile_memtrf_178 }),
  .B({ S3544 }),
  .Y({ S3550 })
);
NAND #() 
NAND_2320_ (
  .A({ S3549 }),
  .B({ S3550 }),
  .Y({ S182 })
);
NAND #() 
NAND_2321_ (
  .A({ datapath_indatatrf_3 }),
  .B({ S3543 }),
  .Y({ S3551 })
);
NAND #() 
NAND_2322_ (
  .A({ datapath_theregisterfile_memtrf_179 }),
  .B({ S3544 }),
  .Y({ S3552 })
);
NAND #() 
NAND_2323_ (
  .A({ S3551 }),
  .B({ S3552 }),
  .Y({ S183 })
);
NAND #() 
NAND_2324_ (
  .A({ datapath_indatatrf_4 }),
  .B({ S3543 }),
  .Y({ S3553 })
);
NAND #() 
NAND_2325_ (
  .A({ datapath_theregisterfile_memtrf_180 }),
  .B({ S3544 }),
  .Y({ S3554 })
);
NAND #() 
NAND_2326_ (
  .A({ S3553 }),
  .B({ S3554 }),
  .Y({ S184 })
);
NAND #() 
NAND_2327_ (
  .A({ datapath_indatatrf_5 }),
  .B({ S3543 }),
  .Y({ S3555 })
);
NAND #() 
NAND_2328_ (
  .A({ datapath_theregisterfile_memtrf_181 }),
  .B({ S3544 }),
  .Y({ S3556 })
);
NAND #() 
NAND_2329_ (
  .A({ S3555 }),
  .B({ S3556 }),
  .Y({ S185 })
);
NAND #() 
NAND_2330_ (
  .A({ datapath_indatatrf_6 }),
  .B({ S3543 }),
  .Y({ S3557 })
);
NAND #() 
NAND_2331_ (
  .A({ datapath_theregisterfile_memtrf_182 }),
  .B({ S3544 }),
  .Y({ S3558 })
);
NAND #() 
NAND_2332_ (
  .A({ S3557 }),
  .B({ S3558 }),
  .Y({ S186 })
);
NAND #() 
NAND_2333_ (
  .A({ datapath_indatatrf_7 }),
  .B({ S3543 }),
  .Y({ S3559 })
);
NAND #() 
NAND_2334_ (
  .A({ datapath_theregisterfile_memtrf_183 }),
  .B({ S3544 }),
  .Y({ S3560 })
);
NAND #() 
NAND_2335_ (
  .A({ S3559 }),
  .B({ S3560 }),
  .Y({ S187 })
);
NAND #() 
NAND_2336_ (
  .A({ datapath_indatatrf_8 }),
  .B({ S3543 }),
  .Y({ S3561 })
);
NAND #() 
NAND_2337_ (
  .A({ datapath_theregisterfile_memtrf_184 }),
  .B({ S3544 }),
  .Y({ S3562 })
);
NAND #() 
NAND_2338_ (
  .A({ S3561 }),
  .B({ S3562 }),
  .Y({ S188 })
);
NAND #() 
NAND_2339_ (
  .A({ datapath_indatatrf_9 }),
  .B({ S3543 }),
  .Y({ S3563 })
);
NAND #() 
NAND_2340_ (
  .A({ datapath_theregisterfile_memtrf_185 }),
  .B({ S3544 }),
  .Y({ S3564 })
);
NAND #() 
NAND_2341_ (
  .A({ S3563 }),
  .B({ S3564 }),
  .Y({ S189 })
);
NAND #() 
NAND_2342_ (
  .A({ datapath_indatatrf_10 }),
  .B({ S3543 }),
  .Y({ S3565 })
);
NAND #() 
NAND_2343_ (
  .A({ datapath_theregisterfile_memtrf_186 }),
  .B({ S3544 }),
  .Y({ S3566 })
);
NAND #() 
NAND_2344_ (
  .A({ S3565 }),
  .B({ S3566 }),
  .Y({ S190 })
);
NAND #() 
NAND_2345_ (
  .A({ datapath_indatatrf_11 }),
  .B({ S3543 }),
  .Y({ S3567 })
);
NAND #() 
NAND_2346_ (
  .A({ datapath_theregisterfile_memtrf_187 }),
  .B({ S3544 }),
  .Y({ S3568 })
);
NAND #() 
NAND_2347_ (
  .A({ S3567 }),
  .B({ S3568 }),
  .Y({ S191 })
);
NAND #() 
NAND_2348_ (
  .A({ datapath_indatatrf_12 }),
  .B({ S3543 }),
  .Y({ S3569 })
);
NAND #() 
NAND_2349_ (
  .A({ datapath_theregisterfile_memtrf_188 }),
  .B({ S3544 }),
  .Y({ S3570 })
);
NAND #() 
NAND_2350_ (
  .A({ S3569 }),
  .B({ S3570 }),
  .Y({ S192 })
);
NAND #() 
NAND_2351_ (
  .A({ datapath_indatatrf_13 }),
  .B({ S3543 }),
  .Y({ S3571 })
);
NAND #() 
NAND_2352_ (
  .A({ datapath_theregisterfile_memtrf_189 }),
  .B({ S3544 }),
  .Y({ S3572 })
);
NAND #() 
NAND_2353_ (
  .A({ S3571 }),
  .B({ S3572 }),
  .Y({ S193 })
);
NAND #() 
NAND_2354_ (
  .A({ datapath_indatatrf_14 }),
  .B({ S3543 }),
  .Y({ S3573 })
);
NAND #() 
NAND_2355_ (
  .A({ datapath_theregisterfile_memtrf_190 }),
  .B({ S3544 }),
  .Y({ S3574 })
);
NAND #() 
NAND_2356_ (
  .A({ S3573 }),
  .B({ S3574 }),
  .Y({ S194 })
);
NAND #() 
NAND_2357_ (
  .A({ datapath_indatatrf_15 }),
  .B({ S3543 }),
  .Y({ S3575 })
);
NAND #() 
NAND_2358_ (
  .A({ datapath_theregisterfile_memtrf_191 }),
  .B({ S3544 }),
  .Y({ S3576 })
);
NAND #() 
NAND_2359_ (
  .A({ S3575 }),
  .B({ S3576 }),
  .Y({ S195 })
);
NOR #() 
NOR_944_ (
  .A({ S1654 }),
  .B({ S1661 }),
  .Y({ S3577 })
);
NAND #() 
NAND_2360_ (
  .A({ S1655 }),
  .B({ S1662 }),
  .Y({ S3578 })
);
NOR #() 
NOR_945_ (
  .A({ S1672 }),
  .B({ S3578 }),
  .Y({ S3579 })
);
NAND #() 
NAND_2361_ (
  .A({ S1671 }),
  .B({ S3577 }),
  .Y({ S3580 })
);
NOR #() 
NOR_946_ (
  .A({ S1687 }),
  .B({ S3580 }),
  .Y({ S3581 })
);
NAND #() 
NAND_2362_ (
  .A({ S1686 }),
  .B({ S3579 }),
  .Y({ S3582 })
);
NAND #() 
NAND_2363_ (
  .A({ datapath_indatatrf_0 }),
  .B({ S3581 }),
  .Y({ S3583 })
);
NAND #() 
NAND_2364_ (
  .A({ datapath_theregisterfile_memtrf_192 }),
  .B({ S3582 }),
  .Y({ S3584 })
);
NAND #() 
NAND_2365_ (
  .A({ S3583 }),
  .B({ S3584 }),
  .Y({ S196 })
);
NAND #() 
NAND_2366_ (
  .A({ datapath_indatatrf_1 }),
  .B({ S3581 }),
  .Y({ S3585 })
);
NAND #() 
NAND_2367_ (
  .A({ datapath_theregisterfile_memtrf_193 }),
  .B({ S3582 }),
  .Y({ S3586 })
);
NAND #() 
NAND_2368_ (
  .A({ S3585 }),
  .B({ S3586 }),
  .Y({ S197 })
);
NAND #() 
NAND_2369_ (
  .A({ datapath_indatatrf_2 }),
  .B({ S3581 }),
  .Y({ S3587 })
);
NAND #() 
NAND_2370_ (
  .A({ datapath_theregisterfile_memtrf_194 }),
  .B({ S3582 }),
  .Y({ S3588 })
);
NAND #() 
NAND_2371_ (
  .A({ S3587 }),
  .B({ S3588 }),
  .Y({ S198 })
);
NAND #() 
NAND_2372_ (
  .A({ datapath_indatatrf_3 }),
  .B({ S3581 }),
  .Y({ S3589 })
);
NAND #() 
NAND_2373_ (
  .A({ datapath_theregisterfile_memtrf_195 }),
  .B({ S3582 }),
  .Y({ S3590 })
);
NAND #() 
NAND_2374_ (
  .A({ S3589 }),
  .B({ S3590 }),
  .Y({ S199 })
);
NAND #() 
NAND_2375_ (
  .A({ datapath_indatatrf_4 }),
  .B({ S3581 }),
  .Y({ S3591 })
);
NAND #() 
NAND_2376_ (
  .A({ datapath_theregisterfile_memtrf_196 }),
  .B({ S3582 }),
  .Y({ S3592 })
);
NAND #() 
NAND_2377_ (
  .A({ S3591 }),
  .B({ S3592 }),
  .Y({ S200 })
);
NAND #() 
NAND_2378_ (
  .A({ datapath_indatatrf_5 }),
  .B({ S3581 }),
  .Y({ S3593 })
);
NAND #() 
NAND_2379_ (
  .A({ datapath_theregisterfile_memtrf_197 }),
  .B({ S3582 }),
  .Y({ S3594 })
);
NAND #() 
NAND_2380_ (
  .A({ S3593 }),
  .B({ S3594 }),
  .Y({ S201 })
);
NAND #() 
NAND_2381_ (
  .A({ datapath_indatatrf_6 }),
  .B({ S3581 }),
  .Y({ S3595 })
);
NAND #() 
NAND_2382_ (
  .A({ datapath_theregisterfile_memtrf_198 }),
  .B({ S3582 }),
  .Y({ S3596 })
);
NAND #() 
NAND_2383_ (
  .A({ S3595 }),
  .B({ S3596 }),
  .Y({ S202 })
);
NAND #() 
NAND_2384_ (
  .A({ datapath_indatatrf_7 }),
  .B({ S3581 }),
  .Y({ S3597 })
);
NAND #() 
NAND_2385_ (
  .A({ datapath_theregisterfile_memtrf_199 }),
  .B({ S3582 }),
  .Y({ S3598 })
);
NAND #() 
NAND_2386_ (
  .A({ S3597 }),
  .B({ S3598 }),
  .Y({ S203 })
);
NAND #() 
NAND_2387_ (
  .A({ datapath_indatatrf_8 }),
  .B({ S3581 }),
  .Y({ S3599 })
);
NAND #() 
NAND_2388_ (
  .A({ datapath_theregisterfile_memtrf_200 }),
  .B({ S3582 }),
  .Y({ S3600 })
);
NAND #() 
NAND_2389_ (
  .A({ S3599 }),
  .B({ S3600 }),
  .Y({ S204 })
);
NAND #() 
NAND_2390_ (
  .A({ datapath_indatatrf_9 }),
  .B({ S3581 }),
  .Y({ S3601 })
);
NAND #() 
NAND_2391_ (
  .A({ datapath_theregisterfile_memtrf_201 }),
  .B({ S3582 }),
  .Y({ S3602 })
);
NAND #() 
NAND_2392_ (
  .A({ S3601 }),
  .B({ S3602 }),
  .Y({ S205 })
);
NAND #() 
NAND_2393_ (
  .A({ datapath_indatatrf_10 }),
  .B({ S3581 }),
  .Y({ S3603 })
);
NAND #() 
NAND_2394_ (
  .A({ datapath_theregisterfile_memtrf_202 }),
  .B({ S3582 }),
  .Y({ S3604 })
);
NAND #() 
NAND_2395_ (
  .A({ S3603 }),
  .B({ S3604 }),
  .Y({ S206 })
);
NAND #() 
NAND_2396_ (
  .A({ datapath_indatatrf_11 }),
  .B({ S3581 }),
  .Y({ S3605 })
);
NAND #() 
NAND_2397_ (
  .A({ datapath_theregisterfile_memtrf_203 }),
  .B({ S3582 }),
  .Y({ S3606 })
);
NAND #() 
NAND_2398_ (
  .A({ S3605 }),
  .B({ S3606 }),
  .Y({ S207 })
);
NAND #() 
NAND_2399_ (
  .A({ datapath_indatatrf_12 }),
  .B({ S3581 }),
  .Y({ S3607 })
);
NAND #() 
NAND_2400_ (
  .A({ datapath_theregisterfile_memtrf_204 }),
  .B({ S3582 }),
  .Y({ S3608 })
);
NAND #() 
NAND_2401_ (
  .A({ S3607 }),
  .B({ S3608 }),
  .Y({ S208 })
);
NAND #() 
NAND_2402_ (
  .A({ datapath_indatatrf_13 }),
  .B({ S3581 }),
  .Y({ S3609 })
);
NAND #() 
NAND_2403_ (
  .A({ datapath_theregisterfile_memtrf_205 }),
  .B({ S3582 }),
  .Y({ S3610 })
);
NAND #() 
NAND_2404_ (
  .A({ S3609 }),
  .B({ S3610 }),
  .Y({ S209 })
);
NAND #() 
NAND_2405_ (
  .A({ datapath_indatatrf_14 }),
  .B({ S3581 }),
  .Y({ S3611 })
);
NAND #() 
NAND_2406_ (
  .A({ datapath_theregisterfile_memtrf_206 }),
  .B({ S3582 }),
  .Y({ S3612 })
);
NAND #() 
NAND_2407_ (
  .A({ S3611 }),
  .B({ S3612 }),
  .Y({ S210 })
);
NAND #() 
NAND_2408_ (
  .A({ datapath_indatatrf_15 }),
  .B({ S3581 }),
  .Y({ S3613 })
);
NAND #() 
NAND_2409_ (
  .A({ datapath_theregisterfile_memtrf_207 }),
  .B({ S3582 }),
  .Y({ S3614 })
);
NAND #() 
NAND_2410_ (
  .A({ S3613 }),
  .B({ S3614 }),
  .Y({ S211 })
);
NOR #() 
NOR_947_ (
  .A({ S3228 }),
  .B({ S3580 }),
  .Y({ S3615 })
);
NAND #() 
NAND_2411_ (
  .A({ S3227 }),
  .B({ S3579 }),
  .Y({ S3616 })
);
NAND #() 
NAND_2412_ (
  .A({ datapath_indatatrf_0 }),
  .B({ S3615 }),
  .Y({ S3617 })
);
NAND #() 
NAND_2413_ (
  .A({ datapath_theregisterfile_memtrf_208 }),
  .B({ S3616 }),
  .Y({ S3618 })
);
NAND #() 
NAND_2414_ (
  .A({ S3617 }),
  .B({ S3618 }),
  .Y({ S212 })
);
NAND #() 
NAND_2415_ (
  .A({ datapath_indatatrf_1 }),
  .B({ S3615 }),
  .Y({ S3619 })
);
NAND #() 
NAND_2416_ (
  .A({ datapath_theregisterfile_memtrf_209 }),
  .B({ S3616 }),
  .Y({ S3620 })
);
NAND #() 
NAND_2417_ (
  .A({ S3619 }),
  .B({ S3620 }),
  .Y({ S213 })
);
NAND #() 
NAND_2418_ (
  .A({ datapath_indatatrf_2 }),
  .B({ S3615 }),
  .Y({ S3621 })
);
NAND #() 
NAND_2419_ (
  .A({ datapath_theregisterfile_memtrf_210 }),
  .B({ S3616 }),
  .Y({ S3622 })
);
NAND #() 
NAND_2420_ (
  .A({ S3621 }),
  .B({ S3622 }),
  .Y({ S214 })
);
NAND #() 
NAND_2421_ (
  .A({ datapath_indatatrf_3 }),
  .B({ S3615 }),
  .Y({ S3623 })
);
NAND #() 
NAND_2422_ (
  .A({ datapath_theregisterfile_memtrf_211 }),
  .B({ S3616 }),
  .Y({ S3624 })
);
NAND #() 
NAND_2423_ (
  .A({ S3623 }),
  .B({ S3624 }),
  .Y({ S215 })
);
NAND #() 
NAND_2424_ (
  .A({ datapath_indatatrf_4 }),
  .B({ S3615 }),
  .Y({ S3625 })
);
NAND #() 
NAND_2425_ (
  .A({ datapath_theregisterfile_memtrf_212 }),
  .B({ S3616 }),
  .Y({ S3626 })
);
NAND #() 
NAND_2426_ (
  .A({ S3625 }),
  .B({ S3626 }),
  .Y({ S216 })
);
NAND #() 
NAND_2427_ (
  .A({ datapath_indatatrf_5 }),
  .B({ S3615 }),
  .Y({ S3627 })
);
NAND #() 
NAND_2428_ (
  .A({ datapath_theregisterfile_memtrf_213 }),
  .B({ S3616 }),
  .Y({ S3628 })
);
NAND #() 
NAND_2429_ (
  .A({ S3627 }),
  .B({ S3628 }),
  .Y({ S217 })
);
NAND #() 
NAND_2430_ (
  .A({ datapath_indatatrf_6 }),
  .B({ S3615 }),
  .Y({ S3629 })
);
NAND #() 
NAND_2431_ (
  .A({ datapath_theregisterfile_memtrf_214 }),
  .B({ S3616 }),
  .Y({ S3630 })
);
NAND #() 
NAND_2432_ (
  .A({ S3629 }),
  .B({ S3630 }),
  .Y({ S218 })
);
NAND #() 
NAND_2433_ (
  .A({ datapath_indatatrf_7 }),
  .B({ S3615 }),
  .Y({ S3631 })
);
NAND #() 
NAND_2434_ (
  .A({ datapath_theregisterfile_memtrf_215 }),
  .B({ S3616 }),
  .Y({ S3632 })
);
NAND #() 
NAND_2435_ (
  .A({ S3631 }),
  .B({ S3632 }),
  .Y({ S219 })
);
NAND #() 
NAND_2436_ (
  .A({ datapath_indatatrf_8 }),
  .B({ S3615 }),
  .Y({ S3633 })
);
NAND #() 
NAND_2437_ (
  .A({ datapath_theregisterfile_memtrf_216 }),
  .B({ S3616 }),
  .Y({ S3634 })
);
NAND #() 
NAND_2438_ (
  .A({ S3633 }),
  .B({ S3634 }),
  .Y({ S220 })
);
NAND #() 
NAND_2439_ (
  .A({ datapath_indatatrf_9 }),
  .B({ S3615 }),
  .Y({ S3635 })
);
NAND #() 
NAND_2440_ (
  .A({ datapath_theregisterfile_memtrf_217 }),
  .B({ S3616 }),
  .Y({ S3636 })
);
NAND #() 
NAND_2441_ (
  .A({ S3635 }),
  .B({ S3636 }),
  .Y({ S221 })
);
NAND #() 
NAND_2442_ (
  .A({ datapath_indatatrf_10 }),
  .B({ S3615 }),
  .Y({ S3637 })
);
NAND #() 
NAND_2443_ (
  .A({ datapath_theregisterfile_memtrf_218 }),
  .B({ S3616 }),
  .Y({ S3638 })
);
NAND #() 
NAND_2444_ (
  .A({ S3637 }),
  .B({ S3638 }),
  .Y({ S222 })
);
NAND #() 
NAND_2445_ (
  .A({ datapath_indatatrf_11 }),
  .B({ S3615 }),
  .Y({ S3639 })
);
NAND #() 
NAND_2446_ (
  .A({ datapath_theregisterfile_memtrf_219 }),
  .B({ S3616 }),
  .Y({ S3640 })
);
NAND #() 
NAND_2447_ (
  .A({ S3639 }),
  .B({ S3640 }),
  .Y({ S223 })
);
NAND #() 
NAND_2448_ (
  .A({ datapath_indatatrf_12 }),
  .B({ S3615 }),
  .Y({ S3641 })
);
NAND #() 
NAND_2449_ (
  .A({ datapath_theregisterfile_memtrf_220 }),
  .B({ S3616 }),
  .Y({ S3642 })
);
NAND #() 
NAND_2450_ (
  .A({ S3641 }),
  .B({ S3642 }),
  .Y({ S224 })
);
NAND #() 
NAND_2451_ (
  .A({ datapath_indatatrf_13 }),
  .B({ S3615 }),
  .Y({ S3643 })
);
NAND #() 
NAND_2452_ (
  .A({ datapath_theregisterfile_memtrf_221 }),
  .B({ S3616 }),
  .Y({ S3644 })
);
NAND #() 
NAND_2453_ (
  .A({ S3643 }),
  .B({ S3644 }),
  .Y({ S225 })
);
NAND #() 
NAND_2454_ (
  .A({ datapath_indatatrf_14 }),
  .B({ S3615 }),
  .Y({ S3645 })
);
NAND #() 
NAND_2455_ (
  .A({ datapath_theregisterfile_memtrf_222 }),
  .B({ S3616 }),
  .Y({ S3646 })
);
NAND #() 
NAND_2456_ (
  .A({ S3645 }),
  .B({ S3646 }),
  .Y({ S226 })
);
NAND #() 
NAND_2457_ (
  .A({ datapath_indatatrf_15 }),
  .B({ S3615 }),
  .Y({ S3647 })
);
NAND #() 
NAND_2458_ (
  .A({ datapath_theregisterfile_memtrf_223 }),
  .B({ S3616 }),
  .Y({ S3648 })
);
NAND #() 
NAND_2459_ (
  .A({ S3647 }),
  .B({ S3648 }),
  .Y({ S227 })
);
NOR #() 
NOR_948_ (
  .A({ S3192 }),
  .B({ S3578 }),
  .Y({ S3649 })
);
NAND #() 
NAND_2460_ (
  .A({ S3191 }),
  .B({ S3577 }),
  .Y({ S3650 })
);
NAND #() 
NAND_2461_ (
  .A({ datapath_indatatrf_0 }),
  .B({ S3649 }),
  .Y({ S3651 })
);
NAND #() 
NAND_2462_ (
  .A({ datapath_theregisterfile_memtrf_224 }),
  .B({ S3650 }),
  .Y({ S3652 })
);
NAND #() 
NAND_2463_ (
  .A({ S3651 }),
  .B({ S3652 }),
  .Y({ S228 })
);
NAND #() 
NAND_2464_ (
  .A({ datapath_indatatrf_1 }),
  .B({ S3649 }),
  .Y({ S3653 })
);
NAND #() 
NAND_2465_ (
  .A({ datapath_theregisterfile_memtrf_225 }),
  .B({ S3650 }),
  .Y({ S3654 })
);
NAND #() 
NAND_2466_ (
  .A({ S3653 }),
  .B({ S3654 }),
  .Y({ S229 })
);
NAND #() 
NAND_2467_ (
  .A({ datapath_indatatrf_2 }),
  .B({ S3649 }),
  .Y({ S3655 })
);
NAND #() 
NAND_2468_ (
  .A({ datapath_theregisterfile_memtrf_226 }),
  .B({ S3650 }),
  .Y({ S3656 })
);
NAND #() 
NAND_2469_ (
  .A({ S3655 }),
  .B({ S3656 }),
  .Y({ S230 })
);
NAND #() 
NAND_2470_ (
  .A({ datapath_indatatrf_3 }),
  .B({ S3649 }),
  .Y({ S3657 })
);
NAND #() 
NAND_2471_ (
  .A({ datapath_theregisterfile_memtrf_227 }),
  .B({ S3650 }),
  .Y({ S3658 })
);
NAND #() 
NAND_2472_ (
  .A({ S3657 }),
  .B({ S3658 }),
  .Y({ S231 })
);
NAND #() 
NAND_2473_ (
  .A({ datapath_indatatrf_4 }),
  .B({ S3649 }),
  .Y({ S3659 })
);
NAND #() 
NAND_2474_ (
  .A({ datapath_theregisterfile_memtrf_228 }),
  .B({ S3650 }),
  .Y({ S3660 })
);
NAND #() 
NAND_2475_ (
  .A({ S3659 }),
  .B({ S3660 }),
  .Y({ S232 })
);
NAND #() 
NAND_2476_ (
  .A({ datapath_indatatrf_5 }),
  .B({ S3649 }),
  .Y({ S3661 })
);
NAND #() 
NAND_2477_ (
  .A({ datapath_theregisterfile_memtrf_229 }),
  .B({ S3650 }),
  .Y({ S3662 })
);
NAND #() 
NAND_2478_ (
  .A({ S3661 }),
  .B({ S3662 }),
  .Y({ S233 })
);
NAND #() 
NAND_2479_ (
  .A({ datapath_indatatrf_6 }),
  .B({ S3649 }),
  .Y({ S3663 })
);
NAND #() 
NAND_2480_ (
  .A({ datapath_theregisterfile_memtrf_230 }),
  .B({ S3650 }),
  .Y({ S3664 })
);
NAND #() 
NAND_2481_ (
  .A({ S3663 }),
  .B({ S3664 }),
  .Y({ S234 })
);
NAND #() 
NAND_2482_ (
  .A({ datapath_indatatrf_7 }),
  .B({ S3649 }),
  .Y({ S3665 })
);
NAND #() 
NAND_2483_ (
  .A({ datapath_theregisterfile_memtrf_231 }),
  .B({ S3650 }),
  .Y({ S3666 })
);
NAND #() 
NAND_2484_ (
  .A({ S3665 }),
  .B({ S3666 }),
  .Y({ S235 })
);
NAND #() 
NAND_2485_ (
  .A({ datapath_indatatrf_8 }),
  .B({ S3649 }),
  .Y({ S3667 })
);
NAND #() 
NAND_2486_ (
  .A({ datapath_theregisterfile_memtrf_232 }),
  .B({ S3650 }),
  .Y({ S3668 })
);
NAND #() 
NAND_2487_ (
  .A({ S3667 }),
  .B({ S3668 }),
  .Y({ S236 })
);
NAND #() 
NAND_2488_ (
  .A({ datapath_indatatrf_9 }),
  .B({ S3649 }),
  .Y({ S3669 })
);
NAND #() 
NAND_2489_ (
  .A({ datapath_theregisterfile_memtrf_233 }),
  .B({ S3650 }),
  .Y({ S3670 })
);
NAND #() 
NAND_2490_ (
  .A({ S3669 }),
  .B({ S3670 }),
  .Y({ S237 })
);
NAND #() 
NAND_2491_ (
  .A({ datapath_indatatrf_10 }),
  .B({ S3649 }),
  .Y({ S3671 })
);
NAND #() 
NAND_2492_ (
  .A({ datapath_theregisterfile_memtrf_234 }),
  .B({ S3650 }),
  .Y({ S3672 })
);
NAND #() 
NAND_2493_ (
  .A({ S3671 }),
  .B({ S3672 }),
  .Y({ S238 })
);
NAND #() 
NAND_2494_ (
  .A({ datapath_indatatrf_11 }),
  .B({ S3649 }),
  .Y({ S3673 })
);
NAND #() 
NAND_2495_ (
  .A({ datapath_theregisterfile_memtrf_235 }),
  .B({ S3650 }),
  .Y({ S3674 })
);
NAND #() 
NAND_2496_ (
  .A({ S3673 }),
  .B({ S3674 }),
  .Y({ S239 })
);
NAND #() 
NAND_2497_ (
  .A({ datapath_indatatrf_12 }),
  .B({ S3649 }),
  .Y({ S3675 })
);
NAND #() 
NAND_2498_ (
  .A({ datapath_theregisterfile_memtrf_236 }),
  .B({ S3650 }),
  .Y({ S3676 })
);
NAND #() 
NAND_2499_ (
  .A({ S3675 }),
  .B({ S3676 }),
  .Y({ S240 })
);
NAND #() 
NAND_2500_ (
  .A({ datapath_indatatrf_13 }),
  .B({ S3649 }),
  .Y({ S3677 })
);
NAND #() 
NAND_2501_ (
  .A({ datapath_theregisterfile_memtrf_237 }),
  .B({ S3650 }),
  .Y({ S3678 })
);
NAND #() 
NAND_2502_ (
  .A({ S3677 }),
  .B({ S3678 }),
  .Y({ S241 })
);
NAND #() 
NAND_2503_ (
  .A({ datapath_indatatrf_14 }),
  .B({ S3649 }),
  .Y({ S3679 })
);
NAND #() 
NAND_2504_ (
  .A({ datapath_theregisterfile_memtrf_238 }),
  .B({ S3650 }),
  .Y({ S3680 })
);
NAND #() 
NAND_2505_ (
  .A({ S3679 }),
  .B({ S3680 }),
  .Y({ S242 })
);
NAND #() 
NAND_2506_ (
  .A({ datapath_indatatrf_15 }),
  .B({ S3649 }),
  .Y({ S3681 })
);
NAND #() 
NAND_2507_ (
  .A({ datapath_theregisterfile_memtrf_239 }),
  .B({ S3650 }),
  .Y({ S3682 })
);
NAND #() 
NAND_2508_ (
  .A({ S3681 }),
  .B({ S3682 }),
  .Y({ S243 })
);
NOR #() 
NOR_949_ (
  .A({ S1857 }),
  .B({ S1962 }),
  .Y({ S3683 })
);
NOT #() 
NOT_318_ (
  .A({ S3683 }),
  .Y({ S3684 })
);
NOR #() 
NOR_950_ (
  .A({ S3046 }),
  .B({ S3150 }),
  .Y({ S3685 })
);
NAND #() 
NAND_2509_ (
  .A({ S2824 }),
  .B({ S3685 }),
  .Y({ S3686 })
);
NOR #() 
NOR_951_ (
  .A({ S2929 }),
  .B({ S3686 }),
  .Y({ S3687 })
);
NAND #() 
NAND_2510_ (
  .A({ S2626 }),
  .B({ S2724 }),
  .Y({ S3688 })
);
NOT #() 
NOT_319_ (
  .A({ S3688 }),
  .Y({ S3689 })
);
NOR #() 
NOR_952_ (
  .A({ S2424 }),
  .B({ S3688 }),
  .Y({ S3690 })
);
NOT #() 
NOT_320_ (
  .A({ S3690 }),
  .Y({ S3691 })
);
NAND #() 
NAND_2511_ (
  .A({ S2525 }),
  .B({ S3687 }),
  .Y({ S3692 })
);
NOR #() 
NOR_953_ (
  .A({ S3691 }),
  .B({ S3692 }),
  .Y({ S3693 })
);
NOR #() 
NOR_954_ (
  .A({ S2011 }),
  .B({ S2113 }),
  .Y({ S3694 })
);
NAND #() 
NAND_2512_ (
  .A({ S1754 }),
  .B({ S3694 }),
  .Y({ S3695 })
);
NAND #() 
NAND_2513_ (
  .A({ S1522 }),
  .B({ S3683 }),
  .Y({ S3696 })
);
NOR #() 
NOR_955_ (
  .A({ S3695 }),
  .B({ S3696 }),
  .Y({ S3697 })
);
NAND #() 
NAND_2514_ (
  .A({ S3693 }),
  .B({ S3697 }),
  .Y({ S3698 })
);
NOR #() 
NOR_956_ (
  .A({ S2435 }),
  .B({ S3698 }),
  .Y({ S3699 })
);
NOR #() 
NOR_957_ (
  .A({ S1405 }),
  .B({ S3699 }),
  .Y({ S3700 })
);
NOR #() 
NOR_958_ (
  .A({ controller_389_B_0 }),
  .B({ S1404 }),
  .Y({ S3701 })
);
NOR #() 
NOR_959_ (
  .A({ S3700 }),
  .B({ S3701 }),
  .Y({ S264 })
);
NAND #() 
NAND_2515_ (
  .A({ controller_389_B_2 }),
  .B({ S1405 }),
  .Y({ S3702 })
);
NAND #() 
NAND_2516_ (
  .A({ S2211 }),
  .B({ S2319 }),
  .Y({ S3703 })
);
NOR #() 
NOR_960_ (
  .A({ S1853 }),
  .B({ S1958 }),
  .Y({ S3704 })
);
NOR #() 
NOR_961_ (
  .A({ S1957 }),
  .B({ S3704 }),
  .Y({ S3705 })
);
NAND #() 
NAND_2517_ (
  .A({ S1521 }),
  .B({ S1752 }),
  .Y({ S3706 })
);
NAND #() 
NAND_2518_ (
  .A({ S1751 }),
  .B({ S3706 }),
  .Y({ S3707 })
);
NOR #() 
NOR_962_ (
  .A({ S3684 }),
  .B({ S3707 }),
  .Y({ S3708 })
);
NOR #() 
NOR_963_ (
  .A({ S3705 }),
  .B({ S3708 }),
  .Y({ S3709 })
);
NOR #() 
NOR_964_ (
  .A({ S2007 }),
  .B({ S3709 }),
  .Y({ S3710 })
);
NAND #() 
NAND_2519_ (
  .A({ S2010 }),
  .B({ S2112 }),
  .Y({ S3711 })
);
NOR #() 
NOR_965_ (
  .A({ S3710 }),
  .B({ S3711 }),
  .Y({ S3712 })
);
NOR #() 
NOR_966_ (
  .A({ S2435 }),
  .B({ S3712 }),
  .Y({ S3713 })
);
NAND #() 
NAND_2520_ (
  .A({ S2111 }),
  .B({ S3713 }),
  .Y({ S3714 })
);
NAND #() 
NAND_2521_ (
  .A({ S2317 }),
  .B({ S3703 }),
  .Y({ S3715 })
);
NAND #() 
NAND_2522_ (
  .A({ S3714 }),
  .B({ S3715 }),
  .Y({ S3716 })
);
NAND #() 
NAND_2523_ (
  .A({ S3693 }),
  .B({ S3716 }),
  .Y({ S3717 })
);
NOT #() 
NOT_321_ (
  .A({ S3717 }),
  .Y({ S3718 })
);
NOR #() 
NOR_967_ (
  .A({ S2422 }),
  .B({ S2524 }),
  .Y({ S3719 })
);
NOR #() 
NOR_968_ (
  .A({ S2523 }),
  .B({ S3719 }),
  .Y({ S3720 })
);
NAND #() 
NAND_2524_ (
  .A({ S3689 }),
  .B({ S3720 }),
  .Y({ S3721 })
);
NOR #() 
NOR_969_ (
  .A({ S2622 }),
  .B({ S2722 }),
  .Y({ S3722 })
);
NOR #() 
NOR_970_ (
  .A({ S2723 }),
  .B({ S3722 }),
  .Y({ S3723 })
);
NAND #() 
NAND_2525_ (
  .A({ S3721 }),
  .B({ S3723 }),
  .Y({ S3724 })
);
NAND #() 
NAND_2526_ (
  .A({ S3687 }),
  .B({ S3724 }),
  .Y({ S3725 })
);
NOR #() 
NOR_971_ (
  .A({ S2823 }),
  .B({ S2927 }),
  .Y({ S3726 })
);
NOR #() 
NOR_972_ (
  .A({ S2925 }),
  .B({ S3726 }),
  .Y({ S3727 })
);
NAND #() 
NAND_2527_ (
  .A({ S3685 }),
  .B({ S3727 }),
  .Y({ S3728 })
);
NOR #() 
NOR_973_ (
  .A({ S3043 }),
  .B({ S3148 }),
  .Y({ S3729 })
);
NOR #() 
NOR_974_ (
  .A({ S3146 }),
  .B({ S3729 }),
  .Y({ S3730 })
);
NAND #() 
NAND_2528_ (
  .A({ S3728 }),
  .B({ S3730 }),
  .Y({ S3731 })
);
NOR #() 
NOR_975_ (
  .A({ S3718 }),
  .B({ S3731 }),
  .Y({ S3732 })
);
NAND #() 
NAND_2529_ (
  .A({ S3725 }),
  .B({ S3732 }),
  .Y({ S3733 })
);
NAND #() 
NAND_2530_ (
  .A({ S3700 }),
  .B({ S3733 }),
  .Y({ S3734 })
);
NAND #() 
NAND_2531_ (
  .A({ S3702 }),
  .B({ S3734 }),
  .Y({ S265 })
);
NAND #() 
NAND_2532_ (
  .A({ datapath_muxmem_in2_0 }),
  .B({ S8580 }),
  .Y({ S3735 })
);
NOR #() 
NOR_976_ (
  .A({ datapath_muxmem_in2_0 }),
  .B({ S1222 }),
  .Y({ S3736 })
);
NOR #() 
NOR_977_ (
  .A({ S364 }),
  .B({ S3736 }),
  .Y({ S3737 })
);
NAND #() 
NAND_2533_ (
  .A({ S1223 }),
  .B({ S3737 }),
  .Y({ S3738 })
);
NOR #() 
NOR_978_ (
  .A({ datapath_muxmem_in2_0 }),
  .B({ S1334 }),
  .Y({ S3739 })
);
NOR #() 
NOR_979_ (
  .A({ S1370 }),
  .B({ S3739 }),
  .Y({ S3740 })
);
NAND #() 
NAND_2534_ (
  .A({ S3738 }),
  .B({ S3740 }),
  .Y({ S3741 })
);
NOR #() 
NOR_980_ (
  .A({ datapath_addsubunit_in1_0 }),
  .B({ S1371 }),
  .Y({ S3742 })
);
NOR #() 
NOR_981_ (
  .A({ S8580 }),
  .B({ S3742 }),
  .Y({ S3743 })
);
NAND #() 
NAND_2535_ (
  .A({ S3741 }),
  .B({ S3743 }),
  .Y({ S3744 })
);
NAND #() 
NAND_2536_ (
  .A({ S3735 }),
  .B({ S3744 }),
  .Y({ S267 })
);
NAND #() 
NAND_2537_ (
  .A({ datapath_muxmem_in2_1 }),
  .B({ S8580 }),
  .Y({ S3745 })
);
NOR #() 
NOR_982_ (
  .A({ S1224 }),
  .B({ S1226 }),
  .Y({ S3746 })
);
NOR #() 
NOR_983_ (
  .A({ S1228 }),
  .B({ S3746 }),
  .Y({ S3747 })
);
NAND #() 
NAND_2538_ (
  .A({ S365 }),
  .B({ S3747 }),
  .Y({ S3748 })
);
NOR #() 
NOR_984_ (
  .A({ S1334 }),
  .B({ S1774 }),
  .Y({ S3749 })
);
NOR #() 
NOR_985_ (
  .A({ S1370 }),
  .B({ S3749 }),
  .Y({ S3750 })
);
NAND #() 
NAND_2539_ (
  .A({ S3748 }),
  .B({ S3750 }),
  .Y({ S3751 })
);
NOR #() 
NOR_986_ (
  .A({ datapath_addsubunit_in1_1 }),
  .B({ S1371 }),
  .Y({ S3752 })
);
NOR #() 
NOR_987_ (
  .A({ S8580 }),
  .B({ S3752 }),
  .Y({ S3753 })
);
NAND #() 
NAND_2540_ (
  .A({ S3751 }),
  .B({ S3753 }),
  .Y({ S3754 })
);
NAND #() 
NAND_2541_ (
  .A({ S3745 }),
  .B({ S3754 }),
  .Y({ S268 })
);
NAND #() 
NAND_2542_ (
  .A({ datapath_muxmem_in2_2 }),
  .B({ S8580 }),
  .Y({ S3755 })
);
NOR #() 
NOR_988_ (
  .A({ S1229 }),
  .B({ S1231 }),
  .Y({ S3756 })
);
NOR #() 
NOR_989_ (
  .A({ S364 }),
  .B({ S3756 }),
  .Y({ S3757 })
);
NAND #() 
NAND_2543_ (
  .A({ S1232 }),
  .B({ S3757 }),
  .Y({ S3758 })
);
NOR #() 
NOR_990_ (
  .A({ S1334 }),
  .B({ S1875 }),
  .Y({ S3759 })
);
NOR #() 
NOR_991_ (
  .A({ S1370 }),
  .B({ S3759 }),
  .Y({ S3760 })
);
NAND #() 
NAND_2544_ (
  .A({ S3758 }),
  .B({ S3760 }),
  .Y({ S3761 })
);
NOR #() 
NOR_992_ (
  .A({ datapath_addsubunit_in1_2 }),
  .B({ S1371 }),
  .Y({ S3762 })
);
NOR #() 
NOR_993_ (
  .A({ S8580 }),
  .B({ S3762 }),
  .Y({ S3763 })
);
NAND #() 
NAND_2545_ (
  .A({ S3761 }),
  .B({ S3763 }),
  .Y({ S3764 })
);
NAND #() 
NAND_2546_ (
  .A({ S3755 }),
  .B({ S3764 }),
  .Y({ S269 })
);
NAND #() 
NAND_2547_ (
  .A({ datapath_muxmem_in2_3 }),
  .B({ S8580 }),
  .Y({ S3765 })
);
NOR #() 
NOR_994_ (
  .A({ S1069 }),
  .B({ S1070 }),
  .Y({ S3766 })
);
NAND #() 
NAND_2548_ (
  .A({ S1233 }),
  .B({ S3766 }),
  .Y({ S3767 })
);
NOR #() 
NOR_995_ (
  .A({ S1233 }),
  .B({ S3766 }),
  .Y({ S3768 })
);
NOR #() 
NOR_996_ (
  .A({ S364 }),
  .B({ S3768 }),
  .Y({ S3769 })
);
NAND #() 
NAND_2549_ (
  .A({ S3767 }),
  .B({ S3769 }),
  .Y({ S3770 })
);
NOR #() 
NOR_997_ (
  .A({ S1334 }),
  .B({ S1978 }),
  .Y({ S3771 })
);
NOR #() 
NOR_998_ (
  .A({ S1370 }),
  .B({ S3771 }),
  .Y({ S3772 })
);
NAND #() 
NAND_2550_ (
  .A({ S3770 }),
  .B({ S3772 }),
  .Y({ S3773 })
);
NOR #() 
NOR_999_ (
  .A({ datapath_addsubunit_in1_3 }),
  .B({ S1371 }),
  .Y({ S3774 })
);
NOR #() 
NOR_1000_ (
  .A({ S8580 }),
  .B({ S3774 }),
  .Y({ S3775 })
);
NAND #() 
NAND_2551_ (
  .A({ S3773 }),
  .B({ S3775 }),
  .Y({ S3776 })
);
NAND #() 
NAND_2552_ (
  .A({ S3765 }),
  .B({ S3776 }),
  .Y({ S270 })
);
NAND #() 
NAND_2553_ (
  .A({ datapath_muxmem_in2_4 }),
  .B({ S8580 }),
  .Y({ S3777 })
);
NOR #() 
NOR_1001_ (
  .A({ S1019 }),
  .B({ S1235 }),
  .Y({ S3778 })
);
NOR #() 
NOR_1002_ (
  .A({ S1334 }),
  .B({ S2029 }),
  .Y({ S3779 })
);
NOR #() 
NOR_1003_ (
  .A({ S364 }),
  .B({ S3778 }),
  .Y({ S3780 })
);
NAND #() 
NAND_2554_ (
  .A({ S1236 }),
  .B({ S3780 }),
  .Y({ S3781 })
);
NOT #() 
NOT_322_ (
  .A({ S3781 }),
  .Y({ S3782 })
);
NOR #() 
NOR_1004_ (
  .A({ S3779 }),
  .B({ S3782 }),
  .Y({ S3783 })
);
NAND #() 
NAND_2555_ (
  .A({ S1371 }),
  .B({ S3783 }),
  .Y({ S3784 })
);
NOR #() 
NOR_1005_ (
  .A({ datapath_addsubunit_in1_4 }),
  .B({ S1371 }),
  .Y({ S3785 })
);
NOR #() 
NOR_1006_ (
  .A({ S8580 }),
  .B({ S3785 }),
  .Y({ S3786 })
);
NAND #() 
NAND_2556_ (
  .A({ S3784 }),
  .B({ S3786 }),
  .Y({ S3787 })
);
NAND #() 
NAND_2557_ (
  .A({ S3777 }),
  .B({ S3787 }),
  .Y({ S271 })
);
NAND #() 
NAND_2558_ (
  .A({ datapath_muxmem_in2_5 }),
  .B({ S8580 }),
  .Y({ S3788 })
);
NOR #() 
NOR_1007_ (
  .A({ S967 }),
  .B({ S968 }),
  .Y({ S3789 })
);
NAND #() 
NAND_2559_ (
  .A({ S1237 }),
  .B({ S3789 }),
  .Y({ S3790 })
);
NOR #() 
NOR_1008_ (
  .A({ S1237 }),
  .B({ S3789 }),
  .Y({ S3791 })
);
NOR #() 
NOR_1009_ (
  .A({ S364 }),
  .B({ S3791 }),
  .Y({ S3792 })
);
NAND #() 
NAND_2560_ (
  .A({ S3790 }),
  .B({ S3792 }),
  .Y({ S3793 })
);
NOR #() 
NOR_1010_ (
  .A({ S1334 }),
  .B({ S2136 }),
  .Y({ S3794 })
);
NOR #() 
NOR_1011_ (
  .A({ S1370 }),
  .B({ S3794 }),
  .Y({ S3795 })
);
NAND #() 
NAND_2561_ (
  .A({ S3793 }),
  .B({ S3795 }),
  .Y({ S3796 })
);
NOR #() 
NOR_1012_ (
  .A({ datapath_addsubunit_in1_5 }),
  .B({ S1371 }),
  .Y({ S3797 })
);
NOR #() 
NOR_1013_ (
  .A({ S8580 }),
  .B({ S3797 }),
  .Y({ S3798 })
);
NAND #() 
NAND_2562_ (
  .A({ S3796 }),
  .B({ S3798 }),
  .Y({ S3799 })
);
NAND #() 
NAND_2563_ (
  .A({ S3788 }),
  .B({ S3799 }),
  .Y({ S272 })
);
NAND #() 
NAND_2564_ (
  .A({ datapath_muxmem_in2_6 }),
  .B({ S8580 }),
  .Y({ S3800 })
);
NOR #() 
NOR_1014_ (
  .A({ S916 }),
  .B({ S1239 }),
  .Y({ S3801 })
);
NOR #() 
NOR_1015_ (
  .A({ S364 }),
  .B({ S3801 }),
  .Y({ S3802 })
);
NAND #() 
NAND_2565_ (
  .A({ S1240 }),
  .B({ S3802 }),
  .Y({ S3803 })
);
NOR #() 
NOR_1016_ (
  .A({ S1334 }),
  .B({ S2235 }),
  .Y({ S3804 })
);
NOR #() 
NOR_1017_ (
  .A({ S1370 }),
  .B({ S3804 }),
  .Y({ S3805 })
);
NAND #() 
NAND_2566_ (
  .A({ S3803 }),
  .B({ S3805 }),
  .Y({ S3806 })
);
NOR #() 
NOR_1018_ (
  .A({ datapath_addsubunit_in1_6 }),
  .B({ S1371 }),
  .Y({ S3807 })
);
NOR #() 
NOR_1019_ (
  .A({ S8580 }),
  .B({ S3807 }),
  .Y({ S3808 })
);
NAND #() 
NAND_2567_ (
  .A({ S3806 }),
  .B({ S3808 }),
  .Y({ S3809 })
);
NAND #() 
NAND_2568_ (
  .A({ S3800 }),
  .B({ S3809 }),
  .Y({ S273 })
);
NAND #() 
NAND_2569_ (
  .A({ datapath_muxmem_in2_7 }),
  .B({ S8580 }),
  .Y({ S3810 })
);
NOR #() 
NOR_1020_ (
  .A({ S862 }),
  .B({ S863 }),
  .Y({ S3811 })
);
NAND #() 
NAND_2570_ (
  .A({ S1241 }),
  .B({ S3811 }),
  .Y({ S3812 })
);
NOR #() 
NOR_1021_ (
  .A({ S1241 }),
  .B({ S3811 }),
  .Y({ S3813 })
);
NOR #() 
NOR_1022_ (
  .A({ S364 }),
  .B({ S3813 }),
  .Y({ S3814 })
);
NAND #() 
NAND_2571_ (
  .A({ S3812 }),
  .B({ S3814 }),
  .Y({ S3815 })
);
NOR #() 
NOR_1023_ (
  .A({ S1334 }),
  .B({ S2331 }),
  .Y({ S3816 })
);
NOR #() 
NOR_1024_ (
  .A({ S1370 }),
  .B({ S3816 }),
  .Y({ S3817 })
);
NAND #() 
NAND_2572_ (
  .A({ S3815 }),
  .B({ S3817 }),
  .Y({ S3818 })
);
NOR #() 
NOR_1025_ (
  .A({ datapath_addsubunit_in1_7 }),
  .B({ S1371 }),
  .Y({ S3819 })
);
NOR #() 
NOR_1026_ (
  .A({ S8580 }),
  .B({ S3819 }),
  .Y({ S3820 })
);
NAND #() 
NAND_2573_ (
  .A({ S3818 }),
  .B({ S3820 }),
  .Y({ S3821 })
);
NAND #() 
NAND_2574_ (
  .A({ S3810 }),
  .B({ S3821 }),
  .Y({ S274 })
);
NAND #() 
NAND_2575_ (
  .A({ datapath_muxmem_in2_8 }),
  .B({ S8580 }),
  .Y({ S3822 })
);
NOR #() 
NOR_1027_ (
  .A({ S811 }),
  .B({ S1243 }),
  .Y({ S3823 })
);
NOR #() 
NOR_1028_ (
  .A({ S364 }),
  .B({ S3823 }),
  .Y({ S3824 })
);
NAND #() 
NAND_2576_ (
  .A({ S1244 }),
  .B({ S3824 }),
  .Y({ S3825 })
);
NOR #() 
NOR_1029_ (
  .A({ S1334 }),
  .B({ S2449 }),
  .Y({ S3826 })
);
NOR #() 
NOR_1030_ (
  .A({ S1370 }),
  .B({ S3826 }),
  .Y({ S3827 })
);
NAND #() 
NAND_2577_ (
  .A({ S3825 }),
  .B({ S3827 }),
  .Y({ S3828 })
);
NOR #() 
NOR_1031_ (
  .A({ datapath_addsubunit_in1_8 }),
  .B({ S1371 }),
  .Y({ S3829 })
);
NOR #() 
NOR_1032_ (
  .A({ S8580 }),
  .B({ S3829 }),
  .Y({ S3830 })
);
NAND #() 
NAND_2578_ (
  .A({ S3828 }),
  .B({ S3830 }),
  .Y({ S3831 })
);
NAND #() 
NAND_2579_ (
  .A({ S3822 }),
  .B({ S3831 }),
  .Y({ S275 })
);
NAND #() 
NAND_2580_ (
  .A({ datapath_muxmem_in2_9 }),
  .B({ S8580 }),
  .Y({ S3832 })
);
NOR #() 
NOR_1033_ (
  .A({ S758 }),
  .B({ S759 }),
  .Y({ S3833 })
);
NAND #() 
NAND_2581_ (
  .A({ S1245 }),
  .B({ S3833 }),
  .Y({ S3834 })
);
NOR #() 
NOR_1034_ (
  .A({ S1245 }),
  .B({ S3833 }),
  .Y({ S3835 })
);
NOR #() 
NOR_1035_ (
  .A({ S364 }),
  .B({ S3835 }),
  .Y({ S3836 })
);
NAND #() 
NAND_2582_ (
  .A({ S3834 }),
  .B({ S3836 }),
  .Y({ S3837 })
);
NOR #() 
NOR_1036_ (
  .A({ S1334 }),
  .B({ S2551 }),
  .Y({ S3838 })
);
NOR #() 
NOR_1037_ (
  .A({ S1370 }),
  .B({ S3838 }),
  .Y({ S3839 })
);
NAND #() 
NAND_2583_ (
  .A({ S3837 }),
  .B({ S3839 }),
  .Y({ S3840 })
);
NOR #() 
NOR_1038_ (
  .A({ datapath_addsubunit_in1_9 }),
  .B({ S1371 }),
  .Y({ S3841 })
);
NOR #() 
NOR_1039_ (
  .A({ S8580 }),
  .B({ S3841 }),
  .Y({ S3842 })
);
NAND #() 
NAND_2584_ (
  .A({ S3840 }),
  .B({ S3842 }),
  .Y({ S3843 })
);
NAND #() 
NAND_2585_ (
  .A({ S3832 }),
  .B({ S3843 }),
  .Y({ S276 })
);
NAND #() 
NAND_2586_ (
  .A({ datapath_muxmem_in2_10 }),
  .B({ S8580 }),
  .Y({ S3844 })
);
NOR #() 
NOR_1040_ (
  .A({ S708 }),
  .B({ S1247 }),
  .Y({ S3845 })
);
NOR #() 
NOR_1041_ (
  .A({ S364 }),
  .B({ S3845 }),
  .Y({ S3846 })
);
NAND #() 
NAND_2587_ (
  .A({ S1248 }),
  .B({ S3846 }),
  .Y({ S3847 })
);
NOR #() 
NOR_1042_ (
  .A({ S1334 }),
  .B({ S2646 }),
  .Y({ S3848 })
);
NOR #() 
NOR_1043_ (
  .A({ S1370 }),
  .B({ S3848 }),
  .Y({ S3849 })
);
NAND #() 
NAND_2588_ (
  .A({ S3847 }),
  .B({ S3849 }),
  .Y({ S3850 })
);
NOR #() 
NOR_1044_ (
  .A({ datapath_addsubunit_in1_10 }),
  .B({ S1371 }),
  .Y({ S3851 })
);
NOR #() 
NOR_1045_ (
  .A({ S8580 }),
  .B({ S3851 }),
  .Y({ S3852 })
);
NAND #() 
NAND_2589_ (
  .A({ S3850 }),
  .B({ S3852 }),
  .Y({ S3853 })
);
NAND #() 
NAND_2590_ (
  .A({ S3844 }),
  .B({ S3853 }),
  .Y({ S277 })
);
NAND #() 
NAND_2591_ (
  .A({ datapath_muxmem_in2_11 }),
  .B({ S8580 }),
  .Y({ S3854 })
);
NOR #() 
NOR_1046_ (
  .A({ S655 }),
  .B({ S656 }),
  .Y({ S3855 })
);
NAND #() 
NAND_2592_ (
  .A({ S1249 }),
  .B({ S3855 }),
  .Y({ S3856 })
);
NOR #() 
NOR_1047_ (
  .A({ S1249 }),
  .B({ S3855 }),
  .Y({ S3857 })
);
NOR #() 
NOR_1048_ (
  .A({ S364 }),
  .B({ S3857 }),
  .Y({ S3858 })
);
NAND #() 
NAND_2593_ (
  .A({ S3856 }),
  .B({ S3858 }),
  .Y({ S3859 })
);
NOR #() 
NOR_1049_ (
  .A({ S1334 }),
  .B({ S2748 }),
  .Y({ S3860 })
);
NOR #() 
NOR_1050_ (
  .A({ S1370 }),
  .B({ S3860 }),
  .Y({ S3861 })
);
NAND #() 
NAND_2594_ (
  .A({ S3859 }),
  .B({ S3861 }),
  .Y({ S3862 })
);
NOR #() 
NOR_1051_ (
  .A({ datapath_addsubunit_in1_11 }),
  .B({ S1371 }),
  .Y({ S3863 })
);
NOR #() 
NOR_1052_ (
  .A({ S8580 }),
  .B({ S3863 }),
  .Y({ S3864 })
);
NAND #() 
NAND_2595_ (
  .A({ S3862 }),
  .B({ S3864 }),
  .Y({ S3865 })
);
NAND #() 
NAND_2596_ (
  .A({ S3854 }),
  .B({ S3865 }),
  .Y({ S278 })
);
NAND #() 
NAND_2597_ (
  .A({ datapath_muxmem_in2_12 }),
  .B({ S8580 }),
  .Y({ S3866 })
);
NOR #() 
NOR_1053_ (
  .A({ S605 }),
  .B({ S1251 }),
  .Y({ S3867 })
);
NOR #() 
NOR_1054_ (
  .A({ S364 }),
  .B({ S3867 }),
  .Y({ S3868 })
);
NAND #() 
NAND_2598_ (
  .A({ S1252 }),
  .B({ S3868 }),
  .Y({ S3869 })
);
NOR #() 
NOR_1055_ (
  .A({ S1334 }),
  .B({ S2847 }),
  .Y({ S3870 })
);
NOR #() 
NOR_1056_ (
  .A({ S1370 }),
  .B({ S3870 }),
  .Y({ S3871 })
);
NAND #() 
NAND_2599_ (
  .A({ S3869 }),
  .B({ S3871 }),
  .Y({ S3872 })
);
NOR #() 
NOR_1057_ (
  .A({ datapath_addsubunit_in1_12 }),
  .B({ S1371 }),
  .Y({ S3873 })
);
NOR #() 
NOR_1058_ (
  .A({ S8580 }),
  .B({ S3873 }),
  .Y({ S3874 })
);
NAND #() 
NAND_2600_ (
  .A({ S3872 }),
  .B({ S3874 }),
  .Y({ S3875 })
);
NAND #() 
NAND_2601_ (
  .A({ S3866 }),
  .B({ S3875 }),
  .Y({ S279 })
);
NAND #() 
NAND_2602_ (
  .A({ datapath_muxmem_in2_13 }),
  .B({ S8580 }),
  .Y({ S3876 })
);
NOR #() 
NOR_1059_ (
  .A({ S552 }),
  .B({ S553 }),
  .Y({ S3877 })
);
NAND #() 
NAND_2603_ (
  .A({ S1253 }),
  .B({ S3877 }),
  .Y({ S3878 })
);
NOR #() 
NOR_1060_ (
  .A({ S1253 }),
  .B({ S3877 }),
  .Y({ S3879 })
);
NOR #() 
NOR_1061_ (
  .A({ S364 }),
  .B({ S3879 }),
  .Y({ S3880 })
);
NAND #() 
NAND_2604_ (
  .A({ S3878 }),
  .B({ S3880 }),
  .Y({ S3881 })
);
NOR #() 
NOR_1062_ (
  .A({ S1334 }),
  .B({ S2956 }),
  .Y({ S3882 })
);
NOR #() 
NOR_1063_ (
  .A({ S1370 }),
  .B({ S3882 }),
  .Y({ S3883 })
);
NAND #() 
NAND_2605_ (
  .A({ S3881 }),
  .B({ S3883 }),
  .Y({ S3884 })
);
NOR #() 
NOR_1064_ (
  .A({ datapath_addsubunit_in1_13 }),
  .B({ S1371 }),
  .Y({ S3885 })
);
NOR #() 
NOR_1065_ (
  .A({ S8580 }),
  .B({ S3885 }),
  .Y({ S3886 })
);
NAND #() 
NAND_2606_ (
  .A({ S3884 }),
  .B({ S3886 }),
  .Y({ S3887 })
);
NAND #() 
NAND_2607_ (
  .A({ S3876 }),
  .B({ S3887 }),
  .Y({ S280 })
);
NAND #() 
NAND_2608_ (
  .A({ datapath_muxmem_in2_14 }),
  .B({ S8580 }),
  .Y({ S3888 })
);
NOR #() 
NOR_1066_ (
  .A({ S502 }),
  .B({ S1255 }),
  .Y({ S3889 })
);
NOR #() 
NOR_1067_ (
  .A({ S364 }),
  .B({ S3889 }),
  .Y({ S3890 })
);
NAND #() 
NAND_2609_ (
  .A({ S1256 }),
  .B({ S3890 }),
  .Y({ S3891 })
);
NOR #() 
NOR_1068_ (
  .A({ S1334 }),
  .B({ S3066 }),
  .Y({ S3892 })
);
NOR #() 
NOR_1069_ (
  .A({ S1370 }),
  .B({ S3892 }),
  .Y({ S3893 })
);
NAND #() 
NAND_2610_ (
  .A({ S3891 }),
  .B({ S3893 }),
  .Y({ S3894 })
);
NOR #() 
NOR_1070_ (
  .A({ datapath_addsubunit_in1_14 }),
  .B({ S1371 }),
  .Y({ S3895 })
);
NOR #() 
NOR_1071_ (
  .A({ S8580 }),
  .B({ S3895 }),
  .Y({ S3896 })
);
NAND #() 
NAND_2611_ (
  .A({ S3894 }),
  .B({ S3896 }),
  .Y({ S3897 })
);
NAND #() 
NAND_2612_ (
  .A({ S3888 }),
  .B({ S3897 }),
  .Y({ S281 })
);
NOR #() 
NOR_1072_ (
  .A({ S8557 }),
  .B({ S377 }),
  .Y({ S3898 })
);
NAND #() 
NAND_2613_ (
  .A({ S8556 }),
  .B({ S376 }),
  .Y({ S3899 })
);
NOR #() 
NOR_1073_ (
  .A({ S3036 }),
  .B({ S3141 }),
  .Y({ S3900 })
);
NAND #() 
NAND_2614_ (
  .A({ S3037 }),
  .B({ S3142 }),
  .Y({ S3901 })
);
NOR #() 
NOR_1074_ (
  .A({ S2919 }),
  .B({ S3901 }),
  .Y({ S3902 })
);
NAND #() 
NAND_2615_ (
  .A({ S2920 }),
  .B({ S3900 }),
  .Y({ S3903 })
);
NOR #() 
NOR_1075_ (
  .A({ S2816 }),
  .B({ S3903 }),
  .Y({ S3904 })
);
NAND #() 
NAND_2616_ (
  .A({ S2817 }),
  .B({ S3902 }),
  .Y({ S3905 })
);
NOR #() 
NOR_1076_ (
  .A({ S2717 }),
  .B({ S3905 }),
  .Y({ S3906 })
);
NAND #() 
NAND_2617_ (
  .A({ S2718 }),
  .B({ S3904 }),
  .Y({ S3907 })
);
NOR #() 
NOR_1077_ (
  .A({ S2617 }),
  .B({ S3907 }),
  .Y({ S3908 })
);
NAND #() 
NAND_2618_ (
  .A({ S2618 }),
  .B({ S3906 }),
  .Y({ S3909 })
);
NOR #() 
NOR_1078_ (
  .A({ S2517 }),
  .B({ S3909 }),
  .Y({ S3910 })
);
NAND #() 
NAND_2619_ (
  .A({ S2518 }),
  .B({ S3908 }),
  .Y({ S3911 })
);
NOR #() 
NOR_1079_ (
  .A({ S2417 }),
  .B({ S3911 }),
  .Y({ S3912 })
);
NAND #() 
NAND_2620_ (
  .A({ S2418 }),
  .B({ S3910 }),
  .Y({ S3913 })
);
NOR #() 
NOR_1080_ (
  .A({ S2311 }),
  .B({ S3913 }),
  .Y({ S3914 })
);
NAND #() 
NAND_2621_ (
  .A({ S2312 }),
  .B({ S3912 }),
  .Y({ S3915 })
);
NOR #() 
NOR_1081_ (
  .A({ S2205 }),
  .B({ S3915 }),
  .Y({ S3916 })
);
NAND #() 
NAND_2622_ (
  .A({ S2206 }),
  .B({ S3914 }),
  .Y({ S3917 })
);
NOR #() 
NOR_1082_ (
  .A({ S2106 }),
  .B({ S3917 }),
  .Y({ S3918 })
);
NAND #() 
NAND_2623_ (
  .A({ S2107 }),
  .B({ S3916 }),
  .Y({ S3919 })
);
NOR #() 
NOR_1083_ (
  .A({ S1597 }),
  .B({ S3919 }),
  .Y({ S3920 })
);
NAND #() 
NAND_2624_ (
  .A({ S1598 }),
  .B({ S3918 }),
  .Y({ S3921 })
);
NOR #() 
NOR_1084_ (
  .A({ S1952 }),
  .B({ S3921 }),
  .Y({ S3922 })
);
NAND #() 
NAND_2625_ (
  .A({ S1953 }),
  .B({ S3920 }),
  .Y({ S3923 })
);
NOR #() 
NOR_1085_ (
  .A({ S1848 }),
  .B({ S3923 }),
  .Y({ S3924 })
);
NAND #() 
NAND_2626_ (
  .A({ S1849 }),
  .B({ S3922 }),
  .Y({ S3925 })
);
NOR #() 
NOR_1086_ (
  .A({ S1745 }),
  .B({ S3925 }),
  .Y({ S3926 })
);
NAND #() 
NAND_2627_ (
  .A({ S1746 }),
  .B({ S3924 }),
  .Y({ S3927 })
);
NOR #() 
NOR_1087_ (
  .A({ S1516 }),
  .B({ S3927 }),
  .Y({ S3928 })
);
NAND #() 
NAND_2628_ (
  .A({ S1515 }),
  .B({ S3926 }),
  .Y({ S3929 })
);
NOR #() 
NOR_1088_ (
  .A({ S1304 }),
  .B({ S3928 }),
  .Y({ S3930 })
);
NAND #() 
NAND_2629_ (
  .A({ datapath_addsubunit_in1_15 }),
  .B({ S3929 }),
  .Y({ S3931 })
);
NOR #() 
NOR_1089_ (
  .A({ S1745 }),
  .B({ S3931 }),
  .Y({ S3932 })
);
NAND #() 
NAND_2630_ (
  .A({ S1746 }),
  .B({ S3930 }),
  .Y({ S3933 })
);
NOR #() 
NOR_1090_ (
  .A({ datapath_addsubunit_in1_15 }),
  .B({ S1746 }),
  .Y({ S3934 })
);
NAND #() 
NAND_2631_ (
  .A({ S1304 }),
  .B({ S1745 }),
  .Y({ S3935 })
);
NOR #() 
NOR_1091_ (
  .A({ S3932 }),
  .B({ S3934 }),
  .Y({ S3936 })
);
NAND #() 
NAND_2632_ (
  .A({ S3933 }),
  .B({ S3935 }),
  .Y({ S3937 })
);
NOR #() 
NOR_1092_ (
  .A({ datapath_addsubunit_in1_14 }),
  .B({ S1516 }),
  .Y({ S3938 })
);
NOT #() 
NOT_323_ (
  .A({ S3938 }),
  .Y({ S3939 })
);
NOR #() 
NOR_1093_ (
  .A({ S3937 }),
  .B({ S3938 }),
  .Y({ S3940 })
);
NAND #() 
NAND_2633_ (
  .A({ S3936 }),
  .B({ S3939 }),
  .Y({ S3941 })
);
NOR #() 
NOR_1094_ (
  .A({ S3932 }),
  .B({ S3940 }),
  .Y({ S3942 })
);
NAND #() 
NAND_2634_ (
  .A({ S3933 }),
  .B({ S3941 }),
  .Y({ S3943 })
);
NOR #() 
NOR_1095_ (
  .A({ S3925 }),
  .B({ S3942 }),
  .Y({ S3944 })
);
NAND #() 
NAND_2635_ (
  .A({ S3924 }),
  .B({ S3943 }),
  .Y({ S3945 })
);
NAND #() 
NAND_2636_ (
  .A({ S3937 }),
  .B({ S3938 }),
  .Y({ S3946 })
);
NAND #() 
NAND_2637_ (
  .A({ S3941 }),
  .B({ S3946 }),
  .Y({ S3947 })
);
NAND #() 
NAND_2638_ (
  .A({ S3930 }),
  .B({ S3945 }),
  .Y({ S3948 })
);
NOT #() 
NOT_324_ (
  .A({ S3948 }),
  .Y({ S3949 })
);
NOR #() 
NOR_1096_ (
  .A({ S3945 }),
  .B({ S3947 }),
  .Y({ S3950 })
);
NOT #() 
NOT_325_ (
  .A({ S3950 }),
  .Y({ S3951 })
);
NAND #() 
NAND_2639_ (
  .A({ S3948 }),
  .B({ S3951 }),
  .Y({ S3952 })
);
NOR #() 
NOR_1097_ (
  .A({ S3949 }),
  .B({ S3950 }),
  .Y({ S3953 })
);
NOR #() 
NOR_1098_ (
  .A({ S1516 }),
  .B({ S3945 }),
  .Y({ S3954 })
);
NAND #() 
NAND_2640_ (
  .A({ S1515 }),
  .B({ S3944 }),
  .Y({ S3955 })
);
NOR #() 
NOR_1099_ (
  .A({ S492 }),
  .B({ S3954 }),
  .Y({ S3956 })
);
NAND #() 
NAND_2641_ (
  .A({ datapath_addsubunit_in1_14 }),
  .B({ S3955 }),
  .Y({ S3957 })
);
NOR #() 
NOR_1100_ (
  .A({ S1745 }),
  .B({ S3957 }),
  .Y({ S3958 })
);
NAND #() 
NAND_2642_ (
  .A({ S1746 }),
  .B({ S3956 }),
  .Y({ S3959 })
);
NOR #() 
NOR_1101_ (
  .A({ S1746 }),
  .B({ S3956 }),
  .Y({ S3960 })
);
NAND #() 
NAND_2643_ (
  .A({ S1745 }),
  .B({ S3957 }),
  .Y({ S3961 })
);
NOR #() 
NOR_1102_ (
  .A({ S3958 }),
  .B({ S3960 }),
  .Y({ S3962 })
);
NAND #() 
NAND_2644_ (
  .A({ S3959 }),
  .B({ S3961 }),
  .Y({ S3963 })
);
NOR #() 
NOR_1103_ (
  .A({ datapath_addsubunit_in1_13 }),
  .B({ S1516 }),
  .Y({ S3964 })
);
NAND #() 
NAND_2645_ (
  .A({ S548 }),
  .B({ S1515 }),
  .Y({ S3965 })
);
NOR #() 
NOR_1104_ (
  .A({ S3963 }),
  .B({ S3964 }),
  .Y({ S3966 })
);
NAND #() 
NAND_2646_ (
  .A({ S3962 }),
  .B({ S3965 }),
  .Y({ S3967 })
);
NOR #() 
NOR_1105_ (
  .A({ S3958 }),
  .B({ S3966 }),
  .Y({ S3968 })
);
NAND #() 
NAND_2647_ (
  .A({ S3959 }),
  .B({ S3967 }),
  .Y({ S3969 })
);
NOR #() 
NOR_1106_ (
  .A({ S1849 }),
  .B({ S3923 }),
  .Y({ S3970 })
);
NAND #() 
NAND_2648_ (
  .A({ S3969 }),
  .B({ S3970 }),
  .Y({ S3971 })
);
NOR #() 
NOR_1107_ (
  .A({ S3925 }),
  .B({ S3969 }),
  .Y({ S3972 })
);
NAND #() 
NAND_2649_ (
  .A({ S3952 }),
  .B({ S3971 }),
  .Y({ S3973 })
);
NOR #() 
NOR_1108_ (
  .A({ S3972 }),
  .B({ S3973 }),
  .Y({ S3974 })
);
NOT #() 
NOT_326_ (
  .A({ S3974 }),
  .Y({ S3975 })
);
NOR #() 
NOR_1109_ (
  .A({ S1848 }),
  .B({ S3953 }),
  .Y({ S3976 })
);
NAND #() 
NAND_2650_ (
  .A({ S1849 }),
  .B({ S3952 }),
  .Y({ S3977 })
);
NOR #() 
NOR_1110_ (
  .A({ S3969 }),
  .B({ S3976 }),
  .Y({ S3978 })
);
NAND #() 
NAND_2651_ (
  .A({ S3968 }),
  .B({ S3977 }),
  .Y({ S3979 })
);
NOR #() 
NOR_1111_ (
  .A({ datapath_addsubunit_in1_15 }),
  .B({ S1849 }),
  .Y({ S3980 })
);
NAND #() 
NAND_2652_ (
  .A({ S1304 }),
  .B({ S1848 }),
  .Y({ S3981 })
);
NOR #() 
NOR_1112_ (
  .A({ S3923 }),
  .B({ S3980 }),
  .Y({ S3982 })
);
NAND #() 
NAND_2653_ (
  .A({ S3922 }),
  .B({ S3981 }),
  .Y({ S3983 })
);
NOR #() 
NOR_1113_ (
  .A({ S3978 }),
  .B({ S3983 }),
  .Y({ S3984 })
);
NAND #() 
NAND_2654_ (
  .A({ S3979 }),
  .B({ S3982 }),
  .Y({ S3985 })
);
NOR #() 
NOR_1114_ (
  .A({ S3962 }),
  .B({ S3965 }),
  .Y({ S3986 })
);
NOR #() 
NOR_1115_ (
  .A({ S3966 }),
  .B({ S3986 }),
  .Y({ S3987 })
);
NOR #() 
NOR_1116_ (
  .A({ S3985 }),
  .B({ S3987 }),
  .Y({ S3988 })
);
NOT #() 
NOT_327_ (
  .A({ S3988 }),
  .Y({ S3989 })
);
NOR #() 
NOR_1117_ (
  .A({ S3956 }),
  .B({ S3984 }),
  .Y({ S3990 })
);
NAND #() 
NAND_2655_ (
  .A({ S3957 }),
  .B({ S3985 }),
  .Y({ S3991 })
);
NOR #() 
NOR_1118_ (
  .A({ S3988 }),
  .B({ S3990 }),
  .Y({ S3992 })
);
NAND #() 
NAND_2656_ (
  .A({ S3989 }),
  .B({ S3991 }),
  .Y({ S3993 })
);
NOR #() 
NOR_1119_ (
  .A({ S1848 }),
  .B({ S3993 }),
  .Y({ S3994 })
);
NAND #() 
NAND_2657_ (
  .A({ S1849 }),
  .B({ S3992 }),
  .Y({ S3995 })
);
NOR #() 
NOR_1120_ (
  .A({ S1849 }),
  .B({ S3992 }),
  .Y({ S3996 })
);
NAND #() 
NAND_2658_ (
  .A({ S1848 }),
  .B({ S3993 }),
  .Y({ S3997 })
);
NOR #() 
NOR_1121_ (
  .A({ S3994 }),
  .B({ S3996 }),
  .Y({ S3998 })
);
NAND #() 
NAND_2659_ (
  .A({ S3995 }),
  .B({ S3997 }),
  .Y({ S3999 })
);
NOR #() 
NOR_1122_ (
  .A({ S1516 }),
  .B({ S3985 }),
  .Y({ S4000 })
);
NAND #() 
NAND_2660_ (
  .A({ S1515 }),
  .B({ S3984 }),
  .Y({ S4001 })
);
NOR #() 
NOR_1123_ (
  .A({ datapath_addsubunit_in1_13 }),
  .B({ S4000 }),
  .Y({ S4002 })
);
NAND #() 
NAND_2661_ (
  .A({ S548 }),
  .B({ S4001 }),
  .Y({ S4003 })
);
NOR #() 
NOR_1124_ (
  .A({ S548 }),
  .B({ S4001 }),
  .Y({ S4004 })
);
NAND #() 
NAND_2662_ (
  .A({ datapath_addsubunit_in1_13 }),
  .B({ S4000 }),
  .Y({ S4005 })
);
NOR #() 
NOR_1125_ (
  .A({ S4002 }),
  .B({ S4004 }),
  .Y({ S4006 })
);
NAND #() 
NAND_2663_ (
  .A({ S4003 }),
  .B({ S4005 }),
  .Y({ S4007 })
);
NOR #() 
NOR_1126_ (
  .A({ S1745 }),
  .B({ S4007 }),
  .Y({ S4008 })
);
NAND #() 
NAND_2664_ (
  .A({ S1746 }),
  .B({ S4006 }),
  .Y({ S4009 })
);
NOR #() 
NOR_1127_ (
  .A({ datapath_addsubunit_in1_12 }),
  .B({ S1516 }),
  .Y({ S4010 })
);
NAND #() 
NAND_2665_ (
  .A({ S599 }),
  .B({ S1515 }),
  .Y({ S4011 })
);
NOR #() 
NOR_1128_ (
  .A({ S1746 }),
  .B({ S4006 }),
  .Y({ S4012 })
);
NAND #() 
NAND_2666_ (
  .A({ S1745 }),
  .B({ S4007 }),
  .Y({ S4013 })
);
NOR #() 
NOR_1129_ (
  .A({ S4008 }),
  .B({ S4012 }),
  .Y({ S4014 })
);
NAND #() 
NAND_2667_ (
  .A({ S4009 }),
  .B({ S4013 }),
  .Y({ S4015 })
);
NOR #() 
NOR_1130_ (
  .A({ S4010 }),
  .B({ S4015 }),
  .Y({ S4016 })
);
NAND #() 
NAND_2668_ (
  .A({ S4011 }),
  .B({ S4014 }),
  .Y({ S4017 })
);
NOR #() 
NOR_1131_ (
  .A({ S4008 }),
  .B({ S4016 }),
  .Y({ S4018 })
);
NAND #() 
NAND_2669_ (
  .A({ S4009 }),
  .B({ S4017 }),
  .Y({ S4019 })
);
NOR #() 
NOR_1132_ (
  .A({ S3999 }),
  .B({ S4018 }),
  .Y({ S4020 })
);
NAND #() 
NAND_2670_ (
  .A({ S3998 }),
  .B({ S4019 }),
  .Y({ S4021 })
);
NOR #() 
NOR_1133_ (
  .A({ S3994 }),
  .B({ S4020 }),
  .Y({ S4022 })
);
NAND #() 
NAND_2671_ (
  .A({ S3995 }),
  .B({ S4021 }),
  .Y({ S4023 })
);
NOR #() 
NOR_1134_ (
  .A({ S1952 }),
  .B({ S4022 }),
  .Y({ S4024 })
);
NAND #() 
NAND_2672_ (
  .A({ S1953 }),
  .B({ S4023 }),
  .Y({ S4025 })
);
NOR #() 
NOR_1135_ (
  .A({ S1953 }),
  .B({ S4023 }),
  .Y({ S4026 })
);
NAND #() 
NAND_2673_ (
  .A({ S1952 }),
  .B({ S4022 }),
  .Y({ S4027 })
);
NOR #() 
NOR_1136_ (
  .A({ S3921 }),
  .B({ S4026 }),
  .Y({ S4028 })
);
NAND #() 
NAND_2674_ (
  .A({ S3920 }),
  .B({ S4027 }),
  .Y({ S4029 })
);
NAND #() 
NAND_2675_ (
  .A({ S4025 }),
  .B({ S4028 }),
  .Y({ S4030 })
);
NAND #() 
NAND_2676_ (
  .A({ S3974 }),
  .B({ S4030 }),
  .Y({ S4031 })
);
NOR #() 
NOR_1137_ (
  .A({ S3974 }),
  .B({ S4024 }),
  .Y({ S4032 })
);
NAND #() 
NAND_2677_ (
  .A({ S3975 }),
  .B({ S4025 }),
  .Y({ S4033 })
);
NOR #() 
NOR_1138_ (
  .A({ S4029 }),
  .B({ S4032 }),
  .Y({ S4034 })
);
NAND #() 
NAND_2678_ (
  .A({ S4028 }),
  .B({ S4033 }),
  .Y({ S4035 })
);
NOR #() 
NOR_1139_ (
  .A({ S3998 }),
  .B({ S4019 }),
  .Y({ S4036 })
);
NOR #() 
NOR_1140_ (
  .A({ S4020 }),
  .B({ S4036 }),
  .Y({ S4037 })
);
NOR #() 
NOR_1141_ (
  .A({ S4035 }),
  .B({ S4037 }),
  .Y({ S4038 })
);
NOT #() 
NOT_328_ (
  .A({ S4038 }),
  .Y({ S4039 })
);
NOR #() 
NOR_1142_ (
  .A({ S3992 }),
  .B({ S4034 }),
  .Y({ S4040 })
);
NAND #() 
NAND_2679_ (
  .A({ S3993 }),
  .B({ S4035 }),
  .Y({ S4041 })
);
NOR #() 
NOR_1143_ (
  .A({ S4038 }),
  .B({ S4040 }),
  .Y({ S4042 })
);
NAND #() 
NAND_2680_ (
  .A({ S4039 }),
  .B({ S4041 }),
  .Y({ S4043 })
);
NOR #() 
NOR_1144_ (
  .A({ S1952 }),
  .B({ S4043 }),
  .Y({ S4044 })
);
NAND #() 
NAND_2681_ (
  .A({ S1953 }),
  .B({ S4042 }),
  .Y({ S4045 })
);
NOR #() 
NOR_1145_ (
  .A({ S1953 }),
  .B({ S4042 }),
  .Y({ S4046 })
);
NAND #() 
NAND_2682_ (
  .A({ S1952 }),
  .B({ S4043 }),
  .Y({ S4047 })
);
NOR #() 
NOR_1146_ (
  .A({ S4044 }),
  .B({ S4046 }),
  .Y({ S4048 })
);
NAND #() 
NAND_2683_ (
  .A({ S4045 }),
  .B({ S4047 }),
  .Y({ S4049 })
);
NOR #() 
NOR_1147_ (
  .A({ S4011 }),
  .B({ S4014 }),
  .Y({ S4050 })
);
NOR #() 
NOR_1148_ (
  .A({ S4016 }),
  .B({ S4050 }),
  .Y({ S4051 })
);
NOR #() 
NOR_1149_ (
  .A({ S4035 }),
  .B({ S4051 }),
  .Y({ S4052 })
);
NOT #() 
NOT_329_ (
  .A({ S4052 }),
  .Y({ S4053 })
);
NAND #() 
NAND_2684_ (
  .A({ S4007 }),
  .B({ S4035 }),
  .Y({ S4054 })
);
NOT #() 
NOT_330_ (
  .A({ S4054 }),
  .Y({ S4055 })
);
NOR #() 
NOR_1150_ (
  .A({ S4052 }),
  .B({ S4055 }),
  .Y({ S4056 })
);
NAND #() 
NAND_2685_ (
  .A({ S4053 }),
  .B({ S4054 }),
  .Y({ S4057 })
);
NOR #() 
NOR_1151_ (
  .A({ S1848 }),
  .B({ S4057 }),
  .Y({ S4058 })
);
NAND #() 
NAND_2686_ (
  .A({ S1849 }),
  .B({ S4056 }),
  .Y({ S4059 })
);
NOR #() 
NOR_1152_ (
  .A({ S1849 }),
  .B({ S4056 }),
  .Y({ S4060 })
);
NAND #() 
NAND_2687_ (
  .A({ S1848 }),
  .B({ S4057 }),
  .Y({ S4061 })
);
NOR #() 
NOR_1153_ (
  .A({ S4058 }),
  .B({ S4060 }),
  .Y({ S4062 })
);
NAND #() 
NAND_2688_ (
  .A({ S4059 }),
  .B({ S4061 }),
  .Y({ S4063 })
);
NOR #() 
NOR_1154_ (
  .A({ S1516 }),
  .B({ S4035 }),
  .Y({ S4064 })
);
NAND #() 
NAND_2689_ (
  .A({ S1515 }),
  .B({ S4034 }),
  .Y({ S4065 })
);
NOR #() 
NOR_1155_ (
  .A({ S599 }),
  .B({ S4064 }),
  .Y({ S4066 })
);
NAND #() 
NAND_2690_ (
  .A({ datapath_addsubunit_in1_12 }),
  .B({ S4065 }),
  .Y({ S4067 })
);
NOR #() 
NOR_1156_ (
  .A({ S4011 }),
  .B({ S4035 }),
  .Y({ S4068 })
);
NOT #() 
NOT_331_ (
  .A({ S4068 }),
  .Y({ S4069 })
);
NOR #() 
NOR_1157_ (
  .A({ S4066 }),
  .B({ S4068 }),
  .Y({ S4070 })
);
NAND #() 
NAND_2691_ (
  .A({ S4067 }),
  .B({ S4069 }),
  .Y({ S4071 })
);
NOR #() 
NOR_1158_ (
  .A({ S1745 }),
  .B({ S4070 }),
  .Y({ S4072 })
);
NAND #() 
NAND_2692_ (
  .A({ S1746 }),
  .B({ S4071 }),
  .Y({ S4073 })
);
NOR #() 
NOR_1159_ (
  .A({ S1746 }),
  .B({ S4071 }),
  .Y({ S4074 })
);
NAND #() 
NAND_2693_ (
  .A({ S1745 }),
  .B({ S4070 }),
  .Y({ S4075 })
);
NOR #() 
NOR_1160_ (
  .A({ S4072 }),
  .B({ S4074 }),
  .Y({ S4076 })
);
NAND #() 
NAND_2694_ (
  .A({ S4073 }),
  .B({ S4075 }),
  .Y({ S4077 })
);
NOR #() 
NOR_1161_ (
  .A({ datapath_addsubunit_in1_11 }),
  .B({ S1516 }),
  .Y({ S4078 })
);
NAND #() 
NAND_2695_ (
  .A({ S651 }),
  .B({ S1515 }),
  .Y({ S4079 })
);
NOR #() 
NOR_1162_ (
  .A({ S4077 }),
  .B({ S4078 }),
  .Y({ S4080 })
);
NAND #() 
NAND_2696_ (
  .A({ S4076 }),
  .B({ S4079 }),
  .Y({ S4081 })
);
NOR #() 
NOR_1163_ (
  .A({ S4072 }),
  .B({ S4080 }),
  .Y({ S4082 })
);
NAND #() 
NAND_2697_ (
  .A({ S4073 }),
  .B({ S4081 }),
  .Y({ S4083 })
);
NOR #() 
NOR_1164_ (
  .A({ S4063 }),
  .B({ S4082 }),
  .Y({ S4084 })
);
NAND #() 
NAND_2698_ (
  .A({ S4062 }),
  .B({ S4083 }),
  .Y({ S4085 })
);
NOR #() 
NOR_1165_ (
  .A({ S4058 }),
  .B({ S4084 }),
  .Y({ S4086 })
);
NAND #() 
NAND_2699_ (
  .A({ S4059 }),
  .B({ S4085 }),
  .Y({ S4087 })
);
NOR #() 
NOR_1166_ (
  .A({ S4049 }),
  .B({ S4086 }),
  .Y({ S4088 })
);
NAND #() 
NAND_2700_ (
  .A({ S4048 }),
  .B({ S4087 }),
  .Y({ S4089 })
);
NOR #() 
NOR_1167_ (
  .A({ S4044 }),
  .B({ S4088 }),
  .Y({ S4090 })
);
NAND #() 
NAND_2701_ (
  .A({ S4045 }),
  .B({ S4089 }),
  .Y({ S4091 })
);
NAND #() 
NAND_2702_ (
  .A({ S1597 }),
  .B({ S3918 }),
  .Y({ S4092 })
);
NAND #() 
NAND_2703_ (
  .A({ S3920 }),
  .B({ S4090 }),
  .Y({ S4093 })
);
NOR #() 
NOR_1168_ (
  .A({ S4090 }),
  .B({ S4092 }),
  .Y({ S4094 })
);
NOT #() 
NOT_332_ (
  .A({ S4094 }),
  .Y({ S4095 })
);
NOR #() 
NOR_1169_ (
  .A({ S4031 }),
  .B({ S4094 }),
  .Y({ S4096 })
);
NAND #() 
NAND_2704_ (
  .A({ S4093 }),
  .B({ S4095 }),
  .Y({ S4097 })
);
NOR #() 
NOR_1170_ (
  .A({ S4031 }),
  .B({ S4097 }),
  .Y({ S4098 })
);
NAND #() 
NAND_2705_ (
  .A({ S4093 }),
  .B({ S4096 }),
  .Y({ S4099 })
);
NOR #() 
NOR_1171_ (
  .A({ S1597 }),
  .B({ S4031 }),
  .Y({ S4100 })
);
NOT #() 
NOT_333_ (
  .A({ S4100 }),
  .Y({ S4101 })
);
NOR #() 
NOR_1172_ (
  .A({ S4091 }),
  .B({ S4100 }),
  .Y({ S4102 })
);
NAND #() 
NAND_2706_ (
  .A({ S4090 }),
  .B({ S4101 }),
  .Y({ S4103 })
);
NAND #() 
NAND_2707_ (
  .A({ S1597 }),
  .B({ S3975 }),
  .Y({ S4104 })
);
NAND #() 
NAND_2708_ (
  .A({ S3918 }),
  .B({ S4104 }),
  .Y({ S4105 })
);
NOT #() 
NOT_334_ (
  .A({ S4105 }),
  .Y({ S4106 })
);
NOR #() 
NOR_1173_ (
  .A({ S4102 }),
  .B({ S4105 }),
  .Y({ S4107 })
);
NAND #() 
NAND_2709_ (
  .A({ S4103 }),
  .B({ S4106 }),
  .Y({ S4108 })
);
NOR #() 
NOR_1174_ (
  .A({ S4048 }),
  .B({ S4087 }),
  .Y({ S4109 })
);
NOR #() 
NOR_1175_ (
  .A({ S4088 }),
  .B({ S4109 }),
  .Y({ S4110 })
);
NOR #() 
NOR_1176_ (
  .A({ S4108 }),
  .B({ S4110 }),
  .Y({ S4111 })
);
NOT #() 
NOT_335_ (
  .A({ S4111 }),
  .Y({ S4112 })
);
NOR #() 
NOR_1177_ (
  .A({ S4042 }),
  .B({ S4107 }),
  .Y({ S4113 })
);
NAND #() 
NAND_2710_ (
  .A({ S4043 }),
  .B({ S4108 }),
  .Y({ S4114 })
);
NOR #() 
NOR_1178_ (
  .A({ S4111 }),
  .B({ S4113 }),
  .Y({ S4115 })
);
NAND #() 
NAND_2711_ (
  .A({ S4112 }),
  .B({ S4114 }),
  .Y({ S4116 })
);
NOR #() 
NOR_1179_ (
  .A({ S1597 }),
  .B({ S4116 }),
  .Y({ S4117 })
);
NAND #() 
NAND_2712_ (
  .A({ S1598 }),
  .B({ S4115 }),
  .Y({ S4118 })
);
NOR #() 
NOR_1180_ (
  .A({ S1598 }),
  .B({ S4115 }),
  .Y({ S4119 })
);
NAND #() 
NAND_2713_ (
  .A({ S1597 }),
  .B({ S4116 }),
  .Y({ S4120 })
);
NOR #() 
NOR_1181_ (
  .A({ S4117 }),
  .B({ S4119 }),
  .Y({ S4121 })
);
NAND #() 
NAND_2714_ (
  .A({ S4118 }),
  .B({ S4120 }),
  .Y({ S4122 })
);
NOR #() 
NOR_1182_ (
  .A({ S4062 }),
  .B({ S4083 }),
  .Y({ S4123 })
);
NOR #() 
NOR_1183_ (
  .A({ S4084 }),
  .B({ S4123 }),
  .Y({ S4124 })
);
NOR #() 
NOR_1184_ (
  .A({ S4108 }),
  .B({ S4124 }),
  .Y({ S4125 })
);
NOT #() 
NOT_336_ (
  .A({ S4125 }),
  .Y({ S4126 })
);
NOR #() 
NOR_1185_ (
  .A({ S4056 }),
  .B({ S4107 }),
  .Y({ S4127 })
);
NAND #() 
NAND_2715_ (
  .A({ S4057 }),
  .B({ S4108 }),
  .Y({ S4128 })
);
NOR #() 
NOR_1186_ (
  .A({ S4125 }),
  .B({ S4127 }),
  .Y({ S4129 })
);
NAND #() 
NAND_2716_ (
  .A({ S4126 }),
  .B({ S4128 }),
  .Y({ S4130 })
);
NOR #() 
NOR_1187_ (
  .A({ S1952 }),
  .B({ S4130 }),
  .Y({ S4131 })
);
NAND #() 
NAND_2717_ (
  .A({ S1953 }),
  .B({ S4129 }),
  .Y({ S4132 })
);
NOR #() 
NOR_1188_ (
  .A({ S1953 }),
  .B({ S4129 }),
  .Y({ S4133 })
);
NAND #() 
NAND_2718_ (
  .A({ S1952 }),
  .B({ S4130 }),
  .Y({ S4134 })
);
NOR #() 
NOR_1189_ (
  .A({ S4131 }),
  .B({ S4133 }),
  .Y({ S4135 })
);
NAND #() 
NAND_2719_ (
  .A({ S4132 }),
  .B({ S4134 }),
  .Y({ S4136 })
);
NOR #() 
NOR_1190_ (
  .A({ S4076 }),
  .B({ S4079 }),
  .Y({ S4137 })
);
NOR #() 
NOR_1191_ (
  .A({ S4080 }),
  .B({ S4137 }),
  .Y({ S4138 })
);
NOR #() 
NOR_1192_ (
  .A({ S4108 }),
  .B({ S4138 }),
  .Y({ S4139 })
);
NOT #() 
NOT_337_ (
  .A({ S4139 }),
  .Y({ S4140 })
);
NAND #() 
NAND_2720_ (
  .A({ S4070 }),
  .B({ S4108 }),
  .Y({ S4141 })
);
NOT #() 
NOT_338_ (
  .A({ S4141 }),
  .Y({ S4142 })
);
NOR #() 
NOR_1193_ (
  .A({ S4139 }),
  .B({ S4142 }),
  .Y({ S4143 })
);
NAND #() 
NAND_2721_ (
  .A({ S4140 }),
  .B({ S4141 }),
  .Y({ S4144 })
);
NOR #() 
NOR_1194_ (
  .A({ S1848 }),
  .B({ S4144 }),
  .Y({ S4145 })
);
NAND #() 
NAND_2722_ (
  .A({ S1849 }),
  .B({ S4143 }),
  .Y({ S4146 })
);
NOR #() 
NOR_1195_ (
  .A({ S1849 }),
  .B({ S4143 }),
  .Y({ S4147 })
);
NAND #() 
NAND_2723_ (
  .A({ S1848 }),
  .B({ S4144 }),
  .Y({ S4148 })
);
NOR #() 
NOR_1196_ (
  .A({ S4145 }),
  .B({ S4147 }),
  .Y({ S4149 })
);
NAND #() 
NAND_2724_ (
  .A({ S4146 }),
  .B({ S4148 }),
  .Y({ S4150 })
);
NOR #() 
NOR_1197_ (
  .A({ S1516 }),
  .B({ S4108 }),
  .Y({ S4151 })
);
NAND #() 
NAND_2725_ (
  .A({ S1515 }),
  .B({ S4107 }),
  .Y({ S4152 })
);
NOR #() 
NOR_1198_ (
  .A({ S651 }),
  .B({ S4152 }),
  .Y({ S4153 })
);
NAND #() 
NAND_2726_ (
  .A({ datapath_addsubunit_in1_11 }),
  .B({ S4151 }),
  .Y({ S4154 })
);
NOR #() 
NOR_1199_ (
  .A({ datapath_addsubunit_in1_11 }),
  .B({ S4151 }),
  .Y({ S4155 })
);
NAND #() 
NAND_2727_ (
  .A({ S651 }),
  .B({ S4152 }),
  .Y({ S4156 })
);
NAND #() 
NAND_2728_ (
  .A({ S4154 }),
  .B({ S4156 }),
  .Y({ S4157 })
);
NOR #() 
NOR_1200_ (
  .A({ S4153 }),
  .B({ S4155 }),
  .Y({ S4158 })
);
NOR #() 
NOR_1201_ (
  .A({ S1745 }),
  .B({ S4157 }),
  .Y({ S4159 })
);
NAND #() 
NAND_2729_ (
  .A({ S1746 }),
  .B({ S4158 }),
  .Y({ S4160 })
);
NOR #() 
NOR_1202_ (
  .A({ datapath_addsubunit_in1_10 }),
  .B({ S1516 }),
  .Y({ S4161 })
);
NAND #() 
NAND_2730_ (
  .A({ S702 }),
  .B({ S1515 }),
  .Y({ S4162 })
);
NOR #() 
NOR_1203_ (
  .A({ S1746 }),
  .B({ S4158 }),
  .Y({ S4163 })
);
NAND #() 
NAND_2731_ (
  .A({ S1745 }),
  .B({ S4157 }),
  .Y({ S4164 })
);
NOR #() 
NOR_1204_ (
  .A({ S4159 }),
  .B({ S4163 }),
  .Y({ S4165 })
);
NAND #() 
NAND_2732_ (
  .A({ S4160 }),
  .B({ S4164 }),
  .Y({ S4166 })
);
NOR #() 
NOR_1205_ (
  .A({ S4161 }),
  .B({ S4166 }),
  .Y({ S4167 })
);
NAND #() 
NAND_2733_ (
  .A({ S4162 }),
  .B({ S4165 }),
  .Y({ S4168 })
);
NOR #() 
NOR_1206_ (
  .A({ S4159 }),
  .B({ S4167 }),
  .Y({ S4169 })
);
NAND #() 
NAND_2734_ (
  .A({ S4160 }),
  .B({ S4168 }),
  .Y({ S4170 })
);
NOR #() 
NOR_1207_ (
  .A({ S4150 }),
  .B({ S4169 }),
  .Y({ S4171 })
);
NAND #() 
NAND_2735_ (
  .A({ S4149 }),
  .B({ S4170 }),
  .Y({ S4172 })
);
NOR #() 
NOR_1208_ (
  .A({ S4145 }),
  .B({ S4171 }),
  .Y({ S4173 })
);
NAND #() 
NAND_2736_ (
  .A({ S4146 }),
  .B({ S4172 }),
  .Y({ S4174 })
);
NOR #() 
NOR_1209_ (
  .A({ S4136 }),
  .B({ S4173 }),
  .Y({ S4175 })
);
NAND #() 
NAND_2737_ (
  .A({ S4135 }),
  .B({ S4174 }),
  .Y({ S4176 })
);
NOR #() 
NOR_1210_ (
  .A({ S4131 }),
  .B({ S4175 }),
  .Y({ S4177 })
);
NAND #() 
NAND_2738_ (
  .A({ S4132 }),
  .B({ S4176 }),
  .Y({ S4178 })
);
NOR #() 
NOR_1211_ (
  .A({ S4122 }),
  .B({ S4177 }),
  .Y({ S4179 })
);
NAND #() 
NAND_2739_ (
  .A({ S4121 }),
  .B({ S4178 }),
  .Y({ S4180 })
);
NOR #() 
NOR_1212_ (
  .A({ S4117 }),
  .B({ S4179 }),
  .Y({ S4181 })
);
NAND #() 
NAND_2740_ (
  .A({ S4118 }),
  .B({ S4180 }),
  .Y({ S4182 })
);
NOR #() 
NOR_1213_ (
  .A({ S2106 }),
  .B({ S4181 }),
  .Y({ S4183 })
);
NAND #() 
NAND_2741_ (
  .A({ S2107 }),
  .B({ S4182 }),
  .Y({ S4184 })
);
NOR #() 
NOR_1214_ (
  .A({ S2107 }),
  .B({ S4182 }),
  .Y({ S4185 })
);
NAND #() 
NAND_2742_ (
  .A({ S2106 }),
  .B({ S4181 }),
  .Y({ S4186 })
);
NOR #() 
NOR_1215_ (
  .A({ S3917 }),
  .B({ S4185 }),
  .Y({ S4187 })
);
NAND #() 
NAND_2743_ (
  .A({ S3916 }),
  .B({ S4186 }),
  .Y({ S4188 })
);
NOR #() 
NOR_1216_ (
  .A({ S4183 }),
  .B({ S4188 }),
  .Y({ S4189 })
);
NOR #() 
NOR_1217_ (
  .A({ S4099 }),
  .B({ S4189 }),
  .Y({ S4190 })
);
NOT #() 
NOT_339_ (
  .A({ S4190 }),
  .Y({ S4191 })
);
NOR #() 
NOR_1218_ (
  .A({ S4098 }),
  .B({ S4183 }),
  .Y({ S4192 })
);
NAND #() 
NAND_2744_ (
  .A({ S4099 }),
  .B({ S4184 }),
  .Y({ S4193 })
);
NOR #() 
NOR_1219_ (
  .A({ S4188 }),
  .B({ S4192 }),
  .Y({ S4194 })
);
NAND #() 
NAND_2745_ (
  .A({ S4187 }),
  .B({ S4193 }),
  .Y({ S4195 })
);
NOR #() 
NOR_1220_ (
  .A({ S4121 }),
  .B({ S4178 }),
  .Y({ S4196 })
);
NAND #() 
NAND_2746_ (
  .A({ S4122 }),
  .B({ S4177 }),
  .Y({ S4197 })
);
NOR #() 
NOR_1221_ (
  .A({ S4179 }),
  .B({ S4196 }),
  .Y({ S4198 })
);
NAND #() 
NAND_2747_ (
  .A({ S4180 }),
  .B({ S4197 }),
  .Y({ S4199 })
);
NOR #() 
NOR_1222_ (
  .A({ S4195 }),
  .B({ S4198 }),
  .Y({ S4200 })
);
NAND #() 
NAND_2748_ (
  .A({ S4194 }),
  .B({ S4199 }),
  .Y({ S4201 })
);
NOR #() 
NOR_1223_ (
  .A({ S4115 }),
  .B({ S4194 }),
  .Y({ S4202 })
);
NAND #() 
NAND_2749_ (
  .A({ S4116 }),
  .B({ S4195 }),
  .Y({ S4203 })
);
NOR #() 
NOR_1224_ (
  .A({ S4200 }),
  .B({ S4202 }),
  .Y({ S4204 })
);
NAND #() 
NAND_2750_ (
  .A({ S4201 }),
  .B({ S4203 }),
  .Y({ S4205 })
);
NOR #() 
NOR_1225_ (
  .A({ S2106 }),
  .B({ S4205 }),
  .Y({ S4206 })
);
NAND #() 
NAND_2751_ (
  .A({ S2107 }),
  .B({ S4204 }),
  .Y({ S4207 })
);
NOR #() 
NOR_1226_ (
  .A({ S2107 }),
  .B({ S4204 }),
  .Y({ S4208 })
);
NAND #() 
NAND_2752_ (
  .A({ S2106 }),
  .B({ S4205 }),
  .Y({ S4209 })
);
NOR #() 
NOR_1227_ (
  .A({ S4206 }),
  .B({ S4208 }),
  .Y({ S4210 })
);
NAND #() 
NAND_2753_ (
  .A({ S4207 }),
  .B({ S4209 }),
  .Y({ S4211 })
);
NOR #() 
NOR_1228_ (
  .A({ S4135 }),
  .B({ S4174 }),
  .Y({ S4212 })
);
NAND #() 
NAND_2754_ (
  .A({ S4136 }),
  .B({ S4173 }),
  .Y({ S4213 })
);
NOR #() 
NOR_1229_ (
  .A({ S4175 }),
  .B({ S4212 }),
  .Y({ S4214 })
);
NAND #() 
NAND_2755_ (
  .A({ S4176 }),
  .B({ S4213 }),
  .Y({ S4215 })
);
NOR #() 
NOR_1230_ (
  .A({ S4195 }),
  .B({ S4214 }),
  .Y({ S4216 })
);
NAND #() 
NAND_2756_ (
  .A({ S4194 }),
  .B({ S4215 }),
  .Y({ S4217 })
);
NOR #() 
NOR_1231_ (
  .A({ S4129 }),
  .B({ S4194 }),
  .Y({ S4218 })
);
NAND #() 
NAND_2757_ (
  .A({ S4130 }),
  .B({ S4195 }),
  .Y({ S4219 })
);
NOR #() 
NOR_1232_ (
  .A({ S4216 }),
  .B({ S4218 }),
  .Y({ S4220 })
);
NAND #() 
NAND_2758_ (
  .A({ S4217 }),
  .B({ S4219 }),
  .Y({ S4221 })
);
NOR #() 
NOR_1233_ (
  .A({ S1597 }),
  .B({ S4221 }),
  .Y({ S4222 })
);
NAND #() 
NAND_2759_ (
  .A({ S1598 }),
  .B({ S4220 }),
  .Y({ S4223 })
);
NOR #() 
NOR_1234_ (
  .A({ S1598 }),
  .B({ S4220 }),
  .Y({ S4224 })
);
NAND #() 
NAND_2760_ (
  .A({ S1597 }),
  .B({ S4221 }),
  .Y({ S4225 })
);
NOR #() 
NOR_1235_ (
  .A({ S4222 }),
  .B({ S4224 }),
  .Y({ S4226 })
);
NAND #() 
NAND_2761_ (
  .A({ S4223 }),
  .B({ S4225 }),
  .Y({ S4227 })
);
NOR #() 
NOR_1236_ (
  .A({ S4149 }),
  .B({ S4170 }),
  .Y({ S4228 })
);
NAND #() 
NAND_2762_ (
  .A({ S4150 }),
  .B({ S4169 }),
  .Y({ S4229 })
);
NOR #() 
NOR_1237_ (
  .A({ S4171 }),
  .B({ S4228 }),
  .Y({ S4230 })
);
NAND #() 
NAND_2763_ (
  .A({ S4172 }),
  .B({ S4229 }),
  .Y({ S4231 })
);
NOR #() 
NOR_1238_ (
  .A({ S4195 }),
  .B({ S4230 }),
  .Y({ S4232 })
);
NAND #() 
NAND_2764_ (
  .A({ S4194 }),
  .B({ S4231 }),
  .Y({ S4233 })
);
NOR #() 
NOR_1239_ (
  .A({ S4143 }),
  .B({ S4194 }),
  .Y({ S4234 })
);
NAND #() 
NAND_2765_ (
  .A({ S4144 }),
  .B({ S4195 }),
  .Y({ S4235 })
);
NOR #() 
NOR_1240_ (
  .A({ S4232 }),
  .B({ S4234 }),
  .Y({ S4236 })
);
NAND #() 
NAND_2766_ (
  .A({ S4233 }),
  .B({ S4235 }),
  .Y({ S4237 })
);
NOR #() 
NOR_1241_ (
  .A({ S1952 }),
  .B({ S4237 }),
  .Y({ S4238 })
);
NAND #() 
NAND_2767_ (
  .A({ S1953 }),
  .B({ S4236 }),
  .Y({ S4239 })
);
NOR #() 
NOR_1242_ (
  .A({ S1953 }),
  .B({ S4236 }),
  .Y({ S4240 })
);
NAND #() 
NAND_2768_ (
  .A({ S1952 }),
  .B({ S4237 }),
  .Y({ S4241 })
);
NOR #() 
NOR_1243_ (
  .A({ S4238 }),
  .B({ S4240 }),
  .Y({ S4242 })
);
NAND #() 
NAND_2769_ (
  .A({ S4239 }),
  .B({ S4241 }),
  .Y({ S4243 })
);
NOR #() 
NOR_1244_ (
  .A({ S4158 }),
  .B({ S4194 }),
  .Y({ S4244 })
);
NAND #() 
NAND_2770_ (
  .A({ S4157 }),
  .B({ S4195 }),
  .Y({ S4245 })
);
NOR #() 
NOR_1245_ (
  .A({ S4162 }),
  .B({ S4165 }),
  .Y({ S4246 })
);
NAND #() 
NAND_2771_ (
  .A({ S4161 }),
  .B({ S4166 }),
  .Y({ S4247 })
);
NOR #() 
NOR_1246_ (
  .A({ S4167 }),
  .B({ S4246 }),
  .Y({ S4248 })
);
NAND #() 
NAND_2772_ (
  .A({ S4168 }),
  .B({ S4247 }),
  .Y({ S4249 })
);
NOR #() 
NOR_1247_ (
  .A({ S4195 }),
  .B({ S4248 }),
  .Y({ S4250 })
);
NAND #() 
NAND_2773_ (
  .A({ S4194 }),
  .B({ S4249 }),
  .Y({ S4251 })
);
NOR #() 
NOR_1248_ (
  .A({ S4244 }),
  .B({ S4250 }),
  .Y({ S4252 })
);
NAND #() 
NAND_2774_ (
  .A({ S4245 }),
  .B({ S4251 }),
  .Y({ S4253 })
);
NOR #() 
NOR_1249_ (
  .A({ S1848 }),
  .B({ S4253 }),
  .Y({ S4254 })
);
NAND #() 
NAND_2775_ (
  .A({ S1849 }),
  .B({ S4252 }),
  .Y({ S4255 })
);
NOR #() 
NOR_1250_ (
  .A({ S1849 }),
  .B({ S4252 }),
  .Y({ S4256 })
);
NAND #() 
NAND_2776_ (
  .A({ S1848 }),
  .B({ S4253 }),
  .Y({ S4257 })
);
NOR #() 
NOR_1251_ (
  .A({ S4254 }),
  .B({ S4256 }),
  .Y({ S4258 })
);
NAND #() 
NAND_2777_ (
  .A({ S4255 }),
  .B({ S4257 }),
  .Y({ S4259 })
);
NOR #() 
NOR_1252_ (
  .A({ S1516 }),
  .B({ S4195 }),
  .Y({ S4260 })
);
NAND #() 
NAND_2778_ (
  .A({ S1515 }),
  .B({ S4194 }),
  .Y({ S4261 })
);
NOR #() 
NOR_1253_ (
  .A({ S702 }),
  .B({ S4261 }),
  .Y({ S4262 })
);
NAND #() 
NAND_2779_ (
  .A({ datapath_addsubunit_in1_10 }),
  .B({ S4260 }),
  .Y({ S4263 })
);
NOR #() 
NOR_1254_ (
  .A({ datapath_addsubunit_in1_10 }),
  .B({ S4260 }),
  .Y({ S4264 })
);
NAND #() 
NAND_2780_ (
  .A({ S702 }),
  .B({ S4261 }),
  .Y({ S4265 })
);
NOR #() 
NOR_1255_ (
  .A({ S4262 }),
  .B({ S4264 }),
  .Y({ S4266 })
);
NAND #() 
NAND_2781_ (
  .A({ S4263 }),
  .B({ S4265 }),
  .Y({ S4267 })
);
NOR #() 
NOR_1256_ (
  .A({ S1745 }),
  .B({ S4267 }),
  .Y({ S4268 })
);
NAND #() 
NAND_2782_ (
  .A({ S1746 }),
  .B({ S4266 }),
  .Y({ S4269 })
);
NOR #() 
NOR_1257_ (
  .A({ S1746 }),
  .B({ S4266 }),
  .Y({ S4270 })
);
NAND #() 
NAND_2783_ (
  .A({ S1745 }),
  .B({ S4267 }),
  .Y({ S4271 })
);
NOR #() 
NOR_1258_ (
  .A({ S4268 }),
  .B({ S4270 }),
  .Y({ S4272 })
);
NAND #() 
NAND_2784_ (
  .A({ S4269 }),
  .B({ S4271 }),
  .Y({ S4273 })
);
NOR #() 
NOR_1259_ (
  .A({ datapath_addsubunit_in1_9 }),
  .B({ S1516 }),
  .Y({ S4274 })
);
NAND #() 
NAND_2785_ (
  .A({ S754 }),
  .B({ S1515 }),
  .Y({ S4275 })
);
NOR #() 
NOR_1260_ (
  .A({ S4273 }),
  .B({ S4274 }),
  .Y({ S4276 })
);
NAND #() 
NAND_2786_ (
  .A({ S4272 }),
  .B({ S4275 }),
  .Y({ S4277 })
);
NOR #() 
NOR_1261_ (
  .A({ S4268 }),
  .B({ S4276 }),
  .Y({ S4278 })
);
NAND #() 
NAND_2787_ (
  .A({ S4269 }),
  .B({ S4277 }),
  .Y({ S4279 })
);
NOR #() 
NOR_1262_ (
  .A({ S4259 }),
  .B({ S4278 }),
  .Y({ S4280 })
);
NAND #() 
NAND_2788_ (
  .A({ S4258 }),
  .B({ S4279 }),
  .Y({ S4281 })
);
NOR #() 
NOR_1263_ (
  .A({ S4254 }),
  .B({ S4280 }),
  .Y({ S4282 })
);
NAND #() 
NAND_2789_ (
  .A({ S4255 }),
  .B({ S4281 }),
  .Y({ S4283 })
);
NOR #() 
NOR_1264_ (
  .A({ S4243 }),
  .B({ S4282 }),
  .Y({ S4284 })
);
NAND #() 
NAND_2790_ (
  .A({ S4242 }),
  .B({ S4283 }),
  .Y({ S4285 })
);
NOR #() 
NOR_1265_ (
  .A({ S4238 }),
  .B({ S4284 }),
  .Y({ S4286 })
);
NAND #() 
NAND_2791_ (
  .A({ S4239 }),
  .B({ S4285 }),
  .Y({ S4287 })
);
NOR #() 
NOR_1266_ (
  .A({ S4227 }),
  .B({ S4286 }),
  .Y({ S4288 })
);
NAND #() 
NAND_2792_ (
  .A({ S4226 }),
  .B({ S4287 }),
  .Y({ S4289 })
);
NOR #() 
NOR_1267_ (
  .A({ S4222 }),
  .B({ S4288 }),
  .Y({ S4290 })
);
NAND #() 
NAND_2793_ (
  .A({ S4223 }),
  .B({ S4289 }),
  .Y({ S4291 })
);
NOR #() 
NOR_1268_ (
  .A({ S4211 }),
  .B({ S4290 }),
  .Y({ S4292 })
);
NAND #() 
NAND_2794_ (
  .A({ S4210 }),
  .B({ S4291 }),
  .Y({ S4293 })
);
NOR #() 
NOR_1269_ (
  .A({ S4206 }),
  .B({ S4292 }),
  .Y({ S4294 })
);
NAND #() 
NAND_2795_ (
  .A({ S4207 }),
  .B({ S4293 }),
  .Y({ S4295 })
);
NAND #() 
NAND_2796_ (
  .A({ S2206 }),
  .B({ S4295 }),
  .Y({ S4296 })
);
NAND #() 
NAND_2797_ (
  .A({ S3914 }),
  .B({ S4295 }),
  .Y({ S4297 })
);
NAND #() 
NAND_2798_ (
  .A({ S3917 }),
  .B({ S4297 }),
  .Y({ S4298 })
);
NAND #() 
NAND_2799_ (
  .A({ S4296 }),
  .B({ S4298 }),
  .Y({ S4299 })
);
NAND #() 
NAND_2800_ (
  .A({ S4190 }),
  .B({ S4299 }),
  .Y({ S4300 })
);
NOT #() 
NOT_340_ (
  .A({ S4300 }),
  .Y({ S4301 })
);
NOR #() 
NOR_1270_ (
  .A({ S2311 }),
  .B({ S4300 }),
  .Y({ S4302 })
);
NAND #() 
NAND_2801_ (
  .A({ S2312 }),
  .B({ S4301 }),
  .Y({ S4303 })
);
NOR #() 
NOR_1271_ (
  .A({ S2312 }),
  .B({ S4190 }),
  .Y({ S4304 })
);
NOR #() 
NOR_1272_ (
  .A({ S4302 }),
  .B({ S4304 }),
  .Y({ S4305 })
);
NOT #() 
NOT_341_ (
  .A({ S4305 }),
  .Y({ S4306 })
);
NOR #() 
NOR_1273_ (
  .A({ S3917 }),
  .B({ S4191 }),
  .Y({ S4307 })
);
NAND #() 
NAND_2802_ (
  .A({ S3916 }),
  .B({ S4190 }),
  .Y({ S4308 })
);
NOR #() 
NOR_1274_ (
  .A({ S2206 }),
  .B({ S4098 }),
  .Y({ S4309 })
);
NOR #() 
NOR_1275_ (
  .A({ S4294 }),
  .B({ S4309 }),
  .Y({ S4310 })
);
NOR #() 
NOR_1276_ (
  .A({ S4297 }),
  .B({ S4309 }),
  .Y({ S4311 })
);
NAND #() 
NAND_2803_ (
  .A({ S3914 }),
  .B({ S4310 }),
  .Y({ S4312 })
);
NOR #() 
NOR_1277_ (
  .A({ S4307 }),
  .B({ S4311 }),
  .Y({ S4313 })
);
NAND #() 
NAND_2804_ (
  .A({ S4308 }),
  .B({ S4312 }),
  .Y({ S4314 })
);
NOR #() 
NOR_1278_ (
  .A({ S4210 }),
  .B({ S4291 }),
  .Y({ S4315 })
);
NOR #() 
NOR_1279_ (
  .A({ S4292 }),
  .B({ S4315 }),
  .Y({ S4316 })
);
NOR #() 
NOR_1280_ (
  .A({ S4313 }),
  .B({ S4316 }),
  .Y({ S4317 })
);
NOT #() 
NOT_342_ (
  .A({ S4317 }),
  .Y({ S4318 })
);
NOR #() 
NOR_1281_ (
  .A({ S4204 }),
  .B({ S4314 }),
  .Y({ S4319 })
);
NAND #() 
NAND_2805_ (
  .A({ S4205 }),
  .B({ S4313 }),
  .Y({ S4320 })
);
NOR #() 
NOR_1282_ (
  .A({ S4317 }),
  .B({ S4319 }),
  .Y({ S4321 })
);
NAND #() 
NAND_2806_ (
  .A({ S4318 }),
  .B({ S4320 }),
  .Y({ S4322 })
);
NOR #() 
NOR_1283_ (
  .A({ S2205 }),
  .B({ S4322 }),
  .Y({ S4323 })
);
NAND #() 
NAND_2807_ (
  .A({ S2206 }),
  .B({ S4321 }),
  .Y({ S4324 })
);
NOR #() 
NOR_1284_ (
  .A({ S2206 }),
  .B({ S4321 }),
  .Y({ S4325 })
);
NAND #() 
NAND_2808_ (
  .A({ S2205 }),
  .B({ S4322 }),
  .Y({ S4326 })
);
NOR #() 
NOR_1285_ (
  .A({ S4323 }),
  .B({ S4325 }),
  .Y({ S4327 })
);
NAND #() 
NAND_2809_ (
  .A({ S4324 }),
  .B({ S4326 }),
  .Y({ S4328 })
);
NOR #() 
NOR_1286_ (
  .A({ S4226 }),
  .B({ S4287 }),
  .Y({ S4329 })
);
NOR #() 
NOR_1287_ (
  .A({ S4288 }),
  .B({ S4329 }),
  .Y({ S4330 })
);
NOR #() 
NOR_1288_ (
  .A({ S4313 }),
  .B({ S4330 }),
  .Y({ S4331 })
);
NOT #() 
NOT_343_ (
  .A({ S4331 }),
  .Y({ S4332 })
);
NOR #() 
NOR_1289_ (
  .A({ S4220 }),
  .B({ S4314 }),
  .Y({ S4333 })
);
NAND #() 
NAND_2810_ (
  .A({ S4221 }),
  .B({ S4313 }),
  .Y({ S4334 })
);
NOR #() 
NOR_1290_ (
  .A({ S4331 }),
  .B({ S4333 }),
  .Y({ S4335 })
);
NAND #() 
NAND_2811_ (
  .A({ S4332 }),
  .B({ S4334 }),
  .Y({ S4336 })
);
NOR #() 
NOR_1291_ (
  .A({ S2106 }),
  .B({ S4336 }),
  .Y({ S4337 })
);
NAND #() 
NAND_2812_ (
  .A({ S2107 }),
  .B({ S4335 }),
  .Y({ S4338 })
);
NOR #() 
NOR_1292_ (
  .A({ S2107 }),
  .B({ S4335 }),
  .Y({ S4339 })
);
NAND #() 
NAND_2813_ (
  .A({ S2106 }),
  .B({ S4336 }),
  .Y({ S4340 })
);
NOR #() 
NOR_1293_ (
  .A({ S4337 }),
  .B({ S4339 }),
  .Y({ S4341 })
);
NAND #() 
NAND_2814_ (
  .A({ S4338 }),
  .B({ S4340 }),
  .Y({ S4342 })
);
NOR #() 
NOR_1294_ (
  .A({ S4242 }),
  .B({ S4283 }),
  .Y({ S4343 })
);
NOR #() 
NOR_1295_ (
  .A({ S4284 }),
  .B({ S4343 }),
  .Y({ S4344 })
);
NOR #() 
NOR_1296_ (
  .A({ S4313 }),
  .B({ S4344 }),
  .Y({ S4345 })
);
NOT #() 
NOT_344_ (
  .A({ S4345 }),
  .Y({ S4346 })
);
NOR #() 
NOR_1297_ (
  .A({ S4236 }),
  .B({ S4314 }),
  .Y({ S4347 })
);
NAND #() 
NAND_2815_ (
  .A({ S4237 }),
  .B({ S4313 }),
  .Y({ S4348 })
);
NOR #() 
NOR_1298_ (
  .A({ S4345 }),
  .B({ S4347 }),
  .Y({ S4349 })
);
NAND #() 
NAND_2816_ (
  .A({ S4346 }),
  .B({ S4348 }),
  .Y({ S4350 })
);
NOR #() 
NOR_1299_ (
  .A({ S1597 }),
  .B({ S4350 }),
  .Y({ S4351 })
);
NAND #() 
NAND_2817_ (
  .A({ S1598 }),
  .B({ S4349 }),
  .Y({ S4352 })
);
NOR #() 
NOR_1300_ (
  .A({ S1598 }),
  .B({ S4349 }),
  .Y({ S4353 })
);
NAND #() 
NAND_2818_ (
  .A({ S1597 }),
  .B({ S4350 }),
  .Y({ S4354 })
);
NOR #() 
NOR_1301_ (
  .A({ S4351 }),
  .B({ S4353 }),
  .Y({ S4355 })
);
NAND #() 
NAND_2819_ (
  .A({ S4352 }),
  .B({ S4354 }),
  .Y({ S4356 })
);
NOR #() 
NOR_1302_ (
  .A({ S4258 }),
  .B({ S4279 }),
  .Y({ S4357 })
);
NOR #() 
NOR_1303_ (
  .A({ S4280 }),
  .B({ S4357 }),
  .Y({ S4358 })
);
NOR #() 
NOR_1304_ (
  .A({ S4313 }),
  .B({ S4358 }),
  .Y({ S4359 })
);
NOT #() 
NOT_345_ (
  .A({ S4359 }),
  .Y({ S4360 })
);
NAND #() 
NAND_2820_ (
  .A({ S4253 }),
  .B({ S4313 }),
  .Y({ S4361 })
);
NOT #() 
NOT_346_ (
  .A({ S4361 }),
  .Y({ S4362 })
);
NOR #() 
NOR_1305_ (
  .A({ S4359 }),
  .B({ S4362 }),
  .Y({ S4363 })
);
NAND #() 
NAND_2821_ (
  .A({ S4360 }),
  .B({ S4361 }),
  .Y({ S4364 })
);
NOR #() 
NOR_1306_ (
  .A({ S1952 }),
  .B({ S4364 }),
  .Y({ S4365 })
);
NAND #() 
NAND_2822_ (
  .A({ S1953 }),
  .B({ S4363 }),
  .Y({ S4366 })
);
NOR #() 
NOR_1307_ (
  .A({ S1953 }),
  .B({ S4363 }),
  .Y({ S4367 })
);
NAND #() 
NAND_2823_ (
  .A({ S1952 }),
  .B({ S4364 }),
  .Y({ S4368 })
);
NOR #() 
NOR_1308_ (
  .A({ S4365 }),
  .B({ S4367 }),
  .Y({ S4369 })
);
NAND #() 
NAND_2824_ (
  .A({ S4366 }),
  .B({ S4368 }),
  .Y({ S4370 })
);
NOR #() 
NOR_1309_ (
  .A({ S4272 }),
  .B({ S4275 }),
  .Y({ S4371 })
);
NOR #() 
NOR_1310_ (
  .A({ S4276 }),
  .B({ S4371 }),
  .Y({ S4372 })
);
NOR #() 
NOR_1311_ (
  .A({ S4313 }),
  .B({ S4372 }),
  .Y({ S4373 })
);
NOT #() 
NOT_347_ (
  .A({ S4373 }),
  .Y({ S4374 })
);
NOR #() 
NOR_1312_ (
  .A({ S4266 }),
  .B({ S4314 }),
  .Y({ S4375 })
);
NAND #() 
NAND_2825_ (
  .A({ S4267 }),
  .B({ S4313 }),
  .Y({ S4376 })
);
NOR #() 
NOR_1313_ (
  .A({ S4373 }),
  .B({ S4375 }),
  .Y({ S4377 })
);
NAND #() 
NAND_2826_ (
  .A({ S4374 }),
  .B({ S4376 }),
  .Y({ S4378 })
);
NOR #() 
NOR_1314_ (
  .A({ S1848 }),
  .B({ S4378 }),
  .Y({ S4379 })
);
NAND #() 
NAND_2827_ (
  .A({ S1849 }),
  .B({ S4377 }),
  .Y({ S4380 })
);
NOR #() 
NOR_1315_ (
  .A({ S1849 }),
  .B({ S4377 }),
  .Y({ S4381 })
);
NAND #() 
NAND_2828_ (
  .A({ S1848 }),
  .B({ S4378 }),
  .Y({ S4382 })
);
NOR #() 
NOR_1316_ (
  .A({ S4379 }),
  .B({ S4381 }),
  .Y({ S4383 })
);
NAND #() 
NAND_2829_ (
  .A({ S4380 }),
  .B({ S4382 }),
  .Y({ S4384 })
);
NOR #() 
NOR_1317_ (
  .A({ S1516 }),
  .B({ S4313 }),
  .Y({ S4385 })
);
NAND #() 
NAND_2830_ (
  .A({ S1515 }),
  .B({ S4314 }),
  .Y({ S4386 })
);
NOR #() 
NOR_1318_ (
  .A({ S754 }),
  .B({ S4386 }),
  .Y({ S4387 })
);
NAND #() 
NAND_2831_ (
  .A({ datapath_addsubunit_in1_9 }),
  .B({ S4385 }),
  .Y({ S4388 })
);
NOR #() 
NOR_1319_ (
  .A({ datapath_addsubunit_in1_9 }),
  .B({ S4385 }),
  .Y({ S4389 })
);
NAND #() 
NAND_2832_ (
  .A({ S754 }),
  .B({ S4386 }),
  .Y({ S4390 })
);
NOR #() 
NOR_1320_ (
  .A({ S4387 }),
  .B({ S4389 }),
  .Y({ S4391 })
);
NAND #() 
NAND_2833_ (
  .A({ S4388 }),
  .B({ S4390 }),
  .Y({ S4392 })
);
NOR #() 
NOR_1321_ (
  .A({ S1745 }),
  .B({ S4392 }),
  .Y({ S4393 })
);
NAND #() 
NAND_2834_ (
  .A({ S1746 }),
  .B({ S4391 }),
  .Y({ S4394 })
);
NOR #() 
NOR_1322_ (
  .A({ datapath_addsubunit_in1_8 }),
  .B({ S1516 }),
  .Y({ S4395 })
);
NAND #() 
NAND_2835_ (
  .A({ S805 }),
  .B({ S1515 }),
  .Y({ S4396 })
);
NOR #() 
NOR_1323_ (
  .A({ S1746 }),
  .B({ S4391 }),
  .Y({ S4397 })
);
NAND #() 
NAND_2836_ (
  .A({ S1745 }),
  .B({ S4392 }),
  .Y({ S4398 })
);
NOR #() 
NOR_1324_ (
  .A({ S4393 }),
  .B({ S4397 }),
  .Y({ S4399 })
);
NAND #() 
NAND_2837_ (
  .A({ S4394 }),
  .B({ S4398 }),
  .Y({ S4400 })
);
NOR #() 
NOR_1325_ (
  .A({ S4395 }),
  .B({ S4400 }),
  .Y({ S4401 })
);
NAND #() 
NAND_2838_ (
  .A({ S4396 }),
  .B({ S4399 }),
  .Y({ S4402 })
);
NOR #() 
NOR_1326_ (
  .A({ S4393 }),
  .B({ S4401 }),
  .Y({ S4403 })
);
NAND #() 
NAND_2839_ (
  .A({ S4394 }),
  .B({ S4402 }),
  .Y({ S4404 })
);
NOR #() 
NOR_1327_ (
  .A({ S4384 }),
  .B({ S4403 }),
  .Y({ S4405 })
);
NAND #() 
NAND_2840_ (
  .A({ S4383 }),
  .B({ S4404 }),
  .Y({ S4406 })
);
NOR #() 
NOR_1328_ (
  .A({ S4379 }),
  .B({ S4405 }),
  .Y({ S4407 })
);
NAND #() 
NAND_2841_ (
  .A({ S4380 }),
  .B({ S4406 }),
  .Y({ S4408 })
);
NOR #() 
NOR_1329_ (
  .A({ S4370 }),
  .B({ S4407 }),
  .Y({ S4409 })
);
NAND #() 
NAND_2842_ (
  .A({ S4369 }),
  .B({ S4408 }),
  .Y({ S4410 })
);
NOR #() 
NOR_1330_ (
  .A({ S4365 }),
  .B({ S4409 }),
  .Y({ S4411 })
);
NAND #() 
NAND_2843_ (
  .A({ S4366 }),
  .B({ S4410 }),
  .Y({ S4412 })
);
NOR #() 
NOR_1331_ (
  .A({ S4356 }),
  .B({ S4411 }),
  .Y({ S4413 })
);
NAND #() 
NAND_2844_ (
  .A({ S4355 }),
  .B({ S4412 }),
  .Y({ S4414 })
);
NOR #() 
NOR_1332_ (
  .A({ S4351 }),
  .B({ S4413 }),
  .Y({ S4415 })
);
NAND #() 
NAND_2845_ (
  .A({ S4352 }),
  .B({ S4414 }),
  .Y({ S4416 })
);
NOR #() 
NOR_1333_ (
  .A({ S4342 }),
  .B({ S4415 }),
  .Y({ S4417 })
);
NAND #() 
NAND_2846_ (
  .A({ S4341 }),
  .B({ S4416 }),
  .Y({ S4418 })
);
NOR #() 
NOR_1334_ (
  .A({ S4337 }),
  .B({ S4417 }),
  .Y({ S4419 })
);
NAND #() 
NAND_2847_ (
  .A({ S4338 }),
  .B({ S4418 }),
  .Y({ S4420 })
);
NOR #() 
NOR_1335_ (
  .A({ S4328 }),
  .B({ S4419 }),
  .Y({ S4421 })
);
NAND #() 
NAND_2848_ (
  .A({ S4327 }),
  .B({ S4420 }),
  .Y({ S4422 })
);
NOR #() 
NOR_1336_ (
  .A({ S4323 }),
  .B({ S4421 }),
  .Y({ S4423 })
);
NAND #() 
NAND_2849_ (
  .A({ S4324 }),
  .B({ S4422 }),
  .Y({ S4424 })
);
NOR #() 
NOR_1337_ (
  .A({ S4306 }),
  .B({ S4423 }),
  .Y({ S4425 })
);
NAND #() 
NAND_2850_ (
  .A({ S4305 }),
  .B({ S4424 }),
  .Y({ S4426 })
);
NOR #() 
NOR_1338_ (
  .A({ S4302 }),
  .B({ S4425 }),
  .Y({ S4427 })
);
NAND #() 
NAND_2851_ (
  .A({ S4303 }),
  .B({ S4426 }),
  .Y({ S4428 })
);
NOR #() 
NOR_1339_ (
  .A({ S3913 }),
  .B({ S4427 }),
  .Y({ S4429 })
);
NAND #() 
NAND_2852_ (
  .A({ S3912 }),
  .B({ S4428 }),
  .Y({ S4430 })
);
NOR #() 
NOR_1340_ (
  .A({ S4327 }),
  .B({ S4420 }),
  .Y({ S4431 })
);
NAND #() 
NAND_2853_ (
  .A({ S4328 }),
  .B({ S4419 }),
  .Y({ S4432 })
);
NOR #() 
NOR_1341_ (
  .A({ S4421 }),
  .B({ S4431 }),
  .Y({ S4433 })
);
NAND #() 
NAND_2854_ (
  .A({ S4422 }),
  .B({ S4432 }),
  .Y({ S4434 })
);
NOR #() 
NOR_1342_ (
  .A({ S4430 }),
  .B({ S4433 }),
  .Y({ S4435 })
);
NAND #() 
NAND_2855_ (
  .A({ S4429 }),
  .B({ S4434 }),
  .Y({ S4436 })
);
NOR #() 
NOR_1343_ (
  .A({ S4321 }),
  .B({ S4429 }),
  .Y({ S4437 })
);
NAND #() 
NAND_2856_ (
  .A({ S4322 }),
  .B({ S4430 }),
  .Y({ S4438 })
);
NOR #() 
NOR_1344_ (
  .A({ S4435 }),
  .B({ S4437 }),
  .Y({ S4439 })
);
NAND #() 
NAND_2857_ (
  .A({ S4436 }),
  .B({ S4438 }),
  .Y({ S4440 })
);
NOR #() 
NOR_1345_ (
  .A({ S2311 }),
  .B({ S4440 }),
  .Y({ S4441 })
);
NAND #() 
NAND_2858_ (
  .A({ S2312 }),
  .B({ S4439 }),
  .Y({ S4442 })
);
NOR #() 
NOR_1346_ (
  .A({ S2312 }),
  .B({ S4439 }),
  .Y({ S4443 })
);
NAND #() 
NAND_2859_ (
  .A({ S2311 }),
  .B({ S4440 }),
  .Y({ S4444 })
);
NOR #() 
NOR_1347_ (
  .A({ S4441 }),
  .B({ S4443 }),
  .Y({ S4445 })
);
NAND #() 
NAND_2860_ (
  .A({ S4442 }),
  .B({ S4444 }),
  .Y({ S4446 })
);
NAND #() 
NAND_2861_ (
  .A({ S4342 }),
  .B({ S4415 }),
  .Y({ S4447 })
);
NAND #() 
NAND_2862_ (
  .A({ S4418 }),
  .B({ S4447 }),
  .Y({ S4448 })
);
NAND #() 
NAND_2863_ (
  .A({ S4429 }),
  .B({ S4448 }),
  .Y({ S4449 })
);
NAND #() 
NAND_2864_ (
  .A({ S4336 }),
  .B({ S4430 }),
  .Y({ S4450 })
);
NAND #() 
NAND_2865_ (
  .A({ S4449 }),
  .B({ S4450 }),
  .Y({ S4451 })
);
NOT #() 
NOT_348_ (
  .A({ S4451 }),
  .Y({ S4452 })
);
NAND #() 
NAND_2866_ (
  .A({ S2206 }),
  .B({ S4452 }),
  .Y({ S4453 })
);
NAND #() 
NAND_2867_ (
  .A({ S2205 }),
  .B({ S4451 }),
  .Y({ S4454 })
);
NAND #() 
NAND_2868_ (
  .A({ S4356 }),
  .B({ S4411 }),
  .Y({ S4455 })
);
NAND #() 
NAND_2869_ (
  .A({ S4414 }),
  .B({ S4455 }),
  .Y({ S4456 })
);
NAND #() 
NAND_2870_ (
  .A({ S4429 }),
  .B({ S4456 }),
  .Y({ S4457 })
);
NAND #() 
NAND_2871_ (
  .A({ S4350 }),
  .B({ S4430 }),
  .Y({ S4458 })
);
NAND #() 
NAND_2872_ (
  .A({ S4457 }),
  .B({ S4458 }),
  .Y({ S4459 })
);
NOT #() 
NOT_349_ (
  .A({ S4459 }),
  .Y({ S4460 })
);
NOR #() 
NOR_1348_ (
  .A({ S2106 }),
  .B({ S4459 }),
  .Y({ S4461 })
);
NAND #() 
NAND_2873_ (
  .A({ S2107 }),
  .B({ S4460 }),
  .Y({ S4462 })
);
NAND #() 
NAND_2874_ (
  .A({ S2106 }),
  .B({ S4459 }),
  .Y({ S4463 })
);
NOT #() 
NOT_350_ (
  .A({ S4463 }),
  .Y({ S4464 })
);
NOR #() 
NOR_1349_ (
  .A({ S4461 }),
  .B({ S4464 }),
  .Y({ S4465 })
);
NOT #() 
NOT_351_ (
  .A({ S4465 }),
  .Y({ S4466 })
);
NOR #() 
NOR_1350_ (
  .A({ S4363 }),
  .B({ S4429 }),
  .Y({ S4467 })
);
NAND #() 
NAND_2875_ (
  .A({ S4364 }),
  .B({ S4430 }),
  .Y({ S4468 })
);
NOR #() 
NOR_1351_ (
  .A({ S4369 }),
  .B({ S4408 }),
  .Y({ S4469 })
);
NAND #() 
NAND_2876_ (
  .A({ S4370 }),
  .B({ S4407 }),
  .Y({ S4470 })
);
NOR #() 
NOR_1352_ (
  .A({ S4409 }),
  .B({ S4469 }),
  .Y({ S4471 })
);
NAND #() 
NAND_2877_ (
  .A({ S4410 }),
  .B({ S4470 }),
  .Y({ S4472 })
);
NOR #() 
NOR_1353_ (
  .A({ S4430 }),
  .B({ S4471 }),
  .Y({ S4473 })
);
NAND #() 
NAND_2878_ (
  .A({ S4429 }),
  .B({ S4472 }),
  .Y({ S4474 })
);
NOR #() 
NOR_1354_ (
  .A({ S4467 }),
  .B({ S4473 }),
  .Y({ S4475 })
);
NAND #() 
NAND_2879_ (
  .A({ S4468 }),
  .B({ S4474 }),
  .Y({ S4476 })
);
NOR #() 
NOR_1355_ (
  .A({ S1597 }),
  .B({ S4476 }),
  .Y({ S4477 })
);
NAND #() 
NAND_2880_ (
  .A({ S1598 }),
  .B({ S4475 }),
  .Y({ S4478 })
);
NOR #() 
NOR_1356_ (
  .A({ S1598 }),
  .B({ S4475 }),
  .Y({ S4479 })
);
NAND #() 
NAND_2881_ (
  .A({ S1597 }),
  .B({ S4476 }),
  .Y({ S4480 })
);
NOR #() 
NOR_1357_ (
  .A({ S4477 }),
  .B({ S4479 }),
  .Y({ S4481 })
);
NAND #() 
NAND_2882_ (
  .A({ S4478 }),
  .B({ S4480 }),
  .Y({ S4482 })
);
NOR #() 
NOR_1358_ (
  .A({ S4383 }),
  .B({ S4404 }),
  .Y({ S4483 })
);
NAND #() 
NAND_2883_ (
  .A({ S4384 }),
  .B({ S4403 }),
  .Y({ S4484 })
);
NOR #() 
NOR_1359_ (
  .A({ S4405 }),
  .B({ S4483 }),
  .Y({ S4485 })
);
NAND #() 
NAND_2884_ (
  .A({ S4406 }),
  .B({ S4484 }),
  .Y({ S4486 })
);
NOR #() 
NOR_1360_ (
  .A({ S4430 }),
  .B({ S4485 }),
  .Y({ S4487 })
);
NAND #() 
NAND_2885_ (
  .A({ S4429 }),
  .B({ S4486 }),
  .Y({ S4488 })
);
NOR #() 
NOR_1361_ (
  .A({ S4377 }),
  .B({ S4429 }),
  .Y({ S4489 })
);
NAND #() 
NAND_2886_ (
  .A({ S4378 }),
  .B({ S4430 }),
  .Y({ S4490 })
);
NOR #() 
NOR_1362_ (
  .A({ S4487 }),
  .B({ S4489 }),
  .Y({ S4491 })
);
NAND #() 
NAND_2887_ (
  .A({ S4488 }),
  .B({ S4490 }),
  .Y({ S4492 })
);
NOR #() 
NOR_1363_ (
  .A({ S1952 }),
  .B({ S4492 }),
  .Y({ S4493 })
);
NAND #() 
NAND_2888_ (
  .A({ S1953 }),
  .B({ S4491 }),
  .Y({ S4494 })
);
NOR #() 
NOR_1364_ (
  .A({ S1953 }),
  .B({ S4491 }),
  .Y({ S4495 })
);
NAND #() 
NAND_2889_ (
  .A({ S1952 }),
  .B({ S4492 }),
  .Y({ S4496 })
);
NOR #() 
NOR_1365_ (
  .A({ S4493 }),
  .B({ S4495 }),
  .Y({ S4497 })
);
NAND #() 
NAND_2890_ (
  .A({ S4494 }),
  .B({ S4496 }),
  .Y({ S4498 })
);
NOR #() 
NOR_1366_ (
  .A({ S4396 }),
  .B({ S4399 }),
  .Y({ S4499 })
);
NAND #() 
NAND_2891_ (
  .A({ S4395 }),
  .B({ S4400 }),
  .Y({ S4500 })
);
NOR #() 
NOR_1367_ (
  .A({ S4401 }),
  .B({ S4499 }),
  .Y({ S4501 })
);
NAND #() 
NAND_2892_ (
  .A({ S4402 }),
  .B({ S4500 }),
  .Y({ S4502 })
);
NOR #() 
NOR_1368_ (
  .A({ S4430 }),
  .B({ S4501 }),
  .Y({ S4503 })
);
NAND #() 
NAND_2893_ (
  .A({ S4429 }),
  .B({ S4502 }),
  .Y({ S4504 })
);
NOR #() 
NOR_1369_ (
  .A({ S4391 }),
  .B({ S4429 }),
  .Y({ S4505 })
);
NAND #() 
NAND_2894_ (
  .A({ S4392 }),
  .B({ S4430 }),
  .Y({ S4506 })
);
NOR #() 
NOR_1370_ (
  .A({ S4503 }),
  .B({ S4505 }),
  .Y({ S4507 })
);
NAND #() 
NAND_2895_ (
  .A({ S4504 }),
  .B({ S4506 }),
  .Y({ S4508 })
);
NOR #() 
NOR_1371_ (
  .A({ S1848 }),
  .B({ S4508 }),
  .Y({ S4509 })
);
NAND #() 
NAND_2896_ (
  .A({ S1849 }),
  .B({ S4507 }),
  .Y({ S4510 })
);
NOR #() 
NOR_1372_ (
  .A({ S1849 }),
  .B({ S4507 }),
  .Y({ S4511 })
);
NAND #() 
NAND_2897_ (
  .A({ S1848 }),
  .B({ S4508 }),
  .Y({ S4512 })
);
NOR #() 
NOR_1373_ (
  .A({ S4509 }),
  .B({ S4511 }),
  .Y({ S4513 })
);
NAND #() 
NAND_2898_ (
  .A({ S4510 }),
  .B({ S4512 }),
  .Y({ S4514 })
);
NOR #() 
NOR_1374_ (
  .A({ S1516 }),
  .B({ S4430 }),
  .Y({ S4515 })
);
NAND #() 
NAND_2899_ (
  .A({ S1515 }),
  .B({ S4429 }),
  .Y({ S4516 })
);
NOR #() 
NOR_1375_ (
  .A({ S805 }),
  .B({ S4515 }),
  .Y({ S4517 })
);
NAND #() 
NAND_2900_ (
  .A({ datapath_addsubunit_in1_8 }),
  .B({ S4516 }),
  .Y({ S4518 })
);
NOR #() 
NOR_1376_ (
  .A({ S4396 }),
  .B({ S4430 }),
  .Y({ S4519 })
);
NAND #() 
NAND_2901_ (
  .A({ S4395 }),
  .B({ S4429 }),
  .Y({ S4520 })
);
NOR #() 
NOR_1377_ (
  .A({ S4517 }),
  .B({ S4519 }),
  .Y({ S4521 })
);
NAND #() 
NAND_2902_ (
  .A({ S4518 }),
  .B({ S4520 }),
  .Y({ S4522 })
);
NOR #() 
NOR_1378_ (
  .A({ S1745 }),
  .B({ S4521 }),
  .Y({ S4523 })
);
NAND #() 
NAND_2903_ (
  .A({ S1746 }),
  .B({ S4522 }),
  .Y({ S4524 })
);
NAND #() 
NAND_2904_ (
  .A({ S858 }),
  .B({ S1515 }),
  .Y({ S4525 })
);
NOT #() 
NOT_352_ (
  .A({ S4525 }),
  .Y({ S4526 })
);
NOR #() 
NOR_1379_ (
  .A({ S1746 }),
  .B({ S4522 }),
  .Y({ S4527 })
);
NAND #() 
NAND_2905_ (
  .A({ S1745 }),
  .B({ S4521 }),
  .Y({ S4528 })
);
NOR #() 
NOR_1380_ (
  .A({ S4523 }),
  .B({ S4527 }),
  .Y({ S4529 })
);
NAND #() 
NAND_2906_ (
  .A({ S4524 }),
  .B({ S4528 }),
  .Y({ S4530 })
);
NOR #() 
NOR_1381_ (
  .A({ S4526 }),
  .B({ S4530 }),
  .Y({ S4531 })
);
NAND #() 
NAND_2907_ (
  .A({ S4525 }),
  .B({ S4529 }),
  .Y({ S4532 })
);
NOR #() 
NOR_1382_ (
  .A({ S4523 }),
  .B({ S4531 }),
  .Y({ S4533 })
);
NAND #() 
NAND_2908_ (
  .A({ S4524 }),
  .B({ S4532 }),
  .Y({ S4534 })
);
NOR #() 
NOR_1383_ (
  .A({ S4514 }),
  .B({ S4533 }),
  .Y({ S4535 })
);
NAND #() 
NAND_2909_ (
  .A({ S4513 }),
  .B({ S4534 }),
  .Y({ S4536 })
);
NOR #() 
NOR_1384_ (
  .A({ S4509 }),
  .B({ S4535 }),
  .Y({ S4537 })
);
NAND #() 
NAND_2910_ (
  .A({ S4510 }),
  .B({ S4536 }),
  .Y({ S4538 })
);
NOR #() 
NOR_1385_ (
  .A({ S4498 }),
  .B({ S4537 }),
  .Y({ S4539 })
);
NAND #() 
NAND_2911_ (
  .A({ S4497 }),
  .B({ S4538 }),
  .Y({ S4540 })
);
NOR #() 
NOR_1386_ (
  .A({ S4493 }),
  .B({ S4539 }),
  .Y({ S4541 })
);
NAND #() 
NAND_2912_ (
  .A({ S4494 }),
  .B({ S4540 }),
  .Y({ S4542 })
);
NOR #() 
NOR_1387_ (
  .A({ S4482 }),
  .B({ S4541 }),
  .Y({ S4543 })
);
NAND #() 
NAND_2913_ (
  .A({ S4481 }),
  .B({ S4542 }),
  .Y({ S4544 })
);
NOR #() 
NOR_1388_ (
  .A({ S4477 }),
  .B({ S4543 }),
  .Y({ S4545 })
);
NAND #() 
NAND_2914_ (
  .A({ S4478 }),
  .B({ S4544 }),
  .Y({ S4546 })
);
NOR #() 
NOR_1389_ (
  .A({ S4466 }),
  .B({ S4545 }),
  .Y({ S4547 })
);
NAND #() 
NAND_2915_ (
  .A({ S4465 }),
  .B({ S4546 }),
  .Y({ S4548 })
);
NOR #() 
NOR_1390_ (
  .A({ S4461 }),
  .B({ S4547 }),
  .Y({ S4549 })
);
NAND #() 
NAND_2916_ (
  .A({ S4462 }),
  .B({ S4548 }),
  .Y({ S4550 })
);
NAND #() 
NAND_2917_ (
  .A({ S4454 }),
  .B({ S4550 }),
  .Y({ S4551 })
);
NAND #() 
NAND_2918_ (
  .A({ S4453 }),
  .B({ S4549 }),
  .Y({ S4552 })
);
NAND #() 
NAND_2919_ (
  .A({ S4454 }),
  .B({ S4552 }),
  .Y({ S4553 })
);
NAND #() 
NAND_2920_ (
  .A({ S4453 }),
  .B({ S4551 }),
  .Y({ S4554 })
);
NOR #() 
NOR_1391_ (
  .A({ S4446 }),
  .B({ S4553 }),
  .Y({ S4555 })
);
NAND #() 
NAND_2921_ (
  .A({ S4445 }),
  .B({ S4554 }),
  .Y({ S4556 })
);
NOR #() 
NOR_1392_ (
  .A({ S4441 }),
  .B({ S4555 }),
  .Y({ S4557 })
);
NAND #() 
NAND_2922_ (
  .A({ S4442 }),
  .B({ S4556 }),
  .Y({ S4558 })
);
NOR #() 
NOR_1393_ (
  .A({ S4300 }),
  .B({ S4429 }),
  .Y({ S4559 })
);
NOR #() 
NOR_1394_ (
  .A({ S3950 }),
  .B({ S4559 }),
  .Y({ S4560 })
);
NOT #() 
NOT_353_ (
  .A({ S4560 }),
  .Y({ S4561 })
);
NOR #() 
NOR_1395_ (
  .A({ S2417 }),
  .B({ S4560 }),
  .Y({ S4562 })
);
NAND #() 
NAND_2923_ (
  .A({ S2418 }),
  .B({ S4561 }),
  .Y({ S4563 })
);
NOR #() 
NOR_1396_ (
  .A({ S4558 }),
  .B({ S4562 }),
  .Y({ S4564 })
);
NAND #() 
NAND_2924_ (
  .A({ S4557 }),
  .B({ S4563 }),
  .Y({ S4565 })
);
NOR #() 
NOR_1397_ (
  .A({ S2418 }),
  .B({ S4561 }),
  .Y({ S4566 })
);
NAND #() 
NAND_2925_ (
  .A({ S2417 }),
  .B({ S4560 }),
  .Y({ S4567 })
);
NOR #() 
NOR_1398_ (
  .A({ S3911 }),
  .B({ S4566 }),
  .Y({ S4568 })
);
NAND #() 
NAND_2926_ (
  .A({ S3910 }),
  .B({ S4567 }),
  .Y({ S4569 })
);
NOR #() 
NOR_1399_ (
  .A({ S4564 }),
  .B({ S4569 }),
  .Y({ S4570 })
);
NAND #() 
NAND_2927_ (
  .A({ S4565 }),
  .B({ S4568 }),
  .Y({ S4571 })
);
NOR #() 
NOR_1400_ (
  .A({ S4445 }),
  .B({ S4554 }),
  .Y({ S4572 })
);
NOR #() 
NOR_1401_ (
  .A({ S4555 }),
  .B({ S4572 }),
  .Y({ S4573 })
);
NOR #() 
NOR_1402_ (
  .A({ S4571 }),
  .B({ S4573 }),
  .Y({ S4574 })
);
NOR #() 
NOR_1403_ (
  .A({ S4439 }),
  .B({ S4570 }),
  .Y({ S4575 })
);
NOR #() 
NOR_1404_ (
  .A({ S4574 }),
  .B({ S4575 }),
  .Y({ S4576 })
);
NOT #() 
NOT_354_ (
  .A({ S4576 }),
  .Y({ S4577 })
);
NOR #() 
NOR_1405_ (
  .A({ S2417 }),
  .B({ S4577 }),
  .Y({ S4578 })
);
NAND #() 
NAND_2928_ (
  .A({ S2418 }),
  .B({ S4576 }),
  .Y({ S4579 })
);
NOR #() 
NOR_1406_ (
  .A({ S2418 }),
  .B({ S4576 }),
  .Y({ S4580 })
);
NOT #() 
NOT_355_ (
  .A({ S4580 }),
  .Y({ S4581 })
);
NAND #() 
NAND_2929_ (
  .A({ S4579 }),
  .B({ S4581 }),
  .Y({ S4582 })
);
NOT #() 
NOT_356_ (
  .A({ S4582 }),
  .Y({ S4583 })
);
NAND #() 
NAND_2930_ (
  .A({ S4453 }),
  .B({ S4454 }),
  .Y({ S4584 })
);
NAND #() 
NAND_2931_ (
  .A({ S4549 }),
  .B({ S4584 }),
  .Y({ S4585 })
);
NOT #() 
NOT_357_ (
  .A({ S4585 }),
  .Y({ S4586 })
);
NOR #() 
NOR_1407_ (
  .A({ S4549 }),
  .B({ S4584 }),
  .Y({ S4587 })
);
NOR #() 
NOR_1408_ (
  .A({ S4586 }),
  .B({ S4587 }),
  .Y({ S4588 })
);
NOR #() 
NOR_1409_ (
  .A({ S4571 }),
  .B({ S4588 }),
  .Y({ S4589 })
);
NOR #() 
NOR_1410_ (
  .A({ S4452 }),
  .B({ S4570 }),
  .Y({ S4590 })
);
NOR #() 
NOR_1411_ (
  .A({ S4589 }),
  .B({ S4590 }),
  .Y({ S4591 })
);
NOT #() 
NOT_358_ (
  .A({ S4591 }),
  .Y({ S4592 })
);
NOR #() 
NOR_1412_ (
  .A({ S2311 }),
  .B({ S4592 }),
  .Y({ S4593 })
);
NOR #() 
NOR_1413_ (
  .A({ S2312 }),
  .B({ S4591 }),
  .Y({ S4594 })
);
NOR #() 
NOR_1414_ (
  .A({ S4465 }),
  .B({ S4546 }),
  .Y({ S4595 })
);
NOR #() 
NOR_1415_ (
  .A({ S4547 }),
  .B({ S4595 }),
  .Y({ S4596 })
);
NOR #() 
NOR_1416_ (
  .A({ S4571 }),
  .B({ S4596 }),
  .Y({ S4597 })
);
NOR #() 
NOR_1417_ (
  .A({ S4460 }),
  .B({ S4570 }),
  .Y({ S4598 })
);
NOR #() 
NOR_1418_ (
  .A({ S4597 }),
  .B({ S4598 }),
  .Y({ S4599 })
);
NOT #() 
NOT_359_ (
  .A({ S4599 }),
  .Y({ S4600 })
);
NOR #() 
NOR_1419_ (
  .A({ S2205 }),
  .B({ S4600 }),
  .Y({ S4601 })
);
NAND #() 
NAND_2932_ (
  .A({ S2206 }),
  .B({ S4599 }),
  .Y({ S4602 })
);
NAND #() 
NAND_2933_ (
  .A({ S2205 }),
  .B({ S4600 }),
  .Y({ S4603 })
);
NAND #() 
NAND_2934_ (
  .A({ S4602 }),
  .B({ S4603 }),
  .Y({ S4604 })
);
NOT #() 
NOT_360_ (
  .A({ S4604 }),
  .Y({ S4605 })
);
NOR #() 
NOR_1420_ (
  .A({ S4481 }),
  .B({ S4542 }),
  .Y({ S4606 })
);
NOR #() 
NOR_1421_ (
  .A({ S4543 }),
  .B({ S4606 }),
  .Y({ S4607 })
);
NOR #() 
NOR_1422_ (
  .A({ S4571 }),
  .B({ S4607 }),
  .Y({ S4608 })
);
NOR #() 
NOR_1423_ (
  .A({ S4475 }),
  .B({ S4570 }),
  .Y({ S4609 })
);
NOR #() 
NOR_1424_ (
  .A({ S4608 }),
  .B({ S4609 }),
  .Y({ S4610 })
);
NOT #() 
NOT_361_ (
  .A({ S4610 }),
  .Y({ S4611 })
);
NOR #() 
NOR_1425_ (
  .A({ S2106 }),
  .B({ S4611 }),
  .Y({ S4612 })
);
NAND #() 
NAND_2935_ (
  .A({ S2107 }),
  .B({ S4610 }),
  .Y({ S4613 })
);
NAND #() 
NAND_2936_ (
  .A({ S2106 }),
  .B({ S4611 }),
  .Y({ S4614 })
);
NAND #() 
NAND_2937_ (
  .A({ S4613 }),
  .B({ S4614 }),
  .Y({ S4615 })
);
NOT #() 
NOT_362_ (
  .A({ S4615 }),
  .Y({ S4616 })
);
NOR #() 
NOR_1426_ (
  .A({ S4491 }),
  .B({ S4570 }),
  .Y({ S4617 })
);
NOR #() 
NOR_1427_ (
  .A({ S4497 }),
  .B({ S4538 }),
  .Y({ S4618 })
);
NOR #() 
NOR_1428_ (
  .A({ S4539 }),
  .B({ S4618 }),
  .Y({ S4619 })
);
NOR #() 
NOR_1429_ (
  .A({ S4571 }),
  .B({ S4619 }),
  .Y({ S4620 })
);
NOR #() 
NOR_1430_ (
  .A({ S4617 }),
  .B({ S4620 }),
  .Y({ S4621 })
);
NOT #() 
NOT_363_ (
  .A({ S4621 }),
  .Y({ S4622 })
);
NOR #() 
NOR_1431_ (
  .A({ S1597 }),
  .B({ S4622 }),
  .Y({ S4623 })
);
NAND #() 
NAND_2938_ (
  .A({ S1598 }),
  .B({ S4621 }),
  .Y({ S4624 })
);
NAND #() 
NAND_2939_ (
  .A({ S1597 }),
  .B({ S4622 }),
  .Y({ S4625 })
);
NAND #() 
NAND_2940_ (
  .A({ S4624 }),
  .B({ S4625 }),
  .Y({ S4626 })
);
NOT #() 
NOT_364_ (
  .A({ S4626 }),
  .Y({ S4627 })
);
NOR #() 
NOR_1432_ (
  .A({ S4513 }),
  .B({ S4534 }),
  .Y({ S4628 })
);
NOR #() 
NOR_1433_ (
  .A({ S4535 }),
  .B({ S4628 }),
  .Y({ S4629 })
);
NOR #() 
NOR_1434_ (
  .A({ S4571 }),
  .B({ S4629 }),
  .Y({ S4630 })
);
NOR #() 
NOR_1435_ (
  .A({ S4507 }),
  .B({ S4570 }),
  .Y({ S4631 })
);
NOR #() 
NOR_1436_ (
  .A({ S4630 }),
  .B({ S4631 }),
  .Y({ S4632 })
);
NOT #() 
NOT_365_ (
  .A({ S4632 }),
  .Y({ S4633 })
);
NAND #() 
NAND_2941_ (
  .A({ S1953 }),
  .B({ S4632 }),
  .Y({ S4634 })
);
NAND #() 
NAND_2942_ (
  .A({ S1952 }),
  .B({ S4633 }),
  .Y({ S4635 })
);
NOR #() 
NOR_1437_ (
  .A({ S4525 }),
  .B({ S4529 }),
  .Y({ S4636 })
);
NOR #() 
NOR_1438_ (
  .A({ S4531 }),
  .B({ S4636 }),
  .Y({ S4637 })
);
NOR #() 
NOR_1439_ (
  .A({ S4571 }),
  .B({ S4637 }),
  .Y({ S4638 })
);
NOR #() 
NOR_1440_ (
  .A({ S4522 }),
  .B({ S4570 }),
  .Y({ S4639 })
);
NOR #() 
NOR_1441_ (
  .A({ S4638 }),
  .B({ S4639 }),
  .Y({ S4640 })
);
NOT #() 
NOT_366_ (
  .A({ S4640 }),
  .Y({ S4641 })
);
NOR #() 
NOR_1442_ (
  .A({ S1848 }),
  .B({ S4641 }),
  .Y({ S4642 })
);
NAND #() 
NAND_2943_ (
  .A({ S1849 }),
  .B({ S4640 }),
  .Y({ S4643 })
);
NOR #() 
NOR_1443_ (
  .A({ S1516 }),
  .B({ S4571 }),
  .Y({ S4644 })
);
NAND #() 
NAND_2944_ (
  .A({ S1515 }),
  .B({ S4570 }),
  .Y({ S4645 })
);
NOR #() 
NOR_1444_ (
  .A({ S858 }),
  .B({ S4644 }),
  .Y({ S4646 })
);
NAND #() 
NAND_2945_ (
  .A({ datapath_addsubunit_in1_7 }),
  .B({ S4645 }),
  .Y({ S4647 })
);
NOR #() 
NOR_1445_ (
  .A({ datapath_addsubunit_in1_7 }),
  .B({ S4645 }),
  .Y({ S4648 })
);
NAND #() 
NAND_2946_ (
  .A({ S858 }),
  .B({ S4644 }),
  .Y({ S4649 })
);
NOR #() 
NOR_1446_ (
  .A({ S4646 }),
  .B({ S4648 }),
  .Y({ S4650 })
);
NAND #() 
NAND_2947_ (
  .A({ S4647 }),
  .B({ S4649 }),
  .Y({ S4651 })
);
NOR #() 
NOR_1447_ (
  .A({ S1745 }),
  .B({ S4650 }),
  .Y({ S4652 })
);
NAND #() 
NAND_2948_ (
  .A({ S1746 }),
  .B({ S4651 }),
  .Y({ S4653 })
);
NAND #() 
NAND_2949_ (
  .A({ S910 }),
  .B({ S1515 }),
  .Y({ S4654 })
);
NOT #() 
NOT_367_ (
  .A({ S4654 }),
  .Y({ S4655 })
);
NOR #() 
NOR_1448_ (
  .A({ S1746 }),
  .B({ S4651 }),
  .Y({ S4656 })
);
NAND #() 
NAND_2950_ (
  .A({ S1745 }),
  .B({ S4650 }),
  .Y({ S4657 })
);
NOR #() 
NOR_1449_ (
  .A({ S4652 }),
  .B({ S4656 }),
  .Y({ S4658 })
);
NAND #() 
NAND_2951_ (
  .A({ S4653 }),
  .B({ S4657 }),
  .Y({ S4659 })
);
NOR #() 
NOR_1450_ (
  .A({ S4655 }),
  .B({ S4659 }),
  .Y({ S4660 })
);
NAND #() 
NAND_2952_ (
  .A({ S4654 }),
  .B({ S4658 }),
  .Y({ S4661 })
);
NOR #() 
NOR_1451_ (
  .A({ S4652 }),
  .B({ S4660 }),
  .Y({ S4662 })
);
NAND #() 
NAND_2953_ (
  .A({ S4653 }),
  .B({ S4661 }),
  .Y({ S4663 })
);
NAND #() 
NAND_2954_ (
  .A({ S1848 }),
  .B({ S4641 }),
  .Y({ S4664 })
);
NAND #() 
NAND_2955_ (
  .A({ S4643 }),
  .B({ S4664 }),
  .Y({ S4665 })
);
NOT #() 
NOT_368_ (
  .A({ S4665 }),
  .Y({ S4666 })
);
NOR #() 
NOR_1452_ (
  .A({ S4662 }),
  .B({ S4665 }),
  .Y({ S4667 })
);
NAND #() 
NAND_2956_ (
  .A({ S4663 }),
  .B({ S4666 }),
  .Y({ S4668 })
);
NOR #() 
NOR_1453_ (
  .A({ S4642 }),
  .B({ S4667 }),
  .Y({ S4669 })
);
NAND #() 
NAND_2957_ (
  .A({ S4643 }),
  .B({ S4668 }),
  .Y({ S4670 })
);
NAND #() 
NAND_2958_ (
  .A({ S4635 }),
  .B({ S4670 }),
  .Y({ S4671 })
);
NAND #() 
NAND_2959_ (
  .A({ S4634 }),
  .B({ S4669 }),
  .Y({ S4672 })
);
NAND #() 
NAND_2960_ (
  .A({ S4635 }),
  .B({ S4672 }),
  .Y({ S4673 })
);
NAND #() 
NAND_2961_ (
  .A({ S4634 }),
  .B({ S4671 }),
  .Y({ S4674 })
);
NOR #() 
NOR_1454_ (
  .A({ S4626 }),
  .B({ S4673 }),
  .Y({ S4675 })
);
NAND #() 
NAND_2962_ (
  .A({ S4627 }),
  .B({ S4674 }),
  .Y({ S4676 })
);
NOR #() 
NOR_1455_ (
  .A({ S4623 }),
  .B({ S4675 }),
  .Y({ S4677 })
);
NAND #() 
NAND_2963_ (
  .A({ S4624 }),
  .B({ S4676 }),
  .Y({ S4678 })
);
NOR #() 
NOR_1456_ (
  .A({ S4615 }),
  .B({ S4677 }),
  .Y({ S4679 })
);
NAND #() 
NAND_2964_ (
  .A({ S4616 }),
  .B({ S4678 }),
  .Y({ S4680 })
);
NOR #() 
NOR_1457_ (
  .A({ S4612 }),
  .B({ S4679 }),
  .Y({ S4681 })
);
NAND #() 
NAND_2965_ (
  .A({ S4613 }),
  .B({ S4680 }),
  .Y({ S4682 })
);
NOR #() 
NOR_1458_ (
  .A({ S4604 }),
  .B({ S4681 }),
  .Y({ S4683 })
);
NAND #() 
NAND_2966_ (
  .A({ S4605 }),
  .B({ S4682 }),
  .Y({ S4684 })
);
NOR #() 
NOR_1459_ (
  .A({ S4601 }),
  .B({ S4683 }),
  .Y({ S4685 })
);
NAND #() 
NAND_2967_ (
  .A({ S4602 }),
  .B({ S4684 }),
  .Y({ S4686 })
);
NOR #() 
NOR_1460_ (
  .A({ S4594 }),
  .B({ S4685 }),
  .Y({ S4687 })
);
NOR #() 
NOR_1461_ (
  .A({ S4593 }),
  .B({ S4686 }),
  .Y({ S4688 })
);
NOR #() 
NOR_1462_ (
  .A({ S4593 }),
  .B({ S4687 }),
  .Y({ S4689 })
);
NOR #() 
NOR_1463_ (
  .A({ S4594 }),
  .B({ S4688 }),
  .Y({ S4690 })
);
NOR #() 
NOR_1464_ (
  .A({ S4582 }),
  .B({ S4689 }),
  .Y({ S4691 })
);
NAND #() 
NAND_2968_ (
  .A({ S4583 }),
  .B({ S4690 }),
  .Y({ S4692 })
);
NOR #() 
NOR_1465_ (
  .A({ S4578 }),
  .B({ S4691 }),
  .Y({ S4693 })
);
NAND #() 
NAND_2969_ (
  .A({ S4579 }),
  .B({ S4692 }),
  .Y({ S4694 })
);
NOR #() 
NOR_1466_ (
  .A({ S2418 }),
  .B({ S3911 }),
  .Y({ S4695 })
);
NOR #() 
NOR_1467_ (
  .A({ S4557 }),
  .B({ S4695 }),
  .Y({ S4696 })
);
NOR #() 
NOR_1468_ (
  .A({ S3912 }),
  .B({ S4558 }),
  .Y({ S4697 })
);
NOR #() 
NOR_1469_ (
  .A({ S4696 }),
  .B({ S4697 }),
  .Y({ S4698 })
);
NOR #() 
NOR_1470_ (
  .A({ S4560 }),
  .B({ S4698 }),
  .Y({ S4699 })
);
NOT #() 
NOT_369_ (
  .A({ S4699 }),
  .Y({ S4700 })
);
NOR #() 
NOR_1471_ (
  .A({ S2517 }),
  .B({ S4700 }),
  .Y({ S4701 })
);
NAND #() 
NAND_2970_ (
  .A({ S2518 }),
  .B({ S4699 }),
  .Y({ S4702 })
);
NOR #() 
NOR_1472_ (
  .A({ S4694 }),
  .B({ S4701 }),
  .Y({ S4703 })
);
NAND #() 
NAND_2971_ (
  .A({ S4693 }),
  .B({ S4702 }),
  .Y({ S4704 })
);
NAND #() 
NAND_2972_ (
  .A({ S2517 }),
  .B({ S4560 }),
  .Y({ S4705 })
);
NAND #() 
NAND_2973_ (
  .A({ S3908 }),
  .B({ S4705 }),
  .Y({ S4706 })
);
NOT #() 
NOT_370_ (
  .A({ S4706 }),
  .Y({ S4707 })
);
NOR #() 
NOR_1473_ (
  .A({ S4703 }),
  .B({ S4706 }),
  .Y({ S4708 })
);
NAND #() 
NAND_2974_ (
  .A({ S4704 }),
  .B({ S4707 }),
  .Y({ S4709 })
);
NAND #() 
NAND_2975_ (
  .A({ S4582 }),
  .B({ S4689 }),
  .Y({ S4710 })
);
NAND #() 
NAND_2976_ (
  .A({ S4692 }),
  .B({ S4710 }),
  .Y({ S4711 })
);
NAND #() 
NAND_2977_ (
  .A({ S4708 }),
  .B({ S4711 }),
  .Y({ S4712 })
);
NOT #() 
NOT_371_ (
  .A({ S4712 }),
  .Y({ S4713 })
);
NOR #() 
NOR_1474_ (
  .A({ S4576 }),
  .B({ S4708 }),
  .Y({ S4714 })
);
NOT #() 
NOT_372_ (
  .A({ S4714 }),
  .Y({ S4715 })
);
NOR #() 
NOR_1475_ (
  .A({ S4713 }),
  .B({ S4714 }),
  .Y({ S4716 })
);
NAND #() 
NAND_2978_ (
  .A({ S4712 }),
  .B({ S4715 }),
  .Y({ S4717 })
);
NOR #() 
NOR_1476_ (
  .A({ S2517 }),
  .B({ S4717 }),
  .Y({ S4718 })
);
NAND #() 
NAND_2979_ (
  .A({ S2518 }),
  .B({ S4716 }),
  .Y({ S4719 })
);
NOR #() 
NOR_1477_ (
  .A({ S2518 }),
  .B({ S4716 }),
  .Y({ S4720 })
);
NAND #() 
NAND_2980_ (
  .A({ S2517 }),
  .B({ S4717 }),
  .Y({ S4721 })
);
NOR #() 
NOR_1478_ (
  .A({ S4718 }),
  .B({ S4720 }),
  .Y({ S4722 })
);
NAND #() 
NAND_2981_ (
  .A({ S4719 }),
  .B({ S4721 }),
  .Y({ S4723 })
);
NOR #() 
NOR_1479_ (
  .A({ S4593 }),
  .B({ S4594 }),
  .Y({ S4724 })
);
NOR #() 
NOR_1480_ (
  .A({ S4686 }),
  .B({ S4724 }),
  .Y({ S4725 })
);
NOT #() 
NOT_373_ (
  .A({ S4725 }),
  .Y({ S4726 })
);
NAND #() 
NAND_2982_ (
  .A({ S4686 }),
  .B({ S4724 }),
  .Y({ S4727 })
);
NAND #() 
NAND_2983_ (
  .A({ S4726 }),
  .B({ S4727 }),
  .Y({ S4728 })
);
NAND #() 
NAND_2984_ (
  .A({ S4708 }),
  .B({ S4728 }),
  .Y({ S4729 })
);
NOT #() 
NOT_374_ (
  .A({ S4729 }),
  .Y({ S4730 })
);
NOR #() 
NOR_1481_ (
  .A({ S4591 }),
  .B({ S4708 }),
  .Y({ S4731 })
);
NOT #() 
NOT_375_ (
  .A({ S4731 }),
  .Y({ S4732 })
);
NOR #() 
NOR_1482_ (
  .A({ S4730 }),
  .B({ S4731 }),
  .Y({ S4733 })
);
NAND #() 
NAND_2985_ (
  .A({ S4729 }),
  .B({ S4732 }),
  .Y({ S4734 })
);
NOR #() 
NOR_1483_ (
  .A({ S2417 }),
  .B({ S4734 }),
  .Y({ S4735 })
);
NAND #() 
NAND_2986_ (
  .A({ S2418 }),
  .B({ S4733 }),
  .Y({ S4736 })
);
NOR #() 
NOR_1484_ (
  .A({ S2418 }),
  .B({ S4733 }),
  .Y({ S4737 })
);
NAND #() 
NAND_2987_ (
  .A({ S2417 }),
  .B({ S4734 }),
  .Y({ S4738 })
);
NAND #() 
NAND_2988_ (
  .A({ S4604 }),
  .B({ S4681 }),
  .Y({ S4739 })
);
NAND #() 
NAND_2989_ (
  .A({ S4684 }),
  .B({ S4739 }),
  .Y({ S4740 })
);
NAND #() 
NAND_2990_ (
  .A({ S4708 }),
  .B({ S4740 }),
  .Y({ S4741 })
);
NOT #() 
NOT_376_ (
  .A({ S4741 }),
  .Y({ S4742 })
);
NOR #() 
NOR_1485_ (
  .A({ S4599 }),
  .B({ S4708 }),
  .Y({ S4743 })
);
NOT #() 
NOT_377_ (
  .A({ S4743 }),
  .Y({ S4744 })
);
NOR #() 
NOR_1486_ (
  .A({ S4742 }),
  .B({ S4743 }),
  .Y({ S4745 })
);
NAND #() 
NAND_2991_ (
  .A({ S4741 }),
  .B({ S4744 }),
  .Y({ S4746 })
);
NOR #() 
NOR_1487_ (
  .A({ S2311 }),
  .B({ S4746 }),
  .Y({ S4747 })
);
NAND #() 
NAND_2992_ (
  .A({ S2312 }),
  .B({ S4745 }),
  .Y({ S4748 })
);
NOR #() 
NOR_1488_ (
  .A({ S2312 }),
  .B({ S4745 }),
  .Y({ S4749 })
);
NAND #() 
NAND_2993_ (
  .A({ S2311 }),
  .B({ S4746 }),
  .Y({ S4750 })
);
NOR #() 
NOR_1489_ (
  .A({ S4747 }),
  .B({ S4749 }),
  .Y({ S4751 })
);
NAND #() 
NAND_2994_ (
  .A({ S4748 }),
  .B({ S4750 }),
  .Y({ S4752 })
);
NAND #() 
NAND_2995_ (
  .A({ S4615 }),
  .B({ S4677 }),
  .Y({ S4753 })
);
NAND #() 
NAND_2996_ (
  .A({ S4680 }),
  .B({ S4753 }),
  .Y({ S4754 })
);
NAND #() 
NAND_2997_ (
  .A({ S4708 }),
  .B({ S4754 }),
  .Y({ S4755 })
);
NOT #() 
NOT_378_ (
  .A({ S4755 }),
  .Y({ S4756 })
);
NOR #() 
NOR_1490_ (
  .A({ S4610 }),
  .B({ S4708 }),
  .Y({ S4757 })
);
NOT #() 
NOT_379_ (
  .A({ S4757 }),
  .Y({ S4758 })
);
NOR #() 
NOR_1491_ (
  .A({ S4756 }),
  .B({ S4757 }),
  .Y({ S4759 })
);
NAND #() 
NAND_2998_ (
  .A({ S4755 }),
  .B({ S4758 }),
  .Y({ S4760 })
);
NOR #() 
NOR_1492_ (
  .A({ S2205 }),
  .B({ S4760 }),
  .Y({ S4761 })
);
NAND #() 
NAND_2999_ (
  .A({ S2206 }),
  .B({ S4759 }),
  .Y({ S4762 })
);
NOR #() 
NOR_1493_ (
  .A({ S2206 }),
  .B({ S4759 }),
  .Y({ S4763 })
);
NAND #() 
NAND_3000_ (
  .A({ S2205 }),
  .B({ S4760 }),
  .Y({ S4764 })
);
NOR #() 
NOR_1494_ (
  .A({ S4761 }),
  .B({ S4763 }),
  .Y({ S4765 })
);
NAND #() 
NAND_3001_ (
  .A({ S4762 }),
  .B({ S4764 }),
  .Y({ S4766 })
);
NAND #() 
NAND_3002_ (
  .A({ S4626 }),
  .B({ S4673 }),
  .Y({ S4767 })
);
NAND #() 
NAND_3003_ (
  .A({ S4676 }),
  .B({ S4767 }),
  .Y({ S4768 })
);
NAND #() 
NAND_3004_ (
  .A({ S4708 }),
  .B({ S4768 }),
  .Y({ S4769 })
);
NOT #() 
NOT_380_ (
  .A({ S4769 }),
  .Y({ S4770 })
);
NOR #() 
NOR_1495_ (
  .A({ S4621 }),
  .B({ S4708 }),
  .Y({ S4771 })
);
NOT #() 
NOT_381_ (
  .A({ S4771 }),
  .Y({ S4772 })
);
NOR #() 
NOR_1496_ (
  .A({ S4770 }),
  .B({ S4771 }),
  .Y({ S4773 })
);
NAND #() 
NAND_3005_ (
  .A({ S4769 }),
  .B({ S4772 }),
  .Y({ S4774 })
);
NOR #() 
NOR_1497_ (
  .A({ S2106 }),
  .B({ S4774 }),
  .Y({ S4775 })
);
NAND #() 
NAND_3006_ (
  .A({ S2107 }),
  .B({ S4773 }),
  .Y({ S4776 })
);
NOR #() 
NOR_1498_ (
  .A({ S2107 }),
  .B({ S4773 }),
  .Y({ S4777 })
);
NAND #() 
NAND_3007_ (
  .A({ S2106 }),
  .B({ S4774 }),
  .Y({ S4778 })
);
NOR #() 
NOR_1499_ (
  .A({ S4775 }),
  .B({ S4777 }),
  .Y({ S4779 })
);
NAND #() 
NAND_3008_ (
  .A({ S4776 }),
  .B({ S4778 }),
  .Y({ S4780 })
);
NAND #() 
NAND_3009_ (
  .A({ S4634 }),
  .B({ S4635 }),
  .Y({ S4781 })
);
NOR #() 
NOR_1500_ (
  .A({ S4670 }),
  .B({ S4781 }),
  .Y({ S4782 })
);
NAND #() 
NAND_3010_ (
  .A({ S4670 }),
  .B({ S4781 }),
  .Y({ S4783 })
);
NOT #() 
NOT_382_ (
  .A({ S4783 }),
  .Y({ S4784 })
);
NOR #() 
NOR_1501_ (
  .A({ S4782 }),
  .B({ S4784 }),
  .Y({ S4785 })
);
NAND #() 
NAND_3011_ (
  .A({ S4708 }),
  .B({ S4785 }),
  .Y({ S4786 })
);
NOT #() 
NOT_383_ (
  .A({ S4786 }),
  .Y({ S4787 })
);
NOR #() 
NOR_1502_ (
  .A({ S4632 }),
  .B({ S4708 }),
  .Y({ S4788 })
);
NOT #() 
NOT_384_ (
  .A({ S4788 }),
  .Y({ S4789 })
);
NOR #() 
NOR_1503_ (
  .A({ S4787 }),
  .B({ S4788 }),
  .Y({ S4790 })
);
NAND #() 
NAND_3012_ (
  .A({ S4786 }),
  .B({ S4789 }),
  .Y({ S4791 })
);
NOR #() 
NOR_1504_ (
  .A({ S1597 }),
  .B({ S4791 }),
  .Y({ S4792 })
);
NAND #() 
NAND_3013_ (
  .A({ S1598 }),
  .B({ S4790 }),
  .Y({ S4793 })
);
NOR #() 
NOR_1505_ (
  .A({ S1598 }),
  .B({ S4790 }),
  .Y({ S4794 })
);
NAND #() 
NAND_3014_ (
  .A({ S1597 }),
  .B({ S4791 }),
  .Y({ S4795 })
);
NOR #() 
NOR_1506_ (
  .A({ S4792 }),
  .B({ S4794 }),
  .Y({ S4796 })
);
NAND #() 
NAND_3015_ (
  .A({ S4793 }),
  .B({ S4795 }),
  .Y({ S4797 })
);
NOR #() 
NOR_1507_ (
  .A({ S4640 }),
  .B({ S4708 }),
  .Y({ S4798 })
);
NOT #() 
NOT_385_ (
  .A({ S4798 }),
  .Y({ S4799 })
);
NAND #() 
NAND_3016_ (
  .A({ S4662 }),
  .B({ S4665 }),
  .Y({ S4800 })
);
NAND #() 
NAND_3017_ (
  .A({ S4668 }),
  .B({ S4800 }),
  .Y({ S4801 })
);
NAND #() 
NAND_3018_ (
  .A({ S4708 }),
  .B({ S4801 }),
  .Y({ S4802 })
);
NOT #() 
NOT_386_ (
  .A({ S4802 }),
  .Y({ S4803 })
);
NOR #() 
NOR_1508_ (
  .A({ S4798 }),
  .B({ S4803 }),
  .Y({ S4804 })
);
NAND #() 
NAND_3019_ (
  .A({ S4799 }),
  .B({ S4802 }),
  .Y({ S4805 })
);
NOR #() 
NOR_1509_ (
  .A({ S1952 }),
  .B({ S4805 }),
  .Y({ S4806 })
);
NAND #() 
NAND_3020_ (
  .A({ S1953 }),
  .B({ S4804 }),
  .Y({ S4807 })
);
NOR #() 
NOR_1510_ (
  .A({ S4654 }),
  .B({ S4658 }),
  .Y({ S4808 })
);
NOR #() 
NOR_1511_ (
  .A({ S4660 }),
  .B({ S4808 }),
  .Y({ S4809 })
);
NAND #() 
NAND_3021_ (
  .A({ S4708 }),
  .B({ S4809 }),
  .Y({ S4810 })
);
NOT #() 
NOT_387_ (
  .A({ S4810 }),
  .Y({ S4811 })
);
NOR #() 
NOR_1512_ (
  .A({ S4650 }),
  .B({ S4708 }),
  .Y({ S4812 })
);
NOT #() 
NOT_388_ (
  .A({ S4812 }),
  .Y({ S4813 })
);
NOR #() 
NOR_1513_ (
  .A({ S4811 }),
  .B({ S4812 }),
  .Y({ S4814 })
);
NAND #() 
NAND_3022_ (
  .A({ S4810 }),
  .B({ S4813 }),
  .Y({ S4815 })
);
NOR #() 
NOR_1514_ (
  .A({ S1848 }),
  .B({ S4814 }),
  .Y({ S4816 })
);
NAND #() 
NAND_3023_ (
  .A({ S1849 }),
  .B({ S4815 }),
  .Y({ S4817 })
);
NOR #() 
NOR_1515_ (
  .A({ S1849 }),
  .B({ S4815 }),
  .Y({ S4818 })
);
NAND #() 
NAND_3024_ (
  .A({ S1848 }),
  .B({ S4814 }),
  .Y({ S4819 })
);
NOR #() 
NOR_1516_ (
  .A({ S4816 }),
  .B({ S4818 }),
  .Y({ S4820 })
);
NAND #() 
NAND_3025_ (
  .A({ S4817 }),
  .B({ S4819 }),
  .Y({ S4821 })
);
NOR #() 
NOR_1517_ (
  .A({ S1516 }),
  .B({ S4709 }),
  .Y({ S4822 })
);
NAND #() 
NAND_3026_ (
  .A({ S1515 }),
  .B({ S4708 }),
  .Y({ S4823 })
);
NOR #() 
NOR_1518_ (
  .A({ S910 }),
  .B({ S4822 }),
  .Y({ S4824 })
);
NAND #() 
NAND_3027_ (
  .A({ datapath_addsubunit_in1_6 }),
  .B({ S4823 }),
  .Y({ S4825 })
);
NOR #() 
NOR_1519_ (
  .A({ datapath_addsubunit_in1_6 }),
  .B({ S4823 }),
  .Y({ S4826 })
);
NAND #() 
NAND_3028_ (
  .A({ S910 }),
  .B({ S4822 }),
  .Y({ S4827 })
);
NOR #() 
NOR_1520_ (
  .A({ S4824 }),
  .B({ S4826 }),
  .Y({ S4828 })
);
NAND #() 
NAND_3029_ (
  .A({ S4825 }),
  .B({ S4827 }),
  .Y({ S4829 })
);
NOR #() 
NOR_1521_ (
  .A({ S1745 }),
  .B({ S4828 }),
  .Y({ S4830 })
);
NAND #() 
NAND_3030_ (
  .A({ S1746 }),
  .B({ S4829 }),
  .Y({ S4831 })
);
NOR #() 
NOR_1522_ (
  .A({ S1746 }),
  .B({ S4829 }),
  .Y({ S4832 })
);
NAND #() 
NAND_3031_ (
  .A({ S1745 }),
  .B({ S4828 }),
  .Y({ S4833 })
);
NOR #() 
NOR_1523_ (
  .A({ S4830 }),
  .B({ S4832 }),
  .Y({ S4834 })
);
NAND #() 
NAND_3032_ (
  .A({ S4831 }),
  .B({ S4833 }),
  .Y({ S4835 })
);
NOR #() 
NOR_1524_ (
  .A({ datapath_addsubunit_in1_5 }),
  .B({ S1516 }),
  .Y({ S4836 })
);
NAND #() 
NAND_3033_ (
  .A({ S963 }),
  .B({ S1515 }),
  .Y({ S4837 })
);
NOR #() 
NOR_1525_ (
  .A({ S4835 }),
  .B({ S4836 }),
  .Y({ S4838 })
);
NAND #() 
NAND_3034_ (
  .A({ S4834 }),
  .B({ S4837 }),
  .Y({ S4839 })
);
NOR #() 
NOR_1526_ (
  .A({ S4830 }),
  .B({ S4838 }),
  .Y({ S4840 })
);
NAND #() 
NAND_3035_ (
  .A({ S4831 }),
  .B({ S4839 }),
  .Y({ S4841 })
);
NOR #() 
NOR_1527_ (
  .A({ S4821 }),
  .B({ S4840 }),
  .Y({ S4842 })
);
NAND #() 
NAND_3036_ (
  .A({ S4820 }),
  .B({ S4841 }),
  .Y({ S4843 })
);
NOR #() 
NOR_1528_ (
  .A({ S4816 }),
  .B({ S4842 }),
  .Y({ S4844 })
);
NAND #() 
NAND_3037_ (
  .A({ S4817 }),
  .B({ S4843 }),
  .Y({ S4845 })
);
NOR #() 
NOR_1529_ (
  .A({ S1953 }),
  .B({ S4804 }),
  .Y({ S4846 })
);
NAND #() 
NAND_3038_ (
  .A({ S1952 }),
  .B({ S4805 }),
  .Y({ S4847 })
);
NOR #() 
NOR_1530_ (
  .A({ S4806 }),
  .B({ S4846 }),
  .Y({ S4848 })
);
NAND #() 
NAND_3039_ (
  .A({ S4807 }),
  .B({ S4847 }),
  .Y({ S4849 })
);
NOR #() 
NOR_1531_ (
  .A({ S4844 }),
  .B({ S4849 }),
  .Y({ S4850 })
);
NAND #() 
NAND_3040_ (
  .A({ S4845 }),
  .B({ S4848 }),
  .Y({ S4851 })
);
NOR #() 
NOR_1532_ (
  .A({ S4806 }),
  .B({ S4850 }),
  .Y({ S4852 })
);
NAND #() 
NAND_3041_ (
  .A({ S4807 }),
  .B({ S4851 }),
  .Y({ S4853 })
);
NOR #() 
NOR_1533_ (
  .A({ S4797 }),
  .B({ S4852 }),
  .Y({ S4854 })
);
NAND #() 
NAND_3042_ (
  .A({ S4796 }),
  .B({ S4853 }),
  .Y({ S4855 })
);
NOR #() 
NOR_1534_ (
  .A({ S4792 }),
  .B({ S4854 }),
  .Y({ S4856 })
);
NAND #() 
NAND_3043_ (
  .A({ S4793 }),
  .B({ S4855 }),
  .Y({ S4857 })
);
NOR #() 
NOR_1535_ (
  .A({ S4780 }),
  .B({ S4856 }),
  .Y({ S4858 })
);
NAND #() 
NAND_3044_ (
  .A({ S4779 }),
  .B({ S4857 }),
  .Y({ S4859 })
);
NOR #() 
NOR_1536_ (
  .A({ S4775 }),
  .B({ S4858 }),
  .Y({ S4860 })
);
NAND #() 
NAND_3045_ (
  .A({ S4776 }),
  .B({ S4859 }),
  .Y({ S4861 })
);
NOR #() 
NOR_1537_ (
  .A({ S4766 }),
  .B({ S4860 }),
  .Y({ S4862 })
);
NAND #() 
NAND_3046_ (
  .A({ S4765 }),
  .B({ S4861 }),
  .Y({ S4863 })
);
NOR #() 
NOR_1538_ (
  .A({ S4761 }),
  .B({ S4862 }),
  .Y({ S4864 })
);
NAND #() 
NAND_3047_ (
  .A({ S4762 }),
  .B({ S4863 }),
  .Y({ S4865 })
);
NOR #() 
NOR_1539_ (
  .A({ S4752 }),
  .B({ S4864 }),
  .Y({ S4866 })
);
NAND #() 
NAND_3048_ (
  .A({ S4751 }),
  .B({ S4865 }),
  .Y({ S4867 })
);
NOR #() 
NOR_1540_ (
  .A({ S4747 }),
  .B({ S4866 }),
  .Y({ S4868 })
);
NAND #() 
NAND_3049_ (
  .A({ S4748 }),
  .B({ S4867 }),
  .Y({ S4869 })
);
NOR #() 
NOR_1541_ (
  .A({ S4737 }),
  .B({ S4868 }),
  .Y({ S4870 })
);
NAND #() 
NAND_3050_ (
  .A({ S4738 }),
  .B({ S4869 }),
  .Y({ S4871 })
);
NOR #() 
NOR_1542_ (
  .A({ S4735 }),
  .B({ S4870 }),
  .Y({ S4872 })
);
NAND #() 
NAND_3051_ (
  .A({ S4736 }),
  .B({ S4871 }),
  .Y({ S4873 })
);
NOR #() 
NOR_1543_ (
  .A({ S4723 }),
  .B({ S4872 }),
  .Y({ S4874 })
);
NAND #() 
NAND_3052_ (
  .A({ S4722 }),
  .B({ S4873 }),
  .Y({ S4875 })
);
NAND #() 
NAND_3053_ (
  .A({ S2517 }),
  .B({ S3908 }),
  .Y({ S4876 })
);
NOT #() 
NOT_389_ (
  .A({ S4876 }),
  .Y({ S4877 })
);
NOR #() 
NOR_1544_ (
  .A({ S4693 }),
  .B({ S4877 }),
  .Y({ S4878 })
);
NOR #() 
NOR_1545_ (
  .A({ S3910 }),
  .B({ S4694 }),
  .Y({ S4879 })
);
NOR #() 
NOR_1546_ (
  .A({ S4878 }),
  .B({ S4879 }),
  .Y({ S4880 })
);
NOR #() 
NOR_1547_ (
  .A({ S4700 }),
  .B({ S4880 }),
  .Y({ S4881 })
);
NOT #() 
NOT_390_ (
  .A({ S4881 }),
  .Y({ S4882 })
);
NOR #() 
NOR_1548_ (
  .A({ S2617 }),
  .B({ S4882 }),
  .Y({ S4883 })
);
NAND #() 
NAND_3054_ (
  .A({ S2618 }),
  .B({ S4881 }),
  .Y({ S4884 })
);
NOR #() 
NOR_1549_ (
  .A({ S4718 }),
  .B({ S4883 }),
  .Y({ S4885 })
);
NAND #() 
NAND_3055_ (
  .A({ S4719 }),
  .B({ S4884 }),
  .Y({ S4886 })
);
NOR #() 
NOR_1550_ (
  .A({ S4874 }),
  .B({ S4886 }),
  .Y({ S4887 })
);
NAND #() 
NAND_3056_ (
  .A({ S4875 }),
  .B({ S4885 }),
  .Y({ S4888 })
);
NOR #() 
NOR_1551_ (
  .A({ S2618 }),
  .B({ S4699 }),
  .Y({ S4889 })
);
NAND #() 
NAND_3057_ (
  .A({ S2617 }),
  .B({ S4700 }),
  .Y({ S4890 })
);
NOR #() 
NOR_1552_ (
  .A({ S3907 }),
  .B({ S4889 }),
  .Y({ S4891 })
);
NAND #() 
NAND_3058_ (
  .A({ S3906 }),
  .B({ S4890 }),
  .Y({ S4892 })
);
NOR #() 
NOR_1553_ (
  .A({ S4883 }),
  .B({ S4889 }),
  .Y({ S4893 })
);
NAND #() 
NAND_3059_ (
  .A({ S4884 }),
  .B({ S4890 }),
  .Y({ S4894 })
);
NOR #() 
NOR_1554_ (
  .A({ S4887 }),
  .B({ S4892 }),
  .Y({ S4895 })
);
NAND #() 
NAND_3060_ (
  .A({ S4888 }),
  .B({ S4891 }),
  .Y({ S4896 })
);
NOR #() 
NOR_1555_ (
  .A({ S4722 }),
  .B({ S4873 }),
  .Y({ S4897 })
);
NAND #() 
NAND_3061_ (
  .A({ S4723 }),
  .B({ S4872 }),
  .Y({ S4898 })
);
NOR #() 
NOR_1556_ (
  .A({ S4874 }),
  .B({ S4897 }),
  .Y({ S4899 })
);
NAND #() 
NAND_3062_ (
  .A({ S4875 }),
  .B({ S4898 }),
  .Y({ S4900 })
);
NOR #() 
NOR_1557_ (
  .A({ S4896 }),
  .B({ S4899 }),
  .Y({ S4901 })
);
NAND #() 
NAND_3063_ (
  .A({ S4895 }),
  .B({ S4900 }),
  .Y({ S4902 })
);
NOR #() 
NOR_1558_ (
  .A({ S4716 }),
  .B({ S4895 }),
  .Y({ S4903 })
);
NAND #() 
NAND_3064_ (
  .A({ S4717 }),
  .B({ S4896 }),
  .Y({ S4904 })
);
NOR #() 
NOR_1559_ (
  .A({ S4901 }),
  .B({ S4903 }),
  .Y({ S4905 })
);
NAND #() 
NAND_3065_ (
  .A({ S4902 }),
  .B({ S4904 }),
  .Y({ S4906 })
);
NOR #() 
NOR_1560_ (
  .A({ S2617 }),
  .B({ S4906 }),
  .Y({ S4907 })
);
NAND #() 
NAND_3066_ (
  .A({ S2618 }),
  .B({ S4905 }),
  .Y({ S4908 })
);
NOR #() 
NOR_1561_ (
  .A({ S2618 }),
  .B({ S4905 }),
  .Y({ S4909 })
);
NAND #() 
NAND_3067_ (
  .A({ S2617 }),
  .B({ S4906 }),
  .Y({ S4910 })
);
NOR #() 
NOR_1562_ (
  .A({ S4907 }),
  .B({ S4909 }),
  .Y({ S4911 })
);
NAND #() 
NAND_3068_ (
  .A({ S4908 }),
  .B({ S4910 }),
  .Y({ S4912 })
);
NOR #() 
NOR_1563_ (
  .A({ S4735 }),
  .B({ S4737 }),
  .Y({ S4913 })
);
NAND #() 
NAND_3069_ (
  .A({ S4736 }),
  .B({ S4738 }),
  .Y({ S4914 })
);
NOR #() 
NOR_1564_ (
  .A({ S4869 }),
  .B({ S4913 }),
  .Y({ S4915 })
);
NAND #() 
NAND_3070_ (
  .A({ S4868 }),
  .B({ S4914 }),
  .Y({ S4916 })
);
NOR #() 
NOR_1565_ (
  .A({ S4868 }),
  .B({ S4914 }),
  .Y({ S4917 })
);
NAND #() 
NAND_3071_ (
  .A({ S4869 }),
  .B({ S4913 }),
  .Y({ S4918 })
);
NOR #() 
NOR_1566_ (
  .A({ S4915 }),
  .B({ S4917 }),
  .Y({ S4919 })
);
NAND #() 
NAND_3072_ (
  .A({ S4916 }),
  .B({ S4918 }),
  .Y({ S4920 })
);
NOR #() 
NOR_1567_ (
  .A({ S4896 }),
  .B({ S4919 }),
  .Y({ S4921 })
);
NAND #() 
NAND_3073_ (
  .A({ S4895 }),
  .B({ S4920 }),
  .Y({ S4922 })
);
NOR #() 
NOR_1568_ (
  .A({ S4733 }),
  .B({ S4895 }),
  .Y({ S4923 })
);
NAND #() 
NAND_3074_ (
  .A({ S4734 }),
  .B({ S4896 }),
  .Y({ S4924 })
);
NOR #() 
NOR_1569_ (
  .A({ S4921 }),
  .B({ S4923 }),
  .Y({ S4925 })
);
NAND #() 
NAND_3075_ (
  .A({ S4922 }),
  .B({ S4924 }),
  .Y({ S4926 })
);
NOR #() 
NOR_1570_ (
  .A({ S2518 }),
  .B({ S4925 }),
  .Y({ S4927 })
);
NAND #() 
NAND_3076_ (
  .A({ S2517 }),
  .B({ S4926 }),
  .Y({ S4928 })
);
NOR #() 
NOR_1571_ (
  .A({ S2517 }),
  .B({ S4926 }),
  .Y({ S4929 })
);
NAND #() 
NAND_3077_ (
  .A({ S2518 }),
  .B({ S4925 }),
  .Y({ S4930 })
);
NOR #() 
NOR_1572_ (
  .A({ S4751 }),
  .B({ S4865 }),
  .Y({ S4931 })
);
NAND #() 
NAND_3078_ (
  .A({ S4752 }),
  .B({ S4864 }),
  .Y({ S4932 })
);
NOR #() 
NOR_1573_ (
  .A({ S4866 }),
  .B({ S4931 }),
  .Y({ S4933 })
);
NAND #() 
NAND_3079_ (
  .A({ S4867 }),
  .B({ S4932 }),
  .Y({ S4934 })
);
NOR #() 
NOR_1574_ (
  .A({ S4896 }),
  .B({ S4933 }),
  .Y({ S4935 })
);
NAND #() 
NAND_3080_ (
  .A({ S4895 }),
  .B({ S4934 }),
  .Y({ S4936 })
);
NOR #() 
NOR_1575_ (
  .A({ S4745 }),
  .B({ S4895 }),
  .Y({ S4937 })
);
NAND #() 
NAND_3081_ (
  .A({ S4746 }),
  .B({ S4896 }),
  .Y({ S4938 })
);
NOR #() 
NOR_1576_ (
  .A({ S4935 }),
  .B({ S4937 }),
  .Y({ S4939 })
);
NAND #() 
NAND_3082_ (
  .A({ S4936 }),
  .B({ S4938 }),
  .Y({ S4940 })
);
NOR #() 
NOR_1577_ (
  .A({ S2417 }),
  .B({ S4940 }),
  .Y({ S4941 })
);
NAND #() 
NAND_3083_ (
  .A({ S2418 }),
  .B({ S4939 }),
  .Y({ S4942 })
);
NOR #() 
NOR_1578_ (
  .A({ S2418 }),
  .B({ S4939 }),
  .Y({ S4943 })
);
NAND #() 
NAND_3084_ (
  .A({ S2417 }),
  .B({ S4940 }),
  .Y({ S4944 })
);
NOR #() 
NOR_1579_ (
  .A({ S4941 }),
  .B({ S4943 }),
  .Y({ S4945 })
);
NAND #() 
NAND_3085_ (
  .A({ S4942 }),
  .B({ S4944 }),
  .Y({ S4946 })
);
NOR #() 
NOR_1580_ (
  .A({ S4765 }),
  .B({ S4861 }),
  .Y({ S4947 })
);
NAND #() 
NAND_3086_ (
  .A({ S4766 }),
  .B({ S4860 }),
  .Y({ S4948 })
);
NOR #() 
NOR_1581_ (
  .A({ S4862 }),
  .B({ S4947 }),
  .Y({ S4949 })
);
NAND #() 
NAND_3087_ (
  .A({ S4863 }),
  .B({ S4948 }),
  .Y({ S4950 })
);
NOR #() 
NOR_1582_ (
  .A({ S4896 }),
  .B({ S4949 }),
  .Y({ S4951 })
);
NAND #() 
NAND_3088_ (
  .A({ S4895 }),
  .B({ S4950 }),
  .Y({ S4952 })
);
NOR #() 
NOR_1583_ (
  .A({ S4759 }),
  .B({ S4895 }),
  .Y({ S4953 })
);
NAND #() 
NAND_3089_ (
  .A({ S4760 }),
  .B({ S4896 }),
  .Y({ S4954 })
);
NOR #() 
NOR_1584_ (
  .A({ S4951 }),
  .B({ S4953 }),
  .Y({ S4955 })
);
NAND #() 
NAND_3090_ (
  .A({ S4952 }),
  .B({ S4954 }),
  .Y({ S4956 })
);
NOR #() 
NOR_1585_ (
  .A({ S2311 }),
  .B({ S4956 }),
  .Y({ S4957 })
);
NAND #() 
NAND_3091_ (
  .A({ S2312 }),
  .B({ S4955 }),
  .Y({ S4958 })
);
NOR #() 
NOR_1586_ (
  .A({ S2312 }),
  .B({ S4955 }),
  .Y({ S4959 })
);
NAND #() 
NAND_3092_ (
  .A({ S2311 }),
  .B({ S4956 }),
  .Y({ S4960 })
);
NOR #() 
NOR_1587_ (
  .A({ S4773 }),
  .B({ S4895 }),
  .Y({ S4961 })
);
NAND #() 
NAND_3093_ (
  .A({ S4774 }),
  .B({ S4896 }),
  .Y({ S4962 })
);
NOR #() 
NOR_1588_ (
  .A({ S4779 }),
  .B({ S4857 }),
  .Y({ S4963 })
);
NAND #() 
NAND_3094_ (
  .A({ S4780 }),
  .B({ S4856 }),
  .Y({ S4964 })
);
NOR #() 
NOR_1589_ (
  .A({ S4858 }),
  .B({ S4963 }),
  .Y({ S4965 })
);
NAND #() 
NAND_3095_ (
  .A({ S4859 }),
  .B({ S4964 }),
  .Y({ S4966 })
);
NOR #() 
NOR_1590_ (
  .A({ S4896 }),
  .B({ S4965 }),
  .Y({ S4967 })
);
NAND #() 
NAND_3096_ (
  .A({ S4895 }),
  .B({ S4966 }),
  .Y({ S4968 })
);
NOR #() 
NOR_1591_ (
  .A({ S4961 }),
  .B({ S4967 }),
  .Y({ S4969 })
);
NAND #() 
NAND_3097_ (
  .A({ S4962 }),
  .B({ S4968 }),
  .Y({ S4970 })
);
NOR #() 
NOR_1592_ (
  .A({ S2205 }),
  .B({ S4970 }),
  .Y({ S4971 })
);
NAND #() 
NAND_3098_ (
  .A({ S2206 }),
  .B({ S4969 }),
  .Y({ S4972 })
);
NOR #() 
NOR_1593_ (
  .A({ S2206 }),
  .B({ S4969 }),
  .Y({ S4973 })
);
NAND #() 
NAND_3099_ (
  .A({ S2205 }),
  .B({ S4970 }),
  .Y({ S4974 })
);
NOR #() 
NOR_1594_ (
  .A({ S4971 }),
  .B({ S4973 }),
  .Y({ S4975 })
);
NAND #() 
NAND_3100_ (
  .A({ S4972 }),
  .B({ S4974 }),
  .Y({ S4976 })
);
NOR #() 
NOR_1595_ (
  .A({ S4796 }),
  .B({ S4853 }),
  .Y({ S4977 })
);
NAND #() 
NAND_3101_ (
  .A({ S4797 }),
  .B({ S4852 }),
  .Y({ S4978 })
);
NOR #() 
NOR_1596_ (
  .A({ S4854 }),
  .B({ S4977 }),
  .Y({ S4979 })
);
NAND #() 
NAND_3102_ (
  .A({ S4855 }),
  .B({ S4978 }),
  .Y({ S4980 })
);
NOR #() 
NOR_1597_ (
  .A({ S4896 }),
  .B({ S4979 }),
  .Y({ S4981 })
);
NAND #() 
NAND_3103_ (
  .A({ S4895 }),
  .B({ S4980 }),
  .Y({ S4982 })
);
NOR #() 
NOR_1598_ (
  .A({ S4790 }),
  .B({ S4895 }),
  .Y({ S4983 })
);
NAND #() 
NAND_3104_ (
  .A({ S4791 }),
  .B({ S4896 }),
  .Y({ S4984 })
);
NOR #() 
NOR_1599_ (
  .A({ S4981 }),
  .B({ S4983 }),
  .Y({ S4985 })
);
NAND #() 
NAND_3105_ (
  .A({ S4982 }),
  .B({ S4984 }),
  .Y({ S4986 })
);
NOR #() 
NOR_1600_ (
  .A({ S2106 }),
  .B({ S4986 }),
  .Y({ S4987 })
);
NAND #() 
NAND_3106_ (
  .A({ S2107 }),
  .B({ S4985 }),
  .Y({ S4988 })
);
NOR #() 
NOR_1601_ (
  .A({ S2107 }),
  .B({ S4985 }),
  .Y({ S4989 })
);
NAND #() 
NAND_3107_ (
  .A({ S2106 }),
  .B({ S4986 }),
  .Y({ S4990 })
);
NOR #() 
NOR_1602_ (
  .A({ S4804 }),
  .B({ S4895 }),
  .Y({ S4991 })
);
NAND #() 
NAND_3108_ (
  .A({ S4805 }),
  .B({ S4896 }),
  .Y({ S4992 })
);
NOR #() 
NOR_1603_ (
  .A({ S4845 }),
  .B({ S4848 }),
  .Y({ S4993 })
);
NAND #() 
NAND_3109_ (
  .A({ S4844 }),
  .B({ S4849 }),
  .Y({ S4994 })
);
NOR #() 
NOR_1604_ (
  .A({ S4850 }),
  .B({ S4993 }),
  .Y({ S4995 })
);
NAND #() 
NAND_3110_ (
  .A({ S4851 }),
  .B({ S4994 }),
  .Y({ S4996 })
);
NOR #() 
NOR_1605_ (
  .A({ S4896 }),
  .B({ S4995 }),
  .Y({ S4997 })
);
NAND #() 
NAND_3111_ (
  .A({ S4895 }),
  .B({ S4996 }),
  .Y({ S4998 })
);
NOR #() 
NOR_1606_ (
  .A({ S4991 }),
  .B({ S4997 }),
  .Y({ S4999 })
);
NAND #() 
NAND_3112_ (
  .A({ S4992 }),
  .B({ S4998 }),
  .Y({ S5000 })
);
NOR #() 
NOR_1607_ (
  .A({ S1597 }),
  .B({ S5000 }),
  .Y({ S5001 })
);
NAND #() 
NAND_3113_ (
  .A({ S1598 }),
  .B({ S4999 }),
  .Y({ S5002 })
);
NOR #() 
NOR_1608_ (
  .A({ S4815 }),
  .B({ S4895 }),
  .Y({ S5003 })
);
NAND #() 
NAND_3114_ (
  .A({ S4814 }),
  .B({ S4896 }),
  .Y({ S5004 })
);
NOR #() 
NOR_1609_ (
  .A({ S4820 }),
  .B({ S4841 }),
  .Y({ S5005 })
);
NAND #() 
NAND_3115_ (
  .A({ S4821 }),
  .B({ S4840 }),
  .Y({ S5006 })
);
NOR #() 
NOR_1610_ (
  .A({ S4842 }),
  .B({ S5005 }),
  .Y({ S5007 })
);
NAND #() 
NAND_3116_ (
  .A({ S4843 }),
  .B({ S5006 }),
  .Y({ S5008 })
);
NOR #() 
NOR_1611_ (
  .A({ S4896 }),
  .B({ S5007 }),
  .Y({ S5009 })
);
NAND #() 
NAND_3117_ (
  .A({ S4895 }),
  .B({ S5008 }),
  .Y({ S5010 })
);
NOR #() 
NOR_1612_ (
  .A({ S5003 }),
  .B({ S5009 }),
  .Y({ S5011 })
);
NAND #() 
NAND_3118_ (
  .A({ S5004 }),
  .B({ S5010 }),
  .Y({ S5012 })
);
NOR #() 
NOR_1613_ (
  .A({ S1952 }),
  .B({ S5012 }),
  .Y({ S5013 })
);
NAND #() 
NAND_3119_ (
  .A({ S1953 }),
  .B({ S5011 }),
  .Y({ S5014 })
);
NOR #() 
NOR_1614_ (
  .A({ S1953 }),
  .B({ S5011 }),
  .Y({ S5015 })
);
NAND #() 
NAND_3120_ (
  .A({ S1952 }),
  .B({ S5012 }),
  .Y({ S5016 })
);
NOR #() 
NOR_1615_ (
  .A({ S5013 }),
  .B({ S5015 }),
  .Y({ S5017 })
);
NAND #() 
NAND_3121_ (
  .A({ S5014 }),
  .B({ S5016 }),
  .Y({ S5018 })
);
NOR #() 
NOR_1616_ (
  .A({ S4834 }),
  .B({ S4837 }),
  .Y({ S5019 })
);
NAND #() 
NAND_3122_ (
  .A({ S4835 }),
  .B({ S4836 }),
  .Y({ S5020 })
);
NOR #() 
NOR_1617_ (
  .A({ S4838 }),
  .B({ S5019 }),
  .Y({ S5021 })
);
NAND #() 
NAND_3123_ (
  .A({ S4839 }),
  .B({ S5020 }),
  .Y({ S5022 })
);
NOR #() 
NOR_1618_ (
  .A({ S4896 }),
  .B({ S5021 }),
  .Y({ S5023 })
);
NAND #() 
NAND_3124_ (
  .A({ S4895 }),
  .B({ S5022 }),
  .Y({ S5024 })
);
NOR #() 
NOR_1619_ (
  .A({ S4829 }),
  .B({ S4895 }),
  .Y({ S5025 })
);
NAND #() 
NAND_3125_ (
  .A({ S4828 }),
  .B({ S4896 }),
  .Y({ S5026 })
);
NOR #() 
NOR_1620_ (
  .A({ S5023 }),
  .B({ S5025 }),
  .Y({ S5027 })
);
NAND #() 
NAND_3126_ (
  .A({ S5024 }),
  .B({ S5026 }),
  .Y({ S5028 })
);
NOR #() 
NOR_1621_ (
  .A({ S1848 }),
  .B({ S5028 }),
  .Y({ S5029 })
);
NAND #() 
NAND_3127_ (
  .A({ S1849 }),
  .B({ S5027 }),
  .Y({ S5030 })
);
NOR #() 
NOR_1622_ (
  .A({ S1849 }),
  .B({ S5027 }),
  .Y({ S5031 })
);
NAND #() 
NAND_3128_ (
  .A({ S1848 }),
  .B({ S5028 }),
  .Y({ S5032 })
);
NOR #() 
NOR_1623_ (
  .A({ S5029 }),
  .B({ S5031 }),
  .Y({ S5033 })
);
NAND #() 
NAND_3129_ (
  .A({ S5030 }),
  .B({ S5032 }),
  .Y({ S5034 })
);
NOR #() 
NOR_1624_ (
  .A({ S1516 }),
  .B({ S4896 }),
  .Y({ S5035 })
);
NAND #() 
NAND_3130_ (
  .A({ S1515 }),
  .B({ S4895 }),
  .Y({ S5036 })
);
NOR #() 
NOR_1625_ (
  .A({ S963 }),
  .B({ S5035 }),
  .Y({ S5037 })
);
NAND #() 
NAND_3131_ (
  .A({ datapath_addsubunit_in1_5 }),
  .B({ S5036 }),
  .Y({ S5038 })
);
NOR #() 
NOR_1626_ (
  .A({ datapath_addsubunit_in1_5 }),
  .B({ S5036 }),
  .Y({ S5039 })
);
NAND #() 
NAND_3132_ (
  .A({ S963 }),
  .B({ S5035 }),
  .Y({ S5040 })
);
NOR #() 
NOR_1627_ (
  .A({ S5037 }),
  .B({ S5039 }),
  .Y({ S5041 })
);
NAND #() 
NAND_3133_ (
  .A({ S5038 }),
  .B({ S5040 }),
  .Y({ S5042 })
);
NOR #() 
NOR_1628_ (
  .A({ S1745 }),
  .B({ S5041 }),
  .Y({ S5043 })
);
NAND #() 
NAND_3134_ (
  .A({ S1746 }),
  .B({ S5042 }),
  .Y({ S5044 })
);
NOR #() 
NOR_1629_ (
  .A({ datapath_addsubunit_in1_4 }),
  .B({ S1516 }),
  .Y({ S5045 })
);
NAND #() 
NAND_3135_ (
  .A({ S1013 }),
  .B({ S1515 }),
  .Y({ S5046 })
);
NOR #() 
NOR_1630_ (
  .A({ S1746 }),
  .B({ S5042 }),
  .Y({ S5047 })
);
NAND #() 
NAND_3136_ (
  .A({ S1745 }),
  .B({ S5041 }),
  .Y({ S5048 })
);
NOR #() 
NOR_1631_ (
  .A({ S5043 }),
  .B({ S5047 }),
  .Y({ S5049 })
);
NAND #() 
NAND_3137_ (
  .A({ S5044 }),
  .B({ S5048 }),
  .Y({ S5050 })
);
NOR #() 
NOR_1632_ (
  .A({ S5045 }),
  .B({ S5050 }),
  .Y({ S5051 })
);
NAND #() 
NAND_3138_ (
  .A({ S5046 }),
  .B({ S5049 }),
  .Y({ S5052 })
);
NOR #() 
NOR_1633_ (
  .A({ S5043 }),
  .B({ S5051 }),
  .Y({ S5053 })
);
NAND #() 
NAND_3139_ (
  .A({ S5044 }),
  .B({ S5052 }),
  .Y({ S5054 })
);
NOR #() 
NOR_1634_ (
  .A({ S5034 }),
  .B({ S5053 }),
  .Y({ S5055 })
);
NAND #() 
NAND_3140_ (
  .A({ S5033 }),
  .B({ S5054 }),
  .Y({ S5056 })
);
NOR #() 
NOR_1635_ (
  .A({ S5029 }),
  .B({ S5055 }),
  .Y({ S5057 })
);
NAND #() 
NAND_3141_ (
  .A({ S5030 }),
  .B({ S5056 }),
  .Y({ S5058 })
);
NOR #() 
NOR_1636_ (
  .A({ S5018 }),
  .B({ S5057 }),
  .Y({ S5059 })
);
NAND #() 
NAND_3142_ (
  .A({ S5017 }),
  .B({ S5058 }),
  .Y({ S5060 })
);
NOR #() 
NOR_1637_ (
  .A({ S5013 }),
  .B({ S5059 }),
  .Y({ S5061 })
);
NAND #() 
NAND_3143_ (
  .A({ S5014 }),
  .B({ S5060 }),
  .Y({ S5062 })
);
NOR #() 
NOR_1638_ (
  .A({ S1598 }),
  .B({ S4999 }),
  .Y({ S5063 })
);
NAND #() 
NAND_3144_ (
  .A({ S1597 }),
  .B({ S5000 }),
  .Y({ S5064 })
);
NOR #() 
NOR_1639_ (
  .A({ S5001 }),
  .B({ S5063 }),
  .Y({ S5065 })
);
NAND #() 
NAND_3145_ (
  .A({ S5002 }),
  .B({ S5064 }),
  .Y({ S5066 })
);
NOR #() 
NOR_1640_ (
  .A({ S5061 }),
  .B({ S5066 }),
  .Y({ S5067 })
);
NAND #() 
NAND_3146_ (
  .A({ S5062 }),
  .B({ S5065 }),
  .Y({ S5068 })
);
NOR #() 
NOR_1641_ (
  .A({ S5001 }),
  .B({ S5067 }),
  .Y({ S5069 })
);
NAND #() 
NAND_3147_ (
  .A({ S5002 }),
  .B({ S5068 }),
  .Y({ S5070 })
);
NOR #() 
NOR_1642_ (
  .A({ S4989 }),
  .B({ S5069 }),
  .Y({ S5071 })
);
NAND #() 
NAND_3148_ (
  .A({ S4990 }),
  .B({ S5070 }),
  .Y({ S5072 })
);
NOR #() 
NOR_1643_ (
  .A({ S4987 }),
  .B({ S5071 }),
  .Y({ S5073 })
);
NAND #() 
NAND_3149_ (
  .A({ S4988 }),
  .B({ S5072 }),
  .Y({ S5074 })
);
NOR #() 
NOR_1644_ (
  .A({ S4976 }),
  .B({ S5073 }),
  .Y({ S5075 })
);
NAND #() 
NAND_3150_ (
  .A({ S4975 }),
  .B({ S5074 }),
  .Y({ S5076 })
);
NOR #() 
NOR_1645_ (
  .A({ S4971 }),
  .B({ S5075 }),
  .Y({ S5077 })
);
NAND #() 
NAND_3151_ (
  .A({ S4972 }),
  .B({ S5076 }),
  .Y({ S5078 })
);
NOR #() 
NOR_1646_ (
  .A({ S4959 }),
  .B({ S5077 }),
  .Y({ S5079 })
);
NAND #() 
NAND_3152_ (
  .A({ S4960 }),
  .B({ S5078 }),
  .Y({ S5080 })
);
NOR #() 
NOR_1647_ (
  .A({ S4957 }),
  .B({ S5079 }),
  .Y({ S5081 })
);
NAND #() 
NAND_3153_ (
  .A({ S4958 }),
  .B({ S5080 }),
  .Y({ S5082 })
);
NOR #() 
NOR_1648_ (
  .A({ S4946 }),
  .B({ S5081 }),
  .Y({ S5083 })
);
NAND #() 
NAND_3154_ (
  .A({ S4945 }),
  .B({ S5082 }),
  .Y({ S5084 })
);
NOR #() 
NOR_1649_ (
  .A({ S4941 }),
  .B({ S5083 }),
  .Y({ S5085 })
);
NAND #() 
NAND_3155_ (
  .A({ S4942 }),
  .B({ S5084 }),
  .Y({ S5086 })
);
NOR #() 
NOR_1650_ (
  .A({ S4929 }),
  .B({ S5086 }),
  .Y({ S5087 })
);
NAND #() 
NAND_3156_ (
  .A({ S4930 }),
  .B({ S5085 }),
  .Y({ S5088 })
);
NOR #() 
NOR_1651_ (
  .A({ S4927 }),
  .B({ S5087 }),
  .Y({ S5089 })
);
NAND #() 
NAND_3157_ (
  .A({ S4928 }),
  .B({ S5088 }),
  .Y({ S5090 })
);
NOR #() 
NOR_1652_ (
  .A({ S4912 }),
  .B({ S5090 }),
  .Y({ S5091 })
);
NAND #() 
NAND_3158_ (
  .A({ S4911 }),
  .B({ S5089 }),
  .Y({ S5092 })
);
NOR #() 
NOR_1653_ (
  .A({ S4881 }),
  .B({ S4895 }),
  .Y({ S5093 })
);
NOR #() 
NOR_1654_ (
  .A({ S4718 }),
  .B({ S4874 }),
  .Y({ S5094 })
);
NAND #() 
NAND_3159_ (
  .A({ S4719 }),
  .B({ S4875 }),
  .Y({ S5095 })
);
NOR #() 
NOR_1655_ (
  .A({ S4894 }),
  .B({ S5094 }),
  .Y({ S5096 })
);
NOR #() 
NOR_1656_ (
  .A({ S4893 }),
  .B({ S5095 }),
  .Y({ S5097 })
);
NOR #() 
NOR_1657_ (
  .A({ S5096 }),
  .B({ S5097 }),
  .Y({ S5098 })
);
NOR #() 
NOR_1658_ (
  .A({ S4896 }),
  .B({ S5098 }),
  .Y({ S5099 })
);
NOR #() 
NOR_1659_ (
  .A({ S5093 }),
  .B({ S5099 }),
  .Y({ S5100 })
);
NOT #() 
NOT_391_ (
  .A({ S5100 }),
  .Y({ S5101 })
);
NOR #() 
NOR_1660_ (
  .A({ S2717 }),
  .B({ S5101 }),
  .Y({ S5102 })
);
NAND #() 
NAND_3160_ (
  .A({ S2718 }),
  .B({ S5100 }),
  .Y({ S5103 })
);
NOR #() 
NOR_1661_ (
  .A({ S4907 }),
  .B({ S5102 }),
  .Y({ S5104 })
);
NAND #() 
NAND_3161_ (
  .A({ S4908 }),
  .B({ S5103 }),
  .Y({ S5105 })
);
NOR #() 
NOR_1662_ (
  .A({ S5091 }),
  .B({ S5105 }),
  .Y({ S5106 })
);
NAND #() 
NAND_3162_ (
  .A({ S5092 }),
  .B({ S5104 }),
  .Y({ S5107 })
);
NOR #() 
NOR_1663_ (
  .A({ S2718 }),
  .B({ S5100 }),
  .Y({ S5108 })
);
NAND #() 
NAND_3163_ (
  .A({ S2717 }),
  .B({ S5101 }),
  .Y({ S5109 })
);
NOR #() 
NOR_1664_ (
  .A({ S3905 }),
  .B({ S5108 }),
  .Y({ S5110 })
);
NAND #() 
NAND_3164_ (
  .A({ S3904 }),
  .B({ S5109 }),
  .Y({ S5111 })
);
NOR #() 
NOR_1665_ (
  .A({ S5106 }),
  .B({ S5111 }),
  .Y({ S5112 })
);
NAND #() 
NAND_3165_ (
  .A({ S5107 }),
  .B({ S5110 }),
  .Y({ S5113 })
);
NOR #() 
NOR_1666_ (
  .A({ S5102 }),
  .B({ S5108 }),
  .Y({ S5114 })
);
NAND #() 
NAND_3166_ (
  .A({ S5103 }),
  .B({ S5109 }),
  .Y({ S5115 })
);
NOR #() 
NOR_1667_ (
  .A({ S4907 }),
  .B({ S5091 }),
  .Y({ S5116 })
);
NAND #() 
NAND_3167_ (
  .A({ S4908 }),
  .B({ S5092 }),
  .Y({ S5117 })
);
NOR #() 
NOR_1668_ (
  .A({ S5114 }),
  .B({ S5117 }),
  .Y({ S5118 })
);
NOR #() 
NOR_1669_ (
  .A({ S5115 }),
  .B({ S5116 }),
  .Y({ S5119 })
);
NOR #() 
NOR_1670_ (
  .A({ S5118 }),
  .B({ S5119 }),
  .Y({ S5120 })
);
NAND #() 
NAND_3168_ (
  .A({ S5112 }),
  .B({ S5120 }),
  .Y({ S5121 })
);
NAND #() 
NAND_3169_ (
  .A({ S5100 }),
  .B({ S5113 }),
  .Y({ S5122 })
);
NAND #() 
NAND_3170_ (
  .A({ S5121 }),
  .B({ S5122 }),
  .Y({ S5123 })
);
NOR #() 
NOR_1671_ (
  .A({ S4911 }),
  .B({ S5089 }),
  .Y({ S5124 })
);
NAND #() 
NAND_3171_ (
  .A({ S4912 }),
  .B({ S5090 }),
  .Y({ S5125 })
);
NOR #() 
NOR_1672_ (
  .A({ S5091 }),
  .B({ S5124 }),
  .Y({ S5126 })
);
NAND #() 
NAND_3172_ (
  .A({ S5092 }),
  .B({ S5125 }),
  .Y({ S5127 })
);
NOR #() 
NOR_1673_ (
  .A({ S5113 }),
  .B({ S5126 }),
  .Y({ S5128 })
);
NAND #() 
NAND_3173_ (
  .A({ S5112 }),
  .B({ S5127 }),
  .Y({ S5129 })
);
NOR #() 
NOR_1674_ (
  .A({ S4905 }),
  .B({ S5112 }),
  .Y({ S5130 })
);
NAND #() 
NAND_3174_ (
  .A({ S4906 }),
  .B({ S5113 }),
  .Y({ S5131 })
);
NOR #() 
NOR_1675_ (
  .A({ S5128 }),
  .B({ S5130 }),
  .Y({ S5132 })
);
NAND #() 
NAND_3175_ (
  .A({ S5129 }),
  .B({ S5131 }),
  .Y({ S5133 })
);
NOR #() 
NOR_1676_ (
  .A({ S2717 }),
  .B({ S5133 }),
  .Y({ S5134 })
);
NAND #() 
NAND_3176_ (
  .A({ S2718 }),
  .B({ S5132 }),
  .Y({ S5135 })
);
NAND #() 
NAND_3177_ (
  .A({ S2717 }),
  .B({ S5133 }),
  .Y({ S5136 })
);
NAND #() 
NAND_3178_ (
  .A({ S5135 }),
  .B({ S5136 }),
  .Y({ S5137 })
);
NOT #() 
NOT_392_ (
  .A({ S5137 }),
  .Y({ S5138 })
);
NOR #() 
NOR_1677_ (
  .A({ S4927 }),
  .B({ S4929 }),
  .Y({ S5139 })
);
NAND #() 
NAND_3179_ (
  .A({ S4928 }),
  .B({ S4930 }),
  .Y({ S5140 })
);
NOR #() 
NOR_1678_ (
  .A({ S5086 }),
  .B({ S5139 }),
  .Y({ S5141 })
);
NOR #() 
NOR_1679_ (
  .A({ S5085 }),
  .B({ S5140 }),
  .Y({ S5142 })
);
NOR #() 
NOR_1680_ (
  .A({ S5141 }),
  .B({ S5142 }),
  .Y({ S5143 })
);
NOR #() 
NOR_1681_ (
  .A({ S5113 }),
  .B({ S5143 }),
  .Y({ S5144 })
);
NOR #() 
NOR_1682_ (
  .A({ S4925 }),
  .B({ S5112 }),
  .Y({ S5145 })
);
NOR #() 
NOR_1683_ (
  .A({ S5144 }),
  .B({ S5145 }),
  .Y({ S5146 })
);
NOT #() 
NOT_393_ (
  .A({ S5146 }),
  .Y({ S5147 })
);
NAND #() 
NAND_3180_ (
  .A({ S2617 }),
  .B({ S5147 }),
  .Y({ S5148 })
);
NAND #() 
NAND_3181_ (
  .A({ S2618 }),
  .B({ S5146 }),
  .Y({ S5149 })
);
NOR #() 
NOR_1684_ (
  .A({ S4945 }),
  .B({ S5082 }),
  .Y({ S5150 })
);
NOR #() 
NOR_1685_ (
  .A({ S5083 }),
  .B({ S5150 }),
  .Y({ S5151 })
);
NOR #() 
NOR_1686_ (
  .A({ S5113 }),
  .B({ S5151 }),
  .Y({ S5152 })
);
NOR #() 
NOR_1687_ (
  .A({ S4939 }),
  .B({ S5112 }),
  .Y({ S5153 })
);
NOR #() 
NOR_1688_ (
  .A({ S5152 }),
  .B({ S5153 }),
  .Y({ S5154 })
);
NOT #() 
NOT_394_ (
  .A({ S5154 }),
  .Y({ S5155 })
);
NOR #() 
NOR_1689_ (
  .A({ S2517 }),
  .B({ S5155 }),
  .Y({ S5156 })
);
NAND #() 
NAND_3182_ (
  .A({ S2518 }),
  .B({ S5154 }),
  .Y({ S5157 })
);
NOR #() 
NOR_1690_ (
  .A({ S2518 }),
  .B({ S5154 }),
  .Y({ S5158 })
);
NOR #() 
NOR_1691_ (
  .A({ S5156 }),
  .B({ S5158 }),
  .Y({ S5159 })
);
NOT #() 
NOT_395_ (
  .A({ S5159 }),
  .Y({ S5160 })
);
NOR #() 
NOR_1692_ (
  .A({ S4957 }),
  .B({ S4959 }),
  .Y({ S5161 })
);
NAND #() 
NAND_3183_ (
  .A({ S4958 }),
  .B({ S4960 }),
  .Y({ S5162 })
);
NOR #() 
NOR_1693_ (
  .A({ S5077 }),
  .B({ S5161 }),
  .Y({ S5163 })
);
NAND #() 
NAND_3184_ (
  .A({ S5078 }),
  .B({ S5162 }),
  .Y({ S5164 })
);
NOR #() 
NOR_1694_ (
  .A({ S5078 }),
  .B({ S5162 }),
  .Y({ S5165 })
);
NAND #() 
NAND_3185_ (
  .A({ S5077 }),
  .B({ S5161 }),
  .Y({ S5166 })
);
NOR #() 
NOR_1695_ (
  .A({ S5163 }),
  .B({ S5165 }),
  .Y({ S5167 })
);
NAND #() 
NAND_3186_ (
  .A({ S5164 }),
  .B({ S5166 }),
  .Y({ S5168 })
);
NOR #() 
NOR_1696_ (
  .A({ S5113 }),
  .B({ S5168 }),
  .Y({ S5169 })
);
NAND #() 
NAND_3187_ (
  .A({ S5112 }),
  .B({ S5167 }),
  .Y({ S5170 })
);
NOR #() 
NOR_1697_ (
  .A({ S4955 }),
  .B({ S5112 }),
  .Y({ S5171 })
);
NAND #() 
NAND_3188_ (
  .A({ S4956 }),
  .B({ S5113 }),
  .Y({ S5172 })
);
NOR #() 
NOR_1698_ (
  .A({ S5169 }),
  .B({ S5171 }),
  .Y({ S5173 })
);
NAND #() 
NAND_3189_ (
  .A({ S5170 }),
  .B({ S5172 }),
  .Y({ S5174 })
);
NOR #() 
NOR_1699_ (
  .A({ S2417 }),
  .B({ S5174 }),
  .Y({ S5175 })
);
NAND #() 
NAND_3190_ (
  .A({ S2418 }),
  .B({ S5173 }),
  .Y({ S5176 })
);
NOR #() 
NOR_1700_ (
  .A({ S2418 }),
  .B({ S5173 }),
  .Y({ S5177 })
);
NAND #() 
NAND_3191_ (
  .A({ S2417 }),
  .B({ S5174 }),
  .Y({ S5178 })
);
NOR #() 
NOR_1701_ (
  .A({ S4975 }),
  .B({ S5074 }),
  .Y({ S5179 })
);
NAND #() 
NAND_3192_ (
  .A({ S4976 }),
  .B({ S5073 }),
  .Y({ S5180 })
);
NOR #() 
NOR_1702_ (
  .A({ S5075 }),
  .B({ S5179 }),
  .Y({ S5181 })
);
NAND #() 
NAND_3193_ (
  .A({ S5076 }),
  .B({ S5180 }),
  .Y({ S5182 })
);
NOR #() 
NOR_1703_ (
  .A({ S5113 }),
  .B({ S5181 }),
  .Y({ S5183 })
);
NAND #() 
NAND_3194_ (
  .A({ S5112 }),
  .B({ S5182 }),
  .Y({ S5184 })
);
NOR #() 
NOR_1704_ (
  .A({ S4969 }),
  .B({ S5112 }),
  .Y({ S5185 })
);
NAND #() 
NAND_3195_ (
  .A({ S4970 }),
  .B({ S5113 }),
  .Y({ S5186 })
);
NOR #() 
NOR_1705_ (
  .A({ S5183 }),
  .B({ S5185 }),
  .Y({ S5187 })
);
NAND #() 
NAND_3196_ (
  .A({ S5184 }),
  .B({ S5186 }),
  .Y({ S5188 })
);
NOR #() 
NOR_1706_ (
  .A({ S2311 }),
  .B({ S5188 }),
  .Y({ S5189 })
);
NAND #() 
NAND_3197_ (
  .A({ S2312 }),
  .B({ S5187 }),
  .Y({ S5190 })
);
NOR #() 
NOR_1707_ (
  .A({ S2312 }),
  .B({ S5187 }),
  .Y({ S5191 })
);
NAND #() 
NAND_3198_ (
  .A({ S2311 }),
  .B({ S5188 }),
  .Y({ S5192 })
);
NOR #() 
NOR_1708_ (
  .A({ S5189 }),
  .B({ S5191 }),
  .Y({ S5193 })
);
NAND #() 
NAND_3199_ (
  .A({ S5190 }),
  .B({ S5192 }),
  .Y({ S5194 })
);
NOR #() 
NOR_1709_ (
  .A({ S4987 }),
  .B({ S4989 }),
  .Y({ S5195 })
);
NAND #() 
NAND_3200_ (
  .A({ S4988 }),
  .B({ S4990 }),
  .Y({ S5196 })
);
NOR #() 
NOR_1710_ (
  .A({ S5070 }),
  .B({ S5195 }),
  .Y({ S5197 })
);
NAND #() 
NAND_3201_ (
  .A({ S5069 }),
  .B({ S5196 }),
  .Y({ S5198 })
);
NOR #() 
NOR_1711_ (
  .A({ S5069 }),
  .B({ S5196 }),
  .Y({ S5199 })
);
NAND #() 
NAND_3202_ (
  .A({ S5070 }),
  .B({ S5195 }),
  .Y({ S5200 })
);
NOR #() 
NOR_1712_ (
  .A({ S5197 }),
  .B({ S5199 }),
  .Y({ S5201 })
);
NAND #() 
NAND_3203_ (
  .A({ S5198 }),
  .B({ S5200 }),
  .Y({ S5202 })
);
NOR #() 
NOR_1713_ (
  .A({ S5113 }),
  .B({ S5201 }),
  .Y({ S5203 })
);
NAND #() 
NAND_3204_ (
  .A({ S5112 }),
  .B({ S5202 }),
  .Y({ S5204 })
);
NOR #() 
NOR_1714_ (
  .A({ S4985 }),
  .B({ S5112 }),
  .Y({ S5205 })
);
NAND #() 
NAND_3205_ (
  .A({ S4986 }),
  .B({ S5113 }),
  .Y({ S5206 })
);
NOR #() 
NOR_1715_ (
  .A({ S5203 }),
  .B({ S5205 }),
  .Y({ S5207 })
);
NAND #() 
NAND_3206_ (
  .A({ S5204 }),
  .B({ S5206 }),
  .Y({ S5208 })
);
NOR #() 
NOR_1716_ (
  .A({ S2205 }),
  .B({ S5208 }),
  .Y({ S5209 })
);
NAND #() 
NAND_3207_ (
  .A({ S2206 }),
  .B({ S5207 }),
  .Y({ S5210 })
);
NOR #() 
NOR_1717_ (
  .A({ S2206 }),
  .B({ S5207 }),
  .Y({ S5211 })
);
NAND #() 
NAND_3208_ (
  .A({ S2205 }),
  .B({ S5208 }),
  .Y({ S5212 })
);
NOR #() 
NOR_1718_ (
  .A({ S5062 }),
  .B({ S5065 }),
  .Y({ S5213 })
);
NAND #() 
NAND_3209_ (
  .A({ S5061 }),
  .B({ S5066 }),
  .Y({ S5214 })
);
NOR #() 
NOR_1719_ (
  .A({ S5067 }),
  .B({ S5213 }),
  .Y({ S5215 })
);
NAND #() 
NAND_3210_ (
  .A({ S5068 }),
  .B({ S5214 }),
  .Y({ S5216 })
);
NOR #() 
NOR_1720_ (
  .A({ S5113 }),
  .B({ S5215 }),
  .Y({ S5217 })
);
NAND #() 
NAND_3211_ (
  .A({ S5112 }),
  .B({ S5216 }),
  .Y({ S5218 })
);
NOR #() 
NOR_1721_ (
  .A({ S4999 }),
  .B({ S5112 }),
  .Y({ S5219 })
);
NAND #() 
NAND_3212_ (
  .A({ S5000 }),
  .B({ S5113 }),
  .Y({ S5220 })
);
NOR #() 
NOR_1722_ (
  .A({ S5217 }),
  .B({ S5219 }),
  .Y({ S5221 })
);
NAND #() 
NAND_3213_ (
  .A({ S5218 }),
  .B({ S5220 }),
  .Y({ S5222 })
);
NOR #() 
NOR_1723_ (
  .A({ S2106 }),
  .B({ S5222 }),
  .Y({ S5223 })
);
NAND #() 
NAND_3214_ (
  .A({ S2107 }),
  .B({ S5221 }),
  .Y({ S5224 })
);
NAND #() 
NAND_3215_ (
  .A({ S5012 }),
  .B({ S5113 }),
  .Y({ S5225 })
);
NAND #() 
NAND_3216_ (
  .A({ S5018 }),
  .B({ S5057 }),
  .Y({ S5226 })
);
NAND #() 
NAND_3217_ (
  .A({ S5060 }),
  .B({ S5226 }),
  .Y({ S5227 })
);
NAND #() 
NAND_3218_ (
  .A({ S5112 }),
  .B({ S5227 }),
  .Y({ S5228 })
);
NAND #() 
NAND_3219_ (
  .A({ S5225 }),
  .B({ S5228 }),
  .Y({ S5229 })
);
NOT #() 
NOT_396_ (
  .A({ S5229 }),
  .Y({ S5230 })
);
NOR #() 
NOR_1724_ (
  .A({ S1597 }),
  .B({ S5229 }),
  .Y({ S5231 })
);
NAND #() 
NAND_3220_ (
  .A({ S1598 }),
  .B({ S5230 }),
  .Y({ S5232 })
);
NAND #() 
NAND_3221_ (
  .A({ S1597 }),
  .B({ S5229 }),
  .Y({ S5233 })
);
NAND #() 
NAND_3222_ (
  .A({ S5232 }),
  .B({ S5233 }),
  .Y({ S5234 })
);
NOT #() 
NOT_397_ (
  .A({ S5234 }),
  .Y({ S5235 })
);
NAND #() 
NAND_3223_ (
  .A({ S5034 }),
  .B({ S5053 }),
  .Y({ S5236 })
);
NAND #() 
NAND_3224_ (
  .A({ S5056 }),
  .B({ S5236 }),
  .Y({ S5237 })
);
NAND #() 
NAND_3225_ (
  .A({ S5112 }),
  .B({ S5237 }),
  .Y({ S5238 })
);
NAND #() 
NAND_3226_ (
  .A({ S5028 }),
  .B({ S5113 }),
  .Y({ S5239 })
);
NAND #() 
NAND_3227_ (
  .A({ S5238 }),
  .B({ S5239 }),
  .Y({ S5240 })
);
NOT #() 
NOT_398_ (
  .A({ S5240 }),
  .Y({ S5241 })
);
NOR #() 
NOR_1725_ (
  .A({ S1952 }),
  .B({ S5240 }),
  .Y({ S5242 })
);
NAND #() 
NAND_3228_ (
  .A({ S1953 }),
  .B({ S5241 }),
  .Y({ S5243 })
);
NAND #() 
NAND_3229_ (
  .A({ S1952 }),
  .B({ S5240 }),
  .Y({ S5244 })
);
NAND #() 
NAND_3230_ (
  .A({ S5243 }),
  .B({ S5244 }),
  .Y({ S5245 })
);
NOT #() 
NOT_399_ (
  .A({ S5245 }),
  .Y({ S5246 })
);
NOR #() 
NOR_1726_ (
  .A({ S5046 }),
  .B({ S5049 }),
  .Y({ S5247 })
);
NOR #() 
NOR_1727_ (
  .A({ S5051 }),
  .B({ S5247 }),
  .Y({ S5248 })
);
NOR #() 
NOR_1728_ (
  .A({ S5113 }),
  .B({ S5248 }),
  .Y({ S5249 })
);
NOR #() 
NOR_1729_ (
  .A({ S5042 }),
  .B({ S5112 }),
  .Y({ S5250 })
);
NOR #() 
NOR_1730_ (
  .A({ S5249 }),
  .B({ S5250 }),
  .Y({ S5251 })
);
NOT #() 
NOT_400_ (
  .A({ S5251 }),
  .Y({ S5252 })
);
NOR #() 
NOR_1731_ (
  .A({ S1848 }),
  .B({ S5252 }),
  .Y({ S5253 })
);
NAND #() 
NAND_3231_ (
  .A({ S1849 }),
  .B({ S5251 }),
  .Y({ S5254 })
);
NOR #() 
NOR_1732_ (
  .A({ S1849 }),
  .B({ S5251 }),
  .Y({ S5255 })
);
NAND #() 
NAND_3232_ (
  .A({ S1848 }),
  .B({ S5252 }),
  .Y({ S5256 })
);
NOR #() 
NOR_1733_ (
  .A({ S1516 }),
  .B({ S5113 }),
  .Y({ S5257 })
);
NAND #() 
NAND_3233_ (
  .A({ S1515 }),
  .B({ S5112 }),
  .Y({ S5258 })
);
NOR #() 
NOR_1734_ (
  .A({ S1013 }),
  .B({ S5257 }),
  .Y({ S5259 })
);
NAND #() 
NAND_3234_ (
  .A({ datapath_addsubunit_in1_4 }),
  .B({ S5258 }),
  .Y({ S5260 })
);
NOR #() 
NOR_1735_ (
  .A({ datapath_addsubunit_in1_4 }),
  .B({ S5258 }),
  .Y({ S5261 })
);
NAND #() 
NAND_3235_ (
  .A({ S1013 }),
  .B({ S5257 }),
  .Y({ S5262 })
);
NOR #() 
NOR_1736_ (
  .A({ S5259 }),
  .B({ S5261 }),
  .Y({ S5263 })
);
NAND #() 
NAND_3236_ (
  .A({ S5260 }),
  .B({ S5262 }),
  .Y({ S5264 })
);
NOR #() 
NOR_1737_ (
  .A({ S1745 }),
  .B({ S5263 }),
  .Y({ S5265 })
);
NAND #() 
NAND_3237_ (
  .A({ S1746 }),
  .B({ S5264 }),
  .Y({ S5266 })
);
NOR #() 
NOR_1738_ (
  .A({ S1746 }),
  .B({ S5264 }),
  .Y({ S5267 })
);
NAND #() 
NAND_3238_ (
  .A({ S1745 }),
  .B({ S5263 }),
  .Y({ S5268 })
);
NOR #() 
NOR_1739_ (
  .A({ S5265 }),
  .B({ S5267 }),
  .Y({ S5269 })
);
NAND #() 
NAND_3239_ (
  .A({ S5266 }),
  .B({ S5268 }),
  .Y({ S5270 })
);
NOR #() 
NOR_1740_ (
  .A({ datapath_addsubunit_in1_3 }),
  .B({ S1516 }),
  .Y({ S5271 })
);
NAND #() 
NAND_3240_ (
  .A({ S1065 }),
  .B({ S1515 }),
  .Y({ S5272 })
);
NOR #() 
NOR_1741_ (
  .A({ S5270 }),
  .B({ S5271 }),
  .Y({ S5273 })
);
NAND #() 
NAND_3241_ (
  .A({ S5269 }),
  .B({ S5272 }),
  .Y({ S5274 })
);
NOR #() 
NOR_1742_ (
  .A({ S5265 }),
  .B({ S5273 }),
  .Y({ S5275 })
);
NAND #() 
NAND_3242_ (
  .A({ S5266 }),
  .B({ S5274 }),
  .Y({ S5276 })
);
NOR #() 
NOR_1743_ (
  .A({ S5255 }),
  .B({ S5275 }),
  .Y({ S5277 })
);
NAND #() 
NAND_3243_ (
  .A({ S5256 }),
  .B({ S5276 }),
  .Y({ S5278 })
);
NOR #() 
NOR_1744_ (
  .A({ S5253 }),
  .B({ S5277 }),
  .Y({ S5279 })
);
NAND #() 
NAND_3244_ (
  .A({ S5254 }),
  .B({ S5278 }),
  .Y({ S5280 })
);
NOR #() 
NOR_1745_ (
  .A({ S5245 }),
  .B({ S5279 }),
  .Y({ S5281 })
);
NAND #() 
NAND_3245_ (
  .A({ S5246 }),
  .B({ S5280 }),
  .Y({ S5282 })
);
NOR #() 
NOR_1746_ (
  .A({ S5242 }),
  .B({ S5281 }),
  .Y({ S5283 })
);
NAND #() 
NAND_3246_ (
  .A({ S5243 }),
  .B({ S5282 }),
  .Y({ S5284 })
);
NOR #() 
NOR_1747_ (
  .A({ S5234 }),
  .B({ S5283 }),
  .Y({ S5285 })
);
NAND #() 
NAND_3247_ (
  .A({ S5235 }),
  .B({ S5284 }),
  .Y({ S5286 })
);
NOR #() 
NOR_1748_ (
  .A({ S5231 }),
  .B({ S5285 }),
  .Y({ S5287 })
);
NAND #() 
NAND_3248_ (
  .A({ S5232 }),
  .B({ S5286 }),
  .Y({ S5288 })
);
NOR #() 
NOR_1749_ (
  .A({ S2107 }),
  .B({ S5221 }),
  .Y({ S5289 })
);
NAND #() 
NAND_3249_ (
  .A({ S2106 }),
  .B({ S5222 }),
  .Y({ S5290 })
);
NOR #() 
NOR_1750_ (
  .A({ S5223 }),
  .B({ S5289 }),
  .Y({ S5291 })
);
NAND #() 
NAND_3250_ (
  .A({ S5224 }),
  .B({ S5290 }),
  .Y({ S5292 })
);
NOR #() 
NOR_1751_ (
  .A({ S5287 }),
  .B({ S5292 }),
  .Y({ S5293 })
);
NAND #() 
NAND_3251_ (
  .A({ S5288 }),
  .B({ S5291 }),
  .Y({ S5294 })
);
NOR #() 
NOR_1752_ (
  .A({ S5223 }),
  .B({ S5293 }),
  .Y({ S5295 })
);
NAND #() 
NAND_3252_ (
  .A({ S5224 }),
  .B({ S5294 }),
  .Y({ S5296 })
);
NOR #() 
NOR_1753_ (
  .A({ S5211 }),
  .B({ S5295 }),
  .Y({ S5297 })
);
NAND #() 
NAND_3253_ (
  .A({ S5212 }),
  .B({ S5296 }),
  .Y({ S5298 })
);
NOR #() 
NOR_1754_ (
  .A({ S5209 }),
  .B({ S5297 }),
  .Y({ S5299 })
);
NAND #() 
NAND_3254_ (
  .A({ S5210 }),
  .B({ S5298 }),
  .Y({ S5300 })
);
NOR #() 
NOR_1755_ (
  .A({ S5194 }),
  .B({ S5299 }),
  .Y({ S5301 })
);
NAND #() 
NAND_3255_ (
  .A({ S5193 }),
  .B({ S5300 }),
  .Y({ S5302 })
);
NOR #() 
NOR_1756_ (
  .A({ S5189 }),
  .B({ S5301 }),
  .Y({ S5303 })
);
NAND #() 
NAND_3256_ (
  .A({ S5190 }),
  .B({ S5302 }),
  .Y({ S5304 })
);
NOR #() 
NOR_1757_ (
  .A({ S5177 }),
  .B({ S5303 }),
  .Y({ S5305 })
);
NAND #() 
NAND_3257_ (
  .A({ S5178 }),
  .B({ S5304 }),
  .Y({ S5306 })
);
NOR #() 
NOR_1758_ (
  .A({ S5175 }),
  .B({ S5305 }),
  .Y({ S5307 })
);
NAND #() 
NAND_3258_ (
  .A({ S5176 }),
  .B({ S5306 }),
  .Y({ S5308 })
);
NOR #() 
NOR_1759_ (
  .A({ S5160 }),
  .B({ S5307 }),
  .Y({ S5309 })
);
NAND #() 
NAND_3259_ (
  .A({ S5159 }),
  .B({ S5308 }),
  .Y({ S5310 })
);
NOR #() 
NOR_1760_ (
  .A({ S5156 }),
  .B({ S5309 }),
  .Y({ S5311 })
);
NAND #() 
NAND_3260_ (
  .A({ S5157 }),
  .B({ S5310 }),
  .Y({ S5312 })
);
NAND #() 
NAND_3261_ (
  .A({ S5149 }),
  .B({ S5311 }),
  .Y({ S5313 })
);
NAND #() 
NAND_3262_ (
  .A({ S5148 }),
  .B({ S5312 }),
  .Y({ S5314 })
);
NAND #() 
NAND_3263_ (
  .A({ S5149 }),
  .B({ S5314 }),
  .Y({ S5315 })
);
NAND #() 
NAND_3264_ (
  .A({ S5148 }),
  .B({ S5313 }),
  .Y({ S5316 })
);
NOR #() 
NOR_1761_ (
  .A({ S5137 }),
  .B({ S5316 }),
  .Y({ S5317 })
);
NAND #() 
NAND_3265_ (
  .A({ S5138 }),
  .B({ S5315 }),
  .Y({ S5318 })
);
NOR #() 
NOR_1762_ (
  .A({ S5134 }),
  .B({ S5317 }),
  .Y({ S5319 })
);
NAND #() 
NAND_3266_ (
  .A({ S5135 }),
  .B({ S5318 }),
  .Y({ S5320 })
);
NOR #() 
NOR_1763_ (
  .A({ S2817 }),
  .B({ S3903 }),
  .Y({ S5321 })
);
NOR #() 
NOR_1764_ (
  .A({ S3905 }),
  .B({ S5320 }),
  .Y({ S5322 })
);
NAND #() 
NAND_3267_ (
  .A({ S5320 }),
  .B({ S5321 }),
  .Y({ S5323 })
);
NAND #() 
NAND_3268_ (
  .A({ S5123 }),
  .B({ S5323 }),
  .Y({ S5324 })
);
NAND #() 
NAND_3269_ (
  .A({ S2817 }),
  .B({ S5123 }),
  .Y({ S5325 })
);
NOT #() 
NOT_401_ (
  .A({ S5325 }),
  .Y({ S5326 })
);
NOR #() 
NOR_1765_ (
  .A({ S5320 }),
  .B({ S5326 }),
  .Y({ S5327 })
);
NAND #() 
NAND_3270_ (
  .A({ S5319 }),
  .B({ S5325 }),
  .Y({ S5328 })
);
NOR #() 
NOR_1766_ (
  .A({ S2817 }),
  .B({ S5123 }),
  .Y({ S5329 })
);
NOR #() 
NOR_1767_ (
  .A({ S3903 }),
  .B({ S5329 }),
  .Y({ S5330 })
);
NOT #() 
NOT_402_ (
  .A({ S5330 }),
  .Y({ S5331 })
);
NOR #() 
NOR_1768_ (
  .A({ S5327 }),
  .B({ S5331 }),
  .Y({ S5332 })
);
NAND #() 
NAND_3271_ (
  .A({ S5328 }),
  .B({ S5330 }),
  .Y({ S5333 })
);
NOR #() 
NOR_1769_ (
  .A({ S5322 }),
  .B({ S5324 }),
  .Y({ S5334 })
);
NAND #() 
NAND_3272_ (
  .A({ S2920 }),
  .B({ S5334 }),
  .Y({ S5335 })
);
NOT #() 
NOT_403_ (
  .A({ S5335 }),
  .Y({ S5336 })
);
NAND #() 
NAND_3273_ (
  .A({ S5137 }),
  .B({ S5316 }),
  .Y({ S5337 })
);
NAND #() 
NAND_3274_ (
  .A({ S5318 }),
  .B({ S5337 }),
  .Y({ S5338 })
);
NAND #() 
NAND_3275_ (
  .A({ S5332 }),
  .B({ S5338 }),
  .Y({ S5339 })
);
NAND #() 
NAND_3276_ (
  .A({ S5133 }),
  .B({ S5333 }),
  .Y({ S5340 })
);
NAND #() 
NAND_3277_ (
  .A({ S5339 }),
  .B({ S5340 }),
  .Y({ S5341 })
);
NOT #() 
NOT_404_ (
  .A({ S5341 }),
  .Y({ S5342 })
);
NOR #() 
NOR_1770_ (
  .A({ S2816 }),
  .B({ S5341 }),
  .Y({ S5343 })
);
NAND #() 
NAND_3278_ (
  .A({ S2817 }),
  .B({ S5342 }),
  .Y({ S5344 })
);
NAND #() 
NAND_3279_ (
  .A({ S2816 }),
  .B({ S5341 }),
  .Y({ S5345 })
);
NAND #() 
NAND_3280_ (
  .A({ S5344 }),
  .B({ S5345 }),
  .Y({ S5346 })
);
NOT #() 
NOT_405_ (
  .A({ S5346 }),
  .Y({ S5347 })
);
NAND #() 
NAND_3281_ (
  .A({ S5148 }),
  .B({ S5149 }),
  .Y({ S5348 })
);
NAND #() 
NAND_3282_ (
  .A({ S5311 }),
  .B({ S5348 }),
  .Y({ S5349 })
);
NOR #() 
NOR_1771_ (
  .A({ S5311 }),
  .B({ S5348 }),
  .Y({ S5350 })
);
NOT #() 
NOT_406_ (
  .A({ S5350 }),
  .Y({ S5351 })
);
NAND #() 
NAND_3283_ (
  .A({ S5349 }),
  .B({ S5351 }),
  .Y({ S5352 })
);
NAND #() 
NAND_3284_ (
  .A({ S5332 }),
  .B({ S5352 }),
  .Y({ S5353 })
);
NOT #() 
NOT_407_ (
  .A({ S5353 }),
  .Y({ S5354 })
);
NOR #() 
NOR_1772_ (
  .A({ S5146 }),
  .B({ S5332 }),
  .Y({ S5355 })
);
NOR #() 
NOR_1773_ (
  .A({ S5354 }),
  .B({ S5355 }),
  .Y({ S5356 })
);
NOT #() 
NOT_408_ (
  .A({ S5356 }),
  .Y({ S5357 })
);
NAND #() 
NAND_3285_ (
  .A({ S2717 }),
  .B({ S5357 }),
  .Y({ S5358 })
);
NAND #() 
NAND_3286_ (
  .A({ S2718 }),
  .B({ S5356 }),
  .Y({ S5359 })
);
NOR #() 
NOR_1774_ (
  .A({ S5159 }),
  .B({ S5308 }),
  .Y({ S5360 })
);
NOR #() 
NOR_1775_ (
  .A({ S5309 }),
  .B({ S5360 }),
  .Y({ S5361 })
);
NOR #() 
NOR_1776_ (
  .A({ S5333 }),
  .B({ S5361 }),
  .Y({ S5362 })
);
NOR #() 
NOR_1777_ (
  .A({ S5154 }),
  .B({ S5332 }),
  .Y({ S5363 })
);
NOR #() 
NOR_1778_ (
  .A({ S5362 }),
  .B({ S5363 }),
  .Y({ S5364 })
);
NOT #() 
NOT_409_ (
  .A({ S5364 }),
  .Y({ S5365 })
);
NOR #() 
NOR_1779_ (
  .A({ S2617 }),
  .B({ S5365 }),
  .Y({ S5366 })
);
NOT #() 
NOT_410_ (
  .A({ S5366 }),
  .Y({ S5367 })
);
NOR #() 
NOR_1780_ (
  .A({ S2618 }),
  .B({ S5364 }),
  .Y({ S5368 })
);
NOR #() 
NOR_1781_ (
  .A({ S5366 }),
  .B({ S5368 }),
  .Y({ S5369 })
);
NOT #() 
NOT_411_ (
  .A({ S5369 }),
  .Y({ S5370 })
);
NOR #() 
NOR_1782_ (
  .A({ S5175 }),
  .B({ S5177 }),
  .Y({ S5371 })
);
NAND #() 
NAND_3287_ (
  .A({ S5176 }),
  .B({ S5178 }),
  .Y({ S5372 })
);
NOR #() 
NOR_1783_ (
  .A({ S5304 }),
  .B({ S5371 }),
  .Y({ S5373 })
);
NOR #() 
NOR_1784_ (
  .A({ S5303 }),
  .B({ S5372 }),
  .Y({ S5374 })
);
NOR #() 
NOR_1785_ (
  .A({ S5373 }),
  .B({ S5374 }),
  .Y({ S5375 })
);
NOR #() 
NOR_1786_ (
  .A({ S5174 }),
  .B({ S5332 }),
  .Y({ S5376 })
);
NAND #() 
NAND_3288_ (
  .A({ S5173 }),
  .B({ S5333 }),
  .Y({ S5377 })
);
NAND #() 
NAND_3289_ (
  .A({ S5332 }),
  .B({ S5375 }),
  .Y({ S5378 })
);
NOT #() 
NOT_412_ (
  .A({ S5378 }),
  .Y({ S5379 })
);
NAND #() 
NAND_3290_ (
  .A({ S5377 }),
  .B({ S5378 }),
  .Y({ S5380 })
);
NOR #() 
NOR_1787_ (
  .A({ S5376 }),
  .B({ S5379 }),
  .Y({ S5381 })
);
NOR #() 
NOR_1788_ (
  .A({ S2518 }),
  .B({ S5380 }),
  .Y({ S5382 })
);
NOR #() 
NOR_1789_ (
  .A({ S2517 }),
  .B({ S5381 }),
  .Y({ S5383 })
);
NAND #() 
NAND_3291_ (
  .A({ S5194 }),
  .B({ S5299 }),
  .Y({ S5384 })
);
NAND #() 
NAND_3292_ (
  .A({ S5302 }),
  .B({ S5384 }),
  .Y({ S5385 })
);
NAND #() 
NAND_3293_ (
  .A({ S5332 }),
  .B({ S5385 }),
  .Y({ S5386 })
);
NAND #() 
NAND_3294_ (
  .A({ S5188 }),
  .B({ S5333 }),
  .Y({ S5387 })
);
NAND #() 
NAND_3295_ (
  .A({ S5386 }),
  .B({ S5387 }),
  .Y({ S5388 })
);
NOT #() 
NOT_413_ (
  .A({ S5388 }),
  .Y({ S5389 })
);
NOR #() 
NOR_1790_ (
  .A({ S2417 }),
  .B({ S5388 }),
  .Y({ S5390 })
);
NAND #() 
NAND_3296_ (
  .A({ S2418 }),
  .B({ S5389 }),
  .Y({ S5391 })
);
NAND #() 
NAND_3297_ (
  .A({ S2417 }),
  .B({ S5388 }),
  .Y({ S5392 })
);
NAND #() 
NAND_3298_ (
  .A({ S5391 }),
  .B({ S5392 }),
  .Y({ S5393 })
);
NOT #() 
NOT_414_ (
  .A({ S5393 }),
  .Y({ S5394 })
);
NOR #() 
NOR_1791_ (
  .A({ S5209 }),
  .B({ S5211 }),
  .Y({ S5395 })
);
NAND #() 
NAND_3299_ (
  .A({ S5210 }),
  .B({ S5212 }),
  .Y({ S5396 })
);
NOR #() 
NOR_1792_ (
  .A({ S5296 }),
  .B({ S5395 }),
  .Y({ S5397 })
);
NOR #() 
NOR_1793_ (
  .A({ S5295 }),
  .B({ S5396 }),
  .Y({ S5398 })
);
NOR #() 
NOR_1794_ (
  .A({ S5397 }),
  .B({ S5398 }),
  .Y({ S5399 })
);
NOR #() 
NOR_1795_ (
  .A({ S5333 }),
  .B({ S5399 }),
  .Y({ S5400 })
);
NOR #() 
NOR_1796_ (
  .A({ S5207 }),
  .B({ S5332 }),
  .Y({ S5401 })
);
NOR #() 
NOR_1797_ (
  .A({ S5400 }),
  .B({ S5401 }),
  .Y({ S5402 })
);
NOT #() 
NOT_415_ (
  .A({ S5402 }),
  .Y({ S5403 })
);
NOR #() 
NOR_1798_ (
  .A({ S2311 }),
  .B({ S5403 }),
  .Y({ S5404 })
);
NOR #() 
NOR_1799_ (
  .A({ S2312 }),
  .B({ S5402 }),
  .Y({ S5405 })
);
NOR #() 
NOR_1800_ (
  .A({ S5288 }),
  .B({ S5291 }),
  .Y({ S5406 })
);
NOT #() 
NOT_416_ (
  .A({ S5406 }),
  .Y({ S5407 })
);
NAND #() 
NAND_3300_ (
  .A({ S5294 }),
  .B({ S5407 }),
  .Y({ S5408 })
);
NAND #() 
NAND_3301_ (
  .A({ S5332 }),
  .B({ S5408 }),
  .Y({ S5409 })
);
NAND #() 
NAND_3302_ (
  .A({ S5222 }),
  .B({ S5333 }),
  .Y({ S5410 })
);
NAND #() 
NAND_3303_ (
  .A({ S5409 }),
  .B({ S5410 }),
  .Y({ S5411 })
);
NOT #() 
NOT_417_ (
  .A({ S5411 }),
  .Y({ S5412 })
);
NOR #() 
NOR_1801_ (
  .A({ S2205 }),
  .B({ S5411 }),
  .Y({ S5413 })
);
NAND #() 
NAND_3304_ (
  .A({ S2206 }),
  .B({ S5412 }),
  .Y({ S5414 })
);
NAND #() 
NAND_3305_ (
  .A({ S5234 }),
  .B({ S5283 }),
  .Y({ S5415 })
);
NAND #() 
NAND_3306_ (
  .A({ S5286 }),
  .B({ S5415 }),
  .Y({ S5416 })
);
NAND #() 
NAND_3307_ (
  .A({ S5332 }),
  .B({ S5416 }),
  .Y({ S5417 })
);
NAND #() 
NAND_3308_ (
  .A({ S5229 }),
  .B({ S5333 }),
  .Y({ S5418 })
);
NAND #() 
NAND_3309_ (
  .A({ S5417 }),
  .B({ S5418 }),
  .Y({ S5419 })
);
NOT #() 
NOT_418_ (
  .A({ S5419 }),
  .Y({ S5420 })
);
NAND #() 
NAND_3310_ (
  .A({ S2107 }),
  .B({ S5420 }),
  .Y({ S5421 })
);
NOT #() 
NOT_419_ (
  .A({ S5421 }),
  .Y({ S5422 })
);
NAND #() 
NAND_3311_ (
  .A({ S2106 }),
  .B({ S5419 }),
  .Y({ S5423 })
);
NAND #() 
NAND_3312_ (
  .A({ S5421 }),
  .B({ S5423 }),
  .Y({ S5424 })
);
NOT #() 
NOT_420_ (
  .A({ S5424 }),
  .Y({ S5425 })
);
NAND #() 
NAND_3313_ (
  .A({ S5245 }),
  .B({ S5279 }),
  .Y({ S5426 })
);
NAND #() 
NAND_3314_ (
  .A({ S5282 }),
  .B({ S5426 }),
  .Y({ S5427 })
);
NAND #() 
NAND_3315_ (
  .A({ S5332 }),
  .B({ S5427 }),
  .Y({ S5428 })
);
NAND #() 
NAND_3316_ (
  .A({ S5240 }),
  .B({ S5333 }),
  .Y({ S5429 })
);
NAND #() 
NAND_3317_ (
  .A({ S5428 }),
  .B({ S5429 }),
  .Y({ S5430 })
);
NOT #() 
NOT_421_ (
  .A({ S5430 }),
  .Y({ S5431 })
);
NAND #() 
NAND_3318_ (
  .A({ S1598 }),
  .B({ S5431 }),
  .Y({ S5432 })
);
NOT #() 
NOT_422_ (
  .A({ S5432 }),
  .Y({ S5433 })
);
NAND #() 
NAND_3319_ (
  .A({ S1597 }),
  .B({ S5430 }),
  .Y({ S5434 })
);
NAND #() 
NAND_3320_ (
  .A({ S5432 }),
  .B({ S5434 }),
  .Y({ S5435 })
);
NOT #() 
NOT_423_ (
  .A({ S5435 }),
  .Y({ S5436 })
);
NOR #() 
NOR_1802_ (
  .A({ S5253 }),
  .B({ S5255 }),
  .Y({ S5437 })
);
NAND #() 
NAND_3321_ (
  .A({ S5254 }),
  .B({ S5256 }),
  .Y({ S5438 })
);
NAND #() 
NAND_3322_ (
  .A({ S5275 }),
  .B({ S5437 }),
  .Y({ S5439 })
);
NAND #() 
NAND_3323_ (
  .A({ S5276 }),
  .B({ S5438 }),
  .Y({ S5440 })
);
NAND #() 
NAND_3324_ (
  .A({ S5439 }),
  .B({ S5440 }),
  .Y({ S5441 })
);
NAND #() 
NAND_3325_ (
  .A({ S5332 }),
  .B({ S5441 }),
  .Y({ S5442 })
);
NAND #() 
NAND_3326_ (
  .A({ S5251 }),
  .B({ S5333 }),
  .Y({ S5443 })
);
NAND #() 
NAND_3327_ (
  .A({ S5442 }),
  .B({ S5443 }),
  .Y({ S5444 })
);
NOT #() 
NOT_424_ (
  .A({ S5444 }),
  .Y({ S5445 })
);
NOR #() 
NOR_1803_ (
  .A({ S1952 }),
  .B({ S5445 }),
  .Y({ S5446 })
);
NAND #() 
NAND_3328_ (
  .A({ S1953 }),
  .B({ S5444 }),
  .Y({ S5447 })
);
NOR #() 
NOR_1804_ (
  .A({ S1953 }),
  .B({ S5444 }),
  .Y({ S5448 })
);
NAND #() 
NAND_3329_ (
  .A({ S1952 }),
  .B({ S5445 }),
  .Y({ S5449 })
);
NOR #() 
NOR_1805_ (
  .A({ S5269 }),
  .B({ S5272 }),
  .Y({ S5450 })
);
NOR #() 
NOR_1806_ (
  .A({ S5273 }),
  .B({ S5450 }),
  .Y({ S5451 })
);
NAND #() 
NAND_3330_ (
  .A({ S5332 }),
  .B({ S5451 }),
  .Y({ S5452 })
);
NOT #() 
NOT_425_ (
  .A({ S5452 }),
  .Y({ S5453 })
);
NOR #() 
NOR_1807_ (
  .A({ S5263 }),
  .B({ S5332 }),
  .Y({ S5454 })
);
NOT #() 
NOT_426_ (
  .A({ S5454 }),
  .Y({ S5455 })
);
NOR #() 
NOR_1808_ (
  .A({ S5453 }),
  .B({ S5454 }),
  .Y({ S5456 })
);
NAND #() 
NAND_3331_ (
  .A({ S5452 }),
  .B({ S5455 }),
  .Y({ S5457 })
);
NOR #() 
NOR_1809_ (
  .A({ S1848 }),
  .B({ S5456 }),
  .Y({ S5458 })
);
NAND #() 
NAND_3332_ (
  .A({ S1849 }),
  .B({ S5457 }),
  .Y({ S5459 })
);
NOR #() 
NOR_1810_ (
  .A({ S1849 }),
  .B({ S5457 }),
  .Y({ S5460 })
);
NAND #() 
NAND_3333_ (
  .A({ S1848 }),
  .B({ S5456 }),
  .Y({ S5461 })
);
NOR #() 
NOR_1811_ (
  .A({ S5458 }),
  .B({ S5460 }),
  .Y({ S5462 })
);
NAND #() 
NAND_3334_ (
  .A({ S5459 }),
  .B({ S5461 }),
  .Y({ S5463 })
);
NOR #() 
NOR_1812_ (
  .A({ S1516 }),
  .B({ S5333 }),
  .Y({ S5464 })
);
NAND #() 
NAND_3335_ (
  .A({ S1515 }),
  .B({ S5332 }),
  .Y({ S5465 })
);
NOR #() 
NOR_1813_ (
  .A({ S1065 }),
  .B({ S5464 }),
  .Y({ S5466 })
);
NAND #() 
NAND_3336_ (
  .A({ datapath_addsubunit_in1_3 }),
  .B({ S5465 }),
  .Y({ S5467 })
);
NAND #() 
NAND_3337_ (
  .A({ S5271 }),
  .B({ S5332 }),
  .Y({ S5468 })
);
NOT #() 
NOT_427_ (
  .A({ S5468 }),
  .Y({ S5469 })
);
NOR #() 
NOR_1814_ (
  .A({ S5466 }),
  .B({ S5469 }),
  .Y({ S5470 })
);
NAND #() 
NAND_3338_ (
  .A({ S5467 }),
  .B({ S5468 }),
  .Y({ S5471 })
);
NOR #() 
NOR_1815_ (
  .A({ S1745 }),
  .B({ S5470 }),
  .Y({ S5472 })
);
NAND #() 
NAND_3339_ (
  .A({ S1746 }),
  .B({ S5471 }),
  .Y({ S5473 })
);
NOR #() 
NOR_1816_ (
  .A({ datapath_addsubunit_in1_2 }),
  .B({ S1516 }),
  .Y({ S5474 })
);
NAND #() 
NAND_3340_ (
  .A({ S1116 }),
  .B({ S1515 }),
  .Y({ S5475 })
);
NOR #() 
NOR_1817_ (
  .A({ S1746 }),
  .B({ S5471 }),
  .Y({ S5476 })
);
NAND #() 
NAND_3341_ (
  .A({ S1745 }),
  .B({ S5470 }),
  .Y({ S5477 })
);
NOR #() 
NOR_1818_ (
  .A({ S5472 }),
  .B({ S5476 }),
  .Y({ S5478 })
);
NAND #() 
NAND_3342_ (
  .A({ S5473 }),
  .B({ S5477 }),
  .Y({ S5479 })
);
NOR #() 
NOR_1819_ (
  .A({ S5474 }),
  .B({ S5479 }),
  .Y({ S5480 })
);
NAND #() 
NAND_3343_ (
  .A({ S5475 }),
  .B({ S5478 }),
  .Y({ S5481 })
);
NOR #() 
NOR_1820_ (
  .A({ S5472 }),
  .B({ S5480 }),
  .Y({ S5482 })
);
NAND #() 
NAND_3344_ (
  .A({ S5473 }),
  .B({ S5481 }),
  .Y({ S5483 })
);
NOR #() 
NOR_1821_ (
  .A({ S5463 }),
  .B({ S5482 }),
  .Y({ S5484 })
);
NAND #() 
NAND_3345_ (
  .A({ S5462 }),
  .B({ S5483 }),
  .Y({ S5485 })
);
NOR #() 
NOR_1822_ (
  .A({ S5458 }),
  .B({ S5484 }),
  .Y({ S5486 })
);
NAND #() 
NAND_3346_ (
  .A({ S5459 }),
  .B({ S5485 }),
  .Y({ S5487 })
);
NOR #() 
NOR_1823_ (
  .A({ S5448 }),
  .B({ S5486 }),
  .Y({ S5488 })
);
NAND #() 
NAND_3347_ (
  .A({ S5449 }),
  .B({ S5487 }),
  .Y({ S5489 })
);
NOR #() 
NOR_1824_ (
  .A({ S5446 }),
  .B({ S5488 }),
  .Y({ S5490 })
);
NAND #() 
NAND_3348_ (
  .A({ S5447 }),
  .B({ S5489 }),
  .Y({ S5491 })
);
NOR #() 
NOR_1825_ (
  .A({ S5435 }),
  .B({ S5490 }),
  .Y({ S5492 })
);
NAND #() 
NAND_3349_ (
  .A({ S5436 }),
  .B({ S5491 }),
  .Y({ S5493 })
);
NOR #() 
NOR_1826_ (
  .A({ S5433 }),
  .B({ S5492 }),
  .Y({ S5494 })
);
NAND #() 
NAND_3350_ (
  .A({ S5432 }),
  .B({ S5493 }),
  .Y({ S5495 })
);
NOR #() 
NOR_1827_ (
  .A({ S5424 }),
  .B({ S5494 }),
  .Y({ S5496 })
);
NAND #() 
NAND_3351_ (
  .A({ S5425 }),
  .B({ S5495 }),
  .Y({ S5497 })
);
NOR #() 
NOR_1828_ (
  .A({ S5422 }),
  .B({ S5496 }),
  .Y({ S5498 })
);
NAND #() 
NAND_3352_ (
  .A({ S5421 }),
  .B({ S5497 }),
  .Y({ S5499 })
);
NAND #() 
NAND_3353_ (
  .A({ S2205 }),
  .B({ S5411 }),
  .Y({ S5500 })
);
NOT #() 
NOT_428_ (
  .A({ S5500 }),
  .Y({ S5501 })
);
NOR #() 
NOR_1829_ (
  .A({ S5413 }),
  .B({ S5501 }),
  .Y({ S5502 })
);
NOT #() 
NOT_429_ (
  .A({ S5502 }),
  .Y({ S5503 })
);
NOR #() 
NOR_1830_ (
  .A({ S5498 }),
  .B({ S5503 }),
  .Y({ S5504 })
);
NAND #() 
NAND_3354_ (
  .A({ S5499 }),
  .B({ S5502 }),
  .Y({ S5505 })
);
NOR #() 
NOR_1831_ (
  .A({ S5413 }),
  .B({ S5504 }),
  .Y({ S5506 })
);
NAND #() 
NAND_3355_ (
  .A({ S5414 }),
  .B({ S5505 }),
  .Y({ S5507 })
);
NOR #() 
NOR_1832_ (
  .A({ S5405 }),
  .B({ S5506 }),
  .Y({ S5508 })
);
NOR #() 
NOR_1833_ (
  .A({ S5404 }),
  .B({ S5507 }),
  .Y({ S5509 })
);
NOR #() 
NOR_1834_ (
  .A({ S5404 }),
  .B({ S5508 }),
  .Y({ S5510 })
);
NOR #() 
NOR_1835_ (
  .A({ S5405 }),
  .B({ S5509 }),
  .Y({ S5511 })
);
NOR #() 
NOR_1836_ (
  .A({ S5393 }),
  .B({ S5510 }),
  .Y({ S5512 })
);
NAND #() 
NAND_3356_ (
  .A({ S5394 }),
  .B({ S5511 }),
  .Y({ S5513 })
);
NOR #() 
NOR_1837_ (
  .A({ S5390 }),
  .B({ S5512 }),
  .Y({ S5514 })
);
NAND #() 
NAND_3357_ (
  .A({ S5391 }),
  .B({ S5513 }),
  .Y({ S5515 })
);
NOR #() 
NOR_1838_ (
  .A({ S5383 }),
  .B({ S5515 }),
  .Y({ S5516 })
);
NOR #() 
NOR_1839_ (
  .A({ S5382 }),
  .B({ S5514 }),
  .Y({ S5517 })
);
NOR #() 
NOR_1840_ (
  .A({ S5382 }),
  .B({ S5516 }),
  .Y({ S5518 })
);
NOR #() 
NOR_1841_ (
  .A({ S5383 }),
  .B({ S5517 }),
  .Y({ S5519 })
);
NOR #() 
NOR_1842_ (
  .A({ S5370 }),
  .B({ S5519 }),
  .Y({ S5520 })
);
NAND #() 
NAND_3358_ (
  .A({ S5369 }),
  .B({ S5518 }),
  .Y({ S5521 })
);
NOR #() 
NOR_1843_ (
  .A({ S5366 }),
  .B({ S5520 }),
  .Y({ S5522 })
);
NAND #() 
NAND_3359_ (
  .A({ S5367 }),
  .B({ S5521 }),
  .Y({ S5523 })
);
NAND #() 
NAND_3360_ (
  .A({ S5359 }),
  .B({ S5522 }),
  .Y({ S5524 })
);
NAND #() 
NAND_3361_ (
  .A({ S5358 }),
  .B({ S5523 }),
  .Y({ S5525 })
);
NAND #() 
NAND_3362_ (
  .A({ S5359 }),
  .B({ S5525 }),
  .Y({ S5526 })
);
NAND #() 
NAND_3363_ (
  .A({ S5358 }),
  .B({ S5524 }),
  .Y({ S5527 })
);
NOR #() 
NOR_1844_ (
  .A({ S5346 }),
  .B({ S5527 }),
  .Y({ S5528 })
);
NAND #() 
NAND_3364_ (
  .A({ S5347 }),
  .B({ S5526 }),
  .Y({ S5529 })
);
NOR #() 
NOR_1845_ (
  .A({ S5343 }),
  .B({ S5528 }),
  .Y({ S5530 })
);
NAND #() 
NAND_3365_ (
  .A({ S5344 }),
  .B({ S5529 }),
  .Y({ S5531 })
);
NOR #() 
NOR_1846_ (
  .A({ S5336 }),
  .B({ S5531 }),
  .Y({ S5532 })
);
NAND #() 
NAND_3366_ (
  .A({ S5335 }),
  .B({ S5530 }),
  .Y({ S5533 })
);
NOR #() 
NOR_1847_ (
  .A({ S2920 }),
  .B({ S5334 }),
  .Y({ S5534 })
);
NOT #() 
NOT_430_ (
  .A({ S5534 }),
  .Y({ S5535 })
);
NOR #() 
NOR_1848_ (
  .A({ S3901 }),
  .B({ S5534 }),
  .Y({ S5536 })
);
NAND #() 
NAND_3367_ (
  .A({ S3900 }),
  .B({ S5535 }),
  .Y({ S5537 })
);
NOR #() 
NOR_1849_ (
  .A({ S5532 }),
  .B({ S5537 }),
  .Y({ S5538 })
);
NAND #() 
NAND_3368_ (
  .A({ S5533 }),
  .B({ S5536 }),
  .Y({ S5539 })
);
NAND #() 
NAND_3369_ (
  .A({ S5346 }),
  .B({ S5527 }),
  .Y({ S5540 })
);
NAND #() 
NAND_3370_ (
  .A({ S5529 }),
  .B({ S5540 }),
  .Y({ S5541 })
);
NAND #() 
NAND_3371_ (
  .A({ S5538 }),
  .B({ S5541 }),
  .Y({ S5542 })
);
NAND #() 
NAND_3372_ (
  .A({ S5341 }),
  .B({ S5539 }),
  .Y({ S5543 })
);
NAND #() 
NAND_3373_ (
  .A({ S5542 }),
  .B({ S5543 }),
  .Y({ S5544 })
);
NOT #() 
NOT_431_ (
  .A({ S5544 }),
  .Y({ S5545 })
);
NAND #() 
NAND_3374_ (
  .A({ S2920 }),
  .B({ S5545 }),
  .Y({ S5546 })
);
NOT #() 
NOT_432_ (
  .A({ S5546 }),
  .Y({ S5547 })
);
NAND #() 
NAND_3375_ (
  .A({ S2919 }),
  .B({ S5544 }),
  .Y({ S5548 })
);
NAND #() 
NAND_3376_ (
  .A({ S5546 }),
  .B({ S5548 }),
  .Y({ S5549 })
);
NOT #() 
NOT_433_ (
  .A({ S5549 }),
  .Y({ S5550 })
);
NAND #() 
NAND_3377_ (
  .A({ S5358 }),
  .B({ S5359 }),
  .Y({ S5551 })
);
NAND #() 
NAND_3378_ (
  .A({ S5522 }),
  .B({ S5551 }),
  .Y({ S5552 })
);
NOT #() 
NOT_434_ (
  .A({ S5552 }),
  .Y({ S5553 })
);
NOR #() 
NOR_1850_ (
  .A({ S5522 }),
  .B({ S5551 }),
  .Y({ S5554 })
);
NOR #() 
NOR_1851_ (
  .A({ S5553 }),
  .B({ S5554 }),
  .Y({ S5555 })
);
NOR #() 
NOR_1852_ (
  .A({ S5539 }),
  .B({ S5555 }),
  .Y({ S5556 })
);
NOR #() 
NOR_1853_ (
  .A({ S5356 }),
  .B({ S5538 }),
  .Y({ S5557 })
);
NOR #() 
NOR_1854_ (
  .A({ S5556 }),
  .B({ S5557 }),
  .Y({ S5558 })
);
NOT #() 
NOT_435_ (
  .A({ S5558 }),
  .Y({ S5559 })
);
NAND #() 
NAND_3379_ (
  .A({ S2817 }),
  .B({ S5558 }),
  .Y({ S5560 })
);
NAND #() 
NAND_3380_ (
  .A({ S2816 }),
  .B({ S5559 }),
  .Y({ S5561 })
);
NOR #() 
NOR_1855_ (
  .A({ S5369 }),
  .B({ S5518 }),
  .Y({ S5562 })
);
NOR #() 
NOR_1856_ (
  .A({ S5520 }),
  .B({ S5562 }),
  .Y({ S5563 })
);
NOR #() 
NOR_1857_ (
  .A({ S5539 }),
  .B({ S5563 }),
  .Y({ S5564 })
);
NOR #() 
NOR_1858_ (
  .A({ S5364 }),
  .B({ S5538 }),
  .Y({ S5565 })
);
NOR #() 
NOR_1859_ (
  .A({ S5564 }),
  .B({ S5565 }),
  .Y({ S5566 })
);
NOT #() 
NOT_436_ (
  .A({ S5566 }),
  .Y({ S5567 })
);
NOR #() 
NOR_1860_ (
  .A({ S2717 }),
  .B({ S5567 }),
  .Y({ S5568 })
);
NOT #() 
NOT_437_ (
  .A({ S5568 }),
  .Y({ S5569 })
);
NOR #() 
NOR_1861_ (
  .A({ S2718 }),
  .B({ S5566 }),
  .Y({ S5570 })
);
NOR #() 
NOR_1862_ (
  .A({ S5568 }),
  .B({ S5570 }),
  .Y({ S5571 })
);
NOT #() 
NOT_438_ (
  .A({ S5571 }),
  .Y({ S5572 })
);
NOR #() 
NOR_1863_ (
  .A({ S5382 }),
  .B({ S5383 }),
  .Y({ S5573 })
);
NOR #() 
NOR_1864_ (
  .A({ S5515 }),
  .B({ S5573 }),
  .Y({ S5574 })
);
NOT #() 
NOT_439_ (
  .A({ S5574 }),
  .Y({ S5575 })
);
NAND #() 
NAND_3381_ (
  .A({ S5515 }),
  .B({ S5573 }),
  .Y({ S5576 })
);
NOT #() 
NOT_440_ (
  .A({ S5576 }),
  .Y({ S5577 })
);
NOR #() 
NOR_1865_ (
  .A({ S5574 }),
  .B({ S5577 }),
  .Y({ S5578 })
);
NAND #() 
NAND_3382_ (
  .A({ S5575 }),
  .B({ S5576 }),
  .Y({ S5579 })
);
NOR #() 
NOR_1866_ (
  .A({ S5539 }),
  .B({ S5578 }),
  .Y({ S5580 })
);
NAND #() 
NAND_3383_ (
  .A({ S5538 }),
  .B({ S5579 }),
  .Y({ S5581 })
);
NOR #() 
NOR_1867_ (
  .A({ S5380 }),
  .B({ S5538 }),
  .Y({ S5582 })
);
NAND #() 
NAND_3384_ (
  .A({ S5381 }),
  .B({ S5539 }),
  .Y({ S5583 })
);
NOR #() 
NOR_1868_ (
  .A({ S5580 }),
  .B({ S5582 }),
  .Y({ S5584 })
);
NAND #() 
NAND_3385_ (
  .A({ S5581 }),
  .B({ S5583 }),
  .Y({ S5585 })
);
NAND #() 
NAND_3386_ (
  .A({ S2618 }),
  .B({ S5584 }),
  .Y({ S5586 })
);
NAND #() 
NAND_3387_ (
  .A({ S2617 }),
  .B({ S5585 }),
  .Y({ S5587 })
);
NAND #() 
NAND_3388_ (
  .A({ S5393 }),
  .B({ S5510 }),
  .Y({ S5588 })
);
NAND #() 
NAND_3389_ (
  .A({ S5513 }),
  .B({ S5588 }),
  .Y({ S5589 })
);
NAND #() 
NAND_3390_ (
  .A({ S5538 }),
  .B({ S5589 }),
  .Y({ S5590 })
);
NAND #() 
NAND_3391_ (
  .A({ S5388 }),
  .B({ S5539 }),
  .Y({ S5591 })
);
NAND #() 
NAND_3392_ (
  .A({ S5590 }),
  .B({ S5591 }),
  .Y({ S5592 })
);
NOT #() 
NOT_441_ (
  .A({ S5592 }),
  .Y({ S5593 })
);
NAND #() 
NAND_3393_ (
  .A({ S2518 }),
  .B({ S5593 }),
  .Y({ S5594 })
);
NOT #() 
NOT_442_ (
  .A({ S5594 }),
  .Y({ S5595 })
);
NAND #() 
NAND_3394_ (
  .A({ S2517 }),
  .B({ S5592 }),
  .Y({ S5596 })
);
NAND #() 
NAND_3395_ (
  .A({ S5594 }),
  .B({ S5596 }),
  .Y({ S5597 })
);
NOT #() 
NOT_443_ (
  .A({ S5597 }),
  .Y({ S5598 })
);
NOR #() 
NOR_1869_ (
  .A({ S5404 }),
  .B({ S5405 }),
  .Y({ S5599 })
);
NOR #() 
NOR_1870_ (
  .A({ S5507 }),
  .B({ S5599 }),
  .Y({ S5600 })
);
NAND #() 
NAND_3396_ (
  .A({ S5507 }),
  .B({ S5599 }),
  .Y({ S5601 })
);
NOT #() 
NOT_444_ (
  .A({ S5601 }),
  .Y({ S5602 })
);
NOR #() 
NOR_1871_ (
  .A({ S5600 }),
  .B({ S5602 }),
  .Y({ S5603 })
);
NOR #() 
NOR_1872_ (
  .A({ S5539 }),
  .B({ S5603 }),
  .Y({ S5604 })
);
NOR #() 
NOR_1873_ (
  .A({ S5402 }),
  .B({ S5538 }),
  .Y({ S5605 })
);
NOR #() 
NOR_1874_ (
  .A({ S5604 }),
  .B({ S5605 }),
  .Y({ S5606 })
);
NOT #() 
NOT_445_ (
  .A({ S5606 }),
  .Y({ S5607 })
);
NOR #() 
NOR_1875_ (
  .A({ S2417 }),
  .B({ S5607 }),
  .Y({ S5608 })
);
NOR #() 
NOR_1876_ (
  .A({ S2418 }),
  .B({ S5606 }),
  .Y({ S5609 })
);
NOR #() 
NOR_1877_ (
  .A({ S5499 }),
  .B({ S5502 }),
  .Y({ S5610 })
);
NOT #() 
NOT_446_ (
  .A({ S5610 }),
  .Y({ S5611 })
);
NAND #() 
NAND_3397_ (
  .A({ S5505 }),
  .B({ S5611 }),
  .Y({ S5612 })
);
NAND #() 
NAND_3398_ (
  .A({ S5538 }),
  .B({ S5612 }),
  .Y({ S5613 })
);
NAND #() 
NAND_3399_ (
  .A({ S5411 }),
  .B({ S5539 }),
  .Y({ S5614 })
);
NAND #() 
NAND_3400_ (
  .A({ S5613 }),
  .B({ S5614 }),
  .Y({ S5615 })
);
NOT #() 
NOT_447_ (
  .A({ S5615 }),
  .Y({ S5616 })
);
NAND #() 
NAND_3401_ (
  .A({ S2312 }),
  .B({ S5616 }),
  .Y({ S5617 })
);
NOT #() 
NOT_448_ (
  .A({ S5617 }),
  .Y({ S5618 })
);
NAND #() 
NAND_3402_ (
  .A({ S2311 }),
  .B({ S5615 }),
  .Y({ S5619 })
);
NAND #() 
NAND_3403_ (
  .A({ S5617 }),
  .B({ S5619 }),
  .Y({ S5620 })
);
NOT #() 
NOT_449_ (
  .A({ S5620 }),
  .Y({ S5621 })
);
NAND #() 
NAND_3404_ (
  .A({ S5424 }),
  .B({ S5494 }),
  .Y({ S5622 })
);
NAND #() 
NAND_3405_ (
  .A({ S5497 }),
  .B({ S5622 }),
  .Y({ S5623 })
);
NAND #() 
NAND_3406_ (
  .A({ S5538 }),
  .B({ S5623 }),
  .Y({ S5624 })
);
NAND #() 
NAND_3407_ (
  .A({ S5419 }),
  .B({ S5539 }),
  .Y({ S5625 })
);
NAND #() 
NAND_3408_ (
  .A({ S5624 }),
  .B({ S5625 }),
  .Y({ S5626 })
);
NOT #() 
NOT_450_ (
  .A({ S5626 }),
  .Y({ S5627 })
);
NOR #() 
NOR_1878_ (
  .A({ S2205 }),
  .B({ S5626 }),
  .Y({ S5628 })
);
NOR #() 
NOR_1879_ (
  .A({ S2206 }),
  .B({ S5627 }),
  .Y({ S5629 })
);
NAND #() 
NAND_3409_ (
  .A({ S5435 }),
  .B({ S5490 }),
  .Y({ S5630 })
);
NAND #() 
NAND_3410_ (
  .A({ S5493 }),
  .B({ S5630 }),
  .Y({ S5631 })
);
NAND #() 
NAND_3411_ (
  .A({ S5538 }),
  .B({ S5631 }),
  .Y({ S5632 })
);
NAND #() 
NAND_3412_ (
  .A({ S5430 }),
  .B({ S5539 }),
  .Y({ S5633 })
);
NAND #() 
NAND_3413_ (
  .A({ S5632 }),
  .B({ S5633 }),
  .Y({ S5634 })
);
NOT #() 
NOT_451_ (
  .A({ S5634 }),
  .Y({ S5635 })
);
NAND #() 
NAND_3414_ (
  .A({ S2107 }),
  .B({ S5635 }),
  .Y({ S5636 })
);
NOT #() 
NOT_452_ (
  .A({ S5636 }),
  .Y({ S5637 })
);
NAND #() 
NAND_3415_ (
  .A({ S2106 }),
  .B({ S5634 }),
  .Y({ S5638 })
);
NAND #() 
NAND_3416_ (
  .A({ S5636 }),
  .B({ S5638 }),
  .Y({ S5639 })
);
NOT #() 
NOT_453_ (
  .A({ S5639 }),
  .Y({ S5640 })
);
NOR #() 
NOR_1880_ (
  .A({ S5446 }),
  .B({ S5448 }),
  .Y({ S5641 })
);
NAND #() 
NAND_3417_ (
  .A({ S5447 }),
  .B({ S5449 }),
  .Y({ S5642 })
);
NOR #() 
NOR_1881_ (
  .A({ S5486 }),
  .B({ S5642 }),
  .Y({ S5643 })
);
NOR #() 
NOR_1882_ (
  .A({ S5487 }),
  .B({ S5641 }),
  .Y({ S5644 })
);
NOR #() 
NOR_1883_ (
  .A({ S5643 }),
  .B({ S5644 }),
  .Y({ S5645 })
);
NAND #() 
NAND_3418_ (
  .A({ S5538 }),
  .B({ S5645 }),
  .Y({ S5646 })
);
NAND #() 
NAND_3419_ (
  .A({ S5444 }),
  .B({ S5539 }),
  .Y({ S5647 })
);
NAND #() 
NAND_3420_ (
  .A({ S5646 }),
  .B({ S5647 }),
  .Y({ S5648 })
);
NOT #() 
NOT_454_ (
  .A({ S5648 }),
  .Y({ S5649 })
);
NOR #() 
NOR_1884_ (
  .A({ S1597 }),
  .B({ S5649 }),
  .Y({ S5650 })
);
NAND #() 
NAND_3421_ (
  .A({ S1598 }),
  .B({ S5648 }),
  .Y({ S5651 })
);
NOR #() 
NOR_1885_ (
  .A({ S1598 }),
  .B({ S5648 }),
  .Y({ S5652 })
);
NAND #() 
NAND_3422_ (
  .A({ S1597 }),
  .B({ S5649 }),
  .Y({ S5653 })
);
NOR #() 
NOR_1886_ (
  .A({ S5462 }),
  .B({ S5483 }),
  .Y({ S5654 })
);
NAND #() 
NAND_3423_ (
  .A({ S5463 }),
  .B({ S5482 }),
  .Y({ S5655 })
);
NOR #() 
NOR_1887_ (
  .A({ S5484 }),
  .B({ S5654 }),
  .Y({ S5656 })
);
NAND #() 
NAND_3424_ (
  .A({ S5485 }),
  .B({ S5655 }),
  .Y({ S5657 })
);
NOR #() 
NOR_1888_ (
  .A({ S5539 }),
  .B({ S5656 }),
  .Y({ S5658 })
);
NAND #() 
NAND_3425_ (
  .A({ S5538 }),
  .B({ S5657 }),
  .Y({ S5659 })
);
NOR #() 
NOR_1889_ (
  .A({ S5457 }),
  .B({ S5538 }),
  .Y({ S5660 })
);
NAND #() 
NAND_3426_ (
  .A({ S5456 }),
  .B({ S5539 }),
  .Y({ S5661 })
);
NOR #() 
NOR_1890_ (
  .A({ S5658 }),
  .B({ S5660 }),
  .Y({ S5662 })
);
NAND #() 
NAND_3427_ (
  .A({ S5659 }),
  .B({ S5661 }),
  .Y({ S5663 })
);
NOR #() 
NOR_1891_ (
  .A({ S1952 }),
  .B({ S5663 }),
  .Y({ S5664 })
);
NAND #() 
NAND_3428_ (
  .A({ S1953 }),
  .B({ S5662 }),
  .Y({ S5665 })
);
NOR #() 
NOR_1892_ (
  .A({ S1953 }),
  .B({ S5662 }),
  .Y({ S5666 })
);
NAND #() 
NAND_3429_ (
  .A({ S1952 }),
  .B({ S5663 }),
  .Y({ S5667 })
);
NOR #() 
NOR_1893_ (
  .A({ S5664 }),
  .B({ S5666 }),
  .Y({ S5668 })
);
NAND #() 
NAND_3430_ (
  .A({ S5665 }),
  .B({ S5667 }),
  .Y({ S5669 })
);
NOR #() 
NOR_1894_ (
  .A({ S5475 }),
  .B({ S5478 }),
  .Y({ S5670 })
);
NAND #() 
NAND_3431_ (
  .A({ S5474 }),
  .B({ S5479 }),
  .Y({ S5671 })
);
NOR #() 
NOR_1895_ (
  .A({ S5480 }),
  .B({ S5670 }),
  .Y({ S5672 })
);
NAND #() 
NAND_3432_ (
  .A({ S5481 }),
  .B({ S5671 }),
  .Y({ S5673 })
);
NOR #() 
NOR_1896_ (
  .A({ S5539 }),
  .B({ S5672 }),
  .Y({ S5674 })
);
NAND #() 
NAND_3433_ (
  .A({ S5538 }),
  .B({ S5673 }),
  .Y({ S5675 })
);
NOR #() 
NOR_1897_ (
  .A({ S5471 }),
  .B({ S5538 }),
  .Y({ S5676 })
);
NAND #() 
NAND_3434_ (
  .A({ S5470 }),
  .B({ S5539 }),
  .Y({ S5677 })
);
NOR #() 
NOR_1898_ (
  .A({ S5674 }),
  .B({ S5676 }),
  .Y({ S5678 })
);
NAND #() 
NAND_3435_ (
  .A({ S5675 }),
  .B({ S5677 }),
  .Y({ S5679 })
);
NOR #() 
NOR_1899_ (
  .A({ S1848 }),
  .B({ S5679 }),
  .Y({ S5680 })
);
NAND #() 
NAND_3436_ (
  .A({ S1849 }),
  .B({ S5678 }),
  .Y({ S5681 })
);
NOR #() 
NOR_1900_ (
  .A({ S1849 }),
  .B({ S5678 }),
  .Y({ S5682 })
);
NAND #() 
NAND_3437_ (
  .A({ S1848 }),
  .B({ S5679 }),
  .Y({ S5683 })
);
NOR #() 
NOR_1901_ (
  .A({ S1516 }),
  .B({ S5539 }),
  .Y({ S5684 })
);
NAND #() 
NAND_3438_ (
  .A({ S1515 }),
  .B({ S5538 }),
  .Y({ S5685 })
);
NOR #() 
NOR_1902_ (
  .A({ S1116 }),
  .B({ S5684 }),
  .Y({ S5686 })
);
NAND #() 
NAND_3439_ (
  .A({ datapath_addsubunit_in1_2 }),
  .B({ S5685 }),
  .Y({ S5687 })
);
NOR #() 
NOR_1903_ (
  .A({ S5475 }),
  .B({ S5539 }),
  .Y({ S5688 })
);
NAND #() 
NAND_3440_ (
  .A({ S5474 }),
  .B({ S5538 }),
  .Y({ S5689 })
);
NOR #() 
NOR_1904_ (
  .A({ S5686 }),
  .B({ S5688 }),
  .Y({ S5690 })
);
NAND #() 
NAND_3441_ (
  .A({ S5687 }),
  .B({ S5689 }),
  .Y({ S5691 })
);
NOR #() 
NOR_1905_ (
  .A({ S1745 }),
  .B({ S5690 }),
  .Y({ S5692 })
);
NAND #() 
NAND_3442_ (
  .A({ S1746 }),
  .B({ S5691 }),
  .Y({ S5693 })
);
NOR #() 
NOR_1906_ (
  .A({ S1746 }),
  .B({ S5691 }),
  .Y({ S5694 })
);
NAND #() 
NAND_3443_ (
  .A({ S1745 }),
  .B({ S5690 }),
  .Y({ S5695 })
);
NOR #() 
NOR_1907_ (
  .A({ S5692 }),
  .B({ S5694 }),
  .Y({ S5696 })
);
NAND #() 
NAND_3444_ (
  .A({ S5693 }),
  .B({ S5695 }),
  .Y({ S5697 })
);
NAND #() 
NAND_3445_ (
  .A({ S1168 }),
  .B({ S1515 }),
  .Y({ S5698 })
);
NOT #() 
NOT_455_ (
  .A({ S5698 }),
  .Y({ S5699 })
);
NOR #() 
NOR_1908_ (
  .A({ S5697 }),
  .B({ S5699 }),
  .Y({ S5700 })
);
NAND #() 
NAND_3446_ (
  .A({ S5696 }),
  .B({ S5698 }),
  .Y({ S5701 })
);
NOR #() 
NOR_1909_ (
  .A({ S5692 }),
  .B({ S5700 }),
  .Y({ S5702 })
);
NAND #() 
NAND_3447_ (
  .A({ S5693 }),
  .B({ S5701 }),
  .Y({ S5703 })
);
NOR #() 
NOR_1910_ (
  .A({ S5682 }),
  .B({ S5702 }),
  .Y({ S5704 })
);
NAND #() 
NAND_3448_ (
  .A({ S5683 }),
  .B({ S5703 }),
  .Y({ S5705 })
);
NOR #() 
NOR_1911_ (
  .A({ S5680 }),
  .B({ S5704 }),
  .Y({ S5706 })
);
NAND #() 
NAND_3449_ (
  .A({ S5681 }),
  .B({ S5705 }),
  .Y({ S5707 })
);
NOR #() 
NOR_1912_ (
  .A({ S5669 }),
  .B({ S5706 }),
  .Y({ S5708 })
);
NAND #() 
NAND_3450_ (
  .A({ S5668 }),
  .B({ S5707 }),
  .Y({ S5709 })
);
NOR #() 
NOR_1913_ (
  .A({ S5664 }),
  .B({ S5708 }),
  .Y({ S5710 })
);
NAND #() 
NAND_3451_ (
  .A({ S5665 }),
  .B({ S5709 }),
  .Y({ S5711 })
);
NOR #() 
NOR_1914_ (
  .A({ S5652 }),
  .B({ S5710 }),
  .Y({ S5712 })
);
NAND #() 
NAND_3452_ (
  .A({ S5653 }),
  .B({ S5711 }),
  .Y({ S5713 })
);
NOR #() 
NOR_1915_ (
  .A({ S5650 }),
  .B({ S5712 }),
  .Y({ S5714 })
);
NAND #() 
NAND_3453_ (
  .A({ S5651 }),
  .B({ S5713 }),
  .Y({ S5715 })
);
NOR #() 
NOR_1916_ (
  .A({ S5639 }),
  .B({ S5714 }),
  .Y({ S5716 })
);
NAND #() 
NAND_3454_ (
  .A({ S5640 }),
  .B({ S5715 }),
  .Y({ S5717 })
);
NOR #() 
NOR_1917_ (
  .A({ S5637 }),
  .B({ S5716 }),
  .Y({ S5718 })
);
NAND #() 
NAND_3455_ (
  .A({ S5636 }),
  .B({ S5717 }),
  .Y({ S5719 })
);
NOR #() 
NOR_1918_ (
  .A({ S5629 }),
  .B({ S5718 }),
  .Y({ S5720 })
);
NOR #() 
NOR_1919_ (
  .A({ S5628 }),
  .B({ S5719 }),
  .Y({ S5721 })
);
NOR #() 
NOR_1920_ (
  .A({ S5628 }),
  .B({ S5720 }),
  .Y({ S5722 })
);
NOR #() 
NOR_1921_ (
  .A({ S5629 }),
  .B({ S5721 }),
  .Y({ S5723 })
);
NOR #() 
NOR_1922_ (
  .A({ S5620 }),
  .B({ S5722 }),
  .Y({ S5724 })
);
NAND #() 
NAND_3456_ (
  .A({ S5621 }),
  .B({ S5723 }),
  .Y({ S5725 })
);
NOR #() 
NOR_1923_ (
  .A({ S5618 }),
  .B({ S5724 }),
  .Y({ S5726 })
);
NAND #() 
NAND_3457_ (
  .A({ S5617 }),
  .B({ S5725 }),
  .Y({ S5727 })
);
NOR #() 
NOR_1924_ (
  .A({ S5609 }),
  .B({ S5726 }),
  .Y({ S5728 })
);
NOR #() 
NOR_1925_ (
  .A({ S5608 }),
  .B({ S5727 }),
  .Y({ S5729 })
);
NOR #() 
NOR_1926_ (
  .A({ S5608 }),
  .B({ S5728 }),
  .Y({ S5730 })
);
NOR #() 
NOR_1927_ (
  .A({ S5609 }),
  .B({ S5729 }),
  .Y({ S5731 })
);
NOR #() 
NOR_1928_ (
  .A({ S5597 }),
  .B({ S5730 }),
  .Y({ S5732 })
);
NAND #() 
NAND_3458_ (
  .A({ S5598 }),
  .B({ S5731 }),
  .Y({ S5733 })
);
NOR #() 
NOR_1929_ (
  .A({ S5595 }),
  .B({ S5732 }),
  .Y({ S5734 })
);
NAND #() 
NAND_3459_ (
  .A({ S5594 }),
  .B({ S5733 }),
  .Y({ S5735 })
);
NAND #() 
NAND_3460_ (
  .A({ S5587 }),
  .B({ S5735 }),
  .Y({ S5736 })
);
NAND #() 
NAND_3461_ (
  .A({ S5586 }),
  .B({ S5734 }),
  .Y({ S5737 })
);
NAND #() 
NAND_3462_ (
  .A({ S5587 }),
  .B({ S5737 }),
  .Y({ S5738 })
);
NAND #() 
NAND_3463_ (
  .A({ S5586 }),
  .B({ S5736 }),
  .Y({ S5739 })
);
NOR #() 
NOR_1930_ (
  .A({ S5572 }),
  .B({ S5738 }),
  .Y({ S5740 })
);
NAND #() 
NAND_3464_ (
  .A({ S5571 }),
  .B({ S5739 }),
  .Y({ S5741 })
);
NOR #() 
NOR_1931_ (
  .A({ S5568 }),
  .B({ S5740 }),
  .Y({ S5742 })
);
NAND #() 
NAND_3465_ (
  .A({ S5569 }),
  .B({ S5741 }),
  .Y({ S5743 })
);
NAND #() 
NAND_3466_ (
  .A({ S5561 }),
  .B({ S5743 }),
  .Y({ S5744 })
);
NAND #() 
NAND_3467_ (
  .A({ S5560 }),
  .B({ S5742 }),
  .Y({ S5745 })
);
NAND #() 
NAND_3468_ (
  .A({ S5561 }),
  .B({ S5745 }),
  .Y({ S5746 })
);
NAND #() 
NAND_3469_ (
  .A({ S5560 }),
  .B({ S5744 }),
  .Y({ S5747 })
);
NOR #() 
NOR_1932_ (
  .A({ S5549 }),
  .B({ S5746 }),
  .Y({ S5748 })
);
NAND #() 
NAND_3470_ (
  .A({ S5550 }),
  .B({ S5747 }),
  .Y({ S5749 })
);
NAND #() 
NAND_3471_ (
  .A({ S5334 }),
  .B({ S5539 }),
  .Y({ S5750 })
);
NOT #() 
NOT_456_ (
  .A({ S5750 }),
  .Y({ S5751 })
);
NOR #() 
NOR_1933_ (
  .A({ S3950 }),
  .B({ S5751 }),
  .Y({ S5752 })
);
NOR #() 
NOR_1934_ (
  .A({ S3036 }),
  .B({ S5752 }),
  .Y({ S5753 })
);
NOT #() 
NOT_457_ (
  .A({ S5753 }),
  .Y({ S5754 })
);
NOR #() 
NOR_1935_ (
  .A({ S5547 }),
  .B({ S5753 }),
  .Y({ S5755 })
);
NAND #() 
NAND_3472_ (
  .A({ S5546 }),
  .B({ S5754 }),
  .Y({ S5756 })
);
NOR #() 
NOR_1936_ (
  .A({ S5748 }),
  .B({ S5756 }),
  .Y({ S5757 })
);
NAND #() 
NAND_3473_ (
  .A({ S5749 }),
  .B({ S5755 }),
  .Y({ S5758 })
);
NAND #() 
NAND_3474_ (
  .A({ S3036 }),
  .B({ S5752 }),
  .Y({ S5759 })
);
NAND #() 
NAND_3475_ (
  .A({ S3142 }),
  .B({ S5759 }),
  .Y({ S5760 })
);
NOT #() 
NOT_458_ (
  .A({ S5760 }),
  .Y({ S5761 })
);
NOR #() 
NOR_1937_ (
  .A({ S5757 }),
  .B({ S5760 }),
  .Y({ S5762 })
);
NAND #() 
NAND_3476_ (
  .A({ S5758 }),
  .B({ S5761 }),
  .Y({ S5763 })
);
NAND #() 
NAND_3477_ (
  .A({ S5639 }),
  .B({ S5714 }),
  .Y({ S5764 })
);
NAND #() 
NAND_3478_ (
  .A({ S5717 }),
  .B({ S5764 }),
  .Y({ S5765 })
);
NAND #() 
NAND_3479_ (
  .A({ S5762 }),
  .B({ S5765 }),
  .Y({ S5766 })
);
NAND #() 
NAND_3480_ (
  .A({ S5634 }),
  .B({ S5763 }),
  .Y({ S5767 })
);
NAND #() 
NAND_3481_ (
  .A({ S5766 }),
  .B({ S5767 }),
  .Y({ S5768 })
);
NAND #() 
NAND_3482_ (
  .A({ S2205 }),
  .B({ S5768 }),
  .Y({ S5769 })
);
NOR #() 
NOR_1938_ (
  .A({ S5650 }),
  .B({ S5652 }),
  .Y({ S5770 })
);
NAND #() 
NAND_3483_ (
  .A({ S5651 }),
  .B({ S5653 }),
  .Y({ S5771 })
);
NOR #() 
NOR_1939_ (
  .A({ S5710 }),
  .B({ S5771 }),
  .Y({ S5772 })
);
NOR #() 
NOR_1940_ (
  .A({ S5711 }),
  .B({ S5770 }),
  .Y({ S5773 })
);
NOR #() 
NOR_1941_ (
  .A({ S5772 }),
  .B({ S5773 }),
  .Y({ S5774 })
);
NAND #() 
NAND_3484_ (
  .A({ S5762 }),
  .B({ S5774 }),
  .Y({ S5775 })
);
NAND #() 
NAND_3485_ (
  .A({ S5648 }),
  .B({ S5763 }),
  .Y({ S5776 })
);
NAND #() 
NAND_3486_ (
  .A({ S5775 }),
  .B({ S5776 }),
  .Y({ S5777 })
);
NAND #() 
NAND_3487_ (
  .A({ S2107 }),
  .B({ S5777 }),
  .Y({ S5778 })
);
NOR #() 
NOR_1942_ (
  .A({ S5696 }),
  .B({ S5698 }),
  .Y({ S5779 })
);
NOR #() 
NOR_1943_ (
  .A({ S5700 }),
  .B({ S5779 }),
  .Y({ S5780 })
);
NOR #() 
NOR_1944_ (
  .A({ S5763 }),
  .B({ S5780 }),
  .Y({ S5781 })
);
NOR #() 
NOR_1945_ (
  .A({ S5691 }),
  .B({ S5762 }),
  .Y({ S5782 })
);
NOR #() 
NOR_1946_ (
  .A({ S5781 }),
  .B({ S5782 }),
  .Y({ S5783 })
);
NAND #() 
NAND_3488_ (
  .A({ S1849 }),
  .B({ S5783 }),
  .Y({ S5784 })
);
NAND #() 
NAND_3489_ (
  .A({ S1515 }),
  .B({ S5762 }),
  .Y({ S5785 })
);
NAND #() 
NAND_3490_ (
  .A({ datapath_addsubunit_in1_1 }),
  .B({ S5785 }),
  .Y({ S5786 })
);
NOR #() 
NOR_1947_ (
  .A({ datapath_addsubunit_in1_0 }),
  .B({ S1516 }),
  .Y({ S5787 })
);
NOR #() 
NOR_1948_ (
  .A({ S1745 }),
  .B({ S5787 }),
  .Y({ S5788 })
);
NOR #() 
NOR_1949_ (
  .A({ S5698 }),
  .B({ S5763 }),
  .Y({ S5789 })
);
NOR #() 
NOR_1950_ (
  .A({ S5788 }),
  .B({ S5789 }),
  .Y({ S5790 })
);
NAND #() 
NAND_3491_ (
  .A({ S5786 }),
  .B({ S5790 }),
  .Y({ S5791 })
);
NAND #() 
NAND_3492_ (
  .A({ S1745 }),
  .B({ S5787 }),
  .Y({ S5792 })
);
NAND #() 
NAND_3493_ (
  .A({ S5791 }),
  .B({ S5792 }),
  .Y({ S5793 })
);
NAND #() 
NAND_3494_ (
  .A({ S5784 }),
  .B({ S5793 }),
  .Y({ S5794 })
);
NOR #() 
NOR_1951_ (
  .A({ S5680 }),
  .B({ S5682 }),
  .Y({ S5795 })
);
NAND #() 
NAND_3495_ (
  .A({ S5681 }),
  .B({ S5683 }),
  .Y({ S5796 })
);
NAND #() 
NAND_3496_ (
  .A({ S5702 }),
  .B({ S5795 }),
  .Y({ S5797 })
);
NAND #() 
NAND_3497_ (
  .A({ S5703 }),
  .B({ S5796 }),
  .Y({ S5798 })
);
NAND #() 
NAND_3498_ (
  .A({ S5797 }),
  .B({ S5798 }),
  .Y({ S5799 })
);
NAND #() 
NAND_3499_ (
  .A({ S5762 }),
  .B({ S5799 }),
  .Y({ S5800 })
);
NOT #() 
NOT_459_ (
  .A({ S5800 }),
  .Y({ S5801 })
);
NOR #() 
NOR_1952_ (
  .A({ S5679 }),
  .B({ S5762 }),
  .Y({ S5802 })
);
NAND #() 
NAND_3500_ (
  .A({ S5678 }),
  .B({ S5763 }),
  .Y({ S5803 })
);
NOR #() 
NOR_1953_ (
  .A({ S5801 }),
  .B({ S5802 }),
  .Y({ S5804 })
);
NAND #() 
NAND_3501_ (
  .A({ S5800 }),
  .B({ S5803 }),
  .Y({ S5805 })
);
NOR #() 
NOR_1954_ (
  .A({ S1953 }),
  .B({ S5805 }),
  .Y({ S5806 })
);
NOR #() 
NOR_1955_ (
  .A({ S1849 }),
  .B({ S5783 }),
  .Y({ S5807 })
);
NOR #() 
NOR_1956_ (
  .A({ S5806 }),
  .B({ S5807 }),
  .Y({ S5808 })
);
NAND #() 
NAND_3502_ (
  .A({ S5794 }),
  .B({ S5808 }),
  .Y({ S5809 })
);
NOR #() 
NOR_1957_ (
  .A({ S1952 }),
  .B({ S5804 }),
  .Y({ S5810 })
);
NAND #() 
NAND_3503_ (
  .A({ S5669 }),
  .B({ S5706 }),
  .Y({ S5811 })
);
NAND #() 
NAND_3504_ (
  .A({ S5709 }),
  .B({ S5811 }),
  .Y({ S5812 })
);
NAND #() 
NAND_3505_ (
  .A({ S5762 }),
  .B({ S5812 }),
  .Y({ S5813 })
);
NOT #() 
NOT_460_ (
  .A({ S5813 }),
  .Y({ S5814 })
);
NOR #() 
NOR_1958_ (
  .A({ S5662 }),
  .B({ S5762 }),
  .Y({ S5815 })
);
NOT #() 
NOT_461_ (
  .A({ S5815 }),
  .Y({ S5816 })
);
NOR #() 
NOR_1959_ (
  .A({ S5814 }),
  .B({ S5815 }),
  .Y({ S5817 })
);
NAND #() 
NAND_3506_ (
  .A({ S5813 }),
  .B({ S5816 }),
  .Y({ S5818 })
);
NOR #() 
NOR_1960_ (
  .A({ S1597 }),
  .B({ S5818 }),
  .Y({ S5819 })
);
NOR #() 
NOR_1961_ (
  .A({ S5810 }),
  .B({ S5819 }),
  .Y({ S5820 })
);
NAND #() 
NAND_3507_ (
  .A({ S5809 }),
  .B({ S5820 }),
  .Y({ S5821 })
);
NOR #() 
NOR_1962_ (
  .A({ S2107 }),
  .B({ S5777 }),
  .Y({ S5822 })
);
NOR #() 
NOR_1963_ (
  .A({ S1598 }),
  .B({ S5817 }),
  .Y({ S5823 })
);
NOR #() 
NOR_1964_ (
  .A({ S5822 }),
  .B({ S5823 }),
  .Y({ S5824 })
);
NAND #() 
NAND_3508_ (
  .A({ S5821 }),
  .B({ S5824 }),
  .Y({ S5825 })
);
NAND #() 
NAND_3509_ (
  .A({ S5778 }),
  .B({ S5825 }),
  .Y({ S5826 })
);
NAND #() 
NAND_3510_ (
  .A({ S5769 }),
  .B({ S5826 }),
  .Y({ S5827 })
);
NOR #() 
NOR_1965_ (
  .A({ S5628 }),
  .B({ S5629 }),
  .Y({ S5828 })
);
NOR #() 
NOR_1966_ (
  .A({ S5719 }),
  .B({ S5828 }),
  .Y({ S5829 })
);
NAND #() 
NAND_3511_ (
  .A({ S5719 }),
  .B({ S5828 }),
  .Y({ S5830 })
);
NOT #() 
NOT_462_ (
  .A({ S5830 }),
  .Y({ S5831 })
);
NOR #() 
NOR_1967_ (
  .A({ S5829 }),
  .B({ S5831 }),
  .Y({ S5832 })
);
NOR #() 
NOR_1968_ (
  .A({ S5626 }),
  .B({ S5762 }),
  .Y({ S5833 })
);
NAND #() 
NAND_3512_ (
  .A({ S5762 }),
  .B({ S5832 }),
  .Y({ S5834 })
);
NOT #() 
NOT_463_ (
  .A({ S5834 }),
  .Y({ S5835 })
);
NOR #() 
NOR_1969_ (
  .A({ S5833 }),
  .B({ S5835 }),
  .Y({ S5836 })
);
NOR #() 
NOR_1970_ (
  .A({ S2311 }),
  .B({ S5836 }),
  .Y({ S5837 })
);
NOR #() 
NOR_1971_ (
  .A({ S2205 }),
  .B({ S5768 }),
  .Y({ S5838 })
);
NOR #() 
NOR_1972_ (
  .A({ S5837 }),
  .B({ S5838 }),
  .Y({ S5839 })
);
NAND #() 
NAND_3513_ (
  .A({ S5827 }),
  .B({ S5839 }),
  .Y({ S5840 })
);
NAND #() 
NAND_3514_ (
  .A({ S5597 }),
  .B({ S5730 }),
  .Y({ S5841 })
);
NAND #() 
NAND_3515_ (
  .A({ S5733 }),
  .B({ S5841 }),
  .Y({ S5842 })
);
NAND #() 
NAND_3516_ (
  .A({ S5762 }),
  .B({ S5842 }),
  .Y({ S5843 })
);
NAND #() 
NAND_3517_ (
  .A({ S5592 }),
  .B({ S5763 }),
  .Y({ S5844 })
);
NAND #() 
NAND_3518_ (
  .A({ S5843 }),
  .B({ S5844 }),
  .Y({ S5845 })
);
NOR #() 
NOR_1973_ (
  .A({ S2617 }),
  .B({ S5845 }),
  .Y({ S5846 })
);
NAND #() 
NAND_3519_ (
  .A({ S5586 }),
  .B({ S5587 }),
  .Y({ S5847 })
);
NAND #() 
NAND_3520_ (
  .A({ S5735 }),
  .B({ S5847 }),
  .Y({ S5848 })
);
NOT #() 
NOT_464_ (
  .A({ S5848 }),
  .Y({ S5849 })
);
NOR #() 
NOR_1974_ (
  .A({ S5735 }),
  .B({ S5847 }),
  .Y({ S5850 })
);
NOR #() 
NOR_1975_ (
  .A({ S5849 }),
  .B({ S5850 }),
  .Y({ S5851 })
);
NAND #() 
NAND_3521_ (
  .A({ S5762 }),
  .B({ S5851 }),
  .Y({ S5852 })
);
NOT #() 
NOT_465_ (
  .A({ S5852 }),
  .Y({ S5853 })
);
NOR #() 
NOR_1976_ (
  .A({ S5584 }),
  .B({ S5762 }),
  .Y({ S5854 })
);
NOT #() 
NOT_466_ (
  .A({ S5854 }),
  .Y({ S5855 })
);
NOR #() 
NOR_1977_ (
  .A({ S5853 }),
  .B({ S5854 }),
  .Y({ S5856 })
);
NAND #() 
NAND_3522_ (
  .A({ S5852 }),
  .B({ S5855 }),
  .Y({ S5857 })
);
NOR #() 
NOR_1978_ (
  .A({ S2717 }),
  .B({ S5857 }),
  .Y({ S5858 })
);
NOR #() 
NOR_1979_ (
  .A({ S5846 }),
  .B({ S5858 }),
  .Y({ S5859 })
);
NOT #() 
NOT_467_ (
  .A({ S5859 }),
  .Y({ S5860 })
);
NAND #() 
NAND_3523_ (
  .A({ S2617 }),
  .B({ S5845 }),
  .Y({ S5861 })
);
NOR #() 
NOR_1980_ (
  .A({ S2718 }),
  .B({ S5856 }),
  .Y({ S5862 })
);
NAND #() 
NAND_3524_ (
  .A({ S2717 }),
  .B({ S5857 }),
  .Y({ S5863 })
);
NAND #() 
NAND_3525_ (
  .A({ S5861 }),
  .B({ S5863 }),
  .Y({ S5864 })
);
NOR #() 
NOR_1981_ (
  .A({ S5860 }),
  .B({ S5864 }),
  .Y({ S5865 })
);
NAND #() 
NAND_3526_ (
  .A({ S5620 }),
  .B({ S5722 }),
  .Y({ S5866 })
);
NAND #() 
NAND_3527_ (
  .A({ S5725 }),
  .B({ S5866 }),
  .Y({ S5867 })
);
NAND #() 
NAND_3528_ (
  .A({ S5762 }),
  .B({ S5867 }),
  .Y({ S5868 })
);
NAND #() 
NAND_3529_ (
  .A({ S5615 }),
  .B({ S5763 }),
  .Y({ S5869 })
);
NAND #() 
NAND_3530_ (
  .A({ S5868 }),
  .B({ S5869 }),
  .Y({ S5870 })
);
NOT #() 
NOT_468_ (
  .A({ S5870 }),
  .Y({ S5871 })
);
NOR #() 
NOR_1982_ (
  .A({ S2417 }),
  .B({ S5870 }),
  .Y({ S5872 })
);
NAND #() 
NAND_3531_ (
  .A({ S2418 }),
  .B({ S5871 }),
  .Y({ S5873 })
);
NAND #() 
NAND_3532_ (
  .A({ S2311 }),
  .B({ S5836 }),
  .Y({ S5874 })
);
NOR #() 
NOR_1983_ (
  .A({ S5608 }),
  .B({ S5609 }),
  .Y({ S5875 })
);
NOR #() 
NOR_1984_ (
  .A({ S5727 }),
  .B({ S5875 }),
  .Y({ S5876 })
);
NOT #() 
NOT_469_ (
  .A({ S5876 }),
  .Y({ S5877 })
);
NAND #() 
NAND_3533_ (
  .A({ S5727 }),
  .B({ S5875 }),
  .Y({ S5878 })
);
NAND #() 
NAND_3534_ (
  .A({ S5877 }),
  .B({ S5878 }),
  .Y({ S5879 })
);
NAND #() 
NAND_3535_ (
  .A({ S5762 }),
  .B({ S5879 }),
  .Y({ S5880 })
);
NOT #() 
NOT_470_ (
  .A({ S5880 }),
  .Y({ S5881 })
);
NOR #() 
NOR_1985_ (
  .A({ S5606 }),
  .B({ S5762 }),
  .Y({ S5882 })
);
NOR #() 
NOR_1986_ (
  .A({ S5881 }),
  .B({ S5882 }),
  .Y({ S5883 })
);
NOT #() 
NOT_471_ (
  .A({ S5883 }),
  .Y({ S5884 })
);
NAND #() 
NAND_3536_ (
  .A({ S2518 }),
  .B({ S5883 }),
  .Y({ S5885 })
);
NOR #() 
NOR_1987_ (
  .A({ S2518 }),
  .B({ S5883 }),
  .Y({ S5886 })
);
NAND #() 
NAND_3537_ (
  .A({ S2517 }),
  .B({ S5884 }),
  .Y({ S5887 })
);
NAND #() 
NAND_3538_ (
  .A({ S2417 }),
  .B({ S5870 }),
  .Y({ S5888 })
);
NAND #() 
NAND_3539_ (
  .A({ S5874 }),
  .B({ S5887 }),
  .Y({ S5889 })
);
NAND #() 
NAND_3540_ (
  .A({ S5885 }),
  .B({ S5888 }),
  .Y({ S5890 })
);
NOR #() 
NOR_1988_ (
  .A({ S5889 }),
  .B({ S5890 }),
  .Y({ S5891 })
);
NAND #() 
NAND_3541_ (
  .A({ S5865 }),
  .B({ S5891 }),
  .Y({ S5892 })
);
NOR #() 
NOR_1989_ (
  .A({ S5872 }),
  .B({ S5892 }),
  .Y({ S5893 })
);
NAND #() 
NAND_3542_ (
  .A({ S5840 }),
  .B({ S5893 }),
  .Y({ S5894 })
);
NAND #() 
NAND_3543_ (
  .A({ S5873 }),
  .B({ S5885 }),
  .Y({ S5895 })
);
NAND #() 
NAND_3544_ (
  .A({ S5865 }),
  .B({ S5895 }),
  .Y({ S5896 })
);
NOR #() 
NOR_1990_ (
  .A({ S5886 }),
  .B({ S5896 }),
  .Y({ S5897 })
);
NOR #() 
NOR_1991_ (
  .A({ S5859 }),
  .B({ S5862 }),
  .Y({ S5898 })
);
NOR #() 
NOR_1992_ (
  .A({ S5897 }),
  .B({ S5898 }),
  .Y({ S5899 })
);
NAND #() 
NAND_3545_ (
  .A({ S5894 }),
  .B({ S5899 }),
  .Y({ S5900 })
);
NOR #() 
NOR_1993_ (
  .A({ S5752 }),
  .B({ S5762 }),
  .Y({ S5901 })
);
NOT #() 
NOT_472_ (
  .A({ S5901 }),
  .Y({ S5902 })
);
NAND #() 
NAND_3546_ (
  .A({ S5121 }),
  .B({ S5902 }),
  .Y({ S5903 })
);
NAND #() 
NAND_3547_ (
  .A({ S3142 }),
  .B({ S5903 }),
  .Y({ S5904 })
);
NAND #() 
NAND_3548_ (
  .A({ S5549 }),
  .B({ S5746 }),
  .Y({ S5905 })
);
NAND #() 
NAND_3549_ (
  .A({ S5749 }),
  .B({ S5905 }),
  .Y({ S5906 })
);
NAND #() 
NAND_3550_ (
  .A({ S5762 }),
  .B({ S5906 }),
  .Y({ S5907 })
);
NAND #() 
NAND_3551_ (
  .A({ S5544 }),
  .B({ S5763 }),
  .Y({ S5908 })
);
NAND #() 
NAND_3552_ (
  .A({ S5907 }),
  .B({ S5908 }),
  .Y({ S5909 })
);
NOR #() 
NOR_1994_ (
  .A({ S3036 }),
  .B({ S5909 }),
  .Y({ S5910 })
);
NOT #() 
NOT_473_ (
  .A({ S5910 }),
  .Y({ S5911 })
);
NAND #() 
NAND_3553_ (
  .A({ S5904 }),
  .B({ S5911 }),
  .Y({ S5912 })
);
NOR #() 
NOR_1995_ (
  .A({ S3142 }),
  .B({ S5903 }),
  .Y({ S5913 })
);
NOT #() 
NOT_474_ (
  .A({ S5913 }),
  .Y({ S5914 })
);
NAND #() 
NAND_3554_ (
  .A({ S3036 }),
  .B({ S5909 }),
  .Y({ S5915 })
);
NAND #() 
NAND_3555_ (
  .A({ S5914 }),
  .B({ S5915 }),
  .Y({ S5916 })
);
NOR #() 
NOR_1996_ (
  .A({ S5912 }),
  .B({ S5916 }),
  .Y({ S5917 })
);
NOR #() 
NOR_1997_ (
  .A({ S5571 }),
  .B({ S5739 }),
  .Y({ S5918 })
);
NOR #() 
NOR_1998_ (
  .A({ S5740 }),
  .B({ S5918 }),
  .Y({ S5919 })
);
NOR #() 
NOR_1999_ (
  .A({ S5763 }),
  .B({ S5919 }),
  .Y({ S5920 })
);
NOR #() 
NOR_2000_ (
  .A({ S5566 }),
  .B({ S5762 }),
  .Y({ S5921 })
);
NOR #() 
NOR_2001_ (
  .A({ S5920 }),
  .B({ S5921 }),
  .Y({ S5922 })
);
NAND #() 
NAND_3556_ (
  .A({ S2817 }),
  .B({ S5922 }),
  .Y({ S5923 })
);
NAND #() 
NAND_3557_ (
  .A({ S5560 }),
  .B({ S5561 }),
  .Y({ S5924 })
);
NAND #() 
NAND_3558_ (
  .A({ S5742 }),
  .B({ S5924 }),
  .Y({ S5925 })
);
NOR #() 
NOR_2002_ (
  .A({ S5742 }),
  .B({ S5924 }),
  .Y({ S5926 })
);
NOT #() 
NOT_475_ (
  .A({ S5926 }),
  .Y({ S5927 })
);
NAND #() 
NAND_3559_ (
  .A({ S5925 }),
  .B({ S5927 }),
  .Y({ S5928 })
);
NAND #() 
NAND_3560_ (
  .A({ S5762 }),
  .B({ S5928 }),
  .Y({ S5929 })
);
NOT #() 
NOT_476_ (
  .A({ S5929 }),
  .Y({ S5930 })
);
NOR #() 
NOR_2003_ (
  .A({ S5558 }),
  .B({ S5762 }),
  .Y({ S5931 })
);
NOR #() 
NOR_2004_ (
  .A({ S5930 }),
  .B({ S5931 }),
  .Y({ S5932 })
);
NAND #() 
NAND_3561_ (
  .A({ S2920 }),
  .B({ S5932 }),
  .Y({ S5933 })
);
NAND #() 
NAND_3562_ (
  .A({ S5923 }),
  .B({ S5933 }),
  .Y({ S5934 })
);
NOR #() 
NOR_2005_ (
  .A({ S2817 }),
  .B({ S5922 }),
  .Y({ S5935 })
);
NOR #() 
NOR_2006_ (
  .A({ S2920 }),
  .B({ S5932 }),
  .Y({ S5936 })
);
NOR #() 
NOR_2007_ (
  .A({ S5934 }),
  .B({ S5936 }),
  .Y({ S5937 })
);
NAND #() 
NAND_3563_ (
  .A({ S5917 }),
  .B({ S5937 }),
  .Y({ S5938 })
);
NOR #() 
NOR_2008_ (
  .A({ S5935 }),
  .B({ S5938 }),
  .Y({ S5939 })
);
NAND #() 
NAND_3564_ (
  .A({ S5900 }),
  .B({ S5939 }),
  .Y({ S5940 })
);
NAND #() 
NAND_3565_ (
  .A({ S5910 }),
  .B({ S5914 }),
  .Y({ S5941 })
);
NAND #() 
NAND_3566_ (
  .A({ S5904 }),
  .B({ S5941 }),
  .Y({ S5942 })
);
NAND #() 
NAND_3567_ (
  .A({ S5917 }),
  .B({ S5934 }),
  .Y({ S5943 })
);
NOR #() 
NOR_2009_ (
  .A({ S5936 }),
  .B({ S5943 }),
  .Y({ S5944 })
);
NOR #() 
NOR_2010_ (
  .A({ S5942 }),
  .B({ S5944 }),
  .Y({ S5945 })
);
NAND #() 
NAND_3568_ (
  .A({ S5940 }),
  .B({ S5945 }),
  .Y({ S5946 })
);
NAND #() 
NAND_3569_ (
  .A({ S3898 }),
  .B({ S5946 }),
  .Y({ S5947 })
);
NOR #() 
NOR_2011_ (
  .A({ S377 }),
  .B({ S1392 }),
  .Y({ S5948 })
);
NAND #() 
NAND_3570_ (
  .A({ S376 }),
  .B({ S1391 }),
  .Y({ S5949 })
);
NAND #() 
NAND_3571_ (
  .A({ S8564 }),
  .B({ S376 }),
  .Y({ S5950 })
);
NAND #() 
NAND_3572_ (
  .A({ datapath_multdivunit_outmdu1_0 }),
  .B({ S5950 }),
  .Y({ S5951 })
);
NOT #() 
NOT_477_ (
  .A({ S5951 }),
  .Y({ S5952 })
);
NAND #() 
NAND_3573_ (
  .A({ S1515 }),
  .B({ S5948 }),
  .Y({ S5953 })
);
NOR #() 
NOR_2012_ (
  .A({ S1220 }),
  .B({ S5953 }),
  .Y({ S5954 })
);
NOR #() 
NOR_2013_ (
  .A({ S5952 }),
  .B({ S5954 }),
  .Y({ S5955 })
);
NAND #() 
NAND_3574_ (
  .A({ S5947 }),
  .B({ S5955 }),
  .Y({ S282 })
);
NAND #() 
NAND_3575_ (
  .A({ S3898 }),
  .B({ S5762 }),
  .Y({ S5956 })
);
NOR #() 
NOR_2014_ (
  .A({ S1168 }),
  .B({ S1516 }),
  .Y({ S5957 })
);
NAND #() 
NAND_3576_ (
  .A({ datapath_addsubunit_in1_0 }),
  .B({ S1745 }),
  .Y({ S5958 })
);
NOT #() 
NOT_478_ (
  .A({ S5958 }),
  .Y({ S5959 })
);
NAND #() 
NAND_3577_ (
  .A({ datapath_addsubunit_in1_1 }),
  .B({ S1745 }),
  .Y({ S5960 })
);
NAND #() 
NAND_3578_ (
  .A({ S5957 }),
  .B({ S5959 }),
  .Y({ S5961 })
);
NOR #() 
NOR_2015_ (
  .A({ S5957 }),
  .B({ S5959 }),
  .Y({ S5962 })
);
NAND #() 
NAND_3579_ (
  .A({ S5948 }),
  .B({ S5961 }),
  .Y({ S5963 })
);
NOR #() 
NOR_2016_ (
  .A({ S5962 }),
  .B({ S5963 }),
  .Y({ S5964 })
);
NAND #() 
NAND_3580_ (
  .A({ datapath_multdivunit_outmdu1_1 }),
  .B({ S5950 }),
  .Y({ S5965 })
);
NOT #() 
NOT_479_ (
  .A({ S5965 }),
  .Y({ S5966 })
);
NOR #() 
NOR_2017_ (
  .A({ S5964 }),
  .B({ S5966 }),
  .Y({ S5967 })
);
NAND #() 
NAND_3581_ (
  .A({ S5956 }),
  .B({ S5967 }),
  .Y({ S283 })
);
NOR #() 
NOR_2018_ (
  .A({ S3899 }),
  .B({ S5539 }),
  .Y({ S5968 })
);
NAND #() 
NAND_3582_ (
  .A({ datapath_multdivunit_outmdu1_2 }),
  .B({ S5950 }),
  .Y({ S5969 })
);
NAND #() 
NAND_3583_ (
  .A({ datapath_addsubunit_in1_0 }),
  .B({ S1848 }),
  .Y({ S5970 })
);
NOT #() 
NOT_480_ (
  .A({ S5970 }),
  .Y({ S5971 })
);
NAND #() 
NAND_3584_ (
  .A({ datapath_addsubunit_in1_2 }),
  .B({ S1515 }),
  .Y({ S5972 })
);
NAND #() 
NAND_3585_ (
  .A({ S5960 }),
  .B({ S5972 }),
  .Y({ S5973 })
);
NOR #() 
NOR_2019_ (
  .A({ S1116 }),
  .B({ S1746 }),
  .Y({ S5974 })
);
NAND #() 
NAND_3586_ (
  .A({ datapath_addsubunit_in1_2 }),
  .B({ S1745 }),
  .Y({ S5975 })
);
NAND #() 
NAND_3587_ (
  .A({ S5957 }),
  .B({ S5974 }),
  .Y({ S5976 })
);
NOT #() 
NOT_481_ (
  .A({ S5976 }),
  .Y({ S5977 })
);
NAND #() 
NAND_3588_ (
  .A({ S5973 }),
  .B({ S5976 }),
  .Y({ S5978 })
);
NOT #() 
NOT_482_ (
  .A({ S5978 }),
  .Y({ S5979 })
);
NAND #() 
NAND_3589_ (
  .A({ S5971 }),
  .B({ S5979 }),
  .Y({ S5980 })
);
NOT #() 
NOT_483_ (
  .A({ S5980 }),
  .Y({ S5981 })
);
NAND #() 
NAND_3590_ (
  .A({ S5970 }),
  .B({ S5978 }),
  .Y({ S5982 })
);
NAND #() 
NAND_3591_ (
  .A({ S5980 }),
  .B({ S5982 }),
  .Y({ S5983 })
);
NOR #() 
NOR_2020_ (
  .A({ S5961 }),
  .B({ S5983 }),
  .Y({ S5984 })
);
NAND #() 
NAND_3592_ (
  .A({ S5961 }),
  .B({ S5983 }),
  .Y({ S5985 })
);
NAND #() 
NAND_3593_ (
  .A({ S5948 }),
  .B({ S5985 }),
  .Y({ S5986 })
);
NOR #() 
NOR_2021_ (
  .A({ S5984 }),
  .B({ S5986 }),
  .Y({ S5987 })
);
NOR #() 
NOR_2022_ (
  .A({ S5968 }),
  .B({ S5987 }),
  .Y({ S5988 })
);
NAND #() 
NAND_3594_ (
  .A({ S5969 }),
  .B({ S5988 }),
  .Y({ S284 })
);
NOR #() 
NOR_2023_ (
  .A({ S3899 }),
  .B({ S5333 }),
  .Y({ S5989 })
);
NAND #() 
NAND_3595_ (
  .A({ datapath_multdivunit_outmdu1_3 }),
  .B({ S5950 }),
  .Y({ S5990 })
);
NOR #() 
NOR_2024_ (
  .A({ S1220 }),
  .B({ S1953 }),
  .Y({ S5991 })
);
NAND #() 
NAND_3596_ (
  .A({ datapath_addsubunit_in1_0 }),
  .B({ S1952 }),
  .Y({ S5992 })
);
NOR #() 
NOR_2025_ (
  .A({ S5977 }),
  .B({ S5981 }),
  .Y({ S5993 })
);
NOR #() 
NOR_2026_ (
  .A({ S1168 }),
  .B({ S1849 }),
  .Y({ S5994 })
);
NAND #() 
NAND_3597_ (
  .A({ datapath_addsubunit_in1_1 }),
  .B({ S1848 }),
  .Y({ S5995 })
);
NOR #() 
NOR_2027_ (
  .A({ S1065 }),
  .B({ S1516 }),
  .Y({ S5996 })
);
NAND #() 
NAND_3598_ (
  .A({ datapath_addsubunit_in1_3 }),
  .B({ S1515 }),
  .Y({ S5997 })
);
NOR #() 
NOR_2028_ (
  .A({ S5974 }),
  .B({ S5996 }),
  .Y({ S5998 })
);
NAND #() 
NAND_3599_ (
  .A({ S5975 }),
  .B({ S5997 }),
  .Y({ S5999 })
);
NOR #() 
NOR_2029_ (
  .A({ S1065 }),
  .B({ S1746 }),
  .Y({ S6000 })
);
NAND #() 
NAND_3600_ (
  .A({ datapath_addsubunit_in1_3 }),
  .B({ S1745 }),
  .Y({ S6001 })
);
NOR #() 
NOR_2030_ (
  .A({ S5975 }),
  .B({ S5997 }),
  .Y({ S6002 })
);
NAND #() 
NAND_3601_ (
  .A({ S5974 }),
  .B({ S5996 }),
  .Y({ S6003 })
);
NOR #() 
NOR_2031_ (
  .A({ S5998 }),
  .B({ S6002 }),
  .Y({ S6004 })
);
NAND #() 
NAND_3602_ (
  .A({ S5999 }),
  .B({ S6003 }),
  .Y({ S6005 })
);
NOR #() 
NOR_2032_ (
  .A({ S5995 }),
  .B({ S6005 }),
  .Y({ S6006 })
);
NAND #() 
NAND_3603_ (
  .A({ S5994 }),
  .B({ S6004 }),
  .Y({ S6007 })
);
NAND #() 
NAND_3604_ (
  .A({ S5995 }),
  .B({ S6005 }),
  .Y({ S6008 })
);
NAND #() 
NAND_3605_ (
  .A({ S6007 }),
  .B({ S6008 }),
  .Y({ S6009 })
);
NOR #() 
NOR_2033_ (
  .A({ S5993 }),
  .B({ S6009 }),
  .Y({ S6010 })
);
NOT #() 
NOT_484_ (
  .A({ S6010 }),
  .Y({ S6011 })
);
NAND #() 
NAND_3606_ (
  .A({ S5993 }),
  .B({ S6009 }),
  .Y({ S6012 })
);
NAND #() 
NAND_3607_ (
  .A({ S6011 }),
  .B({ S6012 }),
  .Y({ S6013 })
);
NOT #() 
NOT_485_ (
  .A({ S6013 }),
  .Y({ S6014 })
);
NAND #() 
NAND_3608_ (
  .A({ S5991 }),
  .B({ S6014 }),
  .Y({ S6015 })
);
NOT #() 
NOT_486_ (
  .A({ S6015 }),
  .Y({ S6016 })
);
NAND #() 
NAND_3609_ (
  .A({ S5992 }),
  .B({ S6013 }),
  .Y({ S6017 })
);
NOT #() 
NOT_487_ (
  .A({ S6017 }),
  .Y({ S6018 })
);
NOR #() 
NOR_2034_ (
  .A({ S6016 }),
  .B({ S6018 }),
  .Y({ S6019 })
);
NAND #() 
NAND_3610_ (
  .A({ S5984 }),
  .B({ S6019 }),
  .Y({ S6020 })
);
NOR #() 
NOR_2035_ (
  .A({ S5984 }),
  .B({ S6019 }),
  .Y({ S6021 })
);
NAND #() 
NAND_3611_ (
  .A({ S5948 }),
  .B({ S6020 }),
  .Y({ S6022 })
);
NOR #() 
NOR_2036_ (
  .A({ S6021 }),
  .B({ S6022 }),
  .Y({ S6023 })
);
NOR #() 
NOR_2037_ (
  .A({ S5989 }),
  .B({ S6023 }),
  .Y({ S6024 })
);
NAND #() 
NAND_3612_ (
  .A({ S5990 }),
  .B({ S6024 }),
  .Y({ S285 })
);
NOR #() 
NOR_2038_ (
  .A({ S3899 }),
  .B({ S5113 }),
  .Y({ S6025 })
);
NOR #() 
NOR_2039_ (
  .A({ S6010 }),
  .B({ S6016 }),
  .Y({ S6026 })
);
NAND #() 
NAND_3613_ (
  .A({ datapath_addsubunit_in1_0 }),
  .B({ S1597 }),
  .Y({ S6027 })
);
NAND #() 
NAND_3614_ (
  .A({ datapath_addsubunit_in1_1 }),
  .B({ S1952 }),
  .Y({ S6028 })
);
NAND #() 
NAND_3615_ (
  .A({ S6027 }),
  .B({ S6028 }),
  .Y({ S6029 })
);
NOR #() 
NOR_2040_ (
  .A({ S1168 }),
  .B({ S1598 }),
  .Y({ S6030 })
);
NAND #() 
NAND_3616_ (
  .A({ datapath_addsubunit_in1_1 }),
  .B({ S1597 }),
  .Y({ S6031 })
);
NOR #() 
NOR_2041_ (
  .A({ S5992 }),
  .B({ S6031 }),
  .Y({ S6032 })
);
NAND #() 
NAND_3617_ (
  .A({ S5991 }),
  .B({ S6030 }),
  .Y({ S6033 })
);
NAND #() 
NAND_3618_ (
  .A({ S6029 }),
  .B({ S6033 }),
  .Y({ S6034 })
);
NOT #() 
NOT_488_ (
  .A({ S6034 }),
  .Y({ S6035 })
);
NOR #() 
NOR_2042_ (
  .A({ S6002 }),
  .B({ S6006 }),
  .Y({ S6036 })
);
NAND #() 
NAND_3619_ (
  .A({ S6003 }),
  .B({ S6007 }),
  .Y({ S6037 })
);
NOR #() 
NOR_2043_ (
  .A({ S1116 }),
  .B({ S1849 }),
  .Y({ S6038 })
);
NAND #() 
NAND_3620_ (
  .A({ datapath_addsubunit_in1_2 }),
  .B({ S1848 }),
  .Y({ S6039 })
);
NOR #() 
NOR_2044_ (
  .A({ S1013 }),
  .B({ S1516 }),
  .Y({ S6040 })
);
NAND #() 
NAND_3621_ (
  .A({ datapath_addsubunit_in1_4 }),
  .B({ S1515 }),
  .Y({ S6041 })
);
NOR #() 
NOR_2045_ (
  .A({ S6000 }),
  .B({ S6040 }),
  .Y({ S6042 })
);
NAND #() 
NAND_3622_ (
  .A({ S6001 }),
  .B({ S6041 }),
  .Y({ S6043 })
);
NOR #() 
NOR_2046_ (
  .A({ S1013 }),
  .B({ S1746 }),
  .Y({ S6044 })
);
NAND #() 
NAND_3623_ (
  .A({ datapath_addsubunit_in1_4 }),
  .B({ S1745 }),
  .Y({ S6045 })
);
NOR #() 
NOR_2047_ (
  .A({ S6001 }),
  .B({ S6041 }),
  .Y({ S6046 })
);
NAND #() 
NAND_3624_ (
  .A({ S6000 }),
  .B({ S6040 }),
  .Y({ S6047 })
);
NOR #() 
NOR_2048_ (
  .A({ S6042 }),
  .B({ S6046 }),
  .Y({ S6048 })
);
NAND #() 
NAND_3625_ (
  .A({ S6043 }),
  .B({ S6047 }),
  .Y({ S6049 })
);
NOR #() 
NOR_2049_ (
  .A({ S6039 }),
  .B({ S6049 }),
  .Y({ S6050 })
);
NAND #() 
NAND_3626_ (
  .A({ S6038 }),
  .B({ S6048 }),
  .Y({ S6051 })
);
NOR #() 
NOR_2050_ (
  .A({ S6038 }),
  .B({ S6048 }),
  .Y({ S6052 })
);
NAND #() 
NAND_3627_ (
  .A({ S6039 }),
  .B({ S6049 }),
  .Y({ S6053 })
);
NOR #() 
NOR_2051_ (
  .A({ S6050 }),
  .B({ S6052 }),
  .Y({ S6054 })
);
NAND #() 
NAND_3628_ (
  .A({ S6051 }),
  .B({ S6053 }),
  .Y({ S6055 })
);
NOR #() 
NOR_2052_ (
  .A({ S6036 }),
  .B({ S6055 }),
  .Y({ S6056 })
);
NAND #() 
NAND_3629_ (
  .A({ S6037 }),
  .B({ S6054 }),
  .Y({ S6057 })
);
NAND #() 
NAND_3630_ (
  .A({ S6036 }),
  .B({ S6055 }),
  .Y({ S6058 })
);
NAND #() 
NAND_3631_ (
  .A({ S6057 }),
  .B({ S6058 }),
  .Y({ S6059 })
);
NOT #() 
NOT_489_ (
  .A({ S6059 }),
  .Y({ S6060 })
);
NAND #() 
NAND_3632_ (
  .A({ S6035 }),
  .B({ S6060 }),
  .Y({ S6061 })
);
NOT #() 
NOT_490_ (
  .A({ S6061 }),
  .Y({ S6062 })
);
NAND #() 
NAND_3633_ (
  .A({ S6034 }),
  .B({ S6059 }),
  .Y({ S6063 })
);
NAND #() 
NAND_3634_ (
  .A({ S6061 }),
  .B({ S6063 }),
  .Y({ S6064 })
);
NAND #() 
NAND_3635_ (
  .A({ S6026 }),
  .B({ S6064 }),
  .Y({ S6065 })
);
NOR #() 
NOR_2053_ (
  .A({ S6026 }),
  .B({ S6064 }),
  .Y({ S6066 })
);
NOT #() 
NOT_491_ (
  .A({ S6066 }),
  .Y({ S6067 })
);
NAND #() 
NAND_3636_ (
  .A({ S6065 }),
  .B({ S6067 }),
  .Y({ S6068 })
);
NAND #() 
NAND_3637_ (
  .A({ S6020 }),
  .B({ S6068 }),
  .Y({ S6069 })
);
NOR #() 
NOR_2054_ (
  .A({ S6020 }),
  .B({ S6068 }),
  .Y({ S6070 })
);
NOR #() 
NOR_2055_ (
  .A({ S5949 }),
  .B({ S6070 }),
  .Y({ S6071 })
);
NAND #() 
NAND_3638_ (
  .A({ S6069 }),
  .B({ S6071 }),
  .Y({ S6072 })
);
NAND #() 
NAND_3639_ (
  .A({ datapath_multdivunit_outmdu1_4 }),
  .B({ S5950 }),
  .Y({ S6073 })
);
NOT #() 
NOT_492_ (
  .A({ S6073 }),
  .Y({ S6074 })
);
NOR #() 
NOR_2056_ (
  .A({ S6025 }),
  .B({ S6074 }),
  .Y({ S6075 })
);
NAND #() 
NAND_3640_ (
  .A({ S6072 }),
  .B({ S6075 }),
  .Y({ S286 })
);
NOR #() 
NOR_2057_ (
  .A({ S3899 }),
  .B({ S4896 }),
  .Y({ S6076 })
);
NAND #() 
NAND_3641_ (
  .A({ datapath_multdivunit_outmdu1_5 }),
  .B({ S5950 }),
  .Y({ S6077 })
);
NOR #() 
NOR_2058_ (
  .A({ S6056 }),
  .B({ S6062 }),
  .Y({ S6078 })
);
NAND #() 
NAND_3642_ (
  .A({ S6057 }),
  .B({ S6061 }),
  .Y({ S6079 })
);
NOR #() 
NOR_2059_ (
  .A({ S1220 }),
  .B({ S2107 }),
  .Y({ S6080 })
);
NAND #() 
NAND_3643_ (
  .A({ datapath_addsubunit_in1_0 }),
  .B({ S2106 }),
  .Y({ S6081 })
);
NOR #() 
NOR_2060_ (
  .A({ S1116 }),
  .B({ S1953 }),
  .Y({ S6082 })
);
NAND #() 
NAND_3644_ (
  .A({ datapath_addsubunit_in1_2 }),
  .B({ S1952 }),
  .Y({ S6083 })
);
NOR #() 
NOR_2061_ (
  .A({ S6030 }),
  .B({ S6082 }),
  .Y({ S6084 })
);
NAND #() 
NAND_3645_ (
  .A({ S6031 }),
  .B({ S6083 }),
  .Y({ S6085 })
);
NOR #() 
NOR_2062_ (
  .A({ S1116 }),
  .B({ S1598 }),
  .Y({ S6086 })
);
NAND #() 
NAND_3646_ (
  .A({ datapath_addsubunit_in1_2 }),
  .B({ S1597 }),
  .Y({ S6087 })
);
NOR #() 
NOR_2063_ (
  .A({ S6031 }),
  .B({ S6083 }),
  .Y({ S6088 })
);
NAND #() 
NAND_3647_ (
  .A({ S6030 }),
  .B({ S6082 }),
  .Y({ S6089 })
);
NOR #() 
NOR_2064_ (
  .A({ S6084 }),
  .B({ S6088 }),
  .Y({ S6090 })
);
NAND #() 
NAND_3648_ (
  .A({ S6085 }),
  .B({ S6089 }),
  .Y({ S6091 })
);
NOR #() 
NOR_2065_ (
  .A({ S6081 }),
  .B({ S6091 }),
  .Y({ S6092 })
);
NAND #() 
NAND_3649_ (
  .A({ S6080 }),
  .B({ S6090 }),
  .Y({ S6093 })
);
NOR #() 
NOR_2066_ (
  .A({ S6080 }),
  .B({ S6090 }),
  .Y({ S6094 })
);
NAND #() 
NAND_3650_ (
  .A({ S6081 }),
  .B({ S6091 }),
  .Y({ S6095 })
);
NOR #() 
NOR_2067_ (
  .A({ S6092 }),
  .B({ S6094 }),
  .Y({ S6096 })
);
NAND #() 
NAND_3651_ (
  .A({ S6093 }),
  .B({ S6095 }),
  .Y({ S6097 })
);
NOR #() 
NOR_2068_ (
  .A({ S6046 }),
  .B({ S6050 }),
  .Y({ S6098 })
);
NAND #() 
NAND_3652_ (
  .A({ S6047 }),
  .B({ S6051 }),
  .Y({ S6099 })
);
NOR #() 
NOR_2069_ (
  .A({ S1065 }),
  .B({ S1849 }),
  .Y({ S6100 })
);
NAND #() 
NAND_3653_ (
  .A({ datapath_addsubunit_in1_3 }),
  .B({ S1848 }),
  .Y({ S6101 })
);
NOR #() 
NOR_2070_ (
  .A({ S963 }),
  .B({ S1516 }),
  .Y({ S6102 })
);
NAND #() 
NAND_3654_ (
  .A({ datapath_addsubunit_in1_5 }),
  .B({ S1515 }),
  .Y({ S6103 })
);
NOR #() 
NOR_2071_ (
  .A({ S6044 }),
  .B({ S6102 }),
  .Y({ S6104 })
);
NAND #() 
NAND_3655_ (
  .A({ S6045 }),
  .B({ S6103 }),
  .Y({ S6105 })
);
NOR #() 
NOR_2072_ (
  .A({ S963 }),
  .B({ S1746 }),
  .Y({ S6106 })
);
NAND #() 
NAND_3656_ (
  .A({ datapath_addsubunit_in1_5 }),
  .B({ S1745 }),
  .Y({ S6107 })
);
NOR #() 
NOR_2073_ (
  .A({ S6045 }),
  .B({ S6103 }),
  .Y({ S6108 })
);
NAND #() 
NAND_3657_ (
  .A({ S6044 }),
  .B({ S6102 }),
  .Y({ S6109 })
);
NOR #() 
NOR_2074_ (
  .A({ S6104 }),
  .B({ S6108 }),
  .Y({ S6110 })
);
NAND #() 
NAND_3658_ (
  .A({ S6105 }),
  .B({ S6109 }),
  .Y({ S6111 })
);
NOR #() 
NOR_2075_ (
  .A({ S6101 }),
  .B({ S6111 }),
  .Y({ S6112 })
);
NAND #() 
NAND_3659_ (
  .A({ S6100 }),
  .B({ S6110 }),
  .Y({ S6113 })
);
NOR #() 
NOR_2076_ (
  .A({ S6100 }),
  .B({ S6110 }),
  .Y({ S6114 })
);
NAND #() 
NAND_3660_ (
  .A({ S6101 }),
  .B({ S6111 }),
  .Y({ S6115 })
);
NOR #() 
NOR_2077_ (
  .A({ S6112 }),
  .B({ S6114 }),
  .Y({ S6116 })
);
NAND #() 
NAND_3661_ (
  .A({ S6113 }),
  .B({ S6115 }),
  .Y({ S6117 })
);
NOR #() 
NOR_2078_ (
  .A({ S6098 }),
  .B({ S6117 }),
  .Y({ S6118 })
);
NAND #() 
NAND_3662_ (
  .A({ S6099 }),
  .B({ S6116 }),
  .Y({ S6119 })
);
NOR #() 
NOR_2079_ (
  .A({ S6099 }),
  .B({ S6116 }),
  .Y({ S6120 })
);
NAND #() 
NAND_3663_ (
  .A({ S6098 }),
  .B({ S6117 }),
  .Y({ S6121 })
);
NOR #() 
NOR_2080_ (
  .A({ S6118 }),
  .B({ S6120 }),
  .Y({ S6122 })
);
NAND #() 
NAND_3664_ (
  .A({ S6119 }),
  .B({ S6121 }),
  .Y({ S6123 })
);
NOR #() 
NOR_2081_ (
  .A({ S6097 }),
  .B({ S6123 }),
  .Y({ S6124 })
);
NAND #() 
NAND_3665_ (
  .A({ S6096 }),
  .B({ S6122 }),
  .Y({ S6125 })
);
NOR #() 
NOR_2082_ (
  .A({ S6096 }),
  .B({ S6122 }),
  .Y({ S6126 })
);
NAND #() 
NAND_3666_ (
  .A({ S6097 }),
  .B({ S6123 }),
  .Y({ S6127 })
);
NOR #() 
NOR_2083_ (
  .A({ S6124 }),
  .B({ S6126 }),
  .Y({ S6128 })
);
NAND #() 
NAND_3667_ (
  .A({ S6125 }),
  .B({ S6127 }),
  .Y({ S6129 })
);
NOR #() 
NOR_2084_ (
  .A({ S6078 }),
  .B({ S6129 }),
  .Y({ S6130 })
);
NOR #() 
NOR_2085_ (
  .A({ S6079 }),
  .B({ S6128 }),
  .Y({ S6131 })
);
NOR #() 
NOR_2086_ (
  .A({ S6130 }),
  .B({ S6131 }),
  .Y({ S6132 })
);
NOT #() 
NOT_493_ (
  .A({ S6132 }),
  .Y({ S6133 })
);
NOR #() 
NOR_2087_ (
  .A({ S6033 }),
  .B({ S6133 }),
  .Y({ S6134 })
);
NOR #() 
NOR_2088_ (
  .A({ S6032 }),
  .B({ S6132 }),
  .Y({ S6135 })
);
NOR #() 
NOR_2089_ (
  .A({ S6134 }),
  .B({ S6135 }),
  .Y({ S6136 })
);
NAND #() 
NAND_3668_ (
  .A({ S6066 }),
  .B({ S6136 }),
  .Y({ S6137 })
);
NOT #() 
NOT_494_ (
  .A({ S6137 }),
  .Y({ S6138 })
);
NOR #() 
NOR_2090_ (
  .A({ S6066 }),
  .B({ S6136 }),
  .Y({ S6139 })
);
NOR #() 
NOR_2091_ (
  .A({ S6138 }),
  .B({ S6139 }),
  .Y({ S6140 })
);
NAND #() 
NAND_3669_ (
  .A({ S6070 }),
  .B({ S6140 }),
  .Y({ S6141 })
);
NOR #() 
NOR_2092_ (
  .A({ S6070 }),
  .B({ S6140 }),
  .Y({ S6142 })
);
NAND #() 
NAND_3670_ (
  .A({ S5948 }),
  .B({ S6141 }),
  .Y({ S6143 })
);
NOR #() 
NOR_2093_ (
  .A({ S6142 }),
  .B({ S6143 }),
  .Y({ S6144 })
);
NOR #() 
NOR_2094_ (
  .A({ S6076 }),
  .B({ S6144 }),
  .Y({ S6145 })
);
NAND #() 
NAND_3671_ (
  .A({ S6077 }),
  .B({ S6145 }),
  .Y({ S287 })
);
NOR #() 
NOR_2095_ (
  .A({ S3899 }),
  .B({ S4709 }),
  .Y({ S6146 })
);
NAND #() 
NAND_3672_ (
  .A({ datapath_multdivunit_outmdu1_6 }),
  .B({ S5950 }),
  .Y({ S6147 })
);
NOR #() 
NOR_2096_ (
  .A({ S6130 }),
  .B({ S6134 }),
  .Y({ S6148 })
);
NOT #() 
NOT_495_ (
  .A({ S6148 }),
  .Y({ S6149 })
);
NOR #() 
NOR_2097_ (
  .A({ S1220 }),
  .B({ S2206 }),
  .Y({ S6150 })
);
NAND #() 
NAND_3673_ (
  .A({ datapath_addsubunit_in1_0 }),
  .B({ S2205 }),
  .Y({ S6151 })
);
NOR #() 
NOR_2098_ (
  .A({ S6088 }),
  .B({ S6092 }),
  .Y({ S6152 })
);
NAND #() 
NAND_3674_ (
  .A({ S6089 }),
  .B({ S6093 }),
  .Y({ S6153 })
);
NOR #() 
NOR_2099_ (
  .A({ S6151 }),
  .B({ S6152 }),
  .Y({ S6154 })
);
NAND #() 
NAND_3675_ (
  .A({ S6150 }),
  .B({ S6153 }),
  .Y({ S6155 })
);
NAND #() 
NAND_3676_ (
  .A({ S6151 }),
  .B({ S6152 }),
  .Y({ S6156 })
);
NAND #() 
NAND_3677_ (
  .A({ S6155 }),
  .B({ S6156 }),
  .Y({ S6157 })
);
NOT #() 
NOT_496_ (
  .A({ S6157 }),
  .Y({ S6158 })
);
NOR #() 
NOR_2100_ (
  .A({ S6118 }),
  .B({ S6124 }),
  .Y({ S6159 })
);
NAND #() 
NAND_3678_ (
  .A({ S6119 }),
  .B({ S6125 }),
  .Y({ S6160 })
);
NOR #() 
NOR_2101_ (
  .A({ S1168 }),
  .B({ S2107 }),
  .Y({ S6161 })
);
NAND #() 
NAND_3679_ (
  .A({ datapath_addsubunit_in1_1 }),
  .B({ S2106 }),
  .Y({ S6162 })
);
NOR #() 
NOR_2102_ (
  .A({ S1065 }),
  .B({ S1953 }),
  .Y({ S6163 })
);
NAND #() 
NAND_3680_ (
  .A({ datapath_addsubunit_in1_3 }),
  .B({ S1952 }),
  .Y({ S6164 })
);
NOR #() 
NOR_2103_ (
  .A({ S6086 }),
  .B({ S6163 }),
  .Y({ S6165 })
);
NAND #() 
NAND_3681_ (
  .A({ S6087 }),
  .B({ S6164 }),
  .Y({ S6166 })
);
NOR #() 
NOR_2104_ (
  .A({ S1065 }),
  .B({ S1598 }),
  .Y({ S6167 })
);
NAND #() 
NAND_3682_ (
  .A({ datapath_addsubunit_in1_3 }),
  .B({ S1597 }),
  .Y({ S6168 })
);
NOR #() 
NOR_2105_ (
  .A({ S6087 }),
  .B({ S6164 }),
  .Y({ S6169 })
);
NAND #() 
NAND_3683_ (
  .A({ S6086 }),
  .B({ S6163 }),
  .Y({ S6170 })
);
NOR #() 
NOR_2106_ (
  .A({ S6165 }),
  .B({ S6169 }),
  .Y({ S6171 })
);
NAND #() 
NAND_3684_ (
  .A({ S6166 }),
  .B({ S6170 }),
  .Y({ S6172 })
);
NOR #() 
NOR_2107_ (
  .A({ S6162 }),
  .B({ S6172 }),
  .Y({ S6173 })
);
NAND #() 
NAND_3685_ (
  .A({ S6161 }),
  .B({ S6171 }),
  .Y({ S6174 })
);
NOR #() 
NOR_2108_ (
  .A({ S6161 }),
  .B({ S6171 }),
  .Y({ S6175 })
);
NAND #() 
NAND_3686_ (
  .A({ S6162 }),
  .B({ S6172 }),
  .Y({ S6176 })
);
NOR #() 
NOR_2109_ (
  .A({ S6173 }),
  .B({ S6175 }),
  .Y({ S6177 })
);
NAND #() 
NAND_3687_ (
  .A({ S6174 }),
  .B({ S6176 }),
  .Y({ S6178 })
);
NOR #() 
NOR_2110_ (
  .A({ S6108 }),
  .B({ S6112 }),
  .Y({ S6179 })
);
NAND #() 
NAND_3688_ (
  .A({ S6109 }),
  .B({ S6113 }),
  .Y({ S6180 })
);
NOR #() 
NOR_2111_ (
  .A({ S1013 }),
  .B({ S1849 }),
  .Y({ S6181 })
);
NAND #() 
NAND_3689_ (
  .A({ datapath_addsubunit_in1_4 }),
  .B({ S1848 }),
  .Y({ S6182 })
);
NOR #() 
NOR_2112_ (
  .A({ S910 }),
  .B({ S1516 }),
  .Y({ S6183 })
);
NAND #() 
NAND_3690_ (
  .A({ datapath_addsubunit_in1_6 }),
  .B({ S1515 }),
  .Y({ S6184 })
);
NOR #() 
NOR_2113_ (
  .A({ S6106 }),
  .B({ S6183 }),
  .Y({ S6185 })
);
NAND #() 
NAND_3691_ (
  .A({ S6107 }),
  .B({ S6184 }),
  .Y({ S6186 })
);
NOR #() 
NOR_2114_ (
  .A({ S910 }),
  .B({ S1746 }),
  .Y({ S6187 })
);
NAND #() 
NAND_3692_ (
  .A({ datapath_addsubunit_in1_6 }),
  .B({ S1745 }),
  .Y({ S6188 })
);
NOR #() 
NOR_2115_ (
  .A({ S6107 }),
  .B({ S6184 }),
  .Y({ S6189 })
);
NAND #() 
NAND_3693_ (
  .A({ S6106 }),
  .B({ S6183 }),
  .Y({ S6190 })
);
NOR #() 
NOR_2116_ (
  .A({ S6185 }),
  .B({ S6189 }),
  .Y({ S6191 })
);
NAND #() 
NAND_3694_ (
  .A({ S6186 }),
  .B({ S6190 }),
  .Y({ S6192 })
);
NOR #() 
NOR_2117_ (
  .A({ S6182 }),
  .B({ S6192 }),
  .Y({ S6193 })
);
NAND #() 
NAND_3695_ (
  .A({ S6181 }),
  .B({ S6191 }),
  .Y({ S6194 })
);
NOR #() 
NOR_2118_ (
  .A({ S6181 }),
  .B({ S6191 }),
  .Y({ S6195 })
);
NAND #() 
NAND_3696_ (
  .A({ S6182 }),
  .B({ S6192 }),
  .Y({ S6196 })
);
NOR #() 
NOR_2119_ (
  .A({ S6193 }),
  .B({ S6195 }),
  .Y({ S6197 })
);
NAND #() 
NAND_3697_ (
  .A({ S6194 }),
  .B({ S6196 }),
  .Y({ S6198 })
);
NOR #() 
NOR_2120_ (
  .A({ S6179 }),
  .B({ S6198 }),
  .Y({ S6199 })
);
NAND #() 
NAND_3698_ (
  .A({ S6180 }),
  .B({ S6197 }),
  .Y({ S6200 })
);
NOR #() 
NOR_2121_ (
  .A({ S6180 }),
  .B({ S6197 }),
  .Y({ S6201 })
);
NAND #() 
NAND_3699_ (
  .A({ S6179 }),
  .B({ S6198 }),
  .Y({ S6202 })
);
NOR #() 
NOR_2122_ (
  .A({ S6199 }),
  .B({ S6201 }),
  .Y({ S6203 })
);
NAND #() 
NAND_3700_ (
  .A({ S6200 }),
  .B({ S6202 }),
  .Y({ S6204 })
);
NOR #() 
NOR_2123_ (
  .A({ S6178 }),
  .B({ S6204 }),
  .Y({ S6205 })
);
NAND #() 
NAND_3701_ (
  .A({ S6177 }),
  .B({ S6203 }),
  .Y({ S6206 })
);
NOR #() 
NOR_2124_ (
  .A({ S6177 }),
  .B({ S6203 }),
  .Y({ S6207 })
);
NAND #() 
NAND_3702_ (
  .A({ S6178 }),
  .B({ S6204 }),
  .Y({ S6208 })
);
NOR #() 
NOR_2125_ (
  .A({ S6205 }),
  .B({ S6207 }),
  .Y({ S6209 })
);
NAND #() 
NAND_3703_ (
  .A({ S6206 }),
  .B({ S6208 }),
  .Y({ S6210 })
);
NOR #() 
NOR_2126_ (
  .A({ S6159 }),
  .B({ S6210 }),
  .Y({ S6211 })
);
NAND #() 
NAND_3704_ (
  .A({ S6160 }),
  .B({ S6209 }),
  .Y({ S6212 })
);
NAND #() 
NAND_3705_ (
  .A({ S6159 }),
  .B({ S6210 }),
  .Y({ S6213 })
);
NAND #() 
NAND_3706_ (
  .A({ S6212 }),
  .B({ S6213 }),
  .Y({ S6214 })
);
NOT #() 
NOT_497_ (
  .A({ S6214 }),
  .Y({ S6215 })
);
NAND #() 
NAND_3707_ (
  .A({ S6158 }),
  .B({ S6215 }),
  .Y({ S6216 })
);
NOT #() 
NOT_498_ (
  .A({ S6216 }),
  .Y({ S6217 })
);
NAND #() 
NAND_3708_ (
  .A({ S6157 }),
  .B({ S6214 }),
  .Y({ S6218 })
);
NAND #() 
NAND_3709_ (
  .A({ S6216 }),
  .B({ S6218 }),
  .Y({ S6219 })
);
NOT #() 
NOT_499_ (
  .A({ S6219 }),
  .Y({ S6220 })
);
NAND #() 
NAND_3710_ (
  .A({ S6148 }),
  .B({ S6219 }),
  .Y({ S6221 })
);
NAND #() 
NAND_3711_ (
  .A({ S6149 }),
  .B({ S6220 }),
  .Y({ S6222 })
);
NOT #() 
NOT_500_ (
  .A({ S6222 }),
  .Y({ S6223 })
);
NAND #() 
NAND_3712_ (
  .A({ S6221 }),
  .B({ S6222 }),
  .Y({ S6224 })
);
NOR #() 
NOR_2127_ (
  .A({ S6137 }),
  .B({ S6224 }),
  .Y({ S6225 })
);
NOT #() 
NOT_501_ (
  .A({ S6225 }),
  .Y({ S6226 })
);
NAND #() 
NAND_3713_ (
  .A({ S6137 }),
  .B({ S6224 }),
  .Y({ S6227 })
);
NAND #() 
NAND_3714_ (
  .A({ S6226 }),
  .B({ S6227 }),
  .Y({ S6228 })
);
NOR #() 
NOR_2128_ (
  .A({ S6141 }),
  .B({ S6228 }),
  .Y({ S6229 })
);
NAND #() 
NAND_3715_ (
  .A({ S6141 }),
  .B({ S6228 }),
  .Y({ S6230 })
);
NAND #() 
NAND_3716_ (
  .A({ S5948 }),
  .B({ S6230 }),
  .Y({ S6231 })
);
NOR #() 
NOR_2129_ (
  .A({ S6229 }),
  .B({ S6231 }),
  .Y({ S6232 })
);
NOR #() 
NOR_2130_ (
  .A({ S6146 }),
  .B({ S6232 }),
  .Y({ S6233 })
);
NAND #() 
NAND_3717_ (
  .A({ S6147 }),
  .B({ S6233 }),
  .Y({ S288 })
);
NOR #() 
NOR_2131_ (
  .A({ S3899 }),
  .B({ S4571 }),
  .Y({ S6234 })
);
NAND #() 
NAND_3718_ (
  .A({ datapath_multdivunit_outmdu1_7 }),
  .B({ S5950 }),
  .Y({ S6235 })
);
NOR #() 
NOR_2132_ (
  .A({ S6211 }),
  .B({ S6217 }),
  .Y({ S6236 })
);
NAND #() 
NAND_3719_ (
  .A({ S6212 }),
  .B({ S6216 }),
  .Y({ S6237 })
);
NOR #() 
NOR_2133_ (
  .A({ S1220 }),
  .B({ S2312 }),
  .Y({ S6238 })
);
NAND #() 
NAND_3720_ (
  .A({ datapath_addsubunit_in1_0 }),
  .B({ S2311 }),
  .Y({ S6239 })
);
NOR #() 
NOR_2134_ (
  .A({ S1168 }),
  .B({ S2206 }),
  .Y({ S6240 })
);
NAND #() 
NAND_3721_ (
  .A({ datapath_addsubunit_in1_1 }),
  .B({ S2205 }),
  .Y({ S6241 })
);
NOR #() 
NOR_2135_ (
  .A({ S6238 }),
  .B({ S6240 }),
  .Y({ S6242 })
);
NAND #() 
NAND_3722_ (
  .A({ S6239 }),
  .B({ S6241 }),
  .Y({ S6243 })
);
NOR #() 
NOR_2136_ (
  .A({ S1168 }),
  .B({ S2312 }),
  .Y({ S6244 })
);
NAND #() 
NAND_3723_ (
  .A({ datapath_addsubunit_in1_1 }),
  .B({ S2311 }),
  .Y({ S6245 })
);
NOR #() 
NOR_2137_ (
  .A({ S6151 }),
  .B({ S6245 }),
  .Y({ S6246 })
);
NAND #() 
NAND_3724_ (
  .A({ S6150 }),
  .B({ S6244 }),
  .Y({ S6247 })
);
NOR #() 
NOR_2138_ (
  .A({ S6242 }),
  .B({ S6246 }),
  .Y({ S6248 })
);
NAND #() 
NAND_3725_ (
  .A({ S6243 }),
  .B({ S6247 }),
  .Y({ S6249 })
);
NOR #() 
NOR_2139_ (
  .A({ S6169 }),
  .B({ S6173 }),
  .Y({ S6250 })
);
NAND #() 
NAND_3726_ (
  .A({ S6170 }),
  .B({ S6174 }),
  .Y({ S6251 })
);
NOR #() 
NOR_2140_ (
  .A({ S6248 }),
  .B({ S6251 }),
  .Y({ S6252 })
);
NAND #() 
NAND_3727_ (
  .A({ S6249 }),
  .B({ S6250 }),
  .Y({ S6253 })
);
NOR #() 
NOR_2141_ (
  .A({ S6249 }),
  .B({ S6250 }),
  .Y({ S6254 })
);
NAND #() 
NAND_3728_ (
  .A({ S6248 }),
  .B({ S6251 }),
  .Y({ S6255 })
);
NOR #() 
NOR_2142_ (
  .A({ S6252 }),
  .B({ S6254 }),
  .Y({ S6256 })
);
NAND #() 
NAND_3729_ (
  .A({ S6253 }),
  .B({ S6255 }),
  .Y({ S6257 })
);
NOR #() 
NOR_2143_ (
  .A({ S6199 }),
  .B({ S6205 }),
  .Y({ S6258 })
);
NAND #() 
NAND_3730_ (
  .A({ S6200 }),
  .B({ S6206 }),
  .Y({ S6259 })
);
NOR #() 
NOR_2144_ (
  .A({ S1116 }),
  .B({ S2107 }),
  .Y({ S6260 })
);
NAND #() 
NAND_3731_ (
  .A({ datapath_addsubunit_in1_2 }),
  .B({ S2106 }),
  .Y({ S6261 })
);
NOR #() 
NOR_2145_ (
  .A({ S1013 }),
  .B({ S1953 }),
  .Y({ S6262 })
);
NAND #() 
NAND_3732_ (
  .A({ datapath_addsubunit_in1_4 }),
  .B({ S1952 }),
  .Y({ S6263 })
);
NOR #() 
NOR_2146_ (
  .A({ S6167 }),
  .B({ S6262 }),
  .Y({ S6264 })
);
NAND #() 
NAND_3733_ (
  .A({ S6168 }),
  .B({ S6263 }),
  .Y({ S6265 })
);
NOR #() 
NOR_2147_ (
  .A({ S1013 }),
  .B({ S1598 }),
  .Y({ S6266 })
);
NAND #() 
NAND_3734_ (
  .A({ datapath_addsubunit_in1_4 }),
  .B({ S1597 }),
  .Y({ S6267 })
);
NOR #() 
NOR_2148_ (
  .A({ S6168 }),
  .B({ S6263 }),
  .Y({ S6268 })
);
NAND #() 
NAND_3735_ (
  .A({ S6167 }),
  .B({ S6262 }),
  .Y({ S6269 })
);
NOR #() 
NOR_2149_ (
  .A({ S6264 }),
  .B({ S6268 }),
  .Y({ S6270 })
);
NAND #() 
NAND_3736_ (
  .A({ S6265 }),
  .B({ S6269 }),
  .Y({ S6271 })
);
NOR #() 
NOR_2150_ (
  .A({ S6261 }),
  .B({ S6271 }),
  .Y({ S6272 })
);
NAND #() 
NAND_3737_ (
  .A({ S6260 }),
  .B({ S6270 }),
  .Y({ S6273 })
);
NOR #() 
NOR_2151_ (
  .A({ S6260 }),
  .B({ S6270 }),
  .Y({ S6274 })
);
NAND #() 
NAND_3738_ (
  .A({ S6261 }),
  .B({ S6271 }),
  .Y({ S6275 })
);
NOR #() 
NOR_2152_ (
  .A({ S6272 }),
  .B({ S6274 }),
  .Y({ S6276 })
);
NAND #() 
NAND_3739_ (
  .A({ S6273 }),
  .B({ S6275 }),
  .Y({ S6277 })
);
NOR #() 
NOR_2153_ (
  .A({ S6189 }),
  .B({ S6193 }),
  .Y({ S6278 })
);
NAND #() 
NAND_3740_ (
  .A({ S6190 }),
  .B({ S6194 }),
  .Y({ S6279 })
);
NOR #() 
NOR_2154_ (
  .A({ S963 }),
  .B({ S1849 }),
  .Y({ S6280 })
);
NAND #() 
NAND_3741_ (
  .A({ datapath_addsubunit_in1_5 }),
  .B({ S1848 }),
  .Y({ S6281 })
);
NOR #() 
NOR_2155_ (
  .A({ S858 }),
  .B({ S1516 }),
  .Y({ S6282 })
);
NAND #() 
NAND_3742_ (
  .A({ datapath_addsubunit_in1_7 }),
  .B({ S1515 }),
  .Y({ S6283 })
);
NOR #() 
NOR_2156_ (
  .A({ S6187 }),
  .B({ S6282 }),
  .Y({ S6284 })
);
NAND #() 
NAND_3743_ (
  .A({ S6188 }),
  .B({ S6283 }),
  .Y({ S6285 })
);
NOR #() 
NOR_2157_ (
  .A({ S858 }),
  .B({ S1746 }),
  .Y({ S6286 })
);
NAND #() 
NAND_3744_ (
  .A({ datapath_addsubunit_in1_7 }),
  .B({ S1745 }),
  .Y({ S6287 })
);
NOR #() 
NOR_2158_ (
  .A({ S6188 }),
  .B({ S6283 }),
  .Y({ S6288 })
);
NAND #() 
NAND_3745_ (
  .A({ S6187 }),
  .B({ S6282 }),
  .Y({ S6289 })
);
NOR #() 
NOR_2159_ (
  .A({ S6284 }),
  .B({ S6288 }),
  .Y({ S6290 })
);
NAND #() 
NAND_3746_ (
  .A({ S6285 }),
  .B({ S6289 }),
  .Y({ S6291 })
);
NOR #() 
NOR_2160_ (
  .A({ S6281 }),
  .B({ S6291 }),
  .Y({ S6292 })
);
NAND #() 
NAND_3747_ (
  .A({ S6280 }),
  .B({ S6290 }),
  .Y({ S6293 })
);
NOR #() 
NOR_2161_ (
  .A({ S6280 }),
  .B({ S6290 }),
  .Y({ S6294 })
);
NAND #() 
NAND_3748_ (
  .A({ S6281 }),
  .B({ S6291 }),
  .Y({ S6295 })
);
NOR #() 
NOR_2162_ (
  .A({ S6292 }),
  .B({ S6294 }),
  .Y({ S6296 })
);
NAND #() 
NAND_3749_ (
  .A({ S6293 }),
  .B({ S6295 }),
  .Y({ S6297 })
);
NOR #() 
NOR_2163_ (
  .A({ S6278 }),
  .B({ S6297 }),
  .Y({ S6298 })
);
NAND #() 
NAND_3750_ (
  .A({ S6279 }),
  .B({ S6296 }),
  .Y({ S6299 })
);
NOR #() 
NOR_2164_ (
  .A({ S6279 }),
  .B({ S6296 }),
  .Y({ S6300 })
);
NAND #() 
NAND_3751_ (
  .A({ S6278 }),
  .B({ S6297 }),
  .Y({ S6301 })
);
NOR #() 
NOR_2165_ (
  .A({ S6298 }),
  .B({ S6300 }),
  .Y({ S6302 })
);
NAND #() 
NAND_3752_ (
  .A({ S6299 }),
  .B({ S6301 }),
  .Y({ S6303 })
);
NOR #() 
NOR_2166_ (
  .A({ S6277 }),
  .B({ S6303 }),
  .Y({ S6304 })
);
NAND #() 
NAND_3753_ (
  .A({ S6276 }),
  .B({ S6302 }),
  .Y({ S6305 })
);
NOR #() 
NOR_2167_ (
  .A({ S6276 }),
  .B({ S6302 }),
  .Y({ S6306 })
);
NAND #() 
NAND_3754_ (
  .A({ S6277 }),
  .B({ S6303 }),
  .Y({ S6307 })
);
NOR #() 
NOR_2168_ (
  .A({ S6304 }),
  .B({ S6306 }),
  .Y({ S6308 })
);
NAND #() 
NAND_3755_ (
  .A({ S6305 }),
  .B({ S6307 }),
  .Y({ S6309 })
);
NOR #() 
NOR_2169_ (
  .A({ S6258 }),
  .B({ S6309 }),
  .Y({ S6310 })
);
NAND #() 
NAND_3756_ (
  .A({ S6259 }),
  .B({ S6308 }),
  .Y({ S6311 })
);
NOR #() 
NOR_2170_ (
  .A({ S6259 }),
  .B({ S6308 }),
  .Y({ S6312 })
);
NAND #() 
NAND_3757_ (
  .A({ S6258 }),
  .B({ S6309 }),
  .Y({ S6313 })
);
NOR #() 
NOR_2171_ (
  .A({ S6310 }),
  .B({ S6312 }),
  .Y({ S6314 })
);
NAND #() 
NAND_3758_ (
  .A({ S6311 }),
  .B({ S6313 }),
  .Y({ S6315 })
);
NOR #() 
NOR_2172_ (
  .A({ S6257 }),
  .B({ S6315 }),
  .Y({ S6316 })
);
NAND #() 
NAND_3759_ (
  .A({ S6256 }),
  .B({ S6314 }),
  .Y({ S6317 })
);
NOR #() 
NOR_2173_ (
  .A({ S6256 }),
  .B({ S6314 }),
  .Y({ S6318 })
);
NAND #() 
NAND_3760_ (
  .A({ S6257 }),
  .B({ S6315 }),
  .Y({ S6319 })
);
NOR #() 
NOR_2174_ (
  .A({ S6316 }),
  .B({ S6318 }),
  .Y({ S6320 })
);
NAND #() 
NAND_3761_ (
  .A({ S6317 }),
  .B({ S6319 }),
  .Y({ S6321 })
);
NOR #() 
NOR_2175_ (
  .A({ S6236 }),
  .B({ S6321 }),
  .Y({ S6322 })
);
NAND #() 
NAND_3762_ (
  .A({ S6237 }),
  .B({ S6320 }),
  .Y({ S6323 })
);
NAND #() 
NAND_3763_ (
  .A({ S6236 }),
  .B({ S6321 }),
  .Y({ S6324 })
);
NAND #() 
NAND_3764_ (
  .A({ S6323 }),
  .B({ S6324 }),
  .Y({ S6325 })
);
NOT #() 
NOT_502_ (
  .A({ S6325 }),
  .Y({ S6326 })
);
NAND #() 
NAND_3765_ (
  .A({ S6154 }),
  .B({ S6326 }),
  .Y({ S6327 })
);
NOT #() 
NOT_503_ (
  .A({ S6327 }),
  .Y({ S6328 })
);
NAND #() 
NAND_3766_ (
  .A({ S6155 }),
  .B({ S6325 }),
  .Y({ S6329 })
);
NAND #() 
NAND_3767_ (
  .A({ S6327 }),
  .B({ S6329 }),
  .Y({ S6330 })
);
NOT #() 
NOT_504_ (
  .A({ S6330 }),
  .Y({ S6331 })
);
NAND #() 
NAND_3768_ (
  .A({ S6223 }),
  .B({ S6331 }),
  .Y({ S6332 })
);
NOT #() 
NOT_505_ (
  .A({ S6332 }),
  .Y({ S6333 })
);
NAND #() 
NAND_3769_ (
  .A({ S6222 }),
  .B({ S6330 }),
  .Y({ S6334 })
);
NAND #() 
NAND_3770_ (
  .A({ S6332 }),
  .B({ S6334 }),
  .Y({ S6335 })
);
NOT #() 
NOT_506_ (
  .A({ S6335 }),
  .Y({ S6336 })
);
NAND #() 
NAND_3771_ (
  .A({ S6229 }),
  .B({ S6336 }),
  .Y({ S6337 })
);
NAND #() 
NAND_3772_ (
  .A({ S5948 }),
  .B({ S6337 }),
  .Y({ S6338 })
);
NOR #() 
NOR_2176_ (
  .A({ S6225 }),
  .B({ S6229 }),
  .Y({ S6339 })
);
NAND #() 
NAND_3773_ (
  .A({ S6335 }),
  .B({ S6339 }),
  .Y({ S6340 })
);
NAND #() 
NAND_3774_ (
  .A({ S6225 }),
  .B({ S6336 }),
  .Y({ S6341 })
);
NAND #() 
NAND_3775_ (
  .A({ S6340 }),
  .B({ S6341 }),
  .Y({ S6342 })
);
NOR #() 
NOR_2177_ (
  .A({ S6338 }),
  .B({ S6342 }),
  .Y({ S6343 })
);
NOR #() 
NOR_2178_ (
  .A({ S6234 }),
  .B({ S6343 }),
  .Y({ S6344 })
);
NAND #() 
NAND_3776_ (
  .A({ S6235 }),
  .B({ S6344 }),
  .Y({ S289 })
);
NOR #() 
NOR_2179_ (
  .A({ S3899 }),
  .B({ S4430 }),
  .Y({ S6345 })
);
NAND #() 
NAND_3777_ (
  .A({ datapath_multdivunit_outmdu1_8 }),
  .B({ S5950 }),
  .Y({ S6346 })
);
NOR #() 
NOR_2180_ (
  .A({ S6322 }),
  .B({ S6328 }),
  .Y({ S6347 })
);
NAND #() 
NAND_3778_ (
  .A({ S6323 }),
  .B({ S6327 }),
  .Y({ S6348 })
);
NOR #() 
NOR_2181_ (
  .A({ S6310 }),
  .B({ S6316 }),
  .Y({ S6349 })
);
NAND #() 
NAND_3779_ (
  .A({ S6311 }),
  .B({ S6317 }),
  .Y({ S6350 })
);
NOR #() 
NOR_2182_ (
  .A({ S1220 }),
  .B({ S2418 }),
  .Y({ S6351 })
);
NAND #() 
NAND_3780_ (
  .A({ datapath_addsubunit_in1_0 }),
  .B({ S2417 }),
  .Y({ S6352 })
);
NOR #() 
NOR_2183_ (
  .A({ S1116 }),
  .B({ S2206 }),
  .Y({ S6353 })
);
NAND #() 
NAND_3781_ (
  .A({ datapath_addsubunit_in1_2 }),
  .B({ S2205 }),
  .Y({ S6354 })
);
NOR #() 
NOR_2184_ (
  .A({ S6244 }),
  .B({ S6353 }),
  .Y({ S6355 })
);
NAND #() 
NAND_3782_ (
  .A({ S6245 }),
  .B({ S6354 }),
  .Y({ S6356 })
);
NOR #() 
NOR_2185_ (
  .A({ S1116 }),
  .B({ S2312 }),
  .Y({ S6357 })
);
NAND #() 
NAND_3783_ (
  .A({ datapath_addsubunit_in1_2 }),
  .B({ S2311 }),
  .Y({ S6358 })
);
NOR #() 
NOR_2186_ (
  .A({ S6245 }),
  .B({ S6354 }),
  .Y({ S6359 })
);
NAND #() 
NAND_3784_ (
  .A({ S6244 }),
  .B({ S6353 }),
  .Y({ S6360 })
);
NOR #() 
NOR_2187_ (
  .A({ S6355 }),
  .B({ S6359 }),
  .Y({ S6361 })
);
NAND #() 
NAND_3785_ (
  .A({ S6356 }),
  .B({ S6360 }),
  .Y({ S6362 })
);
NOR #() 
NOR_2188_ (
  .A({ S6352 }),
  .B({ S6362 }),
  .Y({ S6363 })
);
NAND #() 
NAND_3786_ (
  .A({ S6351 }),
  .B({ S6361 }),
  .Y({ S6364 })
);
NOR #() 
NOR_2189_ (
  .A({ S6351 }),
  .B({ S6361 }),
  .Y({ S6365 })
);
NAND #() 
NAND_3787_ (
  .A({ S6352 }),
  .B({ S6362 }),
  .Y({ S6366 })
);
NOR #() 
NOR_2190_ (
  .A({ S6363 }),
  .B({ S6365 }),
  .Y({ S6367 })
);
NAND #() 
NAND_3788_ (
  .A({ S6364 }),
  .B({ S6366 }),
  .Y({ S6368 })
);
NOR #() 
NOR_2191_ (
  .A({ S6268 }),
  .B({ S6272 }),
  .Y({ S6369 })
);
NAND #() 
NAND_3789_ (
  .A({ S6269 }),
  .B({ S6273 }),
  .Y({ S6370 })
);
NOR #() 
NOR_2192_ (
  .A({ S6368 }),
  .B({ S6369 }),
  .Y({ S6371 })
);
NAND #() 
NAND_3790_ (
  .A({ S6367 }),
  .B({ S6370 }),
  .Y({ S6372 })
);
NOR #() 
NOR_2193_ (
  .A({ S6367 }),
  .B({ S6370 }),
  .Y({ S6373 })
);
NAND #() 
NAND_3791_ (
  .A({ S6368 }),
  .B({ S6369 }),
  .Y({ S6374 })
);
NOR #() 
NOR_2194_ (
  .A({ S6371 }),
  .B({ S6373 }),
  .Y({ S6375 })
);
NAND #() 
NAND_3792_ (
  .A({ S6372 }),
  .B({ S6374 }),
  .Y({ S6376 })
);
NOR #() 
NOR_2195_ (
  .A({ S6247 }),
  .B({ S6376 }),
  .Y({ S6377 })
);
NAND #() 
NAND_3793_ (
  .A({ S6246 }),
  .B({ S6375 }),
  .Y({ S6378 })
);
NOR #() 
NOR_2196_ (
  .A({ S6246 }),
  .B({ S6375 }),
  .Y({ S6379 })
);
NAND #() 
NAND_3794_ (
  .A({ S6247 }),
  .B({ S6376 }),
  .Y({ S6380 })
);
NOR #() 
NOR_2197_ (
  .A({ S6377 }),
  .B({ S6379 }),
  .Y({ S6381 })
);
NAND #() 
NAND_3795_ (
  .A({ S6378 }),
  .B({ S6380 }),
  .Y({ S6382 })
);
NOR #() 
NOR_2198_ (
  .A({ S6298 }),
  .B({ S6304 }),
  .Y({ S6383 })
);
NAND #() 
NAND_3796_ (
  .A({ S6299 }),
  .B({ S6305 }),
  .Y({ S6384 })
);
NOR #() 
NOR_2199_ (
  .A({ S1065 }),
  .B({ S2107 }),
  .Y({ S6385 })
);
NAND #() 
NAND_3797_ (
  .A({ datapath_addsubunit_in1_3 }),
  .B({ S2106 }),
  .Y({ S6386 })
);
NOR #() 
NOR_2200_ (
  .A({ S963 }),
  .B({ S1953 }),
  .Y({ S6387 })
);
NAND #() 
NAND_3798_ (
  .A({ datapath_addsubunit_in1_5 }),
  .B({ S1952 }),
  .Y({ S6388 })
);
NOR #() 
NOR_2201_ (
  .A({ S6266 }),
  .B({ S6387 }),
  .Y({ S6389 })
);
NAND #() 
NAND_3799_ (
  .A({ S6267 }),
  .B({ S6388 }),
  .Y({ S6390 })
);
NOR #() 
NOR_2202_ (
  .A({ S963 }),
  .B({ S1598 }),
  .Y({ S6391 })
);
NAND #() 
NAND_3800_ (
  .A({ datapath_addsubunit_in1_5 }),
  .B({ S1597 }),
  .Y({ S6392 })
);
NOR #() 
NOR_2203_ (
  .A({ S6267 }),
  .B({ S6388 }),
  .Y({ S6393 })
);
NAND #() 
NAND_3801_ (
  .A({ S6266 }),
  .B({ S6387 }),
  .Y({ S6394 })
);
NOR #() 
NOR_2204_ (
  .A({ S6389 }),
  .B({ S6393 }),
  .Y({ S6395 })
);
NAND #() 
NAND_3802_ (
  .A({ S6390 }),
  .B({ S6394 }),
  .Y({ S6396 })
);
NOR #() 
NOR_2205_ (
  .A({ S6386 }),
  .B({ S6396 }),
  .Y({ S6397 })
);
NAND #() 
NAND_3803_ (
  .A({ S6385 }),
  .B({ S6395 }),
  .Y({ S6398 })
);
NOR #() 
NOR_2206_ (
  .A({ S6385 }),
  .B({ S6395 }),
  .Y({ S6399 })
);
NAND #() 
NAND_3804_ (
  .A({ S6386 }),
  .B({ S6396 }),
  .Y({ S6400 })
);
NOR #() 
NOR_2207_ (
  .A({ S6397 }),
  .B({ S6399 }),
  .Y({ S6401 })
);
NAND #() 
NAND_3805_ (
  .A({ S6398 }),
  .B({ S6400 }),
  .Y({ S6402 })
);
NOR #() 
NOR_2208_ (
  .A({ S6288 }),
  .B({ S6292 }),
  .Y({ S6403 })
);
NAND #() 
NAND_3806_ (
  .A({ S6289 }),
  .B({ S6293 }),
  .Y({ S6404 })
);
NOR #() 
NOR_2209_ (
  .A({ S910 }),
  .B({ S1849 }),
  .Y({ S6405 })
);
NAND #() 
NAND_3807_ (
  .A({ datapath_addsubunit_in1_6 }),
  .B({ S1848 }),
  .Y({ S6406 })
);
NOR #() 
NOR_2210_ (
  .A({ S805 }),
  .B({ S1516 }),
  .Y({ S6407 })
);
NAND #() 
NAND_3808_ (
  .A({ datapath_addsubunit_in1_8 }),
  .B({ S1515 }),
  .Y({ S6408 })
);
NOR #() 
NOR_2211_ (
  .A({ S6286 }),
  .B({ S6407 }),
  .Y({ S6409 })
);
NAND #() 
NAND_3809_ (
  .A({ S6287 }),
  .B({ S6408 }),
  .Y({ S6410 })
);
NOR #() 
NOR_2212_ (
  .A({ S805 }),
  .B({ S1746 }),
  .Y({ S6411 })
);
NAND #() 
NAND_3810_ (
  .A({ datapath_addsubunit_in1_8 }),
  .B({ S1745 }),
  .Y({ S6412 })
);
NOR #() 
NOR_2213_ (
  .A({ S6287 }),
  .B({ S6408 }),
  .Y({ S6413 })
);
NAND #() 
NAND_3811_ (
  .A({ S6286 }),
  .B({ S6407 }),
  .Y({ S6414 })
);
NOR #() 
NOR_2214_ (
  .A({ S6409 }),
  .B({ S6413 }),
  .Y({ S6415 })
);
NAND #() 
NAND_3812_ (
  .A({ S6410 }),
  .B({ S6414 }),
  .Y({ S6416 })
);
NOR #() 
NOR_2215_ (
  .A({ S6406 }),
  .B({ S6416 }),
  .Y({ S6417 })
);
NAND #() 
NAND_3813_ (
  .A({ S6405 }),
  .B({ S6415 }),
  .Y({ S6418 })
);
NOR #() 
NOR_2216_ (
  .A({ S6405 }),
  .B({ S6415 }),
  .Y({ S6419 })
);
NAND #() 
NAND_3814_ (
  .A({ S6406 }),
  .B({ S6416 }),
  .Y({ S6420 })
);
NOR #() 
NOR_2217_ (
  .A({ S6417 }),
  .B({ S6419 }),
  .Y({ S6421 })
);
NAND #() 
NAND_3815_ (
  .A({ S6418 }),
  .B({ S6420 }),
  .Y({ S6422 })
);
NOR #() 
NOR_2218_ (
  .A({ S6403 }),
  .B({ S6422 }),
  .Y({ S6423 })
);
NAND #() 
NAND_3816_ (
  .A({ S6404 }),
  .B({ S6421 }),
  .Y({ S6424 })
);
NOR #() 
NOR_2219_ (
  .A({ S6404 }),
  .B({ S6421 }),
  .Y({ S6425 })
);
NAND #() 
NAND_3817_ (
  .A({ S6403 }),
  .B({ S6422 }),
  .Y({ S6426 })
);
NOR #() 
NOR_2220_ (
  .A({ S6423 }),
  .B({ S6425 }),
  .Y({ S6427 })
);
NAND #() 
NAND_3818_ (
  .A({ S6424 }),
  .B({ S6426 }),
  .Y({ S6428 })
);
NOR #() 
NOR_2221_ (
  .A({ S6402 }),
  .B({ S6428 }),
  .Y({ S6429 })
);
NAND #() 
NAND_3819_ (
  .A({ S6401 }),
  .B({ S6427 }),
  .Y({ S6430 })
);
NOR #() 
NOR_2222_ (
  .A({ S6401 }),
  .B({ S6427 }),
  .Y({ S6431 })
);
NAND #() 
NAND_3820_ (
  .A({ S6402 }),
  .B({ S6428 }),
  .Y({ S6432 })
);
NOR #() 
NOR_2223_ (
  .A({ S6429 }),
  .B({ S6431 }),
  .Y({ S6433 })
);
NAND #() 
NAND_3821_ (
  .A({ S6430 }),
  .B({ S6432 }),
  .Y({ S6434 })
);
NOR #() 
NOR_2224_ (
  .A({ S6383 }),
  .B({ S6434 }),
  .Y({ S6435 })
);
NAND #() 
NAND_3822_ (
  .A({ S6384 }),
  .B({ S6433 }),
  .Y({ S6436 })
);
NOR #() 
NOR_2225_ (
  .A({ S6384 }),
  .B({ S6433 }),
  .Y({ S6437 })
);
NAND #() 
NAND_3823_ (
  .A({ S6383 }),
  .B({ S6434 }),
  .Y({ S6438 })
);
NOR #() 
NOR_2226_ (
  .A({ S6435 }),
  .B({ S6437 }),
  .Y({ S6439 })
);
NAND #() 
NAND_3824_ (
  .A({ S6436 }),
  .B({ S6438 }),
  .Y({ S6440 })
);
NOR #() 
NOR_2227_ (
  .A({ S6382 }),
  .B({ S6440 }),
  .Y({ S6441 })
);
NAND #() 
NAND_3825_ (
  .A({ S6381 }),
  .B({ S6439 }),
  .Y({ S6442 })
);
NOR #() 
NOR_2228_ (
  .A({ S6381 }),
  .B({ S6439 }),
  .Y({ S6443 })
);
NAND #() 
NAND_3826_ (
  .A({ S6382 }),
  .B({ S6440 }),
  .Y({ S6444 })
);
NOR #() 
NOR_2229_ (
  .A({ S6441 }),
  .B({ S6443 }),
  .Y({ S6445 })
);
NAND #() 
NAND_3827_ (
  .A({ S6442 }),
  .B({ S6444 }),
  .Y({ S6446 })
);
NOR #() 
NOR_2230_ (
  .A({ S6349 }),
  .B({ S6446 }),
  .Y({ S6447 })
);
NAND #() 
NAND_3828_ (
  .A({ S6350 }),
  .B({ S6445 }),
  .Y({ S6448 })
);
NOR #() 
NOR_2231_ (
  .A({ S6350 }),
  .B({ S6445 }),
  .Y({ S6449 })
);
NAND #() 
NAND_3829_ (
  .A({ S6349 }),
  .B({ S6446 }),
  .Y({ S6450 })
);
NOR #() 
NOR_2232_ (
  .A({ S6447 }),
  .B({ S6449 }),
  .Y({ S6451 })
);
NAND #() 
NAND_3830_ (
  .A({ S6448 }),
  .B({ S6450 }),
  .Y({ S6452 })
);
NOR #() 
NOR_2233_ (
  .A({ S6255 }),
  .B({ S6452 }),
  .Y({ S6453 })
);
NAND #() 
NAND_3831_ (
  .A({ S6254 }),
  .B({ S6451 }),
  .Y({ S6454 })
);
NOR #() 
NOR_2234_ (
  .A({ S6254 }),
  .B({ S6451 }),
  .Y({ S6455 })
);
NAND #() 
NAND_3832_ (
  .A({ S6255 }),
  .B({ S6452 }),
  .Y({ S6456 })
);
NOR #() 
NOR_2235_ (
  .A({ S6453 }),
  .B({ S6455 }),
  .Y({ S6457 })
);
NAND #() 
NAND_3833_ (
  .A({ S6454 }),
  .B({ S6456 }),
  .Y({ S6458 })
);
NAND #() 
NAND_3834_ (
  .A({ S6347 }),
  .B({ S6458 }),
  .Y({ S6459 })
);
NOR #() 
NOR_2236_ (
  .A({ S6347 }),
  .B({ S6458 }),
  .Y({ S6460 })
);
NAND #() 
NAND_3835_ (
  .A({ S6348 }),
  .B({ S6457 }),
  .Y({ S6461 })
);
NAND #() 
NAND_3836_ (
  .A({ S6459 }),
  .B({ S6461 }),
  .Y({ S6462 })
);
NOT #() 
NOT_507_ (
  .A({ S6462 }),
  .Y({ S6463 })
);
NAND #() 
NAND_3837_ (
  .A({ S6333 }),
  .B({ S6463 }),
  .Y({ S6464 })
);
NOT #() 
NOT_508_ (
  .A({ S6464 }),
  .Y({ S6465 })
);
NAND #() 
NAND_3838_ (
  .A({ S6332 }),
  .B({ S6462 }),
  .Y({ S6466 })
);
NAND #() 
NAND_3839_ (
  .A({ S6464 }),
  .B({ S6466 }),
  .Y({ S6467 })
);
NOR #() 
NOR_2237_ (
  .A({ S6341 }),
  .B({ S6467 }),
  .Y({ S6468 })
);
NOT #() 
NOT_509_ (
  .A({ S6468 }),
  .Y({ S6469 })
);
NAND #() 
NAND_3840_ (
  .A({ S6341 }),
  .B({ S6467 }),
  .Y({ S6470 })
);
NAND #() 
NAND_3841_ (
  .A({ S6469 }),
  .B({ S6470 }),
  .Y({ S6471 })
);
NOR #() 
NOR_2238_ (
  .A({ S6337 }),
  .B({ S6471 }),
  .Y({ S6472 })
);
NAND #() 
NAND_3842_ (
  .A({ S6337 }),
  .B({ S6471 }),
  .Y({ S6473 })
);
NAND #() 
NAND_3843_ (
  .A({ S5948 }),
  .B({ S6473 }),
  .Y({ S6474 })
);
NOR #() 
NOR_2239_ (
  .A({ S6472 }),
  .B({ S6474 }),
  .Y({ S6475 })
);
NOR #() 
NOR_2240_ (
  .A({ S6345 }),
  .B({ S6475 }),
  .Y({ S6476 })
);
NAND #() 
NAND_3844_ (
  .A({ S6346 }),
  .B({ S6476 }),
  .Y({ S290 })
);
NOR #() 
NOR_2241_ (
  .A({ S3899 }),
  .B({ S4313 }),
  .Y({ S6477 })
);
NAND #() 
NAND_3845_ (
  .A({ datapath_multdivunit_outmdu1_9 }),
  .B({ S5950 }),
  .Y({ S6478 })
);
NOR #() 
NOR_2242_ (
  .A({ S6468 }),
  .B({ S6472 }),
  .Y({ S6479 })
);
NOR #() 
NOR_2243_ (
  .A({ S6447 }),
  .B({ S6453 }),
  .Y({ S6480 })
);
NOR #() 
NOR_2244_ (
  .A({ S1220 }),
  .B({ S2518 }),
  .Y({ S6481 })
);
NAND #() 
NAND_3846_ (
  .A({ datapath_addsubunit_in1_0 }),
  .B({ S2517 }),
  .Y({ S6482 })
);
NOR #() 
NOR_2245_ (
  .A({ S6371 }),
  .B({ S6377 }),
  .Y({ S6483 })
);
NAND #() 
NAND_3847_ (
  .A({ S6372 }),
  .B({ S6378 }),
  .Y({ S6484 })
);
NOR #() 
NOR_2246_ (
  .A({ S6482 }),
  .B({ S6483 }),
  .Y({ S6485 })
);
NOT #() 
NOT_510_ (
  .A({ S6485 }),
  .Y({ S6486 })
);
NOR #() 
NOR_2247_ (
  .A({ S6481 }),
  .B({ S6484 }),
  .Y({ S6487 })
);
NAND #() 
NAND_3848_ (
  .A({ S6482 }),
  .B({ S6483 }),
  .Y({ S6488 })
);
NOR #() 
NOR_2248_ (
  .A({ S6485 }),
  .B({ S6487 }),
  .Y({ S6489 })
);
NAND #() 
NAND_3849_ (
  .A({ S6486 }),
  .B({ S6488 }),
  .Y({ S6490 })
);
NOR #() 
NOR_2249_ (
  .A({ S6435 }),
  .B({ S6441 }),
  .Y({ S6491 })
);
NAND #() 
NAND_3850_ (
  .A({ S6436 }),
  .B({ S6442 }),
  .Y({ S6492 })
);
NOR #() 
NOR_2250_ (
  .A({ S6359 }),
  .B({ S6363 }),
  .Y({ S6493 })
);
NAND #() 
NAND_3851_ (
  .A({ S6360 }),
  .B({ S6364 }),
  .Y({ S6494 })
);
NOR #() 
NOR_2251_ (
  .A({ S1168 }),
  .B({ S2418 }),
  .Y({ S6495 })
);
NAND #() 
NAND_3852_ (
  .A({ datapath_addsubunit_in1_1 }),
  .B({ S2417 }),
  .Y({ S6496 })
);
NOR #() 
NOR_2252_ (
  .A({ S1065 }),
  .B({ S2206 }),
  .Y({ S6497 })
);
NAND #() 
NAND_3853_ (
  .A({ datapath_addsubunit_in1_3 }),
  .B({ S2205 }),
  .Y({ S6498 })
);
NOR #() 
NOR_2253_ (
  .A({ S6357 }),
  .B({ S6497 }),
  .Y({ S6499 })
);
NAND #() 
NAND_3854_ (
  .A({ S6358 }),
  .B({ S6498 }),
  .Y({ S6500 })
);
NOR #() 
NOR_2254_ (
  .A({ S1065 }),
  .B({ S2312 }),
  .Y({ S6501 })
);
NAND #() 
NAND_3855_ (
  .A({ datapath_addsubunit_in1_3 }),
  .B({ S2311 }),
  .Y({ S6502 })
);
NOR #() 
NOR_2255_ (
  .A({ S6358 }),
  .B({ S6498 }),
  .Y({ S6503 })
);
NAND #() 
NAND_3856_ (
  .A({ S6357 }),
  .B({ S6497 }),
  .Y({ S6504 })
);
NOR #() 
NOR_2256_ (
  .A({ S6499 }),
  .B({ S6503 }),
  .Y({ S6505 })
);
NAND #() 
NAND_3857_ (
  .A({ S6500 }),
  .B({ S6504 }),
  .Y({ S6506 })
);
NOR #() 
NOR_2257_ (
  .A({ S6496 }),
  .B({ S6506 }),
  .Y({ S6507 })
);
NAND #() 
NAND_3858_ (
  .A({ S6495 }),
  .B({ S6505 }),
  .Y({ S6508 })
);
NOR #() 
NOR_2258_ (
  .A({ S6495 }),
  .B({ S6505 }),
  .Y({ S6509 })
);
NAND #() 
NAND_3859_ (
  .A({ S6496 }),
  .B({ S6506 }),
  .Y({ S6510 })
);
NOR #() 
NOR_2259_ (
  .A({ S6507 }),
  .B({ S6509 }),
  .Y({ S6511 })
);
NAND #() 
NAND_3860_ (
  .A({ S6508 }),
  .B({ S6510 }),
  .Y({ S6512 })
);
NOR #() 
NOR_2260_ (
  .A({ S6393 }),
  .B({ S6397 }),
  .Y({ S6513 })
);
NAND #() 
NAND_3861_ (
  .A({ S6394 }),
  .B({ S6398 }),
  .Y({ S6514 })
);
NOR #() 
NOR_2261_ (
  .A({ S6512 }),
  .B({ S6513 }),
  .Y({ S6515 })
);
NAND #() 
NAND_3862_ (
  .A({ S6511 }),
  .B({ S6514 }),
  .Y({ S6516 })
);
NOR #() 
NOR_2262_ (
  .A({ S6511 }),
  .B({ S6514 }),
  .Y({ S6517 })
);
NAND #() 
NAND_3863_ (
  .A({ S6512 }),
  .B({ S6513 }),
  .Y({ S6518 })
);
NOR #() 
NOR_2263_ (
  .A({ S6515 }),
  .B({ S6517 }),
  .Y({ S6519 })
);
NAND #() 
NAND_3864_ (
  .A({ S6516 }),
  .B({ S6518 }),
  .Y({ S6520 })
);
NOR #() 
NOR_2264_ (
  .A({ S6494 }),
  .B({ S6519 }),
  .Y({ S6521 })
);
NAND #() 
NAND_3865_ (
  .A({ S6493 }),
  .B({ S6520 }),
  .Y({ S6522 })
);
NOR #() 
NOR_2265_ (
  .A({ S6493 }),
  .B({ S6520 }),
  .Y({ S6523 })
);
NAND #() 
NAND_3866_ (
  .A({ S6494 }),
  .B({ S6519 }),
  .Y({ S6524 })
);
NOR #() 
NOR_2266_ (
  .A({ S6521 }),
  .B({ S6523 }),
  .Y({ S6525 })
);
NAND #() 
NAND_3867_ (
  .A({ S6522 }),
  .B({ S6524 }),
  .Y({ S6526 })
);
NOR #() 
NOR_2267_ (
  .A({ S6423 }),
  .B({ S6429 }),
  .Y({ S6527 })
);
NAND #() 
NAND_3868_ (
  .A({ S6424 }),
  .B({ S6430 }),
  .Y({ S6528 })
);
NOR #() 
NOR_2268_ (
  .A({ S1013 }),
  .B({ S2107 }),
  .Y({ S6529 })
);
NAND #() 
NAND_3869_ (
  .A({ datapath_addsubunit_in1_4 }),
  .B({ S2106 }),
  .Y({ S6530 })
);
NOR #() 
NOR_2269_ (
  .A({ S910 }),
  .B({ S1953 }),
  .Y({ S6531 })
);
NAND #() 
NAND_3870_ (
  .A({ datapath_addsubunit_in1_6 }),
  .B({ S1952 }),
  .Y({ S6532 })
);
NOR #() 
NOR_2270_ (
  .A({ S6391 }),
  .B({ S6531 }),
  .Y({ S6533 })
);
NAND #() 
NAND_3871_ (
  .A({ S6392 }),
  .B({ S6532 }),
  .Y({ S6534 })
);
NOR #() 
NOR_2271_ (
  .A({ S910 }),
  .B({ S1598 }),
  .Y({ S6535 })
);
NAND #() 
NAND_3872_ (
  .A({ datapath_addsubunit_in1_6 }),
  .B({ S1597 }),
  .Y({ S6536 })
);
NOR #() 
NOR_2272_ (
  .A({ S6392 }),
  .B({ S6532 }),
  .Y({ S6537 })
);
NAND #() 
NAND_3873_ (
  .A({ S6391 }),
  .B({ S6531 }),
  .Y({ S6538 })
);
NOR #() 
NOR_2273_ (
  .A({ S6533 }),
  .B({ S6537 }),
  .Y({ S6539 })
);
NAND #() 
NAND_3874_ (
  .A({ S6534 }),
  .B({ S6538 }),
  .Y({ S6540 })
);
NOR #() 
NOR_2274_ (
  .A({ S6530 }),
  .B({ S6540 }),
  .Y({ S6541 })
);
NAND #() 
NAND_3875_ (
  .A({ S6529 }),
  .B({ S6539 }),
  .Y({ S6542 })
);
NOR #() 
NOR_2275_ (
  .A({ S6529 }),
  .B({ S6539 }),
  .Y({ S6543 })
);
NAND #() 
NAND_3876_ (
  .A({ S6530 }),
  .B({ S6540 }),
  .Y({ S6544 })
);
NOR #() 
NOR_2276_ (
  .A({ S6541 }),
  .B({ S6543 }),
  .Y({ S6545 })
);
NAND #() 
NAND_3877_ (
  .A({ S6542 }),
  .B({ S6544 }),
  .Y({ S6546 })
);
NOR #() 
NOR_2277_ (
  .A({ S6413 }),
  .B({ S6417 }),
  .Y({ S6547 })
);
NAND #() 
NAND_3878_ (
  .A({ S6414 }),
  .B({ S6418 }),
  .Y({ S6548 })
);
NOR #() 
NOR_2278_ (
  .A({ S858 }),
  .B({ S1849 }),
  .Y({ S6549 })
);
NAND #() 
NAND_3879_ (
  .A({ datapath_addsubunit_in1_7 }),
  .B({ S1848 }),
  .Y({ S6550 })
);
NOR #() 
NOR_2279_ (
  .A({ S754 }),
  .B({ S1516 }),
  .Y({ S6551 })
);
NAND #() 
NAND_3880_ (
  .A({ datapath_addsubunit_in1_9 }),
  .B({ S1515 }),
  .Y({ S6552 })
);
NOR #() 
NOR_2280_ (
  .A({ S6411 }),
  .B({ S6551 }),
  .Y({ S6553 })
);
NAND #() 
NAND_3881_ (
  .A({ S6412 }),
  .B({ S6552 }),
  .Y({ S6554 })
);
NOR #() 
NOR_2281_ (
  .A({ S754 }),
  .B({ S1746 }),
  .Y({ S6555 })
);
NAND #() 
NAND_3882_ (
  .A({ datapath_addsubunit_in1_9 }),
  .B({ S1745 }),
  .Y({ S6556 })
);
NOR #() 
NOR_2282_ (
  .A({ S6412 }),
  .B({ S6552 }),
  .Y({ S6557 })
);
NAND #() 
NAND_3883_ (
  .A({ S6411 }),
  .B({ S6551 }),
  .Y({ S6558 })
);
NOR #() 
NOR_2283_ (
  .A({ S6553 }),
  .B({ S6557 }),
  .Y({ S6559 })
);
NAND #() 
NAND_3884_ (
  .A({ S6554 }),
  .B({ S6558 }),
  .Y({ S6560 })
);
NOR #() 
NOR_2284_ (
  .A({ S6550 }),
  .B({ S6560 }),
  .Y({ S6561 })
);
NAND #() 
NAND_3885_ (
  .A({ S6549 }),
  .B({ S6559 }),
  .Y({ S6562 })
);
NOR #() 
NOR_2285_ (
  .A({ S6549 }),
  .B({ S6559 }),
  .Y({ S6563 })
);
NAND #() 
NAND_3886_ (
  .A({ S6550 }),
  .B({ S6560 }),
  .Y({ S6564 })
);
NOR #() 
NOR_2286_ (
  .A({ S6561 }),
  .B({ S6563 }),
  .Y({ S6565 })
);
NAND #() 
NAND_3887_ (
  .A({ S6562 }),
  .B({ S6564 }),
  .Y({ S6566 })
);
NOR #() 
NOR_2287_ (
  .A({ S6547 }),
  .B({ S6566 }),
  .Y({ S6567 })
);
NAND #() 
NAND_3888_ (
  .A({ S6548 }),
  .B({ S6565 }),
  .Y({ S6568 })
);
NOR #() 
NOR_2288_ (
  .A({ S6548 }),
  .B({ S6565 }),
  .Y({ S6569 })
);
NAND #() 
NAND_3889_ (
  .A({ S6547 }),
  .B({ S6566 }),
  .Y({ S6570 })
);
NOR #() 
NOR_2289_ (
  .A({ S6567 }),
  .B({ S6569 }),
  .Y({ S6571 })
);
NAND #() 
NAND_3890_ (
  .A({ S6568 }),
  .B({ S6570 }),
  .Y({ S6572 })
);
NOR #() 
NOR_2290_ (
  .A({ S6546 }),
  .B({ S6572 }),
  .Y({ S6573 })
);
NAND #() 
NAND_3891_ (
  .A({ S6545 }),
  .B({ S6571 }),
  .Y({ S6574 })
);
NOR #() 
NOR_2291_ (
  .A({ S6545 }),
  .B({ S6571 }),
  .Y({ S6575 })
);
NAND #() 
NAND_3892_ (
  .A({ S6546 }),
  .B({ S6572 }),
  .Y({ S6576 })
);
NOR #() 
NOR_2292_ (
  .A({ S6573 }),
  .B({ S6575 }),
  .Y({ S6577 })
);
NAND #() 
NAND_3893_ (
  .A({ S6574 }),
  .B({ S6576 }),
  .Y({ S6578 })
);
NOR #() 
NOR_2293_ (
  .A({ S6527 }),
  .B({ S6578 }),
  .Y({ S6579 })
);
NAND #() 
NAND_3894_ (
  .A({ S6528 }),
  .B({ S6577 }),
  .Y({ S6580 })
);
NOR #() 
NOR_2294_ (
  .A({ S6528 }),
  .B({ S6577 }),
  .Y({ S6581 })
);
NAND #() 
NAND_3895_ (
  .A({ S6527 }),
  .B({ S6578 }),
  .Y({ S6582 })
);
NOR #() 
NOR_2295_ (
  .A({ S6579 }),
  .B({ S6581 }),
  .Y({ S6583 })
);
NAND #() 
NAND_3896_ (
  .A({ S6580 }),
  .B({ S6582 }),
  .Y({ S6584 })
);
NOR #() 
NOR_2296_ (
  .A({ S6526 }),
  .B({ S6584 }),
  .Y({ S6585 })
);
NAND #() 
NAND_3897_ (
  .A({ S6525 }),
  .B({ S6583 }),
  .Y({ S6586 })
);
NOR #() 
NOR_2297_ (
  .A({ S6525 }),
  .B({ S6583 }),
  .Y({ S6587 })
);
NAND #() 
NAND_3898_ (
  .A({ S6526 }),
  .B({ S6584 }),
  .Y({ S6588 })
);
NOR #() 
NOR_2298_ (
  .A({ S6585 }),
  .B({ S6587 }),
  .Y({ S6589 })
);
NAND #() 
NAND_3899_ (
  .A({ S6586 }),
  .B({ S6588 }),
  .Y({ S6590 })
);
NOR #() 
NOR_2299_ (
  .A({ S6491 }),
  .B({ S6590 }),
  .Y({ S6591 })
);
NAND #() 
NAND_3900_ (
  .A({ S6492 }),
  .B({ S6589 }),
  .Y({ S6592 })
);
NOR #() 
NOR_2300_ (
  .A({ S6492 }),
  .B({ S6589 }),
  .Y({ S6593 })
);
NAND #() 
NAND_3901_ (
  .A({ S6491 }),
  .B({ S6590 }),
  .Y({ S6594 })
);
NOR #() 
NOR_2301_ (
  .A({ S6591 }),
  .B({ S6593 }),
  .Y({ S6595 })
);
NAND #() 
NAND_3902_ (
  .A({ S6592 }),
  .B({ S6594 }),
  .Y({ S6596 })
);
NOR #() 
NOR_2302_ (
  .A({ S6490 }),
  .B({ S6596 }),
  .Y({ S6597 })
);
NAND #() 
NAND_3903_ (
  .A({ S6489 }),
  .B({ S6595 }),
  .Y({ S6598 })
);
NAND #() 
NAND_3904_ (
  .A({ S6490 }),
  .B({ S6596 }),
  .Y({ S6599 })
);
NAND #() 
NAND_3905_ (
  .A({ S6598 }),
  .B({ S6599 }),
  .Y({ S6600 })
);
NAND #() 
NAND_3906_ (
  .A({ S6480 }),
  .B({ S6600 }),
  .Y({ S6601 })
);
NOT #() 
NOT_511_ (
  .A({ S6601 }),
  .Y({ S6602 })
);
NOR #() 
NOR_2303_ (
  .A({ S6480 }),
  .B({ S6600 }),
  .Y({ S6603 })
);
NOT #() 
NOT_512_ (
  .A({ S6603 }),
  .Y({ S6604 })
);
NOR #() 
NOR_2304_ (
  .A({ S6602 }),
  .B({ S6603 }),
  .Y({ S6605 })
);
NAND #() 
NAND_3907_ (
  .A({ S6601 }),
  .B({ S6604 }),
  .Y({ S6606 })
);
NOR #() 
NOR_2305_ (
  .A({ S6461 }),
  .B({ S6606 }),
  .Y({ S6607 })
);
NAND #() 
NAND_3908_ (
  .A({ S6460 }),
  .B({ S6605 }),
  .Y({ S6608 })
);
NOR #() 
NOR_2306_ (
  .A({ S6460 }),
  .B({ S6605 }),
  .Y({ S6609 })
);
NAND #() 
NAND_3909_ (
  .A({ S6461 }),
  .B({ S6606 }),
  .Y({ S6610 })
);
NOR #() 
NOR_2307_ (
  .A({ S6607 }),
  .B({ S6609 }),
  .Y({ S6611 })
);
NAND #() 
NAND_3910_ (
  .A({ S6608 }),
  .B({ S6610 }),
  .Y({ S6612 })
);
NAND #() 
NAND_3911_ (
  .A({ S6465 }),
  .B({ S6611 }),
  .Y({ S6613 })
);
NAND #() 
NAND_3912_ (
  .A({ S6464 }),
  .B({ S6612 }),
  .Y({ S6614 })
);
NAND #() 
NAND_3913_ (
  .A({ S6613 }),
  .B({ S6614 }),
  .Y({ S6615 })
);
NOR #() 
NOR_2308_ (
  .A({ S6479 }),
  .B({ S6615 }),
  .Y({ S6616 })
);
NOT #() 
NOT_513_ (
  .A({ S6616 }),
  .Y({ S6617 })
);
NAND #() 
NAND_3914_ (
  .A({ S6479 }),
  .B({ S6615 }),
  .Y({ S6618 })
);
NAND #() 
NAND_3915_ (
  .A({ S5948 }),
  .B({ S6618 }),
  .Y({ S6619 })
);
NOR #() 
NOR_2309_ (
  .A({ S6616 }),
  .B({ S6619 }),
  .Y({ S6620 })
);
NOR #() 
NOR_2310_ (
  .A({ S6477 }),
  .B({ S6620 }),
  .Y({ S6621 })
);
NAND #() 
NAND_3916_ (
  .A({ S6478 }),
  .B({ S6621 }),
  .Y({ S291 })
);
NOR #() 
NOR_2311_ (
  .A({ S3899 }),
  .B({ S4195 }),
  .Y({ S6622 })
);
NAND #() 
NAND_3917_ (
  .A({ datapath_multdivunit_outmdu1_10 }),
  .B({ S5950 }),
  .Y({ S6623 })
);
NAND #() 
NAND_3918_ (
  .A({ S6613 }),
  .B({ S6617 }),
  .Y({ S6624 })
);
NOR #() 
NOR_2312_ (
  .A({ S6591 }),
  .B({ S6597 }),
  .Y({ S6625 })
);
NAND #() 
NAND_3919_ (
  .A({ S6592 }),
  .B({ S6598 }),
  .Y({ S6626 })
);
NOR #() 
NOR_2313_ (
  .A({ S1220 }),
  .B({ S2618 }),
  .Y({ S6627 })
);
NAND #() 
NAND_3920_ (
  .A({ datapath_addsubunit_in1_0 }),
  .B({ S2617 }),
  .Y({ S6628 })
);
NOR #() 
NOR_2314_ (
  .A({ S1168 }),
  .B({ S2518 }),
  .Y({ S6629 })
);
NAND #() 
NAND_3921_ (
  .A({ datapath_addsubunit_in1_1 }),
  .B({ S2517 }),
  .Y({ S6630 })
);
NOR #() 
NOR_2315_ (
  .A({ S6627 }),
  .B({ S6629 }),
  .Y({ S6631 })
);
NAND #() 
NAND_3922_ (
  .A({ S6628 }),
  .B({ S6630 }),
  .Y({ S6632 })
);
NOR #() 
NOR_2316_ (
  .A({ S1168 }),
  .B({ S2618 }),
  .Y({ S6633 })
);
NAND #() 
NAND_3923_ (
  .A({ datapath_addsubunit_in1_1 }),
  .B({ S2617 }),
  .Y({ S6634 })
);
NOR #() 
NOR_2317_ (
  .A({ S6482 }),
  .B({ S6634 }),
  .Y({ S6635 })
);
NAND #() 
NAND_3924_ (
  .A({ S6481 }),
  .B({ S6633 }),
  .Y({ S6636 })
);
NOR #() 
NOR_2318_ (
  .A({ S6631 }),
  .B({ S6635 }),
  .Y({ S6637 })
);
NAND #() 
NAND_3925_ (
  .A({ S6632 }),
  .B({ S6636 }),
  .Y({ S6638 })
);
NOR #() 
NOR_2319_ (
  .A({ S6515 }),
  .B({ S6523 }),
  .Y({ S6639 })
);
NAND #() 
NAND_3926_ (
  .A({ S6516 }),
  .B({ S6524 }),
  .Y({ S6640 })
);
NOR #() 
NOR_2320_ (
  .A({ S6637 }),
  .B({ S6640 }),
  .Y({ S6641 })
);
NAND #() 
NAND_3927_ (
  .A({ S6638 }),
  .B({ S6639 }),
  .Y({ S6642 })
);
NOR #() 
NOR_2321_ (
  .A({ S6638 }),
  .B({ S6639 }),
  .Y({ S6643 })
);
NAND #() 
NAND_3928_ (
  .A({ S6637 }),
  .B({ S6640 }),
  .Y({ S6644 })
);
NOR #() 
NOR_2322_ (
  .A({ S6641 }),
  .B({ S6643 }),
  .Y({ S6645 })
);
NAND #() 
NAND_3929_ (
  .A({ S6642 }),
  .B({ S6644 }),
  .Y({ S6646 })
);
NOR #() 
NOR_2323_ (
  .A({ S6579 }),
  .B({ S6585 }),
  .Y({ S6647 })
);
NAND #() 
NAND_3930_ (
  .A({ S6580 }),
  .B({ S6586 }),
  .Y({ S6648 })
);
NOR #() 
NOR_2324_ (
  .A({ S6503 }),
  .B({ S6507 }),
  .Y({ S6649 })
);
NAND #() 
NAND_3931_ (
  .A({ S6504 }),
  .B({ S6508 }),
  .Y({ S6650 })
);
NOR #() 
NOR_2325_ (
  .A({ S1116 }),
  .B({ S2418 }),
  .Y({ S6651 })
);
NAND #() 
NAND_3932_ (
  .A({ datapath_addsubunit_in1_2 }),
  .B({ S2417 }),
  .Y({ S6652 })
);
NOR #() 
NOR_2326_ (
  .A({ S1013 }),
  .B({ S2206 }),
  .Y({ S6653 })
);
NAND #() 
NAND_3933_ (
  .A({ datapath_addsubunit_in1_4 }),
  .B({ S2205 }),
  .Y({ S6654 })
);
NOR #() 
NOR_2327_ (
  .A({ S6501 }),
  .B({ S6653 }),
  .Y({ S6655 })
);
NAND #() 
NAND_3934_ (
  .A({ S6502 }),
  .B({ S6654 }),
  .Y({ S6656 })
);
NOR #() 
NOR_2328_ (
  .A({ S1013 }),
  .B({ S2312 }),
  .Y({ S6657 })
);
NAND #() 
NAND_3935_ (
  .A({ datapath_addsubunit_in1_4 }),
  .B({ S2311 }),
  .Y({ S6658 })
);
NOR #() 
NOR_2329_ (
  .A({ S6502 }),
  .B({ S6654 }),
  .Y({ S6659 })
);
NAND #() 
NAND_3936_ (
  .A({ S6501 }),
  .B({ S6653 }),
  .Y({ S6660 })
);
NOR #() 
NOR_2330_ (
  .A({ S6655 }),
  .B({ S6659 }),
  .Y({ S6661 })
);
NAND #() 
NAND_3937_ (
  .A({ S6656 }),
  .B({ S6660 }),
  .Y({ S6662 })
);
NOR #() 
NOR_2331_ (
  .A({ S6652 }),
  .B({ S6662 }),
  .Y({ S6663 })
);
NAND #() 
NAND_3938_ (
  .A({ S6651 }),
  .B({ S6661 }),
  .Y({ S6664 })
);
NOR #() 
NOR_2332_ (
  .A({ S6651 }),
  .B({ S6661 }),
  .Y({ S6665 })
);
NAND #() 
NAND_3939_ (
  .A({ S6652 }),
  .B({ S6662 }),
  .Y({ S6666 })
);
NOR #() 
NOR_2333_ (
  .A({ S6663 }),
  .B({ S6665 }),
  .Y({ S6667 })
);
NAND #() 
NAND_3940_ (
  .A({ S6664 }),
  .B({ S6666 }),
  .Y({ S6668 })
);
NOR #() 
NOR_2334_ (
  .A({ S6537 }),
  .B({ S6541 }),
  .Y({ S6669 })
);
NAND #() 
NAND_3941_ (
  .A({ S6538 }),
  .B({ S6542 }),
  .Y({ S6670 })
);
NOR #() 
NOR_2335_ (
  .A({ S6668 }),
  .B({ S6669 }),
  .Y({ S6671 })
);
NAND #() 
NAND_3942_ (
  .A({ S6667 }),
  .B({ S6670 }),
  .Y({ S6672 })
);
NOR #() 
NOR_2336_ (
  .A({ S6667 }),
  .B({ S6670 }),
  .Y({ S6673 })
);
NAND #() 
NAND_3943_ (
  .A({ S6668 }),
  .B({ S6669 }),
  .Y({ S6674 })
);
NOR #() 
NOR_2337_ (
  .A({ S6671 }),
  .B({ S6673 }),
  .Y({ S6675 })
);
NAND #() 
NAND_3944_ (
  .A({ S6672 }),
  .B({ S6674 }),
  .Y({ S6676 })
);
NOR #() 
NOR_2338_ (
  .A({ S6650 }),
  .B({ S6675 }),
  .Y({ S6677 })
);
NAND #() 
NAND_3945_ (
  .A({ S6649 }),
  .B({ S6676 }),
  .Y({ S6678 })
);
NOR #() 
NOR_2339_ (
  .A({ S6649 }),
  .B({ S6676 }),
  .Y({ S6679 })
);
NAND #() 
NAND_3946_ (
  .A({ S6650 }),
  .B({ S6675 }),
  .Y({ S6680 })
);
NOR #() 
NOR_2340_ (
  .A({ S6677 }),
  .B({ S6679 }),
  .Y({ S6681 })
);
NAND #() 
NAND_3947_ (
  .A({ S6678 }),
  .B({ S6680 }),
  .Y({ S6682 })
);
NOR #() 
NOR_2341_ (
  .A({ S6567 }),
  .B({ S6573 }),
  .Y({ S6683 })
);
NAND #() 
NAND_3948_ (
  .A({ S6568 }),
  .B({ S6574 }),
  .Y({ S6684 })
);
NOR #() 
NOR_2342_ (
  .A({ S963 }),
  .B({ S2107 }),
  .Y({ S6685 })
);
NAND #() 
NAND_3949_ (
  .A({ datapath_addsubunit_in1_5 }),
  .B({ S2106 }),
  .Y({ S6686 })
);
NOR #() 
NOR_2343_ (
  .A({ S858 }),
  .B({ S1953 }),
  .Y({ S6687 })
);
NAND #() 
NAND_3950_ (
  .A({ datapath_addsubunit_in1_7 }),
  .B({ S1952 }),
  .Y({ S6688 })
);
NOR #() 
NOR_2344_ (
  .A({ S6535 }),
  .B({ S6687 }),
  .Y({ S6689 })
);
NAND #() 
NAND_3951_ (
  .A({ S6536 }),
  .B({ S6688 }),
  .Y({ S6690 })
);
NOR #() 
NOR_2345_ (
  .A({ S858 }),
  .B({ S1598 }),
  .Y({ S6691 })
);
NAND #() 
NAND_3952_ (
  .A({ datapath_addsubunit_in1_7 }),
  .B({ S1597 }),
  .Y({ S6692 })
);
NOR #() 
NOR_2346_ (
  .A({ S6536 }),
  .B({ S6688 }),
  .Y({ S6693 })
);
NAND #() 
NAND_3953_ (
  .A({ S6535 }),
  .B({ S6687 }),
  .Y({ S6694 })
);
NOR #() 
NOR_2347_ (
  .A({ S6689 }),
  .B({ S6693 }),
  .Y({ S6695 })
);
NAND #() 
NAND_3954_ (
  .A({ S6690 }),
  .B({ S6694 }),
  .Y({ S6696 })
);
NOR #() 
NOR_2348_ (
  .A({ S6686 }),
  .B({ S6696 }),
  .Y({ S6697 })
);
NAND #() 
NAND_3955_ (
  .A({ S6685 }),
  .B({ S6695 }),
  .Y({ S6698 })
);
NOR #() 
NOR_2349_ (
  .A({ S6685 }),
  .B({ S6695 }),
  .Y({ S6699 })
);
NAND #() 
NAND_3956_ (
  .A({ S6686 }),
  .B({ S6696 }),
  .Y({ S6700 })
);
NOR #() 
NOR_2350_ (
  .A({ S6697 }),
  .B({ S6699 }),
  .Y({ S6701 })
);
NAND #() 
NAND_3957_ (
  .A({ S6698 }),
  .B({ S6700 }),
  .Y({ S6702 })
);
NOR #() 
NOR_2351_ (
  .A({ S6557 }),
  .B({ S6561 }),
  .Y({ S6703 })
);
NAND #() 
NAND_3958_ (
  .A({ S6558 }),
  .B({ S6562 }),
  .Y({ S6704 })
);
NOR #() 
NOR_2352_ (
  .A({ S805 }),
  .B({ S1849 }),
  .Y({ S6705 })
);
NAND #() 
NAND_3959_ (
  .A({ datapath_addsubunit_in1_8 }),
  .B({ S1848 }),
  .Y({ S6706 })
);
NOR #() 
NOR_2353_ (
  .A({ S702 }),
  .B({ S1516 }),
  .Y({ S6707 })
);
NAND #() 
NAND_3960_ (
  .A({ datapath_addsubunit_in1_10 }),
  .B({ S1515 }),
  .Y({ S6708 })
);
NOR #() 
NOR_2354_ (
  .A({ S6555 }),
  .B({ S6707 }),
  .Y({ S6709 })
);
NAND #() 
NAND_3961_ (
  .A({ S6556 }),
  .B({ S6708 }),
  .Y({ S6710 })
);
NOR #() 
NOR_2355_ (
  .A({ S702 }),
  .B({ S1746 }),
  .Y({ S6711 })
);
NAND #() 
NAND_3962_ (
  .A({ datapath_addsubunit_in1_10 }),
  .B({ S1745 }),
  .Y({ S6712 })
);
NOR #() 
NOR_2356_ (
  .A({ S6556 }),
  .B({ S6708 }),
  .Y({ S6713 })
);
NAND #() 
NAND_3963_ (
  .A({ S6555 }),
  .B({ S6707 }),
  .Y({ S6714 })
);
NOR #() 
NOR_2357_ (
  .A({ S6709 }),
  .B({ S6713 }),
  .Y({ S6715 })
);
NAND #() 
NAND_3964_ (
  .A({ S6710 }),
  .B({ S6714 }),
  .Y({ S6716 })
);
NOR #() 
NOR_2358_ (
  .A({ S6706 }),
  .B({ S6716 }),
  .Y({ S6717 })
);
NAND #() 
NAND_3965_ (
  .A({ S6705 }),
  .B({ S6715 }),
  .Y({ S6718 })
);
NOR #() 
NOR_2359_ (
  .A({ S6705 }),
  .B({ S6715 }),
  .Y({ S6719 })
);
NAND #() 
NAND_3966_ (
  .A({ S6706 }),
  .B({ S6716 }),
  .Y({ S6720 })
);
NOR #() 
NOR_2360_ (
  .A({ S6717 }),
  .B({ S6719 }),
  .Y({ S6721 })
);
NAND #() 
NAND_3967_ (
  .A({ S6718 }),
  .B({ S6720 }),
  .Y({ S6722 })
);
NOR #() 
NOR_2361_ (
  .A({ S6703 }),
  .B({ S6722 }),
  .Y({ S6723 })
);
NAND #() 
NAND_3968_ (
  .A({ S6704 }),
  .B({ S6721 }),
  .Y({ S6724 })
);
NOR #() 
NOR_2362_ (
  .A({ S6704 }),
  .B({ S6721 }),
  .Y({ S6725 })
);
NAND #() 
NAND_3969_ (
  .A({ S6703 }),
  .B({ S6722 }),
  .Y({ S6726 })
);
NOR #() 
NOR_2363_ (
  .A({ S6723 }),
  .B({ S6725 }),
  .Y({ S6727 })
);
NAND #() 
NAND_3970_ (
  .A({ S6724 }),
  .B({ S6726 }),
  .Y({ S6728 })
);
NOR #() 
NOR_2364_ (
  .A({ S6702 }),
  .B({ S6728 }),
  .Y({ S6729 })
);
NAND #() 
NAND_3971_ (
  .A({ S6701 }),
  .B({ S6727 }),
  .Y({ S6730 })
);
NOR #() 
NOR_2365_ (
  .A({ S6701 }),
  .B({ S6727 }),
  .Y({ S6731 })
);
NAND #() 
NAND_3972_ (
  .A({ S6702 }),
  .B({ S6728 }),
  .Y({ S6732 })
);
NOR #() 
NOR_2366_ (
  .A({ S6729 }),
  .B({ S6731 }),
  .Y({ S6733 })
);
NAND #() 
NAND_3973_ (
  .A({ S6730 }),
  .B({ S6732 }),
  .Y({ S6734 })
);
NOR #() 
NOR_2367_ (
  .A({ S6683 }),
  .B({ S6734 }),
  .Y({ S6735 })
);
NAND #() 
NAND_3974_ (
  .A({ S6684 }),
  .B({ S6733 }),
  .Y({ S6736 })
);
NOR #() 
NOR_2368_ (
  .A({ S6684 }),
  .B({ S6733 }),
  .Y({ S6737 })
);
NAND #() 
NAND_3975_ (
  .A({ S6683 }),
  .B({ S6734 }),
  .Y({ S6738 })
);
NOR #() 
NOR_2369_ (
  .A({ S6735 }),
  .B({ S6737 }),
  .Y({ S6739 })
);
NAND #() 
NAND_3976_ (
  .A({ S6736 }),
  .B({ S6738 }),
  .Y({ S6740 })
);
NOR #() 
NOR_2370_ (
  .A({ S6682 }),
  .B({ S6740 }),
  .Y({ S6741 })
);
NAND #() 
NAND_3977_ (
  .A({ S6681 }),
  .B({ S6739 }),
  .Y({ S6742 })
);
NOR #() 
NOR_2371_ (
  .A({ S6681 }),
  .B({ S6739 }),
  .Y({ S6743 })
);
NAND #() 
NAND_3978_ (
  .A({ S6682 }),
  .B({ S6740 }),
  .Y({ S6744 })
);
NOR #() 
NOR_2372_ (
  .A({ S6741 }),
  .B({ S6743 }),
  .Y({ S6745 })
);
NAND #() 
NAND_3979_ (
  .A({ S6742 }),
  .B({ S6744 }),
  .Y({ S6746 })
);
NOR #() 
NOR_2373_ (
  .A({ S6647 }),
  .B({ S6746 }),
  .Y({ S6747 })
);
NAND #() 
NAND_3980_ (
  .A({ S6648 }),
  .B({ S6745 }),
  .Y({ S6748 })
);
NOR #() 
NOR_2374_ (
  .A({ S6648 }),
  .B({ S6745 }),
  .Y({ S6749 })
);
NAND #() 
NAND_3981_ (
  .A({ S6647 }),
  .B({ S6746 }),
  .Y({ S6750 })
);
NOR #() 
NOR_2375_ (
  .A({ S6747 }),
  .B({ S6749 }),
  .Y({ S6751 })
);
NAND #() 
NAND_3982_ (
  .A({ S6748 }),
  .B({ S6750 }),
  .Y({ S6752 })
);
NOR #() 
NOR_2376_ (
  .A({ S6646 }),
  .B({ S6752 }),
  .Y({ S6753 })
);
NAND #() 
NAND_3983_ (
  .A({ S6645 }),
  .B({ S6751 }),
  .Y({ S6754 })
);
NOR #() 
NOR_2377_ (
  .A({ S6645 }),
  .B({ S6751 }),
  .Y({ S6755 })
);
NAND #() 
NAND_3984_ (
  .A({ S6646 }),
  .B({ S6752 }),
  .Y({ S6756 })
);
NOR #() 
NOR_2378_ (
  .A({ S6753 }),
  .B({ S6755 }),
  .Y({ S6757 })
);
NAND #() 
NAND_3985_ (
  .A({ S6754 }),
  .B({ S6756 }),
  .Y({ S6758 })
);
NOR #() 
NOR_2379_ (
  .A({ S6625 }),
  .B({ S6758 }),
  .Y({ S6759 })
);
NAND #() 
NAND_3986_ (
  .A({ S6626 }),
  .B({ S6757 }),
  .Y({ S6760 })
);
NOR #() 
NOR_2380_ (
  .A({ S6626 }),
  .B({ S6757 }),
  .Y({ S6761 })
);
NOR #() 
NOR_2381_ (
  .A({ S6759 }),
  .B({ S6761 }),
  .Y({ S6762 })
);
NOT #() 
NOT_514_ (
  .A({ S6762 }),
  .Y({ S6763 })
);
NOR #() 
NOR_2382_ (
  .A({ S6486 }),
  .B({ S6763 }),
  .Y({ S6764 })
);
NOT #() 
NOT_515_ (
  .A({ S6764 }),
  .Y({ S6765 })
);
NOR #() 
NOR_2383_ (
  .A({ S6485 }),
  .B({ S6762 }),
  .Y({ S6766 })
);
NOR #() 
NOR_2384_ (
  .A({ S6764 }),
  .B({ S6766 }),
  .Y({ S6767 })
);
NAND #() 
NAND_3987_ (
  .A({ S6603 }),
  .B({ S6767 }),
  .Y({ S6768 })
);
NOT #() 
NOT_516_ (
  .A({ S6768 }),
  .Y({ S6769 })
);
NOR #() 
NOR_2385_ (
  .A({ S6603 }),
  .B({ S6767 }),
  .Y({ S6770 })
);
NOT #() 
NOT_517_ (
  .A({ S6770 }),
  .Y({ S6771 })
);
NOR #() 
NOR_2386_ (
  .A({ S6769 }),
  .B({ S6770 }),
  .Y({ S6772 })
);
NAND #() 
NAND_3988_ (
  .A({ S6768 }),
  .B({ S6771 }),
  .Y({ S6773 })
);
NOR #() 
NOR_2387_ (
  .A({ S6608 }),
  .B({ S6773 }),
  .Y({ S6774 })
);
NOR #() 
NOR_2388_ (
  .A({ S6607 }),
  .B({ S6772 }),
  .Y({ S6775 })
);
NOR #() 
NOR_2389_ (
  .A({ S6774 }),
  .B({ S6775 }),
  .Y({ S6776 })
);
NAND #() 
NAND_3989_ (
  .A({ S6624 }),
  .B({ S6776 }),
  .Y({ S6777 })
);
NOT #() 
NOT_518_ (
  .A({ S6777 }),
  .Y({ S6778 })
);
NOR #() 
NOR_2390_ (
  .A({ S6624 }),
  .B({ S6776 }),
  .Y({ S6779 })
);
NAND #() 
NAND_3990_ (
  .A({ S5948 }),
  .B({ S6777 }),
  .Y({ S6780 })
);
NOR #() 
NOR_2391_ (
  .A({ S6779 }),
  .B({ S6780 }),
  .Y({ S6781 })
);
NOR #() 
NOR_2392_ (
  .A({ S6622 }),
  .B({ S6781 }),
  .Y({ S6782 })
);
NAND #() 
NAND_3991_ (
  .A({ S6623 }),
  .B({ S6782 }),
  .Y({ S292 })
);
NOR #() 
NOR_2393_ (
  .A({ S3899 }),
  .B({ S4108 }),
  .Y({ S6783 })
);
NAND #() 
NAND_3992_ (
  .A({ datapath_multdivunit_outmdu1_11 }),
  .B({ S5950 }),
  .Y({ S6784 })
);
NOR #() 
NOR_2394_ (
  .A({ S6774 }),
  .B({ S6778 }),
  .Y({ S6785 })
);
NOR #() 
NOR_2395_ (
  .A({ S6759 }),
  .B({ S6764 }),
  .Y({ S6786 })
);
NAND #() 
NAND_3993_ (
  .A({ S6760 }),
  .B({ S6765 }),
  .Y({ S6787 })
);
NOR #() 
NOR_2396_ (
  .A({ S6747 }),
  .B({ S6753 }),
  .Y({ S6788 })
);
NAND #() 
NAND_3994_ (
  .A({ S6748 }),
  .B({ S6754 }),
  .Y({ S6789 })
);
NOR #() 
NOR_2397_ (
  .A({ S1220 }),
  .B({ S2718 }),
  .Y({ S6790 })
);
NAND #() 
NAND_3995_ (
  .A({ datapath_addsubunit_in1_0 }),
  .B({ S2717 }),
  .Y({ S6791 })
);
NOR #() 
NOR_2398_ (
  .A({ S1116 }),
  .B({ S2518 }),
  .Y({ S6792 })
);
NAND #() 
NAND_3996_ (
  .A({ datapath_addsubunit_in1_2 }),
  .B({ S2517 }),
  .Y({ S6793 })
);
NOR #() 
NOR_2399_ (
  .A({ S6633 }),
  .B({ S6792 }),
  .Y({ S6794 })
);
NAND #() 
NAND_3997_ (
  .A({ S6634 }),
  .B({ S6793 }),
  .Y({ S6795 })
);
NOR #() 
NOR_2400_ (
  .A({ S1116 }),
  .B({ S2618 }),
  .Y({ S6796 })
);
NAND #() 
NAND_3998_ (
  .A({ datapath_addsubunit_in1_2 }),
  .B({ S2617 }),
  .Y({ S6797 })
);
NOR #() 
NOR_2401_ (
  .A({ S6634 }),
  .B({ S6793 }),
  .Y({ S6798 })
);
NAND #() 
NAND_3999_ (
  .A({ S6633 }),
  .B({ S6792 }),
  .Y({ S6799 })
);
NOR #() 
NOR_2402_ (
  .A({ S6794 }),
  .B({ S6798 }),
  .Y({ S6800 })
);
NAND #() 
NAND_4000_ (
  .A({ S6795 }),
  .B({ S6799 }),
  .Y({ S6801 })
);
NOR #() 
NOR_2403_ (
  .A({ S6791 }),
  .B({ S6801 }),
  .Y({ S6802 })
);
NAND #() 
NAND_4001_ (
  .A({ S6790 }),
  .B({ S6800 }),
  .Y({ S6803 })
);
NOR #() 
NOR_2404_ (
  .A({ S6790 }),
  .B({ S6800 }),
  .Y({ S6804 })
);
NAND #() 
NAND_4002_ (
  .A({ S6791 }),
  .B({ S6801 }),
  .Y({ S6805 })
);
NOR #() 
NOR_2405_ (
  .A({ S6802 }),
  .B({ S6804 }),
  .Y({ S6806 })
);
NAND #() 
NAND_4003_ (
  .A({ S6803 }),
  .B({ S6805 }),
  .Y({ S6807 })
);
NOR #() 
NOR_2406_ (
  .A({ S6636 }),
  .B({ S6807 }),
  .Y({ S6808 })
);
NAND #() 
NAND_4004_ (
  .A({ S6635 }),
  .B({ S6806 }),
  .Y({ S6809 })
);
NOR #() 
NOR_2407_ (
  .A({ S6635 }),
  .B({ S6806 }),
  .Y({ S6810 })
);
NAND #() 
NAND_4005_ (
  .A({ S6636 }),
  .B({ S6807 }),
  .Y({ S6811 })
);
NOR #() 
NOR_2408_ (
  .A({ S6808 }),
  .B({ S6810 }),
  .Y({ S6812 })
);
NAND #() 
NAND_4006_ (
  .A({ S6809 }),
  .B({ S6811 }),
  .Y({ S6813 })
);
NOR #() 
NOR_2409_ (
  .A({ S6671 }),
  .B({ S6679 }),
  .Y({ S6814 })
);
NAND #() 
NAND_4007_ (
  .A({ S6672 }),
  .B({ S6680 }),
  .Y({ S6815 })
);
NOR #() 
NOR_2410_ (
  .A({ S6812 }),
  .B({ S6815 }),
  .Y({ S6816 })
);
NAND #() 
NAND_4008_ (
  .A({ S6813 }),
  .B({ S6814 }),
  .Y({ S6817 })
);
NOR #() 
NOR_2411_ (
  .A({ S6813 }),
  .B({ S6814 }),
  .Y({ S6818 })
);
NAND #() 
NAND_4009_ (
  .A({ S6812 }),
  .B({ S6815 }),
  .Y({ S6819 })
);
NOR #() 
NOR_2412_ (
  .A({ S6816 }),
  .B({ S6818 }),
  .Y({ S6820 })
);
NAND #() 
NAND_4010_ (
  .A({ S6817 }),
  .B({ S6819 }),
  .Y({ S6821 })
);
NOR #() 
NOR_2413_ (
  .A({ S6735 }),
  .B({ S6741 }),
  .Y({ S6822 })
);
NAND #() 
NAND_4011_ (
  .A({ S6736 }),
  .B({ S6742 }),
  .Y({ S6823 })
);
NOR #() 
NOR_2414_ (
  .A({ S6659 }),
  .B({ S6663 }),
  .Y({ S6824 })
);
NAND #() 
NAND_4012_ (
  .A({ S6660 }),
  .B({ S6664 }),
  .Y({ S6825 })
);
NOR #() 
NOR_2415_ (
  .A({ S1065 }),
  .B({ S2418 }),
  .Y({ S6826 })
);
NAND #() 
NAND_4013_ (
  .A({ datapath_addsubunit_in1_3 }),
  .B({ S2417 }),
  .Y({ S6827 })
);
NOR #() 
NOR_2416_ (
  .A({ S963 }),
  .B({ S2206 }),
  .Y({ S6828 })
);
NAND #() 
NAND_4014_ (
  .A({ datapath_addsubunit_in1_5 }),
  .B({ S2205 }),
  .Y({ S6829 })
);
NOR #() 
NOR_2417_ (
  .A({ S6657 }),
  .B({ S6828 }),
  .Y({ S6830 })
);
NAND #() 
NAND_4015_ (
  .A({ S6658 }),
  .B({ S6829 }),
  .Y({ S6831 })
);
NOR #() 
NOR_2418_ (
  .A({ S963 }),
  .B({ S2312 }),
  .Y({ S6832 })
);
NAND #() 
NAND_4016_ (
  .A({ datapath_addsubunit_in1_5 }),
  .B({ S2311 }),
  .Y({ S6833 })
);
NOR #() 
NOR_2419_ (
  .A({ S6658 }),
  .B({ S6829 }),
  .Y({ S6834 })
);
NAND #() 
NAND_4017_ (
  .A({ S6657 }),
  .B({ S6828 }),
  .Y({ S6835 })
);
NOR #() 
NOR_2420_ (
  .A({ S6830 }),
  .B({ S6834 }),
  .Y({ S6836 })
);
NAND #() 
NAND_4018_ (
  .A({ S6831 }),
  .B({ S6835 }),
  .Y({ S6837 })
);
NOR #() 
NOR_2421_ (
  .A({ S6827 }),
  .B({ S6837 }),
  .Y({ S6838 })
);
NAND #() 
NAND_4019_ (
  .A({ S6826 }),
  .B({ S6836 }),
  .Y({ S6839 })
);
NOR #() 
NOR_2422_ (
  .A({ S6826 }),
  .B({ S6836 }),
  .Y({ S6840 })
);
NAND #() 
NAND_4020_ (
  .A({ S6827 }),
  .B({ S6837 }),
  .Y({ S6841 })
);
NOR #() 
NOR_2423_ (
  .A({ S6838 }),
  .B({ S6840 }),
  .Y({ S6842 })
);
NAND #() 
NAND_4021_ (
  .A({ S6839 }),
  .B({ S6841 }),
  .Y({ S6843 })
);
NOR #() 
NOR_2424_ (
  .A({ S6693 }),
  .B({ S6697 }),
  .Y({ S6844 })
);
NAND #() 
NAND_4022_ (
  .A({ S6694 }),
  .B({ S6698 }),
  .Y({ S6845 })
);
NOR #() 
NOR_2425_ (
  .A({ S6843 }),
  .B({ S6844 }),
  .Y({ S6846 })
);
NAND #() 
NAND_4023_ (
  .A({ S6842 }),
  .B({ S6845 }),
  .Y({ S6847 })
);
NOR #() 
NOR_2426_ (
  .A({ S6842 }),
  .B({ S6845 }),
  .Y({ S6848 })
);
NAND #() 
NAND_4024_ (
  .A({ S6843 }),
  .B({ S6844 }),
  .Y({ S6849 })
);
NOR #() 
NOR_2427_ (
  .A({ S6846 }),
  .B({ S6848 }),
  .Y({ S6850 })
);
NAND #() 
NAND_4025_ (
  .A({ S6847 }),
  .B({ S6849 }),
  .Y({ S6851 })
);
NOR #() 
NOR_2428_ (
  .A({ S6825 }),
  .B({ S6850 }),
  .Y({ S6852 })
);
NAND #() 
NAND_4026_ (
  .A({ S6824 }),
  .B({ S6851 }),
  .Y({ S6853 })
);
NOR #() 
NOR_2429_ (
  .A({ S6824 }),
  .B({ S6851 }),
  .Y({ S6854 })
);
NAND #() 
NAND_4027_ (
  .A({ S6825 }),
  .B({ S6850 }),
  .Y({ S6855 })
);
NOR #() 
NOR_2430_ (
  .A({ S6852 }),
  .B({ S6854 }),
  .Y({ S6856 })
);
NAND #() 
NAND_4028_ (
  .A({ S6853 }),
  .B({ S6855 }),
  .Y({ S6857 })
);
NOR #() 
NOR_2431_ (
  .A({ S6723 }),
  .B({ S6729 }),
  .Y({ S6858 })
);
NAND #() 
NAND_4029_ (
  .A({ S6724 }),
  .B({ S6730 }),
  .Y({ S6859 })
);
NOR #() 
NOR_2432_ (
  .A({ S910 }),
  .B({ S2107 }),
  .Y({ S6860 })
);
NAND #() 
NAND_4030_ (
  .A({ datapath_addsubunit_in1_6 }),
  .B({ S2106 }),
  .Y({ S6861 })
);
NOR #() 
NOR_2433_ (
  .A({ S805 }),
  .B({ S1953 }),
  .Y({ S6862 })
);
NAND #() 
NAND_4031_ (
  .A({ datapath_addsubunit_in1_8 }),
  .B({ S1952 }),
  .Y({ S6863 })
);
NOR #() 
NOR_2434_ (
  .A({ S6691 }),
  .B({ S6862 }),
  .Y({ S6864 })
);
NAND #() 
NAND_4032_ (
  .A({ S6692 }),
  .B({ S6863 }),
  .Y({ S6865 })
);
NOR #() 
NOR_2435_ (
  .A({ S805 }),
  .B({ S1598 }),
  .Y({ S6866 })
);
NAND #() 
NAND_4033_ (
  .A({ datapath_addsubunit_in1_8 }),
  .B({ S1597 }),
  .Y({ S6867 })
);
NOR #() 
NOR_2436_ (
  .A({ S6692 }),
  .B({ S6863 }),
  .Y({ S6868 })
);
NAND #() 
NAND_4034_ (
  .A({ S6691 }),
  .B({ S6862 }),
  .Y({ S6869 })
);
NOR #() 
NOR_2437_ (
  .A({ S6864 }),
  .B({ S6868 }),
  .Y({ S6870 })
);
NAND #() 
NAND_4035_ (
  .A({ S6865 }),
  .B({ S6869 }),
  .Y({ S6871 })
);
NOR #() 
NOR_2438_ (
  .A({ S6861 }),
  .B({ S6871 }),
  .Y({ S6872 })
);
NAND #() 
NAND_4036_ (
  .A({ S6860 }),
  .B({ S6870 }),
  .Y({ S6873 })
);
NOR #() 
NOR_2439_ (
  .A({ S6860 }),
  .B({ S6870 }),
  .Y({ S6874 })
);
NAND #() 
NAND_4037_ (
  .A({ S6861 }),
  .B({ S6871 }),
  .Y({ S6875 })
);
NOR #() 
NOR_2440_ (
  .A({ S6872 }),
  .B({ S6874 }),
  .Y({ S6876 })
);
NAND #() 
NAND_4038_ (
  .A({ S6873 }),
  .B({ S6875 }),
  .Y({ S6877 })
);
NOR #() 
NOR_2441_ (
  .A({ S6713 }),
  .B({ S6717 }),
  .Y({ S6878 })
);
NAND #() 
NAND_4039_ (
  .A({ S6714 }),
  .B({ S6718 }),
  .Y({ S6879 })
);
NOR #() 
NOR_2442_ (
  .A({ S754 }),
  .B({ S1849 }),
  .Y({ S6880 })
);
NAND #() 
NAND_4040_ (
  .A({ datapath_addsubunit_in1_9 }),
  .B({ S1848 }),
  .Y({ S6881 })
);
NOR #() 
NOR_2443_ (
  .A({ S651 }),
  .B({ S1516 }),
  .Y({ S6882 })
);
NAND #() 
NAND_4041_ (
  .A({ datapath_addsubunit_in1_11 }),
  .B({ S1515 }),
  .Y({ S6883 })
);
NOR #() 
NOR_2444_ (
  .A({ S6711 }),
  .B({ S6882 }),
  .Y({ S6884 })
);
NAND #() 
NAND_4042_ (
  .A({ S6712 }),
  .B({ S6883 }),
  .Y({ S6885 })
);
NOR #() 
NOR_2445_ (
  .A({ S651 }),
  .B({ S1746 }),
  .Y({ S6886 })
);
NAND #() 
NAND_4043_ (
  .A({ datapath_addsubunit_in1_11 }),
  .B({ S1745 }),
  .Y({ S6887 })
);
NOR #() 
NOR_2446_ (
  .A({ S6712 }),
  .B({ S6883 }),
  .Y({ S6888 })
);
NAND #() 
NAND_4044_ (
  .A({ S6711 }),
  .B({ S6882 }),
  .Y({ S6889 })
);
NOR #() 
NOR_2447_ (
  .A({ S6884 }),
  .B({ S6888 }),
  .Y({ S6890 })
);
NAND #() 
NAND_4045_ (
  .A({ S6885 }),
  .B({ S6889 }),
  .Y({ S6891 })
);
NOR #() 
NOR_2448_ (
  .A({ S6881 }),
  .B({ S6891 }),
  .Y({ S6892 })
);
NAND #() 
NAND_4046_ (
  .A({ S6880 }),
  .B({ S6890 }),
  .Y({ S6893 })
);
NOR #() 
NOR_2449_ (
  .A({ S6880 }),
  .B({ S6890 }),
  .Y({ S6894 })
);
NAND #() 
NAND_4047_ (
  .A({ S6881 }),
  .B({ S6891 }),
  .Y({ S6895 })
);
NOR #() 
NOR_2450_ (
  .A({ S6892 }),
  .B({ S6894 }),
  .Y({ S6896 })
);
NAND #() 
NAND_4048_ (
  .A({ S6893 }),
  .B({ S6895 }),
  .Y({ S6897 })
);
NOR #() 
NOR_2451_ (
  .A({ S6878 }),
  .B({ S6897 }),
  .Y({ S6898 })
);
NAND #() 
NAND_4049_ (
  .A({ S6879 }),
  .B({ S6896 }),
  .Y({ S6899 })
);
NOR #() 
NOR_2452_ (
  .A({ S6879 }),
  .B({ S6896 }),
  .Y({ S6900 })
);
NAND #() 
NAND_4050_ (
  .A({ S6878 }),
  .B({ S6897 }),
  .Y({ S6901 })
);
NOR #() 
NOR_2453_ (
  .A({ S6898 }),
  .B({ S6900 }),
  .Y({ S6902 })
);
NAND #() 
NAND_4051_ (
  .A({ S6899 }),
  .B({ S6901 }),
  .Y({ S6903 })
);
NOR #() 
NOR_2454_ (
  .A({ S6877 }),
  .B({ S6903 }),
  .Y({ S6904 })
);
NAND #() 
NAND_4052_ (
  .A({ S6876 }),
  .B({ S6902 }),
  .Y({ S6905 })
);
NOR #() 
NOR_2455_ (
  .A({ S6876 }),
  .B({ S6902 }),
  .Y({ S6906 })
);
NAND #() 
NAND_4053_ (
  .A({ S6877 }),
  .B({ S6903 }),
  .Y({ S6907 })
);
NOR #() 
NOR_2456_ (
  .A({ S6904 }),
  .B({ S6906 }),
  .Y({ S6908 })
);
NAND #() 
NAND_4054_ (
  .A({ S6905 }),
  .B({ S6907 }),
  .Y({ S6909 })
);
NOR #() 
NOR_2457_ (
  .A({ S6858 }),
  .B({ S6909 }),
  .Y({ S6910 })
);
NAND #() 
NAND_4055_ (
  .A({ S6859 }),
  .B({ S6908 }),
  .Y({ S6911 })
);
NOR #() 
NOR_2458_ (
  .A({ S6859 }),
  .B({ S6908 }),
  .Y({ S6912 })
);
NAND #() 
NAND_4056_ (
  .A({ S6858 }),
  .B({ S6909 }),
  .Y({ S6913 })
);
NOR #() 
NOR_2459_ (
  .A({ S6910 }),
  .B({ S6912 }),
  .Y({ S6914 })
);
NAND #() 
NAND_4057_ (
  .A({ S6911 }),
  .B({ S6913 }),
  .Y({ S6915 })
);
NOR #() 
NOR_2460_ (
  .A({ S6857 }),
  .B({ S6915 }),
  .Y({ S6916 })
);
NAND #() 
NAND_4058_ (
  .A({ S6856 }),
  .B({ S6914 }),
  .Y({ S6917 })
);
NOR #() 
NOR_2461_ (
  .A({ S6856 }),
  .B({ S6914 }),
  .Y({ S6918 })
);
NAND #() 
NAND_4059_ (
  .A({ S6857 }),
  .B({ S6915 }),
  .Y({ S6919 })
);
NOR #() 
NOR_2462_ (
  .A({ S6916 }),
  .B({ S6918 }),
  .Y({ S6920 })
);
NAND #() 
NAND_4060_ (
  .A({ S6917 }),
  .B({ S6919 }),
  .Y({ S6921 })
);
NOR #() 
NOR_2463_ (
  .A({ S6822 }),
  .B({ S6921 }),
  .Y({ S6922 })
);
NAND #() 
NAND_4061_ (
  .A({ S6823 }),
  .B({ S6920 }),
  .Y({ S6923 })
);
NOR #() 
NOR_2464_ (
  .A({ S6823 }),
  .B({ S6920 }),
  .Y({ S6924 })
);
NAND #() 
NAND_4062_ (
  .A({ S6822 }),
  .B({ S6921 }),
  .Y({ S6925 })
);
NOR #() 
NOR_2465_ (
  .A({ S6922 }),
  .B({ S6924 }),
  .Y({ S6926 })
);
NAND #() 
NAND_4063_ (
  .A({ S6923 }),
  .B({ S6925 }),
  .Y({ S6927 })
);
NOR #() 
NOR_2466_ (
  .A({ S6821 }),
  .B({ S6927 }),
  .Y({ S6928 })
);
NAND #() 
NAND_4064_ (
  .A({ S6820 }),
  .B({ S6926 }),
  .Y({ S6929 })
);
NOR #() 
NOR_2467_ (
  .A({ S6820 }),
  .B({ S6926 }),
  .Y({ S6930 })
);
NAND #() 
NAND_4065_ (
  .A({ S6821 }),
  .B({ S6927 }),
  .Y({ S6931 })
);
NOR #() 
NOR_2468_ (
  .A({ S6928 }),
  .B({ S6930 }),
  .Y({ S6932 })
);
NAND #() 
NAND_4066_ (
  .A({ S6929 }),
  .B({ S6931 }),
  .Y({ S6933 })
);
NOR #() 
NOR_2469_ (
  .A({ S6788 }),
  .B({ S6933 }),
  .Y({ S6934 })
);
NAND #() 
NAND_4067_ (
  .A({ S6789 }),
  .B({ S6932 }),
  .Y({ S6935 })
);
NOR #() 
NOR_2470_ (
  .A({ S6789 }),
  .B({ S6932 }),
  .Y({ S6936 })
);
NAND #() 
NAND_4068_ (
  .A({ S6788 }),
  .B({ S6933 }),
  .Y({ S6937 })
);
NOR #() 
NOR_2471_ (
  .A({ S6934 }),
  .B({ S6936 }),
  .Y({ S6938 })
);
NAND #() 
NAND_4069_ (
  .A({ S6935 }),
  .B({ S6937 }),
  .Y({ S6939 })
);
NOR #() 
NOR_2472_ (
  .A({ S6644 }),
  .B({ S6939 }),
  .Y({ S6940 })
);
NAND #() 
NAND_4070_ (
  .A({ S6643 }),
  .B({ S6938 }),
  .Y({ S6941 })
);
NOR #() 
NOR_2473_ (
  .A({ S6643 }),
  .B({ S6938 }),
  .Y({ S6942 })
);
NAND #() 
NAND_4071_ (
  .A({ S6644 }),
  .B({ S6939 }),
  .Y({ S6943 })
);
NOR #() 
NOR_2474_ (
  .A({ S6940 }),
  .B({ S6942 }),
  .Y({ S6944 })
);
NAND #() 
NAND_4072_ (
  .A({ S6941 }),
  .B({ S6943 }),
  .Y({ S6945 })
);
NAND #() 
NAND_4073_ (
  .A({ S6786 }),
  .B({ S6945 }),
  .Y({ S6946 })
);
NAND #() 
NAND_4074_ (
  .A({ S6787 }),
  .B({ S6944 }),
  .Y({ S6947 })
);
NAND #() 
NAND_4075_ (
  .A({ S6946 }),
  .B({ S6947 }),
  .Y({ S6948 })
);
NOR #() 
NOR_2475_ (
  .A({ S6768 }),
  .B({ S6948 }),
  .Y({ S6949 })
);
NOT #() 
NOT_519_ (
  .A({ S6949 }),
  .Y({ S6950 })
);
NAND #() 
NAND_4076_ (
  .A({ S6768 }),
  .B({ S6948 }),
  .Y({ S6951 })
);
NAND #() 
NAND_4077_ (
  .A({ S6950 }),
  .B({ S6951 }),
  .Y({ S6952 })
);
NOR #() 
NOR_2476_ (
  .A({ S6785 }),
  .B({ S6952 }),
  .Y({ S6953 })
);
NAND #() 
NAND_4078_ (
  .A({ S6785 }),
  .B({ S6952 }),
  .Y({ S6954 })
);
NAND #() 
NAND_4079_ (
  .A({ S5948 }),
  .B({ S6954 }),
  .Y({ S6955 })
);
NOR #() 
NOR_2477_ (
  .A({ S6953 }),
  .B({ S6955 }),
  .Y({ S6956 })
);
NOR #() 
NOR_2478_ (
  .A({ S6783 }),
  .B({ S6956 }),
  .Y({ S6957 })
);
NAND #() 
NAND_4080_ (
  .A({ S6784 }),
  .B({ S6957 }),
  .Y({ S293 })
);
NOR #() 
NOR_2479_ (
  .A({ S3899 }),
  .B({ S4035 }),
  .Y({ S6958 })
);
NAND #() 
NAND_4081_ (
  .A({ datapath_multdivunit_outmdu1_12 }),
  .B({ S5950 }),
  .Y({ S6959 })
);
NOR #() 
NOR_2480_ (
  .A({ S6949 }),
  .B({ S6953 }),
  .Y({ S6960 })
);
NOR #() 
NOR_2481_ (
  .A({ S6934 }),
  .B({ S6940 }),
  .Y({ S6961 })
);
NAND #() 
NAND_4082_ (
  .A({ S6935 }),
  .B({ S6941 }),
  .Y({ S6962 })
);
NOR #() 
NOR_2482_ (
  .A({ S6922 }),
  .B({ S6928 }),
  .Y({ S6963 })
);
NAND #() 
NAND_4083_ (
  .A({ S6923 }),
  .B({ S6929 }),
  .Y({ S6964 })
);
NOR #() 
NOR_2483_ (
  .A({ S1220 }),
  .B({ S2817 }),
  .Y({ S6965 })
);
NAND #() 
NAND_4084_ (
  .A({ datapath_addsubunit_in1_0 }),
  .B({ S2816 }),
  .Y({ S6966 })
);
NOR #() 
NOR_2484_ (
  .A({ S6798 }),
  .B({ S6802 }),
  .Y({ S6967 })
);
NAND #() 
NAND_4085_ (
  .A({ S6799 }),
  .B({ S6803 }),
  .Y({ S6968 })
);
NOR #() 
NOR_2485_ (
  .A({ S1168 }),
  .B({ S2718 }),
  .Y({ S6969 })
);
NAND #() 
NAND_4086_ (
  .A({ datapath_addsubunit_in1_1 }),
  .B({ S2717 }),
  .Y({ S6970 })
);
NOR #() 
NOR_2486_ (
  .A({ S1065 }),
  .B({ S2518 }),
  .Y({ S6971 })
);
NAND #() 
NAND_4087_ (
  .A({ datapath_addsubunit_in1_3 }),
  .B({ S2517 }),
  .Y({ S6972 })
);
NOR #() 
NOR_2487_ (
  .A({ S6796 }),
  .B({ S6971 }),
  .Y({ S6973 })
);
NAND #() 
NAND_4088_ (
  .A({ S6797 }),
  .B({ S6972 }),
  .Y({ S6974 })
);
NOR #() 
NOR_2488_ (
  .A({ S1065 }),
  .B({ S2618 }),
  .Y({ S6975 })
);
NAND #() 
NAND_4089_ (
  .A({ datapath_addsubunit_in1_3 }),
  .B({ S2617 }),
  .Y({ S6976 })
);
NOR #() 
NOR_2489_ (
  .A({ S6797 }),
  .B({ S6972 }),
  .Y({ S6977 })
);
NAND #() 
NAND_4090_ (
  .A({ S6796 }),
  .B({ S6971 }),
  .Y({ S6978 })
);
NOR #() 
NOR_2490_ (
  .A({ S6973 }),
  .B({ S6977 }),
  .Y({ S6979 })
);
NAND #() 
NAND_4091_ (
  .A({ S6974 }),
  .B({ S6978 }),
  .Y({ S6980 })
);
NOR #() 
NOR_2491_ (
  .A({ S6970 }),
  .B({ S6980 }),
  .Y({ S6981 })
);
NAND #() 
NAND_4092_ (
  .A({ S6969 }),
  .B({ S6979 }),
  .Y({ S6982 })
);
NOR #() 
NOR_2492_ (
  .A({ S6969 }),
  .B({ S6979 }),
  .Y({ S6983 })
);
NAND #() 
NAND_4093_ (
  .A({ S6970 }),
  .B({ S6980 }),
  .Y({ S6984 })
);
NOR #() 
NOR_2493_ (
  .A({ S6981 }),
  .B({ S6983 }),
  .Y({ S6985 })
);
NAND #() 
NAND_4094_ (
  .A({ S6982 }),
  .B({ S6984 }),
  .Y({ S6986 })
);
NOR #() 
NOR_2494_ (
  .A({ S6967 }),
  .B({ S6986 }),
  .Y({ S6987 })
);
NAND #() 
NAND_4095_ (
  .A({ S6968 }),
  .B({ S6985 }),
  .Y({ S6988 })
);
NOR #() 
NOR_2495_ (
  .A({ S6968 }),
  .B({ S6985 }),
  .Y({ S6989 })
);
NAND #() 
NAND_4096_ (
  .A({ S6967 }),
  .B({ S6986 }),
  .Y({ S6990 })
);
NOR #() 
NOR_2496_ (
  .A({ S6987 }),
  .B({ S6989 }),
  .Y({ S6991 })
);
NAND #() 
NAND_4097_ (
  .A({ S6988 }),
  .B({ S6990 }),
  .Y({ S6992 })
);
NOR #() 
NOR_2497_ (
  .A({ S6966 }),
  .B({ S6992 }),
  .Y({ S6993 })
);
NAND #() 
NAND_4098_ (
  .A({ S6965 }),
  .B({ S6991 }),
  .Y({ S6994 })
);
NOR #() 
NOR_2498_ (
  .A({ S6965 }),
  .B({ S6991 }),
  .Y({ S6995 })
);
NAND #() 
NAND_4099_ (
  .A({ S6966 }),
  .B({ S6992 }),
  .Y({ S6996 })
);
NOR #() 
NOR_2499_ (
  .A({ S6993 }),
  .B({ S6995 }),
  .Y({ S6997 })
);
NAND #() 
NAND_4100_ (
  .A({ S6994 }),
  .B({ S6996 }),
  .Y({ S6998 })
);
NOR #() 
NOR_2500_ (
  .A({ S6846 }),
  .B({ S6854 }),
  .Y({ S6999 })
);
NAND #() 
NAND_4101_ (
  .A({ S6847 }),
  .B({ S6855 }),
  .Y({ S7000 })
);
NOR #() 
NOR_2501_ (
  .A({ S6998 }),
  .B({ S6999 }),
  .Y({ S7001 })
);
NAND #() 
NAND_4102_ (
  .A({ S6997 }),
  .B({ S7000 }),
  .Y({ S7002 })
);
NOR #() 
NOR_2502_ (
  .A({ S6997 }),
  .B({ S7000 }),
  .Y({ S7003 })
);
NAND #() 
NAND_4103_ (
  .A({ S6998 }),
  .B({ S6999 }),
  .Y({ S7004 })
);
NOR #() 
NOR_2503_ (
  .A({ S7001 }),
  .B({ S7003 }),
  .Y({ S7005 })
);
NAND #() 
NAND_4104_ (
  .A({ S7002 }),
  .B({ S7004 }),
  .Y({ S7006 })
);
NOR #() 
NOR_2504_ (
  .A({ S6809 }),
  .B({ S7006 }),
  .Y({ S7007 })
);
NAND #() 
NAND_4105_ (
  .A({ S6808 }),
  .B({ S7005 }),
  .Y({ S7008 })
);
NOR #() 
NOR_2505_ (
  .A({ S6808 }),
  .B({ S7005 }),
  .Y({ S7009 })
);
NAND #() 
NAND_4106_ (
  .A({ S6809 }),
  .B({ S7006 }),
  .Y({ S7010 })
);
NOR #() 
NOR_2506_ (
  .A({ S7007 }),
  .B({ S7009 }),
  .Y({ S7011 })
);
NAND #() 
NAND_4107_ (
  .A({ S7008 }),
  .B({ S7010 }),
  .Y({ S7012 })
);
NOR #() 
NOR_2507_ (
  .A({ S6910 }),
  .B({ S6916 }),
  .Y({ S7013 })
);
NAND #() 
NAND_4108_ (
  .A({ S6911 }),
  .B({ S6917 }),
  .Y({ S7014 })
);
NOR #() 
NOR_2508_ (
  .A({ S6834 }),
  .B({ S6838 }),
  .Y({ S7015 })
);
NAND #() 
NAND_4109_ (
  .A({ S6835 }),
  .B({ S6839 }),
  .Y({ S7016 })
);
NOR #() 
NOR_2509_ (
  .A({ S1013 }),
  .B({ S2418 }),
  .Y({ S7017 })
);
NAND #() 
NAND_4110_ (
  .A({ datapath_addsubunit_in1_4 }),
  .B({ S2417 }),
  .Y({ S7018 })
);
NOR #() 
NOR_2510_ (
  .A({ S910 }),
  .B({ S2206 }),
  .Y({ S7019 })
);
NAND #() 
NAND_4111_ (
  .A({ datapath_addsubunit_in1_6 }),
  .B({ S2205 }),
  .Y({ S7020 })
);
NOR #() 
NOR_2511_ (
  .A({ S6832 }),
  .B({ S7019 }),
  .Y({ S7021 })
);
NAND #() 
NAND_4112_ (
  .A({ S6833 }),
  .B({ S7020 }),
  .Y({ S7022 })
);
NOR #() 
NOR_2512_ (
  .A({ S910 }),
  .B({ S2312 }),
  .Y({ S7023 })
);
NAND #() 
NAND_4113_ (
  .A({ datapath_addsubunit_in1_6 }),
  .B({ S2311 }),
  .Y({ S7024 })
);
NOR #() 
NOR_2513_ (
  .A({ S6833 }),
  .B({ S7020 }),
  .Y({ S7025 })
);
NAND #() 
NAND_4114_ (
  .A({ S6832 }),
  .B({ S7019 }),
  .Y({ S7026 })
);
NOR #() 
NOR_2514_ (
  .A({ S7021 }),
  .B({ S7025 }),
  .Y({ S7027 })
);
NAND #() 
NAND_4115_ (
  .A({ S7022 }),
  .B({ S7026 }),
  .Y({ S7028 })
);
NOR #() 
NOR_2515_ (
  .A({ S7018 }),
  .B({ S7028 }),
  .Y({ S7029 })
);
NAND #() 
NAND_4116_ (
  .A({ S7017 }),
  .B({ S7027 }),
  .Y({ S7030 })
);
NOR #() 
NOR_2516_ (
  .A({ S7017 }),
  .B({ S7027 }),
  .Y({ S7031 })
);
NAND #() 
NAND_4117_ (
  .A({ S7018 }),
  .B({ S7028 }),
  .Y({ S7032 })
);
NOR #() 
NOR_2517_ (
  .A({ S7029 }),
  .B({ S7031 }),
  .Y({ S7033 })
);
NAND #() 
NAND_4118_ (
  .A({ S7030 }),
  .B({ S7032 }),
  .Y({ S7034 })
);
NOR #() 
NOR_2518_ (
  .A({ S6868 }),
  .B({ S6872 }),
  .Y({ S7035 })
);
NAND #() 
NAND_4119_ (
  .A({ S6869 }),
  .B({ S6873 }),
  .Y({ S7036 })
);
NOR #() 
NOR_2519_ (
  .A({ S7034 }),
  .B({ S7035 }),
  .Y({ S7037 })
);
NAND #() 
NAND_4120_ (
  .A({ S7033 }),
  .B({ S7036 }),
  .Y({ S7038 })
);
NOR #() 
NOR_2520_ (
  .A({ S7033 }),
  .B({ S7036 }),
  .Y({ S7039 })
);
NAND #() 
NAND_4121_ (
  .A({ S7034 }),
  .B({ S7035 }),
  .Y({ S7040 })
);
NOR #() 
NOR_2521_ (
  .A({ S7037 }),
  .B({ S7039 }),
  .Y({ S7041 })
);
NAND #() 
NAND_4122_ (
  .A({ S7038 }),
  .B({ S7040 }),
  .Y({ S7042 })
);
NOR #() 
NOR_2522_ (
  .A({ S7016 }),
  .B({ S7041 }),
  .Y({ S7043 })
);
NAND #() 
NAND_4123_ (
  .A({ S7015 }),
  .B({ S7042 }),
  .Y({ S7044 })
);
NOR #() 
NOR_2523_ (
  .A({ S7015 }),
  .B({ S7042 }),
  .Y({ S7045 })
);
NAND #() 
NAND_4124_ (
  .A({ S7016 }),
  .B({ S7041 }),
  .Y({ S7046 })
);
NOR #() 
NOR_2524_ (
  .A({ S7043 }),
  .B({ S7045 }),
  .Y({ S7047 })
);
NAND #() 
NAND_4125_ (
  .A({ S7044 }),
  .B({ S7046 }),
  .Y({ S7048 })
);
NOR #() 
NOR_2525_ (
  .A({ S6898 }),
  .B({ S6904 }),
  .Y({ S7049 })
);
NAND #() 
NAND_4126_ (
  .A({ S6899 }),
  .B({ S6905 }),
  .Y({ S7050 })
);
NOR #() 
NOR_2526_ (
  .A({ S858 }),
  .B({ S2107 }),
  .Y({ S7051 })
);
NAND #() 
NAND_4127_ (
  .A({ datapath_addsubunit_in1_7 }),
  .B({ S2106 }),
  .Y({ S7052 })
);
NOR #() 
NOR_2527_ (
  .A({ S754 }),
  .B({ S1953 }),
  .Y({ S7053 })
);
NAND #() 
NAND_4128_ (
  .A({ datapath_addsubunit_in1_9 }),
  .B({ S1952 }),
  .Y({ S7054 })
);
NOR #() 
NOR_2528_ (
  .A({ S6866 }),
  .B({ S7053 }),
  .Y({ S7055 })
);
NAND #() 
NAND_4129_ (
  .A({ S6867 }),
  .B({ S7054 }),
  .Y({ S7056 })
);
NOR #() 
NOR_2529_ (
  .A({ S754 }),
  .B({ S1598 }),
  .Y({ S7057 })
);
NAND #() 
NAND_4130_ (
  .A({ datapath_addsubunit_in1_9 }),
  .B({ S1597 }),
  .Y({ S7058 })
);
NOR #() 
NOR_2530_ (
  .A({ S6867 }),
  .B({ S7054 }),
  .Y({ S7059 })
);
NAND #() 
NAND_4131_ (
  .A({ S6866 }),
  .B({ S7053 }),
  .Y({ S7060 })
);
NOR #() 
NOR_2531_ (
  .A({ S7055 }),
  .B({ S7059 }),
  .Y({ S7061 })
);
NAND #() 
NAND_4132_ (
  .A({ S7056 }),
  .B({ S7060 }),
  .Y({ S7062 })
);
NOR #() 
NOR_2532_ (
  .A({ S7052 }),
  .B({ S7062 }),
  .Y({ S7063 })
);
NAND #() 
NAND_4133_ (
  .A({ S7051 }),
  .B({ S7061 }),
  .Y({ S7064 })
);
NOR #() 
NOR_2533_ (
  .A({ S7051 }),
  .B({ S7061 }),
  .Y({ S7065 })
);
NAND #() 
NAND_4134_ (
  .A({ S7052 }),
  .B({ S7062 }),
  .Y({ S7066 })
);
NOR #() 
NOR_2534_ (
  .A({ S7063 }),
  .B({ S7065 }),
  .Y({ S7067 })
);
NAND #() 
NAND_4135_ (
  .A({ S7064 }),
  .B({ S7066 }),
  .Y({ S7068 })
);
NOR #() 
NOR_2535_ (
  .A({ S6888 }),
  .B({ S6892 }),
  .Y({ S7069 })
);
NAND #() 
NAND_4136_ (
  .A({ S6889 }),
  .B({ S6893 }),
  .Y({ S7070 })
);
NOR #() 
NOR_2536_ (
  .A({ S702 }),
  .B({ S1849 }),
  .Y({ S7071 })
);
NAND #() 
NAND_4137_ (
  .A({ datapath_addsubunit_in1_10 }),
  .B({ S1848 }),
  .Y({ S7072 })
);
NOR #() 
NOR_2537_ (
  .A({ S599 }),
  .B({ S1516 }),
  .Y({ S7073 })
);
NAND #() 
NAND_4138_ (
  .A({ datapath_addsubunit_in1_12 }),
  .B({ S1515 }),
  .Y({ S7074 })
);
NOR #() 
NOR_2538_ (
  .A({ S6886 }),
  .B({ S7073 }),
  .Y({ S7075 })
);
NAND #() 
NAND_4139_ (
  .A({ S6887 }),
  .B({ S7074 }),
  .Y({ S7076 })
);
NOR #() 
NOR_2539_ (
  .A({ S599 }),
  .B({ S1746 }),
  .Y({ S7077 })
);
NAND #() 
NAND_4140_ (
  .A({ datapath_addsubunit_in1_12 }),
  .B({ S1745 }),
  .Y({ S7078 })
);
NOR #() 
NOR_2540_ (
  .A({ S6887 }),
  .B({ S7074 }),
  .Y({ S7079 })
);
NAND #() 
NAND_4141_ (
  .A({ S6886 }),
  .B({ S7073 }),
  .Y({ S7080 })
);
NOR #() 
NOR_2541_ (
  .A({ S7075 }),
  .B({ S7079 }),
  .Y({ S7081 })
);
NAND #() 
NAND_4142_ (
  .A({ S7076 }),
  .B({ S7080 }),
  .Y({ S7082 })
);
NOR #() 
NOR_2542_ (
  .A({ S7072 }),
  .B({ S7082 }),
  .Y({ S7083 })
);
NAND #() 
NAND_4143_ (
  .A({ S7071 }),
  .B({ S7081 }),
  .Y({ S7084 })
);
NOR #() 
NOR_2543_ (
  .A({ S7071 }),
  .B({ S7081 }),
  .Y({ S7085 })
);
NAND #() 
NAND_4144_ (
  .A({ S7072 }),
  .B({ S7082 }),
  .Y({ S7086 })
);
NOR #() 
NOR_2544_ (
  .A({ S7083 }),
  .B({ S7085 }),
  .Y({ S7087 })
);
NAND #() 
NAND_4145_ (
  .A({ S7084 }),
  .B({ S7086 }),
  .Y({ S7088 })
);
NOR #() 
NOR_2545_ (
  .A({ S7069 }),
  .B({ S7088 }),
  .Y({ S7089 })
);
NAND #() 
NAND_4146_ (
  .A({ S7070 }),
  .B({ S7087 }),
  .Y({ S7090 })
);
NOR #() 
NOR_2546_ (
  .A({ S7070 }),
  .B({ S7087 }),
  .Y({ S7091 })
);
NAND #() 
NAND_4147_ (
  .A({ S7069 }),
  .B({ S7088 }),
  .Y({ S7092 })
);
NOR #() 
NOR_2547_ (
  .A({ S7089 }),
  .B({ S7091 }),
  .Y({ S7093 })
);
NAND #() 
NAND_4148_ (
  .A({ S7090 }),
  .B({ S7092 }),
  .Y({ S7094 })
);
NOR #() 
NOR_2548_ (
  .A({ S7068 }),
  .B({ S7094 }),
  .Y({ S7095 })
);
NAND #() 
NAND_4149_ (
  .A({ S7067 }),
  .B({ S7093 }),
  .Y({ S7096 })
);
NOR #() 
NOR_2549_ (
  .A({ S7067 }),
  .B({ S7093 }),
  .Y({ S7097 })
);
NAND #() 
NAND_4150_ (
  .A({ S7068 }),
  .B({ S7094 }),
  .Y({ S7098 })
);
NOR #() 
NOR_2550_ (
  .A({ S7095 }),
  .B({ S7097 }),
  .Y({ S7099 })
);
NAND #() 
NAND_4151_ (
  .A({ S7096 }),
  .B({ S7098 }),
  .Y({ S7100 })
);
NOR #() 
NOR_2551_ (
  .A({ S7049 }),
  .B({ S7100 }),
  .Y({ S7101 })
);
NAND #() 
NAND_4152_ (
  .A({ S7050 }),
  .B({ S7099 }),
  .Y({ S7102 })
);
NOR #() 
NOR_2552_ (
  .A({ S7050 }),
  .B({ S7099 }),
  .Y({ S7103 })
);
NAND #() 
NAND_4153_ (
  .A({ S7049 }),
  .B({ S7100 }),
  .Y({ S7104 })
);
NOR #() 
NOR_2553_ (
  .A({ S7101 }),
  .B({ S7103 }),
  .Y({ S7105 })
);
NAND #() 
NAND_4154_ (
  .A({ S7102 }),
  .B({ S7104 }),
  .Y({ S7106 })
);
NOR #() 
NOR_2554_ (
  .A({ S7048 }),
  .B({ S7106 }),
  .Y({ S7107 })
);
NAND #() 
NAND_4155_ (
  .A({ S7047 }),
  .B({ S7105 }),
  .Y({ S7108 })
);
NOR #() 
NOR_2555_ (
  .A({ S7047 }),
  .B({ S7105 }),
  .Y({ S7109 })
);
NAND #() 
NAND_4156_ (
  .A({ S7048 }),
  .B({ S7106 }),
  .Y({ S7110 })
);
NOR #() 
NOR_2556_ (
  .A({ S7107 }),
  .B({ S7109 }),
  .Y({ S7111 })
);
NAND #() 
NAND_4157_ (
  .A({ S7108 }),
  .B({ S7110 }),
  .Y({ S7112 })
);
NOR #() 
NOR_2557_ (
  .A({ S7013 }),
  .B({ S7112 }),
  .Y({ S7113 })
);
NAND #() 
NAND_4158_ (
  .A({ S7014 }),
  .B({ S7111 }),
  .Y({ S7114 })
);
NOR #() 
NOR_2558_ (
  .A({ S7014 }),
  .B({ S7111 }),
  .Y({ S7115 })
);
NAND #() 
NAND_4159_ (
  .A({ S7013 }),
  .B({ S7112 }),
  .Y({ S7116 })
);
NOR #() 
NOR_2559_ (
  .A({ S7113 }),
  .B({ S7115 }),
  .Y({ S7117 })
);
NAND #() 
NAND_4160_ (
  .A({ S7114 }),
  .B({ S7116 }),
  .Y({ S7118 })
);
NOR #() 
NOR_2560_ (
  .A({ S7012 }),
  .B({ S7118 }),
  .Y({ S7119 })
);
NAND #() 
NAND_4161_ (
  .A({ S7011 }),
  .B({ S7117 }),
  .Y({ S7120 })
);
NOR #() 
NOR_2561_ (
  .A({ S7011 }),
  .B({ S7117 }),
  .Y({ S7121 })
);
NAND #() 
NAND_4162_ (
  .A({ S7012 }),
  .B({ S7118 }),
  .Y({ S7122 })
);
NOR #() 
NOR_2562_ (
  .A({ S7119 }),
  .B({ S7121 }),
  .Y({ S7123 })
);
NAND #() 
NAND_4163_ (
  .A({ S7120 }),
  .B({ S7122 }),
  .Y({ S7124 })
);
NOR #() 
NOR_2563_ (
  .A({ S6963 }),
  .B({ S7124 }),
  .Y({ S7125 })
);
NAND #() 
NAND_4164_ (
  .A({ S6964 }),
  .B({ S7123 }),
  .Y({ S7126 })
);
NOR #() 
NOR_2564_ (
  .A({ S6964 }),
  .B({ S7123 }),
  .Y({ S7127 })
);
NAND #() 
NAND_4165_ (
  .A({ S6963 }),
  .B({ S7124 }),
  .Y({ S7128 })
);
NOR #() 
NOR_2565_ (
  .A({ S7125 }),
  .B({ S7127 }),
  .Y({ S7129 })
);
NAND #() 
NAND_4166_ (
  .A({ S7126 }),
  .B({ S7128 }),
  .Y({ S7130 })
);
NOR #() 
NOR_2566_ (
  .A({ S6819 }),
  .B({ S7130 }),
  .Y({ S7131 })
);
NAND #() 
NAND_4167_ (
  .A({ S6818 }),
  .B({ S7129 }),
  .Y({ S7132 })
);
NOR #() 
NOR_2567_ (
  .A({ S6818 }),
  .B({ S7129 }),
  .Y({ S7133 })
);
NAND #() 
NAND_4168_ (
  .A({ S6819 }),
  .B({ S7130 }),
  .Y({ S7134 })
);
NOR #() 
NOR_2568_ (
  .A({ S7131 }),
  .B({ S7133 }),
  .Y({ S7135 })
);
NAND #() 
NAND_4169_ (
  .A({ S7132 }),
  .B({ S7134 }),
  .Y({ S7136 })
);
NAND #() 
NAND_4170_ (
  .A({ S6961 }),
  .B({ S7136 }),
  .Y({ S7137 })
);
NAND #() 
NAND_4171_ (
  .A({ S6962 }),
  .B({ S7135 }),
  .Y({ S7138 })
);
NAND #() 
NAND_4172_ (
  .A({ S7137 }),
  .B({ S7138 }),
  .Y({ S7139 })
);
NOR #() 
NOR_2569_ (
  .A({ S6947 }),
  .B({ S7139 }),
  .Y({ S7140 })
);
NOT #() 
NOT_520_ (
  .A({ S7140 }),
  .Y({ S7141 })
);
NAND #() 
NAND_4173_ (
  .A({ S6947 }),
  .B({ S7139 }),
  .Y({ S7142 })
);
NAND #() 
NAND_4174_ (
  .A({ S7141 }),
  .B({ S7142 }),
  .Y({ S7143 })
);
NOR #() 
NOR_2570_ (
  .A({ S6960 }),
  .B({ S7143 }),
  .Y({ S7144 })
);
NAND #() 
NAND_4175_ (
  .A({ S6960 }),
  .B({ S7143 }),
  .Y({ S7145 })
);
NAND #() 
NAND_4176_ (
  .A({ S5948 }),
  .B({ S7145 }),
  .Y({ S7146 })
);
NOR #() 
NOR_2571_ (
  .A({ S7144 }),
  .B({ S7146 }),
  .Y({ S7147 })
);
NOR #() 
NOR_2572_ (
  .A({ S6958 }),
  .B({ S7147 }),
  .Y({ S7148 })
);
NAND #() 
NAND_4177_ (
  .A({ S6959 }),
  .B({ S7148 }),
  .Y({ S294 })
);
NOR #() 
NOR_2573_ (
  .A({ S7140 }),
  .B({ S7144 }),
  .Y({ S7149 })
);
NOR #() 
NOR_2574_ (
  .A({ S7125 }),
  .B({ S7131 }),
  .Y({ S7150 })
);
NAND #() 
NAND_4178_ (
  .A({ S7126 }),
  .B({ S7132 }),
  .Y({ S7151 })
);
NOR #() 
NOR_2575_ (
  .A({ S7001 }),
  .B({ S7007 }),
  .Y({ S7152 })
);
NAND #() 
NAND_4179_ (
  .A({ S7002 }),
  .B({ S7008 }),
  .Y({ S7153 })
);
NOR #() 
NOR_2576_ (
  .A({ S7113 }),
  .B({ S7119 }),
  .Y({ S7154 })
);
NAND #() 
NAND_4180_ (
  .A({ S7114 }),
  .B({ S7120 }),
  .Y({ S7155 })
);
NOR #() 
NOR_2577_ (
  .A({ S6987 }),
  .B({ S6993 }),
  .Y({ S7156 })
);
NAND #() 
NAND_4181_ (
  .A({ S6988 }),
  .B({ S6994 }),
  .Y({ S7157 })
);
NOR #() 
NOR_2578_ (
  .A({ S1220 }),
  .B({ S2920 }),
  .Y({ S7158 })
);
NOR #() 
NOR_2579_ (
  .A({ S1168 }),
  .B({ S2817 }),
  .Y({ S7159 })
);
NAND #() 
NAND_4182_ (
  .A({ datapath_addsubunit_in1_1 }),
  .B({ S2816 }),
  .Y({ S7160 })
);
NOR #() 
NOR_2580_ (
  .A({ S7158 }),
  .B({ S7159 }),
  .Y({ S7161 })
);
NOT #() 
NOT_521_ (
  .A({ S7161 }),
  .Y({ S7162 })
);
NOR #() 
NOR_2581_ (
  .A({ S1168 }),
  .B({ S2920 }),
  .Y({ S7163 })
);
NAND #() 
NAND_4183_ (
  .A({ datapath_addsubunit_in1_1 }),
  .B({ S2919 }),
  .Y({ S7164 })
);
NOR #() 
NOR_2582_ (
  .A({ S6966 }),
  .B({ S7164 }),
  .Y({ S7165 })
);
NAND #() 
NAND_4184_ (
  .A({ S6965 }),
  .B({ S7163 }),
  .Y({ S7166 })
);
NOR #() 
NOR_2583_ (
  .A({ S7161 }),
  .B({ S7165 }),
  .Y({ S7167 })
);
NAND #() 
NAND_4185_ (
  .A({ S7162 }),
  .B({ S7166 }),
  .Y({ S7168 })
);
NOR #() 
NOR_2584_ (
  .A({ S6977 }),
  .B({ S6981 }),
  .Y({ S7169 })
);
NAND #() 
NAND_4186_ (
  .A({ S6978 }),
  .B({ S6982 }),
  .Y({ S7170 })
);
NOR #() 
NOR_2585_ (
  .A({ S1116 }),
  .B({ S2718 }),
  .Y({ S7171 })
);
NAND #() 
NAND_4187_ (
  .A({ datapath_addsubunit_in1_2 }),
  .B({ S2717 }),
  .Y({ S7172 })
);
NOR #() 
NOR_2586_ (
  .A({ S1013 }),
  .B({ S2518 }),
  .Y({ S7173 })
);
NAND #() 
NAND_4188_ (
  .A({ datapath_addsubunit_in1_4 }),
  .B({ S2517 }),
  .Y({ S7174 })
);
NOR #() 
NOR_2587_ (
  .A({ S6975 }),
  .B({ S7173 }),
  .Y({ S7175 })
);
NAND #() 
NAND_4189_ (
  .A({ S6976 }),
  .B({ S7174 }),
  .Y({ S7176 })
);
NOR #() 
NOR_2588_ (
  .A({ S1013 }),
  .B({ S2618 }),
  .Y({ S7177 })
);
NAND #() 
NAND_4190_ (
  .A({ datapath_addsubunit_in1_4 }),
  .B({ S2617 }),
  .Y({ S7178 })
);
NOR #() 
NOR_2589_ (
  .A({ S6976 }),
  .B({ S7174 }),
  .Y({ S7179 })
);
NAND #() 
NAND_4191_ (
  .A({ S6975 }),
  .B({ S7173 }),
  .Y({ S7180 })
);
NOR #() 
NOR_2590_ (
  .A({ S7175 }),
  .B({ S7179 }),
  .Y({ S7181 })
);
NAND #() 
NAND_4192_ (
  .A({ S7176 }),
  .B({ S7180 }),
  .Y({ S7182 })
);
NOR #() 
NOR_2591_ (
  .A({ S7172 }),
  .B({ S7182 }),
  .Y({ S7183 })
);
NAND #() 
NAND_4193_ (
  .A({ S7171 }),
  .B({ S7181 }),
  .Y({ S7184 })
);
NOR #() 
NOR_2592_ (
  .A({ S7171 }),
  .B({ S7181 }),
  .Y({ S7185 })
);
NAND #() 
NAND_4194_ (
  .A({ S7172 }),
  .B({ S7182 }),
  .Y({ S7186 })
);
NOR #() 
NOR_2593_ (
  .A({ S7183 }),
  .B({ S7185 }),
  .Y({ S7187 })
);
NAND #() 
NAND_4195_ (
  .A({ S7184 }),
  .B({ S7186 }),
  .Y({ S7188 })
);
NOR #() 
NOR_2594_ (
  .A({ S7169 }),
  .B({ S7188 }),
  .Y({ S7189 })
);
NAND #() 
NAND_4196_ (
  .A({ S7170 }),
  .B({ S7187 }),
  .Y({ S7190 })
);
NOR #() 
NOR_2595_ (
  .A({ S7170 }),
  .B({ S7187 }),
  .Y({ S7191 })
);
NAND #() 
NAND_4197_ (
  .A({ S7169 }),
  .B({ S7188 }),
  .Y({ S7192 })
);
NOR #() 
NOR_2596_ (
  .A({ S7189 }),
  .B({ S7191 }),
  .Y({ S7193 })
);
NAND #() 
NAND_4198_ (
  .A({ S7190 }),
  .B({ S7192 }),
  .Y({ S7194 })
);
NOR #() 
NOR_2597_ (
  .A({ S7167 }),
  .B({ S7193 }),
  .Y({ S7195 })
);
NAND #() 
NAND_4199_ (
  .A({ S7168 }),
  .B({ S7194 }),
  .Y({ S7196 })
);
NOR #() 
NOR_2598_ (
  .A({ S7168 }),
  .B({ S7194 }),
  .Y({ S7197 })
);
NAND #() 
NAND_4200_ (
  .A({ S7167 }),
  .B({ S7193 }),
  .Y({ S7198 })
);
NOR #() 
NOR_2599_ (
  .A({ S7195 }),
  .B({ S7197 }),
  .Y({ S7199 })
);
NAND #() 
NAND_4201_ (
  .A({ S7196 }),
  .B({ S7198 }),
  .Y({ S7200 })
);
NOR #() 
NOR_2600_ (
  .A({ S7037 }),
  .B({ S7045 }),
  .Y({ S7201 })
);
NAND #() 
NAND_4202_ (
  .A({ S7038 }),
  .B({ S7046 }),
  .Y({ S7202 })
);
NOR #() 
NOR_2601_ (
  .A({ S7200 }),
  .B({ S7201 }),
  .Y({ S7203 })
);
NAND #() 
NAND_4203_ (
  .A({ S7199 }),
  .B({ S7202 }),
  .Y({ S7204 })
);
NOR #() 
NOR_2602_ (
  .A({ S7199 }),
  .B({ S7202 }),
  .Y({ S7205 })
);
NAND #() 
NAND_4204_ (
  .A({ S7200 }),
  .B({ S7201 }),
  .Y({ S7206 })
);
NOR #() 
NOR_2603_ (
  .A({ S7203 }),
  .B({ S7205 }),
  .Y({ S7207 })
);
NAND #() 
NAND_4205_ (
  .A({ S7204 }),
  .B({ S7206 }),
  .Y({ S7208 })
);
NOR #() 
NOR_2604_ (
  .A({ S7157 }),
  .B({ S7207 }),
  .Y({ S7209 })
);
NAND #() 
NAND_4206_ (
  .A({ S7156 }),
  .B({ S7208 }),
  .Y({ S7210 })
);
NOR #() 
NOR_2605_ (
  .A({ S7156 }),
  .B({ S7208 }),
  .Y({ S7211 })
);
NAND #() 
NAND_4207_ (
  .A({ S7157 }),
  .B({ S7207 }),
  .Y({ S7212 })
);
NOR #() 
NOR_2606_ (
  .A({ S7209 }),
  .B({ S7211 }),
  .Y({ S7213 })
);
NAND #() 
NAND_4208_ (
  .A({ S7210 }),
  .B({ S7212 }),
  .Y({ S7214 })
);
NOR #() 
NOR_2607_ (
  .A({ S7101 }),
  .B({ S7107 }),
  .Y({ S7215 })
);
NAND #() 
NAND_4209_ (
  .A({ S7102 }),
  .B({ S7108 }),
  .Y({ S7216 })
);
NOR #() 
NOR_2608_ (
  .A({ S7025 }),
  .B({ S7029 }),
  .Y({ S7217 })
);
NAND #() 
NAND_4210_ (
  .A({ S7026 }),
  .B({ S7030 }),
  .Y({ S7218 })
);
NOR #() 
NOR_2609_ (
  .A({ S963 }),
  .B({ S2418 }),
  .Y({ S7219 })
);
NAND #() 
NAND_4211_ (
  .A({ datapath_addsubunit_in1_5 }),
  .B({ S2417 }),
  .Y({ S7220 })
);
NOR #() 
NOR_2610_ (
  .A({ S858 }),
  .B({ S2206 }),
  .Y({ S7221 })
);
NAND #() 
NAND_4212_ (
  .A({ datapath_addsubunit_in1_7 }),
  .B({ S2205 }),
  .Y({ S7222 })
);
NOR #() 
NOR_2611_ (
  .A({ S7023 }),
  .B({ S7221 }),
  .Y({ S7223 })
);
NAND #() 
NAND_4213_ (
  .A({ S7024 }),
  .B({ S7222 }),
  .Y({ S7224 })
);
NOR #() 
NOR_2612_ (
  .A({ S858 }),
  .B({ S2312 }),
  .Y({ S7225 })
);
NAND #() 
NAND_4214_ (
  .A({ datapath_addsubunit_in1_7 }),
  .B({ S2311 }),
  .Y({ S7226 })
);
NOR #() 
NOR_2613_ (
  .A({ S7024 }),
  .B({ S7222 }),
  .Y({ S7227 })
);
NAND #() 
NAND_4215_ (
  .A({ S7023 }),
  .B({ S7221 }),
  .Y({ S7228 })
);
NOR #() 
NOR_2614_ (
  .A({ S7223 }),
  .B({ S7227 }),
  .Y({ S7229 })
);
NAND #() 
NAND_4216_ (
  .A({ S7224 }),
  .B({ S7228 }),
  .Y({ S7230 })
);
NOR #() 
NOR_2615_ (
  .A({ S7220 }),
  .B({ S7230 }),
  .Y({ S7231 })
);
NAND #() 
NAND_4217_ (
  .A({ S7219 }),
  .B({ S7229 }),
  .Y({ S7232 })
);
NOR #() 
NOR_2616_ (
  .A({ S7219 }),
  .B({ S7229 }),
  .Y({ S7233 })
);
NAND #() 
NAND_4218_ (
  .A({ S7220 }),
  .B({ S7230 }),
  .Y({ S7234 })
);
NOR #() 
NOR_2617_ (
  .A({ S7231 }),
  .B({ S7233 }),
  .Y({ S7235 })
);
NAND #() 
NAND_4219_ (
  .A({ S7232 }),
  .B({ S7234 }),
  .Y({ S7236 })
);
NOR #() 
NOR_2618_ (
  .A({ S7059 }),
  .B({ S7063 }),
  .Y({ S7237 })
);
NAND #() 
NAND_4220_ (
  .A({ S7060 }),
  .B({ S7064 }),
  .Y({ S7238 })
);
NOR #() 
NOR_2619_ (
  .A({ S7236 }),
  .B({ S7237 }),
  .Y({ S7239 })
);
NAND #() 
NAND_4221_ (
  .A({ S7235 }),
  .B({ S7238 }),
  .Y({ S7240 })
);
NOR #() 
NOR_2620_ (
  .A({ S7235 }),
  .B({ S7238 }),
  .Y({ S7241 })
);
NAND #() 
NAND_4222_ (
  .A({ S7236 }),
  .B({ S7237 }),
  .Y({ S7242 })
);
NOR #() 
NOR_2621_ (
  .A({ S7239 }),
  .B({ S7241 }),
  .Y({ S7243 })
);
NAND #() 
NAND_4223_ (
  .A({ S7240 }),
  .B({ S7242 }),
  .Y({ S7244 })
);
NOR #() 
NOR_2622_ (
  .A({ S7218 }),
  .B({ S7243 }),
  .Y({ S7245 })
);
NAND #() 
NAND_4224_ (
  .A({ S7217 }),
  .B({ S7244 }),
  .Y({ S7246 })
);
NOR #() 
NOR_2623_ (
  .A({ S7217 }),
  .B({ S7244 }),
  .Y({ S7247 })
);
NAND #() 
NAND_4225_ (
  .A({ S7218 }),
  .B({ S7243 }),
  .Y({ S7248 })
);
NOR #() 
NOR_2624_ (
  .A({ S7245 }),
  .B({ S7247 }),
  .Y({ S7249 })
);
NAND #() 
NAND_4226_ (
  .A({ S7246 }),
  .B({ S7248 }),
  .Y({ S7250 })
);
NOR #() 
NOR_2625_ (
  .A({ S7089 }),
  .B({ S7095 }),
  .Y({ S7251 })
);
NAND #() 
NAND_4227_ (
  .A({ S7090 }),
  .B({ S7096 }),
  .Y({ S7252 })
);
NOR #() 
NOR_2626_ (
  .A({ S805 }),
  .B({ S2107 }),
  .Y({ S7253 })
);
NAND #() 
NAND_4228_ (
  .A({ datapath_addsubunit_in1_8 }),
  .B({ S2106 }),
  .Y({ S7254 })
);
NOR #() 
NOR_2627_ (
  .A({ S702 }),
  .B({ S1953 }),
  .Y({ S7255 })
);
NAND #() 
NAND_4229_ (
  .A({ datapath_addsubunit_in1_10 }),
  .B({ S1952 }),
  .Y({ S7256 })
);
NOR #() 
NOR_2628_ (
  .A({ S7057 }),
  .B({ S7255 }),
  .Y({ S7257 })
);
NAND #() 
NAND_4230_ (
  .A({ S7058 }),
  .B({ S7256 }),
  .Y({ S7258 })
);
NAND #() 
NAND_4231_ (
  .A({ datapath_addsubunit_in1_10 }),
  .B({ S1597 }),
  .Y({ S7259 })
);
NOR #() 
NOR_2629_ (
  .A({ S7058 }),
  .B({ S7256 }),
  .Y({ S7260 })
);
NAND #() 
NAND_4232_ (
  .A({ S7057 }),
  .B({ S7255 }),
  .Y({ S7261 })
);
NOR #() 
NOR_2630_ (
  .A({ S7257 }),
  .B({ S7260 }),
  .Y({ S7262 })
);
NAND #() 
NAND_4233_ (
  .A({ S7258 }),
  .B({ S7261 }),
  .Y({ S7263 })
);
NOR #() 
NOR_2631_ (
  .A({ S7254 }),
  .B({ S7263 }),
  .Y({ S7264 })
);
NAND #() 
NAND_4234_ (
  .A({ S7253 }),
  .B({ S7262 }),
  .Y({ S7265 })
);
NOR #() 
NOR_2632_ (
  .A({ S7253 }),
  .B({ S7262 }),
  .Y({ S7266 })
);
NAND #() 
NAND_4235_ (
  .A({ S7254 }),
  .B({ S7263 }),
  .Y({ S7267 })
);
NOR #() 
NOR_2633_ (
  .A({ S7264 }),
  .B({ S7266 }),
  .Y({ S7268 })
);
NAND #() 
NAND_4236_ (
  .A({ S7265 }),
  .B({ S7267 }),
  .Y({ S7269 })
);
NOR #() 
NOR_2634_ (
  .A({ S7079 }),
  .B({ S7083 }),
  .Y({ S7270 })
);
NAND #() 
NAND_4237_ (
  .A({ S7080 }),
  .B({ S7084 }),
  .Y({ S7271 })
);
NOR #() 
NOR_2635_ (
  .A({ S651 }),
  .B({ S1849 }),
  .Y({ S7272 })
);
NAND #() 
NAND_4238_ (
  .A({ datapath_addsubunit_in1_11 }),
  .B({ S1848 }),
  .Y({ S7273 })
);
NOR #() 
NOR_2636_ (
  .A({ S548 }),
  .B({ S1516 }),
  .Y({ S7274 })
);
NAND #() 
NAND_4239_ (
  .A({ datapath_addsubunit_in1_13 }),
  .B({ S1515 }),
  .Y({ S7275 })
);
NOR #() 
NOR_2637_ (
  .A({ S7077 }),
  .B({ S7274 }),
  .Y({ S7276 })
);
NAND #() 
NAND_4240_ (
  .A({ S7078 }),
  .B({ S7275 }),
  .Y({ S7277 })
);
NAND #() 
NAND_4241_ (
  .A({ datapath_addsubunit_in1_13 }),
  .B({ S1745 }),
  .Y({ S7278 })
);
NOR #() 
NOR_2638_ (
  .A({ S7078 }),
  .B({ S7275 }),
  .Y({ S7279 })
);
NAND #() 
NAND_4242_ (
  .A({ S7077 }),
  .B({ S7274 }),
  .Y({ S7280 })
);
NOR #() 
NOR_2639_ (
  .A({ S7276 }),
  .B({ S7279 }),
  .Y({ S7281 })
);
NAND #() 
NAND_4243_ (
  .A({ S7277 }),
  .B({ S7280 }),
  .Y({ S7282 })
);
NOR #() 
NOR_2640_ (
  .A({ S7273 }),
  .B({ S7282 }),
  .Y({ S7283 })
);
NAND #() 
NAND_4244_ (
  .A({ S7272 }),
  .B({ S7281 }),
  .Y({ S7284 })
);
NOR #() 
NOR_2641_ (
  .A({ S7272 }),
  .B({ S7281 }),
  .Y({ S7285 })
);
NAND #() 
NAND_4245_ (
  .A({ S7273 }),
  .B({ S7282 }),
  .Y({ S7286 })
);
NOR #() 
NOR_2642_ (
  .A({ S7283 }),
  .B({ S7285 }),
  .Y({ S7287 })
);
NAND #() 
NAND_4246_ (
  .A({ S7284 }),
  .B({ S7286 }),
  .Y({ S7288 })
);
NOR #() 
NOR_2643_ (
  .A({ S7270 }),
  .B({ S7288 }),
  .Y({ S7289 })
);
NAND #() 
NAND_4247_ (
  .A({ S7271 }),
  .B({ S7287 }),
  .Y({ S7290 })
);
NOR #() 
NOR_2644_ (
  .A({ S7271 }),
  .B({ S7287 }),
  .Y({ S7291 })
);
NAND #() 
NAND_4248_ (
  .A({ S7270 }),
  .B({ S7288 }),
  .Y({ S7292 })
);
NOR #() 
NOR_2645_ (
  .A({ S7289 }),
  .B({ S7291 }),
  .Y({ S7293 })
);
NAND #() 
NAND_4249_ (
  .A({ S7290 }),
  .B({ S7292 }),
  .Y({ S7294 })
);
NOR #() 
NOR_2646_ (
  .A({ S7269 }),
  .B({ S7294 }),
  .Y({ S7295 })
);
NAND #() 
NAND_4250_ (
  .A({ S7268 }),
  .B({ S7293 }),
  .Y({ S7296 })
);
NOR #() 
NOR_2647_ (
  .A({ S7268 }),
  .B({ S7293 }),
  .Y({ S7297 })
);
NAND #() 
NAND_4251_ (
  .A({ S7269 }),
  .B({ S7294 }),
  .Y({ S7298 })
);
NOR #() 
NOR_2648_ (
  .A({ S7295 }),
  .B({ S7297 }),
  .Y({ S7299 })
);
NAND #() 
NAND_4252_ (
  .A({ S7296 }),
  .B({ S7298 }),
  .Y({ S7300 })
);
NOR #() 
NOR_2649_ (
  .A({ S7251 }),
  .B({ S7300 }),
  .Y({ S7301 })
);
NAND #() 
NAND_4253_ (
  .A({ S7252 }),
  .B({ S7299 }),
  .Y({ S7302 })
);
NOR #() 
NOR_2650_ (
  .A({ S7252 }),
  .B({ S7299 }),
  .Y({ S7303 })
);
NAND #() 
NAND_4254_ (
  .A({ S7251 }),
  .B({ S7300 }),
  .Y({ S7304 })
);
NOR #() 
NOR_2651_ (
  .A({ S7301 }),
  .B({ S7303 }),
  .Y({ S7305 })
);
NAND #() 
NAND_4255_ (
  .A({ S7302 }),
  .B({ S7304 }),
  .Y({ S7306 })
);
NOR #() 
NOR_2652_ (
  .A({ S7250 }),
  .B({ S7306 }),
  .Y({ S7307 })
);
NAND #() 
NAND_4256_ (
  .A({ S7249 }),
  .B({ S7305 }),
  .Y({ S7308 })
);
NOR #() 
NOR_2653_ (
  .A({ S7249 }),
  .B({ S7305 }),
  .Y({ S7309 })
);
NAND #() 
NAND_4257_ (
  .A({ S7250 }),
  .B({ S7306 }),
  .Y({ S7310 })
);
NOR #() 
NOR_2654_ (
  .A({ S7307 }),
  .B({ S7309 }),
  .Y({ S7311 })
);
NAND #() 
NAND_4258_ (
  .A({ S7308 }),
  .B({ S7310 }),
  .Y({ S7312 })
);
NOR #() 
NOR_2655_ (
  .A({ S7215 }),
  .B({ S7312 }),
  .Y({ S7313 })
);
NAND #() 
NAND_4259_ (
  .A({ S7216 }),
  .B({ S7311 }),
  .Y({ S7314 })
);
NOR #() 
NOR_2656_ (
  .A({ S7216 }),
  .B({ S7311 }),
  .Y({ S7315 })
);
NAND #() 
NAND_4260_ (
  .A({ S7215 }),
  .B({ S7312 }),
  .Y({ S7316 })
);
NOR #() 
NOR_2657_ (
  .A({ S7313 }),
  .B({ S7315 }),
  .Y({ S7317 })
);
NAND #() 
NAND_4261_ (
  .A({ S7314 }),
  .B({ S7316 }),
  .Y({ S7318 })
);
NOR #() 
NOR_2658_ (
  .A({ S7214 }),
  .B({ S7318 }),
  .Y({ S7319 })
);
NAND #() 
NAND_4262_ (
  .A({ S7213 }),
  .B({ S7317 }),
  .Y({ S7320 })
);
NOR #() 
NOR_2659_ (
  .A({ S7213 }),
  .B({ S7317 }),
  .Y({ S7321 })
);
NAND #() 
NAND_4263_ (
  .A({ S7214 }),
  .B({ S7318 }),
  .Y({ S7322 })
);
NOR #() 
NOR_2660_ (
  .A({ S7319 }),
  .B({ S7321 }),
  .Y({ S7323 })
);
NAND #() 
NAND_4264_ (
  .A({ S7320 }),
  .B({ S7322 }),
  .Y({ S7324 })
);
NOR #() 
NOR_2661_ (
  .A({ S7154 }),
  .B({ S7324 }),
  .Y({ S7325 })
);
NOT #() 
NOT_522_ (
  .A({ S7325 }),
  .Y({ S7326 })
);
NOR #() 
NOR_2662_ (
  .A({ S7155 }),
  .B({ S7323 }),
  .Y({ S7327 })
);
NAND #() 
NAND_4265_ (
  .A({ S7154 }),
  .B({ S7324 }),
  .Y({ S7328 })
);
NOR #() 
NOR_2663_ (
  .A({ S7325 }),
  .B({ S7327 }),
  .Y({ S7329 })
);
NAND #() 
NAND_4266_ (
  .A({ S7326 }),
  .B({ S7328 }),
  .Y({ S7330 })
);
NOR #() 
NOR_2664_ (
  .A({ S7152 }),
  .B({ S7330 }),
  .Y({ S7331 })
);
NOR #() 
NOR_2665_ (
  .A({ S7153 }),
  .B({ S7329 }),
  .Y({ S7332 })
);
NOR #() 
NOR_2666_ (
  .A({ S7331 }),
  .B({ S7332 }),
  .Y({ S7333 })
);
NOT #() 
NOT_523_ (
  .A({ S7333 }),
  .Y({ S7334 })
);
NAND #() 
NAND_4267_ (
  .A({ S7150 }),
  .B({ S7334 }),
  .Y({ S7335 })
);
NAND #() 
NAND_4268_ (
  .A({ S7151 }),
  .B({ S7333 }),
  .Y({ S7336 })
);
NAND #() 
NAND_4269_ (
  .A({ S7335 }),
  .B({ S7336 }),
  .Y({ S7337 })
);
NOR #() 
NOR_2667_ (
  .A({ S7138 }),
  .B({ S7337 }),
  .Y({ S7338 })
);
NOT #() 
NOT_524_ (
  .A({ S7338 }),
  .Y({ S7339 })
);
NAND #() 
NAND_4270_ (
  .A({ S7138 }),
  .B({ S7337 }),
  .Y({ S7340 })
);
NAND #() 
NAND_4271_ (
  .A({ S7339 }),
  .B({ S7340 }),
  .Y({ S7341 })
);
NOR #() 
NOR_2668_ (
  .A({ S7149 }),
  .B({ S7341 }),
  .Y({ S7342 })
);
NAND #() 
NAND_4272_ (
  .A({ S7149 }),
  .B({ S7341 }),
  .Y({ S7343 })
);
NOR #() 
NOR_2669_ (
  .A({ S5949 }),
  .B({ S7342 }),
  .Y({ S7344 })
);
NAND #() 
NAND_4273_ (
  .A({ S7343 }),
  .B({ S7344 }),
  .Y({ S7345 })
);
NAND #() 
NAND_4274_ (
  .A({ datapath_multdivunit_outmdu1_13 }),
  .B({ S5950 }),
  .Y({ S7346 })
);
NOT #() 
NOT_525_ (
  .A({ S7346 }),
  .Y({ S7347 })
);
NOR #() 
NOR_2670_ (
  .A({ S3899 }),
  .B({ S3985 }),
  .Y({ S7348 })
);
NOR #() 
NOR_2671_ (
  .A({ S7347 }),
  .B({ S7348 }),
  .Y({ S7349 })
);
NAND #() 
NAND_4275_ (
  .A({ S7345 }),
  .B({ S7349 }),
  .Y({ S295 })
);
NOR #() 
NOR_2672_ (
  .A({ S7325 }),
  .B({ S7331 }),
  .Y({ S7350 })
);
NOT #() 
NOT_526_ (
  .A({ S7350 }),
  .Y({ S7351 })
);
NOR #() 
NOR_2673_ (
  .A({ S7203 }),
  .B({ S7211 }),
  .Y({ S7352 })
);
NOR #() 
NOR_2674_ (
  .A({ S7166 }),
  .B({ S7352 }),
  .Y({ S7353 })
);
NOT #() 
NOT_527_ (
  .A({ S7353 }),
  .Y({ S7354 })
);
NAND #() 
NAND_4276_ (
  .A({ S7166 }),
  .B({ S7352 }),
  .Y({ S7355 })
);
NAND #() 
NAND_4277_ (
  .A({ S7354 }),
  .B({ S7355 }),
  .Y({ S7356 })
);
NOT #() 
NOT_528_ (
  .A({ S7356 }),
  .Y({ S7357 })
);
NOR #() 
NOR_2675_ (
  .A({ S7313 }),
  .B({ S7319 }),
  .Y({ S7358 })
);
NAND #() 
NAND_4278_ (
  .A({ S7314 }),
  .B({ S7320 }),
  .Y({ S7359 })
);
NOR #() 
NOR_2676_ (
  .A({ S7189 }),
  .B({ S7197 }),
  .Y({ S7360 })
);
NAND #() 
NAND_4279_ (
  .A({ S7190 }),
  .B({ S7198 }),
  .Y({ S7361 })
);
NAND #() 
NAND_4280_ (
  .A({ datapath_addsubunit_in1_0 }),
  .B({ S3036 }),
  .Y({ S7362 })
);
NOT #() 
NOT_529_ (
  .A({ S7362 }),
  .Y({ S7363 })
);
NOR #() 
NOR_2677_ (
  .A({ S1116 }),
  .B({ S2817 }),
  .Y({ S7364 })
);
NOR #() 
NOR_2678_ (
  .A({ S7163 }),
  .B({ S7364 }),
  .Y({ S7365 })
);
NOT #() 
NOT_530_ (
  .A({ S7365 }),
  .Y({ S7366 })
);
NOR #() 
NOR_2679_ (
  .A({ S1116 }),
  .B({ S2920 }),
  .Y({ S7367 })
);
NAND #() 
NAND_4281_ (
  .A({ datapath_addsubunit_in1_2 }),
  .B({ S2919 }),
  .Y({ S7368 })
);
NOR #() 
NOR_2680_ (
  .A({ S7160 }),
  .B({ S7368 }),
  .Y({ S7369 })
);
NAND #() 
NAND_4282_ (
  .A({ S7159 }),
  .B({ S7367 }),
  .Y({ S7370 })
);
NOR #() 
NOR_2681_ (
  .A({ S7365 }),
  .B({ S7369 }),
  .Y({ S7371 })
);
NAND #() 
NAND_4283_ (
  .A({ S7366 }),
  .B({ S7370 }),
  .Y({ S7372 })
);
NOR #() 
NOR_2682_ (
  .A({ S7362 }),
  .B({ S7372 }),
  .Y({ S7373 })
);
NAND #() 
NAND_4284_ (
  .A({ S7363 }),
  .B({ S7371 }),
  .Y({ S7374 })
);
NOR #() 
NOR_2683_ (
  .A({ S7363 }),
  .B({ S7371 }),
  .Y({ S7375 })
);
NAND #() 
NAND_4285_ (
  .A({ S7362 }),
  .B({ S7372 }),
  .Y({ S7376 })
);
NOR #() 
NOR_2684_ (
  .A({ S7373 }),
  .B({ S7375 }),
  .Y({ S7377 })
);
NAND #() 
NAND_4286_ (
  .A({ S7374 }),
  .B({ S7376 }),
  .Y({ S7378 })
);
NOR #() 
NOR_2685_ (
  .A({ S7179 }),
  .B({ S7183 }),
  .Y({ S7379 })
);
NAND #() 
NAND_4287_ (
  .A({ S7180 }),
  .B({ S7184 }),
  .Y({ S7380 })
);
NOR #() 
NOR_2686_ (
  .A({ S1065 }),
  .B({ S2718 }),
  .Y({ S7381 })
);
NAND #() 
NAND_4288_ (
  .A({ datapath_addsubunit_in1_3 }),
  .B({ S2717 }),
  .Y({ S7382 })
);
NOR #() 
NOR_2687_ (
  .A({ S963 }),
  .B({ S2518 }),
  .Y({ S7383 })
);
NAND #() 
NAND_4289_ (
  .A({ datapath_addsubunit_in1_5 }),
  .B({ S2517 }),
  .Y({ S7384 })
);
NOR #() 
NOR_2688_ (
  .A({ S7177 }),
  .B({ S7383 }),
  .Y({ S7385 })
);
NAND #() 
NAND_4290_ (
  .A({ S7178 }),
  .B({ S7384 }),
  .Y({ S7386 })
);
NOR #() 
NOR_2689_ (
  .A({ S963 }),
  .B({ S2618 }),
  .Y({ S7387 })
);
NAND #() 
NAND_4291_ (
  .A({ datapath_addsubunit_in1_5 }),
  .B({ S2617 }),
  .Y({ S7388 })
);
NOR #() 
NOR_2690_ (
  .A({ S7174 }),
  .B({ S7388 }),
  .Y({ S7389 })
);
NAND #() 
NAND_4292_ (
  .A({ S7173 }),
  .B({ S7387 }),
  .Y({ S7390 })
);
NOR #() 
NOR_2691_ (
  .A({ S7385 }),
  .B({ S7389 }),
  .Y({ S7391 })
);
NAND #() 
NAND_4293_ (
  .A({ S7386 }),
  .B({ S7390 }),
  .Y({ S7392 })
);
NOR #() 
NOR_2692_ (
  .A({ S7382 }),
  .B({ S7392 }),
  .Y({ S7393 })
);
NAND #() 
NAND_4294_ (
  .A({ S7381 }),
  .B({ S7391 }),
  .Y({ S7394 })
);
NOR #() 
NOR_2693_ (
  .A({ S7381 }),
  .B({ S7391 }),
  .Y({ S7395 })
);
NAND #() 
NAND_4295_ (
  .A({ S7382 }),
  .B({ S7392 }),
  .Y({ S7396 })
);
NOR #() 
NOR_2694_ (
  .A({ S7393 }),
  .B({ S7395 }),
  .Y({ S7397 })
);
NAND #() 
NAND_4296_ (
  .A({ S7394 }),
  .B({ S7396 }),
  .Y({ S7398 })
);
NOR #() 
NOR_2695_ (
  .A({ S7379 }),
  .B({ S7398 }),
  .Y({ S7399 })
);
NAND #() 
NAND_4297_ (
  .A({ S7380 }),
  .B({ S7397 }),
  .Y({ S7400 })
);
NOR #() 
NOR_2696_ (
  .A({ S7380 }),
  .B({ S7397 }),
  .Y({ S7401 })
);
NAND #() 
NAND_4298_ (
  .A({ S7379 }),
  .B({ S7398 }),
  .Y({ S7402 })
);
NOR #() 
NOR_2697_ (
  .A({ S7399 }),
  .B({ S7401 }),
  .Y({ S7403 })
);
NAND #() 
NAND_4299_ (
  .A({ S7400 }),
  .B({ S7402 }),
  .Y({ S7404 })
);
NOR #() 
NOR_2698_ (
  .A({ S7377 }),
  .B({ S7403 }),
  .Y({ S7405 })
);
NAND #() 
NAND_4300_ (
  .A({ S7378 }),
  .B({ S7404 }),
  .Y({ S7406 })
);
NOR #() 
NOR_2699_ (
  .A({ S7378 }),
  .B({ S7404 }),
  .Y({ S7407 })
);
NAND #() 
NAND_4301_ (
  .A({ S7377 }),
  .B({ S7403 }),
  .Y({ S7408 })
);
NOR #() 
NOR_2700_ (
  .A({ S7405 }),
  .B({ S7407 }),
  .Y({ S7409 })
);
NAND #() 
NAND_4302_ (
  .A({ S7406 }),
  .B({ S7408 }),
  .Y({ S7410 })
);
NOR #() 
NOR_2701_ (
  .A({ S7239 }),
  .B({ S7247 }),
  .Y({ S7411 })
);
NAND #() 
NAND_4303_ (
  .A({ S7240 }),
  .B({ S7248 }),
  .Y({ S7412 })
);
NOR #() 
NOR_2702_ (
  .A({ S7410 }),
  .B({ S7411 }),
  .Y({ S7413 })
);
NAND #() 
NAND_4304_ (
  .A({ S7409 }),
  .B({ S7412 }),
  .Y({ S7414 })
);
NOR #() 
NOR_2703_ (
  .A({ S7409 }),
  .B({ S7412 }),
  .Y({ S7415 })
);
NAND #() 
NAND_4305_ (
  .A({ S7410 }),
  .B({ S7411 }),
  .Y({ S7416 })
);
NOR #() 
NOR_2704_ (
  .A({ S7413 }),
  .B({ S7415 }),
  .Y({ S7417 })
);
NAND #() 
NAND_4306_ (
  .A({ S7414 }),
  .B({ S7416 }),
  .Y({ S7418 })
);
NOR #() 
NOR_2705_ (
  .A({ S7361 }),
  .B({ S7417 }),
  .Y({ S7419 })
);
NAND #() 
NAND_4307_ (
  .A({ S7360 }),
  .B({ S7418 }),
  .Y({ S7420 })
);
NOR #() 
NOR_2706_ (
  .A({ S7360 }),
  .B({ S7418 }),
  .Y({ S7421 })
);
NAND #() 
NAND_4308_ (
  .A({ S7361 }),
  .B({ S7417 }),
  .Y({ S7422 })
);
NOR #() 
NOR_2707_ (
  .A({ S7419 }),
  .B({ S7421 }),
  .Y({ S7423 })
);
NAND #() 
NAND_4309_ (
  .A({ S7420 }),
  .B({ S7422 }),
  .Y({ S7424 })
);
NOR #() 
NOR_2708_ (
  .A({ S7301 }),
  .B({ S7307 }),
  .Y({ S7425 })
);
NAND #() 
NAND_4310_ (
  .A({ S7302 }),
  .B({ S7308 }),
  .Y({ S7426 })
);
NOR #() 
NOR_2709_ (
  .A({ S7227 }),
  .B({ S7231 }),
  .Y({ S7427 })
);
NAND #() 
NAND_4311_ (
  .A({ S7228 }),
  .B({ S7232 }),
  .Y({ S7428 })
);
NOR #() 
NOR_2710_ (
  .A({ S910 }),
  .B({ S2418 }),
  .Y({ S7429 })
);
NAND #() 
NAND_4312_ (
  .A({ datapath_addsubunit_in1_6 }),
  .B({ S2417 }),
  .Y({ S7430 })
);
NOR #() 
NOR_2711_ (
  .A({ S805 }),
  .B({ S2206 }),
  .Y({ S7431 })
);
NAND #() 
NAND_4313_ (
  .A({ datapath_addsubunit_in1_8 }),
  .B({ S2205 }),
  .Y({ S7432 })
);
NOR #() 
NOR_2712_ (
  .A({ S7225 }),
  .B({ S7431 }),
  .Y({ S7433 })
);
NAND #() 
NAND_4314_ (
  .A({ S7226 }),
  .B({ S7432 }),
  .Y({ S7434 })
);
NOR #() 
NOR_2713_ (
  .A({ S805 }),
  .B({ S2312 }),
  .Y({ S7435 })
);
NAND #() 
NAND_4315_ (
  .A({ datapath_addsubunit_in1_8 }),
  .B({ S2311 }),
  .Y({ S7436 })
);
NOR #() 
NOR_2714_ (
  .A({ S7222 }),
  .B({ S7436 }),
  .Y({ S7437 })
);
NAND #() 
NAND_4316_ (
  .A({ S7221 }),
  .B({ S7435 }),
  .Y({ S7438 })
);
NOR #() 
NOR_2715_ (
  .A({ S7433 }),
  .B({ S7437 }),
  .Y({ S7439 })
);
NAND #() 
NAND_4317_ (
  .A({ S7434 }),
  .B({ S7438 }),
  .Y({ S7440 })
);
NOR #() 
NOR_2716_ (
  .A({ S7430 }),
  .B({ S7440 }),
  .Y({ S7441 })
);
NAND #() 
NAND_4318_ (
  .A({ S7429 }),
  .B({ S7439 }),
  .Y({ S7442 })
);
NOR #() 
NOR_2717_ (
  .A({ S7429 }),
  .B({ S7439 }),
  .Y({ S7443 })
);
NAND #() 
NAND_4319_ (
  .A({ S7430 }),
  .B({ S7440 }),
  .Y({ S7444 })
);
NOR #() 
NOR_2718_ (
  .A({ S7441 }),
  .B({ S7443 }),
  .Y({ S7445 })
);
NAND #() 
NAND_4320_ (
  .A({ S7442 }),
  .B({ S7444 }),
  .Y({ S7446 })
);
NOR #() 
NOR_2719_ (
  .A({ S7260 }),
  .B({ S7264 }),
  .Y({ S7447 })
);
NAND #() 
NAND_4321_ (
  .A({ S7261 }),
  .B({ S7265 }),
  .Y({ S7448 })
);
NOR #() 
NOR_2720_ (
  .A({ S7446 }),
  .B({ S7447 }),
  .Y({ S7449 })
);
NAND #() 
NAND_4322_ (
  .A({ S7445 }),
  .B({ S7448 }),
  .Y({ S7450 })
);
NOR #() 
NOR_2721_ (
  .A({ S7445 }),
  .B({ S7448 }),
  .Y({ S7451 })
);
NAND #() 
NAND_4323_ (
  .A({ S7446 }),
  .B({ S7447 }),
  .Y({ S7452 })
);
NOR #() 
NOR_2722_ (
  .A({ S7449 }),
  .B({ S7451 }),
  .Y({ S7453 })
);
NAND #() 
NAND_4324_ (
  .A({ S7450 }),
  .B({ S7452 }),
  .Y({ S7454 })
);
NOR #() 
NOR_2723_ (
  .A({ S7428 }),
  .B({ S7453 }),
  .Y({ S7455 })
);
NAND #() 
NAND_4325_ (
  .A({ S7427 }),
  .B({ S7454 }),
  .Y({ S7456 })
);
NOR #() 
NOR_2724_ (
  .A({ S7427 }),
  .B({ S7454 }),
  .Y({ S7457 })
);
NAND #() 
NAND_4326_ (
  .A({ S7428 }),
  .B({ S7453 }),
  .Y({ S7458 })
);
NOR #() 
NOR_2725_ (
  .A({ S7455 }),
  .B({ S7457 }),
  .Y({ S7459 })
);
NAND #() 
NAND_4327_ (
  .A({ S7456 }),
  .B({ S7458 }),
  .Y({ S7460 })
);
NOR #() 
NOR_2726_ (
  .A({ S7289 }),
  .B({ S7295 }),
  .Y({ S7461 })
);
NAND #() 
NAND_4328_ (
  .A({ S7290 }),
  .B({ S7296 }),
  .Y({ S7462 })
);
NOR #() 
NOR_2727_ (
  .A({ S754 }),
  .B({ S2107 }),
  .Y({ S7463 })
);
NAND #() 
NAND_4329_ (
  .A({ datapath_addsubunit_in1_9 }),
  .B({ S2106 }),
  .Y({ S7464 })
);
NAND #() 
NAND_4330_ (
  .A({ datapath_addsubunit_in1_11 }),
  .B({ S1952 }),
  .Y({ S7465 })
);
NAND #() 
NAND_4331_ (
  .A({ S7259 }),
  .B({ S7465 }),
  .Y({ S7466 })
);
NOT #() 
NOT_531_ (
  .A({ S7466 }),
  .Y({ S7467 })
);
NOR #() 
NOR_2728_ (
  .A({ S651 }),
  .B({ S1598 }),
  .Y({ S7468 })
);
NAND #() 
NAND_4332_ (
  .A({ datapath_addsubunit_in1_11 }),
  .B({ S1597 }),
  .Y({ S7469 })
);
NOR #() 
NOR_2729_ (
  .A({ S7256 }),
  .B({ S7469 }),
  .Y({ S7470 })
);
NAND #() 
NAND_4333_ (
  .A({ S7255 }),
  .B({ S7468 }),
  .Y({ S7471 })
);
NOR #() 
NOR_2730_ (
  .A({ S7467 }),
  .B({ S7470 }),
  .Y({ S7472 })
);
NAND #() 
NAND_4334_ (
  .A({ S7466 }),
  .B({ S7471 }),
  .Y({ S7473 })
);
NOR #() 
NOR_2731_ (
  .A({ S7464 }),
  .B({ S7473 }),
  .Y({ S7474 })
);
NAND #() 
NAND_4335_ (
  .A({ S7463 }),
  .B({ S7472 }),
  .Y({ S7475 })
);
NOR #() 
NOR_2732_ (
  .A({ S7463 }),
  .B({ S7472 }),
  .Y({ S7477 })
);
NAND #() 
NAND_4336_ (
  .A({ S7464 }),
  .B({ S7473 }),
  .Y({ S7478 })
);
NOR #() 
NOR_2733_ (
  .A({ S7474 }),
  .B({ S7477 }),
  .Y({ S7479 })
);
NAND #() 
NAND_4337_ (
  .A({ S7475 }),
  .B({ S7478 }),
  .Y({ S7480 })
);
NOR #() 
NOR_2734_ (
  .A({ S7279 }),
  .B({ S7283 }),
  .Y({ S7481 })
);
NAND #() 
NAND_4338_ (
  .A({ S7280 }),
  .B({ S7284 }),
  .Y({ S7482 })
);
NOR #() 
NOR_2735_ (
  .A({ S599 }),
  .B({ S1849 }),
  .Y({ S7483 })
);
NAND #() 
NAND_4339_ (
  .A({ datapath_addsubunit_in1_12 }),
  .B({ S1848 }),
  .Y({ S7484 })
);
NAND #() 
NAND_4340_ (
  .A({ datapath_addsubunit_in1_14 }),
  .B({ S1515 }),
  .Y({ S7485 })
);
NAND #() 
NAND_4341_ (
  .A({ S7278 }),
  .B({ S7485 }),
  .Y({ S7486 })
);
NOT #() 
NOT_532_ (
  .A({ S7486 }),
  .Y({ S7488 })
);
NOR #() 
NOR_2736_ (
  .A({ S492 }),
  .B({ S1746 }),
  .Y({ S7489 })
);
NAND #() 
NAND_4342_ (
  .A({ datapath_addsubunit_in1_14 }),
  .B({ S1745 }),
  .Y({ S7490 })
);
NOR #() 
NOR_2737_ (
  .A({ S7275 }),
  .B({ S7490 }),
  .Y({ S7491 })
);
NAND #() 
NAND_4343_ (
  .A({ S7274 }),
  .B({ S7489 }),
  .Y({ S7492 })
);
NOR #() 
NOR_2738_ (
  .A({ S7488 }),
  .B({ S7491 }),
  .Y({ S7493 })
);
NAND #() 
NAND_4344_ (
  .A({ S7486 }),
  .B({ S7492 }),
  .Y({ S7494 })
);
NOR #() 
NOR_2739_ (
  .A({ S7484 }),
  .B({ S7494 }),
  .Y({ S7495 })
);
NAND #() 
NAND_4345_ (
  .A({ S7483 }),
  .B({ S7493 }),
  .Y({ S7496 })
);
NOR #() 
NOR_2740_ (
  .A({ S7483 }),
  .B({ S7493 }),
  .Y({ S7497 })
);
NAND #() 
NAND_4346_ (
  .A({ S7484 }),
  .B({ S7494 }),
  .Y({ S7499 })
);
NOR #() 
NOR_2741_ (
  .A({ S7495 }),
  .B({ S7497 }),
  .Y({ S7500 })
);
NAND #() 
NAND_4347_ (
  .A({ S7496 }),
  .B({ S7499 }),
  .Y({ S7501 })
);
NOR #() 
NOR_2742_ (
  .A({ S7481 }),
  .B({ S7501 }),
  .Y({ S7502 })
);
NAND #() 
NAND_4348_ (
  .A({ S7482 }),
  .B({ S7500 }),
  .Y({ S7503 })
);
NOR #() 
NOR_2743_ (
  .A({ S7482 }),
  .B({ S7500 }),
  .Y({ S7504 })
);
NAND #() 
NAND_4349_ (
  .A({ S7481 }),
  .B({ S7501 }),
  .Y({ S7505 })
);
NOR #() 
NOR_2744_ (
  .A({ S7502 }),
  .B({ S7504 }),
  .Y({ S7506 })
);
NAND #() 
NAND_4350_ (
  .A({ S7503 }),
  .B({ S7505 }),
  .Y({ S7507 })
);
NOR #() 
NOR_2745_ (
  .A({ S7480 }),
  .B({ S7507 }),
  .Y({ S7508 })
);
NAND #() 
NAND_4351_ (
  .A({ S7479 }),
  .B({ S7506 }),
  .Y({ S7510 })
);
NOR #() 
NOR_2746_ (
  .A({ S7479 }),
  .B({ S7506 }),
  .Y({ S7511 })
);
NAND #() 
NAND_4352_ (
  .A({ S7480 }),
  .B({ S7507 }),
  .Y({ S7512 })
);
NOR #() 
NOR_2747_ (
  .A({ S7508 }),
  .B({ S7511 }),
  .Y({ S7513 })
);
NAND #() 
NAND_4353_ (
  .A({ S7510 }),
  .B({ S7512 }),
  .Y({ S7514 })
);
NOR #() 
NOR_2748_ (
  .A({ S7461 }),
  .B({ S7514 }),
  .Y({ S7515 })
);
NAND #() 
NAND_4354_ (
  .A({ S7462 }),
  .B({ S7513 }),
  .Y({ S7516 })
);
NOR #() 
NOR_2749_ (
  .A({ S7462 }),
  .B({ S7513 }),
  .Y({ S7517 })
);
NAND #() 
NAND_4355_ (
  .A({ S7461 }),
  .B({ S7514 }),
  .Y({ S7518 })
);
NOR #() 
NOR_2750_ (
  .A({ S7515 }),
  .B({ S7517 }),
  .Y({ S7519 })
);
NAND #() 
NAND_4356_ (
  .A({ S7516 }),
  .B({ S7518 }),
  .Y({ S7521 })
);
NOR #() 
NOR_2751_ (
  .A({ S7460 }),
  .B({ S7521 }),
  .Y({ S7522 })
);
NAND #() 
NAND_4357_ (
  .A({ S7459 }),
  .B({ S7519 }),
  .Y({ S7523 })
);
NOR #() 
NOR_2752_ (
  .A({ S7459 }),
  .B({ S7519 }),
  .Y({ S7524 })
);
NAND #() 
NAND_4358_ (
  .A({ S7460 }),
  .B({ S7521 }),
  .Y({ S7525 })
);
NOR #() 
NOR_2753_ (
  .A({ S7522 }),
  .B({ S7524 }),
  .Y({ S7526 })
);
NAND #() 
NAND_4359_ (
  .A({ S7523 }),
  .B({ S7525 }),
  .Y({ S7527 })
);
NOR #() 
NOR_2754_ (
  .A({ S7425 }),
  .B({ S7527 }),
  .Y({ S7528 })
);
NAND #() 
NAND_4360_ (
  .A({ S7426 }),
  .B({ S7526 }),
  .Y({ S7529 })
);
NOR #() 
NOR_2755_ (
  .A({ S7426 }),
  .B({ S7526 }),
  .Y({ S7530 })
);
NAND #() 
NAND_4361_ (
  .A({ S7425 }),
  .B({ S7527 }),
  .Y({ S7532 })
);
NOR #() 
NOR_2756_ (
  .A({ S7528 }),
  .B({ S7530 }),
  .Y({ S7533 })
);
NAND #() 
NAND_4362_ (
  .A({ S7529 }),
  .B({ S7532 }),
  .Y({ S7534 })
);
NOR #() 
NOR_2757_ (
  .A({ S7424 }),
  .B({ S7534 }),
  .Y({ S7535 })
);
NAND #() 
NAND_4363_ (
  .A({ S7423 }),
  .B({ S7533 }),
  .Y({ S7536 })
);
NOR #() 
NOR_2758_ (
  .A({ S7423 }),
  .B({ S7533 }),
  .Y({ S7537 })
);
NAND #() 
NAND_4364_ (
  .A({ S7424 }),
  .B({ S7534 }),
  .Y({ S7538 })
);
NOR #() 
NOR_2759_ (
  .A({ S7535 }),
  .B({ S7537 }),
  .Y({ S7539 })
);
NAND #() 
NAND_4365_ (
  .A({ S7536 }),
  .B({ S7538 }),
  .Y({ S7540 })
);
NOR #() 
NOR_2760_ (
  .A({ S7358 }),
  .B({ S7540 }),
  .Y({ S7541 })
);
NAND #() 
NAND_4366_ (
  .A({ S7359 }),
  .B({ S7539 }),
  .Y({ S7543 })
);
NAND #() 
NAND_4367_ (
  .A({ S7358 }),
  .B({ S7540 }),
  .Y({ S7544 })
);
NAND #() 
NAND_4368_ (
  .A({ S7543 }),
  .B({ S7544 }),
  .Y({ S7545 })
);
NOT #() 
NOT_533_ (
  .A({ S7545 }),
  .Y({ S7546 })
);
NAND #() 
NAND_4369_ (
  .A({ S7357 }),
  .B({ S7546 }),
  .Y({ S7547 })
);
NOT #() 
NOT_534_ (
  .A({ S7547 }),
  .Y({ S7548 })
);
NAND #() 
NAND_4370_ (
  .A({ S7356 }),
  .B({ S7545 }),
  .Y({ S7549 })
);
NAND #() 
NAND_4371_ (
  .A({ S7547 }),
  .B({ S7549 }),
  .Y({ S7550 })
);
NOT #() 
NOT_535_ (
  .A({ S7550 }),
  .Y({ S7551 })
);
NAND #() 
NAND_4372_ (
  .A({ S7350 }),
  .B({ S7550 }),
  .Y({ S7552 })
);
NAND #() 
NAND_4373_ (
  .A({ S7351 }),
  .B({ S7551 }),
  .Y({ S7554 })
);
NAND #() 
NAND_4374_ (
  .A({ S7552 }),
  .B({ S7554 }),
  .Y({ S7555 })
);
NOR #() 
NOR_2761_ (
  .A({ S7336 }),
  .B({ S7555 }),
  .Y({ S7556 })
);
NOT #() 
NOT_536_ (
  .A({ S7556 }),
  .Y({ S7557 })
);
NAND #() 
NAND_4375_ (
  .A({ S7336 }),
  .B({ S7555 }),
  .Y({ S7558 })
);
NAND #() 
NAND_4376_ (
  .A({ S7557 }),
  .B({ S7558 }),
  .Y({ S7559 })
);
NOR #() 
NOR_2762_ (
  .A({ S7338 }),
  .B({ S7342 }),
  .Y({ S7560 })
);
NAND #() 
NAND_4377_ (
  .A({ S7559 }),
  .B({ S7560 }),
  .Y({ S7561 })
);
NOR #() 
NOR_2763_ (
  .A({ S7559 }),
  .B({ S7560 }),
  .Y({ S7562 })
);
NOR #() 
NOR_2764_ (
  .A({ S5949 }),
  .B({ S7562 }),
  .Y({ S7563 })
);
NAND #() 
NAND_4378_ (
  .A({ S7561 }),
  .B({ S7563 }),
  .Y({ S7565 })
);
NAND #() 
NAND_4379_ (
  .A({ datapath_multdivunit_outmdu1_14 }),
  .B({ S5950 }),
  .Y({ S7566 })
);
NOT #() 
NOT_537_ (
  .A({ S7566 }),
  .Y({ S7567 })
);
NOR #() 
NOR_2765_ (
  .A({ S3899 }),
  .B({ S3945 }),
  .Y({ S7568 })
);
NOR #() 
NOR_2766_ (
  .A({ S7567 }),
  .B({ S7568 }),
  .Y({ S7569 })
);
NAND #() 
NAND_4380_ (
  .A({ S7565 }),
  .B({ S7569 }),
  .Y({ S296 })
);
NOR #() 
NOR_2767_ (
  .A({ S7556 }),
  .B({ S7562 }),
  .Y({ S7570 })
);
NOR #() 
NOR_2768_ (
  .A({ S7541 }),
  .B({ S7548 }),
  .Y({ S7571 })
);
NAND #() 
NAND_4381_ (
  .A({ S7543 }),
  .B({ S7547 }),
  .Y({ S7572 })
);
NOR #() 
NOR_2769_ (
  .A({ S7449 }),
  .B({ S7457 }),
  .Y({ S7573 })
);
NAND #() 
NAND_4382_ (
  .A({ S7450 }),
  .B({ S7458 }),
  .Y({ S7575 })
);
NOR #() 
NOR_2770_ (
  .A({ S548 }),
  .B({ S1849 }),
  .Y({ S7576 })
);
NAND #() 
NAND_4383_ (
  .A({ datapath_addsubunit_in1_13 }),
  .B({ S1848 }),
  .Y({ S7577 })
);
NOR #() 
NOR_2771_ (
  .A({ S1304 }),
  .B({ S1516 }),
  .Y({ S7578 })
);
NAND #() 
NAND_4384_ (
  .A({ datapath_addsubunit_in1_15 }),
  .B({ S1515 }),
  .Y({ S7579 })
);
NOR #() 
NOR_2772_ (
  .A({ S7490 }),
  .B({ S7578 }),
  .Y({ S7580 })
);
NAND #() 
NAND_4385_ (
  .A({ S7489 }),
  .B({ S7579 }),
  .Y({ S7581 })
);
NOR #() 
NOR_2773_ (
  .A({ S7489 }),
  .B({ S7579 }),
  .Y({ S7582 })
);
NAND #() 
NAND_4386_ (
  .A({ S7490 }),
  .B({ S7578 }),
  .Y({ S7583 })
);
NOR #() 
NOR_2774_ (
  .A({ S7580 }),
  .B({ S7582 }),
  .Y({ S7584 })
);
NAND #() 
NAND_4387_ (
  .A({ S7581 }),
  .B({ S7583 }),
  .Y({ S7586 })
);
NOR #() 
NOR_2775_ (
  .A({ S599 }),
  .B({ S1953 }),
  .Y({ S7587 })
);
NAND #() 
NAND_4388_ (
  .A({ datapath_addsubunit_in1_12 }),
  .B({ S1952 }),
  .Y({ S7588 })
);
NOR #() 
NOR_2776_ (
  .A({ S7469 }),
  .B({ S7587 }),
  .Y({ S7589 })
);
NAND #() 
NAND_4389_ (
  .A({ S7468 }),
  .B({ S7588 }),
  .Y({ S7590 })
);
NOR #() 
NOR_2777_ (
  .A({ S7468 }),
  .B({ S7588 }),
  .Y({ S7591 })
);
NAND #() 
NAND_4390_ (
  .A({ S7469 }),
  .B({ S7587 }),
  .Y({ S7592 })
);
NOR #() 
NOR_2778_ (
  .A({ S7589 }),
  .B({ S7591 }),
  .Y({ S7593 })
);
NAND #() 
NAND_4391_ (
  .A({ S7590 }),
  .B({ S7592 }),
  .Y({ S7594 })
);
NOR #() 
NOR_2779_ (
  .A({ S7584 }),
  .B({ S7593 }),
  .Y({ S7595 })
);
NAND #() 
NAND_4392_ (
  .A({ S7586 }),
  .B({ S7594 }),
  .Y({ S7597 })
);
NOR #() 
NOR_2780_ (
  .A({ S7586 }),
  .B({ S7594 }),
  .Y({ S7598 })
);
NAND #() 
NAND_4393_ (
  .A({ S7584 }),
  .B({ S7593 }),
  .Y({ S7599 })
);
NOR #() 
NOR_2781_ (
  .A({ S7595 }),
  .B({ S7598 }),
  .Y({ S7600 })
);
NAND #() 
NAND_4394_ (
  .A({ S7597 }),
  .B({ S7599 }),
  .Y({ S7601 })
);
NOR #() 
NOR_2782_ (
  .A({ S7576 }),
  .B({ S7601 }),
  .Y({ S7602 })
);
NAND #() 
NAND_4395_ (
  .A({ S7577 }),
  .B({ S7600 }),
  .Y({ S7603 })
);
NOR #() 
NOR_2783_ (
  .A({ S7577 }),
  .B({ S7600 }),
  .Y({ S7604 })
);
NAND #() 
NAND_4396_ (
  .A({ S7576 }),
  .B({ S7601 }),
  .Y({ S7605 })
);
NOR #() 
NOR_2784_ (
  .A({ S7602 }),
  .B({ S7604 }),
  .Y({ S7606 })
);
NAND #() 
NAND_4397_ (
  .A({ S7603 }),
  .B({ S7605 }),
  .Y({ S7608 })
);
NOR #() 
NOR_2785_ (
  .A({ S702 }),
  .B({ S2107 }),
  .Y({ S7609 })
);
NAND #() 
NAND_4398_ (
  .A({ datapath_addsubunit_in1_10 }),
  .B({ S2106 }),
  .Y({ S7610 })
);
NOR #() 
NOR_2786_ (
  .A({ S7491 }),
  .B({ S7495 }),
  .Y({ S7611 })
);
NAND #() 
NAND_4399_ (
  .A({ S7492 }),
  .B({ S7496 }),
  .Y({ S7612 })
);
NOR #() 
NOR_2787_ (
  .A({ S7609 }),
  .B({ S7611 }),
  .Y({ S7613 })
);
NAND #() 
NAND_4400_ (
  .A({ S7610 }),
  .B({ S7612 }),
  .Y({ S7614 })
);
NOR #() 
NOR_2788_ (
  .A({ S7610 }),
  .B({ S7612 }),
  .Y({ S7615 })
);
NAND #() 
NAND_4401_ (
  .A({ S7609 }),
  .B({ S7611 }),
  .Y({ S7616 })
);
NOR #() 
NOR_2789_ (
  .A({ S7613 }),
  .B({ S7615 }),
  .Y({ S7617 })
);
NAND #() 
NAND_4402_ (
  .A({ S7614 }),
  .B({ S7616 }),
  .Y({ S7619 })
);
NOR #() 
NOR_2790_ (
  .A({ S7470 }),
  .B({ S7474 }),
  .Y({ S7620 })
);
NAND #() 
NAND_4403_ (
  .A({ S7471 }),
  .B({ S7475 }),
  .Y({ S7621 })
);
NOR #() 
NOR_2791_ (
  .A({ S858 }),
  .B({ S2418 }),
  .Y({ S7622 })
);
NAND #() 
NAND_4404_ (
  .A({ datapath_addsubunit_in1_7 }),
  .B({ S2417 }),
  .Y({ S7623 })
);
NOR #() 
NOR_2792_ (
  .A({ S754 }),
  .B({ S2206 }),
  .Y({ S7624 })
);
NAND #() 
NAND_4405_ (
  .A({ datapath_addsubunit_in1_9 }),
  .B({ S2205 }),
  .Y({ S7625 })
);
NOR #() 
NOR_2793_ (
  .A({ S7435 }),
  .B({ S7625 }),
  .Y({ S7626 })
);
NAND #() 
NAND_4406_ (
  .A({ S7436 }),
  .B({ S7624 }),
  .Y({ S7627 })
);
NOR #() 
NOR_2794_ (
  .A({ S7436 }),
  .B({ S7624 }),
  .Y({ S7628 })
);
NAND #() 
NAND_4407_ (
  .A({ S7435 }),
  .B({ S7625 }),
  .Y({ S7630 })
);
NOR #() 
NOR_2795_ (
  .A({ S7626 }),
  .B({ S7628 }),
  .Y({ S7631 })
);
NAND #() 
NAND_4408_ (
  .A({ S7627 }),
  .B({ S7630 }),
  .Y({ S7632 })
);
NOR #() 
NOR_2796_ (
  .A({ S7623 }),
  .B({ S7632 }),
  .Y({ S7633 })
);
NAND #() 
NAND_4409_ (
  .A({ S7622 }),
  .B({ S7631 }),
  .Y({ S7634 })
);
NOR #() 
NOR_2797_ (
  .A({ S7622 }),
  .B({ S7631 }),
  .Y({ S7635 })
);
NAND #() 
NAND_4410_ (
  .A({ S7623 }),
  .B({ S7632 }),
  .Y({ S7636 })
);
NOR #() 
NOR_2798_ (
  .A({ S7633 }),
  .B({ S7635 }),
  .Y({ S7637 })
);
NAND #() 
NAND_4411_ (
  .A({ S7634 }),
  .B({ S7636 }),
  .Y({ S7638 })
);
NOR #() 
NOR_2799_ (
  .A({ S7620 }),
  .B({ S7637 }),
  .Y({ S7639 })
);
NAND #() 
NAND_4412_ (
  .A({ S7621 }),
  .B({ S7638 }),
  .Y({ S7641 })
);
NOR #() 
NOR_2800_ (
  .A({ S7621 }),
  .B({ S7638 }),
  .Y({ S7642 })
);
NAND #() 
NAND_4413_ (
  .A({ S7620 }),
  .B({ S7637 }),
  .Y({ S7643 })
);
NOR #() 
NOR_2801_ (
  .A({ S7639 }),
  .B({ S7642 }),
  .Y({ S7644 })
);
NAND #() 
NAND_4414_ (
  .A({ S7641 }),
  .B({ S7643 }),
  .Y({ S7645 })
);
NOR #() 
NOR_2802_ (
  .A({ S7617 }),
  .B({ S7645 }),
  .Y({ S7646 })
);
NAND #() 
NAND_4415_ (
  .A({ S7619 }),
  .B({ S7644 }),
  .Y({ S7647 })
);
NOR #() 
NOR_2803_ (
  .A({ S7619 }),
  .B({ S7644 }),
  .Y({ S7648 })
);
NAND #() 
NAND_4416_ (
  .A({ S7617 }),
  .B({ S7645 }),
  .Y({ S7649 })
);
NOR #() 
NOR_2804_ (
  .A({ S7646 }),
  .B({ S7648 }),
  .Y({ S7650 })
);
NAND #() 
NAND_4417_ (
  .A({ S7647 }),
  .B({ S7649 }),
  .Y({ S7652 })
);
NOR #() 
NOR_2805_ (
  .A({ S7606 }),
  .B({ S7650 }),
  .Y({ S7653 })
);
NAND #() 
NAND_4418_ (
  .A({ S7608 }),
  .B({ S7652 }),
  .Y({ S7654 })
);
NOR #() 
NOR_2806_ (
  .A({ S7608 }),
  .B({ S7652 }),
  .Y({ S7655 })
);
NAND #() 
NAND_4419_ (
  .A({ S7606 }),
  .B({ S7650 }),
  .Y({ S7656 })
);
NOR #() 
NOR_2807_ (
  .A({ S7653 }),
  .B({ S7655 }),
  .Y({ S7657 })
);
NAND #() 
NAND_4420_ (
  .A({ S7654 }),
  .B({ S7656 }),
  .Y({ S7658 })
);
NOR #() 
NOR_2808_ (
  .A({ S7573 }),
  .B({ S7657 }),
  .Y({ S7659 })
);
NAND #() 
NAND_4421_ (
  .A({ S7575 }),
  .B({ S7658 }),
  .Y({ S7660 })
);
NOR #() 
NOR_2809_ (
  .A({ S7575 }),
  .B({ S7658 }),
  .Y({ S7661 })
);
NAND #() 
NAND_4422_ (
  .A({ S7573 }),
  .B({ S7657 }),
  .Y({ S7663 })
);
NOR #() 
NOR_2810_ (
  .A({ S7659 }),
  .B({ S7661 }),
  .Y({ S7664 })
);
NAND #() 
NAND_4423_ (
  .A({ S7660 }),
  .B({ S7663 }),
  .Y({ S7665 })
);
NOR #() 
NOR_2811_ (
  .A({ S1065 }),
  .B({ S2817 }),
  .Y({ S7666 })
);
NAND #() 
NAND_4424_ (
  .A({ datapath_addsubunit_in1_3 }),
  .B({ S2816 }),
  .Y({ S7667 })
);
NOR #() 
NOR_2812_ (
  .A({ S7367 }),
  .B({ S7667 }),
  .Y({ S7668 })
);
NAND #() 
NAND_4425_ (
  .A({ S7368 }),
  .B({ S7666 }),
  .Y({ S7669 })
);
NOR #() 
NOR_2813_ (
  .A({ S7368 }),
  .B({ S7666 }),
  .Y({ S7670 })
);
NAND #() 
NAND_4426_ (
  .A({ S7367 }),
  .B({ S7667 }),
  .Y({ S7671 })
);
NOR #() 
NOR_2814_ (
  .A({ S7668 }),
  .B({ S7670 }),
  .Y({ S7672 })
);
NAND #() 
NAND_4427_ (
  .A({ S7669 }),
  .B({ S7671 }),
  .Y({ S7674 })
);
NOR #() 
NOR_2815_ (
  .A({ S910 }),
  .B({ S2518 }),
  .Y({ S7675 })
);
NAND #() 
NAND_4428_ (
  .A({ datapath_addsubunit_in1_6 }),
  .B({ S2517 }),
  .Y({ S7676 })
);
NOR #() 
NOR_2816_ (
  .A({ S7387 }),
  .B({ S7675 }),
  .Y({ S7677 })
);
NAND #() 
NAND_4429_ (
  .A({ S7388 }),
  .B({ S7676 }),
  .Y({ S7678 })
);
NOR #() 
NOR_2817_ (
  .A({ S7388 }),
  .B({ S7676 }),
  .Y({ S7679 })
);
NAND #() 
NAND_4430_ (
  .A({ S7387 }),
  .B({ S7675 }),
  .Y({ S7680 })
);
NOR #() 
NOR_2818_ (
  .A({ S7677 }),
  .B({ S7679 }),
  .Y({ S7681 })
);
NAND #() 
NAND_4431_ (
  .A({ S7678 }),
  .B({ S7680 }),
  .Y({ S7682 })
);
NOR #() 
NOR_2819_ (
  .A({ S1013 }),
  .B({ S2718 }),
  .Y({ S7683 })
);
NAND #() 
NAND_4432_ (
  .A({ datapath_addsubunit_in1_4 }),
  .B({ S2717 }),
  .Y({ S7685 })
);
NOR #() 
NOR_2820_ (
  .A({ S7672 }),
  .B({ S7685 }),
  .Y({ S7686 })
);
NAND #() 
NAND_4433_ (
  .A({ S7674 }),
  .B({ S7683 }),
  .Y({ S7687 })
);
NOR #() 
NOR_2821_ (
  .A({ S7674 }),
  .B({ S7683 }),
  .Y({ S7688 })
);
NAND #() 
NAND_4434_ (
  .A({ S7672 }),
  .B({ S7685 }),
  .Y({ S7689 })
);
NOR #() 
NOR_2822_ (
  .A({ S7686 }),
  .B({ S7688 }),
  .Y({ S7690 })
);
NAND #() 
NAND_4435_ (
  .A({ S7687 }),
  .B({ S7689 }),
  .Y({ S7691 })
);
NOR #() 
NOR_2823_ (
  .A({ S7682 }),
  .B({ S7691 }),
  .Y({ S7692 })
);
NAND #() 
NAND_4436_ (
  .A({ S7681 }),
  .B({ S7690 }),
  .Y({ S7693 })
);
NOR #() 
NOR_2824_ (
  .A({ S7681 }),
  .B({ S7690 }),
  .Y({ S7694 })
);
NAND #() 
NAND_4437_ (
  .A({ S7682 }),
  .B({ S7691 }),
  .Y({ S7696 })
);
NAND #() 
NAND_4438_ (
  .A({ S7693 }),
  .B({ S7696 }),
  .Y({ S7697 })
);
NOR #() 
NOR_2825_ (
  .A({ S7692 }),
  .B({ S7694 }),
  .Y({ S7698 })
);
NAND #() 
NAND_4439_ (
  .A({ datapath_addsubunit_in1_1 }),
  .B({ S3036 }),
  .Y({ S7699 })
);
NOT #() 
NOT_538_ (
  .A({ S7699 }),
  .Y({ S7700 })
);
NOR #() 
NOR_2826_ (
  .A({ S7389 }),
  .B({ S7393 }),
  .Y({ S7701 })
);
NAND #() 
NAND_4440_ (
  .A({ S7390 }),
  .B({ S7394 }),
  .Y({ S7702 })
);
NOR #() 
NOR_2827_ (
  .A({ S7699 }),
  .B({ S7702 }),
  .Y({ S7703 })
);
NAND #() 
NAND_4441_ (
  .A({ S7700 }),
  .B({ S7701 }),
  .Y({ S7704 })
);
NOR #() 
NOR_2828_ (
  .A({ S7700 }),
  .B({ S7701 }),
  .Y({ S7705 })
);
NAND #() 
NAND_4442_ (
  .A({ S7699 }),
  .B({ S7702 }),
  .Y({ S7707 })
);
NOR #() 
NOR_2829_ (
  .A({ S7703 }),
  .B({ S7705 }),
  .Y({ S7708 })
);
NAND #() 
NAND_4443_ (
  .A({ S7704 }),
  .B({ S7707 }),
  .Y({ S7709 })
);
NOR #() 
NOR_2830_ (
  .A({ S7697 }),
  .B({ S7709 }),
  .Y({ S7710 })
);
NAND #() 
NAND_4444_ (
  .A({ S7698 }),
  .B({ S7708 }),
  .Y({ S7711 })
);
NOR #() 
NOR_2831_ (
  .A({ S7698 }),
  .B({ S7708 }),
  .Y({ S7712 })
);
NAND #() 
NAND_4445_ (
  .A({ S7697 }),
  .B({ S7709 }),
  .Y({ S7713 })
);
NOR #() 
NOR_2832_ (
  .A({ S7710 }),
  .B({ S7712 }),
  .Y({ S7714 })
);
NAND #() 
NAND_4446_ (
  .A({ S7711 }),
  .B({ S7713 }),
  .Y({ S7715 })
);
NOR #() 
NOR_2833_ (
  .A({ S7437 }),
  .B({ S7441 }),
  .Y({ S7716 })
);
NAND #() 
NAND_4447_ (
  .A({ S7438 }),
  .B({ S7442 }),
  .Y({ S7718 })
);
NOR #() 
NOR_2834_ (
  .A({ S7502 }),
  .B({ S7508 }),
  .Y({ S7719 })
);
NAND #() 
NAND_4448_ (
  .A({ S7503 }),
  .B({ S7510 }),
  .Y({ S7720 })
);
NOR #() 
NOR_2835_ (
  .A({ S7718 }),
  .B({ S7720 }),
  .Y({ S7721 })
);
NAND #() 
NAND_4449_ (
  .A({ S7716 }),
  .B({ S7719 }),
  .Y({ S7722 })
);
NOR #() 
NOR_2836_ (
  .A({ S7716 }),
  .B({ S7719 }),
  .Y({ S7723 })
);
NAND #() 
NAND_4450_ (
  .A({ S7718 }),
  .B({ S7720 }),
  .Y({ S7724 })
);
NOR #() 
NOR_2837_ (
  .A({ S7721 }),
  .B({ S7723 }),
  .Y({ S7725 })
);
NAND #() 
NAND_4451_ (
  .A({ S7722 }),
  .B({ S7724 }),
  .Y({ S7726 })
);
NOR #() 
NOR_2838_ (
  .A({ S7714 }),
  .B({ S7726 }),
  .Y({ S7727 })
);
NAND #() 
NAND_4452_ (
  .A({ S7715 }),
  .B({ S7725 }),
  .Y({ S7729 })
);
NOR #() 
NOR_2839_ (
  .A({ S7715 }),
  .B({ S7725 }),
  .Y({ S7730 })
);
NAND #() 
NAND_4453_ (
  .A({ S7714 }),
  .B({ S7726 }),
  .Y({ S7731 })
);
NOR #() 
NOR_2840_ (
  .A({ S7727 }),
  .B({ S7730 }),
  .Y({ S7732 })
);
NAND #() 
NAND_4454_ (
  .A({ S7729 }),
  .B({ S7731 }),
  .Y({ S7733 })
);
NOR #() 
NOR_2841_ (
  .A({ S7664 }),
  .B({ S7733 }),
  .Y({ S7734 })
);
NAND #() 
NAND_4455_ (
  .A({ S7665 }),
  .B({ S7732 }),
  .Y({ S7735 })
);
NOR #() 
NOR_2842_ (
  .A({ S7665 }),
  .B({ S7732 }),
  .Y({ S7736 })
);
NAND #() 
NAND_4456_ (
  .A({ S7664 }),
  .B({ S7733 }),
  .Y({ S7737 })
);
NOR #() 
NOR_2843_ (
  .A({ S7734 }),
  .B({ S7736 }),
  .Y({ S7738 })
);
NAND #() 
NAND_4457_ (
  .A({ S7735 }),
  .B({ S7737 }),
  .Y({ S7740 })
);
NOR #() 
NOR_2844_ (
  .A({ S7528 }),
  .B({ S7535 }),
  .Y({ S7741 })
);
NAND #() 
NAND_4458_ (
  .A({ S7529 }),
  .B({ S7536 }),
  .Y({ S7742 })
);
NOR #() 
NOR_2845_ (
  .A({ S7515 }),
  .B({ S7522 }),
  .Y({ S7743 })
);
NAND #() 
NAND_4459_ (
  .A({ S7516 }),
  .B({ S7523 }),
  .Y({ S7744 })
);
NOR #() 
NOR_2846_ (
  .A({ S1220 }),
  .B({ S3142 }),
  .Y({ S7745 })
);
NAND #() 
NAND_4460_ (
  .A({ datapath_addsubunit_in1_0 }),
  .B({ S3141 }),
  .Y({ S7746 })
);
NOR #() 
NOR_2847_ (
  .A({ S7369 }),
  .B({ S7373 }),
  .Y({ S7747 })
);
NAND #() 
NAND_4461_ (
  .A({ S7370 }),
  .B({ S7374 }),
  .Y({ S7748 })
);
NOR #() 
NOR_2848_ (
  .A({ S7745 }),
  .B({ S7748 }),
  .Y({ S7749 })
);
NAND #() 
NAND_4462_ (
  .A({ S7746 }),
  .B({ S7747 }),
  .Y({ S7751 })
);
NOR #() 
NOR_2849_ (
  .A({ S7746 }),
  .B({ S7747 }),
  .Y({ S7752 })
);
NAND #() 
NAND_4463_ (
  .A({ S7745 }),
  .B({ S7748 }),
  .Y({ S7753 })
);
NOR #() 
NOR_2850_ (
  .A({ S7749 }),
  .B({ S7752 }),
  .Y({ S7754 })
);
NAND #() 
NAND_4464_ (
  .A({ S7751 }),
  .B({ S7753 }),
  .Y({ S7755 })
);
NOR #() 
NOR_2851_ (
  .A({ S7399 }),
  .B({ S7407 }),
  .Y({ S7756 })
);
NAND #() 
NAND_4465_ (
  .A({ S7400 }),
  .B({ S7408 }),
  .Y({ S7757 })
);
NOR #() 
NOR_2852_ (
  .A({ S7755 }),
  .B({ S7757 }),
  .Y({ S7758 })
);
NAND #() 
NAND_4466_ (
  .A({ S7754 }),
  .B({ S7756 }),
  .Y({ S7759 })
);
NOR #() 
NOR_2853_ (
  .A({ S7754 }),
  .B({ S7756 }),
  .Y({ S7760 })
);
NAND #() 
NAND_4467_ (
  .A({ S7755 }),
  .B({ S7757 }),
  .Y({ S7762 })
);
NOR #() 
NOR_2854_ (
  .A({ S7758 }),
  .B({ S7760 }),
  .Y({ S7763 })
);
NAND #() 
NAND_4468_ (
  .A({ S7759 }),
  .B({ S7762 }),
  .Y({ S7764 })
);
NOR #() 
NOR_2855_ (
  .A({ S7743 }),
  .B({ S7764 }),
  .Y({ S7765 })
);
NAND #() 
NAND_4469_ (
  .A({ S7744 }),
  .B({ S7763 }),
  .Y({ S7766 })
);
NOR #() 
NOR_2856_ (
  .A({ S7744 }),
  .B({ S7763 }),
  .Y({ S7767 })
);
NAND #() 
NAND_4470_ (
  .A({ S7743 }),
  .B({ S7764 }),
  .Y({ S7768 })
);
NOR #() 
NOR_2857_ (
  .A({ S7765 }),
  .B({ S7767 }),
  .Y({ S7769 })
);
NAND #() 
NAND_4471_ (
  .A({ S7766 }),
  .B({ S7768 }),
  .Y({ S7770 })
);
NOR #() 
NOR_2858_ (
  .A({ S7413 }),
  .B({ S7421 }),
  .Y({ S7771 })
);
NAND #() 
NAND_4472_ (
  .A({ S7414 }),
  .B({ S7422 }),
  .Y({ S7773 })
);
NOR #() 
NOR_2859_ (
  .A({ S7770 }),
  .B({ S7773 }),
  .Y({ S7774 })
);
NAND #() 
NAND_4473_ (
  .A({ S7769 }),
  .B({ S7771 }),
  .Y({ S7775 })
);
NOR #() 
NOR_2860_ (
  .A({ S7769 }),
  .B({ S7771 }),
  .Y({ S7776 })
);
NAND #() 
NAND_4474_ (
  .A({ S7770 }),
  .B({ S7773 }),
  .Y({ S7777 })
);
NOR #() 
NOR_2861_ (
  .A({ S7774 }),
  .B({ S7776 }),
  .Y({ S7778 })
);
NAND #() 
NAND_4475_ (
  .A({ S7775 }),
  .B({ S7777 }),
  .Y({ S7779 })
);
NOR #() 
NOR_2862_ (
  .A({ S7741 }),
  .B({ S7778 }),
  .Y({ S7780 })
);
NAND #() 
NAND_4476_ (
  .A({ S7742 }),
  .B({ S7779 }),
  .Y({ S7781 })
);
NOR #() 
NOR_2863_ (
  .A({ S7742 }),
  .B({ S7779 }),
  .Y({ S7782 })
);
NAND #() 
NAND_4477_ (
  .A({ S7741 }),
  .B({ S7778 }),
  .Y({ S7784 })
);
NOR #() 
NOR_2864_ (
  .A({ S7780 }),
  .B({ S7782 }),
  .Y({ S7785 })
);
NAND #() 
NAND_4478_ (
  .A({ S7781 }),
  .B({ S7784 }),
  .Y({ S7786 })
);
NOR #() 
NOR_2865_ (
  .A({ S7738 }),
  .B({ S7785 }),
  .Y({ S7787 })
);
NAND #() 
NAND_4479_ (
  .A({ S7740 }),
  .B({ S7786 }),
  .Y({ S7788 })
);
NOR #() 
NOR_2866_ (
  .A({ S7740 }),
  .B({ S7786 }),
  .Y({ S7789 })
);
NAND #() 
NAND_4480_ (
  .A({ S7738 }),
  .B({ S7785 }),
  .Y({ S7790 })
);
NOR #() 
NOR_2867_ (
  .A({ S7787 }),
  .B({ S7789 }),
  .Y({ S7791 })
);
NAND #() 
NAND_4481_ (
  .A({ S7788 }),
  .B({ S7790 }),
  .Y({ S7792 })
);
NOR #() 
NOR_2868_ (
  .A({ S7571 }),
  .B({ S7792 }),
  .Y({ S7793 })
);
NAND #() 
NAND_4482_ (
  .A({ S7572 }),
  .B({ S7791 }),
  .Y({ S7795 })
);
NOR #() 
NOR_2869_ (
  .A({ S7572 }),
  .B({ S7791 }),
  .Y({ S7796 })
);
NAND #() 
NAND_4483_ (
  .A({ S7571 }),
  .B({ S7792 }),
  .Y({ S7797 })
);
NOR #() 
NOR_2870_ (
  .A({ S7793 }),
  .B({ S7796 }),
  .Y({ S7798 })
);
NAND #() 
NAND_4484_ (
  .A({ S7795 }),
  .B({ S7797 }),
  .Y({ S7799 })
);
NAND #() 
NAND_4485_ (
  .A({ S7353 }),
  .B({ S7554 }),
  .Y({ S7800 })
);
NOT #() 
NOT_539_ (
  .A({ S7800 }),
  .Y({ S7801 })
);
NOR #() 
NOR_2871_ (
  .A({ S7353 }),
  .B({ S7554 }),
  .Y({ S7802 })
);
NOT #() 
NOT_540_ (
  .A({ S7802 }),
  .Y({ S7803 })
);
NOR #() 
NOR_2872_ (
  .A({ S7801 }),
  .B({ S7802 }),
  .Y({ S7804 })
);
NAND #() 
NAND_4486_ (
  .A({ S7800 }),
  .B({ S7803 }),
  .Y({ S7806 })
);
NAND #() 
NAND_4487_ (
  .A({ S7798 }),
  .B({ S7806 }),
  .Y({ S7807 })
);
NAND #() 
NAND_4488_ (
  .A({ S7799 }),
  .B({ S7804 }),
  .Y({ S7808 })
);
NAND #() 
NAND_4489_ (
  .A({ S7807 }),
  .B({ S7808 }),
  .Y({ S7809 })
);
NOR #() 
NOR_2873_ (
  .A({ S7570 }),
  .B({ S7809 }),
  .Y({ S7810 })
);
NAND #() 
NAND_4490_ (
  .A({ S7570 }),
  .B({ S7809 }),
  .Y({ S7811 })
);
NOR #() 
NOR_2874_ (
  .A({ S5949 }),
  .B({ S7810 }),
  .Y({ S7812 })
);
NAND #() 
NAND_4491_ (
  .A({ S7811 }),
  .B({ S7812 }),
  .Y({ S7813 })
);
NAND #() 
NAND_4492_ (
  .A({ datapath_multdivunit_outmdu1_15 }),
  .B({ S5950 }),
  .Y({ S7814 })
);
NOT #() 
NOT_541_ (
  .A({ S7814 }),
  .Y({ S7815 })
);
NOR #() 
NOR_2875_ (
  .A({ datapath_addsubunit_in1_15 }),
  .B({ S1516 }),
  .Y({ S7817 })
);
NOR #() 
NOR_2876_ (
  .A({ S3899 }),
  .B({ S7817 }),
  .Y({ S7818 })
);
NOT #() 
NOT_542_ (
  .A({ S7818 }),
  .Y({ S7819 })
);
NOR #() 
NOR_2877_ (
  .A({ S3927 }),
  .B({ S7819 }),
  .Y({ S7820 })
);
NOR #() 
NOR_2878_ (
  .A({ S7815 }),
  .B({ S7820 }),
  .Y({ S7821 })
);
NAND #() 
NAND_4493_ (
  .A({ S7813 }),
  .B({ S7821 }),
  .Y({ S297 })
);
NOR #() 
NOR_2879_ (
  .A({ S8033 }),
  .B({ S1377 }),
  .Y({ S298 })
);
NOR #() 
NOR_2880_ (
  .A({ S8044 }),
  .B({ S1377 }),
  .Y({ S299 })
);
NOR #() 
NOR_2881_ (
  .A({ S8054 }),
  .B({ S1377 }),
  .Y({ S300 })
);
NOR #() 
NOR_2882_ (
  .A({ S8065 }),
  .B({ S1377 }),
  .Y({ S301 })
);
NOR #() 
NOR_2883_ (
  .A({ S8076 }),
  .B({ S1377 }),
  .Y({ S302 })
);
NOR #() 
NOR_2884_ (
  .A({ S8087 }),
  .B({ S1377 }),
  .Y({ S303 })
);
NOR #() 
NOR_2885_ (
  .A({ S8097 }),
  .B({ S1377 }),
  .Y({ S304 })
);
NOR #() 
NOR_2886_ (
  .A({ S8108 }),
  .B({ S1377 }),
  .Y({ S305 })
);
NOR #() 
NOR_2887_ (
  .A({ S8119 }),
  .B({ S1377 }),
  .Y({ S306 })
);
NOR #() 
NOR_2888_ (
  .A({ S8129 }),
  .B({ S1377 }),
  .Y({ S307 })
);
NOR #() 
NOR_2889_ (
  .A({ S8140 }),
  .B({ S1377 }),
  .Y({ S308 })
);
NOR #() 
NOR_2890_ (
  .A({ S8151 }),
  .B({ S1377 }),
  .Y({ S309 })
);
NOR #() 
NOR_2891_ (
  .A({ S8161 }),
  .B({ S1377 }),
  .Y({ S310 })
);
NOR #() 
NOR_2892_ (
  .A({ S8172 }),
  .B({ S1377 }),
  .Y({ S311 })
);
NOR #() 
NOR_2893_ (
  .A({ S8183 }),
  .B({ S1377 }),
  .Y({ S312 })
);
NAND #() 
NAND_4494_ (
  .A({ datapath_databusin_0 }),
  .B({ controller_1115_S_0 }),
  .Y({ S7824 })
);
NAND #() 
NAND_4495_ (
  .A({ datapath_instruction_0 }),
  .B({ S1379 }),
  .Y({ S7825 })
);
NAND #() 
NAND_4496_ (
  .A({ S7824 }),
  .B({ S7825 }),
  .Y({ S313 })
);
NAND #() 
NAND_4497_ (
  .A({ datapath_databusin_1 }),
  .B({ controller_1115_S_0 }),
  .Y({ S7826 })
);
NAND #() 
NAND_4498_ (
  .A({ datapath_instruction_1 }),
  .B({ S1379 }),
  .Y({ S7827 })
);
NAND #() 
NAND_4499_ (
  .A({ S7826 }),
  .B({ S7827 }),
  .Y({ S314 })
);
NAND #() 
NAND_4500_ (
  .A({ datapath_databusin_2 }),
  .B({ controller_1115_S_0 }),
  .Y({ S7828 })
);
NAND #() 
NAND_4501_ (
  .A({ datapath_instruction_2 }),
  .B({ S1379 }),
  .Y({ S7829 })
);
NAND #() 
NAND_4502_ (
  .A({ S7828 }),
  .B({ S7829 }),
  .Y({ S315 })
);
NAND #() 
NAND_4503_ (
  .A({ datapath_databusin_3 }),
  .B({ controller_1115_S_0 }),
  .Y({ S7831 })
);
NAND #() 
NAND_4504_ (
  .A({ datapath_instruction_3 }),
  .B({ S1379 }),
  .Y({ S7832 })
);
NAND #() 
NAND_4505_ (
  .A({ S7831 }),
  .B({ S7832 }),
  .Y({ S316 })
);
NAND #() 
NAND_4506_ (
  .A({ datapath_databusin_4 }),
  .B({ controller_1115_S_0 }),
  .Y({ S7833 })
);
NAND #() 
NAND_4507_ (
  .A({ controller_fib_0 }),
  .B({ S1379 }),
  .Y({ S7834 })
);
NAND #() 
NAND_4508_ (
  .A({ S7833 }),
  .B({ S7834 }),
  .Y({ S317 })
);
NAND #() 
NAND_4509_ (
  .A({ datapath_databusin_5 }),
  .B({ controller_1115_S_0 }),
  .Y({ S7835 })
);
NAND #() 
NAND_4510_ (
  .A({ controller_fib_1 }),
  .B({ S1379 }),
  .Y({ S7836 })
);
NAND #() 
NAND_4511_ (
  .A({ S7835 }),
  .B({ S7836 }),
  .Y({ S318 })
);
NAND #() 
NAND_4512_ (
  .A({ datapath_databusin_6 }),
  .B({ controller_1115_S_0 }),
  .Y({ S7837 })
);
NAND #() 
NAND_4513_ (
  .A({ controller_fib_2 }),
  .B({ S1379 }),
  .Y({ S7839 })
);
NAND #() 
NAND_4514_ (
  .A({ S7837 }),
  .B({ S7839 }),
  .Y({ S319 })
);
NAND #() 
NAND_4515_ (
  .A({ datapath_databusin_7 }),
  .B({ controller_1115_S_0 }),
  .Y({ S7840 })
);
NAND #() 
NAND_4516_ (
  .A({ controller_fib_3 }),
  .B({ S1379 }),
  .Y({ S7841 })
);
NAND #() 
NAND_4517_ (
  .A({ S7840 }),
  .B({ S7841 }),
  .Y({ S320 })
);
NAND #() 
NAND_4518_ (
  .A({ datapath_databusin_8 }),
  .B({ controller_1115_S_0 }),
  .Y({ S7842 })
);
NAND #() 
NAND_4519_ (
  .A({ controller_fib_4 }),
  .B({ S1379 }),
  .Y({ S7843 })
);
NAND #() 
NAND_4520_ (
  .A({ S7842 }),
  .B({ S7843 }),
  .Y({ S321 })
);
NAND #() 
NAND_4521_ (
  .A({ datapath_databusin_9 }),
  .B({ controller_1115_S_0 }),
  .Y({ S7844 })
);
NAND #() 
NAND_4522_ (
  .A({ controller_216_B_0 }),
  .B({ S1379 }),
  .Y({ S7845 })
);
NAND #() 
NAND_4523_ (
  .A({ S7844 }),
  .B({ S7845 }),
  .Y({ S322 })
);
NAND #() 
NAND_4524_ (
  .A({ datapath_databusin_10 }),
  .B({ controller_1115_S_0 }),
  .Y({ S7847 })
);
NAND #() 
NAND_4525_ (
  .A({ controller_opcode_2 }),
  .B({ S1379 }),
  .Y({ S7848 })
);
NAND #() 
NAND_4526_ (
  .A({ S7847 }),
  .B({ S7848 }),
  .Y({ S323 })
);
NAND #() 
NAND_4527_ (
  .A({ datapath_databusin_11 }),
  .B({ controller_1115_S_0 }),
  .Y({ S7849 })
);
NAND #() 
NAND_4528_ (
  .A({ controller_opcode_3 }),
  .B({ S1379 }),
  .Y({ S7850 })
);
NAND #() 
NAND_4529_ (
  .A({ S7849 }),
  .B({ S7850 }),
  .Y({ S324 })
);
NAND #() 
NAND_4530_ (
  .A({ datapath_databusin_12 }),
  .B({ controller_1115_S_0 }),
  .Y({ S7851 })
);
NAND #() 
NAND_4531_ (
  .A({ controller_opcode_4 }),
  .B({ S1379 }),
  .Y({ S7852 })
);
NAND #() 
NAND_4532_ (
  .A({ S7851 }),
  .B({ S7852 }),
  .Y({ S325 })
);
NAND #() 
NAND_4533_ (
  .A({ datapath_databusin_13 }),
  .B({ controller_1115_S_0 }),
  .Y({ S7854 })
);
NAND #() 
NAND_4534_ (
  .A({ controller_opcode_5 }),
  .B({ S1379 }),
  .Y({ S7855 })
);
NAND #() 
NAND_4535_ (
  .A({ S7854 }),
  .B({ S7855 }),
  .Y({ S326 })
);
NAND #() 
NAND_4536_ (
  .A({ datapath_databusin_14 }),
  .B({ controller_1115_S_0 }),
  .Y({ S7856 })
);
NAND #() 
NAND_4537_ (
  .A({ controller_opcode_6 }),
  .B({ S1379 }),
  .Y({ S7857 })
);
NAND #() 
NAND_4538_ (
  .A({ S7856 }),
  .B({ S7857 }),
  .Y({ S327 })
);
NAND #() 
NAND_4539_ (
  .A({ datapath_adr_outreg_0 }),
  .B({ S1383 }),
  .Y({ S7858 })
);
NAND #() 
NAND_4540_ (
  .A({ S1222 }),
  .B({ S1382 }),
  .Y({ S7859 })
);
NAND #() 
NAND_4541_ (
  .A({ S7858 }),
  .B({ S7859 }),
  .Y({ S328 })
);
NAND #() 
NAND_4542_ (
  .A({ datapath_adr_outreg_1 }),
  .B({ S1383 }),
  .Y({ S7860 })
);
NAND #() 
NAND_4543_ (
  .A({ S1170 }),
  .B({ S1382 }),
  .Y({ S7862 })
);
NAND #() 
NAND_4544_ (
  .A({ S7860 }),
  .B({ S7862 }),
  .Y({ S329 })
);
NAND #() 
NAND_4545_ (
  .A({ datapath_adr_outreg_2 }),
  .B({ S1383 }),
  .Y({ S7863 })
);
NAND #() 
NAND_4546_ (
  .A({ S1118 }),
  .B({ S1382 }),
  .Y({ S7864 })
);
NAND #() 
NAND_4547_ (
  .A({ S7863 }),
  .B({ S7864 }),
  .Y({ S330 })
);
NAND #() 
NAND_4548_ (
  .A({ datapath_adr_outreg_3 }),
  .B({ S1383 }),
  .Y({ S7865 })
);
NAND #() 
NAND_4549_ (
  .A({ S1067 }),
  .B({ S1382 }),
  .Y({ S7866 })
);
NAND #() 
NAND_4550_ (
  .A({ S7865 }),
  .B({ S7866 }),
  .Y({ S331 })
);
NAND #() 
NAND_4551_ (
  .A({ datapath_adr_outreg_4 }),
  .B({ S1383 }),
  .Y({ S7867 })
);
NAND #() 
NAND_4552_ (
  .A({ S1015 }),
  .B({ S1382 }),
  .Y({ S7868 })
);
NAND #() 
NAND_4553_ (
  .A({ S7867 }),
  .B({ S7868 }),
  .Y({ S332 })
);
NAND #() 
NAND_4554_ (
  .A({ datapath_adr_outreg_5 }),
  .B({ S1383 }),
  .Y({ S7870 })
);
NAND #() 
NAND_4555_ (
  .A({ S965 }),
  .B({ S1382 }),
  .Y({ S7871 })
);
NAND #() 
NAND_4556_ (
  .A({ S7870 }),
  .B({ S7871 }),
  .Y({ S333 })
);
NAND #() 
NAND_4557_ (
  .A({ datapath_adr_outreg_6 }),
  .B({ S1383 }),
  .Y({ S7872 })
);
NAND #() 
NAND_4558_ (
  .A({ S912 }),
  .B({ S1382 }),
  .Y({ S7873 })
);
NAND #() 
NAND_4559_ (
  .A({ S7872 }),
  .B({ S7873 }),
  .Y({ S334 })
);
NAND #() 
NAND_4560_ (
  .A({ datapath_adr_outreg_7 }),
  .B({ S1383 }),
  .Y({ S7874 })
);
NAND #() 
NAND_4561_ (
  .A({ S860 }),
  .B({ S1382 }),
  .Y({ S7875 })
);
NAND #() 
NAND_4562_ (
  .A({ S7874 }),
  .B({ S7875 }),
  .Y({ S335 })
);
NAND #() 
NAND_4563_ (
  .A({ datapath_adr_outreg_8 }),
  .B({ S1383 }),
  .Y({ S7877 })
);
NAND #() 
NAND_4564_ (
  .A({ S807 }),
  .B({ S1382 }),
  .Y({ S7878 })
);
NAND #() 
NAND_4565_ (
  .A({ S7877 }),
  .B({ S7878 }),
  .Y({ S336 })
);
NAND #() 
NAND_4566_ (
  .A({ datapath_adr_outreg_9 }),
  .B({ S1383 }),
  .Y({ S7879 })
);
NAND #() 
NAND_4567_ (
  .A({ S756 }),
  .B({ S1382 }),
  .Y({ S7880 })
);
NAND #() 
NAND_4568_ (
  .A({ S7879 }),
  .B({ S7880 }),
  .Y({ S337 })
);
NAND #() 
NAND_4569_ (
  .A({ datapath_adr_outreg_10 }),
  .B({ S1383 }),
  .Y({ S7881 })
);
NAND #() 
NAND_4570_ (
  .A({ S704 }),
  .B({ S1382 }),
  .Y({ S7882 })
);
NAND #() 
NAND_4571_ (
  .A({ S7881 }),
  .B({ S7882 }),
  .Y({ S338 })
);
NAND #() 
NAND_4572_ (
  .A({ datapath_adr_outreg_11 }),
  .B({ S1383 }),
  .Y({ S7883 })
);
NAND #() 
NAND_4573_ (
  .A({ S653 }),
  .B({ S1382 }),
  .Y({ S7885 })
);
NAND #() 
NAND_4574_ (
  .A({ S7883 }),
  .B({ S7885 }),
  .Y({ S339 })
);
NAND #() 
NAND_4575_ (
  .A({ datapath_adr_outreg_12 }),
  .B({ S1383 }),
  .Y({ S7886 })
);
NAND #() 
NAND_4576_ (
  .A({ S601 }),
  .B({ S1382 }),
  .Y({ S7887 })
);
NAND #() 
NAND_4577_ (
  .A({ S7886 }),
  .B({ S7887 }),
  .Y({ S340 })
);
NAND #() 
NAND_4578_ (
  .A({ datapath_adr_outreg_13 }),
  .B({ S1383 }),
  .Y({ S7888 })
);
NAND #() 
NAND_4579_ (
  .A({ S550 }),
  .B({ S1382 }),
  .Y({ S7889 })
);
NAND #() 
NAND_4580_ (
  .A({ S7888 }),
  .B({ S7889 }),
  .Y({ S341 })
);
NAND #() 
NAND_4581_ (
  .A({ datapath_adr_outreg_14 }),
  .B({ S1383 }),
  .Y({ S7890 })
);
NAND #() 
NAND_4582_ (
  .A({ S498 }),
  .B({ S1382 }),
  .Y({ S7891 })
);
NAND #() 
NAND_4583_ (
  .A({ S7890 }),
  .B({ S7891 }),
  .Y({ S342 })
);
NOR #() 
NOR_2894_ (
  .A({ controller_216_B_0 }),
  .B({ S1628 }),
  .Y({ controller_readmem })
);
NOR #() 
NOR_2895_ (
  .A({ controller_216_B_0 }),
  .B({ S403 }),
  .Y({ controller_writemem })
);
NAND #() 
NAND_4584_ (
  .A({ controller_216_B_0 }),
  .B({ S1627 }),
  .Y({ S7893 })
);
NOT #() 
NOT_543_ (
  .A({ S7893 }),
  .Y({ controller_readio })
);
NOR #() 
NOR_2896_ (
  .A({ S8278 }),
  .B({ S403 }),
  .Y({ controller_writeio })
);
NOR #() 
NOR_2897_ (
  .A({ S1377 }),
  .B({ controller_1115_S_0 }),
  .Y({ S7894 })
);
NOT #() 
NOT_544_ (
  .A({ S7894 }),
  .Y({ controller_1405_Y_0 })
);
NAND #() 
NAND_4585_ (
  .A({ S8572 }),
  .B({ S8576 }),
  .Y({ S7895 })
);
NOT #() 
NOT_545_ (
  .A({ S7895 }),
  .Y({ S7896 })
);
NAND #() 
NAND_4586_ (
  .A({ S1383 }),
  .B({ S5950 }),
  .Y({ S7898 })
);
NOR #() 
NOR_2898_ (
  .A({ S7896 }),
  .B({ S7898 }),
  .Y({ S7899 })
);
NAND #() 
NAND_4587_ (
  .A({ S1378 }),
  .B({ S7899 }),
  .Y({ controller_1405_Y_1 })
);
NAND #() 
NAND_4588_ (
  .A({ datapath_muxmem_in2_0 }),
  .B({ controller_1115_S_0 }),
  .Y({ S7900 })
);
NAND #() 
NAND_4589_ (
  .A({ datapath_adr_outreg_0 }),
  .B({ S8576 }),
  .Y({ S7901 })
);
NAND #() 
NAND_4590_ (
  .A({ S7900 }),
  .B({ S7901 }),
  .Y({ datapath_addrbus_0 })
);
NAND #() 
NAND_4591_ (
  .A({ datapath_muxmem_in2_1 }),
  .B({ controller_1115_S_0 }),
  .Y({ S7902 })
);
NAND #() 
NAND_4592_ (
  .A({ datapath_adr_outreg_1 }),
  .B({ S8576 }),
  .Y({ S7903 })
);
NAND #() 
NAND_4593_ (
  .A({ S7902 }),
  .B({ S7903 }),
  .Y({ datapath_addrbus_1 })
);
NAND #() 
NAND_4594_ (
  .A({ datapath_muxmem_in2_2 }),
  .B({ controller_1115_S_0 }),
  .Y({ S7904 })
);
NAND #() 
NAND_4595_ (
  .A({ datapath_adr_outreg_2 }),
  .B({ S8576 }),
  .Y({ S7906 })
);
NAND #() 
NAND_4596_ (
  .A({ S7904 }),
  .B({ S7906 }),
  .Y({ datapath_addrbus_2 })
);
NAND #() 
NAND_4597_ (
  .A({ datapath_muxmem_in2_3 }),
  .B({ controller_1115_S_0 }),
  .Y({ S7907 })
);
NAND #() 
NAND_4598_ (
  .A({ datapath_adr_outreg_3 }),
  .B({ S8576 }),
  .Y({ S7908 })
);
NAND #() 
NAND_4599_ (
  .A({ S7907 }),
  .B({ S7908 }),
  .Y({ datapath_addrbus_3 })
);
NAND #() 
NAND_4600_ (
  .A({ datapath_muxmem_in2_4 }),
  .B({ controller_1115_S_0 }),
  .Y({ S7909 })
);
NAND #() 
NAND_4601_ (
  .A({ datapath_adr_outreg_4 }),
  .B({ S8576 }),
  .Y({ S7910 })
);
NAND #() 
NAND_4602_ (
  .A({ S7909 }),
  .B({ S7910 }),
  .Y({ datapath_addrbus_4 })
);
NAND #() 
NAND_4603_ (
  .A({ datapath_muxmem_in2_5 }),
  .B({ controller_1115_S_0 }),
  .Y({ S7911 })
);
NAND #() 
NAND_4604_ (
  .A({ datapath_adr_outreg_5 }),
  .B({ S8576 }),
  .Y({ S7912 })
);
NAND #() 
NAND_4605_ (
  .A({ S7911 }),
  .B({ S7912 }),
  .Y({ datapath_addrbus_5 })
);
NAND #() 
NAND_4606_ (
  .A({ datapath_muxmem_in2_6 }),
  .B({ controller_1115_S_0 }),
  .Y({ S7914 })
);
NAND #() 
NAND_4607_ (
  .A({ datapath_adr_outreg_6 }),
  .B({ S8576 }),
  .Y({ S7915 })
);
NAND #() 
NAND_4608_ (
  .A({ S7914 }),
  .B({ S7915 }),
  .Y({ datapath_addrbus_6 })
);
NAND #() 
NAND_4609_ (
  .A({ datapath_muxmem_in2_7 }),
  .B({ controller_1115_S_0 }),
  .Y({ S7916 })
);
NAND #() 
NAND_4610_ (
  .A({ datapath_adr_outreg_7 }),
  .B({ S8576 }),
  .Y({ S7917 })
);
NAND #() 
NAND_4611_ (
  .A({ S7916 }),
  .B({ S7917 }),
  .Y({ datapath_addrbus_7 })
);
NAND #() 
NAND_4612_ (
  .A({ datapath_muxmem_in2_8 }),
  .B({ controller_1115_S_0 }),
  .Y({ S7918 })
);
NAND #() 
NAND_4613_ (
  .A({ datapath_adr_outreg_8 }),
  .B({ S8576 }),
  .Y({ S7919 })
);
NAND #() 
NAND_4614_ (
  .A({ S7918 }),
  .B({ S7919 }),
  .Y({ datapath_addrbus_8 })
);
NAND #() 
NAND_4615_ (
  .A({ datapath_muxmem_in2_9 }),
  .B({ controller_1115_S_0 }),
  .Y({ S7921 })
);
NAND #() 
NAND_4616_ (
  .A({ datapath_adr_outreg_9 }),
  .B({ S8576 }),
  .Y({ S7922 })
);
NAND #() 
NAND_4617_ (
  .A({ S7921 }),
  .B({ S7922 }),
  .Y({ datapath_addrbus_9 })
);
NAND #() 
NAND_4618_ (
  .A({ datapath_muxmem_in2_10 }),
  .B({ controller_1115_S_0 }),
  .Y({ S7923 })
);
NAND #() 
NAND_4619_ (
  .A({ datapath_adr_outreg_10 }),
  .B({ S8576 }),
  .Y({ S7924 })
);
NAND #() 
NAND_4620_ (
  .A({ S7923 }),
  .B({ S7924 }),
  .Y({ datapath_addrbus_10 })
);
NAND #() 
NAND_4621_ (
  .A({ datapath_muxmem_in2_11 }),
  .B({ controller_1115_S_0 }),
  .Y({ S7925 })
);
NAND #() 
NAND_4622_ (
  .A({ datapath_adr_outreg_11 }),
  .B({ S8576 }),
  .Y({ S7926 })
);
NAND #() 
NAND_4623_ (
  .A({ S7925 }),
  .B({ S7926 }),
  .Y({ datapath_addrbus_11 })
);
NAND #() 
NAND_4624_ (
  .A({ datapath_muxmem_in2_12 }),
  .B({ controller_1115_S_0 }),
  .Y({ S7927 })
);
NAND #() 
NAND_4625_ (
  .A({ datapath_adr_outreg_12 }),
  .B({ S8576 }),
  .Y({ S7929 })
);
NAND #() 
NAND_4626_ (
  .A({ S7927 }),
  .B({ S7929 }),
  .Y({ datapath_addrbus_12 })
);
NAND #() 
NAND_4627_ (
  .A({ datapath_muxmem_in2_13 }),
  .B({ controller_1115_S_0 }),
  .Y({ S7930 })
);
NAND #() 
NAND_4628_ (
  .A({ datapath_adr_outreg_13 }),
  .B({ S8576 }),
  .Y({ S7931 })
);
NAND #() 
NAND_4629_ (
  .A({ S7930 }),
  .B({ S7931 }),
  .Y({ datapath_addrbus_13 })
);
NAND #() 
NAND_4630_ (
  .A({ datapath_muxmem_in2_14 }),
  .B({ controller_1115_S_0 }),
  .Y({ S7932 })
);
NAND #() 
NAND_4631_ (
  .A({ datapath_adr_outreg_14 }),
  .B({ S8576 }),
  .Y({ S7933 })
);
NAND #() 
NAND_4632_ (
  .A({ S7932 }),
  .B({ S7933 }),
  .Y({ datapath_addrbus_14 })
);
NAND #() 
NAND_4633_ (
  .A({ datapath_muxmem_in2_15 }),
  .B({ controller_1115_S_0 }),
  .Y({ S7934 })
);
NAND #() 
NAND_4634_ (
  .A({ datapath_adr_outreg_15 }),
  .B({ S8576 }),
  .Y({ S7935 })
);
NAND #() 
NAND_4635_ (
  .A({ S7934 }),
  .B({ S7935 }),
  .Y({ datapath_addrbus_15 })
);
NOR #() 
NOR_2899_ (
  .A({ S1604 }),
  .B({ S1746 }),
  .Y({ S7937 })
);
NAND #() 
NAND_4636_ (
  .A({ S1605 }),
  .B({ S1745 }),
  .Y({ S7938 })
);
NAND #() 
NAND_4637_ (
  .A({ controller_fib_1 }),
  .B({ S1607 }),
  .Y({ S7939 })
);
NOT #() 
NOT_546_ (
  .A({ S7939 }),
  .Y({ S7940 })
);
NOR #() 
NOR_2900_ (
  .A({ S7937 }),
  .B({ S7940 }),
  .Y({ S7941 })
);
NAND #() 
NAND_4638_ (
  .A({ S7938 }),
  .B({ S7939 }),
  .Y({ S7942 })
);
NOR #() 
NOR_2901_ (
  .A({ S1516 }),
  .B({ S1604 }),
  .Y({ S7943 })
);
NAND #() 
NAND_4639_ (
  .A({ S1515 }),
  .B({ S1605 }),
  .Y({ S7944 })
);
NAND #() 
NAND_4640_ (
  .A({ controller_fib_0 }),
  .B({ S1607 }),
  .Y({ S7945 })
);
NOT #() 
NOT_547_ (
  .A({ S7945 }),
  .Y({ S7947 })
);
NOR #() 
NOR_2902_ (
  .A({ S7943 }),
  .B({ S7947 }),
  .Y({ S7948 })
);
NAND #() 
NAND_4641_ (
  .A({ S7944 }),
  .B({ S7945 }),
  .Y({ S7949 })
);
NOR #() 
NOR_2903_ (
  .A({ S7942 }),
  .B({ S7949 }),
  .Y({ S7950 })
);
NAND #() 
NAND_4642_ (
  .A({ S7941 }),
  .B({ S7948 }),
  .Y({ S7951 })
);
NOR #() 
NOR_2904_ (
  .A({ S1604 }),
  .B({ S1953 }),
  .Y({ S7952 })
);
NAND #() 
NAND_4643_ (
  .A({ S1605 }),
  .B({ S1952 }),
  .Y({ S7953 })
);
NAND #() 
NAND_4644_ (
  .A({ controller_fib_3 }),
  .B({ S1607 }),
  .Y({ S7954 })
);
NOT #() 
NOT_548_ (
  .A({ S7954 }),
  .Y({ S7955 })
);
NOR #() 
NOR_2905_ (
  .A({ S7952 }),
  .B({ S7955 }),
  .Y({ S7956 })
);
NAND #() 
NAND_4645_ (
  .A({ S7953 }),
  .B({ S7954 }),
  .Y({ S7958 })
);
NOR #() 
NOR_2906_ (
  .A({ S1604 }),
  .B({ S1849 }),
  .Y({ S7959 })
);
NAND #() 
NAND_4646_ (
  .A({ S1605 }),
  .B({ S1848 }),
  .Y({ S7960 })
);
NAND #() 
NAND_4647_ (
  .A({ controller_fib_2 }),
  .B({ S1607 }),
  .Y({ S7961 })
);
NOT #() 
NOT_549_ (
  .A({ S7961 }),
  .Y({ S7962 })
);
NOR #() 
NOR_2907_ (
  .A({ S7959 }),
  .B({ S7962 }),
  .Y({ S7963 })
);
NAND #() 
NAND_4648_ (
  .A({ S7960 }),
  .B({ S7961 }),
  .Y({ S7964 })
);
NOR #() 
NOR_2908_ (
  .A({ S7958 }),
  .B({ S7964 }),
  .Y({ S7965 })
);
NAND #() 
NAND_4649_ (
  .A({ S7956 }),
  .B({ S7963 }),
  .Y({ S7966 })
);
NOR #() 
NOR_2909_ (
  .A({ S7951 }),
  .B({ S7966 }),
  .Y({ S7967 })
);
NAND #() 
NAND_4650_ (
  .A({ S7950 }),
  .B({ S7965 }),
  .Y({ S7969 })
);
NAND #() 
NAND_4651_ (
  .A({ datapath_addsubunit_in1_0 }),
  .B({ S7967 }),
  .Y({ S7970 })
);
NOT #() 
NOT_550_ (
  .A({ S7970 }),
  .Y({ datapath_shiftunit_2439_A })
);
NOR #() 
NOR_2910_ (
  .A({ S7941 }),
  .B({ S7948 }),
  .Y({ S7971 })
);
NAND #() 
NAND_4652_ (
  .A({ S7942 }),
  .B({ S7949 }),
  .Y({ S7972 })
);
NOR #() 
NOR_2911_ (
  .A({ S7966 }),
  .B({ S7972 }),
  .Y({ S7973 })
);
NAND #() 
NAND_4653_ (
  .A({ S7965 }),
  .B({ S7971 }),
  .Y({ S7974 })
);
NAND #() 
NAND_4654_ (
  .A({ datapath_addsubunit_in1_3 }),
  .B({ S7973 }),
  .Y({ S7975 })
);
NOR #() 
NOR_2912_ (
  .A({ S7956 }),
  .B({ S7964 }),
  .Y({ S7976 })
);
NAND #() 
NAND_4655_ (
  .A({ S7958 }),
  .B({ S7963 }),
  .Y({ S7977 })
);
NOR #() 
NOR_2913_ (
  .A({ S7941 }),
  .B({ S7949 }),
  .Y({ S7979 })
);
NAND #() 
NAND_4656_ (
  .A({ S7942 }),
  .B({ S7948 }),
  .Y({ S7980 })
);
NAND #() 
NAND_4657_ (
  .A({ S7976 }),
  .B({ S7979 }),
  .Y({ S7981 })
);
NOT #() 
NOT_551_ (
  .A({ S7981 }),
  .Y({ S7982 })
);
NAND #() 
NAND_4658_ (
  .A({ datapath_addsubunit_in1_10 }),
  .B({ S7982 }),
  .Y({ S7983 })
);
NOR #() 
NOR_2914_ (
  .A({ S7951 }),
  .B({ S7977 }),
  .Y({ S7984 })
);
NAND #() 
NAND_4659_ (
  .A({ S7950 }),
  .B({ S7976 }),
  .Y({ S7985 })
);
NAND #() 
NAND_4660_ (
  .A({ datapath_addsubunit_in1_8 }),
  .B({ S7984 }),
  .Y({ S7986 })
);
NOR #() 
NOR_2915_ (
  .A({ S7942 }),
  .B({ S7948 }),
  .Y({ S7987 })
);
NAND #() 
NAND_4661_ (
  .A({ S7941 }),
  .B({ S7949 }),
  .Y({ S7988 })
);
NOR #() 
NOR_2916_ (
  .A({ S7956 }),
  .B({ S7963 }),
  .Y({ S7990 })
);
NAND #() 
NAND_4662_ (
  .A({ S7958 }),
  .B({ S7964 }),
  .Y({ S7991 })
);
NAND #() 
NAND_4663_ (
  .A({ S7987 }),
  .B({ S7990 }),
  .Y({ S7992 })
);
NOT #() 
NOT_552_ (
  .A({ S7992 }),
  .Y({ S7993 })
);
NAND #() 
NAND_4664_ (
  .A({ datapath_addsubunit_in1_13 }),
  .B({ S7993 }),
  .Y({ S7994 })
);
NOR #() 
NOR_2917_ (
  .A({ S7951 }),
  .B({ S7991 }),
  .Y({ S7995 })
);
NAND #() 
NAND_4665_ (
  .A({ S7950 }),
  .B({ S7990 }),
  .Y({ S7996 })
);
NAND #() 
NAND_4666_ (
  .A({ datapath_addsubunit_in1_12 }),
  .B({ S7995 }),
  .Y({ S7997 })
);
NAND #() 
NAND_4667_ (
  .A({ S7994 }),
  .B({ S7997 }),
  .Y({ S7998 })
);
NOR #() 
NOR_2918_ (
  .A({ S7958 }),
  .B({ S7963 }),
  .Y({ S7999 })
);
NAND #() 
NAND_4668_ (
  .A({ S7956 }),
  .B({ S7964 }),
  .Y({ S8001 })
);
NOR #() 
NOR_2919_ (
  .A({ S7951 }),
  .B({ S8001 }),
  .Y({ S8002 })
);
NAND #() 
NAND_4669_ (
  .A({ S7950 }),
  .B({ S7999 }),
  .Y({ S8003 })
);
NOR #() 
NOR_2920_ (
  .A({ S1013 }),
  .B({ S8003 }),
  .Y({ S8004 })
);
NAND #() 
NAND_4670_ (
  .A({ datapath_addsubunit_in1_4 }),
  .B({ S8002 }),
  .Y({ S8005 })
);
NOR #() 
NOR_2921_ (
  .A({ S7972 }),
  .B({ S7977 }),
  .Y({ S8006 })
);
NAND #() 
NAND_4671_ (
  .A({ S7971 }),
  .B({ S7976 }),
  .Y({ S8007 })
);
NAND #() 
NAND_4672_ (
  .A({ datapath_addsubunit_in1_11 }),
  .B({ S8006 }),
  .Y({ S8008 })
);
NOR #() 
NOR_2922_ (
  .A({ S7966 }),
  .B({ S7988 }),
  .Y({ S8009 })
);
NAND #() 
NAND_4673_ (
  .A({ S7965 }),
  .B({ S7987 }),
  .Y({ S8010 })
);
NOR #() 
NOR_2923_ (
  .A({ S1168 }),
  .B({ S8010 }),
  .Y({ S8012 })
);
NAND #() 
NAND_4674_ (
  .A({ datapath_addsubunit_in1_1 }),
  .B({ S8009 }),
  .Y({ S8013 })
);
NOR #() 
NOR_2924_ (
  .A({ S7966 }),
  .B({ S7980 }),
  .Y({ S8014 })
);
NAND #() 
NAND_4675_ (
  .A({ S7965 }),
  .B({ S7979 }),
  .Y({ S8015 })
);
NAND #() 
NAND_4676_ (
  .A({ datapath_addsubunit_in1_2 }),
  .B({ S8014 }),
  .Y({ S8016 })
);
NOR #() 
NOR_2925_ (
  .A({ S7980 }),
  .B({ S8001 }),
  .Y({ S8017 })
);
NAND #() 
NAND_4677_ (
  .A({ S7979 }),
  .B({ S7999 }),
  .Y({ S8018 })
);
NOR #() 
NOR_2926_ (
  .A({ S910 }),
  .B({ S8018 }),
  .Y({ S8019 })
);
NOR #() 
NOR_2927_ (
  .A({ S7977 }),
  .B({ S7988 }),
  .Y({ S8020 })
);
NAND #() 
NAND_4678_ (
  .A({ S7976 }),
  .B({ S7987 }),
  .Y({ S8021 })
);
NAND #() 
NAND_4679_ (
  .A({ datapath_addsubunit_in1_9 }),
  .B({ S8020 }),
  .Y({ S8023 })
);
NOR #() 
NOR_2928_ (
  .A({ S7988 }),
  .B({ S8001 }),
  .Y({ S8024 })
);
NAND #() 
NAND_4680_ (
  .A({ S7987 }),
  .B({ S7999 }),
  .Y({ S8025 })
);
NOR #() 
NOR_2929_ (
  .A({ S963 }),
  .B({ S8025 }),
  .Y({ S8026 })
);
NOR #() 
NOR_2930_ (
  .A({ S7980 }),
  .B({ S7991 }),
  .Y({ S8027 })
);
NAND #() 
NAND_4681_ (
  .A({ datapath_addsubunit_in1_14 }),
  .B({ S8027 }),
  .Y({ S8028 })
);
NAND #() 
NAND_4682_ (
  .A({ S7964 }),
  .B({ S7971 }),
  .Y({ S8029 })
);
NOR #() 
NOR_2931_ (
  .A({ S7972 }),
  .B({ S8001 }),
  .Y({ S8030 })
);
NAND #() 
NAND_4683_ (
  .A({ S7971 }),
  .B({ S7999 }),
  .Y({ S8031 })
);
NOR #() 
NOR_2932_ (
  .A({ S858 }),
  .B({ S8031 }),
  .Y({ S8032 })
);
NAND #() 
NAND_4684_ (
  .A({ datapath_addsubunit_in1_7 }),
  .B({ S8030 }),
  .Y({ S8034 })
);
NOR #() 
NOR_2933_ (
  .A({ S7956 }),
  .B({ S8029 }),
  .Y({ S8035 })
);
NAND #() 
NAND_4685_ (
  .A({ datapath_addsubunit_in1_15 }),
  .B({ S8035 }),
  .Y({ S8036 })
);
NOR #() 
NOR_2934_ (
  .A({ S8004 }),
  .B({ S8032 }),
  .Y({ S8037 })
);
NAND #() 
NAND_4686_ (
  .A({ S7971 }),
  .B({ S7990 }),
  .Y({ S8038 })
);
NAND #() 
NAND_4687_ (
  .A({ S7986 }),
  .B({ S8023 }),
  .Y({ S8039 })
);
NAND #() 
NAND_4688_ (
  .A({ S7970 }),
  .B({ S8013 }),
  .Y({ S8040 })
);
NAND #() 
NAND_4689_ (
  .A({ S7975 }),
  .B({ S8016 }),
  .Y({ S8041 })
);
NOR #() 
NOR_2935_ (
  .A({ S8040 }),
  .B({ S8041 }),
  .Y({ S8042 })
);
NAND #() 
NAND_4690_ (
  .A({ S7983 }),
  .B({ S8042 }),
  .Y({ S8043 })
);
NOR #() 
NOR_2936_ (
  .A({ S7998 }),
  .B({ S8043 }),
  .Y({ S8045 })
);
NOR #() 
NOR_2937_ (
  .A({ S8019 }),
  .B({ S8026 }),
  .Y({ S8046 })
);
NAND #() 
NAND_4691_ (
  .A({ S8037 }),
  .B({ S8046 }),
  .Y({ S8047 })
);
NAND #() 
NAND_4692_ (
  .A({ S8008 }),
  .B({ S8028 }),
  .Y({ S8048 })
);
NOR #() 
NOR_2938_ (
  .A({ S8039 }),
  .B({ S8048 }),
  .Y({ S8049 })
);
NAND #() 
NAND_4693_ (
  .A({ S8036 }),
  .B({ S8049 }),
  .Y({ S8050 })
);
NOR #() 
NOR_2939_ (
  .A({ S8047 }),
  .B({ S8050 }),
  .Y({ S8051 })
);
NAND #() 
NAND_4694_ (
  .A({ S8045 }),
  .B({ S8051 }),
  .Y({ datapath_shiftunit_2135_A })
);
NOR #() 
NOR_2940_ (
  .A({ S910 }),
  .B({ S8025 }),
  .Y({ S8052 })
);
NAND #() 
NAND_4695_ (
  .A({ datapath_addsubunit_in1_6 }),
  .B({ S8024 }),
  .Y({ S8053 })
);
NOR #() 
NOR_2941_ (
  .A({ S1116 }),
  .B({ S8010 }),
  .Y({ S8055 })
);
NAND #() 
NAND_4696_ (
  .A({ datapath_addsubunit_in1_2 }),
  .B({ S8009 }),
  .Y({ S8056 })
);
NOR #() 
NOR_2942_ (
  .A({ S548 }),
  .B({ S7996 }),
  .Y({ S8057 })
);
NAND #() 
NAND_4697_ (
  .A({ datapath_addsubunit_in1_5 }),
  .B({ S8002 }),
  .Y({ S8058 })
);
NAND #() 
NAND_4698_ (
  .A({ datapath_addsubunit_in1_9 }),
  .B({ S7984 }),
  .Y({ S8059 })
);
NAND #() 
NAND_4699_ (
  .A({ datapath_addsubunit_in1_3 }),
  .B({ S8014 }),
  .Y({ S8060 })
);
NOR #() 
NOR_2943_ (
  .A({ S858 }),
  .B({ S8018 }),
  .Y({ S8061 })
);
NAND #() 
NAND_4700_ (
  .A({ datapath_addsubunit_in1_10 }),
  .B({ S8020 }),
  .Y({ S8062 })
);
NOR #() 
NOR_2944_ (
  .A({ S1013 }),
  .B({ S7974 }),
  .Y({ S8063 })
);
NAND #() 
NAND_4701_ (
  .A({ datapath_addsubunit_in1_4 }),
  .B({ S7973 }),
  .Y({ S8064 })
);
NAND #() 
NAND_4702_ (
  .A({ datapath_addsubunit_in1_11 }),
  .B({ S7982 }),
  .Y({ S8066 })
);
NAND #() 
NAND_4703_ (
  .A({ datapath_addsubunit_in1_1 }),
  .B({ S7967 }),
  .Y({ S8067 })
);
NAND #() 
NAND_4704_ (
  .A({ datapath_addsubunit_in1_12 }),
  .B({ S8006 }),
  .Y({ S8068 })
);
NAND #() 
NAND_4705_ (
  .A({ datapath_addsubunit_in1_14 }),
  .B({ S7993 }),
  .Y({ S8069 })
);
NAND #() 
NAND_4706_ (
  .A({ datapath_addsubunit_in1_8 }),
  .B({ S8030 }),
  .Y({ S8070 })
);
NAND #() 
NAND_4707_ (
  .A({ datapath_addsubunit_in1_15 }),
  .B({ S8027 }),
  .Y({ S8071 })
);
NAND #() 
NAND_4708_ (
  .A({ S8062 }),
  .B({ S8070 }),
  .Y({ S8072 })
);
NAND #() 
NAND_4709_ (
  .A({ S8056 }),
  .B({ S8069 }),
  .Y({ S8073 })
);
NOR #() 
NOR_2945_ (
  .A({ S8072 }),
  .B({ S8073 }),
  .Y({ S8074 })
);
NOR #() 
NOR_2946_ (
  .A({ S8052 }),
  .B({ S8057 }),
  .Y({ S8075 })
);
NAND #() 
NAND_4710_ (
  .A({ S8058 }),
  .B({ S8059 }),
  .Y({ S8077 })
);
NOR #() 
NOR_2947_ (
  .A({ S1304 }),
  .B({ S1612 }),
  .Y({ S8078 })
);
NAND #() 
NAND_4711_ (
  .A({ datapath_addsubunit_in1_15 }),
  .B({ S1611 }),
  .Y({ S8079 })
);
NOR #() 
NOR_2948_ (
  .A({ S8038 }),
  .B({ S8079 }),
  .Y({ S8080 })
);
NOR #() 
NOR_2949_ (
  .A({ S8077 }),
  .B({ S8080 }),
  .Y({ S8081 })
);
NAND #() 
NAND_4712_ (
  .A({ S8075 }),
  .B({ S8081 }),
  .Y({ S8082 })
);
NAND #() 
NAND_4713_ (
  .A({ S8068 }),
  .B({ S8071 }),
  .Y({ S8083 })
);
NOR #() 
NOR_2950_ (
  .A({ S8061 }),
  .B({ S8083 }),
  .Y({ S8084 })
);
NAND #() 
NAND_4714_ (
  .A({ S8060 }),
  .B({ S8067 }),
  .Y({ S8085 })
);
NAND #() 
NAND_4715_ (
  .A({ S8064 }),
  .B({ S8066 }),
  .Y({ S8086 })
);
NOR #() 
NOR_2951_ (
  .A({ S8085 }),
  .B({ S8086 }),
  .Y({ S8088 })
);
NAND #() 
NAND_4716_ (
  .A({ S8084 }),
  .B({ S8088 }),
  .Y({ S8089 })
);
NOR #() 
NOR_2952_ (
  .A({ S8082 }),
  .B({ S8089 }),
  .Y({ S8090 })
);
NAND #() 
NAND_4717_ (
  .A({ S8074 }),
  .B({ S8090 }),
  .Y({ datapath_shiftunit_2153_A })
);
NAND #() 
NAND_4718_ (
  .A({ datapath_addsubunit_in1_4 }),
  .B({ S8014 }),
  .Y({ S8091 })
);
NAND #() 
NAND_4719_ (
  .A({ datapath_addsubunit_in1_5 }),
  .B({ S7973 }),
  .Y({ S8092 })
);
NAND #() 
NAND_4720_ (
  .A({ S8091 }),
  .B({ S8092 }),
  .Y({ S8093 })
);
NOR #() 
NOR_2953_ (
  .A({ S599 }),
  .B({ S7981 }),
  .Y({ S8094 })
);
NOR #() 
NOR_2954_ (
  .A({ S1304 }),
  .B({ S7992 }),
  .Y({ S8095 })
);
NOR #() 
NOR_2955_ (
  .A({ S8094 }),
  .B({ S8095 }),
  .Y({ S8096 })
);
NOR #() 
NOR_2956_ (
  .A({ S858 }),
  .B({ S8025 }),
  .Y({ S8098 })
);
NOR #() 
NOR_2957_ (
  .A({ S548 }),
  .B({ S8007 }),
  .Y({ S8099 })
);
NOR #() 
NOR_2958_ (
  .A({ S8098 }),
  .B({ S8099 }),
  .Y({ S8100 })
);
NAND #() 
NAND_4721_ (
  .A({ S8096 }),
  .B({ S8100 }),
  .Y({ S8101 })
);
NOR #() 
NOR_2959_ (
  .A({ S8093 }),
  .B({ S8101 }),
  .Y({ S8102 })
);
NOR #() 
NOR_2960_ (
  .A({ S7941 }),
  .B({ S8079 }),
  .Y({ S8103 })
);
NAND #() 
NAND_4722_ (
  .A({ S7942 }),
  .B({ S8078 }),
  .Y({ S8104 })
);
NOR #() 
NOR_2961_ (
  .A({ S7991 }),
  .B({ S8104 }),
  .Y({ S8105 })
);
NOR #() 
NOR_2962_ (
  .A({ S805 }),
  .B({ S8018 }),
  .Y({ S8106 })
);
NAND #() 
NAND_4723_ (
  .A({ datapath_addsubunit_in1_8 }),
  .B({ S8017 }),
  .Y({ S8107 })
);
NOR #() 
NOR_2963_ (
  .A({ S910 }),
  .B({ S8003 }),
  .Y({ S8109 })
);
NAND #() 
NAND_4724_ (
  .A({ datapath_addsubunit_in1_6 }),
  .B({ S8002 }),
  .Y({ S8110 })
);
NAND #() 
NAND_4725_ (
  .A({ S8107 }),
  .B({ S8110 }),
  .Y({ S8111 })
);
NAND #() 
NAND_4726_ (
  .A({ datapath_addsubunit_in1_2 }),
  .B({ S7967 }),
  .Y({ S8112 })
);
NAND #() 
NAND_4727_ (
  .A({ datapath_addsubunit_in1_14 }),
  .B({ S7995 }),
  .Y({ S8113 })
);
NAND #() 
NAND_4728_ (
  .A({ S8112 }),
  .B({ S8113 }),
  .Y({ S8114 })
);
NOR #() 
NOR_2964_ (
  .A({ S8111 }),
  .B({ S8114 }),
  .Y({ S8115 })
);
NAND #() 
NAND_4729_ (
  .A({ datapath_addsubunit_in1_10 }),
  .B({ S7984 }),
  .Y({ S8116 })
);
NAND #() 
NAND_4730_ (
  .A({ datapath_addsubunit_in1_11 }),
  .B({ S8020 }),
  .Y({ S8117 })
);
NAND #() 
NAND_4731_ (
  .A({ S8116 }),
  .B({ S8117 }),
  .Y({ S8118 })
);
NAND #() 
NAND_4732_ (
  .A({ datapath_addsubunit_in1_3 }),
  .B({ S8009 }),
  .Y({ S8120 })
);
NAND #() 
NAND_4733_ (
  .A({ datapath_addsubunit_in1_9 }),
  .B({ S8030 }),
  .Y({ S8121 })
);
NAND #() 
NAND_4734_ (
  .A({ S8120 }),
  .B({ S8121 }),
  .Y({ S8122 })
);
NOR #() 
NOR_2965_ (
  .A({ S8118 }),
  .B({ S8122 }),
  .Y({ S8123 })
);
NAND #() 
NAND_4735_ (
  .A({ S8115 }),
  .B({ S8123 }),
  .Y({ S8124 })
);
NOR #() 
NOR_2966_ (
  .A({ S8105 }),
  .B({ S8124 }),
  .Y({ S8125 })
);
NAND #() 
NAND_4736_ (
  .A({ S7958 }),
  .B({ S8078 }),
  .Y({ S8126 })
);
NOR #() 
NOR_2967_ (
  .A({ S7991 }),
  .B({ S8079 }),
  .Y({ S8127 })
);
NAND #() 
NAND_4737_ (
  .A({ S8102 }),
  .B({ S8125 }),
  .Y({ datapath_shiftunit_2171_A })
);
NAND #() 
NAND_4738_ (
  .A({ datapath_addsubunit_in1_7 }),
  .B({ S8002 }),
  .Y({ S8128 })
);
NAND #() 
NAND_4739_ (
  .A({ datapath_addsubunit_in1_10 }),
  .B({ S8030 }),
  .Y({ S8130 })
);
NAND #() 
NAND_4740_ (
  .A({ S8128 }),
  .B({ S8130 }),
  .Y({ S8131 })
);
NOR #() 
NOR_2968_ (
  .A({ S1065 }),
  .B({ S7969 }),
  .Y({ S8132 })
);
NAND #() 
NAND_4741_ (
  .A({ datapath_addsubunit_in1_3 }),
  .B({ S7967 }),
  .Y({ S8133 })
);
NAND #() 
NAND_4742_ (
  .A({ datapath_addsubunit_in1_11 }),
  .B({ S7984 }),
  .Y({ S8134 })
);
NAND #() 
NAND_4743_ (
  .A({ S8133 }),
  .B({ S8134 }),
  .Y({ S8135 })
);
NAND #() 
NAND_4744_ (
  .A({ datapath_addsubunit_in1_14 }),
  .B({ S8006 }),
  .Y({ S8136 })
);
NOR #() 
NOR_2969_ (
  .A({ S1611 }),
  .B({ S7950 }),
  .Y({ S8137 })
);
NOR #() 
NOR_2970_ (
  .A({ S7991 }),
  .B({ S8137 }),
  .Y({ S8138 })
);
NAND #() 
NAND_4745_ (
  .A({ datapath_addsubunit_in1_15 }),
  .B({ S8138 }),
  .Y({ S8139 })
);
NAND #() 
NAND_4746_ (
  .A({ S8136 }),
  .B({ S8139 }),
  .Y({ S8141 })
);
NOR #() 
NOR_2971_ (
  .A({ S8135 }),
  .B({ S8141 }),
  .Y({ S8142 })
);
NOT #() 
NOT_553_ (
  .A({ S8142 }),
  .Y({ S8143 })
);
NOR #() 
NOR_2972_ (
  .A({ S8131 }),
  .B({ S8143 }),
  .Y({ S8144 })
);
NAND #() 
NAND_4747_ (
  .A({ datapath_addsubunit_in1_4 }),
  .B({ S8009 }),
  .Y({ S8145 })
);
NOR #() 
NOR_2973_ (
  .A({ S599 }),
  .B({ S8021 }),
  .Y({ S8146 })
);
NOR #() 
NOR_2974_ (
  .A({ S910 }),
  .B({ S7974 }),
  .Y({ S8147 })
);
NAND #() 
NAND_4748_ (
  .A({ datapath_addsubunit_in1_6 }),
  .B({ S7973 }),
  .Y({ S8148 })
);
NOR #() 
NOR_2975_ (
  .A({ S8146 }),
  .B({ S8147 }),
  .Y({ S8149 })
);
NAND #() 
NAND_4749_ (
  .A({ S8145 }),
  .B({ S8149 }),
  .Y({ S8150 })
);
NOR #() 
NOR_2976_ (
  .A({ S805 }),
  .B({ S8025 }),
  .Y({ S8152 })
);
NOR #() 
NOR_2977_ (
  .A({ S963 }),
  .B({ S8015 }),
  .Y({ S8153 })
);
NOR #() 
NOR_2978_ (
  .A({ S8152 }),
  .B({ S8153 }),
  .Y({ S8154 })
);
NOR #() 
NOR_2979_ (
  .A({ S548 }),
  .B({ S7981 }),
  .Y({ S8155 })
);
NOR #() 
NOR_2980_ (
  .A({ S754 }),
  .B({ S8018 }),
  .Y({ S8156 })
);
NAND #() 
NAND_4750_ (
  .A({ datapath_addsubunit_in1_9 }),
  .B({ S8017 }),
  .Y({ S8157 })
);
NOR #() 
NOR_2981_ (
  .A({ S8155 }),
  .B({ S8156 }),
  .Y({ S8158 })
);
NAND #() 
NAND_4751_ (
  .A({ S8154 }),
  .B({ S8158 }),
  .Y({ S8159 })
);
NOR #() 
NOR_2982_ (
  .A({ S8150 }),
  .B({ S8159 }),
  .Y({ S8160 })
);
NAND #() 
NAND_4752_ (
  .A({ S8144 }),
  .B({ S8160 }),
  .Y({ datapath_shiftunit_2189_A })
);
NOR #() 
NOR_2983_ (
  .A({ S805 }),
  .B({ S8003 }),
  .Y({ S8162 })
);
NOR #() 
NOR_2984_ (
  .A({ S1304 }),
  .B({ S8007 }),
  .Y({ S8163 })
);
NOR #() 
NOR_2985_ (
  .A({ S8162 }),
  .B({ S8163 }),
  .Y({ S8164 })
);
NOR #() 
NOR_2986_ (
  .A({ S754 }),
  .B({ S8025 }),
  .Y({ S8165 })
);
NAND #() 
NAND_4753_ (
  .A({ datapath_addsubunit_in1_9 }),
  .B({ S8024 }),
  .Y({ S8166 })
);
NOR #() 
NOR_2987_ (
  .A({ S651 }),
  .B({ S8031 }),
  .Y({ S8167 })
);
NOR #() 
NOR_2988_ (
  .A({ S8165 }),
  .B({ S8167 }),
  .Y({ S8168 })
);
NAND #() 
NAND_4754_ (
  .A({ S8164 }),
  .B({ S8168 }),
  .Y({ S8169 })
);
NOR #() 
NOR_2989_ (
  .A({ S8127 }),
  .B({ S8169 }),
  .Y({ S8170 })
);
NOR #() 
NOR_2990_ (
  .A({ S858 }),
  .B({ S7974 }),
  .Y({ S8171 })
);
NOR #() 
NOR_2991_ (
  .A({ S910 }),
  .B({ S8015 }),
  .Y({ S8173 })
);
NOR #() 
NOR_2992_ (
  .A({ S8171 }),
  .B({ S8173 }),
  .Y({ S8174 })
);
NOR #() 
NOR_2993_ (
  .A({ S963 }),
  .B({ S8010 }),
  .Y({ S8175 })
);
NAND #() 
NAND_4755_ (
  .A({ datapath_addsubunit_in1_5 }),
  .B({ S8009 }),
  .Y({ S8176 })
);
NOR #() 
NOR_2994_ (
  .A({ S1013 }),
  .B({ S7969 }),
  .Y({ S8177 })
);
NAND #() 
NAND_4756_ (
  .A({ datapath_addsubunit_in1_4 }),
  .B({ S7967 }),
  .Y({ S8178 })
);
NOR #() 
NOR_2995_ (
  .A({ S8175 }),
  .B({ S8177 }),
  .Y({ S8179 })
);
NAND #() 
NAND_4757_ (
  .A({ S8174 }),
  .B({ S8179 }),
  .Y({ S8180 })
);
NOR #() 
NOR_2996_ (
  .A({ S548 }),
  .B({ S8021 }),
  .Y({ S8181 })
);
NOR #() 
NOR_2997_ (
  .A({ S702 }),
  .B({ S8018 }),
  .Y({ S8182 })
);
NOR #() 
NOR_2998_ (
  .A({ S8181 }),
  .B({ S8182 }),
  .Y({ S8184 })
);
NOR #() 
NOR_2999_ (
  .A({ S492 }),
  .B({ S7981 }),
  .Y({ S8185 })
);
NOR #() 
NOR_3000_ (
  .A({ S599 }),
  .B({ S7985 }),
  .Y({ S8186 })
);
NOR #() 
NOR_3001_ (
  .A({ S8185 }),
  .B({ S8186 }),
  .Y({ S8187 })
);
NAND #() 
NAND_4758_ (
  .A({ S8184 }),
  .B({ S8187 }),
  .Y({ S8188 })
);
NOR #() 
NOR_3002_ (
  .A({ S8180 }),
  .B({ S8188 }),
  .Y({ S8189 })
);
NAND #() 
NAND_4759_ (
  .A({ S8170 }),
  .B({ S8189 }),
  .Y({ datapath_shiftunit_2207_A })
);
NOR #() 
NOR_3003_ (
  .A({ S7990 }),
  .B({ S8006 }),
  .Y({ S8190 })
);
NOR #() 
NOR_3004_ (
  .A({ S8079 }),
  .B({ S8190 }),
  .Y({ S8191 })
);
NOR #() 
NOR_3005_ (
  .A({ S492 }),
  .B({ S8021 }),
  .Y({ S8192 })
);
NOR #() 
NOR_3006_ (
  .A({ S910 }),
  .B({ S8010 }),
  .Y({ S8194 })
);
NOR #() 
NOR_3007_ (
  .A({ S8192 }),
  .B({ S8194 }),
  .Y({ S8195 })
);
NOR #() 
NOR_3008_ (
  .A({ S651 }),
  .B({ S8018 }),
  .Y({ S8196 })
);
NOR #() 
NOR_3009_ (
  .A({ S805 }),
  .B({ S7974 }),
  .Y({ S8197 })
);
NOR #() 
NOR_3010_ (
  .A({ S8196 }),
  .B({ S8197 }),
  .Y({ S8198 })
);
NAND #() 
NAND_4760_ (
  .A({ S8195 }),
  .B({ S8198 }),
  .Y({ S8199 })
);
NOR #() 
NOR_3011_ (
  .A({ S8191 }),
  .B({ S8199 }),
  .Y({ S8200 })
);
NAND #() 
NAND_4761_ (
  .A({ datapath_addsubunit_in1_10 }),
  .B({ S8024 }),
  .Y({ S8201 })
);
NOR #() 
NOR_3012_ (
  .A({ S858 }),
  .B({ S8015 }),
  .Y({ S8202 })
);
NOR #() 
NOR_3013_ (
  .A({ S754 }),
  .B({ S8003 }),
  .Y({ S8203 })
);
NOR #() 
NOR_3014_ (
  .A({ S8202 }),
  .B({ S8203 }),
  .Y({ S8205 })
);
NAND #() 
NAND_4762_ (
  .A({ S8201 }),
  .B({ S8205 }),
  .Y({ S8206 })
);
NOR #() 
NOR_3015_ (
  .A({ S1304 }),
  .B({ S7981 }),
  .Y({ S8207 })
);
NOR #() 
NOR_3016_ (
  .A({ S599 }),
  .B({ S8031 }),
  .Y({ S8208 })
);
NOR #() 
NOR_3017_ (
  .A({ S8207 }),
  .B({ S8208 }),
  .Y({ S8209 })
);
NOR #() 
NOR_3018_ (
  .A({ S963 }),
  .B({ S7969 }),
  .Y({ S8210 })
);
NOR #() 
NOR_3019_ (
  .A({ S548 }),
  .B({ S7985 }),
  .Y({ S8211 })
);
NOR #() 
NOR_3020_ (
  .A({ S8210 }),
  .B({ S8211 }),
  .Y({ S8212 })
);
NAND #() 
NAND_4763_ (
  .A({ S8209 }),
  .B({ S8212 }),
  .Y({ S8213 })
);
NOR #() 
NOR_3021_ (
  .A({ S8206 }),
  .B({ S8213 }),
  .Y({ S8214 })
);
NAND #() 
NAND_4764_ (
  .A({ S8200 }),
  .B({ S8214 }),
  .Y({ datapath_shiftunit_2225_A })
);
NOR #() 
NOR_3022_ (
  .A({ S548 }),
  .B({ S8031 }),
  .Y({ S8216 })
);
NOR #() 
NOR_3023_ (
  .A({ S651 }),
  .B({ S8025 }),
  .Y({ S8217 })
);
NOR #() 
NOR_3024_ (
  .A({ S805 }),
  .B({ S8015 }),
  .Y({ S8218 })
);
NAND #() 
NAND_4765_ (
  .A({ datapath_addsubunit_in1_15 }),
  .B({ S8020 }),
  .Y({ S8219 })
);
NOR #() 
NOR_3025_ (
  .A({ S858 }),
  .B({ S8010 }),
  .Y({ S8220 })
);
NAND #() 
NAND_4766_ (
  .A({ datapath_addsubunit_in1_7 }),
  .B({ S8009 }),
  .Y({ S8221 })
);
NAND #() 
NAND_4767_ (
  .A({ datapath_addsubunit_in1_9 }),
  .B({ S7973 }),
  .Y({ S8222 })
);
NAND #() 
NAND_4768_ (
  .A({ S7981 }),
  .B({ S8190 }),
  .Y({ S8223 })
);
NAND #() 
NAND_4769_ (
  .A({ S8078 }),
  .B({ S8223 }),
  .Y({ S8224 })
);
NOR #() 
NOR_3026_ (
  .A({ S492 }),
  .B({ S7985 }),
  .Y({ S8226 })
);
NOR #() 
NOR_3027_ (
  .A({ S599 }),
  .B({ S8018 }),
  .Y({ S8227 })
);
NAND #() 
NAND_4770_ (
  .A({ datapath_addsubunit_in1_10 }),
  .B({ S8002 }),
  .Y({ S8228 })
);
NOR #() 
NOR_3028_ (
  .A({ S910 }),
  .B({ S7969 }),
  .Y({ S8229 })
);
NAND #() 
NAND_4771_ (
  .A({ datapath_addsubunit_in1_6 }),
  .B({ S7967 }),
  .Y({ S8230 })
);
NOR #() 
NOR_3029_ (
  .A({ S8217 }),
  .B({ S8218 }),
  .Y({ S8231 })
);
NOR #() 
NOR_3030_ (
  .A({ S8216 }),
  .B({ S8226 }),
  .Y({ S8232 })
);
NAND #() 
NAND_4772_ (
  .A({ S8221 }),
  .B({ S8232 }),
  .Y({ S8233 })
);
NAND #() 
NAND_4773_ (
  .A({ S8224 }),
  .B({ S8231 }),
  .Y({ S8234 })
);
NOR #() 
NOR_3031_ (
  .A({ S8233 }),
  .B({ S8234 }),
  .Y({ S8235 })
);
NAND #() 
NAND_4774_ (
  .A({ S8219 }),
  .B({ S8228 }),
  .Y({ S8237 })
);
NOR #() 
NOR_3032_ (
  .A({ S8227 }),
  .B({ S8229 }),
  .Y({ S8238 })
);
NAND #() 
NAND_4775_ (
  .A({ S8222 }),
  .B({ S8238 }),
  .Y({ S8239 })
);
NOR #() 
NOR_3033_ (
  .A({ S8237 }),
  .B({ S8239 }),
  .Y({ S8240 })
);
NAND #() 
NAND_4776_ (
  .A({ S8235 }),
  .B({ S8240 }),
  .Y({ datapath_shiftunit_2243_A })
);
NOR #() 
NOR_3034_ (
  .A({ S702 }),
  .B({ S7974 }),
  .Y({ S8241 })
);
NAND #() 
NAND_4777_ (
  .A({ datapath_addsubunit_in1_10 }),
  .B({ S7973 }),
  .Y({ S8242 })
);
NOR #() 
NOR_3035_ (
  .A({ S548 }),
  .B({ S8018 }),
  .Y({ S8243 })
);
NOR #() 
NOR_3036_ (
  .A({ S754 }),
  .B({ S8015 }),
  .Y({ S8244 })
);
NAND #() 
NAND_4778_ (
  .A({ datapath_addsubunit_in1_11 }),
  .B({ S8002 }),
  .Y({ S8245 })
);
NOR #() 
NOR_3037_ (
  .A({ S858 }),
  .B({ S7969 }),
  .Y({ S8247 })
);
NOR #() 
NOR_3038_ (
  .A({ S1304 }),
  .B({ S7985 }),
  .Y({ S8248 })
);
NOR #() 
NOR_3039_ (
  .A({ S599 }),
  .B({ S8025 }),
  .Y({ S8249 })
);
NOR #() 
NOR_3040_ (
  .A({ S492 }),
  .B({ S8031 }),
  .Y({ S8250 })
);
NOR #() 
NOR_3041_ (
  .A({ S805 }),
  .B({ S8010 }),
  .Y({ S8251 })
);
NOR #() 
NOR_3042_ (
  .A({ S8247 }),
  .B({ S8249 }),
  .Y({ S8252 })
);
NOR #() 
NOR_3043_ (
  .A({ S8241 }),
  .B({ S8251 }),
  .Y({ S8253 })
);
NAND #() 
NAND_4779_ (
  .A({ S8252 }),
  .B({ S8253 }),
  .Y({ S8254 })
);
NOR #() 
NOR_3044_ (
  .A({ S8021 }),
  .B({ S8079 }),
  .Y({ S8255 })
);
NOR #() 
NOR_3045_ (
  .A({ S8254 }),
  .B({ S8255 }),
  .Y({ S8256 })
);
NOR #() 
NOR_3046_ (
  .A({ S8243 }),
  .B({ S8248 }),
  .Y({ S8258 })
);
NAND #() 
NAND_4780_ (
  .A({ S8245 }),
  .B({ S8258 }),
  .Y({ S8259 })
);
NOR #() 
NOR_3047_ (
  .A({ S8244 }),
  .B({ S8250 }),
  .Y({ S8260 })
);
NAND #() 
NAND_4781_ (
  .A({ S8224 }),
  .B({ S8260 }),
  .Y({ S8261 })
);
NOR #() 
NOR_3048_ (
  .A({ S8259 }),
  .B({ S8261 }),
  .Y({ S8262 })
);
NAND #() 
NAND_4782_ (
  .A({ S8256 }),
  .B({ S8262 }),
  .Y({ datapath_shiftunit_2261_A })
);
NOR #() 
NOR_3049_ (
  .A({ S1304 }),
  .B({ S8031 }),
  .Y({ S8263 })
);
NOR #() 
NOR_3050_ (
  .A({ S548 }),
  .B({ S8025 }),
  .Y({ S8264 })
);
NOR #() 
NOR_3051_ (
  .A({ S754 }),
  .B({ S8010 }),
  .Y({ S8265 })
);
NOR #() 
NOR_3052_ (
  .A({ S599 }),
  .B({ S8003 }),
  .Y({ S8266 })
);
NOR #() 
NOR_3053_ (
  .A({ S492 }),
  .B({ S8018 }),
  .Y({ S8268 })
);
NOR #() 
NOR_3054_ (
  .A({ S651 }),
  .B({ S7974 }),
  .Y({ S8269 })
);
NOR #() 
NOR_3055_ (
  .A({ S805 }),
  .B({ S7969 }),
  .Y({ S8270 })
);
NOR #() 
NOR_3056_ (
  .A({ S702 }),
  .B({ S8015 }),
  .Y({ S8271 })
);
NAND #() 
NAND_4783_ (
  .A({ datapath_addsubunit_in1_10 }),
  .B({ S8014 }),
  .Y({ S8272 })
);
NOR #() 
NOR_3057_ (
  .A({ S8265 }),
  .B({ S8268 }),
  .Y({ S8273 })
);
NOR #() 
NOR_3058_ (
  .A({ S8266 }),
  .B({ S8270 }),
  .Y({ S8274 })
);
NAND #() 
NAND_4784_ (
  .A({ S8126 }),
  .B({ S8274 }),
  .Y({ S8275 })
);
NOR #() 
NOR_3059_ (
  .A({ S8263 }),
  .B({ S8269 }),
  .Y({ S8276 })
);
NOR #() 
NOR_3060_ (
  .A({ S8264 }),
  .B({ S8271 }),
  .Y({ S8277 })
);
NAND #() 
NAND_4785_ (
  .A({ S8276 }),
  .B({ S8277 }),
  .Y({ S8279 })
);
NOR #() 
NOR_3061_ (
  .A({ S8275 }),
  .B({ S8279 }),
  .Y({ S8280 })
);
NAND #() 
NAND_4786_ (
  .A({ S8273 }),
  .B({ S8280 }),
  .Y({ datapath_shiftunit_2279_A })
);
NAND #() 
NAND_4787_ (
  .A({ datapath_addsubunit_in1_12 }),
  .B({ S7973 }),
  .Y({ S8281 })
);
NAND #() 
NAND_4788_ (
  .A({ datapath_addsubunit_in1_13 }),
  .B({ S8002 }),
  .Y({ S8282 })
);
NAND #() 
NAND_4789_ (
  .A({ datapath_addsubunit_in1_14 }),
  .B({ S8024 }),
  .Y({ S8283 })
);
NOR #() 
NOR_3062_ (
  .A({ S7941 }),
  .B({ S7963 }),
  .Y({ S8284 })
);
NOR #() 
NOR_3063_ (
  .A({ S7958 }),
  .B({ S8284 }),
  .Y({ S8285 })
);
NAND #() 
NAND_4790_ (
  .A({ S1612 }),
  .B({ S8018 }),
  .Y({ S8286 })
);
NAND #() 
NAND_4791_ (
  .A({ datapath_addsubunit_in1_15 }),
  .B({ S8286 }),
  .Y({ S8287 })
);
NOR #() 
NOR_3064_ (
  .A({ S8285 }),
  .B({ S8287 }),
  .Y({ S8289 })
);
NAND #() 
NAND_4792_ (
  .A({ datapath_addsubunit_in1_10 }),
  .B({ S8009 }),
  .Y({ S8290 })
);
NAND #() 
NAND_4793_ (
  .A({ datapath_addsubunit_in1_11 }),
  .B({ S8014 }),
  .Y({ S8291 })
);
NOR #() 
NOR_3065_ (
  .A({ S754 }),
  .B({ S7969 }),
  .Y({ S8292 })
);
NAND #() 
NAND_4794_ (
  .A({ datapath_addsubunit_in1_9 }),
  .B({ S7967 }),
  .Y({ S8293 })
);
NAND #() 
NAND_4795_ (
  .A({ S8283 }),
  .B({ S8293 }),
  .Y({ S8294 })
);
NAND #() 
NAND_4796_ (
  .A({ S8281 }),
  .B({ S8290 }),
  .Y({ S8295 })
);
NOR #() 
NOR_3066_ (
  .A({ S8294 }),
  .B({ S8295 }),
  .Y({ S8296 })
);
NAND #() 
NAND_4797_ (
  .A({ S8282 }),
  .B({ S8291 }),
  .Y({ S8297 })
);
NOR #() 
NOR_3067_ (
  .A({ S8289 }),
  .B({ S8297 }),
  .Y({ S8298 })
);
NAND #() 
NAND_4798_ (
  .A({ S8296 }),
  .B({ S8298 }),
  .Y({ datapath_shiftunit_2297_A })
);
NOR #() 
NOR_3068_ (
  .A({ S651 }),
  .B({ S8010 }),
  .Y({ S8300 })
);
NAND #() 
NAND_4799_ (
  .A({ datapath_addsubunit_in1_11 }),
  .B({ S8009 }),
  .Y({ S8301 })
);
NOR #() 
NOR_3069_ (
  .A({ S702 }),
  .B({ S7969 }),
  .Y({ S8302 })
);
NAND #() 
NAND_4800_ (
  .A({ datapath_addsubunit_in1_10 }),
  .B({ S7967 }),
  .Y({ S8303 })
);
NAND #() 
NAND_4801_ (
  .A({ S8301 }),
  .B({ S8303 }),
  .Y({ S8304 })
);
NAND #() 
NAND_4802_ (
  .A({ datapath_addsubunit_in1_13 }),
  .B({ S7973 }),
  .Y({ S8305 })
);
NAND #() 
NAND_4803_ (
  .A({ datapath_addsubunit_in1_15 }),
  .B({ S8024 }),
  .Y({ S8306 })
);
NAND #() 
NAND_4804_ (
  .A({ S8305 }),
  .B({ S8306 }),
  .Y({ S8307 })
);
NOR #() 
NOR_3070_ (
  .A({ S8304 }),
  .B({ S8307 }),
  .Y({ S8308 })
);
NAND #() 
NAND_4805_ (
  .A({ datapath_addsubunit_in1_12 }),
  .B({ S8014 }),
  .Y({ S8310 })
);
NAND #() 
NAND_4806_ (
  .A({ datapath_addsubunit_in1_14 }),
  .B({ S8002 }),
  .Y({ S8311 })
);
NAND #() 
NAND_4807_ (
  .A({ S8310 }),
  .B({ S8311 }),
  .Y({ S8312 })
);
NOR #() 
NOR_3071_ (
  .A({ S8079 }),
  .B({ S8285 }),
  .Y({ S8313 })
);
NOR #() 
NOR_3072_ (
  .A({ S8312 }),
  .B({ S8313 }),
  .Y({ S8314 })
);
NAND #() 
NAND_4808_ (
  .A({ S8308 }),
  .B({ S8314 }),
  .Y({ datapath_shiftunit_2315_A })
);
NAND #() 
NAND_4809_ (
  .A({ datapath_addsubunit_in1_15 }),
  .B({ S8002 }),
  .Y({ S8315 })
);
NAND #() 
NAND_4810_ (
  .A({ datapath_addsubunit_in1_13 }),
  .B({ S8014 }),
  .Y({ S8316 })
);
NOR #() 
NOR_3073_ (
  .A({ S492 }),
  .B({ S7974 }),
  .Y({ S8317 })
);
NOR #() 
NOR_3074_ (
  .A({ S8025 }),
  .B({ S8079 }),
  .Y({ S8318 })
);
NAND #() 
NAND_4811_ (
  .A({ datapath_addsubunit_in1_11 }),
  .B({ S7967 }),
  .Y({ S8320 })
);
NOR #() 
NOR_3075_ (
  .A({ S599 }),
  .B({ S8010 }),
  .Y({ S8321 })
);
NAND #() 
NAND_4812_ (
  .A({ S8315 }),
  .B({ S8316 }),
  .Y({ S8322 })
);
NOR #() 
NOR_3076_ (
  .A({ S8313 }),
  .B({ S8322 }),
  .Y({ S8323 })
);
NOR #() 
NOR_3077_ (
  .A({ S8317 }),
  .B({ S8321 }),
  .Y({ S8324 })
);
NAND #() 
NAND_4813_ (
  .A({ S8320 }),
  .B({ S8324 }),
  .Y({ S8325 })
);
NOR #() 
NOR_3078_ (
  .A({ S8318 }),
  .B({ S8325 }),
  .Y({ S8326 })
);
NAND #() 
NAND_4814_ (
  .A({ S8323 }),
  .B({ S8326 }),
  .Y({ datapath_shiftunit_2333_A })
);
NAND #() 
NAND_4815_ (
  .A({ S7966 }),
  .B({ S8078 }),
  .Y({ S8327 })
);
NOR #() 
NOR_3079_ (
  .A({ S599 }),
  .B({ S7969 }),
  .Y({ S8328 })
);
NAND #() 
NAND_4816_ (
  .A({ datapath_addsubunit_in1_12 }),
  .B({ S7967 }),
  .Y({ S8330 })
);
NAND #() 
NAND_4817_ (
  .A({ datapath_addsubunit_in1_15 }),
  .B({ S7973 }),
  .Y({ S8331 })
);
NAND #() 
NAND_4818_ (
  .A({ S8330 }),
  .B({ S8331 }),
  .Y({ S8332 })
);
NAND #() 
NAND_4819_ (
  .A({ datapath_addsubunit_in1_13 }),
  .B({ S8009 }),
  .Y({ S8333 })
);
NAND #() 
NAND_4820_ (
  .A({ datapath_addsubunit_in1_14 }),
  .B({ S8014 }),
  .Y({ S8334 })
);
NAND #() 
NAND_4821_ (
  .A({ S8333 }),
  .B({ S8334 }),
  .Y({ S8335 })
);
NOR #() 
NOR_3080_ (
  .A({ S8332 }),
  .B({ S8335 }),
  .Y({ S8336 })
);
NAND #() 
NAND_4822_ (
  .A({ S8327 }),
  .B({ S8336 }),
  .Y({ datapath_shiftunit_2351_A })
);
NOR #() 
NOR_3081_ (
  .A({ S7966 }),
  .B({ S7971 }),
  .Y({ S8337 })
);
NOR #() 
NOR_3082_ (
  .A({ S8079 }),
  .B({ S8337 }),
  .Y({ S8338 })
);
NAND #() 
NAND_4823_ (
  .A({ datapath_addsubunit_in1_14 }),
  .B({ S8009 }),
  .Y({ S8340 })
);
NOR #() 
NOR_3083_ (
  .A({ S548 }),
  .B({ S7969 }),
  .Y({ S8341 })
);
NAND #() 
NAND_4824_ (
  .A({ datapath_addsubunit_in1_13 }),
  .B({ S7967 }),
  .Y({ S8342 })
);
NAND #() 
NAND_4825_ (
  .A({ datapath_addsubunit_in1_15 }),
  .B({ S8014 }),
  .Y({ S8343 })
);
NAND #() 
NAND_4826_ (
  .A({ S8340 }),
  .B({ S8342 }),
  .Y({ S8344 })
);
NOR #() 
NOR_3084_ (
  .A({ S8338 }),
  .B({ S8344 }),
  .Y({ S8345 })
);
NAND #() 
NAND_4827_ (
  .A({ S8343 }),
  .B({ S8345 }),
  .Y({ datapath_shiftunit_2369_A })
);
NAND #() 
NAND_4828_ (
  .A({ datapath_addsubunit_in1_15 }),
  .B({ S8009 }),
  .Y({ S8346 })
);
NAND #() 
NAND_4829_ (
  .A({ datapath_addsubunit_in1_14 }),
  .B({ S7967 }),
  .Y({ S8347 })
);
NAND #() 
NAND_4830_ (
  .A({ S8346 }),
  .B({ S8347 }),
  .Y({ S8348 })
);
NOR #() 
NOR_3085_ (
  .A({ S8103 }),
  .B({ S8348 }),
  .Y({ S8350 })
);
NAND #() 
NAND_4831_ (
  .A({ S8327 }),
  .B({ S8350 }),
  .Y({ datapath_shiftunit_2387_A })
);
NAND #() 
NAND_4832_ (
  .A({ datapath_addsubunit_in1_15 }),
  .B({ S7967 }),
  .Y({ S8351 })
);
NAND #() 
NAND_4833_ (
  .A({ S8079 }),
  .B({ S8351 }),
  .Y({ datapath_shiftunit_2405_A })
);
NAND #() 
NAND_4834_ (
  .A({ datapath_addsubunit_in1_0 }),
  .B({ S8009 }),
  .Y({ S8352 })
);
NAND #() 
NAND_4835_ (
  .A({ S8067 }),
  .B({ S8352 }),
  .Y({ datapath_shiftunit_2457_A })
);
NOR #() 
NOR_3086_ (
  .A({ S1220 }),
  .B({ S8015 }),
  .Y({ S8353 })
);
NOR #() 
NOR_3087_ (
  .A({ S8012 }),
  .B({ S8353 }),
  .Y({ S8354 })
);
NAND #() 
NAND_4836_ (
  .A({ S8112 }),
  .B({ S8354 }),
  .Y({ datapath_shiftunit_2475_A })
);
NOR #() 
NOR_3088_ (
  .A({ S8055 }),
  .B({ S8132 }),
  .Y({ S8355 })
);
NOR #() 
NOR_3089_ (
  .A({ S1220 }),
  .B({ S7974 }),
  .Y({ S8357 })
);
NOR #() 
NOR_3090_ (
  .A({ S1168 }),
  .B({ S8015 }),
  .Y({ S8358 })
);
NOR #() 
NOR_3091_ (
  .A({ S8357 }),
  .B({ S8358 }),
  .Y({ S8359 })
);
NAND #() 
NAND_4837_ (
  .A({ S8355 }),
  .B({ S8359 }),
  .Y({ datapath_shiftunit_2493_A })
);
NAND #() 
NAND_4838_ (
  .A({ S8016 }),
  .B({ S8120 }),
  .Y({ S8360 })
);
NAND #() 
NAND_4839_ (
  .A({ datapath_addsubunit_in1_1 }),
  .B({ S7973 }),
  .Y({ S8361 })
);
NAND #() 
NAND_4840_ (
  .A({ datapath_addsubunit_in1_0 }),
  .B({ S8002 }),
  .Y({ S8362 })
);
NAND #() 
NAND_4841_ (
  .A({ S8178 }),
  .B({ S8362 }),
  .Y({ S8363 })
);
NOR #() 
NOR_3092_ (
  .A({ S8360 }),
  .B({ S8363 }),
  .Y({ S8364 })
);
NAND #() 
NAND_4842_ (
  .A({ S8361 }),
  .B({ S8364 }),
  .Y({ datapath_shiftunit_2511_A })
);
NAND #() 
NAND_4843_ (
  .A({ S8060 }),
  .B({ S8145 }),
  .Y({ S8366 })
);
NAND #() 
NAND_4844_ (
  .A({ datapath_addsubunit_in1_0 }),
  .B({ S8024 }),
  .Y({ S8367 })
);
NAND #() 
NAND_4845_ (
  .A({ datapath_addsubunit_in1_2 }),
  .B({ S7973 }),
  .Y({ S8368 })
);
NOR #() 
NOR_3093_ (
  .A({ S1168 }),
  .B({ S8003 }),
  .Y({ S8369 })
);
NOR #() 
NOR_3094_ (
  .A({ S8210 }),
  .B({ S8369 }),
  .Y({ S8370 })
);
NAND #() 
NAND_4846_ (
  .A({ S8367 }),
  .B({ S8368 }),
  .Y({ S8371 })
);
NOR #() 
NOR_3095_ (
  .A({ S8366 }),
  .B({ S8371 }),
  .Y({ S8372 })
);
NAND #() 
NAND_4847_ (
  .A({ S8370 }),
  .B({ S8372 }),
  .Y({ datapath_shiftunit_2529_A })
);
NOR #() 
NOR_3096_ (
  .A({ S1116 }),
  .B({ S8003 }),
  .Y({ S8373 })
);
NAND #() 
NAND_4848_ (
  .A({ datapath_addsubunit_in1_1 }),
  .B({ S8024 }),
  .Y({ S8374 })
);
NAND #() 
NAND_4849_ (
  .A({ datapath_addsubunit_in1_0 }),
  .B({ S8017 }),
  .Y({ S8376 })
);
NAND #() 
NAND_4850_ (
  .A({ S8374 }),
  .B({ S8376 }),
  .Y({ S8377 })
);
NOR #() 
NOR_3097_ (
  .A({ S8373 }),
  .B({ S8377 }),
  .Y({ S8378 })
);
NAND #() 
NAND_4851_ (
  .A({ S7975 }),
  .B({ S8091 }),
  .Y({ S8379 })
);
NAND #() 
NAND_4852_ (
  .A({ S8176 }),
  .B({ S8230 }),
  .Y({ S8380 })
);
NOR #() 
NOR_3098_ (
  .A({ S8379 }),
  .B({ S8380 }),
  .Y({ S8381 })
);
NAND #() 
NAND_4853_ (
  .A({ S8378 }),
  .B({ S8381 }),
  .Y({ datapath_shiftunit_2547_A })
);
NOR #() 
NOR_3099_ (
  .A({ S8153 }),
  .B({ S8194 }),
  .Y({ S8382 })
);
NOR #() 
NOR_3100_ (
  .A({ S8063 }),
  .B({ S8247 }),
  .Y({ S8383 })
);
NAND #() 
NAND_4854_ (
  .A({ S8382 }),
  .B({ S8383 }),
  .Y({ S8384 })
);
NAND #() 
NAND_4855_ (
  .A({ datapath_addsubunit_in1_1 }),
  .B({ S8017 }),
  .Y({ S8386 })
);
NOR #() 
NOR_3101_ (
  .A({ S1220 }),
  .B({ S8031 }),
  .Y({ S8387 })
);
NAND #() 
NAND_4856_ (
  .A({ datapath_addsubunit_in1_2 }),
  .B({ S8024 }),
  .Y({ S8388 })
);
NOR #() 
NOR_3102_ (
  .A({ S1065 }),
  .B({ S8003 }),
  .Y({ S8389 })
);
NAND #() 
NAND_4857_ (
  .A({ S8386 }),
  .B({ S8388 }),
  .Y({ S8390 })
);
NOR #() 
NOR_3103_ (
  .A({ S8389 }),
  .B({ S8390 }),
  .Y({ S8391 })
);
NOR #() 
NOR_3104_ (
  .A({ S8384 }),
  .B({ S8387 }),
  .Y({ S8392 })
);
NAND #() 
NAND_4858_ (
  .A({ S8391 }),
  .B({ S8392 }),
  .Y({ datapath_shiftunit_2565_A })
);
NOR #() 
NOR_3105_ (
  .A({ S1220 }),
  .B({ S7985 }),
  .Y({ S8393 })
);
NAND #() 
NAND_4859_ (
  .A({ datapath_addsubunit_in1_2 }),
  .B({ S8017 }),
  .Y({ S8394 })
);
NAND #() 
NAND_4860_ (
  .A({ datapath_addsubunit_in1_3 }),
  .B({ S8024 }),
  .Y({ S8396 })
);
NAND #() 
NAND_4861_ (
  .A({ S8394 }),
  .B({ S8396 }),
  .Y({ S8397 })
);
NOR #() 
NOR_3106_ (
  .A({ S8393 }),
  .B({ S8397 }),
  .Y({ S8398 })
);
NAND #() 
NAND_4862_ (
  .A({ S8005 }),
  .B({ S8092 }),
  .Y({ S8399 })
);
NOR #() 
NOR_3107_ (
  .A({ S8173 }),
  .B({ S8220 }),
  .Y({ S8400 })
);
NOR #() 
NOR_3108_ (
  .A({ S1168 }),
  .B({ S8031 }),
  .Y({ S8401 })
);
NOR #() 
NOR_3109_ (
  .A({ S8270 }),
  .B({ S8401 }),
  .Y({ S8402 })
);
NAND #() 
NAND_4863_ (
  .A({ S8400 }),
  .B({ S8402 }),
  .Y({ S8403 })
);
NOR #() 
NOR_3110_ (
  .A({ S8399 }),
  .B({ S8403 }),
  .Y({ S8404 })
);
NAND #() 
NAND_4864_ (
  .A({ S8398 }),
  .B({ S8404 }),
  .Y({ datapath_shiftunit_2583_A })
);
NAND #() 
NAND_4865_ (
  .A({ datapath_addsubunit_in1_1 }),
  .B({ S7984 }),
  .Y({ S8406 })
);
NAND #() 
NAND_4866_ (
  .A({ datapath_addsubunit_in1_0 }),
  .B({ S8020 }),
  .Y({ S8407 })
);
NAND #() 
NAND_4867_ (
  .A({ S8406 }),
  .B({ S8407 }),
  .Y({ S8408 })
);
NAND #() 
NAND_4868_ (
  .A({ datapath_addsubunit_in1_3 }),
  .B({ S8017 }),
  .Y({ S8409 })
);
NAND #() 
NAND_4869_ (
  .A({ datapath_addsubunit_in1_4 }),
  .B({ S8024 }),
  .Y({ S8410 })
);
NAND #() 
NAND_4870_ (
  .A({ S8409 }),
  .B({ S8410 }),
  .Y({ S8411 })
);
NOR #() 
NOR_3111_ (
  .A({ S8408 }),
  .B({ S8411 }),
  .Y({ S8412 })
);
NAND #() 
NAND_4871_ (
  .A({ S8058 }),
  .B({ S8148 }),
  .Y({ S8413 })
);
NOR #() 
NOR_3112_ (
  .A({ S8202 }),
  .B({ S8251 }),
  .Y({ S8414 })
);
NOR #() 
NOR_3113_ (
  .A({ S1116 }),
  .B({ S8031 }),
  .Y({ S8415 })
);
NOR #() 
NOR_3114_ (
  .A({ S8292 }),
  .B({ S8415 }),
  .Y({ S8417 })
);
NAND #() 
NAND_4872_ (
  .A({ S8414 }),
  .B({ S8417 }),
  .Y({ S8418 })
);
NOR #() 
NOR_3115_ (
  .A({ S8413 }),
  .B({ S8418 }),
  .Y({ S8419 })
);
NAND #() 
NAND_4873_ (
  .A({ S8412 }),
  .B({ S8419 }),
  .Y({ datapath_shiftunit_2601_A })
);
NOR #() 
NOR_3116_ (
  .A({ S1220 }),
  .B({ S7981 }),
  .Y({ S8420 })
);
NAND #() 
NAND_4874_ (
  .A({ datapath_addsubunit_in1_2 }),
  .B({ S7984 }),
  .Y({ S8421 })
);
NAND #() 
NAND_4875_ (
  .A({ datapath_addsubunit_in1_1 }),
  .B({ S8020 }),
  .Y({ S8422 })
);
NAND #() 
NAND_4876_ (
  .A({ S8421 }),
  .B({ S8422 }),
  .Y({ S8423 })
);
NOR #() 
NOR_3117_ (
  .A({ S8420 }),
  .B({ S8423 }),
  .Y({ S8424 })
);
NOR #() 
NOR_3118_ (
  .A({ S8265 }),
  .B({ S8302 }),
  .Y({ S8425 })
);
NOR #() 
NOR_3119_ (
  .A({ S1065 }),
  .B({ S8031 }),
  .Y({ S8427 })
);
NOR #() 
NOR_3120_ (
  .A({ S1013 }),
  .B({ S8018 }),
  .Y({ S8428 })
);
NOR #() 
NOR_3121_ (
  .A({ S8427 }),
  .B({ S8428 }),
  .Y({ S8429 })
);
NAND #() 
NAND_4877_ (
  .A({ S8425 }),
  .B({ S8429 }),
  .Y({ S8430 })
);
NOR #() 
NOR_3122_ (
  .A({ S8026 }),
  .B({ S8109 }),
  .Y({ S8431 })
);
NOR #() 
NOR_3123_ (
  .A({ S8171 }),
  .B({ S8218 }),
  .Y({ S8432 })
);
NAND #() 
NAND_4878_ (
  .A({ S8431 }),
  .B({ S8432 }),
  .Y({ S8433 })
);
NOR #() 
NOR_3124_ (
  .A({ S8430 }),
  .B({ S8433 }),
  .Y({ S8434 })
);
NAND #() 
NAND_4879_ (
  .A({ S8424 }),
  .B({ S8434 }),
  .Y({ datapath_shiftunit_2619_A })
);
NOR #() 
NOR_3125_ (
  .A({ S1065 }),
  .B({ S7985 }),
  .Y({ S8435 })
);
NOR #() 
NOR_3126_ (
  .A({ S1116 }),
  .B({ S8021 }),
  .Y({ S8437 })
);
NOR #() 
NOR_3127_ (
  .A({ S1220 }),
  .B({ S8007 }),
  .Y({ S8438 })
);
NOR #() 
NOR_3128_ (
  .A({ S963 }),
  .B({ S8018 }),
  .Y({ S8439 })
);
NOR #() 
NOR_3129_ (
  .A({ S1168 }),
  .B({ S7981 }),
  .Y({ S8440 })
);
NOR #() 
NOR_3130_ (
  .A({ S1013 }),
  .B({ S8031 }),
  .Y({ S8441 })
);
NOR #() 
NOR_3131_ (
  .A({ S8197 }),
  .B({ S8438 }),
  .Y({ S8442 })
);
NOR #() 
NOR_3132_ (
  .A({ S8439 }),
  .B({ S8440 }),
  .Y({ S8443 })
);
NAND #() 
NAND_4880_ (
  .A({ S8442 }),
  .B({ S8443 }),
  .Y({ S8444 })
);
NAND #() 
NAND_4881_ (
  .A({ S8053 }),
  .B({ S8290 }),
  .Y({ S8445 })
);
NOR #() 
NOR_3133_ (
  .A({ S8444 }),
  .B({ S8445 }),
  .Y({ S8446 })
);
NAND #() 
NAND_4882_ (
  .A({ S8128 }),
  .B({ S8320 }),
  .Y({ S8448 })
);
NOR #() 
NOR_3134_ (
  .A({ S8244 }),
  .B({ S8435 }),
  .Y({ S8449 })
);
NOR #() 
NOR_3135_ (
  .A({ S8437 }),
  .B({ S8441 }),
  .Y({ S8450 })
);
NAND #() 
NAND_4883_ (
  .A({ S8449 }),
  .B({ S8450 }),
  .Y({ S8451 })
);
NOR #() 
NOR_3136_ (
  .A({ S8448 }),
  .B({ S8451 }),
  .Y({ S8452 })
);
NAND #() 
NAND_4884_ (
  .A({ S8446 }),
  .B({ S8452 }),
  .Y({ datapath_shiftunit_2637_A })
);
NOR #() 
NOR_3137_ (
  .A({ S8019 }),
  .B({ S8098 }),
  .Y({ S8453 })
);
NOR #() 
NOR_3138_ (
  .A({ S963 }),
  .B({ S8031 }),
  .Y({ S8454 })
);
NOR #() 
NOR_3139_ (
  .A({ S1065 }),
  .B({ S8021 }),
  .Y({ S8455 })
);
NOR #() 
NOR_3140_ (
  .A({ S1013 }),
  .B({ S7985 }),
  .Y({ S8456 })
);
NAND #() 
NAND_4885_ (
  .A({ datapath_addsubunit_in1_0 }),
  .B({ S7995 }),
  .Y({ S8458 })
);
NOR #() 
NOR_3141_ (
  .A({ S1168 }),
  .B({ S8007 }),
  .Y({ S8459 })
);
NOR #() 
NOR_3142_ (
  .A({ S1116 }),
  .B({ S7981 }),
  .Y({ S8460 })
);
NOR #() 
NOR_3143_ (
  .A({ S8162 }),
  .B({ S8300 }),
  .Y({ S8461 })
);
NAND #() 
NAND_4886_ (
  .A({ S8453 }),
  .B({ S8461 }),
  .Y({ S8462 })
);
NOR #() 
NOR_3144_ (
  .A({ S8455 }),
  .B({ S8459 }),
  .Y({ S8463 })
);
NAND #() 
NAND_4887_ (
  .A({ S8458 }),
  .B({ S8463 }),
  .Y({ S8464 })
);
NOR #() 
NOR_3145_ (
  .A({ S8462 }),
  .B({ S8464 }),
  .Y({ S8465 })
);
NAND #() 
NAND_4888_ (
  .A({ S8222 }),
  .B({ S8272 }),
  .Y({ S8466 })
);
NOR #() 
NOR_3146_ (
  .A({ S8456 }),
  .B({ S8460 }),
  .Y({ S8467 })
);
NOR #() 
NOR_3147_ (
  .A({ S8328 }),
  .B({ S8454 }),
  .Y({ S8469 })
);
NAND #() 
NAND_4889_ (
  .A({ S8467 }),
  .B({ S8469 }),
  .Y({ S8470 })
);
NOR #() 
NOR_3148_ (
  .A({ S8466 }),
  .B({ S8470 }),
  .Y({ S8471 })
);
NAND #() 
NAND_4890_ (
  .A({ S8465 }),
  .B({ S8471 }),
  .Y({ datapath_shiftunit_2655_A })
);
NOR #() 
NOR_3149_ (
  .A({ S8061 }),
  .B({ S8152 }),
  .Y({ S8472 })
);
NOR #() 
NOR_3150_ (
  .A({ S1168 }),
  .B({ S7996 }),
  .Y({ S8473 })
);
NOR #() 
NOR_3151_ (
  .A({ S1013 }),
  .B({ S8021 }),
  .Y({ S8474 })
);
NOR #() 
NOR_3152_ (
  .A({ S8473 }),
  .B({ S8474 }),
  .Y({ S8475 })
);
NOR #() 
NOR_3153_ (
  .A({ S1116 }),
  .B({ S8007 }),
  .Y({ S8476 })
);
NOR #() 
NOR_3154_ (
  .A({ S1065 }),
  .B({ S7981 }),
  .Y({ S8477 })
);
NOR #() 
NOR_3155_ (
  .A({ S910 }),
  .B({ S8031 }),
  .Y({ S8479 })
);
NOR #() 
NOR_3156_ (
  .A({ S963 }),
  .B({ S7985 }),
  .Y({ S8480 })
);
NOR #() 
NOR_3157_ (
  .A({ S1220 }),
  .B({ S7992 }),
  .Y({ S8481 })
);
NOR #() 
NOR_3158_ (
  .A({ S8203 }),
  .B({ S8321 }),
  .Y({ S8482 })
);
NAND #() 
NAND_4891_ (
  .A({ S8472 }),
  .B({ S8482 }),
  .Y({ S8483 })
);
NOR #() 
NOR_3159_ (
  .A({ S8479 }),
  .B({ S8480 }),
  .Y({ S8484 })
);
NOR #() 
NOR_3160_ (
  .A({ S8477 }),
  .B({ S8481 }),
  .Y({ S8485 })
);
NAND #() 
NAND_4892_ (
  .A({ S8484 }),
  .B({ S8485 }),
  .Y({ S8486 })
);
NOR #() 
NOR_3161_ (
  .A({ S8483 }),
  .B({ S8486 }),
  .Y({ S8487 })
);
NOR #() 
NOR_3162_ (
  .A({ S8341 }),
  .B({ S8476 }),
  .Y({ S8488 })
);
NAND #() 
NAND_4893_ (
  .A({ S8475 }),
  .B({ S8488 }),
  .Y({ S8490 })
);
NAND #() 
NAND_4894_ (
  .A({ S8242 }),
  .B({ S8291 }),
  .Y({ S8491 })
);
NOR #() 
NOR_3163_ (
  .A({ S8490 }),
  .B({ S8491 }),
  .Y({ S8492 })
);
NAND #() 
NAND_4895_ (
  .A({ S8487 }),
  .B({ S8492 }),
  .Y({ datapath_shiftunit_2673_A })
);
NOR #() 
NOR_3164_ (
  .A({ S963 }),
  .B({ S8021 }),
  .Y({ S8493 })
);
NAND #() 
NAND_4896_ (
  .A({ datapath_addsubunit_in1_6 }),
  .B({ S7984 }),
  .Y({ S8494 })
);
NAND #() 
NAND_4897_ (
  .A({ datapath_addsubunit_in1_3 }),
  .B({ S8006 }),
  .Y({ S8495 })
);
NAND #() 
NAND_4898_ (
  .A({ datapath_addsubunit_in1_0 }),
  .B({ S8027 }),
  .Y({ S8496 })
);
NOR #() 
NOR_3165_ (
  .A({ S1013 }),
  .B({ S7981 }),
  .Y({ S8497 })
);
NAND #() 
NAND_4899_ (
  .A({ datapath_addsubunit_in1_2 }),
  .B({ S7995 }),
  .Y({ S8498 })
);
NOR #() 
NOR_3166_ (
  .A({ S1168 }),
  .B({ S7992 }),
  .Y({ S8500 })
);
NOR #() 
NOR_3167_ (
  .A({ S8106 }),
  .B({ S8269 }),
  .Y({ S8501 })
);
NAND #() 
NAND_4900_ (
  .A({ S8496 }),
  .B({ S8498 }),
  .Y({ S8502 })
);
NOR #() 
NOR_3168_ (
  .A({ S8493 }),
  .B({ S8502 }),
  .Y({ S8503 })
);
NAND #() 
NAND_4901_ (
  .A({ S8034 }),
  .B({ S8166 }),
  .Y({ S8504 })
);
NAND #() 
NAND_4902_ (
  .A({ S8333 }),
  .B({ S8494 }),
  .Y({ S8505 })
);
NOR #() 
NOR_3169_ (
  .A({ S8504 }),
  .B({ S8505 }),
  .Y({ S8506 })
);
NAND #() 
NAND_4903_ (
  .A({ S8503 }),
  .B({ S8506 }),
  .Y({ S8507 })
);
NAND #() 
NAND_4904_ (
  .A({ S8228 }),
  .B({ S8495 }),
  .Y({ S8508 })
);
NOR #() 
NOR_3170_ (
  .A({ S8497 }),
  .B({ S8508 }),
  .Y({ S8509 })
);
NAND #() 
NAND_4905_ (
  .A({ S8310 }),
  .B({ S8347 }),
  .Y({ S8511 })
);
NOR #() 
NOR_3171_ (
  .A({ S8500 }),
  .B({ S8511 }),
  .Y({ S8512 })
);
NAND #() 
NAND_4906_ (
  .A({ S8509 }),
  .B({ S8512 }),
  .Y({ S8513 })
);
NOR #() 
NOR_3172_ (
  .A({ S8507 }),
  .B({ S8513 }),
  .Y({ S8514 })
);
NAND #() 
NAND_4907_ (
  .A({ S8501 }),
  .B({ S8514 }),
  .Y({ datapath_shiftunit_2691_A })
);
NAND #() 
NAND_4908_ (
  .A({ S8281 }),
  .B({ S8316 }),
  .Y({ S8515 })
);
NAND #() 
NAND_4909_ (
  .A({ S8340 }),
  .B({ S8351 }),
  .Y({ S8516 })
);
NOR #() 
NOR_3173_ (
  .A({ S8515 }),
  .B({ S8516 }),
  .Y({ S8517 })
);
NAND #() 
NAND_4910_ (
  .A({ S8070 }),
  .B({ S8157 }),
  .Y({ S8518 })
);
NAND #() 
NAND_4911_ (
  .A({ S8201 }),
  .B({ S8245 }),
  .Y({ S8519 })
);
NOR #() 
NOR_3174_ (
  .A({ S8518 }),
  .B({ S8519 }),
  .Y({ S8521 })
);
NAND #() 
NAND_4912_ (
  .A({ S8517 }),
  .B({ S8521 }),
  .Y({ S8522 })
);
NAND #() 
NAND_4913_ (
  .A({ datapath_addsubunit_in1_2 }),
  .B({ S7993 }),
  .Y({ S8523 })
);
NAND #() 
NAND_4914_ (
  .A({ datapath_addsubunit_in1_7 }),
  .B({ S7984 }),
  .Y({ S8524 })
);
NAND #() 
NAND_4915_ (
  .A({ S8523 }),
  .B({ S8524 }),
  .Y({ S8525 })
);
NAND #() 
NAND_4916_ (
  .A({ datapath_addsubunit_in1_3 }),
  .B({ S7995 }),
  .Y({ S8526 })
);
NAND #() 
NAND_4917_ (
  .A({ datapath_addsubunit_in1_1 }),
  .B({ S8027 }),
  .Y({ S8527 })
);
NAND #() 
NAND_4918_ (
  .A({ S8526 }),
  .B({ S8527 }),
  .Y({ S8528 })
);
NOR #() 
NOR_3175_ (
  .A({ S8525 }),
  .B({ S8528 }),
  .Y({ S8529 })
);
NAND #() 
NAND_4919_ (
  .A({ datapath_addsubunit_in1_6 }),
  .B({ S8020 }),
  .Y({ S8530 })
);
NAND #() 
NAND_4920_ (
  .A({ datapath_addsubunit_in1_4 }),
  .B({ S8006 }),
  .Y({ S8532 })
);
NAND #() 
NAND_4921_ (
  .A({ S8530 }),
  .B({ S8532 }),
  .Y({ S8533 })
);
NOR #() 
NOR_3176_ (
  .A({ S963 }),
  .B({ S7981 }),
  .Y({ S8534 })
);
NOT #() 
NOT_554_ (
  .A({ S8534 }),
  .Y({ S8535 })
);
NAND #() 
NAND_4922_ (
  .A({ datapath_addsubunit_in1_0 }),
  .B({ S8035 }),
  .Y({ S8536 })
);
NAND #() 
NAND_4923_ (
  .A({ S8535 }),
  .B({ S8536 }),
  .Y({ S8537 })
);
NOR #() 
NOR_3177_ (
  .A({ S8533 }),
  .B({ S8537 }),
  .Y({ S8538 })
);
NAND #() 
NAND_4924_ (
  .A({ S8529 }),
  .B({ S8538 }),
  .Y({ S8539 })
);
NOR #() 
NOR_3178_ (
  .A({ S8522 }),
  .B({ S8539 }),
  .Y({ S8540 })
);
NOT #() 
NOT_555_ (
  .A({ S8540 }),
  .Y({ datapath_shiftunit_2708_A })
);
BUF #() 
BUF_1_ (
  .A({ datapath_theregisterfile_memtrf_240 }),
  .Y({ S244 })
);
BUF #() 
BUF_2_ (
  .A({ datapath_theregisterfile_memtrf_241 }),
  .Y({ S245 })
);
BUF #() 
BUF_3_ (
  .A({ datapath_theregisterfile_memtrf_242 }),
  .Y({ S246 })
);
BUF #() 
BUF_4_ (
  .A({ datapath_theregisterfile_memtrf_243 }),
  .Y({ S247 })
);
BUF #() 
BUF_5_ (
  .A({ datapath_theregisterfile_memtrf_244 }),
  .Y({ S248 })
);
BUF #() 
BUF_6_ (
  .A({ datapath_theregisterfile_memtrf_245 }),
  .Y({ S249 })
);
BUF #() 
BUF_7_ (
  .A({ datapath_theregisterfile_memtrf_246 }),
  .Y({ S250 })
);
BUF #() 
BUF_8_ (
  .A({ datapath_theregisterfile_memtrf_247 }),
  .Y({ S251 })
);
BUF #() 
BUF_9_ (
  .A({ datapath_theregisterfile_memtrf_248 }),
  .Y({ S252 })
);
BUF #() 
BUF_10_ (
  .A({ datapath_theregisterfile_memtrf_249 }),
  .Y({ S253 })
);
BUF #() 
BUF_11_ (
  .A({ datapath_theregisterfile_memtrf_250 }),
  .Y({ S254 })
);
BUF #() 
BUF_12_ (
  .A({ datapath_theregisterfile_memtrf_251 }),
  .Y({ S255 })
);
BUF #() 
BUF_13_ (
  .A({ datapath_theregisterfile_memtrf_252 }),
  .Y({ S256 })
);
BUF #() 
BUF_14_ (
  .A({ datapath_theregisterfile_memtrf_253 }),
  .Y({ S257 })
);
BUF #() 
BUF_15_ (
  .A({ datapath_theregisterfile_memtrf_254 }),
  .Y({ S258 })
);
BUF #() 
BUF_16_ (
  .A({ datapath_theregisterfile_memtrf_255 }),
  .Y({ S259 })
);
BUF #() 
BUF_17_ (
  .A({ controller_outflag_0 }),
  .Y({ S260 })
);
BUF #() 
BUF_18_ (
  .A({ controller_outflag_1 }),
  .Y({ S261 })
);
BUF #() 
BUF_19_ (
  .A({ controller_outflag_2 }),
  .Y({ S262 })
);
BUF #() 
BUF_20_ (
  .A({ controller_outflag_3 }),
  .Y({ S263 })
);
BUF #() 
BUF_21_ (
  .A({ controller_outflag_6 }),
  .Y({ S266 })
);
BUF #() 
BUF_22_ (
  .A({ controller_outflag_7 }),
  .Y({ S343 })
);
DFF_PP0 #() 
DFF_PP0_1_ (
  .C({ controller_clk }),
  .D({ controller_1405_Y_0 }),
  .Q({ controller_pstate_0 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_2_ (
  .C({ controller_clk }),
  .D({ controller_1405_Y_1 }),
  .Q({ controller_pstate_1 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_3_ (
  .C({ controller_clk }),
  .D({ S328 }),
  .Q({ datapath_adr_outreg_0 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_4_ (
  .C({ controller_clk }),
  .D({ S329 }),
  .Q({ datapath_adr_outreg_1 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_5_ (
  .C({ controller_clk }),
  .D({ S330 }),
  .Q({ datapath_adr_outreg_2 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_6_ (
  .C({ controller_clk }),
  .D({ S331 }),
  .Q({ datapath_adr_outreg_3 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_7_ (
  .C({ controller_clk }),
  .D({ S332 }),
  .Q({ datapath_adr_outreg_4 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_8_ (
  .C({ controller_clk }),
  .D({ S333 }),
  .Q({ datapath_adr_outreg_5 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_9_ (
  .C({ controller_clk }),
  .D({ S334 }),
  .Q({ datapath_adr_outreg_6 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_10_ (
  .C({ controller_clk }),
  .D({ S335 }),
  .Q({ datapath_adr_outreg_7 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_11_ (
  .C({ controller_clk }),
  .D({ S336 }),
  .Q({ datapath_adr_outreg_8 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_12_ (
  .C({ controller_clk }),
  .D({ S337 }),
  .Q({ datapath_adr_outreg_9 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_13_ (
  .C({ controller_clk }),
  .D({ S338 }),
  .Q({ datapath_adr_outreg_10 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_14_ (
  .C({ controller_clk }),
  .D({ S339 }),
  .Q({ datapath_adr_outreg_11 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_15_ (
  .C({ controller_clk }),
  .D({ S340 }),
  .Q({ datapath_adr_outreg_12 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_16_ (
  .C({ controller_clk }),
  .D({ S341 }),
  .Q({ datapath_adr_outreg_13 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_17_ (
  .C({ controller_clk }),
  .D({ S342 }),
  .Q({ datapath_adr_outreg_14 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_18_ (
  .C({ controller_clk }),
  .D({ S3 }),
  .Q({ datapath_adr_outreg_15 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_19_ (
  .C({ controller_clk }),
  .D({ S313 }),
  .Q({ datapath_instruction_0 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_20_ (
  .C({ controller_clk }),
  .D({ S314 }),
  .Q({ datapath_instruction_1 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_21_ (
  .C({ controller_clk }),
  .D({ S315 }),
  .Q({ datapath_instruction_2 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_22_ (
  .C({ controller_clk }),
  .D({ S316 }),
  .Q({ datapath_instruction_3 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_23_ (
  .C({ controller_clk }),
  .D({ S317 }),
  .Q({ controller_fib_0 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_24_ (
  .C({ controller_clk }),
  .D({ S318 }),
  .Q({ controller_fib_1 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_25_ (
  .C({ controller_clk }),
  .D({ S319 }),
  .Q({ controller_fib_2 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_26_ (
  .C({ controller_clk }),
  .D({ S320 }),
  .Q({ controller_fib_3 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_27_ (
  .C({ controller_clk }),
  .D({ S321 }),
  .Q({ controller_fib_4 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_28_ (
  .C({ controller_clk }),
  .D({ S322 }),
  .Q({ controller_216_B_0 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_29_ (
  .C({ controller_clk }),
  .D({ S323 }),
  .Q({ controller_opcode_2 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_30_ (
  .C({ controller_clk }),
  .D({ S324 }),
  .Q({ controller_opcode_3 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_31_ (
  .C({ controller_clk }),
  .D({ S325 }),
  .Q({ controller_opcode_4 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_32_ (
  .C({ controller_clk }),
  .D({ S326 }),
  .Q({ controller_opcode_5 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_33_ (
  .C({ controller_clk }),
  .D({ S327 }),
  .Q({ controller_opcode_6 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_34_ (
  .C({ controller_clk }),
  .D({ S2 }),
  .Q({ controller_opcode_7 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_35_ (
  .C({ controller_clk }),
  .D({ S282 }),
  .Q({ datapath_multdivunit_outmdu1_0 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_36_ (
  .C({ controller_clk }),
  .D({ S283 }),
  .Q({ datapath_multdivunit_outmdu1_1 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_37_ (
  .C({ controller_clk }),
  .D({ S284 }),
  .Q({ datapath_multdivunit_outmdu1_2 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_38_ (
  .C({ controller_clk }),
  .D({ S285 }),
  .Q({ datapath_multdivunit_outmdu1_3 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_39_ (
  .C({ controller_clk }),
  .D({ S286 }),
  .Q({ datapath_multdivunit_outmdu1_4 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_40_ (
  .C({ controller_clk }),
  .D({ S287 }),
  .Q({ datapath_multdivunit_outmdu1_5 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_41_ (
  .C({ controller_clk }),
  .D({ S288 }),
  .Q({ datapath_multdivunit_outmdu1_6 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_42_ (
  .C({ controller_clk }),
  .D({ S289 }),
  .Q({ datapath_multdivunit_outmdu1_7 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_43_ (
  .C({ controller_clk }),
  .D({ S290 }),
  .Q({ datapath_multdivunit_outmdu1_8 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_44_ (
  .C({ controller_clk }),
  .D({ S291 }),
  .Q({ datapath_multdivunit_outmdu1_9 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_45_ (
  .C({ controller_clk }),
  .D({ S292 }),
  .Q({ datapath_multdivunit_outmdu1_10 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_46_ (
  .C({ controller_clk }),
  .D({ S293 }),
  .Q({ datapath_multdivunit_outmdu1_11 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_47_ (
  .C({ controller_clk }),
  .D({ S294 }),
  .Q({ datapath_multdivunit_outmdu1_12 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_48_ (
  .C({ controller_clk }),
  .D({ S295 }),
  .Q({ datapath_multdivunit_outmdu1_13 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_49_ (
  .C({ controller_clk }),
  .D({ S296 }),
  .Q({ datapath_multdivunit_outmdu1_14 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_50_ (
  .C({ controller_clk }),
  .D({ S297 }),
  .Q({ datapath_multdivunit_outmdu1_15 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_51_ (
  .C({ controller_clk }),
  .D({ S298 }),
  .Q({ datapath_multdivunit_outmdu2_0 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_52_ (
  .C({ controller_clk }),
  .D({ S299 }),
  .Q({ datapath_multdivunit_outmdu2_1 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_53_ (
  .C({ controller_clk }),
  .D({ S300 }),
  .Q({ datapath_multdivunit_outmdu2_2 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_54_ (
  .C({ controller_clk }),
  .D({ S301 }),
  .Q({ datapath_multdivunit_outmdu2_3 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_55_ (
  .C({ controller_clk }),
  .D({ S302 }),
  .Q({ datapath_multdivunit_outmdu2_4 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_56_ (
  .C({ controller_clk }),
  .D({ S303 }),
  .Q({ datapath_multdivunit_outmdu2_5 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_57_ (
  .C({ controller_clk }),
  .D({ S304 }),
  .Q({ datapath_multdivunit_outmdu2_6 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_58_ (
  .C({ controller_clk }),
  .D({ S305 }),
  .Q({ datapath_multdivunit_outmdu2_7 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_59_ (
  .C({ controller_clk }),
  .D({ S306 }),
  .Q({ datapath_multdivunit_outmdu2_8 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_60_ (
  .C({ controller_clk }),
  .D({ S307 }),
  .Q({ datapath_multdivunit_outmdu2_9 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_61_ (
  .C({ controller_clk }),
  .D({ S308 }),
  .Q({ datapath_multdivunit_outmdu2_10 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_62_ (
  .C({ controller_clk }),
  .D({ S309 }),
  .Q({ datapath_multdivunit_outmdu2_11 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_63_ (
  .C({ controller_clk }),
  .D({ S310 }),
  .Q({ datapath_multdivunit_outmdu2_12 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_64_ (
  .C({ controller_clk }),
  .D({ S311 }),
  .Q({ datapath_multdivunit_outmdu2_13 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_65_ (
  .C({ controller_clk }),
  .D({ S312 }),
  .Q({ datapath_multdivunit_outmdu2_14 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_66_ (
  .C({ controller_clk }),
  .D({ S1 }),
  .Q({ datapath_multdivunit_outmdu2_15 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_67_ (
  .C({ controller_clk }),
  .D({ S267 }),
  .Q({ datapath_muxmem_in2_0 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_68_ (
  .C({ controller_clk }),
  .D({ S268 }),
  .Q({ datapath_muxmem_in2_1 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_69_ (
  .C({ controller_clk }),
  .D({ S269 }),
  .Q({ datapath_muxmem_in2_2 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_70_ (
  .C({ controller_clk }),
  .D({ S270 }),
  .Q({ datapath_muxmem_in2_3 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_71_ (
  .C({ controller_clk }),
  .D({ S271 }),
  .Q({ datapath_muxmem_in2_4 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_72_ (
  .C({ controller_clk }),
  .D({ S272 }),
  .Q({ datapath_muxmem_in2_5 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_73_ (
  .C({ controller_clk }),
  .D({ S273 }),
  .Q({ datapath_muxmem_in2_6 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_74_ (
  .C({ controller_clk }),
  .D({ S274 }),
  .Q({ datapath_muxmem_in2_7 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_75_ (
  .C({ controller_clk }),
  .D({ S275 }),
  .Q({ datapath_muxmem_in2_8 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_76_ (
  .C({ controller_clk }),
  .D({ S276 }),
  .Q({ datapath_muxmem_in2_9 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_77_ (
  .C({ controller_clk }),
  .D({ S277 }),
  .Q({ datapath_muxmem_in2_10 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_78_ (
  .C({ controller_clk }),
  .D({ S278 }),
  .Q({ datapath_muxmem_in2_11 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_79_ (
  .C({ controller_clk }),
  .D({ S279 }),
  .Q({ datapath_muxmem_in2_12 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_80_ (
  .C({ controller_clk }),
  .D({ S280 }),
  .Q({ datapath_muxmem_in2_13 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_81_ (
  .C({ controller_clk }),
  .D({ S281 }),
  .Q({ datapath_muxmem_in2_14 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_82_ (
  .C({ controller_clk }),
  .D({ S0 }),
  .Q({ datapath_muxmem_in2_15 }),
  .R({ controller_rst })
);
DFF_NP1 #() 
DFF_NP1_1_ (
  .C({ controller_clk }),
  .D({ S4 }),
  .Q({ datapath_theregisterfile_memtrf_64 }),
  .R({ controller_rst })
);
DFF_NP1 #() 
DFF_NP1_2_ (
  .C({ controller_clk }),
  .D({ S5 }),
  .Q({ datapath_theregisterfile_memtrf_65 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_1_ (
  .C({ controller_clk }),
  .D({ S6 }),
  .Q({ datapath_theregisterfile_memtrf_66 }),
  .R({ controller_rst })
);
DFF_NP1 #() 
DFF_NP1_3_ (
  .C({ controller_clk }),
  .D({ S7 }),
  .Q({ datapath_theregisterfile_memtrf_67 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_2_ (
  .C({ controller_clk }),
  .D({ S8 }),
  .Q({ datapath_theregisterfile_memtrf_68 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_3_ (
  .C({ controller_clk }),
  .D({ S9 }),
  .Q({ datapath_theregisterfile_memtrf_69 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_4_ (
  .C({ controller_clk }),
  .D({ S10 }),
  .Q({ datapath_theregisterfile_memtrf_70 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_5_ (
  .C({ controller_clk }),
  .D({ S11 }),
  .Q({ datapath_theregisterfile_memtrf_71 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_6_ (
  .C({ controller_clk }),
  .D({ S12 }),
  .Q({ datapath_theregisterfile_memtrf_72 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_7_ (
  .C({ controller_clk }),
  .D({ S13 }),
  .Q({ datapath_theregisterfile_memtrf_73 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_8_ (
  .C({ controller_clk }),
  .D({ S14 }),
  .Q({ datapath_theregisterfile_memtrf_74 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_9_ (
  .C({ controller_clk }),
  .D({ S15 }),
  .Q({ datapath_theregisterfile_memtrf_75 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_10_ (
  .C({ controller_clk }),
  .D({ S16 }),
  .Q({ datapath_theregisterfile_memtrf_76 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_11_ (
  .C({ controller_clk }),
  .D({ S17 }),
  .Q({ datapath_theregisterfile_memtrf_77 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_12_ (
  .C({ controller_clk }),
  .D({ S18 }),
  .Q({ datapath_theregisterfile_memtrf_78 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_13_ (
  .C({ controller_clk }),
  .D({ S19 }),
  .Q({ datapath_theregisterfile_memtrf_79 }),
  .R({ controller_rst })
);
DFF_NP1 #() 
DFF_NP1_4_ (
  .C({ controller_clk }),
  .D({ S20 }),
  .Q({ datapath_theregisterfile_memtrf_32 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_14_ (
  .C({ controller_clk }),
  .D({ S21 }),
  .Q({ datapath_theregisterfile_memtrf_33 }),
  .R({ controller_rst })
);
DFF_NP1 #() 
DFF_NP1_5_ (
  .C({ controller_clk }),
  .D({ S22 }),
  .Q({ datapath_theregisterfile_memtrf_34 }),
  .R({ controller_rst })
);
DFF_NP1 #() 
DFF_NP1_6_ (
  .C({ controller_clk }),
  .D({ S23 }),
  .Q({ datapath_theregisterfile_memtrf_35 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_15_ (
  .C({ controller_clk }),
  .D({ S24 }),
  .Q({ datapath_theregisterfile_memtrf_36 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_16_ (
  .C({ controller_clk }),
  .D({ S25 }),
  .Q({ datapath_theregisterfile_memtrf_37 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_17_ (
  .C({ controller_clk }),
  .D({ S26 }),
  .Q({ datapath_theregisterfile_memtrf_38 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_18_ (
  .C({ controller_clk }),
  .D({ S27 }),
  .Q({ datapath_theregisterfile_memtrf_39 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_19_ (
  .C({ controller_clk }),
  .D({ S28 }),
  .Q({ datapath_theregisterfile_memtrf_40 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_20_ (
  .C({ controller_clk }),
  .D({ S29 }),
  .Q({ datapath_theregisterfile_memtrf_41 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_21_ (
  .C({ controller_clk }),
  .D({ S30 }),
  .Q({ datapath_theregisterfile_memtrf_42 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_22_ (
  .C({ controller_clk }),
  .D({ S31 }),
  .Q({ datapath_theregisterfile_memtrf_43 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_23_ (
  .C({ controller_clk }),
  .D({ S32 }),
  .Q({ datapath_theregisterfile_memtrf_44 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_24_ (
  .C({ controller_clk }),
  .D({ S33 }),
  .Q({ datapath_theregisterfile_memtrf_45 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_25_ (
  .C({ controller_clk }),
  .D({ S34 }),
  .Q({ datapath_theregisterfile_memtrf_46 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_26_ (
  .C({ controller_clk }),
  .D({ S35 }),
  .Q({ datapath_theregisterfile_memtrf_47 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_27_ (
  .C({ controller_clk }),
  .D({ S36 }),
  .Q({ datapath_theregisterfile_memtrf_48 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_28_ (
  .C({ controller_clk }),
  .D({ S37 }),
  .Q({ datapath_theregisterfile_memtrf_49 }),
  .R({ controller_rst })
);
DFF_NP1 #() 
DFF_NP1_7_ (
  .C({ controller_clk }),
  .D({ S38 }),
  .Q({ datapath_theregisterfile_memtrf_50 }),
  .R({ controller_rst })
);
DFF_NP1 #() 
DFF_NP1_8_ (
  .C({ controller_clk }),
  .D({ S39 }),
  .Q({ datapath_theregisterfile_memtrf_51 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_29_ (
  .C({ controller_clk }),
  .D({ S40 }),
  .Q({ datapath_theregisterfile_memtrf_52 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_30_ (
  .C({ controller_clk }),
  .D({ S41 }),
  .Q({ datapath_theregisterfile_memtrf_53 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_31_ (
  .C({ controller_clk }),
  .D({ S42 }),
  .Q({ datapath_theregisterfile_memtrf_54 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_32_ (
  .C({ controller_clk }),
  .D({ S43 }),
  .Q({ datapath_theregisterfile_memtrf_55 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_33_ (
  .C({ controller_clk }),
  .D({ S44 }),
  .Q({ datapath_theregisterfile_memtrf_56 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_34_ (
  .C({ controller_clk }),
  .D({ S45 }),
  .Q({ datapath_theregisterfile_memtrf_57 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_35_ (
  .C({ controller_clk }),
  .D({ S46 }),
  .Q({ datapath_theregisterfile_memtrf_58 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_36_ (
  .C({ controller_clk }),
  .D({ S47 }),
  .Q({ datapath_theregisterfile_memtrf_59 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_37_ (
  .C({ controller_clk }),
  .D({ S48 }),
  .Q({ datapath_theregisterfile_memtrf_60 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_38_ (
  .C({ controller_clk }),
  .D({ S49 }),
  .Q({ datapath_theregisterfile_memtrf_61 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_39_ (
  .C({ controller_clk }),
  .D({ S50 }),
  .Q({ datapath_theregisterfile_memtrf_62 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_40_ (
  .C({ controller_clk }),
  .D({ S51 }),
  .Q({ datapath_theregisterfile_memtrf_63 }),
  .R({ controller_rst })
);
DFF_NP1 #() 
DFF_NP1_9_ (
  .C({ controller_clk }),
  .D({ S52 }),
  .Q({ datapath_theregisterfile_memtrf_128 }),
  .R({ controller_rst })
);
DFF_NP1 #() 
DFF_NP1_10_ (
  .C({ controller_clk }),
  .D({ S53 }),
  .Q({ datapath_theregisterfile_memtrf_129 }),
  .R({ controller_rst })
);
DFF_NP1 #() 
DFF_NP1_11_ (
  .C({ controller_clk }),
  .D({ S54 }),
  .Q({ datapath_theregisterfile_memtrf_130 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_41_ (
  .C({ controller_clk }),
  .D({ S55 }),
  .Q({ datapath_theregisterfile_memtrf_131 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_42_ (
  .C({ controller_clk }),
  .D({ S56 }),
  .Q({ datapath_theregisterfile_memtrf_132 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_43_ (
  .C({ controller_clk }),
  .D({ S57 }),
  .Q({ datapath_theregisterfile_memtrf_133 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_44_ (
  .C({ controller_clk }),
  .D({ S58 }),
  .Q({ datapath_theregisterfile_memtrf_134 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_45_ (
  .C({ controller_clk }),
  .D({ S59 }),
  .Q({ datapath_theregisterfile_memtrf_135 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_46_ (
  .C({ controller_clk }),
  .D({ S60 }),
  .Q({ datapath_theregisterfile_memtrf_136 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_47_ (
  .C({ controller_clk }),
  .D({ S61 }),
  .Q({ datapath_theregisterfile_memtrf_137 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_48_ (
  .C({ controller_clk }),
  .D({ S62 }),
  .Q({ datapath_theregisterfile_memtrf_138 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_49_ (
  .C({ controller_clk }),
  .D({ S63 }),
  .Q({ datapath_theregisterfile_memtrf_139 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_50_ (
  .C({ controller_clk }),
  .D({ S64 }),
  .Q({ datapath_theregisterfile_memtrf_140 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_51_ (
  .C({ controller_clk }),
  .D({ S65 }),
  .Q({ datapath_theregisterfile_memtrf_141 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_52_ (
  .C({ controller_clk }),
  .D({ S66 }),
  .Q({ datapath_theregisterfile_memtrf_142 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_53_ (
  .C({ controller_clk }),
  .D({ S67 }),
  .Q({ datapath_theregisterfile_memtrf_143 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_54_ (
  .C({ controller_clk }),
  .D({ S68 }),
  .Q({ datapath_theregisterfile_memtrf_16 }),
  .R({ controller_rst })
);
DFF_NP1 #() 
DFF_NP1_12_ (
  .C({ controller_clk }),
  .D({ S69 }),
  .Q({ datapath_theregisterfile_memtrf_17 }),
  .R({ controller_rst })
);
DFF_NP1 #() 
DFF_NP1_13_ (
  .C({ controller_clk }),
  .D({ S70 }),
  .Q({ datapath_theregisterfile_memtrf_18 }),
  .R({ controller_rst })
);
DFF_NP1 #() 
DFF_NP1_14_ (
  .C({ controller_clk }),
  .D({ S71 }),
  .Q({ datapath_theregisterfile_memtrf_19 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_55_ (
  .C({ controller_clk }),
  .D({ S72 }),
  .Q({ datapath_theregisterfile_memtrf_20 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_56_ (
  .C({ controller_clk }),
  .D({ S73 }),
  .Q({ datapath_theregisterfile_memtrf_21 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_57_ (
  .C({ controller_clk }),
  .D({ S74 }),
  .Q({ datapath_theregisterfile_memtrf_22 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_58_ (
  .C({ controller_clk }),
  .D({ S75 }),
  .Q({ datapath_theregisterfile_memtrf_23 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_59_ (
  .C({ controller_clk }),
  .D({ S76 }),
  .Q({ datapath_theregisterfile_memtrf_24 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_60_ (
  .C({ controller_clk }),
  .D({ S77 }),
  .Q({ datapath_theregisterfile_memtrf_25 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_61_ (
  .C({ controller_clk }),
  .D({ S78 }),
  .Q({ datapath_theregisterfile_memtrf_26 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_62_ (
  .C({ controller_clk }),
  .D({ S79 }),
  .Q({ datapath_theregisterfile_memtrf_27 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_63_ (
  .C({ controller_clk }),
  .D({ S80 }),
  .Q({ datapath_theregisterfile_memtrf_28 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_64_ (
  .C({ controller_clk }),
  .D({ S81 }),
  .Q({ datapath_theregisterfile_memtrf_29 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_65_ (
  .C({ controller_clk }),
  .D({ S82 }),
  .Q({ datapath_theregisterfile_memtrf_30 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_66_ (
  .C({ controller_clk }),
  .D({ S83 }),
  .Q({ datapath_theregisterfile_memtrf_31 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_67_ (
  .C({ controller_clk }),
  .D({ S84 }),
  .Q({ datapath_theregisterfile_memtrf_80 }),
  .R({ controller_rst })
);
DFF_NP1 #() 
DFF_NP1_15_ (
  .C({ controller_clk }),
  .D({ S85 }),
  .Q({ datapath_theregisterfile_memtrf_81 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_68_ (
  .C({ controller_clk }),
  .D({ S86 }),
  .Q({ datapath_theregisterfile_memtrf_82 }),
  .R({ controller_rst })
);
DFF_NP1 #() 
DFF_NP1_16_ (
  .C({ controller_clk }),
  .D({ S87 }),
  .Q({ datapath_theregisterfile_memtrf_83 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_69_ (
  .C({ controller_clk }),
  .D({ S88 }),
  .Q({ datapath_theregisterfile_memtrf_84 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_70_ (
  .C({ controller_clk }),
  .D({ S89 }),
  .Q({ datapath_theregisterfile_memtrf_85 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_71_ (
  .C({ controller_clk }),
  .D({ S90 }),
  .Q({ datapath_theregisterfile_memtrf_86 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_72_ (
  .C({ controller_clk }),
  .D({ S91 }),
  .Q({ datapath_theregisterfile_memtrf_87 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_73_ (
  .C({ controller_clk }),
  .D({ S92 }),
  .Q({ datapath_theregisterfile_memtrf_88 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_74_ (
  .C({ controller_clk }),
  .D({ S93 }),
  .Q({ datapath_theregisterfile_memtrf_89 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_75_ (
  .C({ controller_clk }),
  .D({ S94 }),
  .Q({ datapath_theregisterfile_memtrf_90 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_76_ (
  .C({ controller_clk }),
  .D({ S95 }),
  .Q({ datapath_theregisterfile_memtrf_91 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_77_ (
  .C({ controller_clk }),
  .D({ S96 }),
  .Q({ datapath_theregisterfile_memtrf_92 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_78_ (
  .C({ controller_clk }),
  .D({ S97 }),
  .Q({ datapath_theregisterfile_memtrf_93 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_79_ (
  .C({ controller_clk }),
  .D({ S98 }),
  .Q({ datapath_theregisterfile_memtrf_94 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_80_ (
  .C({ controller_clk }),
  .D({ S99 }),
  .Q({ datapath_theregisterfile_memtrf_95 }),
  .R({ controller_rst })
);
DFF_NP1 #() 
DFF_NP1_17_ (
  .C({ controller_clk }),
  .D({ S100 }),
  .Q({ datapath_theregisterfile_memtrf_96 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_81_ (
  .C({ controller_clk }),
  .D({ S101 }),
  .Q({ datapath_theregisterfile_memtrf_97 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_82_ (
  .C({ controller_clk }),
  .D({ S102 }),
  .Q({ datapath_theregisterfile_memtrf_98 }),
  .R({ controller_rst })
);
DFF_NP1 #() 
DFF_NP1_18_ (
  .C({ controller_clk }),
  .D({ S103 }),
  .Q({ datapath_theregisterfile_memtrf_99 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_83_ (
  .C({ controller_clk }),
  .D({ S104 }),
  .Q({ datapath_theregisterfile_memtrf_100 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_84_ (
  .C({ controller_clk }),
  .D({ S105 }),
  .Q({ datapath_theregisterfile_memtrf_101 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_85_ (
  .C({ controller_clk }),
  .D({ S106 }),
  .Q({ datapath_theregisterfile_memtrf_102 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_86_ (
  .C({ controller_clk }),
  .D({ S107 }),
  .Q({ datapath_theregisterfile_memtrf_103 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_87_ (
  .C({ controller_clk }),
  .D({ S108 }),
  .Q({ datapath_theregisterfile_memtrf_104 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_88_ (
  .C({ controller_clk }),
  .D({ S109 }),
  .Q({ datapath_theregisterfile_memtrf_105 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_89_ (
  .C({ controller_clk }),
  .D({ S110 }),
  .Q({ datapath_theregisterfile_memtrf_106 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_90_ (
  .C({ controller_clk }),
  .D({ S111 }),
  .Q({ datapath_theregisterfile_memtrf_107 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_91_ (
  .C({ controller_clk }),
  .D({ S112 }),
  .Q({ datapath_theregisterfile_memtrf_108 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_92_ (
  .C({ controller_clk }),
  .D({ S113 }),
  .Q({ datapath_theregisterfile_memtrf_109 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_93_ (
  .C({ controller_clk }),
  .D({ S114 }),
  .Q({ datapath_theregisterfile_memtrf_110 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_94_ (
  .C({ controller_clk }),
  .D({ S115 }),
  .Q({ datapath_theregisterfile_memtrf_111 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_95_ (
  .C({ controller_clk }),
  .D({ S116 }),
  .Q({ datapath_theregisterfile_memtrf_112 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_96_ (
  .C({ controller_clk }),
  .D({ S117 }),
  .Q({ datapath_theregisterfile_memtrf_113 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_97_ (
  .C({ controller_clk }),
  .D({ S118 }),
  .Q({ datapath_theregisterfile_memtrf_114 }),
  .R({ controller_rst })
);
DFF_NP1 #() 
DFF_NP1_19_ (
  .C({ controller_clk }),
  .D({ S119 }),
  .Q({ datapath_theregisterfile_memtrf_115 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_98_ (
  .C({ controller_clk }),
  .D({ S120 }),
  .Q({ datapath_theregisterfile_memtrf_116 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_99_ (
  .C({ controller_clk }),
  .D({ S121 }),
  .Q({ datapath_theregisterfile_memtrf_117 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_100_ (
  .C({ controller_clk }),
  .D({ S122 }),
  .Q({ datapath_theregisterfile_memtrf_118 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_101_ (
  .C({ controller_clk }),
  .D({ S123 }),
  .Q({ datapath_theregisterfile_memtrf_119 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_102_ (
  .C({ controller_clk }),
  .D({ S124 }),
  .Q({ datapath_theregisterfile_memtrf_120 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_103_ (
  .C({ controller_clk }),
  .D({ S125 }),
  .Q({ datapath_theregisterfile_memtrf_121 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_104_ (
  .C({ controller_clk }),
  .D({ S126 }),
  .Q({ datapath_theregisterfile_memtrf_122 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_105_ (
  .C({ controller_clk }),
  .D({ S127 }),
  .Q({ datapath_theregisterfile_memtrf_123 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_106_ (
  .C({ controller_clk }),
  .D({ S128 }),
  .Q({ datapath_theregisterfile_memtrf_124 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_107_ (
  .C({ controller_clk }),
  .D({ S129 }),
  .Q({ datapath_theregisterfile_memtrf_125 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_108_ (
  .C({ controller_clk }),
  .D({ S130 }),
  .Q({ datapath_theregisterfile_memtrf_126 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_109_ (
  .C({ controller_clk }),
  .D({ S131 }),
  .Q({ datapath_theregisterfile_memtrf_127 }),
  .R({ controller_rst })
);
DFF_NP1 #() 
DFF_NP1_20_ (
  .C({ controller_clk }),
  .D({ S132 }),
  .Q({ datapath_theregisterfile_memtrf_0 }),
  .R({ controller_rst })
);
DFF_NP1 #() 
DFF_NP1_21_ (
  .C({ controller_clk }),
  .D({ S133 }),
  .Q({ datapath_theregisterfile_memtrf_1 }),
  .R({ controller_rst })
);
DFF_NP1 #() 
DFF_NP1_22_ (
  .C({ controller_clk }),
  .D({ S134 }),
  .Q({ datapath_theregisterfile_memtrf_2 }),
  .R({ controller_rst })
);
DFF_NP1 #() 
DFF_NP1_23_ (
  .C({ controller_clk }),
  .D({ S135 }),
  .Q({ datapath_theregisterfile_memtrf_3 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_110_ (
  .C({ controller_clk }),
  .D({ S136 }),
  .Q({ datapath_theregisterfile_memtrf_4 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_111_ (
  .C({ controller_clk }),
  .D({ S137 }),
  .Q({ datapath_theregisterfile_memtrf_5 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_112_ (
  .C({ controller_clk }),
  .D({ S138 }),
  .Q({ datapath_theregisterfile_memtrf_6 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_113_ (
  .C({ controller_clk }),
  .D({ S139 }),
  .Q({ datapath_theregisterfile_memtrf_7 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_114_ (
  .C({ controller_clk }),
  .D({ S140 }),
  .Q({ datapath_theregisterfile_memtrf_8 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_115_ (
  .C({ controller_clk }),
  .D({ S141 }),
  .Q({ datapath_theregisterfile_memtrf_9 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_116_ (
  .C({ controller_clk }),
  .D({ S142 }),
  .Q({ datapath_theregisterfile_memtrf_10 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_117_ (
  .C({ controller_clk }),
  .D({ S143 }),
  .Q({ datapath_theregisterfile_memtrf_11 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_118_ (
  .C({ controller_clk }),
  .D({ S144 }),
  .Q({ datapath_theregisterfile_memtrf_12 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_119_ (
  .C({ controller_clk }),
  .D({ S145 }),
  .Q({ datapath_theregisterfile_memtrf_13 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_120_ (
  .C({ controller_clk }),
  .D({ S146 }),
  .Q({ datapath_theregisterfile_memtrf_14 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_121_ (
  .C({ controller_clk }),
  .D({ S147 }),
  .Q({ datapath_theregisterfile_memtrf_15 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_122_ (
  .C({ controller_clk }),
  .D({ S148 }),
  .Q({ datapath_theregisterfile_memtrf_144 }),
  .R({ controller_rst })
);
DFF_NP1 #() 
DFF_NP1_24_ (
  .C({ controller_clk }),
  .D({ S149 }),
  .Q({ datapath_theregisterfile_memtrf_145 }),
  .R({ controller_rst })
);
DFF_NP1 #() 
DFF_NP1_25_ (
  .C({ controller_clk }),
  .D({ S150 }),
  .Q({ datapath_theregisterfile_memtrf_146 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_123_ (
  .C({ controller_clk }),
  .D({ S151 }),
  .Q({ datapath_theregisterfile_memtrf_147 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_124_ (
  .C({ controller_clk }),
  .D({ S152 }),
  .Q({ datapath_theregisterfile_memtrf_148 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_125_ (
  .C({ controller_clk }),
  .D({ S153 }),
  .Q({ datapath_theregisterfile_memtrf_149 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_126_ (
  .C({ controller_clk }),
  .D({ S154 }),
  .Q({ datapath_theregisterfile_memtrf_150 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_127_ (
  .C({ controller_clk }),
  .D({ S155 }),
  .Q({ datapath_theregisterfile_memtrf_151 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_128_ (
  .C({ controller_clk }),
  .D({ S156 }),
  .Q({ datapath_theregisterfile_memtrf_152 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_129_ (
  .C({ controller_clk }),
  .D({ S157 }),
  .Q({ datapath_theregisterfile_memtrf_153 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_130_ (
  .C({ controller_clk }),
  .D({ S158 }),
  .Q({ datapath_theregisterfile_memtrf_154 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_131_ (
  .C({ controller_clk }),
  .D({ S159 }),
  .Q({ datapath_theregisterfile_memtrf_155 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_132_ (
  .C({ controller_clk }),
  .D({ S160 }),
  .Q({ datapath_theregisterfile_memtrf_156 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_133_ (
  .C({ controller_clk }),
  .D({ S161 }),
  .Q({ datapath_theregisterfile_memtrf_157 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_134_ (
  .C({ controller_clk }),
  .D({ S162 }),
  .Q({ datapath_theregisterfile_memtrf_158 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_135_ (
  .C({ controller_clk }),
  .D({ S163 }),
  .Q({ datapath_theregisterfile_memtrf_159 }),
  .R({ controller_rst })
);
DFF_NP1 #() 
DFF_NP1_26_ (
  .C({ controller_clk }),
  .D({ S164 }),
  .Q({ datapath_theregisterfile_memtrf_160 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_136_ (
  .C({ controller_clk }),
  .D({ S165 }),
  .Q({ datapath_theregisterfile_memtrf_161 }),
  .R({ controller_rst })
);
DFF_NP1 #() 
DFF_NP1_27_ (
  .C({ controller_clk }),
  .D({ S166 }),
  .Q({ datapath_theregisterfile_memtrf_162 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_137_ (
  .C({ controller_clk }),
  .D({ S167 }),
  .Q({ datapath_theregisterfile_memtrf_163 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_138_ (
  .C({ controller_clk }),
  .D({ S168 }),
  .Q({ datapath_theregisterfile_memtrf_164 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_139_ (
  .C({ controller_clk }),
  .D({ S169 }),
  .Q({ datapath_theregisterfile_memtrf_165 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_140_ (
  .C({ controller_clk }),
  .D({ S170 }),
  .Q({ datapath_theregisterfile_memtrf_166 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_141_ (
  .C({ controller_clk }),
  .D({ S171 }),
  .Q({ datapath_theregisterfile_memtrf_167 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_142_ (
  .C({ controller_clk }),
  .D({ S172 }),
  .Q({ datapath_theregisterfile_memtrf_168 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_143_ (
  .C({ controller_clk }),
  .D({ S173 }),
  .Q({ datapath_theregisterfile_memtrf_169 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_144_ (
  .C({ controller_clk }),
  .D({ S174 }),
  .Q({ datapath_theregisterfile_memtrf_170 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_145_ (
  .C({ controller_clk }),
  .D({ S175 }),
  .Q({ datapath_theregisterfile_memtrf_171 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_146_ (
  .C({ controller_clk }),
  .D({ S176 }),
  .Q({ datapath_theregisterfile_memtrf_172 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_147_ (
  .C({ controller_clk }),
  .D({ S177 }),
  .Q({ datapath_theregisterfile_memtrf_173 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_148_ (
  .C({ controller_clk }),
  .D({ S178 }),
  .Q({ datapath_theregisterfile_memtrf_174 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_149_ (
  .C({ controller_clk }),
  .D({ S179 }),
  .Q({ datapath_theregisterfile_memtrf_175 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_150_ (
  .C({ controller_clk }),
  .D({ S180 }),
  .Q({ datapath_theregisterfile_memtrf_176 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_151_ (
  .C({ controller_clk }),
  .D({ S181 }),
  .Q({ datapath_theregisterfile_memtrf_177 }),
  .R({ controller_rst })
);
DFF_NP1 #() 
DFF_NP1_28_ (
  .C({ controller_clk }),
  .D({ S182 }),
  .Q({ datapath_theregisterfile_memtrf_178 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_152_ (
  .C({ controller_clk }),
  .D({ S183 }),
  .Q({ datapath_theregisterfile_memtrf_179 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_153_ (
  .C({ controller_clk }),
  .D({ S184 }),
  .Q({ datapath_theregisterfile_memtrf_180 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_154_ (
  .C({ controller_clk }),
  .D({ S185 }),
  .Q({ datapath_theregisterfile_memtrf_181 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_155_ (
  .C({ controller_clk }),
  .D({ S186 }),
  .Q({ datapath_theregisterfile_memtrf_182 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_156_ (
  .C({ controller_clk }),
  .D({ S187 }),
  .Q({ datapath_theregisterfile_memtrf_183 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_157_ (
  .C({ controller_clk }),
  .D({ S188 }),
  .Q({ datapath_theregisterfile_memtrf_184 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_158_ (
  .C({ controller_clk }),
  .D({ S189 }),
  .Q({ datapath_theregisterfile_memtrf_185 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_159_ (
  .C({ controller_clk }),
  .D({ S190 }),
  .Q({ datapath_theregisterfile_memtrf_186 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_160_ (
  .C({ controller_clk }),
  .D({ S191 }),
  .Q({ datapath_theregisterfile_memtrf_187 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_161_ (
  .C({ controller_clk }),
  .D({ S192 }),
  .Q({ datapath_theregisterfile_memtrf_188 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_162_ (
  .C({ controller_clk }),
  .D({ S193 }),
  .Q({ datapath_theregisterfile_memtrf_189 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_163_ (
  .C({ controller_clk }),
  .D({ S194 }),
  .Q({ datapath_theregisterfile_memtrf_190 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_164_ (
  .C({ controller_clk }),
  .D({ S195 }),
  .Q({ datapath_theregisterfile_memtrf_191 }),
  .R({ controller_rst })
);
DFF_NP1 #() 
DFF_NP1_29_ (
  .C({ controller_clk }),
  .D({ S196 }),
  .Q({ datapath_theregisterfile_memtrf_192 }),
  .R({ controller_rst })
);
DFF_NP1 #() 
DFF_NP1_30_ (
  .C({ controller_clk }),
  .D({ S197 }),
  .Q({ datapath_theregisterfile_memtrf_193 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_165_ (
  .C({ controller_clk }),
  .D({ S198 }),
  .Q({ datapath_theregisterfile_memtrf_194 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_166_ (
  .C({ controller_clk }),
  .D({ S199 }),
  .Q({ datapath_theregisterfile_memtrf_195 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_167_ (
  .C({ controller_clk }),
  .D({ S200 }),
  .Q({ datapath_theregisterfile_memtrf_196 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_168_ (
  .C({ controller_clk }),
  .D({ S201 }),
  .Q({ datapath_theregisterfile_memtrf_197 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_169_ (
  .C({ controller_clk }),
  .D({ S202 }),
  .Q({ datapath_theregisterfile_memtrf_198 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_170_ (
  .C({ controller_clk }),
  .D({ S203 }),
  .Q({ datapath_theregisterfile_memtrf_199 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_171_ (
  .C({ controller_clk }),
  .D({ S204 }),
  .Q({ datapath_theregisterfile_memtrf_200 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_172_ (
  .C({ controller_clk }),
  .D({ S205 }),
  .Q({ datapath_theregisterfile_memtrf_201 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_173_ (
  .C({ controller_clk }),
  .D({ S206 }),
  .Q({ datapath_theregisterfile_memtrf_202 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_174_ (
  .C({ controller_clk }),
  .D({ S207 }),
  .Q({ datapath_theregisterfile_memtrf_203 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_175_ (
  .C({ controller_clk }),
  .D({ S208 }),
  .Q({ datapath_theregisterfile_memtrf_204 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_176_ (
  .C({ controller_clk }),
  .D({ S209 }),
  .Q({ datapath_theregisterfile_memtrf_205 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_177_ (
  .C({ controller_clk }),
  .D({ S210 }),
  .Q({ datapath_theregisterfile_memtrf_206 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_178_ (
  .C({ controller_clk }),
  .D({ S211 }),
  .Q({ datapath_theregisterfile_memtrf_207 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_179_ (
  .C({ controller_clk }),
  .D({ S212 }),
  .Q({ datapath_theregisterfile_memtrf_208 }),
  .R({ controller_rst })
);
DFF_NP1 #() 
DFF_NP1_31_ (
  .C({ controller_clk }),
  .D({ S213 }),
  .Q({ datapath_theregisterfile_memtrf_209 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_180_ (
  .C({ controller_clk }),
  .D({ S214 }),
  .Q({ datapath_theregisterfile_memtrf_210 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_181_ (
  .C({ controller_clk }),
  .D({ S215 }),
  .Q({ datapath_theregisterfile_memtrf_211 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_182_ (
  .C({ controller_clk }),
  .D({ S216 }),
  .Q({ datapath_theregisterfile_memtrf_212 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_183_ (
  .C({ controller_clk }),
  .D({ S217 }),
  .Q({ datapath_theregisterfile_memtrf_213 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_184_ (
  .C({ controller_clk }),
  .D({ S218 }),
  .Q({ datapath_theregisterfile_memtrf_214 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_185_ (
  .C({ controller_clk }),
  .D({ S219 }),
  .Q({ datapath_theregisterfile_memtrf_215 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_186_ (
  .C({ controller_clk }),
  .D({ S220 }),
  .Q({ datapath_theregisterfile_memtrf_216 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_187_ (
  .C({ controller_clk }),
  .D({ S221 }),
  .Q({ datapath_theregisterfile_memtrf_217 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_188_ (
  .C({ controller_clk }),
  .D({ S222 }),
  .Q({ datapath_theregisterfile_memtrf_218 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_189_ (
  .C({ controller_clk }),
  .D({ S223 }),
  .Q({ datapath_theregisterfile_memtrf_219 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_190_ (
  .C({ controller_clk }),
  .D({ S224 }),
  .Q({ datapath_theregisterfile_memtrf_220 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_191_ (
  .C({ controller_clk }),
  .D({ S225 }),
  .Q({ datapath_theregisterfile_memtrf_221 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_192_ (
  .C({ controller_clk }),
  .D({ S226 }),
  .Q({ datapath_theregisterfile_memtrf_222 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_193_ (
  .C({ controller_clk }),
  .D({ S227 }),
  .Q({ datapath_theregisterfile_memtrf_223 }),
  .R({ controller_rst })
);
DFF_NP1 #() 
DFF_NP1_32_ (
  .C({ controller_clk }),
  .D({ S228 }),
  .Q({ datapath_theregisterfile_memtrf_224 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_194_ (
  .C({ controller_clk }),
  .D({ S229 }),
  .Q({ datapath_theregisterfile_memtrf_225 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_195_ (
  .C({ controller_clk }),
  .D({ S230 }),
  .Q({ datapath_theregisterfile_memtrf_226 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_196_ (
  .C({ controller_clk }),
  .D({ S231 }),
  .Q({ datapath_theregisterfile_memtrf_227 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_197_ (
  .C({ controller_clk }),
  .D({ S232 }),
  .Q({ datapath_theregisterfile_memtrf_228 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_198_ (
  .C({ controller_clk }),
  .D({ S233 }),
  .Q({ datapath_theregisterfile_memtrf_229 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_199_ (
  .C({ controller_clk }),
  .D({ S234 }),
  .Q({ datapath_theregisterfile_memtrf_230 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_200_ (
  .C({ controller_clk }),
  .D({ S235 }),
  .Q({ datapath_theregisterfile_memtrf_231 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_201_ (
  .C({ controller_clk }),
  .D({ S236 }),
  .Q({ datapath_theregisterfile_memtrf_232 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_202_ (
  .C({ controller_clk }),
  .D({ S237 }),
  .Q({ datapath_theregisterfile_memtrf_233 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_203_ (
  .C({ controller_clk }),
  .D({ S238 }),
  .Q({ datapath_theregisterfile_memtrf_234 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_204_ (
  .C({ controller_clk }),
  .D({ S239 }),
  .Q({ datapath_theregisterfile_memtrf_235 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_205_ (
  .C({ controller_clk }),
  .D({ S240 }),
  .Q({ datapath_theregisterfile_memtrf_236 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_206_ (
  .C({ controller_clk }),
  .D({ S241 }),
  .Q({ datapath_theregisterfile_memtrf_237 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_207_ (
  .C({ controller_clk }),
  .D({ S242 }),
  .Q({ datapath_theregisterfile_memtrf_238 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_208_ (
  .C({ controller_clk }),
  .D({ S243 }),
  .Q({ datapath_theregisterfile_memtrf_239 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_209_ (
  .C({ controller_clk }),
  .D({ S244 }),
  .Q({ datapath_theregisterfile_memtrf_240 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_210_ (
  .C({ controller_clk }),
  .D({ S245 }),
  .Q({ datapath_theregisterfile_memtrf_241 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_211_ (
  .C({ controller_clk }),
  .D({ S246 }),
  .Q({ datapath_theregisterfile_memtrf_242 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_212_ (
  .C({ controller_clk }),
  .D({ S247 }),
  .Q({ datapath_theregisterfile_memtrf_243 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_213_ (
  .C({ controller_clk }),
  .D({ S248 }),
  .Q({ datapath_theregisterfile_memtrf_244 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_214_ (
  .C({ controller_clk }),
  .D({ S249 }),
  .Q({ datapath_theregisterfile_memtrf_245 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_215_ (
  .C({ controller_clk }),
  .D({ S250 }),
  .Q({ datapath_theregisterfile_memtrf_246 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_216_ (
  .C({ controller_clk }),
  .D({ S251 }),
  .Q({ datapath_theregisterfile_memtrf_247 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_217_ (
  .C({ controller_clk }),
  .D({ S252 }),
  .Q({ datapath_theregisterfile_memtrf_248 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_218_ (
  .C({ controller_clk }),
  .D({ S253 }),
  .Q({ datapath_theregisterfile_memtrf_249 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_219_ (
  .C({ controller_clk }),
  .D({ S254 }),
  .Q({ datapath_theregisterfile_memtrf_250 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_220_ (
  .C({ controller_clk }),
  .D({ S255 }),
  .Q({ datapath_theregisterfile_memtrf_251 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_221_ (
  .C({ controller_clk }),
  .D({ S256 }),
  .Q({ datapath_theregisterfile_memtrf_252 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_222_ (
  .C({ controller_clk }),
  .D({ S257 }),
  .Q({ datapath_theregisterfile_memtrf_253 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_223_ (
  .C({ controller_clk }),
  .D({ S258 }),
  .Q({ datapath_theregisterfile_memtrf_254 }),
  .R({ controller_rst })
);
DFF_NP0 #() 
DFF_NP0_224_ (
  .C({ controller_clk }),
  .D({ S259 }),
  .Q({ datapath_theregisterfile_memtrf_255 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_83_ (
  .C({ controller_clk }),
  .D({ S260 }),
  .Q({ controller_outflag_0 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_84_ (
  .C({ controller_clk }),
  .D({ S261 }),
  .Q({ controller_outflag_1 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_85_ (
  .C({ controller_clk }),
  .D({ S262 }),
  .Q({ controller_outflag_2 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_86_ (
  .C({ controller_clk }),
  .D({ S263 }),
  .Q({ controller_outflag_3 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_87_ (
  .C({ controller_clk }),
  .D({ S264 }),
  .Q({ controller_389_B_0 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_88_ (
  .C({ controller_clk }),
  .D({ S265 }),
  .Q({ controller_389_B_2 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_89_ (
  .C({ controller_clk }),
  .D({ S266 }),
  .Q({ controller_outflag_6 }),
  .R({ controller_rst })
);
DFF_PP0 #() 
DFF_PP0_90_ (
  .C({ controller_clk }),
  .D({ S343 }),
  .Q({ controller_outflag_7 }),
  .R({ controller_rst })
);
OBUF #() 
OBUF_1_ (
  .I({ datapath_muxmem_in2_0 }),
  .O({ PCout[0] })
);
OBUF #() 
OBUF_2_ (
  .I({ datapath_muxmem_in2_1 }),
  .O({ PCout[1] })
);
OBUF #() 
OBUF_3_ (
  .I({ datapath_muxmem_in2_10 }),
  .O({ PCout[10] })
);
OBUF #() 
OBUF_4_ (
  .I({ datapath_muxmem_in2_11 }),
  .O({ PCout[11] })
);
OBUF #() 
OBUF_5_ (
  .I({ datapath_muxmem_in2_12 }),
  .O({ PCout[12] })
);
OBUF #() 
OBUF_6_ (
  .I({ datapath_muxmem_in2_13 }),
  .O({ PCout[13] })
);
OBUF #() 
OBUF_7_ (
  .I({ datapath_muxmem_in2_14 }),
  .O({ PCout[14] })
);
OBUF #() 
OBUF_8_ (
  .I({ datapath_muxmem_in2_15 }),
  .O({ PCout[15] })
);
OBUF #() 
OBUF_9_ (
  .I({ datapath_muxmem_in2_2 }),
  .O({ PCout[2] })
);
OBUF #() 
OBUF_10_ (
  .I({ datapath_muxmem_in2_3 }),
  .O({ PCout[3] })
);
OBUF #() 
OBUF_11_ (
  .I({ datapath_muxmem_in2_4 }),
  .O({ PCout[4] })
);
OBUF #() 
OBUF_12_ (
  .I({ datapath_muxmem_in2_5 }),
  .O({ PCout[5] })
);
OBUF #() 
OBUF_13_ (
  .I({ datapath_muxmem_in2_6 }),
  .O({ PCout[6] })
);
OBUF #() 
OBUF_14_ (
  .I({ datapath_muxmem_in2_7 }),
  .O({ PCout[7] })
);
OBUF #() 
OBUF_15_ (
  .I({ datapath_muxmem_in2_8 }),
  .O({ PCout[8] })
);
OBUF #() 
OBUF_16_ (
  .I({ datapath_muxmem_in2_9 }),
  .O({ PCout[9] })
);
OBUF #() 
OBUF_17_ (
  .I({ datapath_addrbus_0 }),
  .O({ addrBus[0] })
);
OBUF #() 
OBUF_18_ (
  .I({ datapath_addrbus_1 }),
  .O({ addrBus[1] })
);
OBUF #() 
OBUF_19_ (
  .I({ datapath_addrbus_10 }),
  .O({ addrBus[10] })
);
OBUF #() 
OBUF_20_ (
  .I({ datapath_addrbus_11 }),
  .O({ addrBus[11] })
);
OBUF #() 
OBUF_21_ (
  .I({ datapath_addrbus_12 }),
  .O({ addrBus[12] })
);
OBUF #() 
OBUF_22_ (
  .I({ datapath_addrbus_13 }),
  .O({ addrBus[13] })
);
OBUF #() 
OBUF_23_ (
  .I({ datapath_addrbus_14 }),
  .O({ addrBus[14] })
);
OBUF #() 
OBUF_24_ (
  .I({ datapath_addrbus_15 }),
  .O({ addrBus[15] })
);
OBUF #() 
OBUF_25_ (
  .I({ datapath_addrbus_2 }),
  .O({ addrBus[2] })
);
OBUF #() 
OBUF_26_ (
  .I({ datapath_addrbus_3 }),
  .O({ addrBus[3] })
);
OBUF #() 
OBUF_27_ (
  .I({ datapath_addrbus_4 }),
  .O({ addrBus[4] })
);
OBUF #() 
OBUF_28_ (
  .I({ datapath_addrbus_5 }),
  .O({ addrBus[5] })
);
OBUF #() 
OBUF_29_ (
  .I({ datapath_addrbus_6 }),
  .O({ addrBus[6] })
);
OBUF #() 
OBUF_30_ (
  .I({ datapath_addrbus_7 }),
  .O({ addrBus[7] })
);
OBUF #() 
OBUF_31_ (
  .I({ datapath_addrbus_8 }),
  .O({ addrBus[8] })
);
OBUF #() 
OBUF_32_ (
  .I({ datapath_addrbus_9 }),
  .O({ addrBus[9] })
);
IBUF #() 
IBUF_1_ (
  .I({ clk }),
  .O({ controller_clk })
);
IBUF #() 
IBUF_2_ (
  .I({ dataBusIn[0] }),
  .O({ datapath_databusin_0 })
);
IBUF #() 
IBUF_3_ (
  .I({ dataBusIn[1] }),
  .O({ datapath_databusin_1 })
);
IBUF #() 
IBUF_4_ (
  .I({ dataBusIn[10] }),
  .O({ datapath_databusin_10 })
);
IBUF #() 
IBUF_5_ (
  .I({ dataBusIn[11] }),
  .O({ datapath_databusin_11 })
);
IBUF #() 
IBUF_6_ (
  .I({ dataBusIn[12] }),
  .O({ datapath_databusin_12 })
);
IBUF #() 
IBUF_7_ (
  .I({ dataBusIn[13] }),
  .O({ datapath_databusin_13 })
);
IBUF #() 
IBUF_8_ (
  .I({ dataBusIn[14] }),
  .O({ datapath_databusin_14 })
);
IBUF #() 
IBUF_9_ (
  .I({ dataBusIn[15] }),
  .O({ datapath_databusin_15 })
);
IBUF #() 
IBUF_10_ (
  .I({ dataBusIn[2] }),
  .O({ datapath_databusin_2 })
);
IBUF #() 
IBUF_11_ (
  .I({ dataBusIn[3] }),
  .O({ datapath_databusin_3 })
);
IBUF #() 
IBUF_12_ (
  .I({ dataBusIn[4] }),
  .O({ datapath_databusin_4 })
);
IBUF #() 
IBUF_13_ (
  .I({ dataBusIn[5] }),
  .O({ datapath_databusin_5 })
);
IBUF #() 
IBUF_14_ (
  .I({ dataBusIn[6] }),
  .O({ datapath_databusin_6 })
);
IBUF #() 
IBUF_15_ (
  .I({ dataBusIn[7] }),
  .O({ datapath_databusin_7 })
);
IBUF #() 
IBUF_16_ (
  .I({ dataBusIn[8] }),
  .O({ datapath_databusin_8 })
);
IBUF #() 
IBUF_17_ (
  .I({ dataBusIn[9] }),
  .O({ datapath_databusin_9 })
);
OBUF #() 
OBUF_33_ (
  .I({ datapath_addsubunit_in1_0 }),
  .O({ dataBusOut[0] })
);
OBUF #() 
OBUF_34_ (
  .I({ datapath_addsubunit_in1_1 }),
  .O({ dataBusOut[1] })
);
OBUF #() 
OBUF_35_ (
  .I({ datapath_addsubunit_in1_10 }),
  .O({ dataBusOut[10] })
);
OBUF #() 
OBUF_36_ (
  .I({ datapath_addsubunit_in1_11 }),
  .O({ dataBusOut[11] })
);
OBUF #() 
OBUF_37_ (
  .I({ datapath_addsubunit_in1_12 }),
  .O({ dataBusOut[12] })
);
OBUF #() 
OBUF_38_ (
  .I({ datapath_addsubunit_in1_13 }),
  .O({ dataBusOut[13] })
);
OBUF #() 
OBUF_39_ (
  .I({ datapath_addsubunit_in1_14 }),
  .O({ dataBusOut[14] })
);
OBUF #() 
OBUF_40_ (
  .I({ datapath_addsubunit_in1_15 }),
  .O({ dataBusOut[15] })
);
OBUF #() 
OBUF_41_ (
  .I({ datapath_addsubunit_in1_2 }),
  .O({ dataBusOut[2] })
);
OBUF #() 
OBUF_42_ (
  .I({ datapath_addsubunit_in1_3 }),
  .O({ dataBusOut[3] })
);
OBUF #() 
OBUF_43_ (
  .I({ datapath_addsubunit_in1_4 }),
  .O({ dataBusOut[4] })
);
OBUF #() 
OBUF_44_ (
  .I({ datapath_addsubunit_in1_5 }),
  .O({ dataBusOut[5] })
);
OBUF #() 
OBUF_45_ (
  .I({ datapath_addsubunit_in1_6 }),
  .O({ dataBusOut[6] })
);
OBUF #() 
OBUF_46_ (
  .I({ datapath_addsubunit_in1_7 }),
  .O({ dataBusOut[7] })
);
OBUF #() 
OBUF_47_ (
  .I({ datapath_addsubunit_in1_8 }),
  .O({ dataBusOut[8] })
);
OBUF #() 
OBUF_48_ (
  .I({ datapath_addsubunit_in1_9 }),
  .O({ dataBusOut[9] })
);
OBUF #() 
OBUF_49_ (
  .I({ controller_readio }),
  .O({ readIO })
);
OBUF #() 
OBUF_50_ (
  .I({ controller_1115_S_0 }),
  .O({ readInst })
);
OBUF #() 
OBUF_51_ (
  .I({ controller_readmem }),
  .O({ readMEM })
);
IBUF #() 
IBUF_18_ (
  .I({ readyMEM }),
  .O({ controller_readymem })
);
IBUF #() 
IBUF_19_ (
  .I({ rst }),
  .O({ controller_rst })
);
OBUF #() 
OBUF_52_ (
  .I({ controller_writeio }),
  .O({ writeIO })
);
OBUF #() 
OBUF_53_ (
  .I({ controller_writemem }),
  .O({ writeMEM })
);

endmodule