module counter(clk, rst, en, co, counter);

wire S0;
wire S1;
wire S2;
wire S3;
wire S4;
wire S5;
wire S6;
wire S7;
wire S8;
wire S9;
wire S10;
wire S11;
wire S12;
wire S13;
wire S14;
wire S15;
wire S16;
wire S17;
wire S18;
wire S19;
wire S20;
wire S21;
wire S22;
wire S23;
wire S24;
wire S25;
wire new_counter_reg_0;
wire new_counter_reg_1;
wire new_counter_reg_2;
wire new_counter_reg_3;
input clk;
input rst;
input en;
output co;
output [3:0] counter;
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_0_ (
  .in1({ new_counter_reg_0 }),
  .out1({ S4 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1_ (
  .in1({ new_counter_reg_3 }),
  .out1({ S5 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2_ (
  .in1({ S20 }),
  .out1({ S6 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3_ (
  .in1({ new_counter_reg_1, new_counter_reg_0 }),
  .out1({ S7 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4_ (
  .in1({ new_counter_reg_2, new_counter_reg_3 }),
  .out1({ S8 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5_ (
  .in1({ S8, S7 }),
  .out1({ S19 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6_ (
  .in1({ S6, S4 }),
  .out1({ S9 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_7_ (
  .in1({ S20, new_counter_reg_0 }),
  .out1({ S10 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_8_ (
  .in1({ S10, S9 }),
  .out1({ S0 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_9_ (
  .in1({ S7, S6 }),
  .out1({ S11 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_10_ (
  .in1({ S9, new_counter_reg_1 }),
  .out1({ S12 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_11_ (
  .in1({ S12, S11 }),
  .out1({ S1 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_12_ (
  .in1({ S11, new_counter_reg_2 }),
  .out1({ S13 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_13_ (
  .in1({ S13 }),
  .out1({ S14 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_14_ (
  .in1({ S11, new_counter_reg_2 }),
  .out1({ S15 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_15_ (
  .in1({ S15, S14 }),
  .out1({ S2 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_16_ (
  .in1({ S14, new_counter_reg_3 }),
  .out1({ S16 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_17_ (
  .in1({ S13, S5 }),
  .out1({ S17 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_18_ (
  .in1({ S17, S16 }),
  .out1({ S3 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_19_ (
  .C({ S18 }),
  .CE({ 1'b1 }),
  .CLR({ S21 }),
  .D({ S0 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_counter_reg_0 }),
  .Si({ S22 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_20_ (
  .C({ S18 }),
  .CE({ 1'b1 }),
  .CLR({ S21 }),
  .D({ S1 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_counter_reg_1 }),
  .Si({ S23 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_21_ (
  .C({ S18 }),
  .CE({ 1'b1 }),
  .CLR({ S21 }),
  .D({ S2 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_counter_reg_2 }),
  .Si({ S24 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_22_ (
  .C({ S18 }),
  .CE({ 1'b1 }),
  .CLR({ S21 }),
  .D({ S3 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_counter_reg_3 }),
  .Si({ S25 }),
  .global_reset({ 1'b0 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_23_ (
  .in1({ clk }),
  .out1({ S18 })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_24_ (
  .in1({ S19 }),
  .out1({ co })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_25_ (
  .in1({ new_counter_reg_0 }),
  .out1({ counter[0] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_26_ (
  .in1({ new_counter_reg_1 }),
  .out1({ counter[1] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_27_ (
  .in1({ new_counter_reg_2 }),
  .out1({ counter[2] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_28_ (
  .in1({ new_counter_reg_3 }),
  .out1({ counter[3] })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_29_ (
  .in1({ en }),
  .out1({ S20 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_30_ (
  .in1({ rst }),
  .out1({ S21 })
);

endmodule