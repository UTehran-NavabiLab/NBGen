module PUNEH_Top(clk, rst, writeMEM, readMEM, dataBus_in, dataBus_out, addrBus);

wire S0;
wire S1;
wire S2;
wire S3;
wire S4;
wire S5;
wire S6;
wire S7;
wire S8;
wire S9;
wire S10;
wire S11;
wire S12;
wire S13;
wire S14;
wire S15;
wire S16;
wire S17;
wire S18;
wire S19;
wire S20;
wire S21;
wire S22;
wire S23;
wire S24;
wire S25;
wire S26;
wire S27;
wire S28;
wire S29;
wire S30;
wire S31;
wire S32;
wire S33;
wire S34;
wire S35;
wire S36;
wire S37;
wire S38;
wire S39;
wire S40;
wire S41;
wire S42;
wire S43;
wire S44;
wire S45;
wire S46;
wire S47;
wire S48;
wire S49;
wire S50;
wire S51;
wire S52;
wire S53;
wire S54;
wire S55;
wire S56;
wire S57;
wire S58;
wire S59;
wire S60;
wire S61;
wire S62;
wire S63;
wire S64;
wire S65;
wire S66;
wire S67;
wire S68;
wire S69;
wire S70;
wire S71;
wire S72;
wire S73;
wire S74;
wire S75;
wire S76;
wire S77;
wire S78;
wire S79;
wire S80;
wire S81;
wire S82;
wire S83;
wire S84;
wire S85;
wire S86;
wire S87;
wire S88;
wire S89;
wire S90;
wire S91;
wire S92;
wire S93;
wire S94;
wire S95;
wire S96;
wire S97;
wire S98;
wire S99;
wire S100;
wire S101;
wire S102;
wire S103;
wire S104;
wire S105;
wire S106;
wire S107;
wire S108;
wire S109;
wire S110;
wire S111;
wire S112;
wire S113;
wire S114;
wire S115;
wire S116;
wire S117;
wire S118;
wire S119;
wire S120;
wire S121;
wire S122;
wire S123;
wire S124;
wire S125;
wire S126;
wire S127;
wire S128;
wire S129;
wire S130;
wire S131;
wire S132;
wire S133;
wire S134;
wire S135;
wire S136;
wire S137;
wire S138;
wire S139;
wire S140;
wire S141;
wire S142;
wire S143;
wire S144;
wire S145;
wire S146;
wire S147;
wire S148;
wire S149;
wire S150;
wire S151;
wire S152;
wire S153;
wire S154;
wire S155;
wire S156;
wire S157;
wire S158;
wire S159;
wire S160;
wire S161;
wire S162;
wire S163;
wire S164;
wire S165;
wire S166;
wire S167;
wire S168;
wire S169;
wire S170;
wire S171;
wire S172;
wire S173;
wire S174;
wire S175;
wire S176;
wire S177;
wire S178;
wire S179;
wire S180;
wire S181;
wire S182;
wire S183;
wire S184;
wire S185;
wire S186;
wire S187;
wire S188;
wire S189;
wire S190;
wire S191;
wire S192;
wire S193;
wire S194;
wire S195;
wire S196;
wire S197;
wire S198;
wire S199;
wire S200;
wire S201;
wire S202;
wire S203;
wire S204;
wire S205;
wire S206;
wire S207;
wire S208;
wire S209;
wire S210;
wire S211;
wire S212;
wire S213;
wire S214;
wire S215;
wire S216;
wire S217;
wire S218;
wire S219;
wire S220;
wire S221;
wire S222;
wire S223;
wire S224;
wire S225;
wire S226;
wire S227;
wire S228;
wire S229;
wire S230;
wire S231;
wire S232;
wire S233;
wire S234;
wire S235;
wire S236;
wire S237;
wire S238;
wire S239;
wire S240;
wire S241;
wire S242;
wire S243;
wire S244;
wire S245;
wire S246;
wire S247;
wire S248;
wire S249;
wire S250;
wire S251;
wire S252;
wire S253;
wire S254;
wire S255;
wire S256;
wire S257;
wire S258;
wire S259;
wire S260;
wire S261;
wire S262;
wire S263;
wire S264;
wire S265;
wire S266;
wire S267;
wire S268;
wire S269;
wire S270;
wire S271;
wire S272;
wire S273;
wire S274;
wire S275;
wire S276;
wire S277;
wire S278;
wire S279;
wire S280;
wire S281;
wire S282;
wire S283;
wire S284;
wire S285;
wire S286;
wire S287;
wire S288;
wire S289;
wire S290;
wire S291;
wire S292;
wire S293;
wire S294;
wire S295;
wire S296;
wire S297;
wire S298;
wire S299;
wire S300;
wire S301;
wire S302;
wire S303;
wire S304;
wire S305;
wire S306;
wire S307;
wire S308;
wire S309;
wire S310;
wire S311;
wire S312;
wire S313;
wire S314;
wire S315;
wire S316;
wire S317;
wire S318;
wire S319;
wire S320;
wire S321;
wire S322;
wire S323;
wire S324;
wire S325;
wire S326;
wire S327;
wire S328;
wire S329;
wire S330;
wire S331;
wire S332;
wire S333;
wire S334;
wire S335;
wire S336;
wire S337;
wire S338;
wire S339;
wire S340;
wire S341;
wire S342;
wire S343;
wire S344;
wire S345;
wire S346;
wire S347;
wire S348;
wire S349;
wire S350;
wire S351;
wire S352;
wire S353;
wire S354;
wire S355;
wire S356;
wire S357;
wire S358;
wire S359;
wire S360;
wire S361;
wire S362;
wire S363;
wire S364;
wire S365;
wire S366;
wire S367;
wire S368;
wire S369;
wire S370;
wire S371;
wire S372;
wire S373;
wire S374;
wire S375;
wire S376;
wire S377;
wire S378;
wire S379;
wire S380;
wire S381;
wire S382;
wire S383;
wire S384;
wire S385;
wire S386;
wire S387;
wire S388;
wire S389;
wire S390;
wire S391;
wire S392;
wire S393;
wire S394;
wire S395;
wire S396;
wire S397;
wire S398;
wire S399;
wire S400;
wire S401;
wire S402;
wire S403;
wire S404;
wire S405;
wire S406;
wire S407;
wire S408;
wire S409;
wire S410;
wire S411;
wire S412;
wire S413;
wire S414;
wire S415;
wire S416;
wire S417;
wire S418;
wire S419;
wire S420;
wire S421;
wire S422;
wire S423;
wire S424;
wire S425;
wire S426;
wire S427;
wire S428;
wire S429;
wire S430;
wire S431;
wire S432;
wire S433;
wire S434;
wire S435;
wire S436;
wire S437;
wire S438;
wire S439;
wire S440;
wire S441;
wire S442;
wire S443;
wire S444;
wire S445;
wire S446;
wire S447;
wire S448;
wire S449;
wire S450;
wire S451;
wire S452;
wire S453;
wire S454;
wire S455;
wire S456;
wire S457;
wire S458;
wire S459;
wire S460;
wire S461;
wire S462;
wire S463;
wire S464;
wire S465;
wire S466;
wire S467;
wire S468;
wire S469;
wire S470;
wire S471;
wire S472;
wire S473;
wire S474;
wire S475;
wire S476;
wire S477;
wire S478;
wire S479;
wire S480;
wire S481;
wire S482;
wire S483;
wire S484;
wire S485;
wire S486;
wire S487;
wire S488;
wire S489;
wire S490;
wire S491;
wire S492;
wire S493;
wire S494;
wire S495;
wire S496;
wire S497;
wire S498;
wire S499;
wire S500;
wire S501;
wire S502;
wire S503;
wire S504;
wire S505;
wire S506;
wire S507;
wire S508;
wire S509;
wire S510;
wire S511;
wire S512;
wire S513;
wire S514;
wire S515;
wire S516;
wire S517;
wire S518;
wire S519;
wire S520;
wire S521;
wire S522;
wire S523;
wire S524;
wire S525;
wire S526;
wire S527;
wire S528;
wire S529;
wire S530;
wire S531;
wire S532;
wire S533;
wire S534;
wire S535;
wire S536;
wire S537;
wire S538;
wire S539;
wire S540;
wire S541;
wire S542;
wire S543;
wire S544;
wire S545;
wire S546;
wire S547;
wire S548;
wire S549;
wire S550;
wire S551;
wire S552;
wire S553;
wire S554;
wire S555;
wire S556;
wire S557;
wire S558;
wire S559;
wire S560;
wire S561;
wire S562;
wire S563;
wire S564;
wire S565;
wire S566;
wire S567;
wire S568;
wire S569;
wire S570;
wire S571;
wire S572;
wire S573;
wire S574;
wire S575;
wire S576;
wire S577;
wire S578;
wire S579;
wire S580;
wire S581;
wire S582;
wire S583;
wire S584;
wire S585;
wire S586;
wire S587;
wire S588;
wire S589;
wire S590;
wire S591;
wire S592;
wire S593;
wire S594;
wire S595;
wire S596;
wire S597;
wire S598;
wire S599;
wire S600;
wire S601;
wire S602;
wire S603;
wire S604;
wire S605;
wire S606;
wire S607;
wire S608;
wire S609;
wire S610;
wire S611;
wire S612;
wire S613;
wire S614;
wire S615;
wire S616;
wire S617;
wire S618;
wire S619;
wire S620;
wire S621;
wire S622;
wire S623;
wire S624;
wire S625;
wire S626;
wire S627;
wire S628;
wire S629;
wire S630;
wire S631;
wire S632;
wire S633;
wire S634;
wire S635;
wire S636;
wire S637;
wire S638;
wire S639;
wire S640;
wire S641;
wire S642;
wire S643;
wire S644;
wire S645;
wire S646;
wire S647;
wire S648;
wire S649;
wire S650;
wire S651;
wire S652;
wire S653;
wire S654;
wire S655;
wire S656;
wire S657;
wire S658;
wire S659;
wire S660;
wire S661;
wire S662;
wire S663;
wire S664;
wire S665;
wire S666;
wire S667;
wire S668;
wire S669;
wire S670;
wire S671;
wire S672;
wire S673;
wire S674;
wire S675;
wire S676;
wire S677;
wire S678;
wire S679;
wire S680;
wire S681;
wire S682;
wire S683;
wire S684;
wire S685;
wire S686;
wire S687;
wire S688;
wire S689;
wire S690;
wire S691;
wire S692;
wire S693;
wire S694;
wire S695;
wire S696;
wire S697;
wire S698;
wire S699;
wire S700;
wire S701;
wire S702;
wire S703;
wire S704;
wire S705;
wire S706;
wire S707;
wire S708;
wire S709;
wire S710;
wire S711;
wire S712;
wire S713;
wire S714;
wire S715;
wire S716;
wire S717;
wire S718;
wire S719;
wire S720;
wire S721;
wire S722;
wire S723;
wire S724;
wire S725;
wire S726;
wire S727;
wire S728;
wire S729;
wire S730;
wire S731;
wire S732;
wire S733;
wire S734;
wire S735;
wire S736;
wire S737;
wire S738;
wire S739;
wire S740;
wire S741;
wire S742;
wire S743;
wire S744;
wire S745;
wire S746;
wire S747;
wire S748;
wire S749;
wire S750;
wire S751;
wire S752;
wire S753;
wire S754;
wire S755;
wire S756;
wire S757;
wire S758;
wire S759;
wire S760;
wire S761;
wire S762;
wire S763;
wire S764;
wire S765;
wire S766;
wire S767;
wire S768;
wire S769;
wire S770;
wire S771;
wire S772;
wire S773;
wire S774;
wire S775;
wire S776;
wire S777;
wire S778;
wire S779;
wire S780;
wire S781;
wire S782;
wire S783;
wire S784;
wire S785;
wire S786;
wire S787;
wire S788;
wire S789;
wire S790;
wire S791;
wire S792;
wire S793;
wire S794;
wire S795;
wire S796;
wire S797;
wire S798;
wire S799;
wire S800;
wire S801;
wire S802;
wire S803;
wire S804;
wire S805;
wire S806;
wire S807;
wire S808;
wire S809;
wire S810;
wire S811;
wire S812;
wire S813;
wire S814;
wire S815;
wire S816;
wire S817;
wire S818;
wire S819;
wire S820;
wire S821;
wire S822;
wire S823;
wire S824;
wire S825;
wire S826;
wire S827;
wire S828;
wire S829;
wire S830;
wire S831;
wire S832;
wire S833;
wire S834;
wire S835;
wire S836;
wire S837;
wire S838;
wire S839;
wire S840;
wire S841;
wire S842;
wire S843;
wire S844;
wire S845;
wire S846;
wire S847;
wire S848;
wire S849;
wire S850;
wire S851;
wire S852;
wire S853;
wire S854;
wire S855;
wire S856;
wire S857;
wire S858;
wire S859;
wire S860;
wire S861;
wire S862;
wire S863;
wire S864;
wire S865;
wire S866;
wire S867;
wire S868;
wire S869;
wire S870;
wire S871;
wire S872;
wire S873;
wire S874;
wire S875;
wire S876;
wire S877;
wire S878;
wire S879;
wire S880;
wire S881;
wire S882;
wire S883;
wire S884;
wire S885;
wire S886;
wire S887;
wire S888;
wire S889;
wire S890;
wire S891;
wire S892;
wire S893;
wire S894;
wire S895;
wire S896;
wire S897;
wire S898;
wire S899;
wire S900;
wire S901;
wire S902;
wire S903;
wire S904;
wire S905;
wire S906;
wire S907;
wire S908;
wire S909;
wire S910;
wire S911;
wire S912;
wire S913;
wire S914;
wire S915;
wire S916;
wire S917;
wire S918;
wire S919;
wire S920;
wire S921;
wire S922;
wire S923;
wire S924;
wire S925;
wire S926;
wire S927;
wire S928;
wire S929;
wire S930;
wire S931;
wire S932;
wire S933;
wire S934;
wire S935;
wire S936;
wire S937;
wire S938;
wire S939;
wire S940;
wire S941;
wire S942;
wire S943;
wire S944;
wire S945;
wire S946;
wire S947;
wire S948;
wire S949;
wire S950;
wire S951;
wire S952;
wire S953;
wire S954;
wire S955;
wire S956;
wire S957;
wire S958;
wire S959;
wire S960;
wire S961;
wire S962;
wire S963;
wire S964;
wire S965;
wire S966;
wire S967;
wire S968;
wire S969;
wire S970;
wire S971;
wire S972;
wire S973;
wire S974;
wire S975;
wire S976;
wire S977;
wire S978;
wire S979;
wire S980;
wire S981;
wire S982;
wire S983;
wire S984;
wire S985;
wire S986;
wire S987;
wire S988;
wire S989;
wire S990;
wire S991;
wire S992;
wire S993;
wire S994;
wire S995;
wire S996;
wire S997;
wire S998;
wire S999;
wire S1000;
wire S1001;
wire S1002;
wire S1003;
wire S1004;
wire S1005;
wire S1006;
wire S1007;
wire S1008;
wire S1009;
wire S1010;
wire S1011;
wire S1012;
wire S1013;
wire S1014;
wire S1015;
wire S1016;
wire S1017;
wire S1018;
wire S1019;
wire S1020;
wire S1021;
wire S1022;
wire S1023;
wire S1024;
wire S1025;
wire S1026;
wire S1027;
wire S1028;
wire S1029;
wire S1030;
wire S1031;
wire S1032;
wire S1033;
wire S1034;
wire S1035;
wire S1036;
wire S1037;
wire S1038;
wire S1039;
wire S1040;
wire S1041;
wire S1042;
wire S1043;
wire S1044;
wire S1045;
wire S1046;
wire S1047;
wire S1048;
wire S1049;
wire S1050;
wire S1051;
wire S1052;
wire S1053;
wire S1054;
wire S1055;
wire S1056;
wire S1057;
wire S1058;
wire S1059;
wire S1060;
wire S1061;
wire S1062;
wire S1063;
wire S1064;
wire S1065;
wire S1066;
wire S1067;
wire S1068;
wire S1069;
wire S1070;
wire S1071;
wire S1072;
wire S1073;
wire S1074;
wire S1075;
wire S1076;
wire S1077;
wire S1078;
wire S1079;
wire S1080;
wire S1081;
wire S1082;
wire S1083;
wire S1084;
wire S1085;
wire S1086;
wire S1087;
wire S1088;
wire S1089;
wire S1090;
wire S1091;
wire S1092;
wire S1093;
wire S1094;
wire S1095;
wire S1096;
wire S1097;
wire S1098;
wire S1099;
wire S1100;
wire S1101;
wire S1102;
wire S1103;
wire S1104;
wire S1105;
wire S1106;
wire S1107;
wire S1108;
wire S1109;
wire S1110;
wire S1111;
wire S1112;
wire S1113;
wire S1114;
wire S1115;
wire S1116;
wire S1117;
wire S1118;
wire S1119;
wire S1120;
wire S1121;
wire S1122;
wire S1123;
wire S1124;
wire S1125;
wire S1126;
wire S1127;
wire S1128;
wire S1129;
wire S1130;
wire S1131;
wire S1132;
wire S1133;
wire S1134;
wire S1135;
wire S1136;
wire S1137;
wire S1138;
wire S1139;
wire S1140;
wire S1141;
wire S1142;
wire S1143;
wire S1144;
wire S1145;
wire S1146;
wire S1147;
wire S1148;
wire S1149;
wire S1150;
wire S1151;
wire S1152;
wire S1153;
wire S1154;
wire S1155;
wire S1156;
wire S1157;
wire S1158;
wire S1159;
wire S1160;
wire S1161;
wire S1162;
wire S1163;
wire S1164;
wire S1165;
wire S1166;
wire S1167;
wire S1168;
wire S1169;
wire S1170;
wire S1171;
wire S1172;
wire S1173;
wire S1174;
wire S1175;
wire S1176;
wire S1177;
wire S1178;
wire S1179;
wire S1180;
wire S1181;
wire S1182;
wire S1183;
wire S1184;
wire S1185;
wire S1186;
wire S1187;
wire S1188;
wire S1189;
wire S1190;
wire S1191;
wire S1192;
wire S1193;
wire S1194;
wire S1195;
wire S1196;
wire S1197;
wire S1198;
wire S1199;
wire S1200;
wire S1201;
wire S1202;
wire S1203;
wire S1204;
wire S1205;
wire S1206;
wire S1207;
wire S1208;
wire S1209;
wire S1210;
wire S1211;
wire S1212;
wire S1213;
wire S1214;
wire S1215;
wire S1216;
wire S1217;
wire S1218;
wire S1219;
wire S1220;
wire S1221;
wire S1222;
wire S1223;
wire S1224;
wire S1225;
wire S1226;
wire S1227;
wire S1228;
wire S1229;
wire S1230;
wire S1231;
wire S1232;
wire S1233;
wire S1234;
wire S1235;
wire S1236;
wire S1237;
wire S1238;
wire S1239;
wire S1240;
wire S1241;
wire S1242;
wire S1243;
wire S1244;
wire S1245;
wire S1246;
wire S1247;
wire S1248;
wire S1249;
wire S1250;
wire S1251;
wire S1252;
wire S1253;
wire S1254;
wire S1255;
wire S1256;
wire S1257;
wire S1258;
wire S1259;
wire S1260;
wire S1261;
wire S1262;
wire S1263;
wire S1264;
wire S1265;
wire S1266;
wire S1267;
wire S1268;
wire S1269;
wire S1270;
wire S1271;
wire S1272;
wire S1273;
wire S1274;
wire S1275;
wire S1276;
wire S1277;
wire S1278;
wire S1279;
wire S1280;
wire S1281;
wire S1282;
wire S1283;
wire S1284;
wire S1285;
wire S1286;
wire S1287;
wire S1288;
wire S1289;
wire S1290;
wire S1291;
wire S1292;
wire S1293;
wire S1294;
wire S1295;
wire S1296;
wire S1297;
wire S1298;
wire S1299;
wire S1300;
wire S1301;
wire S1302;
wire S1303;
wire S1304;
wire S1305;
wire S1306;
wire S1307;
wire S1308;
wire S1309;
wire S1310;
wire S1311;
wire S1312;
wire S1313;
wire S1314;
wire S1315;
wire S1316;
wire S1317;
wire S1318;
wire S1319;
wire S1320;
wire S1321;
wire S1322;
wire S1323;
wire S1324;
wire S1325;
wire S1326;
wire S1327;
wire S1328;
wire S1329;
wire S1330;
wire S1331;
wire S1332;
wire S1333;
wire S1334;
wire S1335;
wire S1336;
wire S1337;
wire S1338;
wire S1339;
wire S1340;
wire S1341;
wire S1342;
wire S1343;
wire S1344;
wire S1345;
wire S1346;
wire S1347;
wire S1348;
wire S1349;
wire S1350;
wire S1351;
wire S1352;
wire S1353;
wire S1354;
wire S1355;
wire S1356;
wire S1357;
wire S1358;
wire S1359;
wire S1360;
wire S1361;
wire S1362;
wire S1363;
wire S1364;
wire S1365;
wire S1366;
wire S1367;
wire S1368;
wire S1369;
wire S1370;
wire S1371;
wire S1372;
wire S1373;
wire S1374;
wire S1375;
wire S1376;
wire S1377;
wire S1378;
wire S1379;
wire S1380;
wire S1381;
wire S1382;
wire S1383;
wire S1384;
wire S1385;
wire S1386;
wire S1387;
wire S1388;
wire S1389;
wire S1390;
wire S1391;
wire S1392;
wire S1393;
wire S1394;
wire S1395;
wire S1396;
wire S1397;
wire S1398;
wire S1399;
wire S1400;
wire S1401;
wire S1402;
wire S1403;
wire S1404;
wire S1405;
wire S1406;
wire S1407;
wire S1408;
wire S1409;
wire S1410;
wire S1411;
wire S1412;
wire S1413;
wire S1414;
wire S1415;
wire S1416;
wire S1417;
wire S1418;
wire S1419;
wire S1420;
wire S1421;
wire S1422;
wire S1423;
wire S1424;
wire S1425;
wire S1426;
wire S1427;
wire S1428;
wire S1429;
wire S1430;
wire S1431;
wire S1432;
wire S1433;
wire S1434;
wire S1435;
wire S1436;
wire S1437;
wire S1438;
wire S1439;
wire S1440;
wire S1441;
wire S1442;
wire S1443;
wire S1444;
wire S1445;
wire S1446;
wire S1447;
wire S1448;
wire S1449;
wire S1450;
wire S1451;
wire S1452;
wire S1453;
wire S1454;
wire S1455;
wire S1456;
wire S1457;
wire S1458;
wire S1459;
wire S1460;
wire S1461;
wire S1462;
wire S1463;
wire S1464;
wire S1465;
wire S1466;
wire S1467;
wire S1468;
wire S1469;
wire S1470;
wire S1471;
wire S1472;
wire S1473;
wire S1474;
wire S1475;
wire S1476;
wire S1477;
wire S1478;
wire S1479;
wire S1480;
wire S1481;
wire S1482;
wire S1483;
wire S1484;
wire S1485;
wire S1486;
wire S1487;
wire S1488;
wire S1489;
wire S1490;
wire S1491;
wire S1492;
wire S1493;
wire S1494;
wire S1495;
wire S1496;
wire S1497;
wire S1498;
wire S1499;
wire S1500;
wire S1501;
wire S1502;
wire S1503;
wire S1504;
wire S1505;
wire S1506;
wire S1507;
wire S1508;
wire S1509;
wire S1510;
wire S1511;
wire S1512;
wire S1513;
wire S1514;
wire S1515;
wire S1516;
wire S1517;
wire S1518;
wire S1519;
wire S1520;
wire S1521;
wire S1522;
wire S1523;
wire S1524;
wire S1525;
wire S1526;
wire S1527;
wire S1528;
wire S1529;
wire S1530;
wire S1531;
wire S1532;
wire S1533;
wire S1534;
wire S1535;
wire S1536;
wire S1537;
wire S1538;
wire S1539;
wire S1540;
wire S1541;
wire S1542;
wire S1543;
wire S1544;
wire S1545;
wire S1546;
wire S1547;
wire S1548;
wire S1549;
wire S1550;
wire S1551;
wire S1552;
wire S1553;
wire S1554;
wire S1555;
wire S1556;
wire S1557;
wire S1558;
wire S1559;
wire S1560;
wire S1561;
wire S1562;
wire S1563;
wire S1564;
wire S1565;
wire S1566;
wire S1567;
wire S1568;
wire S1569;
wire S1570;
wire S1571;
wire S1572;
wire S1573;
wire S1574;
wire S1575;
wire S1576;
wire S1577;
wire S1578;
wire S1579;
wire S1580;
wire S1581;
wire S1582;
wire S1583;
wire S1584;
wire S1585;
wire S1586;
wire S1587;
wire S1588;
wire S1589;
wire S1590;
wire S1591;
wire S1592;
wire S1593;
wire S1594;
wire S1595;
wire S1596;
wire S1597;
wire S1598;
wire S1599;
wire S1600;
wire S1601;
wire S1602;
wire S1603;
wire S1604;
wire S1605;
wire S1606;
wire S1607;
wire S1608;
wire S1609;
wire S1610;
wire S1611;
wire S1612;
wire S1613;
wire S1614;
wire S1615;
wire S1616;
wire S1617;
wire S1618;
wire S1619;
wire S1620;
wire S1621;
wire S1622;
wire S1623;
wire S1624;
wire S1625;
wire S1626;
wire S1627;
wire S1628;
wire S1629;
wire S1630;
wire S1631;
wire S1632;
wire S1633;
wire S1634;
wire S1635;
wire S1636;
wire S1637;
wire S1638;
wire S1639;
wire S1640;
wire S1641;
wire S1642;
wire S1643;
wire S1644;
wire S1645;
wire S1646;
wire S1647;
wire S1648;
wire S1649;
wire S1650;
wire S1651;
wire S1652;
wire S1653;
wire S1654;
wire S1655;
wire S1656;
wire S1657;
wire S1658;
wire S1659;
wire S1660;
wire S1661;
wire S1662;
wire S1663;
wire S1664;
wire S1665;
wire S1666;
wire S1667;
wire S1668;
wire S1669;
wire S1670;
wire S1671;
wire S1672;
wire S1673;
wire S1674;
wire S1675;
wire S1676;
wire S1677;
wire S1678;
wire S1679;
wire S1680;
wire S1681;
wire S1682;
wire S1683;
wire S1684;
wire S1685;
wire S1686;
wire S1687;
wire S1688;
wire S1689;
wire S1690;
wire S1691;
wire S1692;
wire S1693;
wire S1694;
wire S1695;
wire S1696;
wire S1697;
wire S1698;
wire S1699;
wire S1700;
wire S1701;
wire S1702;
wire S1703;
wire S1704;
wire S1705;
wire S1706;
wire S1707;
wire S1708;
wire S1709;
wire S1710;
wire S1711;
wire S1712;
wire S1713;
wire S1714;
wire S1715;
wire S1716;
wire S1717;
wire S1718;
wire S1719;
wire S1720;
wire S1721;
wire S1722;
wire S1723;
wire S1724;
wire S1725;
wire S1726;
wire S1727;
wire S1728;
wire S1729;
wire S1730;
wire S1731;
wire S1732;
wire S1733;
wire S1734;
wire S1735;
wire S1736;
wire S1737;
wire S1738;
wire S1739;
wire S1740;
wire S1741;
wire S1742;
wire S1743;
wire S1744;
wire S1745;
wire S1746;
wire S1747;
wire S1748;
wire S1749;
wire S1750;
wire S1751;
wire S1752;
wire S1753;
wire S1754;
wire S1755;
wire S1756;
wire S1757;
wire S1758;
wire S1759;
wire S1760;
wire S1761;
wire S1762;
wire S1763;
wire S1764;
wire S1765;
wire S1766;
wire S1767;
wire S1768;
wire S1769;
wire S1770;
wire S1771;
wire S1772;
wire S1773;
wire S1774;
wire S1775;
wire S1776;
wire S1777;
wire S1778;
wire S1779;
wire S1780;
wire S1781;
wire S1782;
wire S1783;
wire S1784;
wire S1785;
wire S1786;
wire S1787;
wire S1788;
wire S1789;
wire S1790;
wire S1791;
wire S1792;
wire S1793;
wire S1794;
wire S1795;
wire S1796;
wire S1797;
wire S1798;
wire S1799;
wire S1800;
wire S1801;
wire S1802;
wire S1803;
wire S1804;
wire S1805;
wire S1806;
wire S1807;
wire S1808;
wire S1809;
wire S1810;
wire S1811;
wire S1812;
wire S1813;
wire S1814;
wire S1815;
wire S1816;
wire S1817;
wire S1818;
wire S1819;
wire S1820;
wire S1821;
wire S1822;
wire S1823;
wire S1824;
wire S1825;
wire S1826;
wire S1827;
wire S1828;
wire S1829;
wire S1830;
wire S1831;
wire S1832;
wire S1833;
wire S1834;
wire S1835;
wire S1836;
wire S1837;
wire S1838;
wire S1839;
wire S1840;
wire S1841;
wire S1842;
wire S1843;
wire S1844;
wire S1845;
wire S1846;
wire S1847;
wire S1848;
wire S1849;
wire S1850;
wire S1851;
wire S1852;
wire S1853;
wire S1854;
wire S1855;
wire S1856;
wire S1857;
wire S1858;
wire S1859;
wire S1860;
wire S1861;
wire S1862;
wire S1863;
wire S1864;
wire S1865;
wire S1866;
wire S1867;
wire S1868;
wire S1869;
wire S1870;
wire S1871;
wire S1872;
wire S1873;
wire S1874;
wire S1875;
wire S1876;
wire S1877;
wire S1878;
wire S1879;
wire S1880;
wire S1881;
wire S1882;
wire S1883;
wire S1884;
wire S1885;
wire S1886;
wire S1887;
wire S1888;
wire S1889;
wire S1890;
wire S1891;
wire S1892;
wire S1893;
wire S1894;
wire S1895;
wire S1896;
wire S1897;
wire S1898;
wire S1899;
wire S1900;
wire S1901;
wire S1902;
wire S1903;
wire S1904;
wire S1905;
wire S1906;
wire S1907;
wire S1908;
wire S1909;
wire S1910;
wire S1911;
wire S1912;
wire S1913;
wire S1914;
wire S1915;
wire S1916;
wire S1917;
wire S1918;
wire S1919;
wire S1920;
wire S1921;
wire S1922;
wire S1923;
wire S1924;
wire S1925;
wire S1926;
wire S1927;
wire S1928;
wire S1929;
wire S1930;
wire S1931;
wire S1932;
wire S1933;
wire S1934;
wire S1935;
wire S1936;
wire S1937;
wire S1938;
wire S1939;
wire S1940;
wire S1941;
wire S1942;
wire S1943;
wire S1944;
wire S1945;
wire S1946;
wire S1947;
wire S1948;
wire S1949;
wire S1950;
wire S1951;
wire S1952;
wire S1953;
wire S1954;
wire S1955;
wire S1956;
wire S1957;
wire S1958;
wire S1959;
wire S1960;
wire S1961;
wire S1962;
wire S1963;
wire S1964;
wire S1965;
wire S1966;
wire S1967;
wire S1968;
wire S1969;
wire S1970;
wire S1971;
wire S1972;
wire S1973;
wire S1974;
wire S1975;
wire S1976;
wire S1977;
wire S1978;
wire S1979;
wire S1980;
wire S1981;
wire S1982;
wire S1983;
wire S1984;
wire S1985;
wire S1986;
wire S1987;
wire S1988;
wire S1989;
wire S1990;
wire S1991;
wire S1992;
wire S1993;
wire S1994;
wire S1995;
wire S1996;
wire S1997;
wire S1998;
wire S1999;
wire S2000;
wire S2001;
wire S2002;
wire S2003;
wire S2004;
wire S2005;
wire S2006;
wire S2007;
wire S2008;
wire S2009;
wire S2010;
wire S2011;
wire S2012;
wire S2013;
wire S2014;
wire S2015;
wire S2016;
wire S2017;
wire S2018;
wire S2019;
wire S2020;
wire S2021;
wire S2022;
wire S2023;
wire S2024;
wire S2025;
wire S2026;
wire S2027;
wire S2028;
wire S2029;
wire S2030;
wire S2031;
wire S2032;
wire S2033;
wire S2034;
wire S2035;
wire S2036;
wire S2037;
wire S2038;
wire S2039;
wire S2040;
wire S2041;
wire S2042;
wire S2043;
wire S2044;
wire S2045;
wire S2046;
wire S2047;
wire S2048;
wire S2049;
wire S2050;
wire S2051;
wire S2052;
wire S2053;
wire S2054;
wire S2055;
wire S2056;
wire S2057;
wire S2058;
wire S2059;
wire S2060;
wire S2061;
wire S2062;
wire S2063;
wire S2064;
wire S2065;
wire S2066;
wire S2067;
wire S2068;
wire S2069;
wire S2070;
wire S2071;
wire S2072;
wire S2073;
wire S2074;
wire S2075;
wire S2076;
wire S2077;
wire S2078;
wire S2079;
wire S2080;
wire S2081;
wire S2082;
wire S2083;
wire S2084;
wire S2085;
wire S2086;
wire S2087;
wire S2088;
wire S2089;
wire S2090;
wire S2091;
wire S2092;
wire S2093;
wire S2094;
wire S2095;
wire S2096;
wire S2097;
wire S2098;
wire S2099;
wire S2100;
wire S2101;
wire S2102;
wire S2103;
wire S2104;
wire S2105;
wire S2106;
wire S2107;
wire S2108;
wire S2109;
wire S2110;
wire S2111;
wire S2112;
wire S2113;
wire S2114;
wire S2115;
wire S2116;
wire S2117;
wire S2118;
wire S2119;
wire S2120;
wire S2121;
wire S2122;
wire S2123;
wire S2124;
wire S2125;
wire S2126;
wire S2127;
wire S2128;
wire S2129;
wire S2130;
wire S2131;
wire S2132;
wire S2133;
wire S2134;
wire S2135;
wire S2136;
wire S2137;
wire S2138;
wire S2139;
wire S2140;
wire S2141;
wire S2142;
wire S2143;
wire S2144;
wire S2145;
wire S2146;
wire S2147;
wire S2148;
wire S2149;
wire S2150;
wire S2151;
wire S2152;
wire S2153;
wire S2154;
wire S2155;
wire S2156;
wire S2157;
wire S2158;
wire S2159;
wire S2160;
wire S2161;
wire S2162;
wire S2163;
wire S2164;
wire S2165;
wire S2166;
wire S2167;
wire S2168;
wire S2169;
wire S2170;
wire S2171;
wire S2172;
wire S2173;
wire S2174;
wire S2175;
wire S2176;
wire S2177;
wire S2178;
wire S2179;
wire S2180;
wire S2181;
wire S2182;
wire S2183;
wire S2184;
wire S2185;
wire S2186;
wire S2187;
wire S2188;
wire S2189;
wire S2190;
wire S2191;
wire S2192;
wire S2193;
wire S2194;
wire S2195;
wire S2196;
wire S2197;
wire S2198;
wire S2199;
wire S2200;
wire S2201;
wire S2202;
wire S2203;
wire S2204;
wire S2205;
wire S2206;
wire S2207;
wire S2208;
wire S2209;
wire S2210;
wire S2211;
wire S2212;
wire S2213;
wire S2214;
wire S2215;
wire S2216;
wire S2217;
wire S2218;
wire S2219;
wire S2220;
wire S2221;
wire S2222;
wire S2223;
wire S2224;
wire S2225;
wire S2226;
wire S2227;
wire S2228;
wire S2229;
wire S2230;
wire S2231;
wire S2232;
wire S2233;
wire S2234;
wire S2235;
wire S2236;
wire S2237;
wire S2238;
wire S2239;
wire S2240;
wire S2241;
wire S2242;
wire S2243;
wire S2244;
wire S2245;
wire S2246;
wire S2247;
wire S2248;
wire S2249;
wire S2250;
wire S2251;
wire S2252;
wire S2253;
wire S2254;
wire S2255;
wire S2256;
wire S2257;
wire S2258;
wire S2259;
wire S2260;
wire S2261;
wire S2262;
wire S2263;
wire S2264;
wire S2265;
wire S2266;
wire S2267;
wire S2268;
wire S2269;
wire S2270;
wire S2271;
wire S2272;
wire S2273;
wire S2274;
wire S2275;
wire S2276;
wire S2277;
wire S2278;
wire S2279;
wire S2280;
wire S2281;
wire S2282;
wire S2283;
wire S2284;
wire S2285;
wire S2286;
wire S2287;
wire S2288;
wire S2289;
wire S2290;
wire S2291;
wire S2292;
wire S2293;
wire S2294;
wire S2295;
wire S2296;
wire S2297;
wire S2298;
wire S2299;
wire S2300;
wire S2301;
wire S2302;
wire S2303;
wire S2304;
wire S2305;
wire S2306;
wire S2307;
wire S2308;
wire S2309;
wire S2310;
wire S2311;
wire S2312;
wire S2313;
wire S2314;
wire S2315;
wire S2316;
wire S2317;
wire S2318;
wire S2319;
wire S2320;
wire S2321;
wire S2322;
wire S2323;
wire S2324;
wire S2325;
wire S2326;
wire S2327;
wire S2328;
wire S2329;
wire S2330;
wire S2331;
wire S2332;
wire S2333;
wire S2334;
wire S2335;
wire S2336;
wire S2337;
wire S2338;
wire S2339;
wire S2340;
wire S2341;
wire S2342;
wire S2343;
wire S2344;
wire S2345;
wire S2346;
wire S2347;
wire S2348;
wire S2349;
wire S2350;
wire S2351;
wire S2352;
wire S2353;
wire S2354;
wire S2355;
wire S2356;
wire S2357;
wire S2358;
wire S2359;
wire S2360;
wire S2361;
wire S2362;
wire S2363;
wire S2364;
wire S2365;
wire S2366;
wire S2367;
wire S2368;
wire S2369;
wire S2370;
wire S2371;
wire S2372;
wire S2373;
wire S2374;
wire S2375;
wire S2376;
wire S2377;
wire S2378;
wire S2379;
wire S2380;
wire S2381;
wire S2382;
wire S2383;
wire S2384;
wire S2385;
wire S2386;
wire S2387;
wire S2388;
wire S2389;
wire S2390;
wire S2391;
wire S2392;
wire S2393;
wire S2394;
wire S2395;
wire S2396;
wire S2397;
wire S2398;
wire S2399;
wire S2400;
wire S2401;
wire S2402;
wire S2403;
wire S2404;
wire S2405;
wire S2406;
wire S2407;
wire S2408;
wire S2409;
wire S2410;
wire S2411;
wire S2412;
wire S2413;
wire S2414;
wire S2415;
wire S2416;
wire S2417;
wire S2418;
wire S2419;
wire S2420;
wire S2421;
wire S2422;
wire S2423;
wire S2424;
wire S2425;
wire S2426;
wire S2427;
wire S2428;
wire S2429;
wire S2430;
wire S2431;
wire S2432;
wire S2433;
wire S2434;
wire S2435;
wire S2436;
wire S2437;
wire S2438;
wire S2439;
wire S2440;
wire S2441;
wire S2442;
wire S2443;
wire S2444;
wire S2445;
wire S2446;
wire S2447;
wire S2448;
wire S2449;
wire S2450;
wire S2451;
wire S2452;
wire S2453;
wire S2454;
wire S2455;
wire S2456;
wire S2457;
wire S2458;
wire S2459;
wire S2460;
wire S2461;
wire S2462;
wire S2463;
wire S2464;
wire S2465;
wire S2466;
wire S2467;
wire S2468;
wire S2469;
wire S2470;
wire S2471;
wire S2472;
wire S2473;
wire S2474;
wire S2475;
wire S2476;
wire S2477;
wire S2478;
wire S2479;
wire S2480;
wire S2481;
wire S2482;
wire S2483;
wire S2484;
wire S2485;
wire S2486;
wire S2487;
wire S2488;
wire S2489;
wire S2490;
wire S2491;
wire S2492;
wire S2493;
wire S2494;
wire S2495;
wire S2496;
wire S2497;
wire S2498;
wire S2499;
wire S2500;
wire S2501;
wire S2502;
wire S2503;
wire S2504;
wire S2505;
wire S2506;
wire S2507;
wire S2508;
wire S2509;
wire S2510;
wire S2511;
wire S2512;
wire S2513;
wire S2514;
wire S2515;
wire S2516;
wire S2517;
wire S2518;
wire S2519;
wire S2520;
wire S2521;
wire S2522;
wire S2523;
wire S2524;
wire S2525;
wire S2526;
wire S2527;
wire S2528;
wire S2529;
wire S2530;
wire S2531;
wire S2532;
wire S2533;
wire S2534;
wire S2535;
wire S2536;
wire S2537;
wire S2538;
wire S2539;
wire S2540;
wire S2541;
wire S2542;
wire S2543;
wire S2544;
wire S2545;
wire S2546;
wire S2547;
wire S2548;
wire S2549;
wire S2550;
wire S2551;
wire S2552;
wire S2553;
wire S2554;
wire S2555;
wire S2556;
wire S2557;
wire S2558;
wire S2559;
wire S2560;
wire S2561;
wire S2562;
wire S2563;
wire S2564;
wire S2565;
wire S2566;
wire S2567;
wire S2568;
wire S2569;
wire S2570;
wire S2571;
wire S2572;
wire S2573;
wire S2574;
wire S2575;
wire S2576;
wire S2577;
wire S2578;
wire S2579;
wire S2580;
wire S2581;
wire S2582;
wire S2583;
wire S2584;
wire S2585;
wire S2586;
wire S2587;
wire S2588;
wire S2589;
wire S2590;
wire S2591;
wire S2592;
wire S2593;
wire S2594;
wire S2595;
wire S2596;
wire S2597;
wire S2598;
wire S2599;
wire S2600;
wire S2601;
wire S2602;
wire S2603;
wire S2604;
wire S2605;
wire S2606;
wire S2607;
wire S2608;
wire S2609;
wire S2610;
wire S2611;
wire S2612;
wire S2613;
wire S2614;
wire S2615;
wire S2616;
wire CU_inst_0;
wire CU_inst_10;
wire CU_inst_11;
wire CU_inst_12;
wire CU_inst_13;
wire CU_inst_14;
wire CU_inst_15;
wire CU_inst_1;
wire CU_inst_2;
wire CU_inst_3;
wire CU_inst_4;
wire CU_inst_5;
wire CU_inst_6;
wire CU_inst_7;
wire CU_inst_8;
wire CU_inst_9;
wire CU_nstate_0;
wire CU_nstate_1;
wire CU_pstate_0;
wire CU_pstate_1;
wire DP_AC_q_0;
wire DP_AC_q_10;
wire DP_AC_q_11;
wire DP_AC_q_12;
wire DP_AC_q_13;
wire DP_AC_q_14;
wire DP_AC_q_15;
wire DP_AC_q_1;
wire DP_AC_q_2;
wire DP_AC_q_3;
wire DP_AC_q_4;
wire DP_AC_q_5;
wire DP_AC_q_6;
wire DP_AC_q_7;
wire DP_AC_q_8;
wire DP_AC_q_9;
wire DP_IMM1_in1_0;
wire DP_IMM1_in1_1;
wire DP_IMM1_in1_2;
wire DP_IMM1_in1_3;
wire DP_IN_q_0;
wire DP_IN_q_10;
wire DP_IN_q_11;
wire DP_IN_q_12;
wire DP_IN_q_13;
wire DP_IN_q_14;
wire DP_IN_q_15;
wire DP_IN_q_1;
wire DP_IN_q_2;
wire DP_IN_q_3;
wire DP_IN_q_4;
wire DP_IN_q_5;
wire DP_IN_q_6;
wire DP_IN_q_7;
wire DP_IN_q_8;
wire DP_IN_q_9;
wire DP_INC_1_in_0;
wire DP_INC_1_in_10;
wire DP_INC_1_in_11;
wire DP_INC_1_in_12;
wire DP_INC_1_in_13;
wire DP_INC_1_in_14;
wire DP_INC_1_in_15;
wire DP_INC_1_in_1;
wire DP_INC_1_in_2;
wire DP_INC_1_in_3;
wire DP_INC_1_in_4;
wire DP_INC_1_in_5;
wire DP_INC_1_in_6;
wire DP_INC_1_in_7;
wire DP_INC_1_in_8;
wire DP_INC_1_in_9;
wire DP_SR_C_q;
wire DP_SR_N_q;
wire DP_SR_V_q;
wire DP_SR_Z_q;
input clk;
input rst;
output writeMEM;
output readMEM;
input [15:0] dataBus_in;output [15:0] dataBus_out;output [15:0] addrBus;
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1_ (
  .in1({ S1864, S1861 }),
  .out1({ S1865 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_2_ (
  .in1({ S1865, S1775 }),
  .out1({ S1866 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_3_ (
  .in1({ S1866, S1849 }),
  .out1({ S71 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_1_ (
  .in1({ CU_pstate_0 }),
  .out1({ S1063 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_2_ (
  .in1({ CU_pstate_1 }),
  .out1({ S1073 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_3_ (
  .in1({ CU_inst_12 }),
  .out1({ S1083 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_4_ (
  .in1({ CU_inst_13 }),
  .out1({ S1093 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_5_ (
  .in1({ CU_inst_15 }),
  .out1({ S1103 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_6_ (
  .in1({ CU_inst_14 }),
  .out1({ S1113 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_7_ (
  .in1({ CU_inst_9 }),
  .out1({ S1123 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_8_ (
  .in1({ CU_inst_8 }),
  .out1({ S1132 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_9_ (
  .in1({ CU_inst_11 }),
  .out1({ S1143 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_10_ (
  .in1({ CU_inst_10 }),
  .out1({ S1153 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_11_ (
  .in1({ CU_inst_5 }),
  .out1({ S1160 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_12_ (
  .in1({ CU_inst_7 }),
  .out1({ S1168 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_13_ (
  .in1({ CU_inst_0 }),
  .out1({ S1176 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_14_ (
  .in1({ S2538[0] }),
  .out1({ S1183 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_15_ (
  .in1({ DP_AC_q_0 }),
  .out1({ S1191 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_16_ (
  .in1({ DP_AC_q_1 }),
  .out1({ S1202 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_17_ (
  .in1({ DP_AC_q_2 }),
  .out1({ S1213 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_18_ (
  .in1({ DP_AC_q_3 }),
  .out1({ S1224 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_19_ (
  .in1({ DP_AC_q_4 }),
  .out1({ S1235 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_20_ (
  .in1({ DP_AC_q_5 }),
  .out1({ S1246 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_21_ (
  .in1({ DP_AC_q_6 }),
  .out1({ S1257 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_22_ (
  .in1({ DP_AC_q_7 }),
  .out1({ S1268 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_23_ (
  .in1({ S2538[3] }),
  .out1({ S1279 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_24_ (
  .in1({ CU_inst_3 }),
  .out1({ S1290 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_25_ (
  .in1({ DP_AC_q_9 }),
  .out1({ S1301 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_26_ (
  .in1({ DP_AC_q_10 }),
  .out1({ S1312 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_27_ (
  .in1({ DP_AC_q_11 }),
  .out1({ S1323 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_28_ (
  .in1({ DP_AC_q_13 }),
  .out1({ S1334 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_29_ (
  .in1({ DP_AC_q_14 }),
  .out1({ S1345 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_30_ (
  .in1({ DP_AC_q_15 }),
  .out1({ S1356 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_31_ (
  .in1({ CU_inst_4 }),
  .out1({ S1366 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_32_ (
  .in1({ S2538[4] }),
  .out1({ S1377 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_33_ (
  .in1({ S2538[5] }),
  .out1({ S1388 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_34_ (
  .in1({ S2538[6] }),
  .out1({ S1399 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_35_ (
  .in1({ S2538[7] }),
  .out1({ S1410 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_36_ (
  .in1({ S2538[8] }),
  .out1({ S1421 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_37_ (
  .in1({ S2538[10] }),
  .out1({ S1432 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_38_ (
  .in1({ S2538[11] }),
  .out1({ S1443 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_39_ (
  .in1({ DP_IMM1_in1_0 }),
  .out1({ S1453 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_40_ (
  .in1({ S2538[12] }),
  .out1({ S1464 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_41_ (
  .in1({ DP_IMM1_in1_1 }),
  .out1({ S1475 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_42_ (
  .in1({ S2538[13] }),
  .out1({ S1486 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_43_ (
  .in1({ DP_IMM1_in1_2 }),
  .out1({ S1497 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_44_ (
  .in1({ S2538[14] }),
  .out1({ S1508 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_45_ (
  .in1({ DP_IMM1_in1_3 }),
  .out1({ S1519 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_46_ (
  .in1({ S2538[15] }),
  .out1({ S1529 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_47_ (
  .in1({ DP_INC_1_in_12 }),
  .out1({ S1540 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_48_ (
  .in1({ DP_INC_1_in_13 }),
  .out1({ S1551 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_49_ (
  .in1({ DP_INC_1_in_14 }),
  .out1({ S1562 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_50_ (
  .in1({ DP_INC_1_in_15 }),
  .out1({ S1572 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_51_ (
  .in1({ DP_INC_1_in_0 }),
  .out1({ S1583 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_52_ (
  .in1({ DP_INC_1_in_1 }),
  .out1({ S1594 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_53_ (
  .in1({ DP_INC_1_in_2 }),
  .out1({ S1604 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_54_ (
  .in1({ DP_INC_1_in_3 }),
  .out1({ S1615 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_55_ (
  .in1({ DP_INC_1_in_4 }),
  .out1({ S1626 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_56_ (
  .in1({ DP_INC_1_in_5 }),
  .out1({ S1636 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_57_ (
  .in1({ DP_INC_1_in_6 }),
  .out1({ S1647 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_58_ (
  .in1({ DP_INC_1_in_7 }),
  .out1({ S1657 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_59_ (
  .in1({ DP_INC_1_in_8 }),
  .out1({ S1668 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_60_ (
  .in1({ DP_INC_1_in_9 }),
  .out1({ S1679 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_61_ (
  .in1({ DP_INC_1_in_10 }),
  .out1({ S1689 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_62_ (
  .in1({ DP_INC_1_in_11 }),
  .out1({ S1700 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_63_ (
  .in1({ DP_SR_C_q }),
  .out1({ S1710 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_64_ (
  .in1({ DP_SR_N_q }),
  .out1({ S1721 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_4_ (
  .in1({ S1073, S1063 }),
  .out1({ S1731 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_65_ (
  .in1({ S1731 }),
  .out1({ CU_nstate_0 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1_ (
  .in1({ CU_inst_14, CU_inst_15 }),
  .out1({ S1751 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_66_ (
  .in1({ S1751 }),
  .out1({ S1762 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_2_ (
  .in1({ S1093, CU_inst_12 }),
  .out1({ S1772 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_5_ (
  .in1({ CU_inst_13, S1083 }),
  .out1({ S1783 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_3_ (
  .in1({ S1783, S1762 }),
  .out1({ S1794 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_6_ (
  .in1({ S1772, S1751 }),
  .out1({ S1804 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_4_ (
  .in1({ S1073, CU_pstate_0 }),
  .out1({ S1814 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_7_ (
  .in1({ CU_pstate_1, S1063 }),
  .out1({ S1825 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_5_ (
  .in1({ S1825, S1804 }),
  .out1({ S1835 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_8_ (
  .in1({ S1814, S1794 }),
  .out1({ S1846 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_6_ (
  .in1({ S1113, CU_inst_15 }),
  .out1({ S1856 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_9_ (
  .in1({ CU_inst_14, S1103 }),
  .out1({ S1867 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_7_ (
  .in1({ S1867, CU_inst_13 }),
  .out1({ S1868 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_10_ (
  .in1({ S1856, S1093 }),
  .out1({ S1869 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_8_ (
  .in1({ S1869, S1825 }),
  .out1({ S1870 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_11_ (
  .in1({ S1868, S1814 }),
  .out1({ S1871 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_9_ (
  .in1({ S1871, CU_inst_12 }),
  .out1({ S1872 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_12_ (
  .in1({ S1870, S1083 }),
  .out1({ S1873 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_10_ (
  .in1({ S1872, S1835 }),
  .out1({ S1874 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_13_ (
  .in1({ S1873, S1846 }),
  .out1({ S1875 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_11_ (
  .in1({ S1113, S1103 }),
  .out1({ S1876 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_14_ (
  .in1({ CU_inst_14, CU_inst_15 }),
  .out1({ S1877 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_12_ (
  .in1({ CU_inst_14, S1103 }),
  .out1({ S1878 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_15_ (
  .in1({ S1113, CU_inst_15 }),
  .out1({ S1879 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_13_ (
  .in1({ S1103, CU_inst_12 }),
  .out1({ S1880 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_16_ (
  .in1({ S1878, CU_inst_12 }),
  .out1({ S1881 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_14_ (
  .in1({ CU_pstate_1, S1063 }),
  .out1({ S1882 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_17_ (
  .in1({ S1073, CU_pstate_0 }),
  .out1({ S1883 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_15_ (
  .in1({ S1093, S1083 }),
  .out1({ S1884 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_18_ (
  .in1({ CU_inst_13, CU_inst_12 }),
  .out1({ S1885 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_19_ (
  .in1({ S1884, S1103 }),
  .out1({ S1886 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_20_ (
  .in1({ S1886, S1881 }),
  .out1({ S1887 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_16_ (
  .in1({ S1887, S1883 }),
  .out1({ S1888 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_17_ (
  .in1({ S1762, CU_inst_13 }),
  .out1({ S1889 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_21_ (
  .in1({ S1751, S1093 }),
  .out1({ S1890 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_18_ (
  .in1({ CU_inst_13, S1083 }),
  .out1({ S1891 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_19_ (
  .in1({ S1890, S1083 }),
  .out1({ S1892 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_20_ (
  .in1({ S1879, S1783 }),
  .out1({ S1893 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_22_ (
  .in1({ S1878, S1772 }),
  .out1({ S1894 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_23_ (
  .in1({ CU_inst_14, CU_inst_13 }),
  .out1({ S1895 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_67_ (
  .in1({ S1895 }),
  .out1({ S1896 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_21_ (
  .in1({ S1856, S1772 }),
  .out1({ S1897 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_24_ (
  .in1({ S1867, S1783 }),
  .out1({ S1898 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_22_ (
  .in1({ S1895, CU_inst_15 }),
  .out1({ S1899 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_25_ (
  .in1({ S1856, CU_inst_13 }),
  .out1({ S1900 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_23_ (
  .in1({ S1879, CU_inst_13 }),
  .out1({ S1901 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_26_ (
  .in1({ S1878, S1093 }),
  .out1({ S1902 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_24_ (
  .in1({ S1901, S1899 }),
  .out1({ S1903 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_27_ (
  .in1({ S1902, S1900 }),
  .out1({ S1904 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_25_ (
  .in1({ S1903, CU_inst_12 }),
  .out1({ S1905 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_28_ (
  .in1({ S1904, S1083 }),
  .out1({ S1906 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_29_ (
  .in1({ S1906, S1890 }),
  .out1({ S1907 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_30_ (
  .in1({ S1898, S1895 }),
  .out1({ S1908 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_26_ (
  .in1({ S1897, S1896 }),
  .out1({ S1909 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_27_ (
  .in1({ S1909, S1892 }),
  .out1({ S1910 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_31_ (
  .in1({ S1910, S1888 }),
  .out1({ S1911 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_28_ (
  .in1({ S1911, S1876 }),
  .out1({ S1912 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_68_ (
  .in1({ S1912 }),
  .out1({ S1913 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_29_ (
  .in1({ S1871, S1083 }),
  .out1({ S1914 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_32_ (
  .in1({ S1870, CU_inst_12 }),
  .out1({ S1915 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_30_ (
  .in1({ S1885, S1877 }),
  .out1({ S1916 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_33_ (
  .in1({ S1884, S1876 }),
  .out1({ S1917 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_31_ (
  .in1({ S1890, CU_inst_12 }),
  .out1({ S1918 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_34_ (
  .in1({ S1889, S1083 }),
  .out1({ S1919 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_32_ (
  .in1({ S1918, S1883 }),
  .out1({ S1920 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_35_ (
  .in1({ S1919, S1882 }),
  .out1({ S1921 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_33_ (
  .in1({ S1921, S1905 }),
  .out1({ S1922 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_36_ (
  .in1({ S1920, S1906 }),
  .out1({ S1923 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_34_ (
  .in1({ S1923, S1916 }),
  .out1({ S1924 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_37_ (
  .in1({ S1922, S1917 }),
  .out1({ S1925 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_35_ (
  .in1({ S1924, S1914 }),
  .out1({ S1926 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_38_ (
  .in1({ S1925, S1915 }),
  .out1({ S1927 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_36_ (
  .in1({ S1927, S1912 }),
  .out1({ S1928 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_39_ (
  .in1({ S1926, S1913 }),
  .out1({ S1929 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_37_ (
  .in1({ S1917, S1883 }),
  .out1({ S1930 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_40_ (
  .in1({ S1916, S1882 }),
  .out1({ S1931 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_38_ (
  .in1({ CU_inst_8, CU_inst_9 }),
  .out1({ S1932 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_39_ (
  .in1({ S1153, CU_inst_11 }),
  .out1({ S1933 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_41_ (
  .in1({ S1933, S1932 }),
  .out1({ S1934 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_69_ (
  .in1({ S1934 }),
  .out1({ S1935 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_40_ (
  .in1({ CU_inst_10, CU_inst_11 }),
  .out1({ S1936 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_70_ (
  .in1({ S1936 }),
  .out1({ S1937 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_42_ (
  .in1({ S1936, CU_inst_9 }),
  .out1({ S1938 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_71_ (
  .in1({ S1938 }),
  .out1({ S1939 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_41_ (
  .in1({ S1939, S1935 }),
  .out1({ S1940 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_43_ (
  .in1({ S1938, S1934 }),
  .out1({ S1941 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_42_ (
  .in1({ S1940, S1931 }),
  .out1({ S1942 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_44_ (
  .in1({ S1941, S1930 }),
  .out1({ S1943 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_43_ (
  .in1({ S1937, S1931 }),
  .out1({ S1944 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_45_ (
  .in1({ S1944, S1932 }),
  .out1({ S1945 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_72_ (
  .in1({ S1945 }),
  .out1({ S1946 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_44_ (
  .in1({ S1946, S1942 }),
  .out1({ S1947 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_46_ (
  .in1({ S1945, S1943 }),
  .out1({ S1948 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_45_ (
  .in1({ S1948, S1929 }),
  .out1({ S1949 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_47_ (
  .in1({ S1947, S1928 }),
  .out1({ S1950 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_46_ (
  .in1({ S1949, S1176 }),
  .out1({ S1951 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_48_ (
  .in1({ S1950, CU_inst_0 }),
  .out1({ S1952 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_47_ (
  .in1({ S1877, CU_inst_13 }),
  .out1({ S1953 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_49_ (
  .in1({ S1876, S1093 }),
  .out1({ S1954 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_48_ (
  .in1({ S1954, CU_inst_12 }),
  .out1({ S1955 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_50_ (
  .in1({ S1953, S1083 }),
  .out1({ S1956 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_49_ (
  .in1({ S1955, S1926 }),
  .out1({ S1957 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_51_ (
  .in1({ S1956, S1927 }),
  .out1({ S1958 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_50_ (
  .in1({ S1958, S1952 }),
  .out1({ S1959 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_52_ (
  .in1({ S1958, DP_INC_1_in_0 }),
  .out1({ S1960 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_51_ (
  .in1({ S1874, DP_IN_q_0 }),
  .out1({ S1961 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_53_ (
  .in1({ S1960, S1874 }),
  .out1({ S1962 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_52_ (
  .in1({ S1962, S1959 }),
  .out1({ S1963 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_53_ (
  .in1({ S1963, S1961 }),
  .out1({ S2536[0] })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_54_ (
  .in1({ S1950, CU_inst_1 }),
  .out1({ S1964 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_73_ (
  .in1({ S1964 }),
  .out1({ S1965 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_54_ (
  .in1({ S1964, S1958 }),
  .out1({ S1966 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_55_ (
  .in1({ S1958, DP_INC_1_in_1 }),
  .out1({ S1967 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_55_ (
  .in1({ S1874, DP_IN_q_1 }),
  .out1({ S1968 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_56_ (
  .in1({ S1967, S1874 }),
  .out1({ S1969 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_56_ (
  .in1({ S1969, S1966 }),
  .out1({ S1970 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_57_ (
  .in1({ S1970, S1968 }),
  .out1({ S2536[1] })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_57_ (
  .in1({ S1950, CU_inst_2 }),
  .out1({ S1971 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_74_ (
  .in1({ S1971 }),
  .out1({ S1972 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_58_ (
  .in1({ S1971, S1958 }),
  .out1({ S1973 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_58_ (
  .in1({ S1958, DP_INC_1_in_2 }),
  .out1({ S1974 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_59_ (
  .in1({ S1874, DP_IN_q_2 }),
  .out1({ S1975 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_59_ (
  .in1({ S1974, S1874 }),
  .out1({ S1976 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_60_ (
  .in1({ S1976, S1973 }),
  .out1({ S1977 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_61_ (
  .in1({ S1977, S1975 }),
  .out1({ S2536[2] })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_62_ (
  .in1({ S1949, S1290 }),
  .out1({ S1978 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_60_ (
  .in1({ S1950, CU_inst_3 }),
  .out1({ S1979 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_63_ (
  .in1({ S1979, S1958 }),
  .out1({ S1980 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_61_ (
  .in1({ S1958, DP_INC_1_in_3 }),
  .out1({ S1981 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_64_ (
  .in1({ S1874, DP_IN_q_3 }),
  .out1({ S1982 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_62_ (
  .in1({ S1981, S1874 }),
  .out1({ S1983 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_65_ (
  .in1({ S1983, S1980 }),
  .out1({ S1984 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_66_ (
  .in1({ S1984, S1982 }),
  .out1({ S2536[3] })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_67_ (
  .in1({ S1928, S1366 }),
  .out1({ S1985 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_63_ (
  .in1({ S1929, CU_inst_4 }),
  .out1({ S1986 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_68_ (
  .in1({ S1947, S1290 }),
  .out1({ S1987 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_64_ (
  .in1({ S1948, CU_inst_3 }),
  .out1({ S1988 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_69_ (
  .in1({ S1987, S1985 }),
  .out1({ S1989 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_65_ (
  .in1({ S1988, S1986 }),
  .out1({ S1990 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_70_ (
  .in1({ S1958, CU_inst_4 }),
  .out1({ S1991 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_71_ (
  .in1({ S1957, DP_INC_1_in_4 }),
  .out1({ S1992 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_72_ (
  .in1({ S1992, S1991 }),
  .out1({ S1993 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_73_ (
  .in1({ S1993, S1875 }),
  .out1({ S1994 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_74_ (
  .in1({ S1874, DP_IN_q_4 }),
  .out1({ S1995 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_75_ (
  .in1({ S1995, S1994 }),
  .out1({ S2536[4] })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_66_ (
  .in1({ S1929, CU_inst_5 }),
  .out1({ S1996 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_67_ (
  .in1({ S1996, S1988 }),
  .out1({ S1997 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_76_ (
  .in1({ S1997, S1958 }),
  .out1({ S1998 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_77_ (
  .in1({ S1957, DP_INC_1_in_5 }),
  .out1({ S1999 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_78_ (
  .in1({ S1999, S1998 }),
  .out1({ S2000 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_79_ (
  .in1({ S2000, S1875 }),
  .out1({ S2001 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_80_ (
  .in1({ S1874, DP_IN_q_5 }),
  .out1({ S2002 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_81_ (
  .in1({ S2002, S2001 }),
  .out1({ S2536[5] })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_68_ (
  .in1({ S1929, CU_inst_6 }),
  .out1({ S2003 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_69_ (
  .in1({ S2003, S1988 }),
  .out1({ S2004 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_82_ (
  .in1({ S1958, CU_inst_6 }),
  .out1({ S2005 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_83_ (
  .in1({ S1957, DP_INC_1_in_6 }),
  .out1({ S2006 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_84_ (
  .in1({ S2006, S2005 }),
  .out1({ S2007 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_85_ (
  .in1({ S2007, S1875 }),
  .out1({ S2008 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_86_ (
  .in1({ S1874, DP_IN_q_6 }),
  .out1({ S2009 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_87_ (
  .in1({ S2009, S2008 }),
  .out1({ S2536[6] })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_70_ (
  .in1({ S1929, CU_inst_7 }),
  .out1({ S2010 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_71_ (
  .in1({ S2010, S1988 }),
  .out1({ S2011 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_88_ (
  .in1({ S1958, CU_inst_7 }),
  .out1({ S2012 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_89_ (
  .in1({ S1957, DP_INC_1_in_7 }),
  .out1({ S2013 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_90_ (
  .in1({ S2013, S2012 }),
  .out1({ S2014 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_91_ (
  .in1({ S2014, S1875 }),
  .out1({ S2015 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_92_ (
  .in1({ S1874, DP_IN_q_7 }),
  .out1({ S2016 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_93_ (
  .in1({ S2016, S2015 }),
  .out1({ S2536[7] })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_72_ (
  .in1({ S1929, CU_inst_8 }),
  .out1({ S2017 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_73_ (
  .in1({ S2017, S1988 }),
  .out1({ S2018 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_74_ (
  .in1({ S2018, S1957 }),
  .out1({ S2019 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_75_ (
  .in1({ S1958, DP_INC_1_in_8 }),
  .out1({ S2020 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_76_ (
  .in1({ S2020, S2019 }),
  .out1({ S2021 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_77_ (
  .in1({ S2021, S1874 }),
  .out1({ S2022 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_78_ (
  .in1({ S1875, DP_IN_q_8 }),
  .out1({ S2023 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_79_ (
  .in1({ S2023, S2022 }),
  .out1({ S2536[8] })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_80_ (
  .in1({ S1929, CU_inst_9 }),
  .out1({ S2024 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_81_ (
  .in1({ S2024, S1988 }),
  .out1({ S2025 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_82_ (
  .in1({ S2025, S1957 }),
  .out1({ S2026 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_83_ (
  .in1({ S1958, DP_INC_1_in_9 }),
  .out1({ S2027 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_84_ (
  .in1({ S2027, S2026 }),
  .out1({ S2028 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_85_ (
  .in1({ S2028, S1874 }),
  .out1({ S2029 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_86_ (
  .in1({ S1875, DP_IN_q_9 }),
  .out1({ S2030 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_87_ (
  .in1({ S2030, S2029 }),
  .out1({ S2536[9] })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_88_ (
  .in1({ S1929, CU_inst_10 }),
  .out1({ S2031 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_89_ (
  .in1({ S2031, S1988 }),
  .out1({ S2032 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_90_ (
  .in1({ S2032, S1957 }),
  .out1({ S2033 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_91_ (
  .in1({ S1958, DP_INC_1_in_10 }),
  .out1({ S2034 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_92_ (
  .in1({ S2034, S2033 }),
  .out1({ S2035 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_93_ (
  .in1({ S2035, S1874 }),
  .out1({ S2036 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_94_ (
  .in1({ S1875, DP_IN_q_10 }),
  .out1({ S2037 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_95_ (
  .in1({ S2037, S2036 }),
  .out1({ S2536[10] })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_96_ (
  .in1({ S1929, CU_inst_11 }),
  .out1({ S2038 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_97_ (
  .in1({ S2038, S1988 }),
  .out1({ S2039 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_75_ (
  .in1({ S2039 }),
  .out1({ S2040 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_98_ (
  .in1({ S2039, S1957 }),
  .out1({ S2041 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_99_ (
  .in1({ S1958, DP_INC_1_in_11 }),
  .out1({ S2042 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_100_ (
  .in1({ S2042, S2041 }),
  .out1({ S2043 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_101_ (
  .in1({ S2043, S1874 }),
  .out1({ S2044 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_102_ (
  .in1({ S1875, DP_IN_q_11 }),
  .out1({ S2045 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_103_ (
  .in1({ S2045, S2044 }),
  .out1({ S2536[11] })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_94_ (
  .in1({ S1912, DP_IMM1_in1_0 }),
  .out1({ S2046 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_104_ (
  .in1({ S1912, S1143 }),
  .out1({ S2047 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_105_ (
  .in1({ S2047, S1947 }),
  .out1({ S2048 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_95_ (
  .in1({ S2048, S2046 }),
  .out1({ S2049 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_96_ (
  .in1({ S2049, S1987 }),
  .out1({ S2050 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_106_ (
  .in1({ S2050, S1957 }),
  .out1({ S2051 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_97_ (
  .in1({ S1957, DP_INC_1_in_12 }),
  .out1({ S2052 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_107_ (
  .in1({ S1875, DP_IN_q_12 }),
  .out1({ S2053 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_98_ (
  .in1({ S2052, S1875 }),
  .out1({ S2054 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_108_ (
  .in1({ S2054, S2051 }),
  .out1({ S2055 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_109_ (
  .in1({ S2055, S2053 }),
  .out1({ S2536[12] })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_99_ (
  .in1({ S1912, DP_IMM1_in1_1 }),
  .out1({ S2056 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_100_ (
  .in1({ S2056, S2048 }),
  .out1({ S2057 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_101_ (
  .in1({ S2057, S1987 }),
  .out1({ S2058 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_102_ (
  .in1({ S2058, S1958 }),
  .out1({ S2059 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_110_ (
  .in1({ S1958, DP_INC_1_in_13 }),
  .out1({ S2060 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_103_ (
  .in1({ S1874, DP_IN_q_13 }),
  .out1({ S2061 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_111_ (
  .in1({ S2060, S1874 }),
  .out1({ S2062 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_104_ (
  .in1({ S2062, S2059 }),
  .out1({ S2063 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_105_ (
  .in1({ S2063, S2061 }),
  .out1({ S2536[13] })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_106_ (
  .in1({ S1912, DP_IMM1_in1_2 }),
  .out1({ S2064 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_107_ (
  .in1({ S2064, S2048 }),
  .out1({ S2065 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_108_ (
  .in1({ S2065, S1987 }),
  .out1({ S2066 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_76_ (
  .in1({ S2066 }),
  .out1({ S2067 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_112_ (
  .in1({ S2066, S1957 }),
  .out1({ S2068 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_109_ (
  .in1({ S1957, DP_INC_1_in_14 }),
  .out1({ S2069 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_113_ (
  .in1({ S1875, DP_IN_q_14 }),
  .out1({ S2070 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_110_ (
  .in1({ S2069, S1875 }),
  .out1({ S2071 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_114_ (
  .in1({ S2071, S2068 }),
  .out1({ S2072 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_115_ (
  .in1({ S2072, S2070 }),
  .out1({ S2536[14] })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_111_ (
  .in1({ S1912, DP_IMM1_in1_3 }),
  .out1({ S2073 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_112_ (
  .in1({ S2073, S2048 }),
  .out1({ S2074 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_113_ (
  .in1({ S2074, S1987 }),
  .out1({ S2075 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_114_ (
  .in1({ S2075, S1958 }),
  .out1({ S2076 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_116_ (
  .in1({ S1958, DP_INC_1_in_15 }),
  .out1({ S2077 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_115_ (
  .in1({ S1874, DP_IN_q_15 }),
  .out1({ S2078 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_117_ (
  .in1({ S2077, S1874 }),
  .out1({ S2079 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_116_ (
  .in1({ S2079, S2076 }),
  .out1({ S2080 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_117_ (
  .in1({ S2080, S2078 }),
  .out1({ S2536[15] })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_118_ (
  .in1({ S1894, S1825 }),
  .out1({ S2081 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_118_ (
  .in1({ S1893, S1814 }),
  .out1({ S2082 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_119_ (
  .in1({ S2081, S1914 }),
  .out1({ S2083 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_119_ (
  .in1({ S2082, S1915 }),
  .out1({ S2084 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_120_ (
  .in1({ S1895, S1883 }),
  .out1({ S2085 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_77_ (
  .in1({ S2085 }),
  .out1({ S2086 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_120_ (
  .in1({ S1876, S1772 }),
  .out1({ S2087 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_121_ (
  .in1({ S2087, S1883 }),
  .out1({ S2088 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_121_ (
  .in1({ S2085, S1880 }),
  .out1({ S2089 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_122_ (
  .in1({ DP_SR_V_q, S1176 }),
  .out1({ S2090 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_122_ (
  .in1({ DP_SR_V_q, S1176 }),
  .out1({ S2091 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_123_ (
  .in1({ S2090, CU_inst_4 }),
  .out1({ S2092 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_123_ (
  .in1({ S2092, S2091 }),
  .out1({ S2093 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_124_ (
  .in1({ DP_SR_Z_q, S1290 }),
  .out1({ S2094 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_124_ (
  .in1({ DP_SR_Z_q, S1290 }),
  .out1({ S2095 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_125_ (
  .in1({ S2094, CU_inst_7 }),
  .out1({ S2096 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_125_ (
  .in1({ S2096, S2095 }),
  .out1({ S2097 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_126_ (
  .in1({ S2097, S2093 }),
  .out1({ S2098 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_127_ (
  .in1({ S1721, CU_inst_2 }),
  .out1({ S2099 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_126_ (
  .in1({ S1721, CU_inst_2 }),
  .out1({ S2100 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_127_ (
  .in1({ S2100, CU_inst_6 }),
  .out1({ S2101 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_128_ (
  .in1({ S2101, S2099 }),
  .out1({ S2102 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_129_ (
  .in1({ S1710, CU_inst_1 }),
  .out1({ S2103 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_128_ (
  .in1({ S1710, CU_inst_1 }),
  .out1({ S2104 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_129_ (
  .in1({ S2104, CU_inst_5 }),
  .out1({ S2105 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_130_ (
  .in1({ S2105, S2103 }),
  .out1({ S2106 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_131_ (
  .in1({ S2106, S2102 }),
  .out1({ S2107 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_130_ (
  .in1({ S2107, S2098 }),
  .out1({ S2108 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_132_ (
  .in1({ S1132, CU_inst_9 }),
  .out1({ S2109 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_133_ (
  .in1({ CU_inst_10, S1143 }),
  .out1({ S2110 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_131_ (
  .in1({ S2110, S2109 }),
  .out1({ S2111 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_132_ (
  .in1({ S2108, S1930 }),
  .out1({ S2112 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_134_ (
  .in1({ S2112, S2111 }),
  .out1({ S2113 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_78_ (
  .in1({ S2113 }),
  .out1({ S2114 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_133_ (
  .in1({ S2114, S1583 }),
  .out1({ S2115 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_79_ (
  .in1({ S2115 }),
  .out1({ S2116 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_134_ (
  .in1({ S2113, DP_INC_1_in_0 }),
  .out1({ S2117 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_135_ (
  .in1({ S2117, S2115 }),
  .out1({ S2118 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_136_ (
  .in1({ S2118, S2088 }),
  .out1({ S2119 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_137_ (
  .in1({ S2089, DP_AC_q_0 }),
  .out1({ S2120 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_138_ (
  .in1({ S2120, S2119 }),
  .out1({ S2121 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_139_ (
  .in1({ S2121, S2083 }),
  .out1({ S2122 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_140_ (
  .in1({ S2084, DP_IN_q_0 }),
  .out1({ S2123 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_141_ (
  .in1({ S2123, S2122 }),
  .out1({ S2539[0] })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_135_ (
  .in1({ S2116, S1594 }),
  .out1({ S2124 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_80_ (
  .in1({ S2124 }),
  .out1({ S2125 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_136_ (
  .in1({ S2115, DP_INC_1_in_1 }),
  .out1({ S2126 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_137_ (
  .in1({ S2126, S2124 }),
  .out1({ S2127 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_142_ (
  .in1({ S2127, S2088 }),
  .out1({ S2128 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_143_ (
  .in1({ S2089, DP_AC_q_1 }),
  .out1({ S2129 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_144_ (
  .in1({ S2129, S2128 }),
  .out1({ S2130 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_145_ (
  .in1({ S2130, S2083 }),
  .out1({ S2131 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_146_ (
  .in1({ S2084, DP_IN_q_1 }),
  .out1({ S2132 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_147_ (
  .in1({ S2132, S2131 }),
  .out1({ S2539[1] })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_138_ (
  .in1({ S2125, S1604 }),
  .out1({ S2133 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_81_ (
  .in1({ S2133 }),
  .out1({ S2134 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_139_ (
  .in1({ S2124, DP_INC_1_in_2 }),
  .out1({ S2135 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_140_ (
  .in1({ S2135, S2133 }),
  .out1({ S2136 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_141_ (
  .in1({ S2136, S2089 }),
  .out1({ S2137 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_142_ (
  .in1({ S2088, DP_AC_q_2 }),
  .out1({ S2138 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_143_ (
  .in1({ S2138, S2137 }),
  .out1({ S2139 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_144_ (
  .in1({ S2139, S2084 }),
  .out1({ S2140 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_145_ (
  .in1({ S2083, DP_IN_q_2 }),
  .out1({ S2141 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_146_ (
  .in1({ S2141, S2140 }),
  .out1({ S2539[2] })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_147_ (
  .in1({ S2134, S1615 }),
  .out1({ S2142 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_148_ (
  .in1({ S2133, DP_INC_1_in_3 }),
  .out1({ S2143 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_148_ (
  .in1({ S2133, DP_INC_1_in_3 }),
  .out1({ S2144 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_149_ (
  .in1({ S2144, S2142 }),
  .out1({ S2145 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_150_ (
  .in1({ S2145, S2089 }),
  .out1({ S2146 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_151_ (
  .in1({ S2088, DP_AC_q_3 }),
  .out1({ S2147 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_152_ (
  .in1({ S2147, S2146 }),
  .out1({ S2148 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_153_ (
  .in1({ S2148, S2084 }),
  .out1({ S2149 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_154_ (
  .in1({ S2083, DP_IN_q_3 }),
  .out1({ S2150 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_155_ (
  .in1({ S2150, S2149 }),
  .out1({ S2539[3] })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_149_ (
  .in1({ S2084, DP_IN_q_4 }),
  .out1({ S2151 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_156_ (
  .in1({ S2143, S1626 }),
  .out1({ S2152 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_150_ (
  .in1({ S2142, DP_INC_1_in_4 }),
  .out1({ S2153 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_151_ (
  .in1({ S2143, S1626 }),
  .out1({ S2154 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_152_ (
  .in1({ S2154, S2153 }),
  .out1({ S2155 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_153_ (
  .in1({ S2155, S2088 }),
  .out1({ S2156 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_157_ (
  .in1({ S2088, DP_AC_q_4 }),
  .out1({ S2157 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_158_ (
  .in1({ S2157, S2084 }),
  .out1({ S2158 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_154_ (
  .in1({ S2158, S2156 }),
  .out1({ S2159 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_155_ (
  .in1({ S2159, S2151 }),
  .out1({ S2539[4] })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_156_ (
  .in1({ S2084, DP_IN_q_5 }),
  .out1({ S2160 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_157_ (
  .in1({ S2152, DP_INC_1_in_5 }),
  .out1({ S2161 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_82_ (
  .in1({ S2161 }),
  .out1({ S2162 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_158_ (
  .in1({ S2153, S1636 }),
  .out1({ S2163 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_159_ (
  .in1({ S2163, S2161 }),
  .out1({ S2164 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_160_ (
  .in1({ S2164, S2088 }),
  .out1({ S2165 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_159_ (
  .in1({ S2088, DP_AC_q_5 }),
  .out1({ S2166 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_160_ (
  .in1({ S2166, S2084 }),
  .out1({ S2167 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_161_ (
  .in1({ S2167, S2165 }),
  .out1({ S2168 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_162_ (
  .in1({ S2168, S2160 }),
  .out1({ S2539[5] })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_163_ (
  .in1({ S2084, DP_IN_q_6 }),
  .out1({ S2169 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_164_ (
  .in1({ S2162, DP_INC_1_in_6 }),
  .out1({ S2170 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_83_ (
  .in1({ S2170 }),
  .out1({ S2171 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_165_ (
  .in1({ S2161, S1647 }),
  .out1({ S2172 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_166_ (
  .in1({ S2172, S2170 }),
  .out1({ S2173 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_167_ (
  .in1({ S2173, S2088 }),
  .out1({ S2174 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_161_ (
  .in1({ S2088, DP_AC_q_6 }),
  .out1({ S2175 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_162_ (
  .in1({ S2175, S2084 }),
  .out1({ S2176 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_168_ (
  .in1({ S2176, S2174 }),
  .out1({ S2177 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_169_ (
  .in1({ S2177, S2169 }),
  .out1({ S2539[6] })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_170_ (
  .in1({ S2084, DP_IN_q_7 }),
  .out1({ S2178 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_171_ (
  .in1({ S2171, DP_INC_1_in_7 }),
  .out1({ S2179 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_84_ (
  .in1({ S2179 }),
  .out1({ S2180 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_172_ (
  .in1({ S2170, S1657 }),
  .out1({ S2181 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_173_ (
  .in1({ S2181, S2179 }),
  .out1({ S2182 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_174_ (
  .in1({ S2182, S2088 }),
  .out1({ S2183 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_163_ (
  .in1({ S2088, DP_AC_q_7 }),
  .out1({ S2184 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_164_ (
  .in1({ S2184, S2084 }),
  .out1({ S2185 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_175_ (
  .in1({ S2185, S2183 }),
  .out1({ S2186 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_176_ (
  .in1({ S2186, S2178 }),
  .out1({ S2539[7] })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_177_ (
  .in1({ S2084, DP_IN_q_8 }),
  .out1({ S2187 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_178_ (
  .in1({ S2180, DP_INC_1_in_8 }),
  .out1({ S2188 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_85_ (
  .in1({ S2188 }),
  .out1({ S2189 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_179_ (
  .in1({ S2179, S1668 }),
  .out1({ S2190 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_180_ (
  .in1({ S2190, S2188 }),
  .out1({ S2191 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_181_ (
  .in1({ S2191, S2088 }),
  .out1({ S2192 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_165_ (
  .in1({ S2088, DP_AC_q_8 }),
  .out1({ S2193 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_166_ (
  .in1({ S2193, S2084 }),
  .out1({ S2194 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_182_ (
  .in1({ S2194, S2192 }),
  .out1({ S2195 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_183_ (
  .in1({ S2195, S2187 }),
  .out1({ S2539[8] })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_184_ (
  .in1({ S2084, DP_IN_q_9 }),
  .out1({ S2196 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_185_ (
  .in1({ S2189, DP_INC_1_in_9 }),
  .out1({ S2197 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_86_ (
  .in1({ S2197 }),
  .out1({ S2198 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_186_ (
  .in1({ S2188, S1679 }),
  .out1({ S2199 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_187_ (
  .in1({ S2199, S2197 }),
  .out1({ S2200 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_188_ (
  .in1({ S2200, S2088 }),
  .out1({ S2201 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_167_ (
  .in1({ S2088, DP_AC_q_9 }),
  .out1({ S2202 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_168_ (
  .in1({ S2202, S2084 }),
  .out1({ S2203 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_189_ (
  .in1({ S2203, S2201 }),
  .out1({ S2204 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_190_ (
  .in1({ S2204, S2196 }),
  .out1({ S2539[9] })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_191_ (
  .in1({ S2084, DP_IN_q_10 }),
  .out1({ S2205 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_169_ (
  .in1({ S2197, S1689 }),
  .out1({ S2206 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_192_ (
  .in1({ S2198, DP_INC_1_in_10 }),
  .out1({ S2207 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_193_ (
  .in1({ S2197, S1689 }),
  .out1({ S2208 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_194_ (
  .in1({ S2208, S2207 }),
  .out1({ S2209 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_195_ (
  .in1({ S2209, S2088 }),
  .out1({ S2210 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_170_ (
  .in1({ S2088, DP_AC_q_10 }),
  .out1({ S2211 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_171_ (
  .in1({ S2211, S2084 }),
  .out1({ S2212 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_196_ (
  .in1({ S2212, S2210 }),
  .out1({ S2213 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_197_ (
  .in1({ S2213, S2205 }),
  .out1({ S2539[10] })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_198_ (
  .in1({ S2084, DP_IN_q_11 }),
  .out1({ S2214 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_172_ (
  .in1({ S2207, S1700 }),
  .out1({ S2215 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_199_ (
  .in1({ S2206, DP_INC_1_in_11 }),
  .out1({ S2216 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_200_ (
  .in1({ S2207, S1700 }),
  .out1({ S2217 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_201_ (
  .in1({ S2217, S2216 }),
  .out1({ S2218 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_202_ (
  .in1({ S2218, S2088 }),
  .out1({ S2219 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_173_ (
  .in1({ S2088, DP_AC_q_11 }),
  .out1({ S2220 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_174_ (
  .in1({ S2220, S2084 }),
  .out1({ S2221 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_203_ (
  .in1({ S2221, S2219 }),
  .out1({ S2222 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_204_ (
  .in1({ S2222, S2214 }),
  .out1({ S2539[11] })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_205_ (
  .in1({ S2084, DP_IN_q_12 }),
  .out1({ S2223 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_175_ (
  .in1({ S2216, S1540 }),
  .out1({ S2224 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_206_ (
  .in1({ S2215, DP_INC_1_in_12 }),
  .out1({ S2225 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_207_ (
  .in1({ S2216, S1540 }),
  .out1({ S2226 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_208_ (
  .in1({ S2226, S2225 }),
  .out1({ S2227 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_209_ (
  .in1({ S2227, S2088 }),
  .out1({ S2228 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_176_ (
  .in1({ S2088, DP_AC_q_12 }),
  .out1({ S2229 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_177_ (
  .in1({ S2229, S2084 }),
  .out1({ S2230 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_210_ (
  .in1({ S2230, S2228 }),
  .out1({ S2231 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_211_ (
  .in1({ S2231, S2223 }),
  .out1({ S2539[12] })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_212_ (
  .in1({ S2084, DP_IN_q_13 }),
  .out1({ S2232 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_213_ (
  .in1({ S2224, DP_INC_1_in_13 }),
  .out1({ S2233 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_87_ (
  .in1({ S2233 }),
  .out1({ S2234 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_214_ (
  .in1({ S2225, S1551 }),
  .out1({ S2235 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_215_ (
  .in1({ S2235, S2233 }),
  .out1({ S2236 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_216_ (
  .in1({ S2236, S2088 }),
  .out1({ S2237 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_178_ (
  .in1({ S2088, DP_AC_q_13 }),
  .out1({ S2238 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_179_ (
  .in1({ S2238, S2084 }),
  .out1({ S2239 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_217_ (
  .in1({ S2239, S2237 }),
  .out1({ S2240 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_218_ (
  .in1({ S2240, S2232 }),
  .out1({ S2539[13] })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_219_ (
  .in1({ S2084, DP_IN_q_14 }),
  .out1({ S2241 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_220_ (
  .in1({ S2234, DP_INC_1_in_14 }),
  .out1({ S2242 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_221_ (
  .in1({ S2233, S1562 }),
  .out1({ S2243 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_222_ (
  .in1({ S2243, S2242 }),
  .out1({ S2244 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_223_ (
  .in1({ S2244, S2088 }),
  .out1({ S2245 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_180_ (
  .in1({ S2088, DP_AC_q_14 }),
  .out1({ S2246 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_181_ (
  .in1({ S2246, S2084 }),
  .out1({ S2247 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_224_ (
  .in1({ S2247, S2245 }),
  .out1({ S2248 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_225_ (
  .in1({ S2248, S2241 }),
  .out1({ S2539[14] })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_226_ (
  .in1({ S2084, DP_IN_q_15 }),
  .out1({ S2249 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_227_ (
  .in1({ S2242, DP_INC_1_in_15 }),
  .out1({ S2250 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_88_ (
  .in1({ S2250 }),
  .out1({ S2251 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_182_ (
  .in1({ S2242, DP_INC_1_in_15 }),
  .out1({ S2252 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_183_ (
  .in1({ S2252, S2251 }),
  .out1({ S2253 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_228_ (
  .in1({ S2253, S2088 }),
  .out1({ S2254 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_184_ (
  .in1({ S2088, DP_AC_q_15 }),
  .out1({ S2255 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_185_ (
  .in1({ S2255, S2084 }),
  .out1({ S2256 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_229_ (
  .in1({ S2256, S2254 }),
  .out1({ S2257 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_230_ (
  .in1({ S2257, S2249 }),
  .out1({ S2539[15] })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_186_ (
  .in1({ S1885, S1762 }),
  .out1({ S2258 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_231_ (
  .in1({ S2258, S1882 }),
  .out1({ S2259 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_187_ (
  .in1({ S2088, S1870 }),
  .out1({ S2260 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_232_ (
  .in1({ S2260, S2259 }),
  .out1({ S2542 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_233_ (
  .in1({ S1876, S1783 }),
  .out1({ S2261 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_234_ (
  .in1({ S2261, S1888 }),
  .out1({ S2262 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_188_ (
  .in1({ S2262, S1907 }),
  .out1({ CU_nstate_1 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_189_ (
  .in1({ S1891, S1877 }),
  .out1({ S2263 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_190_ (
  .in1({ S2263, S2258 }),
  .out1({ S2264 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_235_ (
  .in1({ S2264, S1922 }),
  .out1({ S2265 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_236_ (
  .in1({ S2082, S1846 }),
  .out1({ S2266 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_191_ (
  .in1({ S2266, CU_nstate_0 }),
  .out1({ S2267 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_237_ (
  .in1({ S2267, S2265 }),
  .out1({ S2540 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_238_ (
  .in1({ S2109, S1936 }),
  .out1({ S2268 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_89_ (
  .in1({ S2268 }),
  .out1({ S2269 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_192_ (
  .in1({ S2268, CU_inst_7 }),
  .out1({ S2270 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_239_ (
  .in1({ S2269, S1168 }),
  .out1({ S2271 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_193_ (
  .in1({ CU_inst_6, CU_inst_5 }),
  .out1({ S2272 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_194_ (
  .in1({ S2271, S1917 }),
  .out1({ S2273 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_195_ (
  .in1({ S2271, S1931 }),
  .out1({ S2274 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_240_ (
  .in1({ S2274, S2272 }),
  .out1({ S2275 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_241_ (
  .in1({ S2275, S1945 }),
  .out1({ S2276 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_196_ (
  .in1({ S2276, S1453 }),
  .out1({ S2277 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_242_ (
  .in1({ S2276, S1951 }),
  .out1({ S2278 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_197_ (
  .in1({ S2275, S1540 }),
  .out1({ S2279 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_198_ (
  .in1({ S2279, S2277 }),
  .out1({ S2280 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_243_ (
  .in1({ S2280, S2278 }),
  .out1({ S0 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_199_ (
  .in1({ S2276, S1475 }),
  .out1({ S2281 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_200_ (
  .in1({ S2275, S1551 }),
  .out1({ S2282 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_201_ (
  .in1({ S2282, S2281 }),
  .out1({ S2283 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_244_ (
  .in1({ S2276, S1965 }),
  .out1({ S2284 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_245_ (
  .in1({ S2284, S2283 }),
  .out1({ S1 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_202_ (
  .in1({ S2276, S1497 }),
  .out1({ S2285 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_203_ (
  .in1({ S2275, S1562 }),
  .out1({ S2286 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_204_ (
  .in1({ S2286, S2285 }),
  .out1({ S2287 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_246_ (
  .in1({ S2276, S1972 }),
  .out1({ S2288 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_247_ (
  .in1({ S2288, S2287 }),
  .out1({ S2 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_205_ (
  .in1({ S2276, S1519 }),
  .out1({ S2289 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_206_ (
  .in1({ S2275, S1572 }),
  .out1({ S2290 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_207_ (
  .in1({ S2290, S2289 }),
  .out1({ S2291 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_248_ (
  .in1({ S2276, S1978 }),
  .out1({ S2292 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_249_ (
  .in1({ S2292, S2291 }),
  .out1({ S3 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_208_ (
  .in1({ S1883, S1083 }),
  .out1({ S2293 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_250_ (
  .in1({ S1882, CU_inst_12 }),
  .out1({ S2294 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_209_ (
  .in1({ S2294, S1869 }),
  .out1({ S2295 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_251_ (
  .in1({ S2293, S1868 }),
  .out1({ S2296 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_210_ (
  .in1({ S2295, S2538[0] }),
  .out1({ S2297 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_211_ (
  .in1({ S1908, S1883 }),
  .out1({ S2298 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_252_ (
  .in1({ S1909, S1882 }),
  .out1({ S2299 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_212_ (
  .in1({ S2296, S1183 }),
  .out1({ S2300 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_213_ (
  .in1({ S2300, S2297 }),
  .out1({ S2301 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_253_ (
  .in1({ S2301, S2298 }),
  .out1({ S2302 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_254_ (
  .in1({ S2299, DP_IN_q_0 }),
  .out1({ S2303 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_255_ (
  .in1({ S2303, S2302 }),
  .out1({ S4 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_214_ (
  .in1({ S2300, S2538[1] }),
  .out1({ S2304 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_256_ (
  .in1({ S2538[1], S2538[0] }),
  .out1({ S2305 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_215_ (
  .in1({ S2305, S2296 }),
  .out1({ S2306 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_216_ (
  .in1({ S2306, S2304 }),
  .out1({ S2307 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_257_ (
  .in1({ S2307, S2298 }),
  .out1({ S2308 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_258_ (
  .in1({ S2299, DP_IN_q_1 }),
  .out1({ S2309 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_259_ (
  .in1({ S2309, S2308 }),
  .out1({ S5 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_217_ (
  .in1({ S2306, S2538[2] }),
  .out1({ S2310 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_260_ (
  .in1({ S2306, S2538[2] }),
  .out1({ S2311 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_261_ (
  .in1({ S2295, S2538[2] }),
  .out1({ S2312 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_218_ (
  .in1({ S2312, S2305 }),
  .out1({ S2313 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_219_ (
  .in1({ S2313, S2310 }),
  .out1({ S2314 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_220_ (
  .in1({ S2314, S2299 }),
  .out1({ S2315 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_221_ (
  .in1({ S2298, DP_IN_q_2 }),
  .out1({ S2316 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_222_ (
  .in1({ S2316, S2315 }),
  .out1({ S6 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_223_ (
  .in1({ S2313, S2538[3] }),
  .out1({ S2317 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_224_ (
  .in1({ S2311, S1279 }),
  .out1({ S2318 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_225_ (
  .in1({ S2318, S2317 }),
  .out1({ S2319 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_226_ (
  .in1({ S2319, S2299 }),
  .out1({ S2320 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_227_ (
  .in1({ S2298, DP_IN_q_3 }),
  .out1({ S2321 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_228_ (
  .in1({ S2321, S2320 }),
  .out1({ S7 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_262_ (
  .in1({ S2318, S2538[4] }),
  .out1({ S2322 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_90_ (
  .in1({ S2322 }),
  .out1({ S2323 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_229_ (
  .in1({ S2318, S2538[4] }),
  .out1({ S2324 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_230_ (
  .in1({ S2324, S2323 }),
  .out1({ S2325 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_231_ (
  .in1({ S2325, S2299 }),
  .out1({ S2326 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_232_ (
  .in1({ S2298, DP_IN_q_4 }),
  .out1({ S2327 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_233_ (
  .in1({ S2327, S2326 }),
  .out1({ S8 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_263_ (
  .in1({ S2322, S1388 }),
  .out1({ S2328 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_234_ (
  .in1({ S2322, S1388 }),
  .out1({ S2329 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_235_ (
  .in1({ S2329, S2299 }),
  .out1({ S2330 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_264_ (
  .in1({ S2330, S2328 }),
  .out1({ S2331 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_265_ (
  .in1({ S2299, DP_IN_q_5 }),
  .out1({ S2332 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_266_ (
  .in1({ S2332, S2331 }),
  .out1({ S9 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_236_ (
  .in1({ S2329, S2538[6] }),
  .out1({ S2333 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_267_ (
  .in1({ S2329, S2538[6] }),
  .out1({ S2334 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_91_ (
  .in1({ S2334 }),
  .out1({ S2335 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_237_ (
  .in1({ S2335, S2333 }),
  .out1({ S2336 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_238_ (
  .in1({ S2336, S2299 }),
  .out1({ S2337 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_239_ (
  .in1({ S2298, DP_IN_q_6 }),
  .out1({ S2338 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_240_ (
  .in1({ S2338, S2337 }),
  .out1({ S10 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_241_ (
  .in1({ S2334, S1410 }),
  .out1({ S2339 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_92_ (
  .in1({ S2339 }),
  .out1({ S2340 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_242_ (
  .in1({ S2335, S2538[7] }),
  .out1({ S2341 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_243_ (
  .in1({ S2341, S2339 }),
  .out1({ S2342 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_268_ (
  .in1({ S2342, S2298 }),
  .out1({ S2343 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_269_ (
  .in1({ S2299, DP_IN_q_7 }),
  .out1({ S2344 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_270_ (
  .in1({ S2344, S2343 }),
  .out1({ S11 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_244_ (
  .in1({ S2339, S2538[8] }),
  .out1({ S2345 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_245_ (
  .in1({ S2340, S1421 }),
  .out1({ S2346 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_271_ (
  .in1({ S2339, S2538[8] }),
  .out1({ S2347 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_246_ (
  .in1({ S2298, DP_IN_q_8 }),
  .out1({ S2348 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_247_ (
  .in1({ S2346, S2345 }),
  .out1({ S2349 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_248_ (
  .in1({ S2349, S2299 }),
  .out1({ S2350 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_249_ (
  .in1({ S2350, S2348 }),
  .out1({ S12 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_272_ (
  .in1({ S2299, DP_IN_q_9 }),
  .out1({ S2351 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_273_ (
  .in1({ S2346, S2538[9] }),
  .out1({ S2352 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_250_ (
  .in1({ S2346, S2538[9] }),
  .out1({ S2353 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_251_ (
  .in1({ S2353, S2299 }),
  .out1({ S2354 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_274_ (
  .in1({ S2354, S2352 }),
  .out1({ S2355 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_275_ (
  .in1({ S2355, S2351 }),
  .out1({ S13 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_276_ (
  .in1({ S2352, S1432 }),
  .out1({ S2356 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_252_ (
  .in1({ S2352, S1432 }),
  .out1({ S2357 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_277_ (
  .in1({ S2538[10], S2538[9] }),
  .out1({ S2358 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_253_ (
  .in1({ S2358, S2347 }),
  .out1({ S2359 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_93_ (
  .in1({ S2359 }),
  .out1({ S2360 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_254_ (
  .in1({ S2359, S2299 }),
  .out1({ S2361 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_278_ (
  .in1({ S2361, S2356 }),
  .out1({ S2362 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_279_ (
  .in1({ S2299, DP_IN_q_10 }),
  .out1({ S2363 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_280_ (
  .in1({ S2363, S2362 }),
  .out1({ S14 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_255_ (
  .in1({ S2359, S2538[11] }),
  .out1({ S2364 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_281_ (
  .in1({ S2357, S2538[11] }),
  .out1({ S2365 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_256_ (
  .in1({ S2298, DP_IN_q_11 }),
  .out1({ S2366 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_257_ (
  .in1({ S2360, S1443 }),
  .out1({ S2367 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_258_ (
  .in1({ S2367, S2364 }),
  .out1({ S2368 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_259_ (
  .in1({ S2368, S2299 }),
  .out1({ S2369 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_260_ (
  .in1({ S2369, S2366 }),
  .out1({ S15 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_261_ (
  .in1({ S2298, DP_IN_q_12 }),
  .out1({ S2370 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_262_ (
  .in1({ S2367, S2538[12] }),
  .out1({ S2371 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_263_ (
  .in1({ S2365, S1464 }),
  .out1({ S2372 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_264_ (
  .in1({ S2372, S2371 }),
  .out1({ S2373 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_265_ (
  .in1({ S2373, S2299 }),
  .out1({ S2374 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_282_ (
  .in1({ S2538[12], S2538[11] }),
  .out1({ S2375 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_94_ (
  .in1({ S2375 }),
  .out1({ S2376 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_283_ (
  .in1({ S2376, S2359 }),
  .out1({ S2377 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_266_ (
  .in1({ S2374, S2370 }),
  .out1({ S16 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_284_ (
  .in1({ S2299, DP_IN_q_13 }),
  .out1({ S2378 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_267_ (
  .in1({ S2372, S2538[13] }),
  .out1({ S2379 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_268_ (
  .in1({ S2377, S1486 }),
  .out1({ S2380 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_269_ (
  .in1({ S2380, S2379 }),
  .out1({ S2381 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_285_ (
  .in1({ S2381, S2298 }),
  .out1({ S2382 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_286_ (
  .in1({ S2382, S2378 }),
  .out1({ S17 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_270_ (
  .in1({ S2298, DP_IN_q_14 }),
  .out1({ S2383 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_271_ (
  .in1({ S2380, S2538[14] }),
  .out1({ S2384 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_287_ (
  .in1({ S2380, S2538[14] }),
  .out1({ S2385 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_95_ (
  .in1({ S2385 }),
  .out1({ S2386 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_272_ (
  .in1({ S2386, S2384 }),
  .out1({ S2387 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_273_ (
  .in1({ S2387, S2299 }),
  .out1({ S2388 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_274_ (
  .in1({ S2388, S2383 }),
  .out1({ S18 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_275_ (
  .in1({ S2298, DP_IN_q_15 }),
  .out1({ S2389 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_276_ (
  .in1({ S2385, S1529 }),
  .out1({ S2390 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_277_ (
  .in1({ S2386, S2538[15] }),
  .out1({ S2391 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_278_ (
  .in1({ S2391, S2390 }),
  .out1({ S2392 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_279_ (
  .in1({ S2392, S2299 }),
  .out1({ S2393 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_280_ (
  .in1({ S2393, S2389 }),
  .out1({ S19 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_288_ (
  .in1({ S2270, CU_inst_6 }),
  .out1({ S2394 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_289_ (
  .in1({ S2273, CU_inst_6 }),
  .out1({ S2395 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_290_ (
  .in1({ S2395, S1903 }),
  .out1({ S2396 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_291_ (
  .in1({ S2396, S1882 }),
  .out1({ S2397 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_281_ (
  .in1({ CU_inst_8, S1123 }),
  .out1({ S2398 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_292_ (
  .in1({ S2398, S1933 }),
  .out1({ S2399 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_282_ (
  .in1({ S2399, S1931 }),
  .out1({ S2400 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_96_ (
  .in1({ S2400 }),
  .out1({ S2401 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_293_ (
  .in1({ S2400, CU_inst_6 }),
  .out1({ S2402 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_97_ (
  .in1({ S2402 }),
  .out1({ S2403 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_283_ (
  .in1({ S2399, S1917 }),
  .out1({ S2404 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_284_ (
  .in1({ S2403, S2081 }),
  .out1({ S2405 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_294_ (
  .in1({ S2405, S2397 }),
  .out1({ S2406 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_285_ (
  .in1({ S2406, DP_SR_N_q }),
  .out1({ S2407 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_295_ (
  .in1({ S2394, S1916 }),
  .out1({ S2408 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_286_ (
  .in1({ S2086, S1880 }),
  .out1({ S2409 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_296_ (
  .in1({ S2409, S2408 }),
  .out1({ S2410 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_297_ (
  .in1({ S2410, S2401 }),
  .out1({ S2411 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_98_ (
  .in1({ S2411 }),
  .out1({ S2412 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_287_ (
  .in1({ S1884, S1877 }),
  .out1({ S2413 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_288_ (
  .in1({ S2413, S1918 }),
  .out1({ S2414 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_289_ (
  .in1({ S2268, S1168 }),
  .out1({ S2415 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_298_ (
  .in1({ S2415, S2272 }),
  .out1({ S2416 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_99_ (
  .in1({ S2416 }),
  .out1({ S2417 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_299_ (
  .in1({ S2416, S1916 }),
  .out1({ S2418 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_300_ (
  .in1({ S1884, S1878 }),
  .out1({ S2419 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_290_ (
  .in1({ S2413, S1883 }),
  .out1({ S2420 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_291_ (
  .in1({ S1909, S1883 }),
  .out1({ S2421 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_100_ (
  .in1({ S2421 }),
  .out1({ S2422 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_292_ (
  .in1({ S2413, S2258 }),
  .out1({ S2423 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_301_ (
  .in1({ S2423, S2421 }),
  .out1({ S2424 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_293_ (
  .in1({ S1899, S1889 }),
  .out1({ S2425 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_302_ (
  .in1({ S2425, S2418 }),
  .out1({ S2426 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_294_ (
  .in1({ S2426, S2424 }),
  .out1({ S2427 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_101_ (
  .in1({ S2427 }),
  .out1({ S2428 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_303_ (
  .in1({ S2427, S2419 }),
  .out1({ S2429 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_102_ (
  .in1({ S2429 }),
  .out1({ S2430 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_295_ (
  .in1({ S2430, S2081 }),
  .out1({ S2431 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_304_ (
  .in1({ S2429, S2082 }),
  .out1({ S2432 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_296_ (
  .in1({ S2416, S1931 }),
  .out1({ S2433 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_305_ (
  .in1({ S2417, S1930 }),
  .out1({ S2434 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_297_ (
  .in1({ S1941, S1917 }),
  .out1({ S2435 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_103_ (
  .in1({ S2435 }),
  .out1({ S2436 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_306_ (
  .in1({ S2436, S2414 }),
  .out1({ S2437 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_298_ (
  .in1({ S2435, S1911 }),
  .out1({ S2438 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_299_ (
  .in1({ S2437, S1911 }),
  .out1({ S2439 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_307_ (
  .in1({ S2438, S2414 }),
  .out1({ S2440 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_300_ (
  .in1({ S2440, S2067 }),
  .out1({ S2441 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_308_ (
  .in1({ S2439, S2066 }),
  .out1({ S2442 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_301_ (
  .in1({ S2439, S2538[15] }),
  .out1({ S2443 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_302_ (
  .in1({ S2443, S2441 }),
  .out1({ S2444 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_309_ (
  .in1({ S2444, S2434 }),
  .out1({ S2445 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_303_ (
  .in1({ S2445, S1356 }),
  .out1({ S2446 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_104_ (
  .in1({ S2446 }),
  .out1({ S2447 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_310_ (
  .in1({ S2445, S1356 }),
  .out1({ S2448 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_311_ (
  .in1({ S2448, S2447 }),
  .out1({ S2449 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_312_ (
  .in1({ S2440, S1508 }),
  .out1({ S2450 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_313_ (
  .in1({ S2450, S2442 }),
  .out1({ S2451 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_304_ (
  .in1({ S2451, S2433 }),
  .out1({ S2452 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_305_ (
  .in1({ S2451, S1345 }),
  .out1({ S2453 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_105_ (
  .in1({ S2453 }),
  .out1({ S2454 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_306_ (
  .in1({ S2454, S2433 }),
  .out1({ S2455 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_307_ (
  .in1({ S2452, DP_AC_q_14 }),
  .out1({ S2456 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_308_ (
  .in1({ S2456, S2455 }),
  .out1({ S2457 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_106_ (
  .in1({ S2457 }),
  .out1({ S2458 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_309_ (
  .in1({ S2439, S2538[13] }),
  .out1({ S2459 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_310_ (
  .in1({ S2459, S2441 }),
  .out1({ S2460 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_107_ (
  .in1({ S2460 }),
  .out1({ S2461 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_314_ (
  .in1({ S2460, S2434 }),
  .out1({ S2462 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_311_ (
  .in1({ S2461, S1334 }),
  .out1({ S2463 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_312_ (
  .in1({ S2462, S1334 }),
  .out1({ S2464 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_315_ (
  .in1({ S2463, S2434 }),
  .out1({ S2465 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_316_ (
  .in1({ S2462, S1334 }),
  .out1({ S2466 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_317_ (
  .in1({ S2466, S2465 }),
  .out1({ S2467 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_108_ (
  .in1({ S2467 }),
  .out1({ S2468 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_313_ (
  .in1({ S2439, S2538[12] }),
  .out1({ S2469 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_314_ (
  .in1({ S2469, S2441 }),
  .out1({ S2470 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_109_ (
  .in1({ S2470 }),
  .out1({ S2471 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_315_ (
  .in1({ S2471, S2433 }),
  .out1({ S2472 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_318_ (
  .in1({ S2472, DP_AC_q_12 }),
  .out1({ S2473 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_110_ (
  .in1({ S2473 }),
  .out1({ S2474 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_316_ (
  .in1({ S2472, DP_AC_q_12 }),
  .out1({ S2475 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_317_ (
  .in1({ S2475, S2474 }),
  .out1({ S2476 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_111_ (
  .in1({ S2476 }),
  .out1({ S2477 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_318_ (
  .in1({ S2439, S2538[11] }),
  .out1({ S2478 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_319_ (
  .in1({ S2478, S2441 }),
  .out1({ S2479 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_112_ (
  .in1({ S2479 }),
  .out1({ S2480 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_320_ (
  .in1({ S2480, S2433 }),
  .out1({ S2481 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_319_ (
  .in1({ S2479, S2434 }),
  .out1({ S2482 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_321_ (
  .in1({ S2482, S1323 }),
  .out1({ S2483 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_322_ (
  .in1({ S2481, DP_AC_q_11 }),
  .out1({ S2484 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_323_ (
  .in1({ S2484, S2483 }),
  .out1({ S2485 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_113_ (
  .in1({ S2485 }),
  .out1({ S2486 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_324_ (
  .in1({ S2440, S2032 }),
  .out1({ S2487 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_325_ (
  .in1({ S2439, S2538[10] }),
  .out1({ S2488 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_326_ (
  .in1({ S2488, S2487 }),
  .out1({ S2489 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_114_ (
  .in1({ S2489 }),
  .out1({ S2490 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_327_ (
  .in1({ S2490, S2433 }),
  .out1({ S2491 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_320_ (
  .in1({ S2489, S2434 }),
  .out1({ S2492 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_328_ (
  .in1({ S2492, S1312 }),
  .out1({ S2493 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_329_ (
  .in1({ S2491, DP_AC_q_10 }),
  .out1({ S2494 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_330_ (
  .in1({ S2494, S2493 }),
  .out1({ S2495 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_331_ (
  .in1({ S2440, S2025 }),
  .out1({ S2496 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_332_ (
  .in1({ S2439, S2538[9] }),
  .out1({ S2497 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_333_ (
  .in1({ S2497, S2496 }),
  .out1({ S2498 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_115_ (
  .in1({ S2498 }),
  .out1({ S2499 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_334_ (
  .in1({ S2499, S2433 }),
  .out1({ S2500 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_321_ (
  .in1({ S2498, S2434 }),
  .out1({ S2501 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_335_ (
  .in1({ S2501, S1301 }),
  .out1({ S2502 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_336_ (
  .in1({ S2500, DP_AC_q_9 }),
  .out1({ S2503 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_337_ (
  .in1({ S2440, S2018 }),
  .out1({ S2504 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_338_ (
  .in1({ S2439, S2538[8] }),
  .out1({ S2505 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_339_ (
  .in1({ S2505, S2504 }),
  .out1({ S2506 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_116_ (
  .in1({ S2506 }),
  .out1({ S2507 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_340_ (
  .in1({ S2507, S2433 }),
  .out1({ S2508 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_322_ (
  .in1({ S2508, DP_AC_q_8 }),
  .out1({ S2509 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_117_ (
  .in1({ S2509 }),
  .out1({ S2510 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_341_ (
  .in1({ S2508, DP_AC_q_8 }),
  .out1({ S2511 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_118_ (
  .in1({ S2511 }),
  .out1({ S2512 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_342_ (
  .in1({ S2511, S2510 }),
  .out1({ S2513 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_323_ (
  .in1({ S2512, S2509 }),
  .out1({ S2514 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_343_ (
  .in1({ S2440, S2011 }),
  .out1({ S2515 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_344_ (
  .in1({ S2439, S2538[7] }),
  .out1({ S2516 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_345_ (
  .in1({ S2516, S2515 }),
  .out1({ S2517 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_119_ (
  .in1({ S2517 }),
  .out1({ S2518 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_346_ (
  .in1({ S2518, S2433 }),
  .out1({ S2519 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_324_ (
  .in1({ S2517, S2434 }),
  .out1({ S2520 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_325_ (
  .in1({ S2517, DP_AC_q_7 }),
  .out1({ S2521 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_347_ (
  .in1({ S2520, S1268 }),
  .out1({ S2522 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_326_ (
  .in1({ S2519, DP_AC_q_7 }),
  .out1({ S2523 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_348_ (
  .in1({ S2519, DP_AC_q_7 }),
  .out1({ S2524 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_349_ (
  .in1({ S2524, S2522 }),
  .out1({ S2525 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_120_ (
  .in1({ S2525 }),
  .out1({ S2526 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_350_ (
  .in1({ S2440, S2004 }),
  .out1({ S2527 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_121_ (
  .in1({ S2527 }),
  .out1({ S2528 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_327_ (
  .in1({ S2440, S1399 }),
  .out1({ S2529 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_328_ (
  .in1({ S2529, S2528 }),
  .out1({ S2530 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_122_ (
  .in1({ S2530 }),
  .out1({ S2531 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_351_ (
  .in1({ S2530, S2433 }),
  .out1({ S2532 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_329_ (
  .in1({ S2531, S2434 }),
  .out1({ S2533 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_352_ (
  .in1({ S2533, S1257 }),
  .out1({ S2534 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_330_ (
  .in1({ S2532, DP_AC_q_6 }),
  .out1({ S2535 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_353_ (
  .in1({ S2532, DP_AC_q_6 }),
  .out1({ S72 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_123_ (
  .in1({ S72 }),
  .out1({ S73 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_354_ (
  .in1({ S72, S2534 }),
  .out1({ S74 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_331_ (
  .in1({ S73, S2535 }),
  .out1({ S75 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_355_ (
  .in1({ S2440, S1997 }),
  .out1({ S76 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_356_ (
  .in1({ S2439, S2538[5] }),
  .out1({ S77 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_357_ (
  .in1({ S77, S76 }),
  .out1({ S78 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_124_ (
  .in1({ S78 }),
  .out1({ S79 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_358_ (
  .in1({ S79, S2433 }),
  .out1({ S80 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_332_ (
  .in1({ S78, S2434 }),
  .out1({ S81 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_333_ (
  .in1({ S78, DP_AC_q_5 }),
  .out1({ S82 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_125_ (
  .in1({ S82 }),
  .out1({ S83 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_359_ (
  .in1({ S81, S1246 }),
  .out1({ S84 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_334_ (
  .in1({ S80, DP_AC_q_5 }),
  .out1({ S85 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_360_ (
  .in1({ S80, DP_AC_q_5 }),
  .out1({ S86 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_335_ (
  .in1({ S2440, S2538[4] }),
  .out1({ S87 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_126_ (
  .in1({ S87 }),
  .out1({ S88 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_361_ (
  .in1({ S2440, S1989 }),
  .out1({ S89 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_336_ (
  .in1({ S2439, S1990 }),
  .out1({ S90 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_337_ (
  .in1({ S90, S87 }),
  .out1({ S91 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_362_ (
  .in1({ S89, S88 }),
  .out1({ S92 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_363_ (
  .in1({ S92, S2433 }),
  .out1({ S93 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_338_ (
  .in1({ S91, S2434 }),
  .out1({ S94 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_364_ (
  .in1({ S92, S1235 }),
  .out1({ S95 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_339_ (
  .in1({ S91, DP_AC_q_4 }),
  .out1({ S96 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_365_ (
  .in1({ S94, S1235 }),
  .out1({ S97 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_340_ (
  .in1({ S93, DP_AC_q_4 }),
  .out1({ S98 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_366_ (
  .in1({ S93, DP_AC_q_4 }),
  .out1({ S99 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_127_ (
  .in1({ S99 }),
  .out1({ S100 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_367_ (
  .in1({ S99, S97 }),
  .out1({ S101 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_341_ (
  .in1({ S100, S98 }),
  .out1({ S102 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_368_ (
  .in1({ S2440, S1979 }),
  .out1({ S103 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_342_ (
  .in1({ S2439, S1978 }),
  .out1({ S104 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_343_ (
  .in1({ S2440, S2538[3] }),
  .out1({ S105 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_128_ (
  .in1({ S105 }),
  .out1({ S106 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_344_ (
  .in1({ S105, S104 }),
  .out1({ S107 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_369_ (
  .in1({ S106, S103 }),
  .out1({ S108 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_370_ (
  .in1({ S108, S2433 }),
  .out1({ S109 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_345_ (
  .in1({ S107, S2434 }),
  .out1({ S110 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_371_ (
  .in1({ S108, S1224 }),
  .out1({ S111 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_346_ (
  .in1({ S107, DP_AC_q_3 }),
  .out1({ S112 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_372_ (
  .in1({ S110, S1224 }),
  .out1({ S113 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_347_ (
  .in1({ S109, DP_AC_q_3 }),
  .out1({ S114 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_373_ (
  .in1({ S109, DP_AC_q_3 }),
  .out1({ S115 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_348_ (
  .in1({ S110, S1224 }),
  .out1({ S116 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_374_ (
  .in1({ S2440, S1971 }),
  .out1({ S117 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_129_ (
  .in1({ S117 }),
  .out1({ S118 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_349_ (
  .in1({ S2440, S2538[2] }),
  .out1({ S119 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_130_ (
  .in1({ S119 }),
  .out1({ S120 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_350_ (
  .in1({ S119, S118 }),
  .out1({ S121 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_375_ (
  .in1({ S120, S117 }),
  .out1({ S122 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_376_ (
  .in1({ S122, S2433 }),
  .out1({ S123 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_351_ (
  .in1({ S121, S2434 }),
  .out1({ S124 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_352_ (
  .in1({ S121, DP_AC_q_2 }),
  .out1({ S125 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_377_ (
  .in1({ S124, S1213 }),
  .out1({ S126 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_353_ (
  .in1({ S123, DP_AC_q_2 }),
  .out1({ S127 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_378_ (
  .in1({ S123, DP_AC_q_2 }),
  .out1({ S128 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_131_ (
  .in1({ S128 }),
  .out1({ S129 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_379_ (
  .in1({ S128, S126 }),
  .out1({ S130 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_354_ (
  .in1({ S129, S127 }),
  .out1({ S131 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_380_ (
  .in1({ S2440, S1964 }),
  .out1({ S132 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_132_ (
  .in1({ S132 }),
  .out1({ S133 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_355_ (
  .in1({ S2440, S2538[1] }),
  .out1({ S134 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_133_ (
  .in1({ S134 }),
  .out1({ S135 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_356_ (
  .in1({ S134, S133 }),
  .out1({ S136 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_381_ (
  .in1({ S135, S132 }),
  .out1({ S137 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_382_ (
  .in1({ S137, S2433 }),
  .out1({ S138 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_357_ (
  .in1({ S136, S2434 }),
  .out1({ S139 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_383_ (
  .in1({ S137, S1202 }),
  .out1({ S140 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_384_ (
  .in1({ S139, S1202 }),
  .out1({ S141 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_358_ (
  .in1({ S138, DP_AC_q_1 }),
  .out1({ S142 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_385_ (
  .in1({ S138, DP_AC_q_1 }),
  .out1({ S143 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_134_ (
  .in1({ S143 }),
  .out1({ S144 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_386_ (
  .in1({ S143, S141 }),
  .out1({ S145 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_359_ (
  .in1({ S144, S142 }),
  .out1({ S146 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_387_ (
  .in1({ S2440, S1952 }),
  .out1({ S147 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_360_ (
  .in1({ S2439, S1951 }),
  .out1({ S148 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_361_ (
  .in1({ S2440, S2538[0] }),
  .out1({ S149 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_135_ (
  .in1({ S149 }),
  .out1({ S150 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_362_ (
  .in1({ S149, S148 }),
  .out1({ S151 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_388_ (
  .in1({ S150, S147 }),
  .out1({ S152 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_389_ (
  .in1({ S151, S2433 }),
  .out1({ S153 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_363_ (
  .in1({ S152, S2434 }),
  .out1({ S154 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_390_ (
  .in1({ S153, S1191 }),
  .out1({ S155 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_364_ (
  .in1({ S154, DP_AC_q_0 }),
  .out1({ S156 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_391_ (
  .in1({ S156, S146 }),
  .out1({ S157 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_365_ (
  .in1({ S155, S145 }),
  .out1({ S158 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_392_ (
  .in1({ S157, S141 }),
  .out1({ S159 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_366_ (
  .in1({ S158, S142 }),
  .out1({ S160 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_393_ (
  .in1({ S159, S131 }),
  .out1({ S161 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_367_ (
  .in1({ S160, S130 }),
  .out1({ S162 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_394_ (
  .in1({ S161, S126 }),
  .out1({ S163 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_368_ (
  .in1({ S162, S127 }),
  .out1({ S164 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_395_ (
  .in1({ S163, S115 }),
  .out1({ S165 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_369_ (
  .in1({ S164, S116 }),
  .out1({ S166 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_396_ (
  .in1({ S165, S113 }),
  .out1({ S167 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_370_ (
  .in1({ S166, S114 }),
  .out1({ S168 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_397_ (
  .in1({ S167, S102 }),
  .out1({ S169 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_398_ (
  .in1({ S169, S97 }),
  .out1({ S170 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_399_ (
  .in1({ S170, S86 }),
  .out1({ S171 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_400_ (
  .in1({ S171, S84 }),
  .out1({ S172 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_136_ (
  .in1({ S172 }),
  .out1({ S173 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_371_ (
  .in1({ S173, S74 }),
  .out1({ S174 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_372_ (
  .in1({ S174, S2535 }),
  .out1({ S175 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_137_ (
  .in1({ S175 }),
  .out1({ S176 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_401_ (
  .in1({ S176, S2526 }),
  .out1({ S177 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_138_ (
  .in1({ S177 }),
  .out1({ S178 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_402_ (
  .in1({ S177, S2522 }),
  .out1({ S179 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_373_ (
  .in1({ S178, S2523 }),
  .out1({ S180 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_374_ (
  .in1({ S180, S2513 }),
  .out1({ S181 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_375_ (
  .in1({ S181, S2509 }),
  .out1({ S182 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_403_ (
  .in1({ S182, S2502 }),
  .out1({ S183 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_404_ (
  .in1({ S183, S2503 }),
  .out1({ S184 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_376_ (
  .in1({ S184, S2495 }),
  .out1({ S185 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_139_ (
  .in1({ S185 }),
  .out1({ S186 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_405_ (
  .in1({ S185, S2486 }),
  .out1({ S187 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_377_ (
  .in1({ S2493, S2485 }),
  .out1({ S188 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_406_ (
  .in1({ S187, S2483 }),
  .out1({ S189 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_378_ (
  .in1({ S189, S188 }),
  .out1({ S190 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_140_ (
  .in1({ S190 }),
  .out1({ S191 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_407_ (
  .in1({ S191, S2477 }),
  .out1({ S192 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_379_ (
  .in1({ S192, S2468 }),
  .out1({ S193 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_408_ (
  .in1({ S2473, S2467 }),
  .out1({ S194 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_409_ (
  .in1({ S194, S2464 }),
  .out1({ S195 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_380_ (
  .in1({ S195, S193 }),
  .out1({ S196 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_141_ (
  .in1({ S196 }),
  .out1({ S197 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_410_ (
  .in1({ S197, S2458 }),
  .out1({ S198 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_411_ (
  .in1({ S198, S2455 }),
  .out1({ S199 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_381_ (
  .in1({ S199, S2449 }),
  .out1({ S200 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_412_ (
  .in1({ S199, S2449 }),
  .out1({ S201 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_142_ (
  .in1({ S201 }),
  .out1({ S202 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_382_ (
  .in1({ S202, S200 }),
  .out1({ S203 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_383_ (
  .in1({ S203, S2432 }),
  .out1({ S204 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_384_ (
  .in1({ S2519, DP_AC_q_5 }),
  .out1({ S205 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_385_ (
  .in1({ S80, DP_AC_q_7 }),
  .out1({ S206 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_413_ (
  .in1({ S85, S2523 }),
  .out1({ S207 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_386_ (
  .in1({ S84, S2522 }),
  .out1({ S208 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_387_ (
  .in1({ S206, S205 }),
  .out1({ S209 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_143_ (
  .in1({ S209 }),
  .out1({ S210 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_414_ (
  .in1({ S210, S207 }),
  .out1({ S211 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_388_ (
  .in1({ S209, S208 }),
  .out1({ S212 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_415_ (
  .in1({ S212, S2535 }),
  .out1({ S213 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_389_ (
  .in1({ S211, S2534 }),
  .out1({ S214 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_390_ (
  .in1({ S212, S2535 }),
  .out1({ S215 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_391_ (
  .in1({ S215, S214 }),
  .out1({ S216 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_392_ (
  .in1({ S2519, DP_AC_q_4 }),
  .out1({ S217 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_393_ (
  .in1({ S80, DP_AC_q_6 }),
  .out1({ S218 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_394_ (
  .in1({ S2519, DP_AC_q_6 }),
  .out1({ S219 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_144_ (
  .in1({ S219 }),
  .out1({ S220 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_416_ (
  .in1({ S81, S1235 }),
  .out1({ S221 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_395_ (
  .in1({ S80, DP_AC_q_4 }),
  .out1({ S222 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_417_ (
  .in1({ S222, S219 }),
  .out1({ S223 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_396_ (
  .in1({ S221, S220 }),
  .out1({ S224 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_397_ (
  .in1({ S2532, DP_AC_q_5 }),
  .out1({ S225 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_145_ (
  .in1({ S225 }),
  .out1({ S226 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_398_ (
  .in1({ S218, S217 }),
  .out1({ S227 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_399_ (
  .in1({ S227, S224 }),
  .out1({ S228 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_146_ (
  .in1({ S228 }),
  .out1({ S229 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_418_ (
  .in1({ S228, S225 }),
  .out1({ S230 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_400_ (
  .in1({ S229, S226 }),
  .out1({ S231 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_419_ (
  .in1({ S230, S223 }),
  .out1({ S232 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_420_ (
  .in1({ S232, S216 }),
  .out1({ S233 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_147_ (
  .in1({ S233 }),
  .out1({ S234 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_401_ (
  .in1({ S232, S216 }),
  .out1({ S235 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_402_ (
  .in1({ S235, S234 }),
  .out1({ S236 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_421_ (
  .in1({ S2520, S1224 }),
  .out1({ S237 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_403_ (
  .in1({ S2519, DP_AC_q_3 }),
  .out1({ S238 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_422_ (
  .in1({ S238, S82 }),
  .out1({ S239 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_404_ (
  .in1({ S237, S83 }),
  .out1({ S240 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_423_ (
  .in1({ S2533, S1235 }),
  .out1({ S241 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_405_ (
  .in1({ S2532, DP_AC_q_4 }),
  .out1({ S242 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_424_ (
  .in1({ S237, S84 }),
  .out1({ S243 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_406_ (
  .in1({ S238, S85 }),
  .out1({ S244 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_425_ (
  .in1({ S243, S239 }),
  .out1({ S245 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_407_ (
  .in1({ S244, S240 }),
  .out1({ S246 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_426_ (
  .in1({ S246, S242 }),
  .out1({ S247 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_408_ (
  .in1({ S245, S241 }),
  .out1({ S248 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_427_ (
  .in1({ S247, S239 }),
  .out1({ S249 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_409_ (
  .in1({ S248, S240 }),
  .out1({ S250 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_410_ (
  .in1({ S228, S225 }),
  .out1({ S251 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_148_ (
  .in1({ S251 }),
  .out1({ S252 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_428_ (
  .in1({ S252, S230 }),
  .out1({ S253 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_411_ (
  .in1({ S251, S231 }),
  .out1({ S254 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_429_ (
  .in1({ S254, S249 }),
  .out1({ S255 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_412_ (
  .in1({ S253, S250 }),
  .out1({ S256 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_430_ (
  .in1({ S94, S1268 }),
  .out1({ S257 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_413_ (
  .in1({ S93, DP_AC_q_7 }),
  .out1({ S258 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_431_ (
  .in1({ S253, S250 }),
  .out1({ S259 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_414_ (
  .in1({ S254, S249 }),
  .out1({ S260 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_432_ (
  .in1({ S259, S255 }),
  .out1({ S261 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_415_ (
  .in1({ S260, S256 }),
  .out1({ S262 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_433_ (
  .in1({ S262, S258 }),
  .out1({ S263 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_416_ (
  .in1({ S261, S257 }),
  .out1({ S264 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_434_ (
  .in1({ S263, S255 }),
  .out1({ S265 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_435_ (
  .in1({ S265, S236 }),
  .out1({ S266 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_149_ (
  .in1({ S266 }),
  .out1({ S267 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_417_ (
  .in1({ S265, S236 }),
  .out1({ S268 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_418_ (
  .in1({ S268, S267 }),
  .out1({ S269 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_150_ (
  .in1({ S269 }),
  .out1({ S270 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_436_ (
  .in1({ S2520, S1213 }),
  .out1({ S271 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_419_ (
  .in1({ S2519, DP_AC_q_2 }),
  .out1({ S272 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_420_ (
  .in1({ S80, DP_AC_q_2 }),
  .out1({ S273 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_437_ (
  .in1({ S272, S222 }),
  .out1({ S274 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_421_ (
  .in1({ S271, S221 }),
  .out1({ S275 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_438_ (
  .in1({ S2533, S1224 }),
  .out1({ S276 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_422_ (
  .in1({ S2532, DP_AC_q_3 }),
  .out1({ S277 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_423_ (
  .in1({ S272, S222 }),
  .out1({ S278 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_151_ (
  .in1({ S278 }),
  .out1({ S279 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_439_ (
  .in1({ S279, S274 }),
  .out1({ S280 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_424_ (
  .in1({ S278, S275 }),
  .out1({ S281 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_440_ (
  .in1({ S281, S277 }),
  .out1({ S282 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_425_ (
  .in1({ S280, S276 }),
  .out1({ S283 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_441_ (
  .in1({ S282, S274 }),
  .out1({ S284 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_426_ (
  .in1({ S283, S275 }),
  .out1({ S285 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_442_ (
  .in1({ S245, S241 }),
  .out1({ S286 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_427_ (
  .in1({ S246, S242 }),
  .out1({ S287 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_443_ (
  .in1({ S286, S247 }),
  .out1({ S288 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_428_ (
  .in1({ S287, S248 }),
  .out1({ S289 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_444_ (
  .in1({ S289, S284 }),
  .out1({ S290 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_429_ (
  .in1({ S288, S285 }),
  .out1({ S291 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_430_ (
  .in1({ S109, DP_AC_q_7 }),
  .out1({ S292 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_431_ (
  .in1({ S93, DP_AC_q_6 }),
  .out1({ S293 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_152_ (
  .in1({ S293 }),
  .out1({ S294 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_432_ (
  .in1({ S109, DP_AC_q_6 }),
  .out1({ S295 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_153_ (
  .in1({ S295 }),
  .out1({ S296 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_445_ (
  .in1({ S295, S258 }),
  .out1({ S297 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_433_ (
  .in1({ S296, S257 }),
  .out1({ S298 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_434_ (
  .in1({ S293, S292 }),
  .out1({ S299 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_154_ (
  .in1({ S299 }),
  .out1({ S300 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_446_ (
  .in1({ S300, S297 }),
  .out1({ S301 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_435_ (
  .in1({ S299, S298 }),
  .out1({ S302 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_447_ (
  .in1({ S288, S285 }),
  .out1({ S303 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_436_ (
  .in1({ S289, S284 }),
  .out1({ S304 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_448_ (
  .in1({ S303, S290 }),
  .out1({ S305 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_437_ (
  .in1({ S304, S291 }),
  .out1({ S306 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_449_ (
  .in1({ S306, S302 }),
  .out1({ S307 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_438_ (
  .in1({ S305, S301 }),
  .out1({ S308 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_450_ (
  .in1({ S307, S290 }),
  .out1({ S309 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_439_ (
  .in1({ S308, S291 }),
  .out1({ S310 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_451_ (
  .in1({ S261, S257 }),
  .out1({ S311 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_440_ (
  .in1({ S262, S258 }),
  .out1({ S312 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_452_ (
  .in1({ S311, S263 }),
  .out1({ S313 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_441_ (
  .in1({ S312, S264 }),
  .out1({ S314 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_453_ (
  .in1({ S314, S309 }),
  .out1({ S315 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_442_ (
  .in1({ S313, S310 }),
  .out1({ S316 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_454_ (
  .in1({ S313, S310 }),
  .out1({ S317 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_443_ (
  .in1({ S314, S309 }),
  .out1({ S318 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_455_ (
  .in1({ S317, S315 }),
  .out1({ S319 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_444_ (
  .in1({ S318, S316 }),
  .out1({ S320 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_456_ (
  .in1({ S320, S298 }),
  .out1({ S321 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_457_ (
  .in1({ S321, S315 }),
  .out1({ S322 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_155_ (
  .in1({ S322 }),
  .out1({ S323 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_445_ (
  .in1({ S323, S270 }),
  .out1({ S324 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_156_ (
  .in1({ S324 }),
  .out1({ S325 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_458_ (
  .in1({ S213, S207 }),
  .out1({ S326 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_446_ (
  .in1({ S214, S208 }),
  .out1({ S327 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_447_ (
  .in1({ S2532, DP_AC_q_7 }),
  .out1({ S328 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_459_ (
  .in1({ S2535, S2523 }),
  .out1({ S329 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_448_ (
  .in1({ S2534, S2522 }),
  .out1({ S330 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_449_ (
  .in1({ S328, S219 }),
  .out1({ S331 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_157_ (
  .in1({ S331 }),
  .out1({ S332 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_460_ (
  .in1({ S332, S329 }),
  .out1({ S333 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_450_ (
  .in1({ S331, S330 }),
  .out1({ S334 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_451_ (
  .in1({ S333, S327 }),
  .out1({ S335 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_158_ (
  .in1({ S335 }),
  .out1({ S336 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_452_ (
  .in1({ S334, S326 }),
  .out1({ S337 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_159_ (
  .in1({ S337 }),
  .out1({ S338 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_461_ (
  .in1({ S338, S336 }),
  .out1({ S339 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_462_ (
  .in1({ S266, S233 }),
  .out1({ S340 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_453_ (
  .in1({ S340, S339 }),
  .out1({ S341 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_160_ (
  .in1({ S341 }),
  .out1({ S342 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_463_ (
  .in1({ S340, S339 }),
  .out1({ S343 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_161_ (
  .in1({ S343 }),
  .out1({ S344 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_454_ (
  .in1({ S337, S233 }),
  .out1({ S345 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_455_ (
  .in1({ S339, S266 }),
  .out1({ S346 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_456_ (
  .in1({ S344, S341 }),
  .out1({ S347 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_464_ (
  .in1({ S343, S342 }),
  .out1({ S348 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_465_ (
  .in1({ S348, S324 }),
  .out1({ S349 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_466_ (
  .in1({ S347, S325 }),
  .out1({ S350 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_467_ (
  .in1({ S350, S349 }),
  .out1({ S351 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_162_ (
  .in1({ S351 }),
  .out1({ S352 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_457_ (
  .in1({ S322, S269 }),
  .out1({ S353 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_458_ (
  .in1({ S353, S324 }),
  .out1({ S354 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_163_ (
  .in1({ S354 }),
  .out1({ S355 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_459_ (
  .in1({ S2519, DP_AC_q_1 }),
  .out1({ S356 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_460_ (
  .in1({ S80, DP_AC_q_3 }),
  .out1({ S357 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_461_ (
  .in1({ S80, DP_AC_q_1 }),
  .out1({ S358 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_164_ (
  .in1({ S358 }),
  .out1({ S359 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_468_ (
  .in1({ S358, S238 }),
  .out1({ S360 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_462_ (
  .in1({ S359, S237 }),
  .out1({ S361 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_463_ (
  .in1({ S2532, DP_AC_q_2 }),
  .out1({ S362 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_165_ (
  .in1({ S362 }),
  .out1({ S363 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_464_ (
  .in1({ S357, S356 }),
  .out1({ S364 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_465_ (
  .in1({ S364, S361 }),
  .out1({ S365 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_166_ (
  .in1({ S365 }),
  .out1({ S366 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_469_ (
  .in1({ S365, S362 }),
  .out1({ S367 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_466_ (
  .in1({ S366, S363 }),
  .out1({ S368 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_470_ (
  .in1({ S367, S360 }),
  .out1({ S369 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_167_ (
  .in1({ S369 }),
  .out1({ S370 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_467_ (
  .in1({ S281, S277 }),
  .out1({ S371 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_468_ (
  .in1({ S371, S283 }),
  .out1({ S372 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_168_ (
  .in1({ S372 }),
  .out1({ S373 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_471_ (
  .in1({ S372, S369 }),
  .out1({ S374 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_469_ (
  .in1({ S373, S370 }),
  .out1({ S375 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_470_ (
  .in1({ S93, DP_AC_q_5 }),
  .out1({ S376 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_472_ (
  .in1({ S110, S1246 }),
  .out1({ S377 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_471_ (
  .in1({ S109, DP_AC_q_5 }),
  .out1({ S378 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_473_ (
  .in1({ S378, S293 }),
  .out1({ S379 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_472_ (
  .in1({ S377, S294 }),
  .out1({ S380 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_473_ (
  .in1({ S376, S295 }),
  .out1({ S381 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_169_ (
  .in1({ S381 }),
  .out1({ S382 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_474_ (
  .in1({ S382, S379 }),
  .out1({ S383 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_474_ (
  .in1({ S381, S380 }),
  .out1({ S384 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_475_ (
  .in1({ S372, S369 }),
  .out1({ S385 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_170_ (
  .in1({ S385 }),
  .out1({ S386 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_475_ (
  .in1({ S386, S374 }),
  .out1({ S387 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_476_ (
  .in1({ S385, S375 }),
  .out1({ S388 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_476_ (
  .in1({ S388, S384 }),
  .out1({ S389 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_477_ (
  .in1({ S387, S383 }),
  .out1({ S390 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_477_ (
  .in1({ S389, S374 }),
  .out1({ S391 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_478_ (
  .in1({ S390, S375 }),
  .out1({ S392 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_478_ (
  .in1({ S305, S301 }),
  .out1({ S393 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_479_ (
  .in1({ S306, S302 }),
  .out1({ S394 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_479_ (
  .in1({ S393, S307 }),
  .out1({ S395 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_480_ (
  .in1({ S394, S308 }),
  .out1({ S396 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_480_ (
  .in1({ S396, S391 }),
  .out1({ S397 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_481_ (
  .in1({ S395, S392 }),
  .out1({ S398 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_481_ (
  .in1({ S395, S392 }),
  .out1({ S399 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_482_ (
  .in1({ S396, S391 }),
  .out1({ S400 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_482_ (
  .in1({ S399, S397 }),
  .out1({ S401 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_483_ (
  .in1({ S400, S398 }),
  .out1({ S402 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_483_ (
  .in1({ S402, S380 }),
  .out1({ S403 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_484_ (
  .in1({ S401, S379 }),
  .out1({ S404 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_485_ (
  .in1({ S404, S398 }),
  .out1({ S405 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_484_ (
  .in1({ S319, S297 }),
  .out1({ S406 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_485_ (
  .in1({ S406, S321 }),
  .out1({ S407 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_486_ (
  .in1({ S407, S405 }),
  .out1({ S408 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_171_ (
  .in1({ S408 }),
  .out1({ S409 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_487_ (
  .in1({ S409, S355 }),
  .out1({ S410 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_172_ (
  .in1({ S410 }),
  .out1({ S411 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_488_ (
  .in1({ S408, S354 }),
  .out1({ S412 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_489_ (
  .in1({ S412, S410 }),
  .out1({ S413 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_490_ (
  .in1({ S365, S362 }),
  .out1({ S414 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_173_ (
  .in1({ S414 }),
  .out1({ S415 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_486_ (
  .in1({ S415, S367 }),
  .out1({ S416 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_491_ (
  .in1({ S414, S368 }),
  .out1({ S417 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_492_ (
  .in1({ S2519, DP_AC_q_0 }),
  .out1({ S418 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_487_ (
  .in1({ S81, S1191 }),
  .out1({ S419 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_493_ (
  .in1({ S80, DP_AC_q_0 }),
  .out1({ S420 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_494_ (
  .in1({ S419, S271 }),
  .out1({ S421 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_174_ (
  .in1({ S421 }),
  .out1({ S422 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_495_ (
  .in1({ S418, S273 }),
  .out1({ S423 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_175_ (
  .in1({ S423 }),
  .out1({ S424 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_488_ (
  .in1({ S2533, S1202 }),
  .out1({ S425 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_496_ (
  .in1({ S2532, DP_AC_q_1 }),
  .out1({ S426 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_497_ (
  .in1({ S425, S423 }),
  .out1({ S427 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_498_ (
  .in1({ S426, S421 }),
  .out1({ S428 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_499_ (
  .in1({ S428, S423 }),
  .out1({ S429 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_500_ (
  .in1({ S427, S421 }),
  .out1({ S430 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_489_ (
  .in1({ S429, S417 }),
  .out1({ S431 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_501_ (
  .in1({ S430, S416 }),
  .out1({ S432 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_490_ (
  .in1({ S139, S1268 }),
  .out1({ S433 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_502_ (
  .in1({ S138, DP_AC_q_7 }),
  .out1({ S434 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_491_ (
  .in1({ S378, S96 }),
  .out1({ S435 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_176_ (
  .in1({ S435 }),
  .out1({ S436 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_492_ (
  .in1({ S377, S97 }),
  .out1({ S437 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_503_ (
  .in1({ S378, S98 }),
  .out1({ S438 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_493_ (
  .in1({ S437, S435 }),
  .out1({ S439 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_504_ (
  .in1({ S438, S436 }),
  .out1({ S440 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_494_ (
  .in1({ S439, S433 }),
  .out1({ S441 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_505_ (
  .in1({ S440, S434 }),
  .out1({ S442 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_495_ (
  .in1({ S440, S434 }),
  .out1({ S443 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_177_ (
  .in1({ S443 }),
  .out1({ S444 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_496_ (
  .in1({ S443, S441 }),
  .out1({ S445 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_506_ (
  .in1({ S444, S442 }),
  .out1({ S446 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_497_ (
  .in1({ S430, S416 }),
  .out1({ S447 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_507_ (
  .in1({ S429, S417 }),
  .out1({ S448 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_498_ (
  .in1({ S447, S431 }),
  .out1({ S449 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_508_ (
  .in1({ S448, S432 }),
  .out1({ S450 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_499_ (
  .in1({ S450, S446 }),
  .out1({ S451 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_509_ (
  .in1({ S449, S445 }),
  .out1({ S452 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_500_ (
  .in1({ S451, S431 }),
  .out1({ S453 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_510_ (
  .in1({ S452, S432 }),
  .out1({ S454 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_501_ (
  .in1({ S387, S383 }),
  .out1({ S455 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_511_ (
  .in1({ S388, S384 }),
  .out1({ S456 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_502_ (
  .in1({ S455, S389 }),
  .out1({ S457 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_512_ (
  .in1({ S456, S390 }),
  .out1({ S458 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_503_ (
  .in1({ S458, S453 }),
  .out1({ S459 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_513_ (
  .in1({ S457, S454 }),
  .out1({ S460 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_514_ (
  .in1({ S123, DP_AC_q_7 }),
  .out1({ S461 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_504_ (
  .in1({ S443, S435 }),
  .out1({ S462 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_505_ (
  .in1({ S462, S461 }),
  .out1({ S463 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_178_ (
  .in1({ S463 }),
  .out1({ S464 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_515_ (
  .in1({ S462, S461 }),
  .out1({ S465 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_179_ (
  .in1({ S465 }),
  .out1({ S466 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_506_ (
  .in1({ S466, S463 }),
  .out1({ S467 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_516_ (
  .in1({ S465, S464 }),
  .out1({ S468 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_507_ (
  .in1({ S457, S454 }),
  .out1({ S469 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_517_ (
  .in1({ S458, S453 }),
  .out1({ S470 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_508_ (
  .in1({ S469, S459 }),
  .out1({ S471 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_518_ (
  .in1({ S470, S460 }),
  .out1({ S472 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_509_ (
  .in1({ S472, S468 }),
  .out1({ S473 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_519_ (
  .in1({ S471, S467 }),
  .out1({ S474 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_510_ (
  .in1({ S473, S459 }),
  .out1({ S475 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_520_ (
  .in1({ S474, S460 }),
  .out1({ S476 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_511_ (
  .in1({ S401, S379 }),
  .out1({ S477 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_521_ (
  .in1({ S402, S380 }),
  .out1({ S478 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_512_ (
  .in1({ S477, S403 }),
  .out1({ S479 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_522_ (
  .in1({ S478, S404 }),
  .out1({ S480 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_513_ (
  .in1({ S480, S475 }),
  .out1({ S481 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_523_ (
  .in1({ S479, S476 }),
  .out1({ S482 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_514_ (
  .in1({ S479, S476 }),
  .out1({ S483 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_515_ (
  .in1({ S483, S481 }),
  .out1({ S484 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_180_ (
  .in1({ S484 }),
  .out1({ S485 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_516_ (
  .in1({ S485, S464 }),
  .out1({ S486 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_181_ (
  .in1({ S486 }),
  .out1({ S487 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_517_ (
  .in1({ S486, S481 }),
  .out1({ S488 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_524_ (
  .in1({ S487, S482 }),
  .out1({ S489 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_518_ (
  .in1({ S407, S405 }),
  .out1({ S490 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_182_ (
  .in1({ S490 }),
  .out1({ S491 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_519_ (
  .in1({ S490, S409 }),
  .out1({ S492 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_525_ (
  .in1({ S491, S408 }),
  .out1({ S493 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_520_ (
  .in1({ S493, S488 }),
  .out1({ S494 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_521_ (
  .in1({ S492, S489 }),
  .out1({ S495 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_522_ (
  .in1({ S495, S494 }),
  .out1({ S496 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_183_ (
  .in1({ S496 }),
  .out1({ S497 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_523_ (
  .in1({ S424, S422 }),
  .out1({ S498 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_526_ (
  .in1({ S423, S421 }),
  .out1({ S499 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_527_ (
  .in1({ S2532, DP_AC_q_0 }),
  .out1({ S500 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_524_ (
  .in1({ S426, S420 }),
  .out1({ S501 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_528_ (
  .in1({ S425, S419 }),
  .out1({ S502 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_529_ (
  .in1({ S501, S499 }),
  .out1({ S503 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_184_ (
  .in1({ S503 }),
  .out1({ S504 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_530_ (
  .in1({ S138, DP_AC_q_6 }),
  .out1({ S505 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_531_ (
  .in1({ S109, DP_AC_q_4 }),
  .out1({ S506 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_532_ (
  .in1({ S93, DP_AC_q_3 }),
  .out1({ S507 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_525_ (
  .in1({ S114, S98 }),
  .out1({ S508 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_533_ (
  .in1({ S113, S97 }),
  .out1({ S509 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_534_ (
  .in1({ S507, S506 }),
  .out1({ S510 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_535_ (
  .in1({ S510, S509 }),
  .out1({ S511 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_536_ (
  .in1({ S511, S505 }),
  .out1({ S512 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_185_ (
  .in1({ S512 }),
  .out1({ S513 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_526_ (
  .in1({ S511, S505 }),
  .out1({ S514 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_186_ (
  .in1({ S514 }),
  .out1({ S515 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_527_ (
  .in1({ S514, S513 }),
  .out1({ S516 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_537_ (
  .in1({ S515, S512 }),
  .out1({ S517 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_528_ (
  .in1({ S426, S419 }),
  .out1({ S518 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_538_ (
  .in1({ S425, S420 }),
  .out1({ S519 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_529_ (
  .in1({ S518, S499 }),
  .out1({ S520 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_539_ (
  .in1({ S519, S498 }),
  .out1({ S521 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_530_ (
  .in1({ S519, S498 }),
  .out1({ S522 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_540_ (
  .in1({ S518, S499 }),
  .out1({ S523 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_531_ (
  .in1({ S522, S520 }),
  .out1({ S524 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_541_ (
  .in1({ S523, S521 }),
  .out1({ S525 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_532_ (
  .in1({ S524, S517 }),
  .out1({ S526 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_542_ (
  .in1({ S525, S516 }),
  .out1({ S527 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_533_ (
  .in1({ S526, S504 }),
  .out1({ S528 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_543_ (
  .in1({ S527, S503 }),
  .out1({ S529 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_534_ (
  .in1({ S449, S445 }),
  .out1({ S530 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_544_ (
  .in1({ S450, S446 }),
  .out1({ S531 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_535_ (
  .in1({ S530, S451 }),
  .out1({ S532 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_545_ (
  .in1({ S531, S452 }),
  .out1({ S533 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_536_ (
  .in1({ S533, S528 }),
  .out1({ S534 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_546_ (
  .in1({ S532, S529 }),
  .out1({ S535 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_547_ (
  .in1({ S123, DP_AC_q_6 }),
  .out1({ S536 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_187_ (
  .in1({ S536 }),
  .out1({ S537 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_537_ (
  .in1({ S514, S508 }),
  .out1({ S538 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_188_ (
  .in1({ S538 }),
  .out1({ S539 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_538_ (
  .in1({ S538, S536 }),
  .out1({ S540 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_548_ (
  .in1({ S539, S537 }),
  .out1({ S541 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_549_ (
  .in1({ S538, S536 }),
  .out1({ S542 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_189_ (
  .in1({ S542 }),
  .out1({ S543 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_539_ (
  .in1({ S543, S540 }),
  .out1({ S544 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_550_ (
  .in1({ S542, S541 }),
  .out1({ S545 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_540_ (
  .in1({ S532, S529 }),
  .out1({ S546 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_551_ (
  .in1({ S533, S528 }),
  .out1({ S547 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_541_ (
  .in1({ S546, S534 }),
  .out1({ S548 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_552_ (
  .in1({ S547, S535 }),
  .out1({ S549 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_542_ (
  .in1({ S549, S545 }),
  .out1({ S550 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_553_ (
  .in1({ S548, S544 }),
  .out1({ S551 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_543_ (
  .in1({ S550, S534 }),
  .out1({ S552 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_554_ (
  .in1({ S551, S535 }),
  .out1({ S553 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_544_ (
  .in1({ S471, S467 }),
  .out1({ S554 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_555_ (
  .in1({ S472, S468 }),
  .out1({ S555 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_545_ (
  .in1({ S554, S473 }),
  .out1({ S556 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_556_ (
  .in1({ S555, S474 }),
  .out1({ S557 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_557_ (
  .in1({ S556, S553 }),
  .out1({ S558 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_190_ (
  .in1({ S558 }),
  .out1({ S559 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_546_ (
  .in1({ S556, S553 }),
  .out1({ S560 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_558_ (
  .in1({ S557, S552 }),
  .out1({ S561 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_547_ (
  .in1({ S560, S559 }),
  .out1({ S562 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_559_ (
  .in1({ S561, S558 }),
  .out1({ S563 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_560_ (
  .in1({ S562, S540 }),
  .out1({ S564 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_561_ (
  .in1({ S564, S558 }),
  .out1({ S565 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_191_ (
  .in1({ S565 }),
  .out1({ S566 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_548_ (
  .in1({ S484, S463 }),
  .out1({ S567 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_549_ (
  .in1({ S567, S486 }),
  .out1({ S568 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_192_ (
  .in1({ S568 }),
  .out1({ S569 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_550_ (
  .in1({ S569, S566 }),
  .out1({ S570 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_193_ (
  .in1({ S570 }),
  .out1({ S571 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_551_ (
  .in1({ S568, S565 }),
  .out1({ S572 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_552_ (
  .in1({ S572, S570 }),
  .out1({ S573 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_194_ (
  .in1({ S573 }),
  .out1({ S574 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_553_ (
  .in1({ S139, S1246 }),
  .out1({ S575 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_562_ (
  .in1({ S138, DP_AC_q_5 }),
  .out1({ S576 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_554_ (
  .in1({ S94, S1213 }),
  .out1({ S577 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_563_ (
  .in1({ S93, DP_AC_q_2 }),
  .out1({ S578 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_555_ (
  .in1({ S578, S112 }),
  .out1({ S579 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_195_ (
  .in1({ S579 }),
  .out1({ S580 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_556_ (
  .in1({ S577, S113 }),
  .out1({ S581 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_564_ (
  .in1({ S578, S114 }),
  .out1({ S582 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_557_ (
  .in1({ S581, S579 }),
  .out1({ S583 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_565_ (
  .in1({ S582, S580 }),
  .out1({ S584 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_558_ (
  .in1({ S583, S575 }),
  .out1({ S585 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_566_ (
  .in1({ S584, S576 }),
  .out1({ S586 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_559_ (
  .in1({ S584, S576 }),
  .out1({ S587 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_196_ (
  .in1({ S587 }),
  .out1({ S588 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_560_ (
  .in1({ S587, S585 }),
  .out1({ S589 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_567_ (
  .in1({ S588, S586 }),
  .out1({ S590 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_568_ (
  .in1({ S500, S358 }),
  .out1({ S591 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_197_ (
  .in1({ S591 }),
  .out1({ S592 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_561_ (
  .in1({ S592, S501 }),
  .out1({ S593 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_569_ (
  .in1({ S591, S502 }),
  .out1({ S594 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_562_ (
  .in1({ S594, S590 }),
  .out1({ S595 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_570_ (
  .in1({ S593, S589 }),
  .out1({ S596 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_563_ (
  .in1({ S525, S516 }),
  .out1({ S597 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_571_ (
  .in1({ S524, S517 }),
  .out1({ S598 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_564_ (
  .in1({ S597, S526 }),
  .out1({ S599 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_572_ (
  .in1({ S598, S527 }),
  .out1({ S600 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_565_ (
  .in1({ S600, S596 }),
  .out1({ S601 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_573_ (
  .in1({ S599, S595 }),
  .out1({ S602 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_566_ (
  .in1({ S153, S1268 }),
  .out1({ S603 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_574_ (
  .in1({ S154, DP_AC_q_7 }),
  .out1({ S604 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_575_ (
  .in1({ S123, DP_AC_q_5 }),
  .out1({ S605 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_198_ (
  .in1({ S605 }),
  .out1({ S606 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_567_ (
  .in1({ S587, S579 }),
  .out1({ S607 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_199_ (
  .in1({ S607 }),
  .out1({ S608 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_568_ (
  .in1({ S607, S605 }),
  .out1({ S609 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_576_ (
  .in1({ S608, S606 }),
  .out1({ S610 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_577_ (
  .in1({ S607, S605 }),
  .out1({ S611 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_200_ (
  .in1({ S611 }),
  .out1({ S612 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_569_ (
  .in1({ S612, S609 }),
  .out1({ S613 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_578_ (
  .in1({ S611, S610 }),
  .out1({ S614 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_570_ (
  .in1({ S613, S603 }),
  .out1({ S615 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_579_ (
  .in1({ S614, S604 }),
  .out1({ S616 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_571_ (
  .in1({ S614, S604 }),
  .out1({ S617 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_580_ (
  .in1({ S613, S603 }),
  .out1({ S618 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_572_ (
  .in1({ S617, S615 }),
  .out1({ S619 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_581_ (
  .in1({ S618, S616 }),
  .out1({ S620 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_573_ (
  .in1({ S599, S595 }),
  .out1({ S621 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_582_ (
  .in1({ S600, S596 }),
  .out1({ S622 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_574_ (
  .in1({ S621, S601 }),
  .out1({ S623 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_583_ (
  .in1({ S622, S602 }),
  .out1({ S624 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_575_ (
  .in1({ S624, S620 }),
  .out1({ S625 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_584_ (
  .in1({ S623, S619 }),
  .out1({ S626 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_576_ (
  .in1({ S625, S601 }),
  .out1({ S627 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_585_ (
  .in1({ S626, S602 }),
  .out1({ S628 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_577_ (
  .in1({ S548, S544 }),
  .out1({ S629 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_586_ (
  .in1({ S549, S545 }),
  .out1({ S630 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_578_ (
  .in1({ S629, S550 }),
  .out1({ S631 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_587_ (
  .in1({ S630, S551 }),
  .out1({ S632 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_579_ (
  .in1({ S632, S627 }),
  .out1({ S633 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_588_ (
  .in1({ S631, S628 }),
  .out1({ S634 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_580_ (
  .in1({ S617, S609 }),
  .out1({ S635 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_589_ (
  .in1({ S618, S610 }),
  .out1({ S636 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_581_ (
  .in1({ S631, S628 }),
  .out1({ S637 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_590_ (
  .in1({ S632, S627 }),
  .out1({ S638 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_582_ (
  .in1({ S637, S633 }),
  .out1({ S639 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_591_ (
  .in1({ S638, S634 }),
  .out1({ S640 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_583_ (
  .in1({ S640, S635 }),
  .out1({ S641 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_592_ (
  .in1({ S639, S636 }),
  .out1({ S642 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_584_ (
  .in1({ S641, S633 }),
  .out1({ S643 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_201_ (
  .in1({ S643 }),
  .out1({ S644 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_593_ (
  .in1({ S563, S541 }),
  .out1({ S645 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_594_ (
  .in1({ S645, S564 }),
  .out1({ S646 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_202_ (
  .in1({ S646 }),
  .out1({ S647 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_595_ (
  .in1({ S647, S644 }),
  .out1({ S648 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_203_ (
  .in1({ S648 }),
  .out1({ S649 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_585_ (
  .in1({ S139, S1235 }),
  .out1({ S650 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_596_ (
  .in1({ S138, DP_AC_q_4 }),
  .out1({ S651 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_586_ (
  .in1({ S110, S1213 }),
  .out1({ S652 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_597_ (
  .in1({ S109, DP_AC_q_2 }),
  .out1({ S653 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_587_ (
  .in1({ S94, S1202 }),
  .out1({ S654 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_598_ (
  .in1({ S93, DP_AC_q_1 }),
  .out1({ S655 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_588_ (
  .in1({ S110, S1202 }),
  .out1({ S656 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_599_ (
  .in1({ S109, DP_AC_q_1 }),
  .out1({ S657 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_589_ (
  .in1({ S655, S653 }),
  .out1({ S658 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_204_ (
  .in1({ S658 }),
  .out1({ S659 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_590_ (
  .in1({ S654, S652 }),
  .out1({ S660 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_600_ (
  .in1({ S655, S653 }),
  .out1({ S661 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_591_ (
  .in1({ S660, S658 }),
  .out1({ S662 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_601_ (
  .in1({ S661, S659 }),
  .out1({ S663 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_592_ (
  .in1({ S662, S650 }),
  .out1({ S664 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_602_ (
  .in1({ S663, S651 }),
  .out1({ S665 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_593_ (
  .in1({ S663, S651 }),
  .out1({ S666 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_205_ (
  .in1({ S666 }),
  .out1({ S667 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_594_ (
  .in1({ S666, S664 }),
  .out1({ S668 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_603_ (
  .in1({ S667, S665 }),
  .out1({ S669 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_595_ (
  .in1({ S669, S420 }),
  .out1({ S670 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_604_ (
  .in1({ S668, S419 }),
  .out1({ S671 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_596_ (
  .in1({ S593, S589 }),
  .out1({ S672 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_605_ (
  .in1({ S594, S590 }),
  .out1({ S673 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_597_ (
  .in1({ S672, S595 }),
  .out1({ S674 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_606_ (
  .in1({ S673, S596 }),
  .out1({ S675 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_598_ (
  .in1({ S675, S671 }),
  .out1({ S676 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_607_ (
  .in1({ S674, S670 }),
  .out1({ S677 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_599_ (
  .in1({ S153, S1257 }),
  .out1({ S678 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_608_ (
  .in1({ S154, DP_AC_q_6 }),
  .out1({ S679 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_609_ (
  .in1({ S123, DP_AC_q_4 }),
  .out1({ S680 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_206_ (
  .in1({ S680 }),
  .out1({ S681 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_600_ (
  .in1({ S666, S658 }),
  .out1({ S682 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_207_ (
  .in1({ S682 }),
  .out1({ S683 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_601_ (
  .in1({ S682, S680 }),
  .out1({ S684 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_610_ (
  .in1({ S683, S681 }),
  .out1({ S685 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_611_ (
  .in1({ S682, S680 }),
  .out1({ S686 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_208_ (
  .in1({ S686 }),
  .out1({ S687 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_602_ (
  .in1({ S687, S684 }),
  .out1({ S688 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_612_ (
  .in1({ S686, S685 }),
  .out1({ S689 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_603_ (
  .in1({ S688, S678 }),
  .out1({ S690 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_613_ (
  .in1({ S689, S679 }),
  .out1({ S691 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_604_ (
  .in1({ S689, S679 }),
  .out1({ S692 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_614_ (
  .in1({ S688, S678 }),
  .out1({ S693 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_605_ (
  .in1({ S692, S690 }),
  .out1({ S694 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_615_ (
  .in1({ S693, S691 }),
  .out1({ S695 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_606_ (
  .in1({ S674, S670 }),
  .out1({ S696 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_616_ (
  .in1({ S675, S671 }),
  .out1({ S697 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_607_ (
  .in1({ S696, S676 }),
  .out1({ S698 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_617_ (
  .in1({ S697, S677 }),
  .out1({ S699 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_608_ (
  .in1({ S699, S695 }),
  .out1({ S700 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_618_ (
  .in1({ S698, S694 }),
  .out1({ S701 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_609_ (
  .in1({ S700, S676 }),
  .out1({ S702 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_619_ (
  .in1({ S701, S677 }),
  .out1({ S703 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_610_ (
  .in1({ S623, S619 }),
  .out1({ S704 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_620_ (
  .in1({ S624, S620 }),
  .out1({ S705 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_611_ (
  .in1({ S704, S625 }),
  .out1({ S706 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_621_ (
  .in1({ S705, S626 }),
  .out1({ S707 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_612_ (
  .in1({ S707, S702 }),
  .out1({ S708 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_622_ (
  .in1({ S706, S703 }),
  .out1({ S709 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_613_ (
  .in1({ S692, S684 }),
  .out1({ S710 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_623_ (
  .in1({ S693, S685 }),
  .out1({ S711 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_614_ (
  .in1({ S706, S703 }),
  .out1({ S712 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_624_ (
  .in1({ S707, S702 }),
  .out1({ S713 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_615_ (
  .in1({ S712, S708 }),
  .out1({ S714 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_625_ (
  .in1({ S713, S709 }),
  .out1({ S715 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_616_ (
  .in1({ S715, S710 }),
  .out1({ S716 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_626_ (
  .in1({ S714, S711 }),
  .out1({ S717 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_617_ (
  .in1({ S716, S708 }),
  .out1({ S718 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_627_ (
  .in1({ S640, S635 }),
  .out1({ S719 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_628_ (
  .in1({ S719, S642 }),
  .out1({ S720 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_618_ (
  .in1({ S720, S718 }),
  .out1({ S721 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_209_ (
  .in1({ S721 }),
  .out1({ S722 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_629_ (
  .in1({ S720, S718 }),
  .out1({ S723 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_210_ (
  .in1({ S723 }),
  .out1({ S724 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_619_ (
  .in1({ S724, S721 }),
  .out1({ S725 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_630_ (
  .in1({ S723, S722 }),
  .out1({ S726 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_620_ (
  .in1({ S153, S1246 }),
  .out1({ S727 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_631_ (
  .in1({ S154, DP_AC_q_5 }),
  .out1({ S728 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_621_ (
  .in1({ S124, S1224 }),
  .out1({ S729 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_632_ (
  .in1({ S123, DP_AC_q_3 }),
  .out1({ S730 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_622_ (
  .in1({ S94, S1191 }),
  .out1({ S731 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_633_ (
  .in1({ S93, DP_AC_q_0 }),
  .out1({ S732 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_634_ (
  .in1({ S109, DP_AC_q_0 }),
  .out1({ S733 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_623_ (
  .in1({ S733, S655 }),
  .out1({ S734 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_635_ (
  .in1({ S731, S656 }),
  .out1({ S735 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_636_ (
  .in1({ S138, DP_AC_q_3 }),
  .out1({ S736 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_211_ (
  .in1({ S736 }),
  .out1({ S737 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_624_ (
  .in1({ S731, S656 }),
  .out1({ S738 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_637_ (
  .in1({ S732, S657 }),
  .out1({ S739 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_625_ (
  .in1({ S738, S734 }),
  .out1({ S740 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_638_ (
  .in1({ S739, S735 }),
  .out1({ S741 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_626_ (
  .in1({ S741, S736 }),
  .out1({ S742 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_639_ (
  .in1({ S740, S737 }),
  .out1({ S743 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_627_ (
  .in1({ S742, S734 }),
  .out1({ S744 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_640_ (
  .in1({ S743, S735 }),
  .out1({ S745 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_628_ (
  .in1({ S744, S730 }),
  .out1({ S746 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_641_ (
  .in1({ S745, S729 }),
  .out1({ S747 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_629_ (
  .in1({ S745, S729 }),
  .out1({ S748 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_642_ (
  .in1({ S744, S730 }),
  .out1({ S749 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_630_ (
  .in1({ S748, S746 }),
  .out1({ S750 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_643_ (
  .in1({ S749, S747 }),
  .out1({ S751 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_631_ (
  .in1({ S750, S727 }),
  .out1({ S752 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_644_ (
  .in1({ S751, S728 }),
  .out1({ S753 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_632_ (
  .in1({ S751, S728 }),
  .out1({ S754 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_645_ (
  .in1({ S750, S727 }),
  .out1({ S755 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_633_ (
  .in1({ S754, S752 }),
  .out1({ S756 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_646_ (
  .in1({ S755, S753 }),
  .out1({ S757 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_634_ (
  .in1({ S668, S419 }),
  .out1({ S758 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_647_ (
  .in1({ S669, S420 }),
  .out1({ S759 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_635_ (
  .in1({ S758, S670 }),
  .out1({ S760 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_648_ (
  .in1({ S759, S671 }),
  .out1({ S761 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_636_ (
  .in1({ S761, S757 }),
  .out1({ S762 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_649_ (
  .in1({ S760, S756 }),
  .out1({ S763 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_637_ (
  .in1({ S698, S694 }),
  .out1({ S764 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_650_ (
  .in1({ S699, S695 }),
  .out1({ S765 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_638_ (
  .in1({ S764, S700 }),
  .out1({ S766 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_651_ (
  .in1({ S765, S701 }),
  .out1({ S767 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_639_ (
  .in1({ S767, S763 }),
  .out1({ S768 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_652_ (
  .in1({ S766, S762 }),
  .out1({ S769 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_640_ (
  .in1({ S754, S746 }),
  .out1({ S770 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_212_ (
  .in1({ S770 }),
  .out1({ S771 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_641_ (
  .in1({ S766, S762 }),
  .out1({ S772 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_653_ (
  .in1({ S767, S763 }),
  .out1({ S773 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_642_ (
  .in1({ S772, S768 }),
  .out1({ S774 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_654_ (
  .in1({ S773, S769 }),
  .out1({ S775 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_643_ (
  .in1({ S775, S770 }),
  .out1({ S776 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_655_ (
  .in1({ S774, S771 }),
  .out1({ S777 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_644_ (
  .in1({ S776, S768 }),
  .out1({ S778 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_656_ (
  .in1({ S777, S769 }),
  .out1({ S779 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_645_ (
  .in1({ S714, S711 }),
  .out1({ S780 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_657_ (
  .in1({ S715, S710 }),
  .out1({ S781 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_646_ (
  .in1({ S780, S716 }),
  .out1({ S782 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_658_ (
  .in1({ S781, S717 }),
  .out1({ S783 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_647_ (
  .in1({ S783, S778 }),
  .out1({ S784 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_659_ (
  .in1({ S782, S779 }),
  .out1({ S785 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_648_ (
  .in1({ S782, S779 }),
  .out1({ S786 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_649_ (
  .in1({ S786, S784 }),
  .out1({ S787 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_213_ (
  .in1({ S787 }),
  .out1({ S788 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_650_ (
  .in1({ S153, S1235 }),
  .out1({ S789 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_660_ (
  .in1({ S154, DP_AC_q_4 }),
  .out1({ S790 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_661_ (
  .in1({ S138, DP_AC_q_2 }),
  .out1({ S791 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_662_ (
  .in1({ S138, DP_AC_q_0 }),
  .out1({ S792 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_214_ (
  .in1({ S792 }),
  .out1({ S793 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_651_ (
  .in1({ S792, S653 }),
  .out1({ S794 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_663_ (
  .in1({ S793, S652 }),
  .out1({ S795 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_652_ (
  .in1({ S795, S124 }),
  .out1({ S796 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_664_ (
  .in1({ S794, S123 }),
  .out1({ S797 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_653_ (
  .in1({ S794, S126 }),
  .out1({ S798 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_665_ (
  .in1({ S795, S127 }),
  .out1({ S799 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_654_ (
  .in1({ S798, S796 }),
  .out1({ S800 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_666_ (
  .in1({ S799, S797 }),
  .out1({ S801 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_655_ (
  .in1({ S800, S789 }),
  .out1({ S802 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_667_ (
  .in1({ S801, S790 }),
  .out1({ S803 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_656_ (
  .in1({ S801, S790 }),
  .out1({ S804 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_668_ (
  .in1({ S800, S789 }),
  .out1({ S805 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_657_ (
  .in1({ S804, S802 }),
  .out1({ S806 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_669_ (
  .in1({ S805, S803 }),
  .out1({ S807 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_670_ (
  .in1({ S741, S736 }),
  .out1({ S808 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_215_ (
  .in1({ S808 }),
  .out1({ S809 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_658_ (
  .in1({ S809, S742 }),
  .out1({ S810 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_216_ (
  .in1({ S810 }),
  .out1({ S811 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_659_ (
  .in1({ S811, S807 }),
  .out1({ S812 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_671_ (
  .in1({ S810, S806 }),
  .out1({ S813 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_660_ (
  .in1({ S760, S756 }),
  .out1({ S814 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_672_ (
  .in1({ S761, S757 }),
  .out1({ S815 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_661_ (
  .in1({ S814, S762 }),
  .out1({ S816 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_673_ (
  .in1({ S815, S763 }),
  .out1({ S817 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_662_ (
  .in1({ S817, S813 }),
  .out1({ S818 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_674_ (
  .in1({ S816, S812 }),
  .out1({ S819 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_663_ (
  .in1({ S804, S796 }),
  .out1({ S820 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_675_ (
  .in1({ S805, S797 }),
  .out1({ S821 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_664_ (
  .in1({ S816, S812 }),
  .out1({ S822 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_676_ (
  .in1({ S817, S813 }),
  .out1({ S823 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_665_ (
  .in1({ S822, S818 }),
  .out1({ S824 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_677_ (
  .in1({ S823, S819 }),
  .out1({ S825 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_666_ (
  .in1({ S825, S820 }),
  .out1({ S826 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_678_ (
  .in1({ S824, S821 }),
  .out1({ S827 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_667_ (
  .in1({ S826, S818 }),
  .out1({ S828 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_679_ (
  .in1({ S827, S819 }),
  .out1({ S829 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_668_ (
  .in1({ S774, S771 }),
  .out1({ S830 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_680_ (
  .in1({ S775, S770 }),
  .out1({ S831 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_669_ (
  .in1({ S830, S776 }),
  .out1({ S832 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_681_ (
  .in1({ S831, S777 }),
  .out1({ S833 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_670_ (
  .in1({ S833, S828 }),
  .out1({ S834 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_682_ (
  .in1({ S832, S829 }),
  .out1({ S835 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_671_ (
  .in1({ S832, S829 }),
  .out1({ S836 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_683_ (
  .in1({ S833, S828 }),
  .out1({ S837 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_672_ (
  .in1({ S836, S834 }),
  .out1({ S838 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_684_ (
  .in1({ S837, S835 }),
  .out1({ S839 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_685_ (
  .in1({ S154, DP_AC_q_3 }),
  .out1({ S840 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_686_ (
  .in1({ S123, DP_AC_q_1 }),
  .out1({ S841 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_687_ (
  .in1({ S154, DP_AC_q_1 }),
  .out1({ S842 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_217_ (
  .in1({ S842 }),
  .out1({ S843 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_673_ (
  .in1({ S842, S730 }),
  .out1({ S844 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_688_ (
  .in1({ S843, S729 }),
  .out1({ S845 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_689_ (
  .in1({ S841, S840 }),
  .out1({ S846 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_218_ (
  .in1({ S846 }),
  .out1({ S847 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_674_ (
  .in1({ S847, S844 }),
  .out1({ S848 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_690_ (
  .in1({ S846, S845 }),
  .out1({ S849 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_691_ (
  .in1({ S791, S733 }),
  .out1({ S850 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_219_ (
  .in1({ S850 }),
  .out1({ S851 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_675_ (
  .in1({ S851, S794 }),
  .out1({ S852 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_692_ (
  .in1({ S850, S795 }),
  .out1({ S853 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_676_ (
  .in1({ S853, S849 }),
  .out1({ S854 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_693_ (
  .in1({ S852, S848 }),
  .out1({ S855 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_677_ (
  .in1({ S810, S806 }),
  .out1({ S856 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_694_ (
  .in1({ S811, S807 }),
  .out1({ S857 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_678_ (
  .in1({ S856, S812 }),
  .out1({ S858 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_695_ (
  .in1({ S857, S813 }),
  .out1({ S859 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_679_ (
  .in1({ S859, S855 }),
  .out1({ S860 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_696_ (
  .in1({ S858, S854 }),
  .out1({ S861 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_680_ (
  .in1({ S858, S854 }),
  .out1({ S862 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_697_ (
  .in1({ S859, S855 }),
  .out1({ S863 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_681_ (
  .in1({ S862, S860 }),
  .out1({ S864 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_698_ (
  .in1({ S863, S861 }),
  .out1({ S865 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_682_ (
  .in1({ S865, S845 }),
  .out1({ S866 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_699_ (
  .in1({ S864, S844 }),
  .out1({ S867 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_683_ (
  .in1({ S866, S860 }),
  .out1({ S868 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_220_ (
  .in1({ S868 }),
  .out1({ S869 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_684_ (
  .in1({ S824, S821 }),
  .out1({ S870 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_700_ (
  .in1({ S825, S820 }),
  .out1({ S871 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_685_ (
  .in1({ S870, S826 }),
  .out1({ S872 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_701_ (
  .in1({ S871, S827 }),
  .out1({ S873 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_702_ (
  .in1({ S872, S869 }),
  .out1({ S874 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_221_ (
  .in1({ S874 }),
  .out1({ S875 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_703_ (
  .in1({ S123, DP_AC_q_0 }),
  .out1({ S876 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_704_ (
  .in1({ S151, DP_AC_q_2 }),
  .out1({ S877 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_705_ (
  .in1({ S151, DP_AC_q_0 }),
  .out1({ S878 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_686_ (
  .in1({ S156, S127 }),
  .out1({ S879 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_706_ (
  .in1({ S155, S126 }),
  .out1({ S880 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_707_ (
  .in1({ S154, DP_AC_q_2 }),
  .out1({ S881 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_708_ (
  .in1({ S881, S876 }),
  .out1({ S882 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_709_ (
  .in1({ S882, S880 }),
  .out1({ S883 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_222_ (
  .in1({ S883 }),
  .out1({ S884 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_687_ (
  .in1({ S883, S142 }),
  .out1({ S885 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_223_ (
  .in1({ S885 }),
  .out1({ S886 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_688_ (
  .in1({ S852, S848 }),
  .out1({ S887 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_710_ (
  .in1({ S853, S849 }),
  .out1({ S888 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_689_ (
  .in1({ S887, S854 }),
  .out1({ S889 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_711_ (
  .in1({ S888, S855 }),
  .out1({ S890 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_690_ (
  .in1({ S890, S886 }),
  .out1({ S891 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_712_ (
  .in1({ S889, S885 }),
  .out1({ S892 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_691_ (
  .in1({ S889, S885 }),
  .out1({ S893 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_713_ (
  .in1({ S890, S886 }),
  .out1({ S894 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_692_ (
  .in1({ S893, S891 }),
  .out1({ S895 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_714_ (
  .in1({ S894, S892 }),
  .out1({ S896 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_693_ (
  .in1({ S896, S880 }),
  .out1({ S897 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_715_ (
  .in1({ S895, S879 }),
  .out1({ S898 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_694_ (
  .in1({ S897, S891 }),
  .out1({ S899 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_716_ (
  .in1({ S898, S892 }),
  .out1({ S900 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_695_ (
  .in1({ S864, S844 }),
  .out1({ S901 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_717_ (
  .in1({ S865, S845 }),
  .out1({ S902 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_696_ (
  .in1({ S901, S866 }),
  .out1({ S903 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_718_ (
  .in1({ S902, S867 }),
  .out1({ S904 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_697_ (
  .in1({ S904, S899 }),
  .out1({ S905 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_719_ (
  .in1({ S903, S900 }),
  .out1({ S906 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_720_ (
  .in1({ S151, DP_AC_q_1 }),
  .out1({ S907 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_698_ (
  .in1({ S156, S142 }),
  .out1({ S908 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_721_ (
  .in1({ S155, S141 }),
  .out1({ S909 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_699_ (
  .in1({ S909, S884 }),
  .out1({ S910 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_722_ (
  .in1({ S908, S883 }),
  .out1({ S911 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_700_ (
  .in1({ S895, S879 }),
  .out1({ S912 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_723_ (
  .in1({ S896, S880 }),
  .out1({ S913 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_701_ (
  .in1({ S912, S897 }),
  .out1({ S914 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_724_ (
  .in1({ S913, S898 }),
  .out1({ S915 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_702_ (
  .in1({ S915, S911 }),
  .out1({ S916 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_725_ (
  .in1({ S914, S910 }),
  .out1({ S917 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_703_ (
  .in1({ S903, S900 }),
  .out1({ S918 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_726_ (
  .in1({ S904, S899 }),
  .out1({ S919 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_704_ (
  .in1({ S918, S905 }),
  .out1({ S920 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_727_ (
  .in1({ S919, S906 }),
  .out1({ S921 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_705_ (
  .in1({ S921, S917 }),
  .out1({ S922 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_706_ (
  .in1({ S922, S905 }),
  .out1({ S923 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_224_ (
  .in1({ S923 }),
  .out1({ S924 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_728_ (
  .in1({ S873, S868 }),
  .out1({ S925 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_729_ (
  .in1({ S925, S874 }),
  .out1({ S926 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_225_ (
  .in1({ S926 }),
  .out1({ S927 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_707_ (
  .in1({ S926, S923 }),
  .out1({ S928 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_730_ (
  .in1({ S927, S924 }),
  .out1({ S929 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_708_ (
  .in1({ S928, S875 }),
  .out1({ S930 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_731_ (
  .in1({ S929, S874 }),
  .out1({ S931 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_709_ (
  .in1({ S930, S839 }),
  .out1({ S932 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_732_ (
  .in1({ S931, S838 }),
  .out1({ S933 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_710_ (
  .in1({ S932, S834 }),
  .out1({ S934 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_733_ (
  .in1({ S933, S835 }),
  .out1({ S935 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_711_ (
  .in1({ S934, S788 }),
  .out1({ S936 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_734_ (
  .in1({ S935, S787 }),
  .out1({ S937 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_712_ (
  .in1({ S936, S784 }),
  .out1({ S938 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_735_ (
  .in1({ S937, S785 }),
  .out1({ S939 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_713_ (
  .in1({ S938, S726 }),
  .out1({ S940 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_714_ (
  .in1({ S940, S721 }),
  .out1({ S941 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_736_ (
  .in1({ S646, S643 }),
  .out1({ S942 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_737_ (
  .in1({ S942, S648 }),
  .out1({ S943 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_715_ (
  .in1({ S943, S941 }),
  .out1({ S944 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_226_ (
  .in1({ S944 }),
  .out1({ S945 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_716_ (
  .in1({ S944, S649 }),
  .out1({ S946 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_738_ (
  .in1({ S945, S648 }),
  .out1({ S947 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_717_ (
  .in1({ S946, S574 }),
  .out1({ S948 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_739_ (
  .in1({ S947, S573 }),
  .out1({ S949 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_718_ (
  .in1({ S948, S570 }),
  .out1({ S950 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_740_ (
  .in1({ S949, S571 }),
  .out1({ S951 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_719_ (
  .in1({ S950, S497 }),
  .out1({ S952 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_741_ (
  .in1({ S951, S496 }),
  .out1({ S953 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_720_ (
  .in1({ S952, S494 }),
  .out1({ S954 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_721_ (
  .in1({ S954, S413 }),
  .out1({ S955 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_227_ (
  .in1({ S955 }),
  .out1({ S956 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_722_ (
  .in1({ S955, S411 }),
  .out1({ S957 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_742_ (
  .in1({ S956, S410 }),
  .out1({ S958 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_723_ (
  .in1({ S957, S352 }),
  .out1({ S959 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_743_ (
  .in1({ S958, S351 }),
  .out1({ S960 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_724_ (
  .in1({ S959, S349 }),
  .out1({ S961 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_744_ (
  .in1({ S345, S335 }),
  .out1({ S962 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_228_ (
  .in1({ S962 }),
  .out1({ S963 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_725_ (
  .in1({ S2534, S2523 }),
  .out1({ S964 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_745_ (
  .in1({ S2535, S2522 }),
  .out1({ S965 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_746_ (
  .in1({ S965, S963 }),
  .out1({ S966 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_747_ (
  .in1({ S964, S962 }),
  .out1({ S967 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_748_ (
  .in1({ S967, S966 }),
  .out1({ S968 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_726_ (
  .in1({ S968, S346 }),
  .out1({ S969 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_229_ (
  .in1({ S969 }),
  .out1({ S970 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_749_ (
  .in1({ S968, S346 }),
  .out1({ S971 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_750_ (
  .in1({ S971, S970 }),
  .out1({ S972 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_727_ (
  .in1({ S972, S961 }),
  .out1({ S973 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_728_ (
  .in1({ S973, S2432 }),
  .out1({ S974 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_751_ (
  .in1({ S962, S2522 }),
  .out1({ S975 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_752_ (
  .in1({ S975, S330 }),
  .out1({ S976 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_729_ (
  .in1({ S976, S969 }),
  .out1({ S977 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_753_ (
  .in1({ S977, S974 }),
  .out1({ S978 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_754_ (
  .in1({ S978, S204 }),
  .out1({ S979 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_230_ (
  .in1({ S979 }),
  .out1({ S980 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_730_ (
  .in1({ S979, S2411 }),
  .out1({ S981 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_755_ (
  .in1({ S2400, CU_inst_2 }),
  .out1({ S982 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_756_ (
  .in1({ S982, S2406 }),
  .out1({ S983 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_731_ (
  .in1({ S983, S981 }),
  .out1({ S984 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_732_ (
  .in1({ S984, S2407 }),
  .out1({ S20 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_733_ (
  .in1({ S2421, S1814 }),
  .out1({ S985 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_757_ (
  .in1({ S2422, S1825 }),
  .out1({ S986 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_758_ (
  .in1({ S985, DP_INC_1_in_0 }),
  .out1({ S987 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_734_ (
  .in1({ S2294, S1954 }),
  .out1({ S988 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_759_ (
  .in1({ S2293, S1953 }),
  .out1({ S989 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_760_ (
  .in1({ S2420, S1908 }),
  .out1({ S990 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_735_ (
  .in1({ CU_inst_6, S1160 }),
  .out1({ S991 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_761_ (
  .in1({ S991, S1916 }),
  .out1({ S992 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_736_ (
  .in1({ S992, S2271 }),
  .out1({ S993 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_737_ (
  .in1({ S993, S990 }),
  .out1({ S994 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_231_ (
  .in1({ S994 }),
  .out1({ S995 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_738_ (
  .in1({ S994, S1814 }),
  .out1({ S996 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_762_ (
  .in1({ S995, S1825 }),
  .out1({ S997 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_763_ (
  .in1({ S989, S1951 }),
  .out1({ S998 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_739_ (
  .in1({ S989, S1183 }),
  .out1({ S999 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_740_ (
  .in1({ S999, S997 }),
  .out1({ S1000 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_764_ (
  .in1({ S1000, S998 }),
  .out1({ S1001 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_741_ (
  .in1({ S996, S2118 }),
  .out1({ S1002 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_742_ (
  .in1({ S1002, S985 }),
  .out1({ S1003 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_765_ (
  .in1({ S1003, S1001 }),
  .out1({ S1004 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_766_ (
  .in1({ S1004, S987 }),
  .out1({ S21 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_767_ (
  .in1({ S985, DP_INC_1_in_1 }),
  .out1({ S1005 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_768_ (
  .in1({ S989, S1964 }),
  .out1({ S1006 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_743_ (
  .in1({ S989, S2538[1] }),
  .out1({ S1007 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_744_ (
  .in1({ S1007, S997 }),
  .out1({ S1008 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_769_ (
  .in1({ S1008, S1006 }),
  .out1({ S1009 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_770_ (
  .in1({ S997, S2127 }),
  .out1({ S1010 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_771_ (
  .in1({ S1010, S1009 }),
  .out1({ S1011 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_772_ (
  .in1({ S1011, S986 }),
  .out1({ S1012 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_773_ (
  .in1({ S1012, S1005 }),
  .out1({ S22 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_774_ (
  .in1({ S985, DP_INC_1_in_2 }),
  .out1({ S1013 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_745_ (
  .in1({ S988, S1971 }),
  .out1({ S1014 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_775_ (
  .in1({ S988, S2538[2] }),
  .out1({ S1015 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_776_ (
  .in1({ S1015, S996 }),
  .out1({ S1016 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_746_ (
  .in1({ S1016, S1014 }),
  .out1({ S1017 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_747_ (
  .in1({ S996, S2136 }),
  .out1({ S1018 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_748_ (
  .in1({ S1018, S1017 }),
  .out1({ S1019 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_777_ (
  .in1({ S1019, S986 }),
  .out1({ S1020 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_778_ (
  .in1({ S1020, S1013 }),
  .out1({ S23 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_749_ (
  .in1({ S986, DP_INC_1_in_3 }),
  .out1({ S1021 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_779_ (
  .in1({ S989, S1979 }),
  .out1({ S1022 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_750_ (
  .in1({ S989, S2538[3] }),
  .out1({ S1023 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_780_ (
  .in1({ S997, S2145 }),
  .out1({ S1024 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_751_ (
  .in1({ S1023, S997 }),
  .out1({ S1025 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_781_ (
  .in1({ S1025, S1022 }),
  .out1({ S1026 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_782_ (
  .in1({ S1026, S1024 }),
  .out1({ S1027 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_752_ (
  .in1({ S1027, S985 }),
  .out1({ S1028 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_753_ (
  .in1({ S1028, S1021 }),
  .out1({ S24 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_783_ (
  .in1({ S985, DP_INC_1_in_4 }),
  .out1({ S1029 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_754_ (
  .in1({ S988, S1989 }),
  .out1({ S1030 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_784_ (
  .in1({ S988, S2538[4] }),
  .out1({ S1031 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_785_ (
  .in1({ S997, S2155 }),
  .out1({ S1032 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_786_ (
  .in1({ S1031, S996 }),
  .out1({ S1033 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_755_ (
  .in1({ S1033, S1030 }),
  .out1({ S1034 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_756_ (
  .in1({ S1034, S985 }),
  .out1({ S1035 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_787_ (
  .in1({ S1035, S1032 }),
  .out1({ S1036 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_788_ (
  .in1({ S1036, S1029 }),
  .out1({ S25 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_789_ (
  .in1({ S985, DP_INC_1_in_5 }),
  .out1({ S1037 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_790_ (
  .in1({ S997, S2164 }),
  .out1({ S1038 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_757_ (
  .in1({ S989, S2538[5] }),
  .out1({ S1039 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_758_ (
  .in1({ S988, S1997 }),
  .out1({ S1040 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_759_ (
  .in1({ S1040, S1039 }),
  .out1({ S1041 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_760_ (
  .in1({ S1041, S997 }),
  .out1({ S1042 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_761_ (
  .in1({ S1042, S985 }),
  .out1({ S1043 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_791_ (
  .in1({ S1043, S1038 }),
  .out1({ S1044 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_792_ (
  .in1({ S1044, S1037 }),
  .out1({ S26 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_762_ (
  .in1({ S986, DP_INC_1_in_6 }),
  .out1({ S1045 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_763_ (
  .in1({ S996, S2173 }),
  .out1({ S1046 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_793_ (
  .in1({ S988, S2538[6] }),
  .out1({ S1047 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_794_ (
  .in1({ S989, S2004 }),
  .out1({ S1048 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_795_ (
  .in1({ S1048, S1047 }),
  .out1({ S1049 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_796_ (
  .in1({ S1049, S996 }),
  .out1({ S1050 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_797_ (
  .in1({ S1050, S986 }),
  .out1({ S1051 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_764_ (
  .in1({ S1051, S1046 }),
  .out1({ S1052 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_765_ (
  .in1({ S1052, S1045 }),
  .out1({ S27 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_766_ (
  .in1({ S986, DP_INC_1_in_7 }),
  .out1({ S1053 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_767_ (
  .in1({ S996, S2182 }),
  .out1({ S1054 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_798_ (
  .in1({ S988, S2538[7] }),
  .out1({ S1055 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_799_ (
  .in1({ S989, S2011 }),
  .out1({ S1056 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_800_ (
  .in1({ S1056, S1055 }),
  .out1({ S1057 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_801_ (
  .in1({ S1057, S996 }),
  .out1({ S1058 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_802_ (
  .in1({ S1058, S986 }),
  .out1({ S1059 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_768_ (
  .in1({ S1059, S1054 }),
  .out1({ S1060 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_769_ (
  .in1({ S1060, S1053 }),
  .out1({ S28 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_770_ (
  .in1({ S986, DP_INC_1_in_8 }),
  .out1({ S1061 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_771_ (
  .in1({ S996, S2191 }),
  .out1({ S1062 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_803_ (
  .in1({ S988, S2538[8] }),
  .out1({ S1064 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_804_ (
  .in1({ S989, S2018 }),
  .out1({ S1065 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_805_ (
  .in1({ S1065, S1064 }),
  .out1({ S1066 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_806_ (
  .in1({ S1066, S996 }),
  .out1({ S1067 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_807_ (
  .in1({ S1067, S986 }),
  .out1({ S1068 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_772_ (
  .in1({ S1068, S1062 }),
  .out1({ S1069 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_773_ (
  .in1({ S1069, S1061 }),
  .out1({ S29 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_774_ (
  .in1({ S986, DP_INC_1_in_9 }),
  .out1({ S1070 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_775_ (
  .in1({ S996, S2200 }),
  .out1({ S1071 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_808_ (
  .in1({ S988, S2538[9] }),
  .out1({ S1072 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_809_ (
  .in1({ S989, S2025 }),
  .out1({ S1074 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_810_ (
  .in1({ S1074, S1072 }),
  .out1({ S1075 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_811_ (
  .in1({ S1075, S996 }),
  .out1({ S1076 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_812_ (
  .in1({ S1076, S986 }),
  .out1({ S1077 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_776_ (
  .in1({ S1077, S1071 }),
  .out1({ S1078 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_777_ (
  .in1({ S1078, S1070 }),
  .out1({ S30 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_813_ (
  .in1({ S985, DP_INC_1_in_10 }),
  .out1({ S1079 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_814_ (
  .in1({ S997, S2209 }),
  .out1({ S1080 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_778_ (
  .in1({ S989, S2538[10] }),
  .out1({ S1081 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_779_ (
  .in1({ S988, S2032 }),
  .out1({ S1082 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_780_ (
  .in1({ S1082, S1081 }),
  .out1({ S1084 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_781_ (
  .in1({ S1084, S997 }),
  .out1({ S1085 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_782_ (
  .in1({ S1085, S985 }),
  .out1({ S1086 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_815_ (
  .in1({ S1086, S1080 }),
  .out1({ S1087 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_816_ (
  .in1({ S1087, S1079 }),
  .out1({ S31 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_817_ (
  .in1({ S985, DP_INC_1_in_11 }),
  .out1({ S1088 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_818_ (
  .in1({ S997, S2218 }),
  .out1({ S1089 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_783_ (
  .in1({ S988, S2040 }),
  .out1({ S1090 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_819_ (
  .in1({ S988, S2538[11] }),
  .out1({ S1091 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_820_ (
  .in1({ S1091, S996 }),
  .out1({ S1092 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_784_ (
  .in1({ S1092, S1090 }),
  .out1({ S1094 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_785_ (
  .in1({ S1094, S985 }),
  .out1({ S1095 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_821_ (
  .in1({ S1095, S1089 }),
  .out1({ S1096 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_822_ (
  .in1({ S1096, S1088 }),
  .out1({ S32 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_823_ (
  .in1({ S985, DP_INC_1_in_12 }),
  .out1({ S1097 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_824_ (
  .in1({ S997, S2227 }),
  .out1({ S1098 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_786_ (
  .in1({ S988, S2050 }),
  .out1({ S1099 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_825_ (
  .in1({ S988, S2538[12] }),
  .out1({ S1100 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_826_ (
  .in1({ S1100, S996 }),
  .out1({ S1101 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_787_ (
  .in1({ S1101, S1099 }),
  .out1({ S1102 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_788_ (
  .in1({ S1102, S985 }),
  .out1({ S1104 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_827_ (
  .in1({ S1104, S1098 }),
  .out1({ S1105 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_828_ (
  .in1({ S1105, S1097 }),
  .out1({ S33 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_829_ (
  .in1({ S985, DP_INC_1_in_13 }),
  .out1({ S1106 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_830_ (
  .in1({ S997, S2236 }),
  .out1({ S1107 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_789_ (
  .in1({ S988, S2058 }),
  .out1({ S1108 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_831_ (
  .in1({ S988, S2538[13] }),
  .out1({ S1109 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_832_ (
  .in1({ S1109, S996 }),
  .out1({ S1110 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_790_ (
  .in1({ S1110, S1108 }),
  .out1({ S1111 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_791_ (
  .in1({ S1111, S985 }),
  .out1({ S1112 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_833_ (
  .in1({ S1112, S1107 }),
  .out1({ S1114 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_834_ (
  .in1({ S1114, S1106 }),
  .out1({ S34 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_835_ (
  .in1({ S985, DP_INC_1_in_14 }),
  .out1({ S1115 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_836_ (
  .in1({ S997, S2244 }),
  .out1({ S1116 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_792_ (
  .in1({ S988, S2066 }),
  .out1({ S1117 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_837_ (
  .in1({ S988, S2538[14] }),
  .out1({ S1118 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_838_ (
  .in1({ S1118, S996 }),
  .out1({ S1119 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_793_ (
  .in1({ S1119, S1117 }),
  .out1({ S1120 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_794_ (
  .in1({ S1120, S985 }),
  .out1({ S1121 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_839_ (
  .in1({ S1121, S1116 }),
  .out1({ S1122 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_840_ (
  .in1({ S1122, S1115 }),
  .out1({ S35 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_841_ (
  .in1({ S985, DP_INC_1_in_15 }),
  .out1({ S1124 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_842_ (
  .in1({ S997, S2253 }),
  .out1({ S1125 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_795_ (
  .in1({ S988, S2075 }),
  .out1({ S1126 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_843_ (
  .in1({ S988, S2538[15] }),
  .out1({ S1127 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_844_ (
  .in1({ S1127, S996 }),
  .out1({ S1128 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_796_ (
  .in1({ S1128, S1126 }),
  .out1({ S1129 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_797_ (
  .in1({ S1129, S985 }),
  .out1({ S1130 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_845_ (
  .in1({ S1130, S1125 }),
  .out1({ S1131 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_846_ (
  .in1({ S1131, S1124 }),
  .out1({ S36 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_798_ (
  .in1({ S1902, S1883 }),
  .out1({ S1133 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_799_ (
  .in1({ S1133, S2081 }),
  .out1({ S1134 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_800_ (
  .in1({ S1883, S1160 }),
  .out1({ S1135 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_847_ (
  .in1({ S1135, S2404 }),
  .out1({ S1136 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_848_ (
  .in1({ S1136, S1134 }),
  .out1({ S1137 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_801_ (
  .in1({ S1137, DP_SR_C_q }),
  .out1({ S1138 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_802_ (
  .in1({ S201, S2446 }),
  .out1({ S1139 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_803_ (
  .in1({ S1139, S2431 }),
  .out1({ S1140 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_849_ (
  .in1({ S2400, CU_inst_1 }),
  .out1({ S1141 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_850_ (
  .in1({ S1141, S1137 }),
  .out1({ S1142 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_804_ (
  .in1({ S1142, S1140 }),
  .out1({ S1144 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_805_ (
  .in1({ S1144, S1138 }),
  .out1({ S37 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_851_ (
  .in1({ S2412, DP_AC_q_15 }),
  .out1({ S1145 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_806_ (
  .in1({ S1145, S980 }),
  .out1({ S1146 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_852_ (
  .in1({ S2400, CU_inst_4 }),
  .out1({ S1147 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_853_ (
  .in1({ S1147, S1134 }),
  .out1({ S1148 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_854_ (
  .in1({ S2400, CU_inst_0 }),
  .out1({ S1149 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_855_ (
  .in1({ S1149, S1148 }),
  .out1({ S1150 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_807_ (
  .in1({ S1150, S1146 }),
  .out1({ S1151 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_808_ (
  .in1({ S1148, DP_SR_V_q }),
  .out1({ S1152 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_809_ (
  .in1({ S1152, S1151 }),
  .out1({ S38 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_856_ (
  .in1({ CU_nstate_0, S2538[0] }),
  .out1({ S1154 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_857_ (
  .in1({ S1731, CU_inst_0 }),
  .out1({ S1155 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_858_ (
  .in1({ S1155, S1154 }),
  .out1({ S39 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_859_ (
  .in1({ CU_nstate_0, S2538[1] }),
  .out1({ S1156 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_860_ (
  .in1({ S1731, CU_inst_1 }),
  .out1({ S1157 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_861_ (
  .in1({ S1157, S1156 }),
  .out1({ S40 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_862_ (
  .in1({ CU_nstate_0, S2538[2] }),
  .out1({ S1158 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_863_ (
  .in1({ S1731, CU_inst_2 }),
  .out1({ S1159 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_864_ (
  .in1({ S1159, S1158 }),
  .out1({ S41 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_865_ (
  .in1({ CU_nstate_0, S2538[3] }),
  .out1({ S1161 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_866_ (
  .in1({ S1731, CU_inst_3 }),
  .out1({ S1162 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_867_ (
  .in1({ S1162, S1161 }),
  .out1({ S42 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_868_ (
  .in1({ CU_nstate_0, S2538[4] }),
  .out1({ S1163 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_869_ (
  .in1({ S1731, CU_inst_4 }),
  .out1({ S1164 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_870_ (
  .in1({ S1164, S1163 }),
  .out1({ S43 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_871_ (
  .in1({ CU_nstate_0, S2538[5] }),
  .out1({ S1165 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_872_ (
  .in1({ S1731, CU_inst_5 }),
  .out1({ S1166 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_873_ (
  .in1({ S1166, S1165 }),
  .out1({ S44 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_874_ (
  .in1({ CU_nstate_0, S2538[6] }),
  .out1({ S1167 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_875_ (
  .in1({ S1731, CU_inst_6 }),
  .out1({ S1169 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_876_ (
  .in1({ S1169, S1167 }),
  .out1({ S45 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_877_ (
  .in1({ CU_nstate_0, S2538[7] }),
  .out1({ S1170 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_878_ (
  .in1({ S1731, CU_inst_7 }),
  .out1({ S1171 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_879_ (
  .in1({ S1171, S1170 }),
  .out1({ S46 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_880_ (
  .in1({ CU_nstate_0, S2538[8] }),
  .out1({ S1172 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_881_ (
  .in1({ S1731, CU_inst_8 }),
  .out1({ S1173 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_882_ (
  .in1({ S1173, S1172 }),
  .out1({ S47 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_883_ (
  .in1({ CU_nstate_0, S2538[9] }),
  .out1({ S1174 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_884_ (
  .in1({ S1731, CU_inst_9 }),
  .out1({ S1175 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_885_ (
  .in1({ S1175, S1174 }),
  .out1({ S48 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_886_ (
  .in1({ CU_nstate_0, S2538[10] }),
  .out1({ S1177 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_887_ (
  .in1({ S1731, CU_inst_10 }),
  .out1({ S1178 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_888_ (
  .in1({ S1178, S1177 }),
  .out1({ S49 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_889_ (
  .in1({ CU_nstate_0, S2538[11] }),
  .out1({ S1179 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_890_ (
  .in1({ S1731, CU_inst_11 }),
  .out1({ S1180 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_891_ (
  .in1({ S1180, S1179 }),
  .out1({ S50 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_892_ (
  .in1({ CU_nstate_0, S2538[12] }),
  .out1({ S1181 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_893_ (
  .in1({ S1731, CU_inst_12 }),
  .out1({ S1182 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_894_ (
  .in1({ S1182, S1181 }),
  .out1({ S51 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_895_ (
  .in1({ CU_nstate_0, S2538[13] }),
  .out1({ S1184 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_896_ (
  .in1({ S1731, CU_inst_13 }),
  .out1({ S1185 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_897_ (
  .in1({ S1185, S1184 }),
  .out1({ S52 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_898_ (
  .in1({ CU_nstate_0, S2538[14] }),
  .out1({ S1186 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_899_ (
  .in1({ S1731, CU_inst_14 }),
  .out1({ S1187 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_900_ (
  .in1({ S1187, S1186 }),
  .out1({ S53 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_901_ (
  .in1({ CU_nstate_0, S2538[15] }),
  .out1({ S1188 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_902_ (
  .in1({ S1731, CU_inst_15 }),
  .out1({ S1189 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_903_ (
  .in1({ S1189, S1188 }),
  .out1({ S54 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_904_ (
  .in1({ S2404, CU_inst_7 }),
  .out1({ S1190 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_905_ (
  .in1({ S1190, S2419 }),
  .out1({ S1192 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_810_ (
  .in1({ S1192, S2396 }),
  .out1({ S1193 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_811_ (
  .in1({ S1193, S1883 }),
  .out1({ S1194 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_812_ (
  .in1({ S1194, S2081 }),
  .out1({ S1195 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_232_ (
  .in1({ S1195 }),
  .out1({ S1196 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_813_ (
  .in1({ S1196, DP_SR_Z_q }),
  .out1({ S1197 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_906_ (
  .in1({ S972, S961 }),
  .out1({ S1198 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_907_ (
  .in1({ S1198, S974 }),
  .out1({ S1199 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_814_ (
  .in1({ S196, S2457 }),
  .out1({ S1200 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_815_ (
  .in1({ S1200, S198 }),
  .out1({ S1201 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_908_ (
  .in1({ S1201, S2432 }),
  .out1({ S1203 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_909_ (
  .in1({ S1203, S1199 }),
  .out1({ S1204 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_910_ (
  .in1({ S2473, S2467 }),
  .out1({ S1205 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_816_ (
  .in1({ S1205, S192 }),
  .out1({ S1206 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_817_ (
  .in1({ S194, S2431 }),
  .out1({ S1207 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_911_ (
  .in1({ S1207, S193 }),
  .out1({ S1208 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_818_ (
  .in1({ S1208, S1206 }),
  .out1({ S1209 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_819_ (
  .in1({ S958, S351 }),
  .out1({ S1210 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_912_ (
  .in1({ S960, S2431 }),
  .out1({ S1211 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_820_ (
  .in1({ S1211, S1210 }),
  .out1({ S1212 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_821_ (
  .in1({ S1212, S1209 }),
  .out1({ S1214 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_822_ (
  .in1({ S190, S2476 }),
  .out1({ S1215 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_823_ (
  .in1({ S1215, S192 }),
  .out1({ S1216 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_913_ (
  .in1({ S1216, S2432 }),
  .out1({ S1217 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_914_ (
  .in1({ S954, S413 }),
  .out1({ S1218 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_824_ (
  .in1({ S955, S2432 }),
  .out1({ S1219 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_915_ (
  .in1({ S1219, S1218 }),
  .out1({ S1220 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_916_ (
  .in1({ S1220, S1217 }),
  .out1({ S1221 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_825_ (
  .in1({ S2493, S2485 }),
  .out1({ S1222 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_917_ (
  .in1({ S1222, S185 }),
  .out1({ S1223 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_918_ (
  .in1({ S188, S2432 }),
  .out1({ S1225 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_826_ (
  .in1({ S1225, S187 }),
  .out1({ S1226 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_919_ (
  .in1({ S1226, S1223 }),
  .out1({ S1227 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_233_ (
  .in1({ S1227 }),
  .out1({ S1228 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_827_ (
  .in1({ S951, S496 }),
  .out1({ S1229 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_920_ (
  .in1({ S953, S2431 }),
  .out1({ S1230 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_828_ (
  .in1({ S1230, S1229 }),
  .out1({ S1231 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_234_ (
  .in1({ S1231 }),
  .out1({ S1232 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_829_ (
  .in1({ S1231, S1228 }),
  .out1({ S1233 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_921_ (
  .in1({ S1232, S1227 }),
  .out1({ S1234 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_922_ (
  .in1({ S946, S574 }),
  .out1({ S1236 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_830_ (
  .in1({ S184, S2495 }),
  .out1({ S1237 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_831_ (
  .in1({ S1237, S186 }),
  .out1({ S1238 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_832_ (
  .in1({ S948, S2432 }),
  .out1({ S1239 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_923_ (
  .in1({ S1239, S1236 }),
  .out1({ S1240 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_924_ (
  .in1({ S1238, S2432 }),
  .out1({ S1241 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_925_ (
  .in1({ S1241, S1240 }),
  .out1({ S1242 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_926_ (
  .in1({ S943, S941 }),
  .out1({ S1243 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_833_ (
  .in1({ S944, S2432 }),
  .out1({ S1244 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_927_ (
  .in1({ S1244, S1243 }),
  .out1({ S1245 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_834_ (
  .in1({ S2503, S2502 }),
  .out1({ S1247 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_928_ (
  .in1({ S1247, S182 }),
  .out1({ S1248 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_835_ (
  .in1({ S1247, S182 }),
  .out1({ S1249 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_836_ (
  .in1({ S1249, S2431 }),
  .out1({ S1250 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_929_ (
  .in1({ S1250, S1248 }),
  .out1({ S1251 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_930_ (
  .in1({ S1251, S1245 }),
  .out1({ S1252 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_837_ (
  .in1({ S939, S725 }),
  .out1({ S1253 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_838_ (
  .in1({ S1253, S940 }),
  .out1({ S1254 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_839_ (
  .in1({ S1254, S2432 }),
  .out1({ S1255 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_235_ (
  .in1({ S1255 }),
  .out1({ S1256 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_931_ (
  .in1({ S179, S2514 }),
  .out1({ S1258 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_932_ (
  .in1({ S1258, S181 }),
  .out1({ S1259 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_933_ (
  .in1({ S1259, S2432 }),
  .out1({ S1260 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_934_ (
  .in1({ S1260, S1256 }),
  .out1({ S1261 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_935_ (
  .in1({ S934, S788 }),
  .out1({ S1262 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_840_ (
  .in1({ S175, S2525 }),
  .out1({ S1263 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_841_ (
  .in1({ S1263, S177 }),
  .out1({ S1264 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_936_ (
  .in1({ S1264, S2432 }),
  .out1({ S1265 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_842_ (
  .in1({ S936, S2432 }),
  .out1({ S1266 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_937_ (
  .in1({ S1266, S1262 }),
  .out1({ S1267 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_938_ (
  .in1({ S1267, S1265 }),
  .out1({ S1269 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_939_ (
  .in1({ S930, S839 }),
  .out1({ S1270 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_940_ (
  .in1({ S1270, S933 }),
  .out1({ S1271 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_941_ (
  .in1({ S1271, S2431 }),
  .out1({ S1272 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_942_ (
  .in1({ S172, S75 }),
  .out1({ S1273 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_943_ (
  .in1({ S1273, S174 }),
  .out1({ S1274 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_944_ (
  .in1({ S1274, S2432 }),
  .out1({ S1275 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_945_ (
  .in1({ S1275, S1272 }),
  .out1({ S1276 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_946_ (
  .in1({ S926, S923 }),
  .out1({ S1277 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_947_ (
  .in1({ S1277, S929 }),
  .out1({ S1278 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_948_ (
  .in1({ S1278, S2431 }),
  .out1({ S1280 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_843_ (
  .in1({ S86, S84 }),
  .out1({ S1281 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_949_ (
  .in1({ S1281, S170 }),
  .out1({ S1282 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_844_ (
  .in1({ S1281, S170 }),
  .out1({ S1283 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_845_ (
  .in1({ S1283, S2431 }),
  .out1({ S1284 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_950_ (
  .in1({ S1284, S1282 }),
  .out1({ S1285 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_951_ (
  .in1({ S1285, S1280 }),
  .out1({ S1286 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_846_ (
  .in1({ S920, S916 }),
  .out1({ S1287 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_847_ (
  .in1({ S1287, S922 }),
  .out1({ S1288 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_848_ (
  .in1({ S1288, S2432 }),
  .out1({ S1289 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_849_ (
  .in1({ S168, S101 }),
  .out1({ S1291 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_850_ (
  .in1({ S1291, S169 }),
  .out1({ S1292 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_851_ (
  .in1({ S1292, S2431 }),
  .out1({ S1293 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_852_ (
  .in1({ S1293, S1289 }),
  .out1({ S1294 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_952_ (
  .in1({ S915, S911 }),
  .out1({ S1295 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_953_ (
  .in1({ S1295, S917 }),
  .out1({ S1296 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_954_ (
  .in1({ S1296, S2431 }),
  .out1({ S1297 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_955_ (
  .in1({ S116, S114 }),
  .out1({ S1298 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_956_ (
  .in1({ S1298, S163 }),
  .out1({ S1299 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_957_ (
  .in1({ S165, S114 }),
  .out1({ S1300 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_958_ (
  .in1({ S1300, S1299 }),
  .out1({ S1302 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_959_ (
  .in1({ S1302, S2432 }),
  .out1({ S1303 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_960_ (
  .in1({ S1303, S1297 }),
  .out1({ S1304 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_961_ (
  .in1({ S156, S141 }),
  .out1({ S1305 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_853_ (
  .in1({ S1305, S883 }),
  .out1({ S1306 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_962_ (
  .in1({ S1305, S883 }),
  .out1({ S1307 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_854_ (
  .in1({ S160, S130 }),
  .out1({ S1308 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_963_ (
  .in1({ S159, S131 }),
  .out1({ S1309 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_855_ (
  .in1({ S1308, S161 }),
  .out1({ S1310 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_964_ (
  .in1({ S1309, S162 }),
  .out1({ S1311 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_965_ (
  .in1({ S1307, S2431 }),
  .out1({ S1313 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_856_ (
  .in1({ S1313, S1306 }),
  .out1({ S1314 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_236_ (
  .in1({ S1314 }),
  .out1({ S1315 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_857_ (
  .in1({ S1311, S2431 }),
  .out1({ S1316 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_966_ (
  .in1({ S1310, S2432 }),
  .out1({ S1317 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_967_ (
  .in1({ S1317, S1315 }),
  .out1({ S1318 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_858_ (
  .in1({ S1316, S1314 }),
  .out1({ S1319 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_968_ (
  .in1({ S842, S792 }),
  .out1({ S1320 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_969_ (
  .in1({ S1320, S909 }),
  .out1({ S1321 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_970_ (
  .in1({ S1321, S2431 }),
  .out1({ S1322 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_971_ (
  .in1({ S156, S146 }),
  .out1({ S1324 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_972_ (
  .in1({ S1324, S158 }),
  .out1({ S1325 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_973_ (
  .in1({ S1325, S2432 }),
  .out1({ S1326 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_974_ (
  .in1({ S1326, S1322 }),
  .out1({ S1327 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_859_ (
  .in1({ S154, DP_AC_q_0 }),
  .out1({ S1328 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_860_ (
  .in1({ S155, S2431 }),
  .out1({ S1329 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_861_ (
  .in1({ S156, S2432 }),
  .out1({ S1330 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_862_ (
  .in1({ S1330, S1329 }),
  .out1({ S1331 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_863_ (
  .in1({ S1331, S1328 }),
  .out1({ S1332 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_864_ (
  .in1({ S1332, S2411 }),
  .out1({ S1333 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_975_ (
  .in1({ S1333, S1327 }),
  .out1({ S1335 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_865_ (
  .in1({ S1335, S1318 }),
  .out1({ S1336 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_976_ (
  .in1({ S1336, S1304 }),
  .out1({ S1337 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_866_ (
  .in1({ S1337, S1294 }),
  .out1({ S1338 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_977_ (
  .in1({ S1338, S1286 }),
  .out1({ S1339 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_237_ (
  .in1({ S1339 }),
  .out1({ S1340 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_978_ (
  .in1({ S1340, S1276 }),
  .out1({ S1341 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_867_ (
  .in1({ S1341, S1269 }),
  .out1({ S1342 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_979_ (
  .in1({ S1342, S1261 }),
  .out1({ S1343 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_868_ (
  .in1({ S1343, S1252 }),
  .out1({ S1344 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_238_ (
  .in1({ S1344 }),
  .out1({ S1346 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_869_ (
  .in1({ S1346, S1242 }),
  .out1({ S1347 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_980_ (
  .in1({ S1347, S1233 }),
  .out1({ S1348 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_870_ (
  .in1({ S1348, S1221 }),
  .out1({ S1349 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_981_ (
  .in1({ S1349, S1214 }),
  .out1({ S1350 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_871_ (
  .in1({ S1350, S1204 }),
  .out1({ S1351 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_982_ (
  .in1({ S1351, S979 }),
  .out1({ S1352 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_983_ (
  .in1({ S2400, CU_inst_3 }),
  .out1({ S1353 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_984_ (
  .in1({ S1353, S1352 }),
  .out1({ S1354 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_872_ (
  .in1({ S1354, S1195 }),
  .out1({ S1355 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_873_ (
  .in1({ S1355, S1197 }),
  .out1({ S55 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_874_ (
  .in1({ S2394, S1931 }),
  .out1({ S1357 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_239_ (
  .in1({ S1357 }),
  .out1({ S1358 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_875_ (
  .in1({ S1358, CU_inst_5 }),
  .out1({ S1359 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_876_ (
  .in1({ S2394, S1160 }),
  .out1({ S1360 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_985_ (
  .in1({ S2435, S2416 }),
  .out1({ S1361 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_877_ (
  .in1({ S1361, S1360 }),
  .out1({ S1362 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_878_ (
  .in1({ S1362, S2424 }),
  .out1({ S1363 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_879_ (
  .in1({ S1363, S2266 }),
  .out1({ S1364 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_240_ (
  .in1({ S1364 }),
  .out1({ S1365 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_880_ (
  .in1({ S1365, S1359 }),
  .out1({ S1367 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_986_ (
  .in1({ S1367, DP_AC_q_0 }),
  .out1({ S1368 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_881_ (
  .in1({ S1919, S1883 }),
  .out1({ S1369 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_987_ (
  .in1({ S1918, S1882 }),
  .out1({ S1370 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_988_ (
  .in1({ S1369, S1951 }),
  .out1({ S1371 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_882_ (
  .in1({ S2294, S1890 }),
  .out1({ S1372 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_989_ (
  .in1({ S1892, S1882 }),
  .out1({ S1373 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_883_ (
  .in1({ S1372, S1835 }),
  .out1({ S1374 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_990_ (
  .in1({ S1373, S1846 }),
  .out1({ S1375 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_884_ (
  .in1({ S2427, S2081 }),
  .out1({ S1376 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_991_ (
  .in1({ S2428, S2082 }),
  .out1({ S1378 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_992_ (
  .in1({ S152, DP_AC_q_0 }),
  .out1({ S1379 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_993_ (
  .in1({ S1379, S907 }),
  .out1({ S1380 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_885_ (
  .in1({ S1380, S136 }),
  .out1({ S1381 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_886_ (
  .in1({ S152, DP_AC_q_3 }),
  .out1({ S1382 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_887_ (
  .in1({ S151, DP_AC_q_2 }),
  .out1({ S1383 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_888_ (
  .in1({ S1383, S1382 }),
  .out1({ S1384 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_889_ (
  .in1({ S1384, S137 }),
  .out1({ S1385 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_890_ (
  .in1({ S1385, S1381 }),
  .out1({ S1386 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_891_ (
  .in1({ S1386, S121 }),
  .out1({ S1387 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_994_ (
  .in1({ S1357, CU_inst_5 }),
  .out1({ S1389 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_241_ (
  .in1({ S1389 }),
  .out1({ S1390 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_892_ (
  .in1({ S1390, S107 }),
  .out1({ S1391 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_995_ (
  .in1({ S1389, S108 }),
  .out1({ S1392 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_893_ (
  .in1({ S152, DP_AC_q_5 }),
  .out1({ S1393 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_894_ (
  .in1({ S151, DP_AC_q_4 }),
  .out1({ S1394 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_895_ (
  .in1({ S1394, S1393 }),
  .out1({ S1395 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_896_ (
  .in1({ S1395, S136 }),
  .out1({ S1396 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_897_ (
  .in1({ S152, DP_AC_q_7 }),
  .out1({ S1397 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_898_ (
  .in1({ S151, DP_AC_q_6 }),
  .out1({ S1398 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_899_ (
  .in1({ S1398, S1397 }),
  .out1({ S1400 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_900_ (
  .in1({ S1400, S137 }),
  .out1({ S1401 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_901_ (
  .in1({ S1401, S1396 }),
  .out1({ S1402 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_242_ (
  .in1({ S1402 }),
  .out1({ S1403 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_996_ (
  .in1({ S1403, S121 }),
  .out1({ S1404 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_997_ (
  .in1({ S1404, S1391 }),
  .out1({ S1405 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_902_ (
  .in1({ S1405, S1387 }),
  .out1({ S1406 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_903_ (
  .in1({ S1390, S108 }),
  .out1({ S1407 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_998_ (
  .in1({ S1389, S107 }),
  .out1({ S1408 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_904_ (
  .in1({ S152, DP_AC_q_9 }),
  .out1({ S1409 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_905_ (
  .in1({ S151, DP_AC_q_8 }),
  .out1({ S1411 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_906_ (
  .in1({ S1411, S1409 }),
  .out1({ S1412 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_907_ (
  .in1({ S1412, S136 }),
  .out1({ S1413 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_908_ (
  .in1({ S152, DP_AC_q_11 }),
  .out1({ S1414 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_909_ (
  .in1({ S151, DP_AC_q_10 }),
  .out1({ S1415 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_910_ (
  .in1({ S1415, S1414 }),
  .out1({ S1416 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_911_ (
  .in1({ S1416, S137 }),
  .out1({ S1417 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_912_ (
  .in1({ S1417, S1413 }),
  .out1({ S1418 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_913_ (
  .in1({ S1418, S121 }),
  .out1({ S1419 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_914_ (
  .in1({ S152, DP_AC_q_13 }),
  .out1({ S1420 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_915_ (
  .in1({ S151, DP_AC_q_12 }),
  .out1({ S1422 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_916_ (
  .in1({ S1422, S1420 }),
  .out1({ S1423 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_243_ (
  .in1({ S1423 }),
  .out1({ S1424 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_917_ (
  .in1({ S1423, S136 }),
  .out1({ S1425 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_918_ (
  .in1({ S152, DP_AC_q_15 }),
  .out1({ S1426 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_919_ (
  .in1({ S151, DP_AC_q_14 }),
  .out1({ S1427 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_920_ (
  .in1({ S1427, S1426 }),
  .out1({ S1428 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_921_ (
  .in1({ S1428, S137 }),
  .out1({ S1429 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_922_ (
  .in1({ S1429, S1425 }),
  .out1({ S1430 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_923_ (
  .in1({ S1430, S122 }),
  .out1({ S1431 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_924_ (
  .in1({ S1431, S1419 }),
  .out1({ S1433 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_999_ (
  .in1({ S1433, S1407 }),
  .out1({ S1434 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_925_ (
  .in1({ S1900, S1883 }),
  .out1({ S1435 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1000_ (
  .in1({ S1899, S1882 }),
  .out1({ S1436 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_926_ (
  .in1({ S1389, DP_AC_q_0 }),
  .out1({ S1437 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_927_ (
  .in1({ S1437, S1435 }),
  .out1({ S1438 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1001_ (
  .in1({ S1438, S1434 }),
  .out1({ S1439 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_928_ (
  .in1({ S1439, S1406 }),
  .out1({ S1440 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1002_ (
  .in1({ S1435, S878 }),
  .out1({ S1441 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1003_ (
  .in1({ S1378, S1332 }),
  .out1({ S1442 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1004_ (
  .in1({ S1441, S1376 }),
  .out1({ S1444 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_929_ (
  .in1({ S1444, S1440 }),
  .out1({ S1445 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1005_ (
  .in1({ S1442, S1374 }),
  .out1({ S1446 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_930_ (
  .in1({ S1446, S1445 }),
  .out1({ S1447 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_931_ (
  .in1({ S1374, S2538[0] }),
  .out1({ S1448 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_932_ (
  .in1({ S1448, S1447 }),
  .out1({ S1449 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1006_ (
  .in1({ S1449, S1370 }),
  .out1({ S1450 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1007_ (
  .in1({ S1450, S1371 }),
  .out1({ S1451 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1008_ (
  .in1({ S1451, S1365 }),
  .out1({ S1452 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1009_ (
  .in1({ S1452, S1368 }),
  .out1({ S56 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1010_ (
  .in1({ S1367, DP_AC_q_1 }),
  .out1({ S1454 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1011_ (
  .in1({ S152, DP_AC_q_1 }),
  .out1({ S1455 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1012_ (
  .in1({ S1455, S877 }),
  .out1({ S1456 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1013_ (
  .in1({ S1456, S137 }),
  .out1({ S1457 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_933_ (
  .in1({ S152, DP_AC_q_4 }),
  .out1({ S1458 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_934_ (
  .in1({ S151, DP_AC_q_3 }),
  .out1({ S1459 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_935_ (
  .in1({ S1459, S1458 }),
  .out1({ S1460 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1014_ (
  .in1({ S1460, S136 }),
  .out1({ S1461 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1015_ (
  .in1({ S1461, S1457 }),
  .out1({ S1462 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1016_ (
  .in1({ S1462, S122 }),
  .out1({ S1463 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_936_ (
  .in1({ S152, DP_AC_q_6 }),
  .out1({ S1465 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_937_ (
  .in1({ S151, DP_AC_q_5 }),
  .out1({ S1466 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_938_ (
  .in1({ S1466, S1465 }),
  .out1({ S1467 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_939_ (
  .in1({ S1467, S136 }),
  .out1({ S1468 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_940_ (
  .in1({ S152, DP_AC_q_8 }),
  .out1({ S1469 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_941_ (
  .in1({ S151, DP_AC_q_7 }),
  .out1({ S1470 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_942_ (
  .in1({ S1470, S1469 }),
  .out1({ S1471 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_943_ (
  .in1({ S1471, S137 }),
  .out1({ S1472 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_944_ (
  .in1({ S1472, S1468 }),
  .out1({ S1473 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1017_ (
  .in1({ S1473, S121 }),
  .out1({ S1474 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1018_ (
  .in1({ S1474, S1463 }),
  .out1({ S1476 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1019_ (
  .in1({ S1476, S1391 }),
  .out1({ S1477 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1020_ (
  .in1({ S151, S1312 }),
  .out1({ S1478 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1021_ (
  .in1({ S152, S1301 }),
  .out1({ S1479 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1022_ (
  .in1({ S1479, S1478 }),
  .out1({ S1480 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_945_ (
  .in1({ S152, DP_AC_q_12 }),
  .out1({ S1481 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_946_ (
  .in1({ S151, DP_AC_q_11 }),
  .out1({ S1482 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_947_ (
  .in1({ S1482, S1481 }),
  .out1({ S1483 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1023_ (
  .in1({ S1483, S136 }),
  .out1({ S1484 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_244_ (
  .in1({ S1484 }),
  .out1({ S1485 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_948_ (
  .in1({ S1480, S136 }),
  .out1({ S1487 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_949_ (
  .in1({ S1487, S1485 }),
  .out1({ S1488 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1024_ (
  .in1({ S1488, S122 }),
  .out1({ S1489 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_950_ (
  .in1({ S152, DP_AC_q_14 }),
  .out1({ S1490 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_951_ (
  .in1({ S151, DP_AC_q_13 }),
  .out1({ S1491 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_952_ (
  .in1({ S1491, S1490 }),
  .out1({ S1492 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_953_ (
  .in1({ S1492, S136 }),
  .out1({ S1493 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_245_ (
  .in1({ S1493 }),
  .out1({ S1494 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1025_ (
  .in1({ S152, DP_AC_q_15 }),
  .out1({ S1495 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1026_ (
  .in1({ S1495, S136 }),
  .out1({ S1496 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1027_ (
  .in1({ S1496, S1494 }),
  .out1({ S1498 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1028_ (
  .in1({ S1498, S121 }),
  .out1({ S1499 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1029_ (
  .in1({ S1499, S1489 }),
  .out1({ S1500 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_954_ (
  .in1({ S1500, S1408 }),
  .out1({ S1501 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_955_ (
  .in1({ S1389, DP_AC_q_1 }),
  .out1({ S1502 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_246_ (
  .in1({ S1502 }),
  .out1({ S1503 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1030_ (
  .in1({ S1503, S1436 }),
  .out1({ S1504 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_956_ (
  .in1({ S1504, S1501 }),
  .out1({ S1505 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1031_ (
  .in1({ S1505, S1477 }),
  .out1({ S1506 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_957_ (
  .in1({ S1436, S140 }),
  .out1({ S1507 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_958_ (
  .in1({ S1374, S2538[1] }),
  .out1({ S1509 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_959_ (
  .in1({ S1376, S1327 }),
  .out1({ S1510 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_960_ (
  .in1({ S1507, S1378 }),
  .out1({ S1511 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1032_ (
  .in1({ S1511, S1506 }),
  .out1({ S1512 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1033_ (
  .in1({ S1512, S1374 }),
  .out1({ S1513 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_961_ (
  .in1({ S1513, S1510 }),
  .out1({ S1514 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_962_ (
  .in1({ S1514, S1509 }),
  .out1({ S1515 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_963_ (
  .in1({ S1515, S1369 }),
  .out1({ S1516 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1034_ (
  .in1({ S1369, S1964 }),
  .out1({ S1517 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_964_ (
  .in1({ S1516, S1364 }),
  .out1({ S1518 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1035_ (
  .in1({ S1518, S1517 }),
  .out1({ S1520 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1036_ (
  .in1({ S1520, S1454 }),
  .out1({ S57 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1037_ (
  .in1({ S1367, DP_AC_q_2 }),
  .out1({ S1521 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_965_ (
  .in1({ S1400, S136 }),
  .out1({ S1522 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_966_ (
  .in1({ S1412, S137 }),
  .out1({ S1523 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_967_ (
  .in1({ S1523, S1522 }),
  .out1({ S1524 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_968_ (
  .in1({ S1524, S122 }),
  .out1({ S1525 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1038_ (
  .in1({ S1384, S137 }),
  .out1({ S1526 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1039_ (
  .in1({ S1395, S136 }),
  .out1({ S1527 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_247_ (
  .in1({ S1527 }),
  .out1({ S1528 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_969_ (
  .in1({ S1528, S121 }),
  .out1({ S1530 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1040_ (
  .in1({ S1530, S1526 }),
  .out1({ S1531 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1041_ (
  .in1({ S1531, S1391 }),
  .out1({ S1532 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_970_ (
  .in1({ S1532, S1525 }),
  .out1({ S1533 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_971_ (
  .in1({ S1416, S136 }),
  .out1({ S1534 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_248_ (
  .in1({ S1534 }),
  .out1({ S1535 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1042_ (
  .in1({ S1424, S136 }),
  .out1({ S1536 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1043_ (
  .in1({ S1536, S1535 }),
  .out1({ S1537 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1044_ (
  .in1({ S1537, S122 }),
  .out1({ S1538 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1045_ (
  .in1({ S1428, S137 }),
  .out1({ S1539 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1046_ (
  .in1({ S1539, S121 }),
  .out1({ S1541 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1047_ (
  .in1({ S1541, S1538 }),
  .out1({ S1542 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_249_ (
  .in1({ S1542 }),
  .out1({ S1543 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1048_ (
  .in1({ S1543, S1407 }),
  .out1({ S1544 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_972_ (
  .in1({ S1389, DP_AC_q_2 }),
  .out1({ S1545 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_973_ (
  .in1({ S1545, S1435 }),
  .out1({ S1546 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1049_ (
  .in1({ S1546, S1544 }),
  .out1({ S1547 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_974_ (
  .in1({ S1547, S1533 }),
  .out1({ S1548 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1050_ (
  .in1({ S1435, S125 }),
  .out1({ S1549 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_975_ (
  .in1({ S1376, S1319 }),
  .out1({ S1550 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1051_ (
  .in1({ S1549, S1376 }),
  .out1({ S1552 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_976_ (
  .in1({ S1552, S1548 }),
  .out1({ S1553 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_977_ (
  .in1({ S1553, S1550 }),
  .out1({ S1554 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_978_ (
  .in1({ S1554, S1375 }),
  .out1({ S1555 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1052_ (
  .in1({ S1375, S2538[2] }),
  .out1({ S1556 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1053_ (
  .in1({ S1556, S1370 }),
  .out1({ S1557 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_979_ (
  .in1({ S1557, S1555 }),
  .out1({ S1558 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_980_ (
  .in1({ S1370, S1972 }),
  .out1({ S1559 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_981_ (
  .in1({ S1559, S1558 }),
  .out1({ S1560 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1054_ (
  .in1({ S1560, S1365 }),
  .out1({ S1561 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1055_ (
  .in1({ S1561, S1521 }),
  .out1({ S58 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1056_ (
  .in1({ S1367, DP_AC_q_3 }),
  .out1({ S1563 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1057_ (
  .in1({ S1378, S1304 }),
  .out1({ S1564 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1058_ (
  .in1({ S1467, S136 }),
  .out1({ S1565 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1059_ (
  .in1({ S1460, S137 }),
  .out1({ S1566 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1060_ (
  .in1({ S1566, S1565 }),
  .out1({ S1567 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_982_ (
  .in1({ S1471, S136 }),
  .out1({ S1568 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_250_ (
  .in1({ S1568 }),
  .out1({ S1569 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1061_ (
  .in1({ S1480, S136 }),
  .out1({ S1570 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1062_ (
  .in1({ S1570, S1569 }),
  .out1({ S1571 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_983_ (
  .in1({ S1567, S121 }),
  .out1({ S1573 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1063_ (
  .in1({ S1571, S121 }),
  .out1({ S1574 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1064_ (
  .in1({ S1574, S1391 }),
  .out1({ S1575 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_984_ (
  .in1({ S1575, S1573 }),
  .out1({ S1576 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_985_ (
  .in1({ S1483, S136 }),
  .out1({ S1577 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_986_ (
  .in1({ S1492, S137 }),
  .out1({ S1578 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_987_ (
  .in1({ S1578, S1577 }),
  .out1({ S1579 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_988_ (
  .in1({ S1579, S121 }),
  .out1({ S1580 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_989_ (
  .in1({ S1495, S136 }),
  .out1({ S1581 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_990_ (
  .in1({ S1581, S122 }),
  .out1({ S1582 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_991_ (
  .in1({ S1582, S1580 }),
  .out1({ S1584 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1065_ (
  .in1({ S1584, S1407 }),
  .out1({ S1585 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1066_ (
  .in1({ S1390, S1224 }),
  .out1({ S1586 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1067_ (
  .in1({ S1586, S1585 }),
  .out1({ S1587 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_992_ (
  .in1({ S1587, S1576 }),
  .out1({ S1588 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_993_ (
  .in1({ S1588, S1435 }),
  .out1({ S1589 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1068_ (
  .in1({ S1435, S111 }),
  .out1({ S1590 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1069_ (
  .in1({ S1590, S1376 }),
  .out1({ S1591 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_994_ (
  .in1({ S1591, S1589 }),
  .out1({ S1592 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_995_ (
  .in1({ S1592, S1375 }),
  .out1({ S1593 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1070_ (
  .in1({ S1593, S1564 }),
  .out1({ S1595 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_996_ (
  .in1({ S1374, S1279 }),
  .out1({ S1596 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_997_ (
  .in1({ S1596, S1369 }),
  .out1({ S1597 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1071_ (
  .in1({ S1597, S1595 }),
  .out1({ S1598 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_998_ (
  .in1({ S1370, S1978 }),
  .out1({ S1599 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_999_ (
  .in1({ S1599, S1364 }),
  .out1({ S1600 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1072_ (
  .in1({ S1600, S1598 }),
  .out1({ S1601 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1073_ (
  .in1({ S1601, S1563 }),
  .out1({ S59 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1074_ (
  .in1({ S1367, DP_AC_q_4 }),
  .out1({ S1602 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1000_ (
  .in1({ S1418, S122 }),
  .out1({ S1603 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1075_ (
  .in1({ S1403, S122 }),
  .out1({ S1605 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1001_ (
  .in1({ S1603, S1392 }),
  .out1({ S1606 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1076_ (
  .in1({ S1606, S1605 }),
  .out1({ S1607 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1077_ (
  .in1({ S1430, S122 }),
  .out1({ S1608 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1002_ (
  .in1({ S1608, S1408 }),
  .out1({ S1609 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1078_ (
  .in1({ S1390, S1235 }),
  .out1({ S1610 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1079_ (
  .in1({ S1610, S1436 }),
  .out1({ S1611 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1003_ (
  .in1({ S1611, S1609 }),
  .out1({ S1612 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1080_ (
  .in1({ S1612, S1607 }),
  .out1({ S1613 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1004_ (
  .in1({ S1436, S95 }),
  .out1({ S1614 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1005_ (
  .in1({ S1614, S1378 }),
  .out1({ S1616 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1081_ (
  .in1({ S1616, S1613 }),
  .out1({ S1617 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1082_ (
  .in1({ S1378, S1294 }),
  .out1({ S1618 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1083_ (
  .in1({ S1618, S1617 }),
  .out1({ S1619 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1084_ (
  .in1({ S1619, S1374 }),
  .out1({ S1620 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1006_ (
  .in1({ S1374, S1377 }),
  .out1({ S1621 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1007_ (
  .in1({ S1621, S1369 }),
  .out1({ S1622 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1085_ (
  .in1({ S1622, S1620 }),
  .out1({ S1623 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1008_ (
  .in1({ S1370, S1990 }),
  .out1({ S1624 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1009_ (
  .in1({ S1624, S1364 }),
  .out1({ S1625 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1086_ (
  .in1({ S1625, S1623 }),
  .out1({ S1627 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1087_ (
  .in1({ S1627, S1602 }),
  .out1({ S60 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1088_ (
  .in1({ S1367, DP_AC_q_5 }),
  .out1({ S1628 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1089_ (
  .in1({ S1378, S1286 }),
  .out1({ S1629 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1090_ (
  .in1({ S1488, S121 }),
  .out1({ S1630 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1010_ (
  .in1({ S1473, S121 }),
  .out1({ S1631 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1091_ (
  .in1({ S1630, S1391 }),
  .out1({ S1632 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1011_ (
  .in1({ S1632, S1631 }),
  .out1({ S1633 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1012_ (
  .in1({ S1498, S121 }),
  .out1({ S1634 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1092_ (
  .in1({ S1634, S1407 }),
  .out1({ S1635 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1013_ (
  .in1({ S1389, DP_AC_q_5 }),
  .out1({ S1637 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1014_ (
  .in1({ S1637, S1435 }),
  .out1({ S1638 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1093_ (
  .in1({ S1638, S1635 }),
  .out1({ S1639 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1015_ (
  .in1({ S1639, S1633 }),
  .out1({ S1640 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1016_ (
  .in1({ S1436, S83 }),
  .out1({ S1641 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1017_ (
  .in1({ S1641, S1640 }),
  .out1({ S1642 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1018_ (
  .in1({ S1642, S1378 }),
  .out1({ S1643 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1019_ (
  .in1({ S1643, S1375 }),
  .out1({ S1644 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1094_ (
  .in1({ S1644, S1629 }),
  .out1({ S1645 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1095_ (
  .in1({ S1375, S2538[5] }),
  .out1({ S1646 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1096_ (
  .in1({ S1646, S1370 }),
  .out1({ S1648 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_251_ (
  .in1({ S1648 }),
  .out1({ S1649 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1097_ (
  .in1({ S1649, S1645 }),
  .out1({ S1650 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1020_ (
  .in1({ S1370, S1997 }),
  .out1({ S1651 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1021_ (
  .in1({ S1651, S1364 }),
  .out1({ S1652 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1098_ (
  .in1({ S1652, S1650 }),
  .out1({ S1653 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1099_ (
  .in1({ S1653, S1628 }),
  .out1({ S61 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1100_ (
  .in1({ S1367, DP_AC_q_6 }),
  .out1({ S1654 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1101_ (
  .in1({ S1378, S1276 }),
  .out1({ S1655 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1022_ (
  .in1({ S1524, S121 }),
  .out1({ S1656 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1102_ (
  .in1({ S1537, S121 }),
  .out1({ S1658 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1103_ (
  .in1({ S1658, S1391 }),
  .out1({ S1659 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1023_ (
  .in1({ S1659, S1656 }),
  .out1({ S1660 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1024_ (
  .in1({ S1539, S121 }),
  .out1({ S1661 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1104_ (
  .in1({ S1661, S1407 }),
  .out1({ S1662 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1025_ (
  .in1({ S1389, DP_AC_q_6 }),
  .out1({ S1663 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_252_ (
  .in1({ S1663 }),
  .out1({ S1664 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1105_ (
  .in1({ S1664, S1662 }),
  .out1({ S1665 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1026_ (
  .in1({ S1665, S1660 }),
  .out1({ S1666 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1027_ (
  .in1({ S1666, S1435 }),
  .out1({ S1667 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1028_ (
  .in1({ S1436, S2530 }),
  .out1({ S1669 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1106_ (
  .in1({ S1669, DP_AC_q_6 }),
  .out1({ S1670 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1107_ (
  .in1({ S1670, S1376 }),
  .out1({ S1671 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1029_ (
  .in1({ S1671, S1667 }),
  .out1({ S1672 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1030_ (
  .in1({ S1672, S1375 }),
  .out1({ S1673 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1108_ (
  .in1({ S1673, S1655 }),
  .out1({ S1674 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1109_ (
  .in1({ S1375, S2538[6] }),
  .out1({ S1675 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1110_ (
  .in1({ S1675, S1370 }),
  .out1({ S1676 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_253_ (
  .in1({ S1676 }),
  .out1({ S1677 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1111_ (
  .in1({ S1677, S1674 }),
  .out1({ S1678 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1031_ (
  .in1({ S1370, S2004 }),
  .out1({ S1680 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1032_ (
  .in1({ S1680, S1364 }),
  .out1({ S1681 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1112_ (
  .in1({ S1681, S1678 }),
  .out1({ S1682 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1113_ (
  .in1({ S1682, S1654 }),
  .out1({ S62 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1114_ (
  .in1({ S1367, DP_AC_q_7 }),
  .out1({ S1683 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1033_ (
  .in1({ S1376, S1269 }),
  .out1({ S1684 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1115_ (
  .in1({ S1571, S122 }),
  .out1({ S1685 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1034_ (
  .in1({ S1579, S122 }),
  .out1({ S1686 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1035_ (
  .in1({ S1686, S1392 }),
  .out1({ S1687 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1116_ (
  .in1({ S1687, S1685 }),
  .out1({ S1688 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1117_ (
  .in1({ S1581, S122 }),
  .out1({ S1690 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1036_ (
  .in1({ S1690, S1408 }),
  .out1({ S1691 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1037_ (
  .in1({ S1389, DP_AC_q_7 }),
  .out1({ S1692 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1038_ (
  .in1({ S1692, S1691 }),
  .out1({ S1693 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1118_ (
  .in1({ S1693, S1688 }),
  .out1({ S1694 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1119_ (
  .in1({ S1694, S1436 }),
  .out1({ S1695 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1039_ (
  .in1({ S1436, S2521 }),
  .out1({ S1696 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1040_ (
  .in1({ S1696, S1378 }),
  .out1({ S1697 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1120_ (
  .in1({ S1697, S1695 }),
  .out1({ S1698 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1041_ (
  .in1({ S1684, S1375 }),
  .out1({ S1699 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1121_ (
  .in1({ S1699, S1698 }),
  .out1({ S1701 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1122_ (
  .in1({ S1375, S2538[7] }),
  .out1({ S1702 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1123_ (
  .in1({ S1702, S1370 }),
  .out1({ S1703 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_254_ (
  .in1({ S1703 }),
  .out1({ S1704 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1124_ (
  .in1({ S1704, S1701 }),
  .out1({ S1705 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1042_ (
  .in1({ S1370, S2011 }),
  .out1({ S1706 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1043_ (
  .in1({ S1706, S1364 }),
  .out1({ S1707 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1125_ (
  .in1({ S1707, S1705 }),
  .out1({ S1708 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1126_ (
  .in1({ S1708, S1683 }),
  .out1({ S63 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1127_ (
  .in1({ S1367, DP_AC_q_8 }),
  .out1({ S1709 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1128_ (
  .in1({ S1378, S1261 }),
  .out1({ S1711 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1129_ (
  .in1({ S1433, S1391 }),
  .out1({ S1712 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1044_ (
  .in1({ S1389, DP_AC_q_8 }),
  .out1({ S1713 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_255_ (
  .in1({ S1713 }),
  .out1({ S1714 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1130_ (
  .in1({ S1714, S1712 }),
  .out1({ S1715 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1131_ (
  .in1({ S1715, S1436 }),
  .out1({ S1716 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1132_ (
  .in1({ S2506, DP_AC_q_8 }),
  .out1({ S1717 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1045_ (
  .in1({ S1717, S1436 }),
  .out1({ S1718 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1133_ (
  .in1({ S1716, S1376 }),
  .out1({ S1719 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1046_ (
  .in1({ S1719, S1718 }),
  .out1({ S1720 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1047_ (
  .in1({ S1720, S1375 }),
  .out1({ S1722 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1134_ (
  .in1({ S1722, S1711 }),
  .out1({ S1723 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1135_ (
  .in1({ S1375, S2538[8] }),
  .out1({ S1724 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1136_ (
  .in1({ S1724, S1370 }),
  .out1({ S1725 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_256_ (
  .in1({ S1725 }),
  .out1({ S1726 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1137_ (
  .in1({ S1726, S1723 }),
  .out1({ S1727 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1048_ (
  .in1({ S1370, S2018 }),
  .out1({ S1728 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1049_ (
  .in1({ S1728, S1364 }),
  .out1({ S1729 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1138_ (
  .in1({ S1729, S1727 }),
  .out1({ S1730 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1139_ (
  .in1({ S1730, S1709 }),
  .out1({ S64 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1140_ (
  .in1({ S1367, DP_AC_q_9 }),
  .out1({ S1732 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1050_ (
  .in1({ S1376, S1252 }),
  .out1({ S1733 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1051_ (
  .in1({ S1500, S1392 }),
  .out1({ S1734 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1052_ (
  .in1({ S1389, DP_AC_q_9 }),
  .out1({ S1735 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1053_ (
  .in1({ S1735, S1734 }),
  .out1({ S1736 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1054_ (
  .in1({ S1736, S1435 }),
  .out1({ S1737 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1055_ (
  .in1({ S1436, S1301 }),
  .out1({ S1738 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1141_ (
  .in1({ S1738, S2498 }),
  .out1({ S1739 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1056_ (
  .in1({ S1737, S1378 }),
  .out1({ S1740 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1142_ (
  .in1({ S1740, S1739 }),
  .out1({ S1741 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1143_ (
  .in1({ S1741, S1374 }),
  .out1({ S1742 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1057_ (
  .in1({ S1742, S1733 }),
  .out1({ S1743 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1144_ (
  .in1({ S1375, S2538[9] }),
  .out1({ S1744 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1145_ (
  .in1({ S1744, S1370 }),
  .out1({ S1745 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1058_ (
  .in1({ S1745, S1743 }),
  .out1({ S1746 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1059_ (
  .in1({ S1370, S2025 }),
  .out1({ S1747 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_257_ (
  .in1({ S1747 }),
  .out1({ S1748 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1060_ (
  .in1({ S1746, S1364 }),
  .out1({ S1749 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1146_ (
  .in1({ S1749, S1748 }),
  .out1({ S1750 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1147_ (
  .in1({ S1750, S1732 }),
  .out1({ S65 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1148_ (
  .in1({ S1367, DP_AC_q_10 }),
  .out1({ S1752 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1061_ (
  .in1({ S1376, S1242 }),
  .out1({ S1753 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1062_ (
  .in1({ S1542, S1392 }),
  .out1({ S1754 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1063_ (
  .in1({ S1389, DP_AC_q_10 }),
  .out1({ S1755 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1064_ (
  .in1({ S1755, S1754 }),
  .out1({ S1756 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1065_ (
  .in1({ S1756, S1435 }),
  .out1({ S1757 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1066_ (
  .in1({ S1436, S1312 }),
  .out1({ S1758 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1149_ (
  .in1({ S1758, S2489 }),
  .out1({ S1759 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1067_ (
  .in1({ S1757, S1378 }),
  .out1({ S1760 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1150_ (
  .in1({ S1760, S1759 }),
  .out1({ S1761 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1151_ (
  .in1({ S1761, S1374 }),
  .out1({ S1763 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1068_ (
  .in1({ S1763, S1753 }),
  .out1({ S1764 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1152_ (
  .in1({ S1375, S2538[10] }),
  .out1({ S1765 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1153_ (
  .in1({ S1765, S1370 }),
  .out1({ S1766 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1069_ (
  .in1({ S1766, S1764 }),
  .out1({ S1767 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1070_ (
  .in1({ S1370, S2032 }),
  .out1({ S1768 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_258_ (
  .in1({ S1768 }),
  .out1({ S1769 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1071_ (
  .in1({ S1767, S1364 }),
  .out1({ S1770 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1154_ (
  .in1({ S1770, S1769 }),
  .out1({ S1771 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1155_ (
  .in1({ S1771, S1752 }),
  .out1({ S66 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1156_ (
  .in1({ S1367, DP_AC_q_11 }),
  .out1({ S1773 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1072_ (
  .in1({ S1370, S2039 }),
  .out1({ S1774 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1073_ (
  .in1({ S1774, S1364 }),
  .out1({ S1775 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1074_ (
  .in1({ S1376, S1234 }),
  .out1({ S1776 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1157_ (
  .in1({ S1584, S1391 }),
  .out1({ S1777 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1075_ (
  .in1({ S1389, DP_AC_q_11 }),
  .out1({ S1778 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_259_ (
  .in1({ S1778 }),
  .out1({ S1779 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1158_ (
  .in1({ S1779, S1777 }),
  .out1({ S1780 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1159_ (
  .in1({ S1780, S1436 }),
  .out1({ S1781 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1160_ (
  .in1({ S2479, DP_AC_q_11 }),
  .out1({ S1782 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1076_ (
  .in1({ S1782, S1436 }),
  .out1({ S1784 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1077_ (
  .in1({ S1784, S1378 }),
  .out1({ S1785 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1161_ (
  .in1({ S1785, S1781 }),
  .out1({ S1786 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1162_ (
  .in1({ S1786, S1374 }),
  .out1({ S1787 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1078_ (
  .in1({ S1787, S1776 }),
  .out1({ S1788 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1163_ (
  .in1({ S1375, S2538[11] }),
  .out1({ S1789 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_260_ (
  .in1({ S1789 }),
  .out1({ S1790 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1079_ (
  .in1({ S1790, S1788 }),
  .out1({ S1791 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1164_ (
  .in1({ S1791, S1370 }),
  .out1({ S1792 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1165_ (
  .in1({ S1792, S1775 }),
  .out1({ S1793 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1166_ (
  .in1({ S1793, S1773 }),
  .out1({ S67 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1167_ (
  .in1({ S1367, DP_AC_q_12 }),
  .out1({ S1795 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1080_ (
  .in1({ S1376, S1221 }),
  .out1({ S1796 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1081_ (
  .in1({ S1608, S1392 }),
  .out1({ S1797 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1082_ (
  .in1({ S1389, DP_AC_q_12 }),
  .out1({ S1798 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1083_ (
  .in1({ S1798, S1797 }),
  .out1({ S1799 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_261_ (
  .in1({ S1799 }),
  .out1({ S1800 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1168_ (
  .in1({ S1800, S1436 }),
  .out1({ S1801 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1169_ (
  .in1({ S2470, DP_AC_q_12 }),
  .out1({ S1802 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1084_ (
  .in1({ S1802, S1436 }),
  .out1({ S1803 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1085_ (
  .in1({ S1803, S1378 }),
  .out1({ S1805 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1170_ (
  .in1({ S1805, S1801 }),
  .out1({ S1806 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1171_ (
  .in1({ S1806, S1374 }),
  .out1({ S1807 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1086_ (
  .in1({ S1807, S1796 }),
  .out1({ S1808 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1172_ (
  .in1({ S1375, S2538[12] }),
  .out1({ S1809 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_262_ (
  .in1({ S1809 }),
  .out1({ S1810 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1087_ (
  .in1({ S1810, S1808 }),
  .out1({ S1811 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1173_ (
  .in1({ S1811, S1370 }),
  .out1({ S1812 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1174_ (
  .in1({ S1812, S1775 }),
  .out1({ S1813 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1175_ (
  .in1({ S1813, S1795 }),
  .out1({ S68 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1176_ (
  .in1({ S1367, DP_AC_q_13 }),
  .out1({ S1815 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1088_ (
  .in1({ S1374, S2538[13] }),
  .out1({ S1816 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1089_ (
  .in1({ S1376, S1214 }),
  .out1({ S1817 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1177_ (
  .in1({ S1634, S1391 }),
  .out1({ S1818 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1090_ (
  .in1({ S1389, DP_AC_q_13 }),
  .out1({ S1819 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1091_ (
  .in1({ S1819, S1435 }),
  .out1({ S1820 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1178_ (
  .in1({ S1820, S1818 }),
  .out1({ S1821 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1092_ (
  .in1({ S1436, S2463 }),
  .out1({ S1822 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1093_ (
  .in1({ S1822, S1378 }),
  .out1({ S1823 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1179_ (
  .in1({ S1823, S1821 }),
  .out1({ S1824 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1180_ (
  .in1({ S1824, S1374 }),
  .out1({ S1826 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1094_ (
  .in1({ S1826, S1817 }),
  .out1({ S1827 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1095_ (
  .in1({ S1827, S1816 }),
  .out1({ S1828 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_263_ (
  .in1({ S1828 }),
  .out1({ S1829 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1181_ (
  .in1({ S1829, S1370 }),
  .out1({ S1830 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1182_ (
  .in1({ S1830, S1775 }),
  .out1({ S1831 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1183_ (
  .in1({ S1831, S1815 }),
  .out1({ S69 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1184_ (
  .in1({ S1367, DP_AC_q_14 }),
  .out1({ S1832 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1185_ (
  .in1({ S1375, S1508 }),
  .out1({ S1833 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1186_ (
  .in1({ S1378, S1204 }),
  .out1({ S1834 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1187_ (
  .in1({ S1661, S1391 }),
  .out1({ S1836 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1096_ (
  .in1({ S1389, DP_AC_q_14 }),
  .out1({ S1837 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1097_ (
  .in1({ S1837, S1435 }),
  .out1({ S1838 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1188_ (
  .in1({ S1838, S1836 }),
  .out1({ S1839 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1098_ (
  .in1({ S1436, S2453 }),
  .out1({ S1840 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1189_ (
  .in1({ S1839, S1376 }),
  .out1({ S1841 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1099_ (
  .in1({ S1841, S1840 }),
  .out1({ S1842 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1100_ (
  .in1({ S1842, S1375 }),
  .out1({ S1843 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1190_ (
  .in1({ S1843, S1834 }),
  .out1({ S1844 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1191_ (
  .in1({ S1844, S1833 }),
  .out1({ S1845 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1192_ (
  .in1({ S1845, S1370 }),
  .out1({ S1847 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1193_ (
  .in1({ S1847, S1775 }),
  .out1({ S1848 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1194_ (
  .in1({ S1848, S1832 }),
  .out1({ S70 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1195_ (
  .in1({ S1367, DP_AC_q_15 }),
  .out1({ S1849 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1196_ (
  .in1({ S1378, S979 }),
  .out1({ S1850 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1101_ (
  .in1({ S1690, S1392 }),
  .out1({ S1851 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1102_ (
  .in1({ S1389, DP_AC_q_15 }),
  .out1({ S1852 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1103_ (
  .in1({ S1852, S1851 }),
  .out1({ S1853 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1104_ (
  .in1({ S1853, S1435 }),
  .out1({ S1854 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1105_ (
  .in1({ S1436, S1356 }),
  .out1({ S1855 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1197_ (
  .in1({ S1855, S2444 }),
  .out1({ S1857 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1198_ (
  .in1({ S1857, S1376 }),
  .out1({ S1858 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1106_ (
  .in1({ S1858, S1854 }),
  .out1({ S1859 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1107_ (
  .in1({ S1859, S1375 }),
  .out1({ S1860 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1199_ (
  .in1({ S1860, S1850 }),
  .out1({ S1861 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1200_ (
  .in1({ S1375, S2538[15] }),
  .out1({ S1862 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1201_ (
  .in1({ S1862, S1370 }),
  .out1({ S1863 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_264_ (
  .in1({ S1863 }),
  .out1({ S1864 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_1_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S0 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IMM1_in1_0 }),
  .Si({ S2543 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_2_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S1 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IMM1_in1_1 }),
  .Si({ S2596 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_3_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S2 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IMM1_in1_2 }),
  .Si({ S2597 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_4_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S3 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IMM1_in1_3 }),
  .Si({ S2595 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_5_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S4 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_q_0 }),
  .Si({ S2544 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_6_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S5 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_q_1 }),
  .Si({ S2593 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_7_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S6 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_q_2 }),
  .Si({ S2594 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_8_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S7 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_q_3 }),
  .Si({ S2591 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_9_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S8 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_q_4 }),
  .Si({ S2592 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_10_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S9 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_q_5 }),
  .Si({ S2590 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_11_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S10 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_q_6 }),
  .Si({ S2589 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_12_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S11 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_q_7 }),
  .Si({ S2588 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_13_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S12 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_q_8 }),
  .Si({ S2586 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_14_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S13 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_q_9 }),
  .Si({ S2587 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_15_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S14 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_q_10 }),
  .Si({ S2585 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_16_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S15 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_q_11 }),
  .Si({ S2583 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_17_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S16 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_q_12 }),
  .Si({ S2584 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_18_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S17 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_q_13 }),
  .Si({ S2581 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_19_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S18 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_q_14 }),
  .Si({ S2582 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_20_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S19 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_q_15 }),
  .Si({ S2580 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_21_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S20 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_SR_N_q }),
  .Si({ S2545 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_22_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S21 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_0 }),
  .Si({ S2546 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_23_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S22 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_1 }),
  .Si({ S2578 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_24_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S23 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_2 }),
  .Si({ S2579 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_25_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S24 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_3 }),
  .Si({ S2576 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_26_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S25 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_4 }),
  .Si({ S2577 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_27_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S26 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_5 }),
  .Si({ S2575 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_28_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S27 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_6 }),
  .Si({ S2574 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_29_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S28 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_7 }),
  .Si({ S2572 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_30_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S29 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_8 }),
  .Si({ S2573 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_31_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S30 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_9 }),
  .Si({ S2571 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_32_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S31 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_10 }),
  .Si({ S2569 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_33_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S32 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_11 }),
  .Si({ S2570 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_34_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S33 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_12 }),
  .Si({ S2567 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_35_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S34 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_13 }),
  .Si({ S2568 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_36_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S35 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_14 }),
  .Si({ S2566 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_37_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S36 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_15 }),
  .Si({ S2564 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_38_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S37 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_SR_C_q }),
  .Si({ S2547 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_39_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S38 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_SR_V_q }),
  .Si({ S2548 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_40_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S39 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_0 }),
  .Si({ S2549 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_41_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S40 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_1 }),
  .Si({ S2565 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_42_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S41 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_2 }),
  .Si({ S2562 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_43_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S42 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_3 }),
  .Si({ S2563 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_44_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S43 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_4 }),
  .Si({ S2561 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_45_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S44 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_5 }),
  .Si({ S2559 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_46_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S45 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_6 }),
  .Si({ S2560 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_47_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S46 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_7 }),
  .Si({ S2557 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_48_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S47 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_8 }),
  .Si({ S2558 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_49_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S48 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_9 }),
  .Si({ S2556 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_50_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S49 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_10 }),
  .Si({ S2554 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_51_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S50 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_11 }),
  .Si({ S2555 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_52_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S51 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_12 }),
  .Si({ S2553 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_53_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S52 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_13 }),
  .Si({ S2552 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_54_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S53 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_14 }),
  .Si({ S2551 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_55_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S54 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_15 }),
  .Si({ S2550 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_56_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S55 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_SR_Z_q }),
  .Si({ S2614 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_57_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S56 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_q_0 }),
  .Si({ S2615 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_58_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S57 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_q_1 }),
  .Si({ S2599 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_59_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S58 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_q_2 }),
  .Si({ S2600 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_60_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S59 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_q_3 }),
  .Si({ S2601 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_61_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S60 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_q_4 }),
  .Si({ S2602 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_62_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S61 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_q_5 }),
  .Si({ S2603 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_63_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S62 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_q_6 }),
  .Si({ S2604 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_64_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S63 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_q_7 }),
  .Si({ S2605 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_65_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S64 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_q_8 }),
  .Si({ S2606 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_66_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S65 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_q_9 }),
  .Si({ S2607 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_67_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S66 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_q_10 }),
  .Si({ S2608 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_68_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S67 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_q_11 }),
  .Si({ S2609 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_69_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S68 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_q_12 }),
  .Si({ S2610 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_70_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S69 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_q_13 }),
  .Si({ S2611 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_71_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S70 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_q_14 }),
  .Si({ S2612 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_72_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ S71 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_q_15 }),
  .Si({ S2613 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_73_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ CU_nstate_0 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_pstate_0 }),
  .Si({ S2616 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_74_ (
  .C({ S2537 }),
  .CE({ 1'b1 }),
  .CLR({ S2541 }),
  .D({ CU_nstate_1 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_pstate_1 }),
  .Si({ S2598 }),
  .global_reset({ 1'b0 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_1_ (
  .in1({ S2536[0] }),
  .out1({ addrBus[0] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_2_ (
  .in1({ S2536[1] }),
  .out1({ addrBus[1] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_3_ (
  .in1({ S2536[10] }),
  .out1({ addrBus[10] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_4_ (
  .in1({ S2536[11] }),
  .out1({ addrBus[11] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_5_ (
  .in1({ S2536[12] }),
  .out1({ addrBus[12] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_6_ (
  .in1({ S2536[13] }),
  .out1({ addrBus[13] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_7_ (
  .in1({ S2536[14] }),
  .out1({ addrBus[14] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_8_ (
  .in1({ S2536[15] }),
  .out1({ addrBus[15] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_9_ (
  .in1({ S2536[2] }),
  .out1({ addrBus[2] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_10_ (
  .in1({ S2536[3] }),
  .out1({ addrBus[3] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_11_ (
  .in1({ S2536[4] }),
  .out1({ addrBus[4] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_12_ (
  .in1({ S2536[5] }),
  .out1({ addrBus[5] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_13_ (
  .in1({ S2536[6] }),
  .out1({ addrBus[6] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_14_ (
  .in1({ S2536[7] }),
  .out1({ addrBus[7] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_15_ (
  .in1({ S2536[8] }),
  .out1({ addrBus[8] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_16_ (
  .in1({ S2536[9] }),
  .out1({ addrBus[9] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_17_ (
  .in1({ clk }),
  .out1({ S2537 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_18_ (
  .in1({ dataBus_in[0] }),
  .out1({ S2538[0] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_19_ (
  .in1({ dataBus_in[1] }),
  .out1({ S2538[1] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_20_ (
  .in1({ dataBus_in[10] }),
  .out1({ S2538[10] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_21_ (
  .in1({ dataBus_in[11] }),
  .out1({ S2538[11] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_22_ (
  .in1({ dataBus_in[12] }),
  .out1({ S2538[12] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_23_ (
  .in1({ dataBus_in[13] }),
  .out1({ S2538[13] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_24_ (
  .in1({ dataBus_in[14] }),
  .out1({ S2538[14] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_25_ (
  .in1({ dataBus_in[15] }),
  .out1({ S2538[15] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_26_ (
  .in1({ dataBus_in[2] }),
  .out1({ S2538[2] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_27_ (
  .in1({ dataBus_in[3] }),
  .out1({ S2538[3] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_28_ (
  .in1({ dataBus_in[4] }),
  .out1({ S2538[4] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_29_ (
  .in1({ dataBus_in[5] }),
  .out1({ S2538[5] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_30_ (
  .in1({ dataBus_in[6] }),
  .out1({ S2538[6] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_31_ (
  .in1({ dataBus_in[7] }),
  .out1({ S2538[7] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_32_ (
  .in1({ dataBus_in[8] }),
  .out1({ S2538[8] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_33_ (
  .in1({ dataBus_in[9] }),
  .out1({ S2538[9] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_34_ (
  .in1({ S2539[0] }),
  .out1({ dataBus_out[0] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_35_ (
  .in1({ S2539[1] }),
  .out1({ dataBus_out[1] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_36_ (
  .in1({ S2539[10] }),
  .out1({ dataBus_out[10] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_37_ (
  .in1({ S2539[11] }),
  .out1({ dataBus_out[11] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_38_ (
  .in1({ S2539[12] }),
  .out1({ dataBus_out[12] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_39_ (
  .in1({ S2539[13] }),
  .out1({ dataBus_out[13] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_40_ (
  .in1({ S2539[14] }),
  .out1({ dataBus_out[14] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_41_ (
  .in1({ S2539[15] }),
  .out1({ dataBus_out[15] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_42_ (
  .in1({ S2539[2] }),
  .out1({ dataBus_out[2] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_43_ (
  .in1({ S2539[3] }),
  .out1({ dataBus_out[3] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_44_ (
  .in1({ S2539[4] }),
  .out1({ dataBus_out[4] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_45_ (
  .in1({ S2539[5] }),
  .out1({ dataBus_out[5] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_46_ (
  .in1({ S2539[6] }),
  .out1({ dataBus_out[6] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_47_ (
  .in1({ S2539[7] }),
  .out1({ dataBus_out[7] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_48_ (
  .in1({ S2539[8] }),
  .out1({ dataBus_out[8] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_49_ (
  .in1({ S2539[9] }),
  .out1({ dataBus_out[9] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_50_ (
  .in1({ S2540 }),
  .out1({ readMEM })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_51_ (
  .in1({ rst }),
  .out1({ S2541 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_52_ (
  .in1({ S2542 }),
  .out1({ writeMEM })
);

endmodule