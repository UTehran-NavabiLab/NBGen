module Circuit432(in4, in17, in30, in43, in56, in69, in82, in95, in108, in1, in11, in24, in37, in50, in63, in76, in89, in102, in8, in21, in34, in47, in60, in73, in86, in99, in112, in14, in27, in40, in53, in66, in79, in92, in105, in115, out223, out329, out370, out421, out430, out431, out432);

wire Ckt432_I_0;
wire Ckt432_I_1;
wire Ckt432_I_2;
wire Ckt432_I_3;
wire Ckt432_I_4;
wire Ckt432_I_5;
wire Ckt432_I_6;
wire Ckt432_I_7;
wire Ckt432_I_8;
wire Ckt432_M1_X1_0;
wire Ckt432_M1_X1_1;
wire Ckt432_M1_X1_2;
wire Ckt432_M1_X1_3;
wire Ckt432_M1_X1_4;
wire Ckt432_M1_X1_5;
wire Ckt432_M1_X1_6;
wire Ckt432_M1_X1_7;
wire Ckt432_M1_X1_8;
wire Ckt432_M1_n1;
wire Ckt432_M1_n10;
wire Ckt432_M1_n11;
wire Ckt432_M1_n12;
wire Ckt432_M1_n13;
wire Ckt432_M1_n14;
wire Ckt432_M1_n15;
wire Ckt432_M1_n2;
wire Ckt432_M1_n3;
wire Ckt432_M1_n4;
wire Ckt432_M1_n5;
wire Ckt432_M1_n6;
wire Ckt432_M1_n7;
wire Ckt432_M1_n8;
wire Ckt432_M1_n9;
wire Ckt432_M2_X2_0;
wire Ckt432_M2_X2_1;
wire Ckt432_M2_X2_2;
wire Ckt432_M2_X2_3;
wire Ckt432_M2_X2_4;
wire Ckt432_M2_X2_5;
wire Ckt432_M2_X2_6;
wire Ckt432_M2_X2_7;
wire Ckt432_M2_X2_8;
wire Ckt432_M2_n1;
wire Ckt432_M2_n10;
wire Ckt432_M2_n11;
wire Ckt432_M2_n12;
wire Ckt432_M2_n13;
wire Ckt432_M2_n14;
wire Ckt432_M2_n15;
wire Ckt432_M2_n16;
wire Ckt432_M2_n17;
wire Ckt432_M2_n18;
wire Ckt432_M2_n19;
wire Ckt432_M2_n2;
wire Ckt432_M2_n20;
wire Ckt432_M2_n3;
wire Ckt432_M2_n4;
wire Ckt432_M2_n5;
wire Ckt432_M2_n6;
wire Ckt432_M2_n7;
wire Ckt432_M2_n8;
wire Ckt432_M2_n9;
wire Ckt432_M3_n1;
wire Ckt432_M3_n10;
wire Ckt432_M3_n11;
wire Ckt432_M3_n12;
wire Ckt432_M3_n13;
wire Ckt432_M3_n14;
wire Ckt432_M3_n15;
wire Ckt432_M3_n16;
wire Ckt432_M3_n17;
wire Ckt432_M3_n18;
wire Ckt432_M3_n19;
wire Ckt432_M3_n2;
wire Ckt432_M3_n20;
wire Ckt432_M3_n3;
wire Ckt432_M3_n4;
wire Ckt432_M3_n5;
wire Ckt432_M3_n6;
wire Ckt432_M3_n7;
wire Ckt432_M3_n8;
wire Ckt432_M3_n9;
wire Ckt432_M4_n1;
wire Ckt432_M4_n10;
wire Ckt432_M4_n11;
wire Ckt432_M4_n12;
wire Ckt432_M4_n13;
wire Ckt432_M4_n14;
wire Ckt432_M4_n15;
wire Ckt432_M4_n16;
wire Ckt432_M4_n17;
wire Ckt432_M4_n18;
wire Ckt432_M4_n2;
wire Ckt432_M4_n3;
wire Ckt432_M4_n4;
wire Ckt432_M4_n5;
wire Ckt432_M4_n6;
wire Ckt432_M4_n7;
wire Ckt432_M4_n8;
wire Ckt432_M4_n9;
wire Ckt432_M5_n1;
wire Ckt432_M5_n2;
wire Ckt432_M5_n3;
wire Ckt432_M5_n4;
wire Ckt432_M5_n5;
wire Ckt432_M5_n6;
wire Ckt432_M5_n7;
wire Ckt432_M5_n8;
wire Ckt432_M5_n9;
input in4;
input in17;
input in30;
input in43;
input in56;
input in69;
input in82;
input in95;
input in108;
input in1;
input in11;
input in24;
input in37;
input in50;
input in63;
input in76;
input in89;
input in102;
input in8;
input in21;
input in34;
input in47;
input in60;
input in73;
input in86;
input in99;
input in112;
input in14;
input in27;
input in40;
input in53;
input in66;
input in79;
input in92;
input in105;
input in115;
output out223;
output out329;
output out370;
output out421;
output out430;
output out431;
output out432;

OAI21_X1 #() 
OAI21_X1_1_ (
  .A({ out223 }),
  .B1({ in1 }),
  .B2({ Ckt432_M1_n1 }),
  .ZN({ Ckt432_M1_X1_8 })
);
OR2_X1 #() 
OR2_X1_1_ (
  .A1({ Ckt432_M1_n10 }),
  .A2({ Ckt432_M1_n11 }),
  .ZN({ out223 })
);
OAI221_X1 #() 
OAI221_X1_1_ (
  .A({ Ckt432_M1_n12 }),
  .B1({ Ckt432_M1_n6 }),
  .B2({ in63 }),
  .C1({ Ckt432_M1_n5 }),
  .C2({ in50 }),
  .ZN({ Ckt432_M1_n11 })
);
INV_X1 #() 
INV_X1_1_ (
  .A({ Ckt432_M1_n13 }),
  .ZN({ Ckt432_M1_n12 })
);
OAI222_X1 #() 
OAI222_X1_1_ (
  .A1({ in89 }),
  .A2({ Ckt432_M1_n8 }),
  .B1({ in102 }),
  .B2({ Ckt432_M1_n9 }),
  .C1({ in76 }),
  .C2({ Ckt432_M1_n7 }),
  .ZN({ Ckt432_M1_n13 })
);
INV_X1 #() 
INV_X1_2_ (
  .A({ in82 }),
  .ZN({ Ckt432_M1_n7 })
);
INV_X1 #() 
INV_X1_3_ (
  .A({ in108 }),
  .ZN({ Ckt432_M1_n9 })
);
INV_X1 #() 
INV_X1_4_ (
  .A({ in95 }),
  .ZN({ Ckt432_M1_n8 })
);
INV_X1 #() 
INV_X1_5_ (
  .A({ in56 }),
  .ZN({ Ckt432_M1_n5 })
);
INV_X1 #() 
INV_X1_6_ (
  .A({ in69 }),
  .ZN({ Ckt432_M1_n6 })
);
OAI221_X1 #() 
OAI221_X1_2_ (
  .A({ Ckt432_M1_n14 }),
  .B1({ Ckt432_M1_n2 }),
  .B2({ in11 }),
  .C1({ Ckt432_M1_n1 }),
  .C2({ in1 }),
  .ZN({ Ckt432_M1_n10 })
);
OAI21_X1 #() 
OAI21_X1_2_ (
  .A({ out223 }),
  .B1({ in11 }),
  .B2({ Ckt432_M1_n2 }),
  .ZN({ Ckt432_M1_X1_7 })
);
INV_X1 #() 
INV_X1_7_ (
  .A({ Ckt432_M1_n15 }),
  .ZN({ Ckt432_M1_n14 })
);
OAI22_X1 #() 
OAI22_X1_1_ (
  .A1({ in24 }),
  .A2({ Ckt432_M1_n3 }),
  .B1({ in37 }),
  .B2({ Ckt432_M1_n4 }),
  .ZN({ Ckt432_M1_n15 })
);
INV_X1 #() 
INV_X1_8_ (
  .A({ in43 }),
  .ZN({ Ckt432_M1_n4 })
);
INV_X1 #() 
INV_X1_9_ (
  .A({ in30 }),
  .ZN({ Ckt432_M1_n3 })
);
INV_X1 #() 
INV_X1_10_ (
  .A({ in4 }),
  .ZN({ Ckt432_M1_n1 })
);
INV_X1 #() 
INV_X1_11_ (
  .A({ in17 }),
  .ZN({ Ckt432_M1_n2 })
);
OAI21_X1 #() 
OAI21_X1_3_ (
  .A({ out223 }),
  .B1({ in24 }),
  .B2({ Ckt432_M1_n3 }),
  .ZN({ Ckt432_M1_X1_6 })
);
OAI21_X1 #() 
OAI21_X1_4_ (
  .A({ out223 }),
  .B1({ in37 }),
  .B2({ Ckt432_M1_n4 }),
  .ZN({ Ckt432_M1_X1_5 })
);
OAI21_X1 #() 
OAI21_X1_5_ (
  .A({ out223 }),
  .B1({ in50 }),
  .B2({ Ckt432_M1_n5 }),
  .ZN({ Ckt432_M1_X1_4 })
);
OAI21_X1 #() 
OAI21_X1_6_ (
  .A({ out223 }),
  .B1({ in63 }),
  .B2({ Ckt432_M1_n6 }),
  .ZN({ Ckt432_M1_X1_3 })
);
OAI21_X1 #() 
OAI21_X1_7_ (
  .A({ out223 }),
  .B1({ in76 }),
  .B2({ Ckt432_M1_n7 }),
  .ZN({ Ckt432_M1_X1_2 })
);
OAI21_X1 #() 
OAI21_X1_8_ (
  .A({ out223 }),
  .B1({ in89 }),
  .B2({ Ckt432_M1_n8 }),
  .ZN({ Ckt432_M1_X1_1 })
);
OAI21_X1 #() 
OAI21_X1_9_ (
  .A({ out223 }),
  .B1({ in102 }),
  .B2({ Ckt432_M1_n9 }),
  .ZN({ Ckt432_M1_X1_0 })
);
NAND2_X1 #() 
NAND2_X1_1_ (
  .A1({ out329 }),
  .A2({ Ckt432_M2_n1 }),
  .ZN({ Ckt432_M2_X2_8 })
);
NAND4_X1 #() 
NAND4_X1_1_ (
  .A1({ Ckt432_M2_n5 }),
  .A2({ Ckt432_M2_n4 }),
  .A3({ Ckt432_M2_n10 }),
  .A4({ Ckt432_M2_n11 }),
  .ZN({ out329 })
);
AND4_X1 #() 
AND4_X1_1_ (
  .A1({ Ckt432_M2_n6 }),
  .A2({ Ckt432_M2_n7 }),
  .A3({ Ckt432_M2_n8 }),
  .A4({ Ckt432_M2_n9 }),
  .ZN({ Ckt432_M2_n11 })
);
NAND3_X1 #() 
NAND3_X1_1_ (
  .A1({ in108 }),
  .A2({ Ckt432_M2_n12 }),
  .A3({ Ckt432_M1_X1_0 }),
  .ZN({ Ckt432_M2_n9 })
);
INV_X1 #() 
INV_X1_12_ (
  .A({ in112 }),
  .ZN({ Ckt432_M2_n12 })
);
NAND3_X1 #() 
NAND3_X1_2_ (
  .A1({ in95 }),
  .A2({ Ckt432_M2_n13 }),
  .A3({ Ckt432_M1_X1_1 }),
  .ZN({ Ckt432_M2_n8 })
);
INV_X1 #() 
INV_X1_13_ (
  .A({ in99 }),
  .ZN({ Ckt432_M2_n13 })
);
NAND3_X1 #() 
NAND3_X1_3_ (
  .A1({ in82 }),
  .A2({ Ckt432_M2_n14 }),
  .A3({ Ckt432_M1_X1_2 }),
  .ZN({ Ckt432_M2_n7 })
);
INV_X1 #() 
INV_X1_14_ (
  .A({ in86 }),
  .ZN({ Ckt432_M2_n14 })
);
NAND3_X1 #() 
NAND3_X1_4_ (
  .A1({ in69 }),
  .A2({ Ckt432_M2_n15 }),
  .A3({ Ckt432_M1_X1_3 }),
  .ZN({ Ckt432_M2_n6 })
);
INV_X1 #() 
INV_X1_15_ (
  .A({ in73 }),
  .ZN({ Ckt432_M2_n15 })
);
NAND2_X1 #() 
NAND2_X1_2_ (
  .A1({ out329 }),
  .A2({ Ckt432_M2_n2 }),
  .ZN({ Ckt432_M2_X2_7 })
);
AND3_X1 #() 
AND3_X1_1_ (
  .A1({ Ckt432_M2_n3 }),
  .A2({ Ckt432_M2_n1 }),
  .A3({ Ckt432_M2_n2 }),
  .ZN({ Ckt432_M2_n10 })
);
NAND3_X1 #() 
NAND3_X1_5_ (
  .A1({ in17 }),
  .A2({ Ckt432_M2_n16 }),
  .A3({ Ckt432_M1_X1_7 }),
  .ZN({ Ckt432_M2_n2 })
);
INV_X1 #() 
INV_X1_16_ (
  .A({ in21 }),
  .ZN({ Ckt432_M2_n16 })
);
NAND3_X1 #() 
NAND3_X1_6_ (
  .A1({ in4 }),
  .A2({ Ckt432_M2_n17 }),
  .A3({ Ckt432_M1_X1_8 }),
  .ZN({ Ckt432_M2_n1 })
);
INV_X1 #() 
INV_X1_17_ (
  .A({ in8 }),
  .ZN({ Ckt432_M2_n17 })
);
NAND3_X1 #() 
NAND3_X1_7_ (
  .A1({ in30 }),
  .A2({ Ckt432_M2_n18 }),
  .A3({ Ckt432_M1_X1_6 }),
  .ZN({ Ckt432_M2_n3 })
);
INV_X1 #() 
INV_X1_18_ (
  .A({ in34 }),
  .ZN({ Ckt432_M2_n18 })
);
NAND3_X1 #() 
NAND3_X1_8_ (
  .A1({ in43 }),
  .A2({ Ckt432_M2_n19 }),
  .A3({ Ckt432_M1_X1_5 }),
  .ZN({ Ckt432_M2_n4 })
);
INV_X1 #() 
INV_X1_19_ (
  .A({ in47 }),
  .ZN({ Ckt432_M2_n19 })
);
NAND3_X1 #() 
NAND3_X1_9_ (
  .A1({ in56 }),
  .A2({ Ckt432_M2_n20 }),
  .A3({ Ckt432_M1_X1_4 }),
  .ZN({ Ckt432_M2_n5 })
);
NAND2_X1 #() 
NAND2_X1_3_ (
  .A1({ out329 }),
  .A2({ Ckt432_M2_n3 }),
  .ZN({ Ckt432_M2_X2_6 })
);
INV_X1 #() 
INV_X1_20_ (
  .A({ in60 }),
  .ZN({ Ckt432_M2_n20 })
);
NAND2_X1 #() 
NAND2_X1_4_ (
  .A1({ out329 }),
  .A2({ Ckt432_M2_n4 }),
  .ZN({ Ckt432_M2_X2_5 })
);
NAND2_X1 #() 
NAND2_X1_5_ (
  .A1({ out329 }),
  .A2({ Ckt432_M2_n5 }),
  .ZN({ Ckt432_M2_X2_4 })
);
NAND2_X1 #() 
NAND2_X1_6_ (
  .A1({ out329 }),
  .A2({ Ckt432_M2_n6 }),
  .ZN({ Ckt432_M2_X2_3 })
);
NAND2_X1 #() 
NAND2_X1_7_ (
  .A1({ out329 }),
  .A2({ Ckt432_M2_n7 }),
  .ZN({ Ckt432_M2_X2_2 })
);
NAND2_X1 #() 
NAND2_X1_8_ (
  .A1({ out329 }),
  .A2({ Ckt432_M2_n8 }),
  .ZN({ Ckt432_M2_X2_1 })
);
NAND2_X1 #() 
NAND2_X1_9_ (
  .A1({ out329 }),
  .A2({ Ckt432_M2_n9 }),
  .ZN({ Ckt432_M2_X2_0 })
);
NAND4_X1 #() 
NAND4_X1_2_ (
  .A1({ Ckt432_M3_n1 }),
  .A2({ Ckt432_M3_n2 }),
  .A3({ Ckt432_M3_n3 }),
  .A4({ Ckt432_M3_n4 }),
  .ZN({ out370 })
);
INV_X1 #() 
INV_X1_21_ (
  .A({ in14 }),
  .ZN({ Ckt432_M3_n12 })
);
AND3_X1 #() 
AND3_X1_2_ (
  .A1({ Ckt432_M3_n13 }),
  .A2({ Ckt432_M3_n14 }),
  .A3({ Ckt432_M3_n15 }),
  .ZN({ Ckt432_M3_n3 })
);
NAND4_X1 #() 
NAND4_X1_3_ (
  .A1({ Ckt432_M2_X2_2 }),
  .A2({ Ckt432_M1_X1_2 }),
  .A3({ in82 }),
  .A4({ Ckt432_M3_n16 }),
  .ZN({ Ckt432_M3_n15 })
);
INV_X1 #() 
INV_X1_22_ (
  .A({ in92 }),
  .ZN({ Ckt432_M3_n16 })
);
NAND4_X1 #() 
NAND4_X1_4_ (
  .A1({ Ckt432_M2_X2_0 }),
  .A2({ Ckt432_M1_X1_0 }),
  .A3({ in108 }),
  .A4({ Ckt432_M3_n17 }),
  .ZN({ Ckt432_M3_n14 })
);
INV_X1 #() 
INV_X1_23_ (
  .A({ in115 }),
  .ZN({ Ckt432_M3_n17 })
);
NAND4_X1 #() 
NAND4_X1_5_ (
  .A1({ Ckt432_M2_X2_1 }),
  .A2({ Ckt432_M1_X1_1 }),
  .A3({ in95 }),
  .A4({ Ckt432_M3_n18 }),
  .ZN({ Ckt432_M3_n13 })
);
INV_X1 #() 
INV_X1_24_ (
  .A({ in105 }),
  .ZN({ Ckt432_M3_n18 })
);
NAND4_X1 #() 
NAND4_X1_6_ (
  .A1({ Ckt432_M2_X2_3 }),
  .A2({ Ckt432_M1_X1_3 }),
  .A3({ in69 }),
  .A4({ Ckt432_M3_n19 }),
  .ZN({ Ckt432_M3_n2 })
);
INV_X1 #() 
INV_X1_25_ (
  .A({ in79 }),
  .ZN({ Ckt432_M3_n19 })
);
AND4_X1 #() 
AND4_X1_2_ (
  .A1({ Ckt432_M3_n5 }),
  .A2({ Ckt432_M3_n6 }),
  .A3({ Ckt432_M3_n7 }),
  .A4({ Ckt432_M3_n8 }),
  .ZN({ Ckt432_M3_n4 })
);
NAND4_X1 #() 
NAND4_X1_7_ (
  .A1({ Ckt432_M2_X2_4 }),
  .A2({ Ckt432_M1_X1_4 }),
  .A3({ in56 }),
  .A4({ Ckt432_M3_n20 }),
  .ZN({ Ckt432_M3_n1 })
);
INV_X1 #() 
INV_X1_26_ (
  .A({ in66 }),
  .ZN({ Ckt432_M3_n20 })
);
NAND4_X1 #() 
NAND4_X1_8_ (
  .A1({ Ckt432_M2_X2_5 }),
  .A2({ Ckt432_M1_X1_5 }),
  .A3({ in43 }),
  .A4({ Ckt432_M3_n9 }),
  .ZN({ Ckt432_M3_n8 })
);
INV_X1 #() 
INV_X1_27_ (
  .A({ in53 }),
  .ZN({ Ckt432_M3_n9 })
);
NAND4_X1 #() 
NAND4_X1_9_ (
  .A1({ Ckt432_M2_X2_6 }),
  .A2({ Ckt432_M1_X1_6 }),
  .A3({ in30 }),
  .A4({ Ckt432_M3_n10 }),
  .ZN({ Ckt432_M3_n7 })
);
INV_X1 #() 
INV_X1_28_ (
  .A({ in40 }),
  .ZN({ Ckt432_M3_n10 })
);
NAND4_X1 #() 
NAND4_X1_10_ (
  .A1({ Ckt432_M2_X2_7 }),
  .A2({ Ckt432_M1_X1_7 }),
  .A3({ in17 }),
  .A4({ Ckt432_M3_n11 }),
  .ZN({ Ckt432_M3_n6 })
);
INV_X1 #() 
INV_X1_29_ (
  .A({ in27 }),
  .ZN({ Ckt432_M3_n11 })
);
NAND4_X1 #() 
NAND4_X1_11_ (
  .A1({ Ckt432_M2_X2_8 }),
  .A2({ Ckt432_M1_X1_8 }),
  .A3({ in4 }),
  .A4({ Ckt432_M3_n12 }),
  .ZN({ Ckt432_M3_n5 })
);
NAND3_X1 #() 
NAND3_X1_10_ (
  .A1({ in4 }),
  .A2({ Ckt432_M4_n1 }),
  .A3({ Ckt432_M4_n2 }),
  .ZN({ Ckt432_I_8 })
);
NAND3_X1 #() 
NAND3_X1_11_ (
  .A1({ in43 }),
  .A2({ Ckt432_M4_n7 }),
  .A3({ Ckt432_M4_n8 }),
  .ZN({ Ckt432_I_5 })
);
AOI22_X1 #() 
AOI22_X1_1_ (
  .A1({ in37 }),
  .A2({ out223 }),
  .B1({ in47 }),
  .B2({ out329 }),
  .ZN({ Ckt432_M4_n8 })
);
NAND2_X1 #() 
NAND2_X1_10_ (
  .A1({ in53 }),
  .A2({ out370 }),
  .ZN({ Ckt432_M4_n7 })
);
NAND3_X1 #() 
NAND3_X1_12_ (
  .A1({ in56 }),
  .A2({ Ckt432_M4_n9 }),
  .A3({ Ckt432_M4_n10 }),
  .ZN({ Ckt432_I_4 })
);
AOI22_X1 #() 
AOI22_X1_2_ (
  .A1({ in50 }),
  .A2({ out223 }),
  .B1({ in60 }),
  .B2({ out329 }),
  .ZN({ Ckt432_M4_n10 })
);
NAND2_X1 #() 
NAND2_X1_11_ (
  .A1({ in66 }),
  .A2({ out370 }),
  .ZN({ Ckt432_M4_n9 })
);
NAND3_X1 #() 
NAND3_X1_13_ (
  .A1({ in69 }),
  .A2({ Ckt432_M4_n11 }),
  .A3({ Ckt432_M4_n12 }),
  .ZN({ Ckt432_I_3 })
);
AOI22_X1 #() 
AOI22_X1_3_ (
  .A1({ in63 }),
  .A2({ out223 }),
  .B1({ in73 }),
  .B2({ out329 }),
  .ZN({ Ckt432_M4_n12 })
);
NAND2_X1 #() 
NAND2_X1_12_ (
  .A1({ in79 }),
  .A2({ out370 }),
  .ZN({ Ckt432_M4_n11 })
);
NAND3_X1 #() 
NAND3_X1_14_ (
  .A1({ in82 }),
  .A2({ Ckt432_M4_n13 }),
  .A3({ Ckt432_M4_n14 }),
  .ZN({ Ckt432_I_2 })
);
AOI22_X1 #() 
AOI22_X1_4_ (
  .A1({ out223 }),
  .A2({ in1 }),
  .B1({ out329 }),
  .B2({ in8 }),
  .ZN({ Ckt432_M4_n2 })
);
AOI22_X1 #() 
AOI22_X1_5_ (
  .A1({ in76 }),
  .A2({ out223 }),
  .B1({ in86 }),
  .B2({ out329 }),
  .ZN({ Ckt432_M4_n14 })
);
NAND2_X1 #() 
NAND2_X1_13_ (
  .A1({ in92 }),
  .A2({ out370 }),
  .ZN({ Ckt432_M4_n13 })
);
NAND3_X1 #() 
NAND3_X1_15_ (
  .A1({ in95 }),
  .A2({ Ckt432_M4_n15 }),
  .A3({ Ckt432_M4_n16 }),
  .ZN({ Ckt432_I_1 })
);
AOI22_X1 #() 
AOI22_X1_6_ (
  .A1({ in89 }),
  .A2({ out223 }),
  .B1({ in99 }),
  .B2({ out329 }),
  .ZN({ Ckt432_M4_n16 })
);
NAND2_X1 #() 
NAND2_X1_14_ (
  .A1({ in105 }),
  .A2({ out370 }),
  .ZN({ Ckt432_M4_n15 })
);
NAND3_X1 #() 
NAND3_X1_16_ (
  .A1({ in108 }),
  .A2({ Ckt432_M4_n17 }),
  .A3({ Ckt432_M4_n18 }),
  .ZN({ Ckt432_I_0 })
);
AOI22_X1 #() 
AOI22_X1_7_ (
  .A1({ in102 }),
  .A2({ out223 }),
  .B1({ in112 }),
  .B2({ out329 }),
  .ZN({ Ckt432_M4_n18 })
);
NAND2_X1 #() 
NAND2_X1_15_ (
  .A1({ in115 }),
  .A2({ out370 }),
  .ZN({ Ckt432_M4_n17 })
);
NAND2_X1 #() 
NAND2_X1_16_ (
  .A1({ out370 }),
  .A2({ in14 }),
  .ZN({ Ckt432_M4_n1 })
);
NAND3_X1 #() 
NAND3_X1_17_ (
  .A1({ in17 }),
  .A2({ Ckt432_M4_n3 }),
  .A3({ Ckt432_M4_n4 }),
  .ZN({ Ckt432_I_7 })
);
AOI22_X1 #() 
AOI22_X1_8_ (
  .A1({ in11 }),
  .A2({ out223 }),
  .B1({ in21 }),
  .B2({ out329 }),
  .ZN({ Ckt432_M4_n4 })
);
NAND2_X1 #() 
NAND2_X1_17_ (
  .A1({ in27 }),
  .A2({ out370 }),
  .ZN({ Ckt432_M4_n3 })
);
NAND3_X1 #() 
NAND3_X1_18_ (
  .A1({ in30 }),
  .A2({ Ckt432_M4_n5 }),
  .A3({ Ckt432_M4_n6 }),
  .ZN({ Ckt432_I_6 })
);
AOI22_X1 #() 
AOI22_X1_9_ (
  .A1({ in24 }),
  .A2({ out223 }),
  .B1({ in34 }),
  .B2({ out329 }),
  .ZN({ Ckt432_M4_n6 })
);
NAND2_X1 #() 
NAND2_X1_18_ (
  .A1({ in40 }),
  .A2({ out370 }),
  .ZN({ Ckt432_M4_n5 })
);
AND2_X1 #() 
AND2_X1_1_ (
  .A1({ Ckt432_I_8 }),
  .A2({ Ckt432_M5_n1 }),
  .ZN({ out421 })
);
AOI221_X1 #() 
AOI221_X1_1_ (
  .A({ Ckt432_M5_n9 }),
  .B1({ Ckt432_I_2 }),
  .B2({ Ckt432_M5_n2 }),
  .C1({ Ckt432_I_4 }),
  .C2({ Ckt432_M5_n8 }),
  .ZN({ Ckt432_M5_n6 })
);
INV_X1 #() 
INV_X1_30_ (
  .A({ Ckt432_I_5 }),
  .ZN({ Ckt432_M5_n9 })
);
INV_X1 #() 
INV_X1_31_ (
  .A({ Ckt432_I_3 }),
  .ZN({ Ckt432_M5_n8 })
);
INV_X1 #() 
INV_X1_32_ (
  .A({ Ckt432_I_1 }),
  .ZN({ Ckt432_M5_n2 })
);
OR4_X1 #() 
OR4_X1_1_ (
  .A1({ Ckt432_M5_n2 }),
  .A2({ Ckt432_M5_n3 }),
  .A3({ Ckt432_M5_n4 }),
  .A4({ out430 }),
  .ZN({ Ckt432_M5_n1 })
);
INV_X1 #() 
INV_X1_33_ (
  .A({ Ckt432_I_0 }),
  .ZN({ Ckt432_M5_n3 })
);
NAND4_X1 #() 
NAND4_X1_12_ (
  .A1({ Ckt432_I_7 }),
  .A2({ Ckt432_I_6 }),
  .A3({ Ckt432_I_5 }),
  .A4({ Ckt432_I_4 }),
  .ZN({ out430 })
);
NAND3_X1 #() 
NAND3_X1_19_ (
  .A1({ Ckt432_I_6 }),
  .A2({ Ckt432_M5_n5 }),
  .A3({ Ckt432_I_7 }),
  .ZN({ out431 })
);
NAND3_X1 #() 
NAND3_X1_20_ (
  .A1({ Ckt432_I_4 }),
  .A2({ Ckt432_M5_n4 }),
  .A3({ Ckt432_I_5 }),
  .ZN({ Ckt432_M5_n5 })
);
NAND2_X1 #() 
NAND2_X1_19_ (
  .A1({ Ckt432_I_3 }),
  .A2({ Ckt432_I_2 }),
  .ZN({ Ckt432_M5_n4 })
);
OAI21_X1 #() 
OAI21_X1_10_ (
  .A({ Ckt432_I_7 }),
  .B1({ Ckt432_M5_n6 }),
  .B2({ Ckt432_M5_n7 }),
  .ZN({ out432 })
);
INV_X1 #() 
INV_X1_34_ (
  .A({ Ckt432_I_6 }),
  .ZN({ Ckt432_M5_n7 })
);

endmodule