module keyExpansion(key, w);

wire S0;
wire S1;
wire S2;
wire S3;
wire S4;
wire S5;
wire S6;
wire S7;
wire S8;
wire S9;
wire S10;
wire S11;
wire S12;
wire S13;
wire S14;
wire S15;
wire S16;
wire S17;
wire S18;
wire S19;
wire S20;
wire S21;
wire S22;
wire S23;
wire S24;
wire S25;
wire S26;
wire S27;
wire S28;
wire S29;
wire S30;
wire S31;
wire S32;
wire S33;
wire S34;
wire S35;
wire S36;
wire S37;
wire S38;
wire S39;
wire S40;
wire S41;
wire S42;
wire S43;
wire S44;
wire S45;
wire S46;
wire S47;
wire S48;
wire S49;
wire S50;
wire S51;
wire S52;
wire S53;
wire S54;
wire S55;
wire S56;
wire S57;
wire S58;
wire S59;
wire S60;
wire S61;
wire S62;
wire S63;
wire S64;
wire S65;
wire S66;
wire S67;
wire S68;
wire S69;
wire S70;
wire S71;
wire S72;
wire S73;
wire S74;
wire S75;
wire S76;
wire S77;
wire S78;
wire S79;
wire S80;
wire S81;
wire S82;
wire S83;
wire S84;
wire S85;
wire S86;
wire S87;
wire S88;
wire S89;
wire S90;
wire S91;
wire S92;
wire S93;
wire S94;
wire S95;
wire S96;
wire S97;
wire S98;
wire S99;
wire S100;
wire S101;
wire S102;
wire S103;
wire S104;
wire S105;
wire S106;
wire S107;
wire S108;
wire S109;
wire S110;
wire S111;
wire S112;
wire S113;
wire S114;
wire S115;
wire S116;
wire S117;
wire S118;
wire S119;
wire S120;
wire S121;
wire S122;
wire S123;
wire S124;
wire S125;
wire S126;
wire S127;
wire S128;
wire S129;
wire S130;
wire S131;
wire S132;
wire S133;
wire S134;
wire S135;
wire S136;
wire S137;
wire S138;
wire S139;
wire S140;
wire S141;
wire S142;
wire S143;
wire S144;
wire S145;
wire S146;
wire S147;
wire S148;
wire S149;
wire S150;
wire S151;
wire S152;
wire S153;
wire S154;
wire S155;
wire S156;
wire S157;
wire S158;
wire S159;
wire S160;
wire S161;
wire S162;
wire S163;
wire S164;
wire S165;
wire S166;
wire S167;
wire S168;
wire S169;
wire S170;
wire S171;
wire S172;
wire S173;
wire S174;
wire S175;
wire S176;
wire S177;
wire S178;
wire S179;
wire S180;
wire S181;
wire S182;
wire S183;
wire S184;
wire S185;
wire S186;
wire S187;
wire S188;
wire S189;
wire S190;
wire S191;
wire S192;
wire S193;
wire S194;
wire S195;
wire S196;
wire S197;
wire S198;
wire S199;
wire S200;
wire S201;
wire S202;
wire S203;
wire S204;
wire S205;
wire S206;
wire S207;
wire S208;
wire S209;
wire S210;
wire S211;
wire S212;
wire S213;
wire S214;
wire S215;
wire S216;
wire S217;
wire S218;
wire S219;
wire S220;
wire S221;
wire S222;
wire S223;
wire S224;
wire S225;
wire S226;
wire S227;
wire S228;
wire S229;
wire S230;
wire S231;
wire S232;
wire S233;
wire S234;
wire S235;
wire S236;
wire S237;
wire S238;
wire S239;
wire S240;
wire S241;
wire S242;
wire S243;
wire S244;
wire S245;
wire S246;
wire S247;
wire S248;
wire S249;
wire S250;
wire S251;
wire S252;
wire S253;
wire S254;
wire S255;
wire S256;
wire S257;
wire S258;
wire S259;
wire S260;
wire S261;
wire S262;
wire S263;
wire S264;
wire S265;
wire S266;
wire S267;
wire S268;
wire S269;
wire S270;
wire S271;
wire S272;
wire S273;
wire S274;
wire S275;
wire S276;
wire S277;
wire S278;
wire S279;
wire S280;
wire S281;
wire S282;
wire S283;
wire S284;
wire S285;
wire S286;
wire S287;
wire S288;
wire S289;
wire S290;
wire S291;
wire S292;
wire S293;
wire S294;
wire S295;
wire S296;
wire S297;
wire S298;
wire S299;
wire S300;
wire S301;
wire S302;
wire S303;
wire S304;
wire S305;
wire S306;
wire S307;
wire S308;
wire S309;
wire S310;
wire S311;
wire S312;
wire S313;
wire S314;
wire S315;
wire S316;
wire S317;
wire S318;
wire S319;
wire S320;
wire S321;
wire S322;
wire S323;
wire S324;
wire S325;
wire S326;
wire S327;
wire S328;
wire S329;
wire S330;
wire S331;
wire S332;
wire S333;
wire S334;
wire S335;
wire S336;
wire S337;
wire S338;
wire S339;
wire S340;
wire S341;
wire S342;
wire S343;
wire S344;
wire S345;
wire S346;
wire S347;
wire S348;
wire S349;
wire S350;
wire S351;
wire S352;
wire S353;
wire S354;
wire S355;
wire S356;
wire S357;
wire S358;
wire S359;
wire S360;
wire S361;
wire S362;
wire S363;
wire S364;
wire S365;
wire S366;
wire S367;
wire S368;
wire S369;
wire S370;
wire S371;
wire S372;
wire S373;
wire S374;
wire S375;
wire S376;
wire S377;
wire S378;
wire S379;
wire S380;
wire S381;
wire S382;
wire S383;
wire S384;
wire S385;
wire S386;
wire S387;
wire S388;
wire S389;
wire S390;
wire S391;
wire S392;
wire S393;
wire S394;
wire S395;
wire S396;
wire S397;
wire S398;
wire S399;
wire S400;
wire S401;
wire S402;
wire S403;
wire S404;
wire S405;
wire S406;
wire S407;
wire S408;
wire S409;
wire S410;
wire S411;
wire S412;
wire S413;
wire S414;
wire S415;
wire S416;
wire S417;
wire S418;
wire S419;
wire S420;
wire S421;
wire S422;
wire S423;
wire S424;
wire S425;
wire S426;
wire S427;
wire S428;
wire S429;
wire S430;
wire S431;
wire S432;
wire S433;
wire S434;
wire S435;
wire S436;
wire S437;
wire S438;
wire S439;
wire S440;
wire S441;
wire S442;
wire S443;
wire S444;
wire S445;
wire S446;
wire S447;
wire S448;
wire S449;
wire S450;
wire S451;
wire S452;
wire S453;
wire S454;
wire S455;
wire S456;
wire S457;
wire S458;
wire S459;
wire S460;
wire S461;
wire S462;
wire S463;
wire S464;
wire S465;
wire S466;
wire S467;
wire S468;
wire S469;
wire S470;
wire S471;
wire S472;
wire S473;
wire S474;
wire S475;
wire S476;
wire S477;
wire S478;
wire S479;
wire S480;
wire S481;
wire S482;
wire S483;
wire S484;
wire S485;
wire S486;
wire S487;
wire S488;
wire S489;
wire S490;
wire S491;
wire S492;
wire S493;
wire S494;
wire S495;
wire S496;
wire S497;
wire S498;
wire S499;
wire S500;
wire S501;
wire S502;
wire S503;
wire S504;
wire S505;
wire S506;
wire S507;
wire S508;
wire S509;
wire S510;
wire S511;
wire S512;
wire S513;
wire S514;
wire S515;
wire S516;
wire S517;
wire S518;
wire S519;
wire S520;
wire S521;
wire S522;
wire S523;
wire S524;
wire S525;
wire S526;
wire S527;
wire S528;
wire S529;
wire S530;
wire S531;
wire S532;
wire S533;
wire S534;
wire S535;
wire S536;
wire S537;
wire S538;
wire S539;
wire S540;
wire S541;
wire S542;
wire S543;
wire S544;
wire S545;
wire S546;
wire S547;
wire S548;
wire S549;
wire S550;
wire S551;
wire S552;
wire S553;
wire S554;
wire S555;
wire S556;
wire S557;
wire S558;
wire S559;
wire S560;
wire S561;
wire S562;
wire S563;
wire S564;
wire S565;
wire S566;
wire S567;
wire S568;
wire S569;
wire S570;
wire S571;
wire S572;
wire S573;
wire S574;
wire S575;
wire S576;
wire S577;
wire S578;
wire S579;
wire S580;
wire S581;
wire S582;
wire S583;
wire S584;
wire S585;
wire S586;
wire S587;
wire S588;
wire S589;
wire S590;
wire S591;
wire S592;
wire S593;
wire S594;
wire S595;
wire S596;
wire S597;
wire S598;
wire S599;
wire S600;
wire S601;
wire S602;
wire S603;
wire S604;
wire S605;
wire S606;
wire S607;
wire S608;
wire S609;
wire S610;
wire S611;
wire S612;
wire S613;
wire S614;
wire S615;
wire S616;
wire S617;
wire S618;
wire S619;
wire S620;
wire S621;
wire S622;
wire S623;
wire S624;
wire S625;
wire S626;
wire S627;
wire S628;
wire S629;
wire S630;
wire S631;
wire S632;
wire S633;
wire S634;
wire S635;
wire S636;
wire S637;
wire S638;
wire S639;
wire S640;
wire S641;
wire S642;
wire S643;
wire S644;
wire S645;
wire S646;
wire S647;
wire S648;
wire S649;
wire S650;
wire S651;
wire S652;
wire S653;
wire S654;
wire S655;
wire S656;
wire S657;
wire S658;
wire S659;
wire S660;
wire S661;
wire S662;
wire S663;
wire S664;
wire S665;
wire S666;
wire S667;
wire S668;
wire S669;
wire S670;
wire S671;
wire S672;
wire S673;
wire S674;
wire S675;
wire S676;
wire S677;
wire S678;
wire S679;
wire S680;
wire S681;
wire S682;
wire S683;
wire S684;
wire S685;
wire S686;
wire S687;
wire S688;
wire S689;
wire S690;
wire S691;
wire S692;
wire S693;
wire S694;
wire S695;
wire S696;
wire S697;
wire S698;
wire S699;
wire S700;
wire S701;
wire S702;
wire S703;
wire S704;
wire S705;
wire S706;
wire S707;
wire S708;
wire S709;
wire S710;
wire S711;
wire S712;
wire S713;
wire S714;
wire S715;
wire S716;
wire S717;
wire S718;
wire S719;
wire S720;
wire S721;
wire S722;
wire S723;
wire S724;
wire S725;
wire S726;
wire S727;
wire S728;
wire S729;
wire S730;
wire S731;
wire S732;
wire S733;
wire S734;
wire S735;
wire S736;
wire S737;
wire S738;
wire S739;
wire S740;
wire S741;
wire S742;
wire S743;
wire S744;
wire S745;
wire S746;
wire S747;
wire S748;
wire S749;
wire S750;
wire S751;
wire S752;
wire S753;
wire S754;
wire S755;
wire S756;
wire S757;
wire S758;
wire S759;
wire S760;
wire S761;
wire S762;
wire S763;
wire S764;
wire S765;
wire S766;
wire S767;
wire S768;
wire S769;
wire S770;
wire S771;
wire S772;
wire S773;
wire S774;
wire S775;
wire S776;
wire S777;
wire S778;
wire S779;
wire S780;
wire S781;
wire S782;
wire S783;
wire S784;
wire S785;
wire S786;
wire S787;
wire S788;
wire S789;
wire S790;
wire S791;
wire S792;
wire S793;
wire S794;
wire S795;
wire S796;
wire S797;
wire S798;
wire S799;
wire S800;
wire S801;
wire S802;
wire S803;
wire S804;
wire S805;
wire S806;
wire S807;
wire S808;
wire S809;
wire S810;
wire S811;
wire S812;
wire S813;
wire S814;
wire S815;
wire S816;
wire S817;
wire S818;
wire S819;
wire S820;
wire S821;
wire S822;
wire S823;
wire S824;
wire S825;
wire S826;
wire S827;
wire S828;
wire S829;
wire S830;
wire S831;
wire S832;
wire S833;
wire S834;
wire S835;
wire S836;
wire S837;
wire S838;
wire S839;
wire S840;
wire S841;
wire S842;
wire S843;
wire S844;
wire S845;
wire S846;
wire S847;
wire S848;
wire S849;
wire S850;
wire S851;
wire S852;
wire S853;
wire S854;
wire S855;
wire S856;
wire S857;
wire S858;
wire S859;
wire S860;
wire S861;
wire S862;
wire S863;
wire S864;
wire S865;
wire S866;
wire S867;
wire S868;
wire S869;
wire S870;
wire S871;
wire S872;
wire S873;
wire S874;
wire S875;
wire S876;
wire S877;
wire S878;
wire S879;
wire S880;
wire S881;
wire S882;
wire S883;
wire S884;
wire S885;
wire S886;
wire S887;
wire S888;
wire S889;
wire S890;
wire S891;
wire S892;
wire S893;
wire S894;
wire S895;
wire S896;
wire S897;
wire S898;
wire S899;
wire S900;
wire S901;
wire S902;
wire S903;
wire S904;
wire S905;
wire S906;
wire S907;
wire S908;
wire S909;
wire S910;
wire S911;
wire S912;
wire S913;
wire S914;
wire S915;
wire S916;
wire S917;
wire S918;
wire S919;
wire S920;
wire S921;
wire S922;
wire S923;
wire S924;
wire S925;
wire S926;
wire S927;
wire S928;
wire S929;
wire S930;
wire S931;
wire S932;
wire S933;
wire S934;
wire S935;
wire S936;
wire S937;
wire S938;
wire S939;
wire S940;
wire S941;
wire S942;
wire S943;
wire S944;
wire S945;
wire S946;
wire S947;
wire S948;
wire S949;
wire S950;
wire S951;
wire S952;
wire S953;
wire S954;
wire S955;
wire S956;
wire S957;
wire S958;
wire S959;
wire S960;
wire S961;
wire S962;
wire S963;
wire S964;
wire S965;
wire S966;
wire S967;
wire S968;
wire S969;
wire S970;
wire S971;
wire S972;
wire S973;
wire S974;
wire S975;
wire S976;
wire S977;
wire S978;
wire S979;
wire S980;
wire S981;
wire S982;
wire S983;
wire S984;
wire S985;
wire S986;
wire S987;
wire S988;
wire S989;
wire S990;
wire S991;
wire S992;
wire S993;
wire S994;
wire S995;
wire S996;
wire S997;
wire S998;
wire S999;
wire S1000;
wire S1001;
wire S1002;
wire S1003;
wire S1004;
wire S1005;
wire S1006;
wire S1007;
wire S1008;
wire S1009;
wire S1010;
wire S1011;
wire S1012;
wire S1013;
wire S1014;
wire S1015;
wire S1016;
wire S1017;
wire S1018;
wire S1019;
wire S1020;
wire S1021;
wire S1022;
wire S1023;
wire S1024;
wire S1025;
wire S1026;
wire S1027;
wire S1028;
wire S1029;
wire S1030;
wire S1031;
wire S1032;
wire S1033;
wire S1034;
wire S1035;
wire S1036;
wire S1037;
wire S1038;
wire S1039;
wire S1040;
wire S1041;
wire S1042;
wire S1043;
wire S1044;
wire S1045;
wire S1046;
wire S1047;
wire S1048;
wire S1049;
wire S1050;
wire S1051;
wire S1052;
wire S1053;
wire S1054;
wire S1055;
wire S1056;
wire S1057;
wire S1058;
wire S1059;
wire S1060;
wire S1061;
wire S1062;
wire S1063;
wire S1064;
wire S1065;
wire S1066;
wire S1067;
wire S1068;
wire S1069;
wire S1070;
wire S1071;
wire S1072;
wire S1073;
wire S1074;
wire S1075;
wire S1076;
wire S1077;
wire S1078;
wire S1079;
wire S1080;
wire S1081;
wire S1082;
wire S1083;
wire S1084;
wire S1085;
wire S1086;
wire S1087;
wire S1088;
wire S1089;
wire S1090;
wire S1091;
wire S1092;
wire S1093;
wire S1094;
wire S1095;
wire S1096;
wire S1097;
wire S1098;
wire S1099;
wire S1100;
wire S1101;
wire S1102;
wire S1103;
wire S1104;
wire S1105;
wire S1106;
wire S1107;
wire S1108;
wire S1109;
wire S1110;
wire S1111;
wire S1112;
wire S1113;
wire S1114;
wire S1115;
wire S1116;
wire S1117;
wire S1118;
wire S1119;
wire S1120;
wire S1121;
wire S1122;
wire S1123;
wire S1124;
wire S1125;
wire S1126;
wire S1127;
wire S1128;
wire S1129;
wire S1130;
wire S1131;
wire S1132;
wire S1133;
wire S1134;
wire S1135;
wire S1136;
wire S1137;
wire S1138;
wire S1139;
wire S1140;
wire S1141;
wire S1142;
wire S1143;
wire S1144;
wire S1145;
wire S1146;
wire S1147;
wire S1148;
wire S1149;
wire S1150;
wire S1151;
wire S1152;
wire S1153;
wire S1154;
wire S1155;
wire S1156;
wire S1157;
wire S1158;
wire S1159;
wire S1160;
wire S1161;
wire S1162;
wire S1163;
wire S1164;
wire S1165;
wire S1166;
wire S1167;
wire S1168;
wire S1169;
wire S1170;
wire S1171;
wire S1172;
wire S1173;
wire S1174;
wire S1175;
wire S1176;
wire S1177;
wire S1178;
wire S1179;
wire S1180;
wire S1181;
wire S1182;
wire S1183;
wire S1184;
wire S1185;
wire S1186;
wire S1187;
wire S1188;
wire S1189;
wire S1190;
wire S1191;
wire S1192;
wire S1193;
wire S1194;
wire S1195;
wire S1196;
wire S1197;
wire S1198;
wire S1199;
wire S1200;
wire S1201;
wire S1202;
wire S1203;
wire S1204;
wire S1205;
wire S1206;
wire S1207;
wire S1208;
wire S1209;
wire S1210;
wire S1211;
wire S1212;
wire S1213;
wire S1214;
wire S1215;
wire S1216;
wire S1217;
wire S1218;
wire S1219;
wire S1220;
wire S1221;
wire S1222;
wire S1223;
wire S1224;
wire S1225;
wire S1226;
wire S1227;
wire S1228;
wire S1229;
wire S1230;
wire S1231;
wire S1232;
wire S1233;
wire S1234;
wire S1235;
wire S1236;
wire S1237;
wire S1238;
wire S1239;
wire S1240;
wire S1241;
wire S1242;
wire S1243;
wire S1244;
wire S1245;
wire S1246;
wire S1247;
wire S1248;
wire S1249;
wire S1250;
wire S1251;
wire S1252;
wire S1253;
wire S1254;
wire S1255;
wire S1256;
wire S1257;
wire S1258;
wire S1259;
wire S1260;
wire S1261;
wire S1262;
wire S1263;
wire S1264;
wire S1265;
wire S1266;
wire S1267;
wire S1268;
wire S1269;
wire S1270;
wire S1271;
wire S1272;
wire S1273;
wire S1274;
wire S1275;
wire S1276;
wire S1277;
wire S1278;
wire S1279;
wire S1280;
wire S1281;
wire S1282;
wire S1283;
wire S1284;
wire S1285;
wire S1286;
wire S1287;
wire S1288;
wire S1289;
wire S1290;
wire S1291;
wire S1292;
wire S1293;
wire S1294;
wire S1295;
wire S1296;
wire S1297;
wire S1298;
wire S1299;
wire S1300;
wire S1301;
wire S1302;
wire S1303;
wire S1304;
wire S1305;
wire S1306;
wire S1307;
wire S1308;
wire S1309;
wire S1310;
wire S1311;
wire S1312;
wire S1313;
wire S1314;
wire S1315;
wire S1316;
wire S1317;
wire S1318;
wire S1319;
wire S1320;
wire S1321;
wire S1322;
wire S1323;
wire S1324;
wire S1325;
wire S1326;
wire S1327;
wire S1328;
wire S1329;
wire S1330;
wire S1331;
wire S1332;
wire S1333;
wire S1334;
wire S1335;
wire S1336;
wire S1337;
wire S1338;
wire S1339;
wire S1340;
wire S1341;
wire S1342;
wire S1343;
wire S1344;
wire S1345;
wire S1346;
wire S1347;
wire S1348;
wire S1349;
wire S1350;
wire S1351;
wire S1352;
wire S1353;
wire S1354;
wire S1355;
wire S1356;
wire S1357;
wire S1358;
wire S1359;
wire S1360;
wire S1361;
wire S1362;
wire S1363;
wire S1364;
wire S1365;
wire S1366;
wire S1367;
wire S1368;
wire S1369;
wire S1370;
wire S1371;
wire S1372;
wire S1373;
wire S1374;
wire S1375;
wire S1376;
wire S1377;
wire S1378;
wire S1379;
wire S1380;
wire S1381;
wire S1382;
wire S1383;
wire S1384;
wire S1385;
wire S1386;
wire S1387;
wire S1388;
wire S1389;
wire S1390;
wire S1391;
wire S1392;
wire S1393;
wire S1394;
wire S1395;
wire S1396;
wire S1397;
wire S1398;
wire S1399;
wire S1400;
wire S1401;
wire S1402;
wire S1403;
wire S1404;
wire S1405;
wire S1406;
wire S1407;
wire S1408;
wire S1409;
wire S1410;
wire S1411;
wire S1412;
wire S1413;
wire S1414;
wire S1415;
wire S1416;
wire S1417;
wire S1418;
wire S1419;
wire S1420;
wire S1421;
wire S1422;
wire S1423;
wire S1424;
wire S1425;
wire S1426;
wire S1427;
wire S1428;
wire S1429;
wire S1430;
wire S1431;
wire S1432;
wire S1433;
wire S1434;
wire S1435;
wire S1436;
wire S1437;
wire S1438;
wire S1439;
wire S1440;
wire S1441;
wire S1442;
wire S1443;
wire S1444;
wire S1445;
wire S1446;
wire S1447;
wire S1448;
wire S1449;
wire S1450;
wire S1451;
wire S1452;
wire S1453;
wire S1454;
wire S1455;
wire S1456;
wire S1457;
wire S1458;
wire S1459;
wire S1460;
wire S1461;
wire S1462;
wire S1463;
wire S1464;
wire S1465;
wire S1466;
wire S1467;
wire S1468;
wire S1469;
wire S1470;
wire S1471;
wire S1472;
wire S1473;
wire S1474;
wire S1475;
wire S1476;
wire S1477;
wire S1478;
wire S1479;
wire S1480;
wire S1481;
wire S1482;
wire S1483;
wire S1484;
wire S1485;
wire S1486;
wire S1487;
wire S1488;
wire S1489;
wire S1490;
wire S1491;
wire S1492;
wire S1493;
wire S1494;
wire S1495;
wire S1496;
wire S1497;
wire S1498;
wire S1499;
wire S1500;
wire S1501;
wire S1502;
wire S1503;
wire S1504;
wire S1505;
wire S1506;
wire S1507;
wire S1508;
wire S1509;
wire S1510;
wire S1511;
wire S1512;
wire S1513;
wire S1514;
wire S1515;
wire S1516;
wire S1517;
wire S1518;
wire S1519;
wire S1520;
wire S1521;
wire S1522;
wire S1523;
wire S1524;
wire S1525;
wire S1526;
wire S1527;
wire S1528;
wire S1529;
wire S1530;
wire S1531;
wire S1532;
wire S1533;
wire S1534;
wire S1535;
wire S1536;
wire S1537;
wire S1538;
wire S1539;
wire S1540;
wire S1541;
wire S1542;
wire S1543;
wire S1544;
wire S1545;
wire S1546;
wire S1547;
wire S1548;
wire S1549;
wire S1550;
wire S1551;
wire S1552;
wire S1553;
wire S1554;
wire S1555;
wire S1556;
wire S1557;
wire S1558;
wire S1559;
wire S1560;
wire S1561;
wire S1562;
wire S1563;
wire S1564;
wire S1565;
wire S1566;
wire S1567;
wire S1568;
wire S1569;
wire S1570;
wire S1571;
wire S1572;
wire S1573;
wire S1574;
wire S1575;
wire S1576;
wire S1577;
wire S1578;
wire S1579;
wire S1580;
wire S1581;
wire S1582;
wire S1583;
wire S1584;
wire S1585;
wire S1586;
wire S1587;
wire S1588;
wire S1589;
wire S1590;
wire S1591;
wire S1592;
wire S1593;
wire S1594;
wire S1595;
wire S1596;
wire S1597;
wire S1598;
wire S1599;
wire S1600;
wire S1601;
wire S1602;
wire S1603;
wire S1604;
wire S1605;
wire S1606;
wire S1607;
wire S1608;
wire S1609;
wire S1610;
wire S1611;
wire S1612;
wire S1613;
wire S1614;
wire S1615;
wire S1616;
wire S1617;
wire S1618;
wire S1619;
wire S1620;
wire S1621;
wire S1622;
wire S1623;
wire S1624;
wire S1625;
wire S1626;
wire S1627;
wire S1628;
wire S1629;
wire S1630;
wire S1631;
wire S1632;
wire S1633;
wire S1634;
wire S1635;
wire S1636;
wire S1637;
wire S1638;
wire S1639;
wire S1640;
wire S1641;
wire S1642;
wire S1643;
wire S1644;
wire S1645;
wire S1646;
wire S1647;
wire S1648;
wire S1649;
wire S1650;
wire S1651;
wire S1652;
wire S1653;
wire S1654;
wire S1655;
wire S1656;
wire S1657;
wire S1658;
wire S1659;
wire S1660;
wire S1661;
wire S1662;
wire S1663;
wire S1664;
wire S1665;
wire S1666;
wire S1667;
wire S1668;
wire S1669;
wire S1670;
wire S1671;
wire S1672;
wire S1673;
wire S1674;
wire S1675;
wire S1676;
wire S1677;
wire S1678;
wire S1679;
wire S1680;
wire S1681;
wire S1682;
wire S1683;
wire S1684;
wire S1685;
wire S1686;
wire S1687;
wire S1688;
wire S1689;
wire S1690;
wire S1691;
wire S1692;
wire S1693;
wire S1694;
wire S1695;
wire S1696;
wire S1697;
wire S1698;
wire S1699;
wire S1700;
wire S1701;
wire S1702;
wire S1703;
wire S1704;
wire S1705;
wire S1706;
wire S1707;
wire S1708;
wire S1709;
wire S1710;
wire S1711;
wire S1712;
wire S1713;
wire S1714;
wire S1715;
wire S1716;
wire S1717;
wire S1718;
wire S1719;
wire S1720;
wire S1721;
wire S1722;
wire S1723;
wire S1724;
wire S1725;
wire S1726;
wire S1727;
wire S1728;
wire S1729;
wire S1730;
wire S1731;
wire S1732;
wire S1733;
wire S1734;
wire S1735;
wire S1736;
wire S1737;
wire S1738;
wire S1739;
wire S1740;
wire S1741;
wire S1742;
wire S1743;
wire S1744;
wire S1745;
wire S1746;
wire S1747;
wire S1748;
wire S1749;
wire S1750;
wire S1751;
wire S1752;
wire S1753;
wire S1754;
wire S1755;
wire S1756;
wire S1757;
wire S1758;
wire S1759;
wire S1760;
wire S1761;
wire S1762;
wire S1763;
wire S1764;
wire S1765;
wire S1766;
wire S1767;
wire S1768;
wire S1769;
wire S1770;
wire S1771;
wire S1772;
wire S1773;
wire S1774;
wire S1775;
wire S1776;
wire S1777;
wire S1778;
wire S1779;
wire S1780;
wire S1781;
wire S1782;
wire S1783;
wire S1784;
wire S1785;
wire S1786;
wire S1787;
wire S1788;
wire S1789;
wire S1790;
wire S1791;
wire S1792;
wire S1793;
wire S1794;
wire S1795;
wire S1796;
wire S1797;
wire S1798;
wire S1799;
wire S1800;
wire S1801;
wire S1802;
wire S1803;
wire S1804;
wire S1805;
wire S1806;
wire S1807;
wire S1808;
wire S1809;
wire S1810;
wire S1811;
wire S1812;
wire S1813;
wire S1814;
wire S1815;
wire S1816;
wire S1817;
wire S1818;
wire S1819;
wire S1820;
wire S1821;
wire S1822;
wire S1823;
wire S1824;
wire S1825;
wire S1826;
wire S1827;
wire S1828;
wire S1829;
wire S1830;
wire S1831;
wire S1832;
wire S1833;
wire S1834;
wire S1835;
wire S1836;
wire S1837;
wire S1838;
wire S1839;
wire S1840;
wire S1841;
wire S1842;
wire S1843;
wire S1844;
wire S1845;
wire S1846;
wire S1847;
wire S1848;
wire S1849;
wire S1850;
wire S1851;
wire S1852;
wire S1853;
wire S1854;
wire S1855;
wire S1856;
wire S1857;
wire S1858;
wire S1859;
wire S1860;
wire S1861;
wire S1862;
wire S1863;
wire S1864;
wire S1865;
wire S1866;
wire S1867;
wire S1868;
wire S1869;
wire S1870;
wire S1871;
wire S1872;
wire S1873;
wire S1874;
wire S1875;
wire S1876;
wire S1877;
wire S1878;
wire S1879;
wire S1880;
wire S1881;
wire S1882;
wire S1883;
wire S1884;
wire S1885;
wire S1886;
wire S1887;
wire S1888;
wire S1889;
wire S1890;
wire S1891;
wire S1892;
wire S1893;
wire S1894;
wire S1895;
wire S1896;
wire S1897;
wire S1898;
wire S1899;
wire S1900;
wire S1901;
wire S1902;
wire S1903;
wire S1904;
wire S1905;
wire S1906;
wire S1907;
wire S1908;
wire S1909;
wire S1910;
wire S1911;
wire S1912;
wire S1913;
wire S1914;
wire S1915;
wire S1916;
wire S1917;
wire S1918;
wire S1919;
wire S1920;
wire S1921;
wire S1922;
wire S1923;
wire S1924;
wire S1925;
wire S1926;
wire S1927;
wire S1928;
wire S1929;
wire S1930;
wire S1931;
wire S1932;
wire S1933;
wire S1934;
wire S1935;
wire S1936;
wire S1937;
wire S1938;
wire S1939;
wire S1940;
wire S1941;
wire S1942;
wire S1943;
wire S1944;
wire S1945;
wire S1946;
wire S1947;
wire S1948;
wire S1949;
wire S1950;
wire S1951;
wire S1952;
wire S1953;
wire S1954;
wire S1955;
wire S1956;
wire S1957;
wire S1958;
wire S1959;
wire S1960;
wire S1961;
wire S1962;
wire S1963;
wire S1964;
wire S1965;
wire S1966;
wire S1967;
wire S1968;
wire S1969;
wire S1970;
wire S1971;
wire S1972;
wire S1973;
wire S1974;
wire S1975;
wire S1976;
wire S1977;
wire S1978;
wire S1979;
wire S1980;
wire S1981;
wire S1982;
wire S1983;
wire S1984;
wire S1985;
wire S1986;
wire S1987;
wire S1988;
wire S1989;
wire S1990;
wire S1991;
wire S1992;
wire S1993;
wire S1994;
wire S1995;
wire S1996;
wire S1997;
wire S1998;
wire S1999;
wire S2000;
wire S2001;
wire S2002;
wire S2003;
wire S2004;
wire S2005;
wire S2006;
wire S2007;
wire S2008;
wire S2009;
wire S2010;
wire S2011;
wire S2012;
wire S2013;
wire S2014;
wire S2015;
wire S2016;
wire S2017;
wire S2018;
wire S2019;
wire S2020;
wire S2021;
wire S2022;
wire S2023;
wire S2024;
wire S2025;
wire S2026;
wire S2027;
wire S2028;
wire S2029;
wire S2030;
wire S2031;
wire S2032;
wire S2033;
wire S2034;
wire S2035;
wire S2036;
wire S2037;
wire S2038;
wire S2039;
wire S2040;
wire S2041;
wire S2042;
wire S2043;
wire S2044;
wire S2045;
wire S2046;
wire S2047;
wire S2048;
wire S2049;
wire S2050;
wire S2051;
wire S2052;
wire S2053;
wire S2054;
wire S2055;
wire S2056;
wire S2057;
wire S2058;
wire S2059;
wire S2060;
wire S2061;
wire S2062;
wire S2063;
wire S2064;
wire S2065;
wire S2066;
wire S2067;
wire S2068;
wire S2069;
wire S2070;
wire S2071;
wire S2072;
wire S2073;
wire S2074;
wire S2075;
wire S2076;
wire S2077;
wire S2078;
wire S2079;
wire S2080;
wire S2081;
wire S2082;
wire S2083;
wire S2084;
wire S2085;
wire S2086;
wire S2087;
wire S2088;
wire S2089;
wire S2090;
wire S2091;
wire S2092;
wire S2093;
wire S2094;
wire S2095;
wire S2096;
wire S2097;
wire S2098;
wire S2099;
wire S2100;
wire S2101;
wire S2102;
wire S2103;
wire S2104;
wire S2105;
wire S2106;
wire S2107;
wire S2108;
wire S2109;
wire S2110;
wire S2111;
wire S2112;
wire S2113;
wire S2114;
wire S2115;
wire S2116;
wire S2117;
wire S2118;
wire S2119;
wire S2120;
wire S2121;
wire S2122;
wire S2123;
wire S2124;
wire S2125;
wire S2126;
wire S2127;
wire S2128;
wire S2129;
wire S2130;
wire S2131;
wire S2132;
wire S2133;
wire S2134;
wire S2135;
wire S2136;
wire S2137;
wire S2138;
wire S2139;
wire S2140;
wire S2141;
wire S2142;
wire S2143;
wire S2144;
wire S2145;
wire S2146;
wire S2147;
wire S2148;
wire S2149;
wire S2150;
wire S2151;
wire S2152;
wire S2153;
wire S2154;
wire S2155;
wire S2156;
wire S2157;
wire S2158;
wire S2159;
wire S2160;
wire S2161;
wire S2162;
wire S2163;
wire S2164;
wire S2165;
wire S2166;
wire S2167;
wire S2168;
wire S2169;
wire S2170;
wire S2171;
wire S2172;
wire S2173;
wire S2174;
wire S2175;
wire S2176;
wire S2177;
wire S2178;
wire S2179;
wire S2180;
wire S2181;
wire S2182;
wire S2183;
wire S2184;
wire S2185;
wire S2186;
wire S2187;
wire S2188;
wire S2189;
wire S2190;
wire S2191;
wire S2192;
wire S2193;
wire S2194;
wire S2195;
wire S2196;
wire S2197;
wire S2198;
wire S2199;
wire S2200;
wire S2201;
wire S2202;
wire S2203;
wire S2204;
wire S2205;
wire S2206;
wire S2207;
wire S2208;
wire S2209;
wire S2210;
wire S2211;
wire S2212;
wire S2213;
wire S2214;
wire S2215;
wire S2216;
wire S2217;
wire S2218;
wire S2219;
wire S2220;
wire S2221;
wire S2222;
wire S2223;
wire S2224;
wire S2225;
wire S2226;
wire S2227;
wire S2228;
wire S2229;
wire S2230;
wire S2231;
wire S2232;
wire S2233;
wire S2234;
wire S2235;
wire S2236;
wire S2237;
wire S2238;
wire S2239;
wire S2240;
wire S2241;
wire S2242;
wire S2243;
wire S2244;
wire S2245;
wire S2246;
wire S2247;
wire S2248;
wire S2249;
wire S2250;
wire S2251;
wire S2252;
wire S2253;
wire S2254;
wire S2255;
wire S2256;
wire S2257;
wire S2258;
wire S2259;
wire S2260;
wire S2261;
wire S2262;
wire S2263;
wire S2264;
wire S2265;
wire S2266;
wire S2267;
wire S2268;
wire S2269;
wire S2270;
wire S2271;
wire S2272;
wire S2273;
wire S2274;
wire S2275;
wire S2276;
wire S2277;
wire S2278;
wire S2279;
wire S2280;
wire S2281;
wire S2282;
wire S2283;
wire S2284;
wire S2285;
wire S2286;
wire S2287;
wire S2288;
wire S2289;
wire S2290;
wire S2291;
wire S2292;
wire S2293;
wire S2294;
wire S2295;
wire S2296;
wire S2297;
wire S2298;
wire S2299;
wire S2300;
wire S2301;
wire S2302;
wire S2303;
wire S2304;
wire S2305;
wire S2306;
wire S2307;
wire S2308;
wire S2309;
wire S2310;
wire S2311;
wire S2312;
wire S2313;
wire S2314;
wire S2315;
wire S2316;
wire S2317;
wire S2318;
wire S2319;
wire S2320;
wire S2321;
wire S2322;
wire S2323;
wire S2324;
wire S2325;
wire S2326;
wire S2327;
wire S2328;
wire S2329;
wire S2330;
wire S2331;
wire S2332;
wire S2333;
wire S2334;
wire S2335;
wire S2336;
wire S2337;
wire S2338;
wire S2339;
wire S2340;
wire S2341;
wire S2342;
wire S2343;
wire S2344;
wire S2345;
wire S2346;
wire S2347;
wire S2348;
wire S2349;
wire S2350;
wire S2351;
wire S2352;
wire S2353;
wire S2354;
wire S2355;
wire S2356;
wire S2357;
wire S2358;
wire S2359;
wire S2360;
wire S2361;
wire S2362;
wire S2363;
wire S2364;
wire S2365;
wire S2366;
wire S2367;
wire S2368;
wire S2369;
wire S2370;
wire S2371;
wire S2372;
wire S2373;
wire S2374;
wire S2375;
wire S2376;
wire S2377;
wire S2378;
wire S2379;
wire S2380;
wire S2381;
wire S2382;
wire S2383;
wire S2384;
wire S2385;
wire S2386;
wire S2387;
wire S2388;
wire S2389;
wire S2390;
wire S2391;
wire S2392;
wire S2393;
wire S2394;
wire S2395;
wire S2396;
wire S2397;
wire S2398;
wire S2399;
wire S2400;
wire S2401;
wire S2402;
wire S2403;
wire S2404;
wire S2405;
wire S2406;
wire S2407;
wire S2408;
wire S2409;
wire S2410;
wire S2411;
wire S2412;
wire S2413;
wire S2414;
wire S2415;
wire S2416;
wire S2417;
wire S2418;
wire S2419;
wire S2420;
wire S2421;
wire S2422;
wire S2423;
wire S2424;
wire S2425;
wire S2426;
wire S2427;
wire S2428;
wire S2429;
wire S2430;
wire S2431;
wire S2432;
wire S2433;
wire S2434;
wire S2435;
wire S2436;
wire S2437;
wire S2438;
wire S2439;
wire S2440;
wire S2441;
wire S2442;
wire S2443;
wire S2444;
wire S2445;
wire S2446;
wire S2447;
wire S2448;
wire S2449;
wire S2450;
wire S2451;
wire S2452;
wire S2453;
wire S2454;
wire S2455;
wire S2456;
wire S2457;
wire S2458;
wire S2459;
wire S2460;
wire S2461;
wire S2462;
wire S2463;
wire S2464;
wire S2465;
wire S2466;
wire S2467;
wire S2468;
wire S2469;
wire S2470;
wire S2471;
wire S2472;
wire S2473;
wire S2474;
wire S2475;
wire S2476;
wire S2477;
wire S2478;
wire S2479;
wire S2480;
wire S2481;
wire S2482;
wire S2483;
wire S2484;
wire S2485;
wire S2486;
wire S2487;
wire S2488;
wire S2489;
wire S2490;
wire S2491;
wire S2492;
wire S2493;
wire S2494;
wire S2495;
wire S2496;
wire S2497;
wire S2498;
wire S2499;
wire S2500;
wire S2501;
wire S2502;
wire S2503;
wire S2504;
wire S2505;
wire S2506;
wire S2507;
wire S2508;
wire S2509;
wire S2510;
wire S2511;
wire S2512;
wire S2513;
wire S2514;
wire S2515;
wire S2516;
wire S2517;
wire S2518;
wire S2519;
wire S2520;
wire S2521;
wire S2522;
wire S2523;
wire S2524;
wire S2525;
wire S2526;
wire S2527;
wire S2528;
wire S2529;
wire S2530;
wire S2531;
wire S2532;
wire S2533;
wire S2534;
wire S2535;
wire S2536;
wire S2537;
wire S2538;
wire S2539;
wire S2540;
wire S2541;
wire S2542;
wire S2543;
wire S2544;
wire S2545;
wire S2546;
wire S2547;
wire S2548;
wire S2549;
wire S2550;
wire S2551;
wire S2552;
wire S2553;
wire S2554;
wire S2555;
wire S2556;
wire S2557;
wire S2558;
wire S2559;
wire S2560;
wire S2561;
wire S2562;
wire S2563;
wire S2564;
wire S2565;
wire S2566;
wire S2567;
wire S2568;
wire S2569;
wire S2570;
wire S2571;
wire S2572;
wire S2573;
wire S2574;
wire S2575;
wire S2576;
wire S2577;
wire S2578;
wire S2579;
wire S2580;
wire S2581;
wire S2582;
wire S2583;
wire S2584;
wire S2585;
wire S2586;
wire S2587;
wire S2588;
wire S2589;
wire S2590;
wire S2591;
wire S2592;
wire S2593;
wire S2594;
wire S2595;
wire S2596;
wire S2597;
wire S2598;
wire S2599;
wire S2600;
wire S2601;
wire S2602;
wire S2603;
wire S2604;
wire S2605;
wire S2606;
wire S2607;
wire S2608;
wire S2609;
wire S2610;
wire S2611;
wire S2612;
wire S2613;
wire S2614;
wire S2615;
wire S2616;
wire S2617;
wire S2618;
wire S2619;
wire S2620;
wire S2621;
wire S2622;
wire S2623;
wire S2624;
wire S2625;
wire S2626;
wire S2627;
wire S2628;
wire S2629;
wire S2630;
wire S2631;
wire S2632;
wire S2633;
wire S2634;
wire S2635;
wire S2636;
wire S2637;
wire S2638;
wire S2639;
wire S2640;
wire S2641;
wire S2642;
wire S2643;
wire S2644;
wire S2645;
wire S2646;
wire S2647;
wire S2648;
wire S2649;
wire S2650;
wire S2651;
wire S2652;
wire S2653;
wire S2654;
wire S2655;
wire S2656;
wire S2657;
wire S2658;
wire S2659;
wire S2660;
wire S2661;
wire S2662;
wire S2663;
wire S2664;
wire S2665;
wire S2666;
wire S2667;
wire S2668;
wire S2669;
wire S2670;
wire S2671;
wire S2672;
wire S2673;
wire S2674;
wire S2675;
wire S2676;
wire S2677;
wire S2678;
wire S2679;
wire S2680;
wire S2681;
wire S2682;
wire S2683;
wire S2684;
wire S2685;
wire S2686;
wire S2687;
wire S2688;
wire S2689;
wire S2690;
wire S2691;
wire S2692;
wire S2693;
wire S2694;
wire S2695;
wire S2696;
wire S2697;
wire S2698;
wire S2699;
wire S2700;
wire S2701;
wire S2702;
wire S2703;
wire S2704;
wire S2705;
wire S2706;
wire S2707;
wire S2708;
wire S2709;
wire S2710;
wire S2711;
wire S2712;
wire S2713;
wire S2714;
wire S2715;
wire S2716;
wire S2717;
wire S2718;
wire S2719;
wire S2720;
wire S2721;
wire S2722;
wire S2723;
wire S2724;
wire S2725;
wire S2726;
wire S2727;
wire S2728;
wire S2729;
wire S2730;
wire S2731;
wire S2732;
wire S2733;
wire S2734;
wire S2735;
wire S2736;
wire S2737;
wire S2738;
wire S2739;
wire S2740;
wire S2741;
wire S2742;
wire S2743;
wire S2744;
wire S2745;
wire S2746;
wire S2747;
wire S2748;
wire S2749;
wire S2750;
wire S2751;
wire S2752;
wire S2753;
wire S2754;
wire S2755;
wire S2756;
wire S2757;
wire S2758;
wire S2759;
wire S2760;
wire S2761;
wire S2762;
wire S2763;
wire S2764;
wire S2765;
wire S2766;
wire S2767;
wire S2768;
wire S2769;
wire S2770;
wire S2771;
wire S2772;
wire S2773;
wire S2774;
wire S2775;
wire S2776;
wire S2777;
wire S2778;
wire S2779;
wire S2780;
wire S2781;
wire S2782;
wire S2783;
wire S2784;
wire S2785;
wire S2786;
wire S2787;
wire S2788;
wire S2789;
wire S2790;
wire S2791;
wire S2792;
wire S2793;
wire S2794;
wire S2795;
wire S2796;
wire S2797;
wire S2798;
wire S2799;
wire S2800;
wire S2801;
wire S2802;
wire S2803;
wire S2804;
wire S2805;
wire S2806;
wire S2807;
wire S2808;
wire S2809;
wire S2810;
wire S2811;
wire S2812;
wire S2813;
wire S2814;
wire S2815;
wire S2816;
wire S2817;
wire S2818;
wire S2819;
wire S2820;
wire S2821;
wire S2822;
wire S2823;
wire S2824;
wire S2825;
wire S2826;
wire S2827;
wire S2828;
wire S2829;
wire S2830;
wire S2831;
wire S2832;
wire S2833;
wire S2834;
wire S2835;
wire S2836;
wire S2837;
wire S2838;
wire S2839;
wire S2840;
wire S2841;
wire S2842;
wire S2843;
wire S2844;
wire S2845;
wire S2846;
wire S2847;
wire S2848;
wire S2849;
wire S2850;
wire S2851;
wire S2852;
wire S2853;
wire S2854;
wire S2855;
wire S2856;
wire S2857;
wire S2858;
wire S2859;
wire S2860;
wire S2861;
wire S2862;
wire S2863;
wire S2864;
wire S2865;
wire S2866;
wire S2867;
wire S2868;
wire S2869;
wire S2870;
wire S2871;
wire S2872;
wire S2873;
wire S2874;
wire S2875;
wire S2876;
wire S2877;
wire S2878;
wire S2879;
wire S2880;
wire S2881;
wire S2882;
wire S2883;
wire S2884;
wire S2885;
wire S2886;
wire S2887;
wire S2888;
wire S2889;
wire S2890;
wire S2891;
wire S2892;
wire S2893;
wire S2894;
wire S2895;
wire S2896;
wire S2897;
wire S2898;
wire S2899;
wire S2900;
wire S2901;
wire S2902;
wire S2903;
wire S2904;
wire S2905;
wire S2906;
wire S2907;
wire S2908;
wire S2909;
wire S2910;
wire S2911;
wire S2912;
wire S2913;
wire S2914;
wire S2915;
wire S2916;
wire S2917;
wire S2918;
wire S2919;
wire S2920;
wire S2921;
wire S2922;
wire S2923;
wire S2924;
wire S2925;
wire S2926;
wire S2927;
wire S2928;
wire S2929;
wire S2930;
wire S2931;
wire S2932;
wire S2933;
wire S2934;
wire S2935;
wire S2936;
wire S2937;
wire S2938;
wire S2939;
wire S2940;
wire S2941;
wire S2942;
wire S2943;
wire S2944;
wire S2945;
wire S2946;
wire S2947;
wire S2948;
wire S2949;
wire S2950;
wire S2951;
wire S2952;
wire S2953;
wire S2954;
wire S2955;
wire S2956;
wire S2957;
wire S2958;
wire S2959;
wire S2960;
wire S2961;
wire S2962;
wire S2963;
wire S2964;
wire S2965;
wire S2966;
wire S2967;
wire S2968;
wire S2969;
wire S2970;
wire S2971;
wire S2972;
wire S2973;
wire S2974;
wire S2975;
wire S2976;
wire S2977;
wire S2978;
wire S2979;
wire S2980;
wire S2981;
wire S2982;
wire S2983;
wire S2984;
wire S2985;
wire S2986;
wire S2987;
wire S2988;
wire S2989;
wire S2990;
wire S2991;
wire S2992;
wire S2993;
wire S2994;
wire S2995;
wire S2996;
wire S2997;
wire S2998;
wire S2999;
wire S3000;
wire S3001;
wire S3002;
wire S3003;
wire S3004;
wire S3005;
wire S3006;
wire S3007;
wire S3008;
wire S3009;
wire S3010;
wire S3011;
wire S3012;
wire S3013;
wire S3014;
wire S3015;
wire S3016;
wire S3017;
wire S3018;
wire S3019;
wire S3020;
wire S3021;
wire S3022;
wire S3023;
wire S3024;
wire S3025;
wire S3026;
wire S3027;
wire S3028;
wire S3029;
wire S3030;
wire S3031;
wire S3032;
wire S3033;
wire S3034;
wire S3035;
wire S3036;
wire S3037;
wire S3038;
wire S3039;
wire S3040;
wire S3041;
wire S3042;
wire S3043;
wire S3044;
wire S3045;
wire S3046;
wire S3047;
wire S3048;
wire S3049;
wire S3050;
wire S3051;
wire S3052;
wire S3053;
wire S3054;
wire S3055;
wire S3056;
wire S3057;
wire S3058;
wire S3059;
wire S3060;
wire S3061;
wire S3062;
wire S3063;
wire S3064;
wire S3065;
wire S3066;
wire S3067;
wire S3068;
wire S3069;
wire S3070;
wire S3071;
wire S3072;
wire S3073;
wire S3074;
wire S3075;
wire S3076;
wire S3077;
wire S3078;
wire S3079;
wire S3080;
wire S3081;
wire S3082;
wire S3083;
wire S3084;
wire S3085;
wire S3086;
wire S3087;
wire S3088;
wire S3089;
wire S3090;
wire S3091;
wire S3092;
wire S3093;
wire S3094;
wire S3095;
wire S3096;
wire S3097;
wire S3098;
wire S3099;
wire S3100;
wire S3101;
wire S3102;
wire S3103;
wire S3104;
wire S3105;
wire S3106;
wire S3107;
wire S3108;
wire S3109;
wire S3110;
wire S3111;
wire S3112;
wire S3113;
wire S3114;
wire S3115;
wire S3116;
wire S3117;
wire S3118;
wire S3119;
wire S3120;
wire S3121;
wire S3122;
wire S3123;
wire S3124;
wire S3125;
wire S3126;
wire S3127;
wire S3128;
wire S3129;
wire S3130;
wire S3131;
wire S3132;
wire S3133;
wire S3134;
wire S3135;
wire S3136;
wire S3137;
wire S3138;
wire S3139;
wire S3140;
wire S3141;
wire S3142;
wire S3143;
wire S3144;
wire S3145;
wire S3146;
wire S3147;
wire S3148;
wire S3149;
wire S3150;
wire S3151;
wire S3152;
wire S3153;
wire S3154;
wire S3155;
wire S3156;
wire S3157;
wire S3158;
wire S3159;
wire S3160;
wire S3161;
wire S3162;
wire S3163;
wire S3164;
wire S3165;
wire S3166;
wire S3167;
wire S3168;
wire S3169;
wire S3170;
wire S3171;
wire S3172;
wire S3173;
wire S3174;
wire S3175;
wire S3176;
wire S3177;
wire S3178;
wire S3179;
wire S3180;
wire S3181;
wire S3182;
wire S3183;
wire S3184;
wire S3185;
wire S3186;
wire S3187;
wire S3188;
wire S3189;
wire S3190;
wire S3191;
wire S3192;
wire S3193;
wire S3194;
wire S3195;
wire S3196;
wire S3197;
wire S3198;
wire S3199;
wire S3200;
wire S3201;
wire S3202;
wire S3203;
wire S3204;
wire S3205;
wire S3206;
wire S3207;
wire S3208;
wire S3209;
wire S3210;
wire S3211;
wire S3212;
wire S3213;
wire S3214;
wire S3215;
wire S3216;
wire S3217;
wire S3218;
wire S3219;
wire S3220;
wire S3221;
wire S3222;
wire S3223;
wire S3224;
wire S3225;
wire S3226;
wire S3227;
wire S3228;
wire S3229;
wire S3230;
wire S3231;
wire S3232;
wire S3233;
wire S3234;
wire S3235;
wire S3236;
wire S3237;
wire S3238;
wire S3239;
wire S3240;
wire S3241;
wire S3242;
wire S3243;
wire S3244;
wire S3245;
wire S3246;
wire S3247;
wire S3248;
wire S3249;
wire S3250;
wire S3251;
wire S3252;
wire S3253;
wire S3254;
wire S3255;
wire S3256;
wire S3257;
wire S3258;
wire S3259;
wire S3260;
wire S3261;
wire S3262;
wire S3263;
wire S3264;
wire S3265;
wire S3266;
wire S3267;
wire S3268;
wire S3269;
wire S3270;
wire S3271;
wire S3272;
wire S3273;
wire S3274;
wire S3275;
wire S3276;
wire S3277;
wire S3278;
wire S3279;
wire S3280;
wire S3281;
wire S3282;
wire S3283;
wire S3284;
wire S3285;
wire S3286;
wire S3287;
wire S3288;
wire S3289;
wire S3290;
wire S3291;
wire S3292;
wire S3293;
wire S3294;
wire S3295;
wire S3296;
wire S3297;
wire S3298;
wire S3299;
wire S3300;
wire S3301;
wire S3302;
wire S3303;
wire S3304;
wire S3305;
wire S3306;
wire S3307;
wire S3308;
wire S3309;
wire S3310;
wire S3311;
wire S3312;
wire S3313;
wire S3314;
wire S3315;
wire S3316;
wire S3317;
wire S3318;
wire S3319;
wire S3320;
wire S3321;
wire S3322;
wire S3323;
wire S3324;
wire S3325;
wire S3326;
wire S3327;
wire S3328;
wire S3329;
wire S3330;
wire S3331;
wire S3332;
wire S3333;
wire S3334;
wire S3335;
wire S3336;
wire S3337;
wire S3338;
wire S3339;
wire S3340;
wire S3341;
wire S3342;
wire S3343;
wire S3344;
wire S3345;
wire S3346;
wire S3347;
wire S3348;
wire S3349;
wire S3350;
wire S3351;
wire S3352;
wire S3353;
wire S3354;
wire S3355;
wire S3356;
wire S3357;
wire S3358;
wire S3359;
wire S3360;
wire S3361;
wire S3362;
wire S3363;
wire S3364;
wire S3365;
wire S3366;
wire S3367;
wire S3368;
wire S3369;
wire S3370;
wire S3371;
wire S3372;
wire S3373;
wire S3374;
wire S3375;
wire S3376;
wire S3377;
wire S3378;
wire S3379;
wire S3380;
wire S3381;
wire S3382;
wire S3383;
wire S3384;
wire S3385;
wire S3386;
wire S3387;
wire S3388;
wire S3389;
wire S3390;
wire S3391;
wire S3392;
wire S3393;
wire S3394;
wire S3395;
wire S3396;
wire S3397;
wire S3398;
wire S3399;
wire S3400;
wire S3401;
wire S3402;
wire S3403;
wire S3404;
wire S3405;
wire S3406;
wire S3407;
wire S3408;
wire S3409;
wire S3410;
wire S3411;
wire S3412;
wire S3413;
wire S3414;
wire S3415;
wire S3416;
wire S3417;
wire S3418;
wire S3419;
wire S3420;
wire S3421;
wire S3422;
wire S3423;
wire S3424;
wire S3425;
wire S3426;
wire S3427;
wire S3428;
wire S3429;
wire S3430;
wire S3431;
wire S3432;
wire S3433;
wire S3434;
wire S3435;
wire S3436;
wire S3437;
wire S3438;
wire S3439;
wire S3440;
wire S3441;
wire S3442;
wire S3443;
wire S3444;
wire S3445;
wire S3446;
wire S3447;
wire S3448;
wire S3449;
wire S3450;
wire S3451;
wire S3452;
wire S3453;
wire S3454;
wire S3455;
wire S3456;
wire S3457;
wire S3458;
wire S3459;
wire S3460;
wire S3461;
wire S3462;
wire S3463;
wire S3464;
wire S3465;
wire S3466;
wire S3467;
wire S3468;
wire S3469;
wire S3470;
wire S3471;
wire S3472;
wire S3473;
wire S3474;
wire S3475;
wire S3476;
wire S3477;
wire S3478;
wire S3479;
wire S3480;
wire S3481;
wire S3482;
wire S3483;
wire S3484;
wire S3485;
wire S3486;
wire S3487;
wire S3488;
wire S3489;
wire S3490;
wire S3491;
wire S3492;
wire S3493;
wire S3494;
wire S3495;
wire S3496;
wire S3497;
wire S3498;
wire S3499;
wire S3500;
wire S3501;
wire S3502;
wire S3503;
wire S3504;
wire S3505;
wire S3506;
wire S3507;
wire S3508;
wire S3509;
wire S3510;
wire S3511;
wire S3512;
wire S3513;
wire S3514;
wire S3515;
wire S3516;
wire S3517;
wire S3518;
wire S3519;
wire S3520;
wire S3521;
wire S3522;
wire S3523;
wire S3524;
wire S3525;
wire S3526;
wire S3527;
wire S3528;
wire S3529;
wire S3530;
wire S3531;
wire S3532;
wire S3533;
wire S3534;
wire S3535;
wire S3536;
wire S3537;
wire S3538;
wire S3539;
wire S3540;
wire S3541;
wire S3542;
wire S3543;
wire S3544;
wire S3545;
wire S3546;
wire S3547;
wire S3548;
wire S3549;
wire S3550;
wire S3551;
wire S3552;
wire S3553;
wire S3554;
wire S3555;
wire S3556;
wire S3557;
wire S3558;
wire S3559;
wire S3560;
wire S3561;
wire S3562;
wire S3563;
wire S3564;
wire S3565;
wire S3566;
wire S3567;
wire S3568;
wire S3569;
wire S3570;
wire S3571;
wire S3572;
wire S3573;
wire S3574;
wire S3575;
wire S3576;
wire S3577;
wire S3578;
wire S3579;
wire S3580;
wire S3581;
wire S3582;
wire S3583;
wire S3584;
wire S3585;
wire S3586;
wire S3587;
wire S3588;
wire S3589;
wire S3590;
wire S3591;
wire S3592;
wire S3593;
wire S3594;
wire S3595;
wire S3596;
wire S3597;
wire S3598;
wire S3599;
wire S3600;
wire S3601;
wire S3602;
wire S3603;
wire S3604;
wire S3605;
wire S3606;
wire S3607;
wire S3608;
wire S3609;
wire S3610;
wire S3611;
wire S3612;
wire S3613;
wire S3614;
wire S3615;
wire S3616;
wire S3617;
wire S3618;
wire S3619;
wire S3620;
wire S3621;
wire S3622;
wire S3623;
wire S3624;
wire S3625;
wire S3626;
wire S3627;
wire S3628;
wire S3629;
wire S3630;
wire S3631;
wire S3632;
wire S3633;
wire S3634;
wire S3635;
wire S3636;
wire S3637;
wire S3638;
wire S3639;
wire S3640;
wire S3641;
wire S3642;
wire S3643;
wire S3644;
wire S3645;
wire S3646;
wire S3647;
wire S3648;
wire S3649;
wire S3650;
wire S3651;
wire S3652;
wire S3653;
wire S3654;
wire S3655;
wire S3656;
wire S3657;
wire S3658;
wire S3659;
wire S3660;
wire S3661;
wire S3662;
wire S3663;
wire S3664;
wire S3665;
wire S3666;
wire S3667;
wire S3668;
wire S3669;
wire S3670;
wire S3671;
wire S3672;
wire S3673;
wire S3674;
wire S3675;
wire S3676;
wire S3677;
wire S3678;
wire S3679;
wire S3680;
wire S3681;
wire S3682;
wire S3683;
wire S3684;
wire S3685;
wire S3686;
wire S3687;
wire S3688;
wire S3689;
wire S3690;
wire S3691;
wire S3692;
wire S3693;
wire S3694;
wire S3695;
wire S3696;
wire S3697;
wire S3698;
wire S3699;
wire S3700;
wire S3701;
wire S3702;
wire S3703;
wire S3704;
wire S3705;
wire S3706;
wire S3707;
wire S3708;
wire S3709;
wire S3710;
wire S3711;
wire S3712;
wire S3713;
wire S3714;
wire S3715;
wire S3716;
wire S3717;
wire S3718;
wire S3719;
wire S3720;
wire S3721;
wire S3722;
wire S3723;
wire S3724;
wire S3725;
wire S3726;
wire S3727;
wire S3728;
wire S3729;
wire S3730;
wire S3731;
wire S3732;
wire S3733;
wire S3734;
wire S3735;
wire S3736;
wire S3737;
wire S3738;
wire S3739;
wire S3740;
wire S3741;
wire S3742;
wire S3743;
wire S3744;
wire S3745;
wire S3746;
wire S3747;
wire S3748;
wire S3749;
wire S3750;
wire S3751;
wire S3752;
wire S3753;
wire S3754;
wire S3755;
wire S3756;
wire S3757;
wire S3758;
wire S3759;
wire S3760;
wire S3761;
wire S3762;
wire S3763;
wire S3764;
wire S3765;
wire S3766;
wire S3767;
wire S3768;
wire S3769;
wire S3770;
wire S3771;
wire S3772;
wire S3773;
wire S3774;
wire S3775;
wire S3776;
wire S3777;
wire S3778;
wire S3779;
wire S3780;
wire S3781;
wire S3782;
wire S3783;
wire S3784;
wire S3785;
wire S3786;
wire S3787;
wire S3788;
wire S3789;
wire S3790;
wire S3791;
wire S3792;
wire S3793;
wire S3794;
wire S3795;
wire S3796;
wire S3797;
wire S3798;
wire S3799;
wire S3800;
wire S3801;
wire S3802;
wire S3803;
wire S3804;
wire S3805;
wire S3806;
wire S3807;
wire S3808;
wire S3809;
wire S3810;
wire S3811;
wire S3812;
wire S3813;
wire S3814;
wire S3815;
wire S3816;
wire S3817;
wire S3818;
wire S3819;
wire S3820;
wire S3821;
wire S3822;
wire S3823;
wire S3824;
wire S3825;
wire S3826;
wire S3827;
wire S3828;
wire S3829;
wire S3830;
wire S3831;
wire S3832;
wire S3833;
wire S3834;
wire S3835;
wire S3836;
wire S3837;
wire S3838;
wire S3839;
wire S3840;
wire S3841;
wire S3842;
wire S3843;
wire S3844;
wire S3845;
wire S3846;
wire S3847;
wire S3848;
wire S3849;
wire S3850;
wire S3851;
wire S3852;
wire S3853;
wire S3854;
wire S3855;
wire S3856;
wire S3857;
wire S3858;
wire S3859;
wire S3860;
wire S3861;
wire S3862;
wire S3863;
wire S3864;
wire S3865;
wire S3866;
wire S3867;
wire S3868;
wire S3869;
wire S3870;
wire S3871;
wire S3872;
wire S3873;
wire S3874;
wire S3875;
wire S3876;
wire S3877;
wire S3878;
wire S3879;
wire S3880;
wire S3881;
wire S3882;
wire S3883;
wire S3884;
wire S3885;
wire S3886;
wire S3887;
wire S3888;
wire S3889;
wire S3890;
wire S3891;
wire S3892;
wire S3893;
wire S3894;
wire S3895;
wire S3896;
wire S3897;
wire S3898;
wire S3899;
wire S3900;
wire S3901;
wire S3902;
wire S3903;
wire S3904;
wire S3905;
wire S3906;
wire S3907;
wire S3908;
wire S3909;
wire S3910;
wire S3911;
wire S3912;
wire S3913;
wire S3914;
wire S3915;
wire S3916;
wire S3917;
wire S3918;
wire S3919;
wire S3920;
wire S3921;
wire S3922;
wire S3923;
wire S3924;
wire S3925;
wire S3926;
wire S3927;
wire S3928;
wire S3929;
wire S3930;
wire S3931;
wire S3932;
wire S3933;
wire S3934;
wire S3935;
wire S3936;
wire S3937;
wire S3938;
wire S3939;
wire S3940;
wire S3941;
wire S3942;
wire S3943;
wire S3944;
wire S3945;
wire S3946;
wire S3947;
wire S3948;
wire S3949;
wire S3950;
wire S3951;
wire S3952;
wire S3953;
wire S3954;
wire S3955;
wire S3956;
wire S3957;
wire S3958;
wire S3959;
wire S3960;
wire S3961;
wire S3962;
wire S3963;
wire S3964;
wire S3965;
wire S3966;
wire S3967;
wire S3968;
wire S3969;
wire S3970;
wire S3971;
wire S3972;
wire S3973;
wire S3974;
wire S3975;
wire S3976;
wire S3977;
wire S3978;
wire S3979;
wire S3980;
wire S3981;
wire S3982;
wire S3983;
wire S3984;
wire S3985;
wire S3986;
wire S3987;
wire S3988;
wire S3989;
wire S3990;
wire S3991;
wire S3992;
wire S3993;
wire S3994;
wire S3995;
wire S3996;
wire S3997;
wire S3998;
wire S3999;
wire S4000;
wire S4001;
wire S4002;
wire S4003;
wire S4004;
wire S4005;
wire S4006;
wire S4007;
wire S4008;
wire S4009;
wire S4010;
wire S4011;
wire S4012;
wire S4013;
wire S4014;
wire S4015;
wire S4016;
wire S4017;
wire S4018;
wire S4019;
wire S4020;
wire S4021;
wire S4022;
wire S4023;
wire S4024;
wire S4025;
wire S4026;
wire S4027;
wire S4028;
wire S4029;
wire S4030;
wire S4031;
wire S4032;
wire S4033;
wire S4034;
wire S4035;
wire S4036;
wire S4037;
wire S4038;
wire S4039;
wire S4040;
wire S4041;
wire S4042;
wire S4043;
wire S4044;
wire S4045;
wire S4046;
wire S4047;
wire S4048;
wire S4049;
wire S4050;
wire S4051;
wire S4052;
wire S4053;
wire S4054;
wire S4055;
wire S4056;
wire S4057;
wire S4058;
wire S4059;
wire S4060;
wire S4061;
wire S4062;
wire S4063;
wire S4064;
wire S4065;
wire S4066;
wire S4067;
wire S4068;
wire S4069;
wire S4070;
wire S4071;
wire S4072;
wire S4073;
wire S4074;
wire S4075;
wire S4076;
wire S4077;
wire S4078;
wire S4079;
wire S4080;
wire S4081;
wire S4082;
wire S4083;
wire S4084;
wire S4085;
wire S4086;
wire S4087;
wire S4088;
wire S4089;
wire S4090;
wire S4091;
wire S4092;
wire S4093;
wire S4094;
wire S4095;
wire S4096;
wire S4097;
wire S4098;
wire S4099;
wire S4100;
wire S4101;
wire S4102;
wire S4103;
wire S4104;
wire S4105;
wire S4106;
wire S4107;
wire S4108;
wire S4109;
wire S4110;
wire S4111;
wire S4112;
wire S4113;
wire S4114;
wire S4115;
wire S4116;
wire S4117;
wire S4118;
wire S4119;
wire S4120;
wire S4121;
wire S4122;
wire S4123;
wire S4124;
wire S4125;
wire S4126;
wire S4127;
wire S4128;
wire S4129;
wire S4130;
wire S4131;
wire S4132;
wire S4133;
wire S4134;
wire S4135;
wire S4136;
wire S4137;
wire S4138;
wire S4139;
wire S4140;
wire S4141;
wire S4142;
wire S4143;
wire S4144;
wire S4145;
wire S4146;
wire S4147;
wire S4148;
wire S4149;
wire S4150;
wire S4151;
wire S4152;
wire S4153;
wire S4154;
wire S4155;
wire S4156;
wire S4157;
wire S4158;
wire S4159;
wire S4160;
wire S4161;
wire S4162;
wire S4163;
wire S4164;
wire S4165;
wire S4166;
wire S4167;
wire S4168;
wire S4169;
wire S4170;
wire S4171;
wire S4172;
wire S4173;
wire S4174;
wire S4175;
wire S4176;
wire S4177;
wire S4178;
wire S4179;
wire S4180;
wire S4181;
wire S4182;
wire S4183;
wire S4184;
wire S4185;
wire S4186;
wire S4187;
wire S4188;
wire S4189;
wire S4190;
wire S4191;
wire S4192;
wire S4193;
wire S4194;
wire S4195;
wire S4196;
wire S4197;
wire S4198;
wire S4199;
wire S4200;
wire S4201;
wire S4202;
wire S4203;
wire S4204;
wire S4205;
wire S4206;
wire S4207;
wire S4208;
wire S4209;
wire S4210;
wire S4211;
wire S4212;
wire S4213;
wire S4214;
wire S4215;
wire S4216;
wire S4217;
wire S4218;
wire S4219;
wire S4220;
wire S4221;
wire S4222;
wire S4223;
wire S4224;
wire S4225;
wire S4226;
wire S4227;
wire S4228;
wire S4229;
wire S4230;
wire S4231;
wire S4232;
wire S4233;
wire S4234;
wire S4235;
wire S4236;
wire S4237;
wire S4238;
wire S4239;
wire S4240;
wire S4241;
wire S4242;
wire S4243;
wire S4244;
wire S4245;
wire S4246;
wire S4247;
wire S4248;
wire S4249;
wire S4250;
wire S4251;
wire S4252;
wire S4253;
wire S4254;
wire S4255;
wire S4256;
wire S4257;
wire S4258;
wire S4259;
wire S4260;
wire S4261;
wire S4262;
wire S4263;
wire S4264;
wire S4265;
wire S4266;
wire S4267;
wire S4268;
wire S4269;
wire S4270;
wire S4271;
wire S4272;
wire S4273;
wire S4274;
wire S4275;
wire S4276;
wire S4277;
wire S4278;
wire S4279;
wire S4280;
wire S4281;
wire S4282;
wire S4283;
wire S4284;
wire S4285;
wire S4286;
wire S4287;
wire S4288;
wire S4289;
wire S4290;
wire S4291;
wire S4292;
wire S4293;
wire S4294;
wire S4295;
wire S4296;
wire S4297;
wire S4298;
wire S4299;
wire S4300;
wire S4301;
wire S4302;
wire S4303;
wire S4304;
wire S4305;
wire S4306;
wire S4307;
wire S4308;
wire S4309;
wire S4310;
wire S4311;
wire S4312;
wire S4313;
wire S4314;
wire S4315;
wire S4316;
wire S4317;
wire S4318;
wire S4319;
wire S4320;
wire S4321;
wire S4322;
wire S4323;
wire S4324;
wire S4325;
wire S4326;
wire S4327;
wire S4328;
wire S4329;
wire S4330;
wire S4331;
wire S4332;
wire S4333;
wire S4334;
wire S4335;
wire S4336;
wire S4337;
wire S4338;
wire S4339;
wire S4340;
wire S4341;
wire S4342;
wire S4343;
wire S4344;
wire S4345;
wire S4346;
wire S4347;
wire S4348;
wire S4349;
wire S4350;
wire S4351;
wire S4352;
wire S4353;
wire S4354;
wire S4355;
wire S4356;
wire S4357;
wire S4358;
wire S4359;
wire S4360;
wire S4361;
wire S4362;
wire S4363;
wire S4364;
wire S4365;
wire S4366;
wire S4367;
wire S4368;
wire S4369;
wire S4370;
wire S4371;
wire S4372;
wire S4373;
wire S4374;
wire S4375;
wire S4376;
wire S4377;
wire S4378;
wire S4379;
wire S4380;
wire S4381;
wire S4382;
wire S4383;
wire S4384;
wire S4385;
wire S4386;
wire S4387;
wire S4388;
wire S4389;
wire S4390;
wire S4391;
wire S4392;
wire S4393;
wire S4394;
wire S4395;
wire S4396;
wire S4397;
wire S4398;
wire S4399;
wire S4400;
wire S4401;
wire S4402;
wire S4403;
wire S4404;
wire S4405;
wire S4406;
wire S4407;
wire S4408;
wire S4409;
wire S4410;
wire S4411;
wire S4412;
wire S4413;
wire S4414;
wire S4415;
wire S4416;
wire S4417;
wire S4418;
wire S4419;
wire S4420;
wire S4421;
wire S4422;
wire S4423;
wire S4424;
wire S4425;
wire S4426;
wire S4427;
wire S4428;
wire S4429;
wire S4430;
wire S4431;
wire S4432;
wire S4433;
wire S4434;
wire S4435;
wire S4436;
wire S4437;
wire S4438;
wire S4439;
wire S4440;
wire S4441;
wire S4442;
wire S4443;
wire S4444;
wire S4445;
wire S4446;
wire S4447;
wire S4448;
wire S4449;
wire S4450;
wire S4451;
wire S4452;
wire S4453;
wire S4454;
wire S4455;
wire S4456;
wire S4457;
wire S4458;
wire S4459;
wire S4460;
wire S4461;
wire S4462;
wire S4463;
wire S4464;
wire S4465;
wire S4466;
wire S4467;
wire S4468;
wire S4469;
wire S4470;
wire S4471;
wire S4472;
wire S4473;
wire S4474;
wire S4475;
wire S4476;
wire S4477;
wire S4478;
wire S4479;
wire S4480;
wire S4481;
wire S4482;
wire S4483;
wire S4484;
wire S4485;
wire S4486;
wire S4487;
wire S4488;
wire S4489;
wire S4490;
wire S4491;
wire S4492;
wire S4493;
wire S4494;
wire S4495;
wire S4496;
wire S4497;
wire S4498;
wire S4499;
wire S4500;
wire S4501;
wire S4502;
wire S4503;
wire S4504;
wire S4505;
wire S4506;
wire S4507;
wire S4508;
wire S4509;
wire S4510;
wire S4511;
wire S4512;
wire S4513;
wire S4514;
wire S4515;
wire S4516;
wire S4517;
wire S4518;
wire S4519;
wire S4520;
wire S4521;
wire S4522;
wire S4523;
wire S4524;
wire S4525;
wire S4526;
wire S4527;
wire S4528;
wire S4529;
wire S4530;
wire S4531;
wire S4532;
wire S4533;
wire S4534;
wire S4535;
wire S4536;
wire S4537;
wire S4538;
wire S4539;
wire S4540;
wire S4541;
wire S4542;
wire S4543;
wire S4544;
wire S4545;
wire S4546;
wire S4547;
wire S4548;
wire S4549;
wire S4550;
wire S4551;
wire S4552;
wire S4553;
wire S4554;
wire S4555;
wire S4556;
wire S4557;
wire S4558;
wire S4559;
wire S4560;
wire S4561;
wire S4562;
wire S4563;
wire S4564;
wire S4565;
wire S4566;
wire S4567;
wire S4568;
wire S4569;
wire S4570;
wire S4571;
wire S4572;
wire S4573;
wire S4574;
wire S4575;
wire S4576;
wire S4577;
wire S4578;
wire S4579;
wire S4580;
wire S4581;
wire S4582;
wire S4583;
wire S4584;
wire S4585;
wire S4586;
wire S4587;
wire S4588;
wire S4589;
wire S4590;
wire S4591;
wire S4592;
wire S4593;
wire S4594;
wire S4595;
wire S4596;
wire S4597;
wire S4598;
wire S4599;
wire S4600;
wire S4601;
wire S4602;
wire S4603;
wire S4604;
wire S4605;
wire S4606;
wire S4607;
wire S4608;
wire S4609;
wire S4610;
wire S4611;
wire S4612;
wire S4613;
wire S4614;
wire S4615;
wire S4616;
wire S4617;
wire S4618;
wire S4619;
wire S4620;
wire S4621;
wire S4622;
wire S4623;
wire S4624;
wire S4625;
wire S4626;
wire S4627;
wire S4628;
wire S4629;
wire S4630;
wire S4631;
wire S4632;
wire S4633;
wire S4634;
wire S4635;
wire S4636;
wire S4637;
wire S4638;
wire S4639;
wire S4640;
wire S4641;
wire S4642;
wire S4643;
wire S4644;
wire S4645;
wire S4646;
wire S4647;
wire S4648;
wire S4649;
wire S4650;
wire S4651;
wire S4652;
wire S4653;
wire S4654;
wire S4655;
wire S4656;
wire S4657;
wire S4658;
wire S4659;
wire S4660;
wire S4661;
wire S4662;
wire S4663;
wire S4664;
wire S4665;
wire S4666;
wire S4667;
wire S4668;
wire S4669;
wire S4670;
wire S4671;
wire S4672;
wire S4673;
wire S4674;
wire S4675;
wire S4676;
wire S4677;
wire S4678;
wire S4679;
wire S4680;
wire S4681;
wire S4682;
wire S4683;
wire S4684;
wire S4685;
wire S4686;
wire S4687;
wire S4688;
wire S4689;
wire S4690;
wire S4691;
wire S4692;
wire S4693;
wire S4694;
wire S4695;
wire S4696;
wire S4697;
wire S4698;
wire S4699;
wire S4700;
wire S4701;
wire S4702;
wire S4703;
wire S4704;
wire S4705;
wire S4706;
wire S4707;
wire S4708;
wire S4709;
wire S4710;
wire S4711;
wire S4712;
wire S4713;
wire S4714;
wire S4715;
wire S4716;
wire S4717;
wire S4718;
wire S4719;
wire S4720;
wire S4721;
wire S4722;
wire S4723;
wire S4724;
wire S4725;
wire S4726;
wire S4727;
wire S4728;
wire S4729;
wire S4730;
wire S4731;
wire S4732;
wire S4733;
wire S4734;
wire S4735;
wire S4736;
wire S4737;
wire S4738;
wire S4739;
wire S4740;
wire S4741;
wire S4742;
wire S4743;
wire S4744;
wire S4745;
wire S4746;
wire S4747;
wire S4748;
wire S4749;
wire S4750;
wire S4751;
wire S4752;
wire S4753;
wire S4754;
wire S4755;
wire S4756;
wire S4757;
wire S4758;
wire S4759;
wire S4760;
wire S4761;
wire S4762;
wire S4763;
wire S4764;
wire S4765;
wire S4766;
wire S4767;
wire S4768;
wire S4769;
wire S4770;
wire S4771;
wire S4772;
wire S4773;
wire S4774;
wire S4775;
wire S4776;
wire S4777;
wire S4778;
wire S4779;
wire S4780;
wire S4781;
wire S4782;
wire S4783;
wire S4784;
wire S4785;
wire S4786;
wire S4787;
wire S4788;
wire S4789;
wire S4790;
wire S4791;
wire S4792;
wire S4793;
wire S4794;
wire S4795;
wire S4796;
wire S4797;
wire S4798;
wire S4799;
wire S4800;
wire S4801;
wire S4802;
wire S4803;
wire S4804;
wire S4805;
wire S4806;
wire S4807;
wire S4808;
wire S4809;
wire S4810;
wire S4811;
wire S4812;
wire S4813;
wire S4814;
wire S4815;
wire S4816;
wire S4817;
wire S4818;
wire S4819;
wire S4820;
wire S4821;
wire S4822;
wire S4823;
wire S4824;
wire S4825;
wire S4826;
wire S4827;
wire S4828;
wire S4829;
wire S4830;
wire S4831;
wire S4832;
wire S4833;
wire S4834;
wire S4835;
wire S4836;
wire S4837;
wire S4838;
wire S4839;
wire S4840;
wire S4841;
wire S4842;
wire S4843;
wire S4844;
wire S4845;
wire S4846;
wire S4847;
wire S4848;
wire S4849;
wire S4850;
wire S4851;
wire S4852;
wire S4853;
wire S4854;
wire S4855;
wire S4856;
wire S4857;
wire S4858;
wire S4859;
wire S4860;
wire S4861;
wire S4862;
wire S4863;
wire S4864;
wire S4865;
wire S4866;
wire S4867;
wire S4868;
wire S4869;
wire S4870;
wire S4871;
wire S4872;
wire S4873;
wire S4874;
wire S4875;
wire S4876;
wire S4877;
wire S4878;
wire S4879;
wire S4880;
wire S4881;
wire S4882;
wire S4883;
wire S4884;
wire S4885;
wire S4886;
wire S4887;
wire S4888;
wire S4889;
wire S4890;
wire S4891;
wire S4892;
wire S4893;
wire S4894;
wire S4895;
wire S4896;
wire S4897;
wire S4898;
wire S4899;
wire S4900;
wire S4901;
wire S4902;
wire S4903;
wire S4904;
wire S4905;
wire S4906;
wire S4907;
wire S4908;
wire S4909;
wire S4910;
wire S4911;
wire S4912;
wire S4913;
wire S4914;
wire S4915;
wire S4916;
wire S4917;
wire S4918;
wire S4919;
wire S4920;
wire S4921;
wire S4922;
wire S4923;
wire S4924;
wire S4925;
wire S4926;
wire S4927;
wire S4928;
wire S4929;
wire S4930;
wire S4931;
wire S4932;
wire S4933;
wire S4934;
wire S4935;
wire S4936;
wire S4937;
wire S4938;
wire S4939;
wire S4940;
wire S4941;
wire S4942;
wire S4943;
wire S4944;
wire S4945;
wire S4946;
wire S4947;
wire S4948;
wire S4949;
wire S4950;
wire S4951;
wire S4952;
wire S4953;
wire S4954;
wire S4955;
wire S4956;
wire S4957;
wire S4958;
wire S4959;
wire S4960;
wire S4961;
wire S4962;
wire S4963;
wire S4964;
wire S4965;
wire S4966;
wire S4967;
wire S4968;
wire S4969;
wire S4970;
wire S4971;
wire S4972;
wire S4973;
wire S4974;
wire S4975;
wire S4976;
wire S4977;
wire S4978;
wire S4979;
wire S4980;
wire S4981;
wire S4982;
wire S4983;
wire S4984;
wire S4985;
wire S4986;
wire S4987;
wire S4988;
wire S4989;
wire S4990;
wire S4991;
wire S4992;
wire S4993;
wire S4994;
wire S4995;
wire S4996;
wire S4997;
wire S4998;
wire S4999;
wire S5000;
wire S5001;
wire S5002;
wire S5003;
wire S5004;
wire S5005;
wire S5006;
wire S5007;
wire S5008;
wire S5009;
wire S5010;
wire S5011;
wire S5012;
wire S5013;
wire S5014;
wire S5015;
wire S5016;
wire S5017;
wire S5018;
wire S5019;
wire S5020;
wire S5021;
wire S5022;
wire S5023;
wire S5024;
wire S5025;
wire S5026;
wire S5027;
wire S5028;
wire S5029;
wire S5030;
wire S5031;
wire S5032;
wire S5033;
wire S5034;
wire S5035;
wire S5036;
wire S5037;
wire S5038;
wire S5039;
wire S5040;
wire S5041;
wire S5042;
wire S5043;
wire S5044;
wire S5045;
wire S5046;
wire S5047;
wire S5048;
wire S5049;
wire S5050;
wire S5051;
wire S5052;
wire S5053;
wire S5054;
wire S5055;
wire S5056;
wire S5057;
wire S5058;
wire S5059;
wire S5060;
wire S5061;
wire S5062;
wire S5063;
wire S5064;
wire S5065;
wire S5066;
wire S5067;
wire S5068;
wire S5069;
wire S5070;
wire S5071;
wire S5072;
wire S5073;
wire S5074;
wire S5075;
wire S5076;
wire S5077;
wire S5078;
wire S5079;
wire S5080;
wire S5081;
wire S5082;
wire S5083;
wire S5084;
wire S5085;
wire S5086;
wire S5087;
wire S5088;
wire S5089;
wire S5090;
wire S5091;
wire S5092;
wire S5093;
wire S5094;
wire S5095;
wire S5096;
wire S5097;
wire S5098;
wire S5099;
wire S5100;
wire S5101;
wire S5102;
wire S5103;
wire S5104;
wire S5105;
wire S5106;
wire S5107;
wire S5108;
wire S5109;
wire S5110;
wire S5111;
wire S5112;
wire S5113;
wire S5114;
wire S5115;
wire S5116;
wire S5117;
wire S5118;
wire S5119;
wire S5120;
wire S5121;
wire S5122;
wire S5123;
wire S5124;
wire S5125;
wire S5126;
wire S5127;
wire S5128;
wire S5129;
wire S5130;
wire S5131;
wire S5132;
wire S5133;
wire S5134;
wire S5135;
wire S5136;
wire S5137;
wire S5138;
wire S5139;
wire S5140;
wire S5141;
wire S5142;
wire S5143;
wire S5144;
wire S5145;
wire S5146;
wire S5147;
wire S5148;
wire S5149;
wire S5150;
wire S5151;
wire S5152;
wire S5153;
wire S5154;
wire S5155;
wire S5156;
wire S5157;
wire S5158;
wire S5159;
wire S5160;
wire S5161;
wire S5162;
wire S5163;
wire S5164;
wire S5165;
wire S5166;
wire S5167;
wire S5168;
wire S5169;
wire S5170;
wire S5171;
wire S5172;
wire S5173;
wire S5174;
wire S5175;
wire S5176;
wire S5177;
wire S5178;
wire S5179;
wire S5180;
wire S5181;
wire S5182;
wire S5183;
wire S5184;
wire S5185;
wire S5186;
wire S5187;
wire S5188;
wire S5189;
wire S5190;
wire S5191;
wire S5192;
wire S5193;
wire S5194;
wire S5195;
wire S5196;
wire S5197;
wire S5198;
wire S5199;
wire S5200;
wire S5201;
wire S5202;
wire S5203;
wire S5204;
wire S5205;
wire S5206;
wire S5207;
wire S5208;
wire S5209;
wire S5210;
wire S5211;
wire S5212;
wire S5213;
wire S5214;
wire S5215;
wire S5216;
wire S5217;
wire S5218;
wire S5219;
wire S5220;
wire S5221;
wire S5222;
wire S5223;
wire S5224;
wire S5225;
wire S5226;
wire S5227;
wire S5228;
wire S5229;
wire S5230;
wire S5231;
wire S5232;
wire S5233;
wire S5234;
wire S5235;
wire S5236;
wire S5237;
wire S5238;
wire S5239;
wire S5240;
wire S5241;
wire S5242;
wire S5243;
wire S5244;
wire S5245;
wire S5246;
wire S5247;
wire S5248;
wire S5249;
wire S5250;
wire S5251;
wire S5252;
wire S5253;
wire S5254;
wire S5255;
wire S5256;
wire S5257;
wire S5258;
wire S5259;
wire S5260;
wire S5261;
wire S5262;
wire S5263;
wire S5264;
wire S5265;
wire S5266;
wire S5267;
wire S5268;
wire S5269;
wire S5270;
wire S5271;
wire S5272;
wire S5273;
wire S5274;
wire S5275;
wire S5276;
wire S5277;
wire S5278;
wire S5279;
wire S5280;
wire S5281;
wire S5282;
wire S5283;
wire S5284;
wire S5285;
wire S5286;
wire S5287;
wire S5288;
wire S5289;
wire S5290;
wire S5291;
wire S5292;
wire S5293;
wire S5294;
wire S5295;
wire S5296;
wire S5297;
wire S5298;
wire S5299;
wire S5300;
wire S5301;
wire S5302;
wire S5303;
wire S5304;
wire S5305;
wire S5306;
wire S5307;
wire S5308;
wire S5309;
wire S5310;
wire S5311;
wire S5312;
wire S5313;
wire S5314;
wire S5315;
wire S5316;
wire S5317;
wire S5318;
wire S5319;
wire S5320;
wire S5321;
wire S5322;
wire S5323;
wire S5324;
wire S5325;
wire S5326;
wire S5327;
wire S5328;
wire S5329;
wire S5330;
wire S5331;
wire S5332;
wire S5333;
wire S5334;
wire S5335;
wire S5336;
wire S5337;
wire S5338;
wire S5339;
wire S5340;
wire S5341;
wire S5342;
wire S5343;
wire S5344;
wire S5345;
wire S5346;
wire S5347;
wire S5348;
wire S5349;
wire S5350;
wire S5351;
wire S5352;
wire S5353;
wire S5354;
wire S5355;
wire S5356;
wire S5357;
wire S5358;
wire S5359;
wire S5360;
wire S5361;
wire S5362;
wire S5363;
wire S5364;
wire S5365;
wire S5366;
wire S5367;
wire S5368;
wire S5369;
wire S5370;
wire S5371;
wire S5372;
wire S5373;
wire S5374;
wire S5375;
wire S5376;
wire S5377;
wire S5378;
wire S5379;
wire S5380;
wire S5381;
wire S5382;
wire S5383;
wire S5384;
wire S5385;
wire S5386;
wire S5387;
wire S5388;
wire S5389;
wire S5390;
wire S5391;
wire S5392;
wire S5393;
wire S5394;
wire S5395;
wire S5396;
wire S5397;
wire S5398;
wire S5399;
wire S5400;
wire S5401;
wire S5402;
wire S5403;
wire S5404;
wire S5405;
wire S5406;
wire S5407;
wire S5408;
wire S5409;
wire S5410;
wire S5411;
wire S5412;
wire S5413;
wire S5414;
wire S5415;
wire S5416;
wire S5417;
wire S5418;
wire S5419;
wire S5420;
wire S5421;
wire S5422;
wire S5423;
wire S5424;
wire S5425;
wire S5426;
wire S5427;
wire S5428;
wire S5429;
wire S5430;
wire S5431;
wire S5432;
wire S5433;
wire S5434;
wire S5435;
wire S5436;
wire S5437;
wire S5438;
wire S5439;
wire S5440;
wire S5441;
wire S5442;
wire S5443;
wire S5444;
wire S5445;
wire S5446;
wire S5447;
wire S5448;
wire S5449;
wire S5450;
wire S5451;
wire S5452;
wire S5453;
wire S5454;
wire S5455;
wire S5456;
wire S5457;
wire S5458;
wire S5459;
wire S5460;
wire S5461;
wire S5462;
wire S5463;
wire S5464;
wire S5465;
wire S5466;
wire S5467;
wire S5468;
wire S5469;
wire S5470;
wire S5471;
wire S5472;
wire S5473;
wire S5474;
wire S5475;
wire S5476;
wire S5477;
wire S5478;
wire S5479;
wire S5480;
wire S5481;
wire S5482;
wire S5483;
wire S5484;
wire S5485;
wire S5486;
wire S5487;
wire S5488;
wire S5489;
wire S5490;
wire S5491;
wire S5492;
wire S5493;
wire S5494;
wire S5495;
wire S5496;
wire S5497;
wire S5498;
wire S5499;
wire S5500;
wire S5501;
wire S5502;
wire S5503;
wire S5504;
wire S5505;
wire S5506;
wire S5507;
wire S5508;
wire S5509;
wire S5510;
wire S5511;
wire S5512;
wire S5513;
wire S5514;
wire S5515;
wire S5516;
wire S5517;
wire S5518;
wire S5519;
wire S5520;
wire S5521;
wire S5522;
wire S5523;
wire S5524;
wire S5525;
wire S5526;
wire S5527;
wire S5528;
wire S5529;
wire S5530;
wire S5531;
wire S5532;
wire S5533;
wire S5534;
wire S5535;
wire S5536;
wire S5537;
wire S5538;
wire S5539;
wire S5540;
wire S5541;
wire S5542;
wire S5543;
wire S5544;
wire S5545;
wire S5546;
wire S5547;
wire S5548;
wire S5549;
wire S5550;
wire S5551;
wire S5552;
wire S5553;
wire S5554;
wire S5555;
wire S5556;
wire S5557;
wire S5558;
wire S5559;
wire S5560;
wire S5561;
wire S5562;
wire S5563;
wire S5564;
wire S5565;
wire S5566;
wire S5567;
wire S5568;
wire S5569;
wire S5570;
wire S5571;
wire S5572;
wire S5573;
wire S5574;
wire S5575;
wire S5576;
wire S5577;
wire S5578;
wire S5579;
wire S5580;
wire S5581;
wire S5582;
wire S5583;
wire S5584;
wire S5585;
wire S5586;
wire S5587;
wire S5588;
wire S5589;
wire S5590;
wire S5591;
wire S5592;
wire S5593;
wire S5594;
wire S5595;
wire S5596;
wire S5597;
wire S5598;
wire S5599;
wire S5600;
wire S5601;
wire S5602;
wire S5603;
wire S5604;
wire S5605;
wire S5606;
wire S5607;
wire S5608;
wire S5609;
wire S5610;
wire S5611;
wire S5612;
wire S5613;
wire S5614;
wire S5615;
wire S5616;
wire S5617;
wire S5618;
wire S5619;
wire S5620;
wire S5621;
wire S5622;
wire S5623;
wire S5624;
wire S5625;
wire S5626;
wire S5627;
wire S5628;
wire S5629;
wire S5630;
wire S5631;
wire S5632;
wire S5633;
wire S5634;
wire S5635;
wire S5636;
wire S5637;
wire S5638;
wire S5639;
wire S5640;
wire S5641;
wire S5642;
wire S5643;
wire S5644;
wire S5645;
wire S5646;
wire S5647;
wire S5648;
wire S5649;
wire S5650;
wire S5651;
wire S5652;
wire S5653;
wire S5654;
wire S5655;
wire S5656;
wire S5657;
wire S5658;
wire S5659;
wire S5660;
wire S5661;
wire S5662;
wire S5663;
wire S5664;
wire S5665;
wire S5666;
wire S5667;
wire S5668;
wire S5669;
wire S5670;
wire S5671;
wire S5672;
wire S5673;
wire S5674;
wire S5675;
wire S5676;
wire S5677;
wire S5678;
wire S5679;
wire S5680;
wire S5681;
wire S5682;
wire S5683;
wire S5684;
wire S5685;
wire S5686;
wire S5687;
wire S5688;
wire S5689;
wire S5690;
wire S5691;
wire S5692;
wire S5693;
wire S5694;
wire S5695;
wire S5696;
wire S5697;
wire S5698;
wire S5699;
wire S5700;
wire S5701;
wire S5702;
wire S5703;
wire S5704;
wire S5705;
wire S5706;
wire S5707;
wire S5708;
wire S5709;
wire S5710;
wire S5711;
wire S5712;
wire S5713;
wire S5714;
wire S5715;
wire S5716;
wire S5717;
wire S5718;
wire S5719;
wire S5720;
wire S5721;
wire S5722;
wire S5723;
wire S5724;
wire S5725;
wire S5726;
wire S5727;
wire S5728;
wire S5729;
wire S5730;
wire S5731;
wire S5732;
wire S5733;
wire S5734;
wire S5735;
wire S5736;
wire S5737;
wire S5738;
wire S5739;
wire S5740;
wire S5741;
wire S5742;
wire S5743;
wire S5744;
wire S5745;
wire S5746;
wire S5747;
wire S5748;
wire S5749;
wire S5750;
wire S5751;
wire S5752;
wire S5753;
wire S5754;
wire S5755;
wire S5756;
wire S5757;
wire S5758;
wire S5759;
wire S5760;
wire S5761;
wire S5762;
wire S5763;
wire S5764;
wire S5765;
wire S5766;
wire S5767;
wire S5768;
wire S5769;
wire S5770;
wire S5771;
wire S5772;
wire S5773;
wire S5774;
wire S5775;
wire S5776;
wire S5777;
wire S5778;
wire S5779;
wire S5780;
wire S5781;
wire S5782;
wire S5783;
wire S5784;
wire S5785;
wire S5786;
wire S5787;
wire S5788;
wire S5789;
wire S5790;
wire S5791;
wire S5792;
wire S5793;
wire S5794;
wire S5795;
wire S5796;
wire S5797;
wire S5798;
wire S5799;
wire S5800;
wire S5801;
wire S5802;
wire S5803;
wire S5804;
wire S5805;
wire S5806;
wire S5807;
wire S5808;
wire S5809;
wire S5810;
wire S5811;
wire S5812;
wire S5813;
wire S5814;
wire S5815;
wire S5816;
wire S5817;
wire S5818;
wire S5819;
wire S5820;
wire S5821;
wire S5822;
wire S5823;
wire S5824;
wire S5825;
wire S5826;
wire S5827;
wire S5828;
wire S5829;
wire S5830;
wire S5831;
wire S5832;
wire S5833;
wire S5834;
wire S5835;
wire S5836;
wire S5837;
wire S5838;
wire S5839;
wire S5840;
wire S5841;
wire S5842;
wire S5843;
wire S5844;
wire S5845;
wire S5846;
wire S5847;
wire S5848;
wire S5849;
wire S5850;
wire S5851;
wire S5852;
wire S5853;
wire S5854;
wire S5855;
wire S5856;
wire S5857;
wire S5858;
wire S5859;
wire S5860;
wire S5861;
wire S5862;
wire S5863;
wire S5864;
wire S5865;
wire S5866;
wire S5867;
wire S5868;
wire S5869;
wire S5870;
wire S5871;
wire S5872;
wire S5873;
wire S5874;
wire S5875;
wire S5876;
wire S5877;
wire S5878;
wire S5879;
wire S5880;
wire S5881;
wire S5882;
wire S5883;
wire S5884;
wire S5885;
wire S5886;
wire S5887;
wire S5888;
wire S5889;
wire S5890;
wire S5891;
wire S5892;
wire S5893;
wire S5894;
wire S5895;
wire S5896;
wire S5897;
wire S5898;
wire S5899;
wire S5900;
wire S5901;
wire S5902;
wire S5903;
wire S5904;
wire S5905;
wire S5906;
wire S5907;
wire S5908;
wire S5909;
wire S5910;
wire S5911;
wire S5912;
wire S5913;
wire S5914;
wire S5915;
wire S5916;
wire S5917;
wire S5918;
wire S5919;
wire S5920;
wire S5921;
wire S5922;
wire S5923;
wire S5924;
wire S5925;
wire S5926;
wire S5927;
wire S5928;
wire S5929;
wire S5930;
wire S5931;
wire S5932;
wire S5933;
wire S5934;
wire S5935;
wire S5936;
wire S5937;
wire S5938;
wire S5939;
wire S5940;
wire S5941;
wire S5942;
wire S5943;
wire S5944;
wire S5945;
wire S5946;
wire S5947;
wire S5948;
wire S5949;
wire S5950;
wire S5951;
wire S5952;
wire S5953;
wire S5954;
wire S5955;
wire S5956;
wire S5957;
wire S5958;
wire S5959;
wire S5960;
wire S5961;
wire S5962;
wire S5963;
wire S5964;
wire S5965;
wire S5966;
wire S5967;
wire S5968;
wire S5969;
wire S5970;
wire S5971;
wire S5972;
wire S5973;
wire S5974;
wire S5975;
wire S5976;
wire S5977;
wire S5978;
wire S5979;
wire S5980;
wire S5981;
wire S5982;
wire S5983;
wire S5984;
wire S5985;
wire S5986;
wire S5987;
wire S5988;
wire S5989;
wire S5990;
wire S5991;
wire S5992;
wire S5993;
wire S5994;
wire S5995;
wire S5996;
wire S5997;
wire S5998;
wire S5999;
wire S6000;
wire S6001;
wire S6002;
wire S6003;
wire S6004;
wire S6005;
wire S6006;
wire S6007;
wire S6008;
wire S6009;
wire S6010;
wire S6011;
wire S6012;
wire S6013;
wire S6014;
wire S6015;
wire S6016;
wire S6017;
wire S6018;
wire S6019;
wire S6020;
wire S6021;
wire S6022;
wire S6023;
wire S6024;
wire S6025;
wire S6026;
wire S6027;
wire S6028;
wire S6029;
wire S6030;
wire S6031;
wire S6032;
wire S6033;
wire S6034;
wire S6035;
wire S6036;
wire S6037;
wire S6038;
wire S6039;
wire S6040;
wire S6041;
wire S6042;
wire S6043;
wire S6044;
wire S6045;
wire S6046;
wire S6047;
wire S6048;
wire S6049;
wire S6050;
wire S6051;
wire S6052;
wire S6053;
wire S6054;
wire S6055;
wire S6056;
wire S6057;
wire S6058;
wire S6059;
wire S6060;
wire S6061;
wire S6062;
wire S6063;
wire S6064;
wire S6065;
wire S6066;
wire S6067;
wire S6068;
wire S6069;
wire S6070;
wire S6071;
wire S6072;
wire S6073;
wire S6074;
wire S6075;
wire S6076;
wire S6077;
wire S6078;
wire S6079;
wire S6080;
wire S6081;
wire S6082;
wire S6083;
wire S6084;
wire S6085;
wire S6086;
wire S6087;
wire S6088;
wire S6089;
wire S6090;
wire S6091;
wire S6092;
wire S6093;
wire S6094;
wire S6095;
wire S6096;
wire S6097;
wire S6098;
wire S6099;
wire S6100;
wire S6101;
wire S6102;
wire S6103;
wire S6104;
wire S6105;
wire S6106;
wire S6107;
wire S6108;
wire S6109;
wire S6110;
wire S6111;
wire S6112;
wire S6113;
wire S6114;
wire S6115;
wire S6116;
wire S6117;
wire S6118;
wire S6119;
wire S6120;
wire S6121;
wire S6122;
wire S6123;
wire S6124;
wire S6125;
wire S6126;
wire S6127;
wire S6128;
wire S6129;
wire S6130;
wire S6131;
wire S6132;
wire S6133;
wire S6134;
wire S6135;
wire S6136;
wire S6137;
wire S6138;
wire S6139;
wire S6140;
wire S6141;
wire S6142;
wire S6143;
wire S6144;
wire S6145;
wire S6146;
wire S6147;
wire S6148;
wire S6149;
wire S6150;
wire S6151;
wire S6152;
wire S6153;
wire S6154;
wire S6155;
wire S6156;
wire S6157;
wire S6158;
wire S6159;
wire S6160;
wire S6161;
wire S6162;
wire S6163;
wire S6164;
wire S6165;
wire S6166;
wire S6167;
wire S6168;
wire S6169;
wire S6170;
wire S6171;
wire S6172;
wire S6173;
wire S6174;
wire S6175;
wire S6176;
wire S6177;
wire S6178;
wire S6179;
wire S6180;
wire S6181;
wire S6182;
wire S6183;
wire S6184;
wire S6185;
wire S6186;
wire S6187;
wire S6188;
wire S6189;
wire S6190;
wire S6191;
wire S6192;
wire S6193;
wire S6194;
wire S6195;
wire S6196;
wire S6197;
wire S6198;
wire S6199;
wire S6200;
wire S6201;
wire S6202;
wire S6203;
wire S6204;
wire S6205;
wire S6206;
wire S6207;
wire S6208;
wire S6209;
wire S6210;
wire S6211;
wire S6212;
wire S6213;
wire S6214;
wire S6215;
wire S6216;
wire S6217;
wire S6218;
wire S6219;
wire S6220;
wire S6221;
wire S6222;
wire S6223;
wire S6224;
wire S6225;
wire S6226;
wire S6227;
wire S6228;
wire S6229;
wire S6230;
wire S6231;
wire S6232;
wire S6233;
wire S6234;
wire S6235;
wire S6236;
wire S6237;
wire S6238;
wire S6239;
wire S6240;
wire S6241;
wire S6242;
wire S6243;
wire S6244;
wire S6245;
wire S6246;
wire S6247;
wire S6248;
wire S6249;
wire S6250;
wire S6251;
wire S6252;
wire S6253;
wire S6254;
wire S6255;
wire S6256;
wire S6257;
wire S6258;
wire S6259;
wire S6260;
wire S6261;
wire S6262;
wire S6263;
wire S6264;
wire S6265;
wire S6266;
wire S6267;
wire S6268;
wire S6269;
wire S6270;
wire S6271;
wire S6272;
wire S6273;
wire S6274;
wire S6275;
wire S6276;
wire S6277;
wire S6278;
wire S6279;
wire S6280;
wire S6281;
wire S6282;
wire S6283;
wire S6284;
wire S6285;
wire S6286;
wire S6287;
wire S6288;
wire S6289;
wire S6290;
wire S6291;
wire S6292;
wire S6293;
wire S6294;
wire S6295;
wire S6296;
wire S6297;
wire S6298;
wire S6299;
wire S6300;
wire S6301;
wire S6302;
wire S6303;
wire S6304;
wire S6305;
wire S6306;
wire S6307;
wire S6308;
wire S6309;
wire S6310;
wire S6311;
wire S6312;
wire S6313;
wire S6314;
wire S6315;
wire S6316;
wire S6317;
wire S6318;
wire S6319;
wire S6320;
wire S6321;
wire S6322;
wire S6323;
wire S6324;
wire S6325;
wire S6326;
wire S6327;
wire S6328;
wire S6329;
wire S6330;
wire S6331;
wire S6332;
wire S6333;
wire S6334;
wire S6335;
wire S6336;
wire S6337;
wire S6338;
wire S6339;
wire S6340;
wire S6341;
wire S6342;
wire S6343;
wire S6344;
wire S6345;
wire S6346;
wire S6347;
wire S6348;
wire S6349;
wire S6350;
wire S6351;
wire S6352;
wire S6353;
wire S6354;
wire S6355;
wire S6356;
wire S6357;
wire S6358;
wire S6359;
wire S6360;
wire S6361;
wire S6362;
wire S6363;
wire S6364;
wire S6365;
wire S6366;
wire S6367;
wire S6368;
wire S6369;
wire S6370;
wire S6371;
wire S6372;
wire S6373;
wire S6374;
wire S6375;
wire S6376;
wire S6377;
wire S6378;
wire S6379;
wire S6380;
wire S6381;
wire S6382;
wire S6383;
wire S6384;
wire S6385;
wire S6386;
wire S6387;
wire S6388;
wire S6389;
wire S6390;
wire S6391;
wire S6392;
wire S6393;
wire S6394;
wire S6395;
wire S6396;
wire S6397;
wire S6398;
wire S6399;
wire S6400;
wire S6401;
wire S6402;
wire S6403;
wire S6404;
wire S6405;
wire S6406;
wire S6407;
wire S6408;
wire S6409;
wire S6410;
wire S6411;
wire S6412;
wire S6413;
wire S6414;
wire S6415;
wire S6416;
wire S6417;
wire S6418;
wire S6419;
wire S6420;
wire S6421;
wire S6422;
wire S6423;
wire S6424;
wire S6425;
wire S6426;
wire S6427;
wire S6428;
wire S6429;
wire S6430;
wire S6431;
wire S6432;
wire S6433;
wire S6434;
wire S6435;
wire S6436;
wire S6437;
wire S6438;
wire S6439;
wire S6440;
wire S6441;
wire S6442;
wire S6443;
wire S6444;
wire S6445;
wire S6446;
wire S6447;
wire S6448;
wire S6449;
wire S6450;
wire S6451;
wire S6452;
wire S6453;
wire S6454;
wire S6455;
wire S6456;
wire S6457;
wire S6458;
wire S6459;
wire S6460;
wire S6461;
wire S6462;
wire S6463;
wire S6464;
wire S6465;
wire S6466;
wire S6467;
wire S6468;
wire S6469;
wire S6470;
wire S6471;
wire S6472;
wire S6473;
wire S6474;
wire S6475;
wire S6476;
wire S6477;
wire S6478;
wire S6479;
wire S6480;
wire S6481;
wire S6482;
wire S6483;
wire S6484;
wire S6485;
wire S6486;
wire S6487;
wire S6488;
wire S6489;
wire S6490;
wire S6491;
wire S6492;
wire S6493;
wire S6494;
wire S6495;
wire S6496;
wire S6497;
wire S6498;
wire S6499;
wire S6500;
wire S6501;
wire S6502;
wire S6503;
wire S6504;
wire S6505;
wire S6506;
wire S6507;
wire S6508;
wire S6509;
wire S6510;
wire S6511;
wire S6512;
wire S6513;
wire S6514;
wire S6515;
wire S6516;
wire S6517;
wire S6518;
wire S6519;
wire S6520;
wire S6521;
wire S6522;
wire S6523;
wire S6524;
wire S6525;
wire S6526;
wire S6527;
wire S6528;
wire S6529;
wire S6530;
wire S6531;
wire S6532;
wire S6533;
wire S6534;
wire S6535;
wire S6536;
wire S6537;
wire S6538;
wire S6539;
wire S6540;
wire S6541;
wire S6542;
wire S6543;
wire S6544;
wire S6545;
wire S6546;
wire S6547;
wire S6548;
wire S6549;
wire S6550;
wire S6551;
wire S6552;
wire S6553;
wire S6554;
wire S6555;
wire S6556;
wire S6557;
wire S6558;
wire S6559;
wire S6560;
wire S6561;
wire S6562;
wire S6563;
wire S6564;
wire S6565;
wire S6566;
wire S6567;
wire S6568;
wire S6569;
wire S6570;
wire S6571;
wire S6572;
wire S6573;
wire S6574;
wire S6575;
wire S6576;
wire S6577;
wire S6578;
wire S6579;
wire S6580;
wire S6581;
wire S6582;
wire S6583;
wire S6584;
wire S6585;
wire S6586;
wire S6587;
wire S6588;
wire S6589;
wire S6590;
wire S6591;
wire S6592;
wire S6593;
wire S6594;
wire S6595;
wire S6596;
wire S6597;
wire S6598;
wire S6599;
wire S6600;
wire S6601;
wire S6602;
wire S6603;
wire S6604;
wire S6605;
wire S6606;
wire S6607;
wire S6608;
wire S6609;
wire S6610;
wire S6611;
wire S6612;
wire S6613;
wire S6614;
wire S6615;
wire S6616;
wire S6617;
wire S6618;
wire S6619;
wire S6620;
wire S6621;
wire S6622;
wire S6623;
wire S6624;
wire S6625;
wire S6626;
wire S6627;
wire S6628;
wire S6629;
wire S6630;
wire S6631;
wire S6632;
wire S6633;
wire S6634;
wire S6635;
wire S6636;
wire S6637;
wire S6638;
wire S6639;
wire S6640;
wire S6641;
wire S6642;
wire S6643;
wire S6644;
wire S6645;
wire S6646;
wire S6647;
wire S6648;
wire S6649;
wire S6650;
wire S6651;
wire S6652;
wire S6653;
wire S6654;
wire S6655;
wire S6656;
wire S6657;
wire S6658;
wire S6659;
wire S6660;
wire S6661;
wire S6662;
wire S6663;
wire S6664;
wire S6665;
wire S6666;
wire S6667;
wire S6668;
wire S6669;
wire S6670;
wire S6671;
wire S6672;
wire S6673;
wire S6674;
wire S6675;
wire S6676;
wire S6677;
wire S6678;
wire S6679;
wire S6680;
wire S6681;
wire S6682;
wire S6683;
wire S6684;
wire S6685;
wire S6686;
wire S6687;
wire S6688;
wire S6689;
wire S6690;
wire S6691;
wire S6692;
wire S6693;
wire S6694;
wire S6695;
wire S6696;
wire S6697;
wire S6698;
wire S6699;
wire S6700;
wire S6701;
wire S6702;
wire S6703;
wire S6704;
wire S6705;
wire S6706;
wire S6707;
wire S6708;
wire S6709;
wire S6710;
wire S6711;
wire S6712;
wire S6713;
wire S6714;
wire S6715;
wire S6716;
wire S6717;
wire S6718;
wire S6719;
wire S6720;
wire S6721;
wire S6722;
wire S6723;
wire S6724;
wire S6725;
wire S6726;
wire S6727;
wire S6728;
wire S6729;
wire S6730;
wire S6731;
wire S6732;
wire S6733;
wire S6734;
wire S6735;
wire S6736;
wire S6737;
wire S6738;
wire S6739;
wire S6740;
wire S6741;
wire S6742;
wire S6743;
wire S6744;
wire S6745;
wire S6746;
wire S6747;
wire S6748;
wire S6749;
wire S6750;
wire S6751;
wire S6752;
wire S6753;
wire S6754;
wire S6755;
wire S6756;
wire S6757;
wire S6758;
wire S6759;
wire S6760;
wire S6761;
wire S6762;
wire S6763;
wire S6764;
wire S6765;
wire S6766;
wire S6767;
wire S6768;
wire S6769;
wire S6770;
wire S6771;
wire S6772;
wire S6773;
wire S6774;
wire S6775;
wire S6776;
wire S6777;
wire S6778;
wire S6779;
wire S6780;
wire S6781;
wire S6782;
wire S6783;
wire S6784;
wire S6785;
wire S6786;
wire S6787;
wire S6788;
wire S6789;
wire S6790;
wire S6791;
wire S6792;
wire S6793;
wire S6794;
wire S6795;
wire S6796;
wire S6797;
wire S6798;
wire S6799;
wire S6800;
wire S6801;
wire S6802;
wire S6803;
wire S6804;
wire S6805;
wire S6806;
wire S6807;
wire S6808;
wire S6809;
wire S6810;
wire S6811;
wire S6812;
wire S6813;
wire S6814;
wire S6815;
wire S6816;
wire S6817;
wire S6818;
wire S6819;
wire S6820;
wire S6821;
wire S6822;
wire S6823;
wire S6824;
wire S6825;
wire S6826;
wire S6827;
wire S6828;
wire S6829;
wire S6830;
wire S6831;
wire S6832;
wire S6833;
wire S6834;
wire S6835;
wire S6836;
wire S6837;
wire S6838;
wire S6839;
wire S6840;
wire S6841;
wire S6842;
wire S6843;
wire S6844;
wire S6845;
wire S6846;
wire S6847;
wire S6848;
wire S6849;
wire S6850;
wire S6851;
wire S6852;
wire S6853;
wire S6854;
wire S6855;
wire S6856;
wire S6857;
wire S6858;
wire S6859;
wire S6860;
wire S6861;
wire S6862;
wire S6863;
wire S6864;
wire S6865;
wire S6866;
wire S6867;
wire S6868;
wire S6869;
wire S6870;
wire S6871;
wire S6872;
wire S6873;
wire S6874;
wire S6875;
wire S6876;
wire S6877;
wire S6878;
wire S6879;
wire S6880;
wire S6881;
wire S6882;
wire S6883;
wire S6884;
wire S6885;
wire S6886;
wire S6887;
wire S6888;
wire S6889;
wire S6890;
wire S6891;
wire S6892;
wire S6893;
wire S6894;
wire S6895;
wire S6896;
wire S6897;
wire S6898;
wire S6899;
wire S6900;
wire S6901;
wire S6902;
wire S6903;
wire S6904;
wire S6905;
wire S6906;
wire S6907;
wire S6908;
wire S6909;
wire S6910;
wire S6911;
wire S6912;
wire S6913;
wire S6914;
wire S6915;
wire S6916;
wire S6917;
wire S6918;
wire S6919;
wire S6920;
wire S6921;
wire S6922;
wire S6923;
wire S6924;
wire S6925;
wire S6926;
wire S6927;
wire S6928;
wire S6929;
wire S6930;
wire S6931;
wire S6932;
wire S6933;
wire S6934;
wire S6935;
wire S6936;
wire S6937;
wire S6938;
wire S6939;
wire S6940;
wire S6941;
wire S6942;
wire S6943;
wire S6944;
wire S6945;
wire S6946;
wire S6947;
wire S6948;
wire S6949;
wire S6950;
wire S6951;
wire S6952;
wire S6953;
wire S6954;
wire S6955;
wire S6956;
wire S6957;
wire S6958;
wire S6959;
wire S6960;
wire S6961;
wire S6962;
wire S6963;
wire S6964;
wire S6965;
wire S6966;
wire S6967;
wire S6968;
wire S6969;
wire S6970;
wire S6971;
wire S6972;
wire S6973;
wire S6974;
wire S6975;
wire S6976;
wire S6977;
wire S6978;
wire S6979;
wire S6980;
wire S6981;
wire S6982;
wire S6983;
wire S6984;
wire S6985;
wire S6986;
wire S6987;
wire S6988;
wire S6989;
wire S6990;
wire S6991;
wire S6992;
wire S6993;
wire S6994;
wire S6995;
wire S6996;
wire S6997;
wire S6998;
wire S6999;
wire S7000;
wire S7001;
wire S7002;
wire S7003;
wire S7004;
wire S7005;
wire S7006;
wire S7007;
wire S7008;
wire S7009;
wire S7010;
wire S7011;
wire S7012;
wire S7013;
wire S7014;
wire S7015;
wire S7016;
wire S7017;
wire S7018;
wire S7019;
wire S7020;
wire S7021;
wire S7022;
wire S7023;
wire S7024;
wire S7025;
wire S7026;
wire S7027;
wire S7028;
wire S7029;
wire S7030;
wire S7031;
wire S7032;
wire S7033;
wire S7034;
wire S7035;
wire S7036;
wire S7037;
wire S7038;
wire S7039;
wire S7040;
wire S7041;
wire S7042;
wire S7043;
wire S7044;
wire S7045;
wire S7046;
wire S7047;
wire S7048;
wire S7049;
wire S7050;
wire S7051;
wire S7052;
wire S7053;
wire S7054;
wire S7055;
wire S7056;
wire S7057;
wire S7058;
wire S7059;
wire S7060;
wire S7061;
wire S7062;
wire S7063;
wire S7064;
wire S7065;
wire S7066;
wire S7067;
wire S7068;
wire S7069;
wire S7070;
wire S7071;
wire S7072;
wire S7073;
wire S7074;
wire S7075;
wire S7076;
wire S7077;
wire S7078;
wire S7079;
wire S7080;
wire S7081;
wire S7082;
wire S7083;
wire S7084;
wire S7085;
wire S7086;
wire S7087;
wire S7088;
wire S7089;
wire S7090;
wire S7091;
wire S7092;
wire S7093;
wire S7094;
wire S7095;
wire S7096;
wire S7097;
wire S7098;
wire S7099;
wire S7100;
wire S7101;
wire S7102;
wire S7103;
wire S7104;
wire S7105;
wire S7106;
wire S7107;
wire S7108;
wire S7109;
wire S7110;
wire S7111;
wire S7112;
wire S7113;
wire S7114;
wire S7115;
wire S7116;
wire S7117;
wire S7118;
wire S7119;
wire S7120;
wire S7121;
wire S7122;
wire S7123;
wire S7124;
wire S7125;
wire S7126;
wire S7127;
wire S7128;
wire S7129;
wire S7130;
wire S7131;
wire S7132;
wire S7133;
wire S7134;
wire S7135;
wire S7136;
wire S7137;
wire S7138;
wire S7139;
wire S7140;
wire S7141;
wire S7142;
wire S7143;
wire S7144;
wire S7145;
wire S7146;
wire S7147;
wire S7148;
wire S7149;
wire S7150;
wire S7151;
wire S7152;
wire S7153;
wire S7154;
wire S7155;
wire S7156;
wire S7157;
wire S7158;
wire S7159;
wire S7160;
wire S7161;
wire S7162;
wire S7163;
wire S7164;
wire S7165;
wire S7166;
wire S7167;
wire S7168;
wire S7169;
wire S7170;
wire S7171;
wire S7172;
wire S7173;
wire S7174;
wire S7175;
wire S7176;
wire S7177;
wire S7178;
wire S7179;
wire S7180;
wire S7181;
wire S7182;
wire S7183;
wire S7184;
wire S7185;
wire S7186;
wire S7187;
wire S7188;
wire S7189;
wire S7190;
wire S7191;
wire S7192;
wire S7193;
wire S7194;
wire S7195;
wire S7196;
wire S7197;
wire S7198;
wire S7199;
wire S7200;
wire S7201;
wire S7202;
wire S7203;
wire S7204;
wire S7205;
wire S7206;
wire S7207;
wire S7208;
wire S7209;
wire S7210;
wire S7211;
wire S7212;
wire S7213;
wire S7214;
wire S7215;
wire S7216;
wire S7217;
wire S7218;
wire S7219;
wire S7220;
wire S7221;
wire S7222;
wire S7223;
wire S7224;
wire S7225;
wire S7226;
wire S7227;
wire S7228;
wire S7229;
wire S7230;
wire S7231;
wire S7232;
wire S7233;
wire S7234;
wire S7235;
wire S7236;
wire S7237;
wire S7238;
wire S7239;
wire S7240;
wire S7241;
wire S7242;
wire S7243;
wire S7244;
wire S7245;
wire S7246;
wire S7247;
wire S7248;
wire S7249;
wire S7250;
wire S7251;
wire S7252;
wire S7253;
wire S7254;
wire S7255;
wire S7256;
wire S7257;
wire S7258;
wire S7259;
wire S7260;
wire S7261;
wire S7262;
wire S7263;
wire S7264;
wire S7265;
wire S7266;
wire S7267;
wire S7268;
wire S7269;
wire S7270;
wire S7271;
wire S7272;
wire S7273;
wire S7274;
wire S7275;
wire S7276;
wire S7277;
wire S7278;
wire S7279;
wire S7280;
wire S7281;
wire S7282;
wire S7283;
wire S7284;
wire S7285;
wire S7286;
wire S7287;
wire S7288;
wire S7289;
wire S7290;
wire S7291;
wire S7292;
wire S7293;
wire S7294;
wire S7295;
wire S7296;
wire S7297;
wire S7298;
wire S7299;
wire S7300;
wire S7301;
wire S7302;
wire S7303;
wire S7304;
wire S7305;
wire S7306;
wire S7307;
wire S7308;
wire S7309;
wire S7310;
wire S7311;
wire S7312;
wire S7313;
wire S7314;
wire S7315;
wire S7316;
wire S7317;
wire S7318;
wire S7319;
wire S7320;
wire S7321;
wire S7322;
wire S7323;
wire S7324;
wire S7325;
wire S7326;
wire S7327;
wire S7328;
wire S7329;
wire S7330;
wire S7331;
wire S7332;
wire S7333;
wire S7334;
wire S7335;
wire S7336;
wire S7337;
wire S7338;
wire S7339;
wire S7340;
wire S7341;
wire S7342;
wire S7343;
wire S7344;
wire S7345;
wire S7346;
wire S7347;
wire S7348;
wire S7349;
wire S7350;
wire S7351;
wire S7352;
wire S7353;
wire S7354;
wire S7355;
wire S7356;
wire S7357;
wire S7358;
wire S7359;
wire S7360;
wire S7361;
wire S7362;
wire S7363;
wire S7364;
wire S7365;
wire S7366;
wire S7367;
wire S7368;
wire S7369;
wire S7370;
wire S7371;
wire S7372;
wire S7373;
wire S7374;
wire S7375;
wire S7376;
wire S7377;
wire S7378;
wire S7379;
wire S7380;
wire S7381;
wire S7382;
wire S7383;
wire S7384;
wire S7385;
wire S7386;
wire S7387;
wire S7388;
wire S7389;
wire S7390;
wire S7391;
wire S7392;
wire S7393;
wire S7394;
wire S7395;
wire S7396;
wire S7397;
wire S7398;
wire S7399;
wire S7400;
wire S7401;
wire S7402;
wire S7403;
wire S7404;
wire S7405;
wire S7406;
wire S7407;
wire S7408;
wire S7409;
wire S7410;
wire S7411;
wire S7412;
wire S7413;
wire S7414;
wire S7415;
wire S7416;
wire S7417;
wire S7418;
wire S7419;
wire S7420;
wire S7421;
wire S7422;
wire S7423;
wire S7424;
wire S7425;
wire S7426;
wire S7427;
wire S7428;
wire S7429;
wire S7430;
wire S7431;
wire S7432;
wire S7433;
wire S7434;
wire S7435;
wire S7436;
wire S7437;
wire S7438;
wire S7439;
wire S7440;
wire S7441;
wire S7442;
wire S7443;
wire S7444;
wire S7445;
wire S7446;
wire S7447;
wire S7448;
wire S7449;
wire S7450;
wire S7451;
wire S7452;
wire S7453;
wire S7454;
wire S7455;
wire S7456;
wire S7457;
wire S7458;
wire S7459;
wire S7460;
wire S7461;
wire S7462;
wire S7463;
wire S7464;
wire S7465;
wire S7466;
wire S7467;
wire S7468;
wire S7469;
wire S7470;
wire S7471;
wire S7472;
wire S7473;
wire S7474;
wire S7475;
wire S7476;
wire S7477;
wire S7478;
wire S7479;
wire S7480;
wire S7481;
wire S7482;
wire S7483;
wire S7484;
wire S7485;
wire S7486;
wire S7487;
wire S7488;
wire S7489;
wire S7490;
wire S7491;
wire S7492;
wire S7493;
wire S7494;
wire S7495;
wire S7496;
wire S7497;
wire S7498;
wire S7499;
wire S7500;
wire S7501;
wire S7502;
wire S7503;
wire S7504;
wire S7505;
wire S7506;
wire S7507;
wire S7508;
wire S7509;
wire S7510;
wire S7511;
wire S7512;
wire S7513;
wire S7514;
wire S7515;
wire S7516;
wire S7517;
wire S7518;
wire S7519;
wire S7520;
wire S7521;
wire S7522;
wire S7523;
wire S7524;
wire S7525;
wire S7526;
wire S7527;
wire S7528;
wire S7529;
wire S7530;
wire S7531;
wire S7532;
wire S7533;
wire S7534;
wire S7535;
wire S7536;
wire S7537;
wire S7538;
wire S7539;
wire S7540;
wire S7541;
wire S7542;
wire S7543;
wire S7544;
wire S7545;
wire S7546;
wire S7547;
wire S7548;
wire S7549;
wire S7550;
wire S7551;
wire S7552;
wire S7553;
wire S7554;
wire S7555;
wire S7556;
wire S7557;
wire S7558;
wire S7559;
wire S7560;
wire S7561;
wire S7562;
wire S7563;
wire S7564;
wire S7565;
wire S7566;
wire S7567;
wire S7568;
wire S7569;
wire S7570;
wire S7571;
wire S7572;
wire S7573;
wire S7574;
wire S7575;
wire S7576;
wire S7577;
wire S7578;
wire S7579;
wire S7580;
wire S7581;
wire S7582;
wire S7583;
wire S7584;
wire S7585;
wire S7586;
wire S7587;
wire S7588;
wire S7589;
wire S7590;
wire S7591;
wire S7592;
wire S7593;
wire S7594;
wire S7595;
wire S7596;
wire S7597;
wire S7598;
wire S7599;
wire S7600;
wire S7601;
wire S7602;
wire S7603;
wire S7604;
wire S7605;
wire S7606;
wire S7607;
wire S7608;
wire S7609;
wire S7610;
wire S7611;
wire S7612;
wire S7613;
wire S7614;
wire S7615;
wire S7616;
wire S7617;
wire S7618;
wire S7619;
wire S7620;
wire S7621;
wire S7622;
wire S7623;
wire S7624;
wire S7625;
wire S7626;
wire S7627;
wire S7628;
wire S7629;
wire S7630;
wire S7631;
wire S7632;
wire S7633;
wire S7634;
wire S7635;
wire S7636;
wire S7637;
wire S7638;
wire S7639;
wire S7640;
wire S7641;
wire S7642;
wire S7643;
wire S7644;
wire S7645;
wire S7646;
wire S7647;
wire S7648;
wire S7649;
wire S7650;
wire S7651;
wire S7652;
wire S7653;
wire S7654;
wire S7655;
wire S7656;
wire S7657;
wire S7658;
wire S7659;
wire S7660;
wire S7661;
wire S7662;
wire S7663;
wire S7664;
wire S7665;
wire S7666;
wire S7667;
wire S7668;
wire S7669;
wire S7670;
wire S7671;
wire S7672;
wire S7673;
wire S7674;
wire S7675;
wire S7676;
wire S7677;
wire S7678;
wire S7679;
wire S7680;
wire S7681;
wire S7682;
wire S7683;
wire S7684;
wire S7685;
wire S7686;
wire S7687;
wire S7688;
wire S7689;
wire S7690;
wire S7691;
wire S7692;
wire S7693;
wire S7694;
wire S7695;
wire S7696;
wire S7697;
wire S7698;
wire S7699;
wire S7700;
wire S7701;
wire S7702;
wire S7703;
wire S7704;
wire S7705;
wire S7706;
wire S7707;
wire S7708;
wire S7709;
wire S7710;
wire S7711;
wire S7712;
wire S7713;
wire S7714;
wire S7715;
wire S7716;
wire S7717;
wire S7718;
wire S7719;
wire S7720;
wire S7721;
wire S7722;
wire S7723;
wire S7724;
wire S7725;
wire S7726;
wire S7727;
wire S7728;
wire S7729;
wire S7730;
wire S7731;
wire S7732;
wire S7733;
wire S7734;
wire S7735;
wire S7736;
wire S7737;
wire S7738;
wire S7739;
wire S7740;
wire S7741;
wire S7742;
wire S7743;
wire S7744;
wire S7745;
wire S7746;
wire S7747;
wire S7748;
wire S7749;
wire S7750;
wire S7751;
wire S7752;
wire S7753;
wire S7754;
wire S7755;
wire S7756;
wire S7757;
wire S7758;
wire S7759;
wire S7760;
wire S7761;
wire S7762;
wire S7763;
wire S7764;
wire S7765;
wire S7766;
wire S7767;
wire S7768;
wire S7769;
wire S7770;
wire S7771;
wire S7772;
wire S7773;
wire S7774;
wire S7775;
wire S7776;
wire S7777;
wire S7778;
wire S7779;
wire S7780;
wire S7781;
wire S7782;
wire S7783;
wire S7784;
wire S7785;
wire S7786;
wire S7787;
wire S7788;
wire S7789;
wire S7790;
wire S7791;
wire S7792;
wire S7793;
wire S7794;
wire S7795;
wire S7796;
wire S7797;
wire S7798;
wire S7799;
wire S7800;
wire S7801;
wire S7802;
wire S7803;
wire S7804;
wire S7805;
wire S7806;
wire S7807;
wire S7808;
wire S7809;
wire S7810;
wire S7811;
wire S7812;
wire S7813;
wire S7814;
wire S7815;
wire S7816;
wire S7817;
wire S7818;
wire S7819;
wire S7820;
wire S7821;
wire S7822;
wire S7823;
wire S7824;
wire S7825;
wire S7826;
wire S7827;
wire S7828;
wire S7829;
wire S7830;
wire S7831;
wire S7832;
wire S7833;
wire S7834;
wire S7835;
wire S7836;
wire S7837;
wire S7838;
wire S7839;
wire S7840;
wire S7841;
wire S7842;
wire S7843;
wire S7844;
wire S7845;
wire S7846;
wire S7847;
wire S7848;
wire S7849;
wire S7850;
wire S7851;
wire S7852;
wire S7853;
wire S7854;
wire S7855;
wire S7856;
wire S7857;
wire S7858;
wire S7859;
wire S7860;
wire S7861;
wire S7862;
wire S7863;
wire S7864;
wire S7865;
wire S7866;
wire S7867;
wire S7868;
wire S7869;
wire S7870;
wire S7871;
wire S7872;
wire S7873;
wire S7874;
wire S7875;
wire S7876;
wire S7877;
wire S7878;
wire S7879;
wire S7880;
wire S7881;
wire S7882;
wire S7883;
wire S7884;
wire S7885;
wire S7886;
wire S7887;
wire S7888;
wire S7889;
wire S7890;
wire S7891;
wire S7892;
wire S7893;
wire S7894;
wire S7895;
wire S7896;
wire S7897;
wire S7898;
wire S7899;
wire S7900;
wire S7901;
wire S7902;
wire S7903;
wire S7904;
wire S7905;
wire S7906;
wire S7907;
wire S7908;
wire S7909;
wire S7910;
wire S7911;
wire S7912;
wire S7913;
wire S7914;
wire S7915;
wire S7916;
wire S7917;
wire S7918;
wire S7919;
wire S7920;
wire S7921;
wire S7922;
wire S7923;
wire S7924;
wire S7925;
wire S7926;
wire S7927;
wire S7928;
wire S7929;
wire S7930;
wire S7931;
wire S7932;
wire S7933;
wire S7934;
wire S7935;
wire S7936;
wire S7937;
wire S7938;
wire S7939;
wire S7940;
wire S7941;
wire S7942;
wire S7943;
wire S7944;
wire S7945;
wire S7946;
wire S7947;
wire S7948;
wire S7949;
wire S7950;
wire S7951;
wire S7952;
wire S7953;
wire S7954;
wire S7955;
wire S7956;
wire S7957;
wire S7958;
wire S7959;
wire S7960;
wire S7961;
wire S7962;
wire S7963;
wire S7964;
wire S7965;
wire S7966;
wire S7967;
wire S7968;
wire S7969;
wire S7970;
wire S7971;
wire S7972;
wire S7973;
wire S7974;
wire S7975;
wire S7976;
wire S7977;
wire S7978;
wire S7979;
wire S7980;
wire S7981;
wire S7982;
wire S7983;
wire S7984;
wire S7985;
wire S7986;
wire S7987;
wire S7988;
wire S7989;
wire S7990;
wire S7991;
wire S7992;
wire S7993;
wire S7994;
wire S7995;
wire S7996;
wire S7997;
wire S7998;
wire S7999;
wire S8000;
wire S8001;
wire S8002;
wire S8003;
wire S8004;
wire S8005;
wire S8006;
wire S8007;
wire S8008;
wire S8009;
wire S8010;
wire S8011;
wire S8012;
wire S8013;
wire S8014;
wire S8015;
wire S8016;
wire S8017;
wire S8018;
wire S8019;
wire S8020;
wire S8021;
wire S8022;
wire S8023;
wire S8024;
wire S8025;
wire S8026;
wire S8027;
wire S8028;
wire S8029;
wire S8030;
wire S8031;
wire S8032;
wire S8033;
wire S8034;
wire S8035;
wire S8036;
wire S8037;
wire S8038;
wire S8039;
wire S8040;
wire S8041;
wire S8042;
wire S8043;
wire S8044;
wire S8045;
wire S8046;
wire S8047;
wire S8048;
wire S8049;
wire S8050;
wire S8051;
wire S8052;
wire S8053;
wire S8054;
wire S8055;
wire S8056;
wire S8057;
wire S8058;
wire S8059;
wire S8060;
wire S8061;
wire S8062;
wire S8063;
wire S8064;
wire S8065;
wire S8066;
wire S8067;
wire S8068;
wire S8069;
wire S8070;
wire S8071;
wire S8072;
wire S8073;
wire S8074;
wire S8075;
wire S8076;
wire S8077;
wire S8078;
wire S8079;
wire S8080;
wire S8081;
wire S8082;
wire S8083;
wire S8084;
wire S8085;
wire S8086;
wire S8087;
wire S8088;
wire S8089;
wire S8090;
wire S8091;
wire S8092;
wire S8093;
wire S8094;
wire S8095;
wire S8096;
wire S8097;
wire S8098;
wire S8099;
wire S8100;
wire S8101;
wire S8102;
wire S8103;
wire S8104;
wire S8105;
wire S8106;
wire S8107;
wire S8108;
wire S8109;
wire S8110;
wire S8111;
wire S8112;
wire S8113;
wire S8114;
wire S8115;
wire S8116;
wire S8117;
wire S8118;
wire S8119;
wire S8120;
wire S8121;
wire S8122;
wire S8123;
wire S8124;
wire S8125;
wire S8126;
wire S8127;
wire S8128;
wire S8129;
wire S8130;
wire S8131;
wire S8132;
wire S8133;
wire S8134;
wire S8135;
wire S8136;
wire S8137;
wire S8138;
wire S8139;
wire S8140;
wire S8141;
wire S8142;
wire S8143;
wire S8144;
wire S8145;
wire S8146;
wire S8147;
wire S8148;
wire S8149;
wire S8150;
wire S8151;
wire S8152;
wire S8153;
wire S8154;
wire S8155;
wire S8156;
wire S8157;
wire S8158;
wire S8159;
wire S8160;
wire S8161;
wire S8162;
wire S8163;
wire S8164;
wire S8165;
wire S8166;
wire S8167;
wire S8168;
wire S8169;
wire S8170;
wire S8171;
wire S8172;
wire S8173;
wire S8174;
wire S8175;
wire S8176;
wire S8177;
wire S8178;
wire S8179;
wire S8180;
wire S8181;
wire S8182;
wire S8183;
wire S8184;
wire S8185;
wire S8186;
wire S8187;
wire S8188;
wire S8189;
wire S8190;
wire S8191;
wire S8192;
wire S8193;
wire S8194;
wire S8195;
wire S8196;
wire S8197;
wire S8198;
wire S8199;
wire S8200;
wire S8201;
wire S8202;
wire S8203;
wire S8204;
wire S8205;
wire S8206;
wire S8207;
wire S8208;
wire S8209;
wire S8210;
wire S8211;
wire S8212;
wire S8213;
wire S8214;
wire S8215;
wire S8216;
wire S8217;
wire S8218;
wire S8219;
wire S8220;
wire S8221;
wire S8222;
wire S8223;
wire S8224;
wire S8225;
wire S8226;
wire S8227;
wire S8228;
wire S8229;
wire S8230;
wire S8231;
wire S8232;
wire S8233;
wire S8234;
wire S8235;
wire S8236;
wire S8237;
wire S8238;
wire S8239;
wire S8240;
wire S8241;
wire S8242;
wire S8243;
wire S8244;
wire S8245;
wire S8246;
wire S8247;
wire S8248;
wire S8249;
wire S8250;
wire S8251;
wire S8252;
wire S8253;
wire S8254;
wire S8255;
wire S8256;
wire S8257;
wire S8258;
wire S8259;
wire S8260;
wire S8261;
wire S8262;
wire S8263;
wire S8264;
wire S8265;
wire S8266;
wire S8267;
wire S8268;
wire S8269;
wire S8270;
wire S8271;
wire S8272;
wire S8273;
wire S8274;
wire S8275;
wire S8276;
wire S8277;
wire S8278;
wire S8279;
wire S8280;
wire S8281;
wire S8282;
wire S8283;
wire S8284;
wire S8285;
wire S8286;
wire S8287;
wire S8288;
wire S8289;
wire S8290;
wire S8291;
wire S8292;
wire S8293;
wire S8294;
wire S8295;
wire S8296;
wire S8297;
wire S8298;
wire S8299;
wire S8300;
wire S8301;
wire S8302;
wire S8303;
wire S8304;
wire S8305;
wire S8306;
wire S8307;
wire S8308;
wire S8309;
wire S8310;
wire S8311;
wire S8312;
wire S8313;
wire S8314;
wire S8315;
wire S8316;
wire S8317;
wire S8318;
wire S8319;
wire S8320;
wire S8321;
wire S8322;
wire S8323;
wire S8324;
wire S8325;
wire S8326;
wire S8327;
wire S8328;
wire S8329;
wire S8330;
wire S8331;
wire S8332;
wire S8333;
wire S8334;
wire S8335;
wire S8336;
wire S8337;
wire S8338;
wire S8339;
wire S8340;
wire S8341;
wire S8342;
wire S8343;
wire S8344;
wire S8345;
wire S8346;
wire S8347;
wire S8348;
wire S8349;
wire S8350;
wire S8351;
wire S8352;
wire S8353;
wire S8354;
wire S8355;
wire S8356;
wire S8357;
wire S8358;
wire S8359;
wire S8360;
wire S8361;
wire S8362;
wire S8363;
wire S8364;
wire S8365;
wire S8366;
wire S8367;
wire S8368;
wire S8369;
wire S8370;
wire S8371;
wire S8372;
wire S8373;
wire S8374;
wire S8375;
wire S8376;
wire S8377;
wire S8378;
wire S8379;
wire S8380;
wire S8381;
wire S8382;
wire S8383;
wire S8384;
wire S8385;
wire S8386;
wire S8387;
wire S8388;
wire S8389;
wire S8390;
wire S8391;
wire S8392;
wire S8393;
wire S8394;
wire S8395;
wire S8396;
wire S8397;
wire S8398;
wire S8399;
wire S8400;
wire S8401;
wire S8402;
wire S8403;
wire S8404;
wire S8405;
wire S8406;
wire S8407;
wire S8408;
wire S8409;
wire S8410;
wire S8411;
wire S8412;
wire S8413;
wire S8414;
wire S8415;
wire S8416;
wire S8417;
wire S8418;
wire S8419;
wire S8420;
wire S8421;
wire S8422;
wire S8423;
wire S8424;
wire S8425;
wire S8426;
wire S8427;
wire S8428;
wire S8429;
wire S8430;
wire S8431;
wire S8432;
wire S8433;
wire S8434;
wire S8435;
wire S8436;
wire S8437;
wire S8438;
wire S8439;
wire S8440;
wire S8441;
wire S8442;
wire S8443;
wire S8444;
wire S8445;
wire S8446;
wire S8447;
wire S8448;
wire S8449;
wire S8450;
wire S8451;
wire S8452;
wire S8453;
wire S8454;
wire S8455;
wire S8456;
wire S8457;
wire S8458;
wire S8459;
wire S8460;
wire S8461;
wire S8462;
wire S8463;
wire S8464;
wire S8465;
wire S8466;
wire S8467;
wire S8468;
wire S8469;
wire S8470;
wire S8471;
wire S8472;
wire S8473;
wire S8474;
wire S8475;
wire S8476;
wire S8477;
wire S8478;
wire S8479;
wire S8480;
wire S8481;
wire S8482;
wire S8483;
wire S8484;
wire S8485;
wire S8486;
wire S8487;
wire S8488;
wire S8489;
wire S8490;
wire S8491;
wire S8492;
wire S8493;
wire S8494;
wire S8495;
wire S8496;
wire S8497;
wire S8498;
wire S8499;
wire S8500;
wire S8501;
wire S8502;
wire S8503;
wire S8504;
wire S8505;
wire S8506;
wire S8507;
wire S8508;
wire S8509;
wire S8510;
wire S8511;
wire S8512;
wire S8513;
wire S8514;
wire S8515;
wire S8516;
wire S8517;
wire S8518;
wire S8519;
wire S8520;
wire S8521;
wire S8522;
wire S8523;
wire S8524;
wire S8525;
wire S8526;
wire S8527;
wire S8528;
wire S8529;
wire S8530;
wire S8531;
wire S8532;
wire S8533;
wire S8534;
wire S8535;
wire S8536;
wire S8537;
wire S8538;
wire S8539;
wire S8540;
wire S8541;
wire S8542;
wire S8543;
wire S8544;
wire S8545;
wire S8546;
wire S8547;
wire S8548;
wire S8549;
wire S8550;
wire S8551;
wire S8552;
wire S8553;
wire S8554;
wire S8555;
wire S8556;
wire S8557;
wire S8558;
wire S8559;
wire S8560;
wire S8561;
wire S8562;
wire S8563;
wire S8564;
wire S8565;
wire S8566;
wire S8567;
wire S8568;
wire S8569;
wire S8570;
wire S8571;
wire S8572;
wire S8573;
wire S8574;
wire S8575;
wire S8576;
wire S8577;
wire S8578;
wire S8579;
wire S8580;
wire S8581;
wire S8582;
wire S8583;
wire S8584;
wire S8585;
wire S8586;
wire S8587;
wire S8588;
wire S8589;
wire S8590;
wire S8591;
wire S8592;
wire S8593;
wire S8594;
wire S8595;
wire S8596;
wire S8597;
wire S8598;
wire S8599;
wire S8600;
wire S8601;
wire S8602;
wire S8603;
wire S8604;
wire S8605;
wire S8606;
wire S8607;
wire S8608;
wire S8609;
wire S8610;
wire S8611;
wire S8612;
wire S8613;
wire S8614;
wire S8615;
wire S8616;
wire S8617;
wire S8618;
wire S8619;
wire S8620;
wire S8621;
wire S8622;
wire S8623;
wire S8624;
wire S8625;
wire S8626;
wire S8627;
wire S8628;
wire S8629;
wire S8630;
wire S8631;
wire S8632;
wire S8633;
wire S8634;
wire S8635;
wire S8636;
wire S8637;
wire S8638;
wire S8639;
wire S8640;
wire S8641;
wire S8642;
wire S8643;
wire S8644;
wire S8645;
wire S8646;
wire S8647;
wire S8648;
wire S8649;
wire S8650;
wire S8651;
wire S8652;
wire S8653;
wire S8654;
wire S8655;
wire S8656;
wire S8657;
wire S8658;
wire S8659;
wire S8660;
wire S8661;
wire S8662;
wire S8663;
wire S8664;
wire S8665;
wire S8666;
wire S8667;
wire S8668;
wire S8669;
wire S8670;
wire S8671;
wire S8672;
wire S8673;
wire S8674;
wire S8675;
wire S8676;
wire S8677;
wire S8678;
wire S8679;
wire S8680;
wire S8681;
wire S8682;
wire S8683;
wire S8684;
wire S8685;
wire S8686;
wire S8687;
wire S8688;
wire S8689;
wire S8690;
wire S8691;
wire S8692;
wire S8693;
wire S8694;
wire S8695;
wire S8696;
wire S8697;
wire S8698;
wire S8699;
wire S8700;
wire S8701;
wire S8702;
wire S8703;
wire S8704;
wire S8705;
wire S8706;
wire S8707;
wire S8708;
wire S8709;
wire S8710;
wire S8711;
wire S8712;
wire S8713;
wire S8714;
wire S8715;
wire S8716;
wire S8717;
wire S8718;
wire S8719;
wire S8720;
wire S8721;
wire S8722;
wire S8723;
wire S8724;
wire S8725;
wire S8726;
wire S8727;
wire S8728;
wire S8729;
wire S8730;
wire S8731;
wire S8732;
wire S8733;
wire S8734;
wire S8735;
wire S8736;
wire S8737;
wire S8738;
wire S8739;
wire S8740;
wire S8741;
wire S8742;
wire S8743;
wire S8744;
wire S8745;
wire S8746;
wire S8747;
wire S8748;
wire S8749;
wire S8750;
wire S8751;
wire S8752;
wire S8753;
wire S8754;
wire S8755;
wire S8756;
wire S8757;
wire S8758;
wire S8759;
wire S8760;
wire S8761;
wire S8762;
wire S8763;
wire S8764;
wire S8765;
wire S8766;
wire S8767;
wire S8768;
wire S8769;
wire S8770;
wire S8771;
wire S8772;
wire S8773;
wire S8774;
wire S8775;
wire S8776;
wire S8777;
wire S8778;
wire S8779;
wire S8780;
wire S8781;
wire S8782;
wire S8783;
wire S8784;
wire S8785;
wire S8786;
wire S8787;
wire S8788;
wire S8789;
wire S8790;
wire S8791;
wire S8792;
wire S8793;
wire S8794;
wire S8795;
wire S8796;
wire S8797;
wire S8798;
wire S8799;
wire S8800;
wire S8801;
wire S8802;
wire S8803;
wire S8804;
wire S8805;
wire S8806;
wire S8807;
wire S8808;
wire S8809;
wire S8810;
wire S8811;
wire S8812;
wire S8813;
wire S8814;
wire S8815;
wire S8816;
wire S8817;
wire S8818;
wire S8819;
wire S8820;
wire S8821;
wire S8822;
wire S8823;
wire S8824;
wire S8825;
wire S8826;
wire S8827;
wire S8828;
wire S8829;
wire S8830;
wire S8831;
wire S8832;
wire S8833;
wire S8834;
wire S8835;
wire S8836;
wire S8837;
wire S8838;
wire S8839;
wire S8840;
wire S8841;
wire S8842;
wire S8843;
wire S8844;
wire S8845;
wire S8846;
wire S8847;
wire S8848;
wire S8849;
wire S8850;
wire S8851;
wire S8852;
wire S8853;
wire S8854;
wire S8855;
wire S8856;
wire S8857;
wire S8858;
wire S8859;
wire S8860;
wire S8861;
wire S8862;
wire S8863;
wire S8864;
wire S8865;
wire S8866;
wire S8867;
wire S8868;
wire S8869;
wire S8870;
wire S8871;
wire S8872;
wire S8873;
wire S8874;
wire S8875;
wire S8876;
wire S8877;
wire S8878;
wire S8879;
wire S8880;
wire S8881;
wire S8882;
wire S8883;
wire S8884;
wire S8885;
wire S8886;
wire S8887;
wire S8888;
wire S8889;
wire S8890;
wire S8891;
wire S8892;
wire S8893;
wire S8894;
wire S8895;
wire S8896;
wire S8897;
wire S8898;
wire S8899;
wire S8900;
wire S8901;
wire S8902;
wire S8903;
wire S8904;
wire S8905;
wire S8906;
wire S8907;
wire S8908;
wire S8909;
wire S8910;
wire S8911;
wire S8912;
wire S8913;
wire S8914;
wire S8915;
wire S8916;
wire S8917;
wire S8918;
wire S8919;
wire S8920;
wire S8921;
wire S8922;
wire S8923;
wire S8924;
wire S8925;
wire S8926;
wire S8927;
wire S8928;
wire S8929;
wire S8930;
wire S8931;
wire S8932;
wire S8933;
wire S8934;
wire S8935;
wire S8936;
wire S8937;
wire S8938;
wire S8939;
wire S8940;
wire S8941;
wire S8942;
wire S8943;
wire S8944;
wire S8945;
wire S8946;
wire S8947;
wire S8948;
wire S8949;
wire S8950;
wire S8951;
wire S8952;
wire S8953;
wire S8954;
wire S8955;
wire S8956;
wire S8957;
wire S8958;
wire S8959;
wire S8960;
wire S8961;
wire S8962;
wire S8963;
wire S8964;
wire S8965;
wire S8966;
wire S8967;
wire S8968;
wire S8969;
wire S8970;
wire S8971;
wire S8972;
wire S8973;
wire S8974;
wire S8975;
wire S8976;
wire S8977;
wire S8978;
wire S8979;
wire S8980;
wire S8981;
wire S8982;
wire S8983;
wire S8984;
wire S8985;
wire S8986;
wire S8987;
wire S8988;
wire S8989;
wire S8990;
wire S8991;
wire S8992;
wire S8993;
wire S8994;
wire S8995;
wire S8996;
wire S8997;
wire S8998;
wire S8999;
wire S9000;
wire S9001;
wire S9002;
wire S9003;
wire S9004;
wire S9005;
wire S9006;
wire S9007;
wire S9008;
wire S9009;
wire S9010;
wire S9011;
wire S9012;
wire S9013;
wire S9014;
wire S9015;
wire S9016;
wire S9017;
wire S9018;
wire S9019;
wire S9020;
wire S9021;
wire S9022;
wire S9023;
wire S9024;
wire S9025;
wire S9026;
wire S9027;
wire S9028;
wire S9029;
wire S9030;
wire S9031;
wire S9032;
wire S9033;
wire S9034;
wire S9035;
wire S9036;
wire S9037;
wire S9038;
wire S9039;
wire S9040;
wire S9041;
wire S9042;
wire S9043;
wire S9044;
wire S9045;
wire S9046;
wire S9047;
wire S9048;
wire S9049;
wire S9050;
wire S9051;
wire S9052;
wire S9053;
wire S9054;
wire S9055;
wire S9056;
wire S9057;
wire S9058;
wire S9059;
wire S9060;
wire S9061;
wire S9062;
wire S9063;
wire S9064;
wire S9065;
wire S9066;
wire S9067;
wire S9068;
wire S9069;
wire S9070;
wire S9071;
wire S9072;
wire S9073;
wire S9074;
wire S9075;
wire S9076;
wire S9077;
wire S9078;
wire S9079;
wire S9080;
wire S9081;
wire S9082;
wire S9083;
wire S9084;
wire S9085;
wire S9086;
wire S9087;
wire S9088;
wire S9089;
wire S9090;
wire S9091;
wire S9092;
wire S9093;
wire S9094;
wire S9095;
wire S9096;
wire S9097;
wire S9098;
wire S9099;
wire S9100;
wire S9101;
wire S9102;
wire S9103;
wire S9104;
wire S9105;
wire S9106;
wire S9107;
wire S9108;
wire S9109;
wire S9110;
wire S9111;
wire S9112;
wire S9113;
wire S9114;
wire S9115;
wire S9116;
wire S9117;
wire S9118;
wire S9119;
wire S9120;
wire S9121;
wire S9122;
wire S9123;
wire S9124;
wire S9125;
wire S9126;
wire S9127;
wire S9128;
wire S9129;
wire S9130;
wire S9131;
wire S9132;
wire S9133;
wire S9134;
wire S9135;
wire S9136;
wire S9137;
wire S9138;
wire S9139;
wire S9140;
wire S9141;
wire S9142;
wire S9143;
wire S9144;
wire S9145;
wire S9146;
wire S9147;
wire S9148;
wire S9149;
wire S9150;
wire S9151;
wire S9152;
wire S9153;
wire S9154;
wire S9155;
wire S9156;
wire S9157;
wire S9158;
wire S9159;
wire S9160;
wire S9161;
wire S9162;
wire S9163;
wire S9164;
wire S9165;
wire S9166;
wire S9167;
wire S9168;
wire S9169;
wire S9170;
wire S9171;
wire S9172;
wire S9173;
wire S9174;
wire S9175;
wire S9176;
wire S9177;
wire S9178;
wire S9179;
wire S9180;
wire S9181;
wire S9182;
wire S9183;
wire S9184;
wire S9185;
wire S9186;
wire S9187;
wire S9188;
wire S9189;
wire S9190;
wire S9191;
wire S9192;
wire S9193;
wire S9194;
wire S9195;
wire S9196;
wire S9197;
wire S9198;
wire S9199;
wire S9200;
wire S9201;
wire S9202;
wire S9203;
wire S9204;
wire S9205;
wire S9206;
wire S9207;
wire S9208;
wire S9209;
wire S9210;
wire S9211;
wire S9212;
wire S9213;
wire S9214;
wire S9215;
wire S9216;
wire S9217;
wire S9218;
wire S9219;
wire S9220;
wire S9221;
wire S9222;
wire S9223;
wire S9224;
wire S9225;
wire S9226;
wire S9227;
wire S9228;
wire S9229;
wire S9230;
wire S9231;
wire S9232;
wire S9233;
wire S9234;
wire S9235;
wire S9236;
wire S9237;
wire S9238;
wire S9239;
wire S9240;
wire S9241;
wire S9242;
wire S9243;
wire S9244;
wire S9245;
wire S9246;
wire S9247;
wire S9248;
wire S9249;
wire S9250;
wire S9251;
wire S9252;
wire S9253;
wire S9254;
wire S9255;
wire S9256;
wire S9257;
wire S9258;
wire S9259;
wire S9260;
wire S9261;
wire S9262;
wire S9263;
wire S9264;
wire S9265;
wire S9266;
wire S9267;
wire S9268;
wire S9269;
wire S9270;
wire S9271;
wire S9272;
wire S9273;
wire S9274;
wire S9275;
wire S9276;
wire S9277;
wire S9278;
wire S9279;
wire S9280;
wire S9281;
wire S9282;
wire S9283;
wire S9284;
wire S9285;
wire S9286;
wire S9287;
wire S9288;
wire S9289;
wire S9290;
wire S9291;
wire S9292;
wire S9293;
wire S9294;
wire S9295;
wire S9296;
wire S9297;
wire S9298;
wire S9299;
wire S9300;
wire S9301;
wire S9302;
wire S9303;
wire S9304;
wire S9305;
wire S9306;
wire S9307;
wire S9308;
wire S9309;
wire S9310;
wire S9311;
wire S9312;
wire S9313;
wire S9314;
wire S9315;
wire S9316;
wire S9317;
wire S9318;
wire S9319;
wire S9320;
wire S9321;
wire S9322;
wire S9323;
wire S9324;
wire S9325;
wire S9326;
wire S9327;
wire S9328;
wire S9329;
wire S9330;
wire S9331;
wire S9332;
wire S9333;
wire S9334;
wire S9335;
wire S9336;
wire S9337;
wire S9338;
wire S9339;
wire S9340;
wire S9341;
wire S9342;
wire S9343;
wire S9344;
wire S9345;
wire S9346;
wire S9347;
wire S9348;
wire S9349;
wire S9350;
wire S9351;
wire S9352;
wire S9353;
wire S9354;
wire S9355;
wire S9356;
wire S9357;
wire S9358;
wire S9359;
wire S9360;
wire S9361;
wire S9362;
wire S9363;
wire S9364;
wire S9365;
wire S9366;
wire S9367;
wire S9368;
wire S9369;
wire S9370;
wire S9371;
wire S9372;
wire S9373;
wire S9374;
wire S9375;
wire S9376;
wire S9377;
wire S9378;
wire S9379;
wire S9380;
wire S9381;
wire S9382;
wire S9383;
wire S9384;
wire S9385;
wire S9386;
wire S9387;
wire S9388;
wire S9389;
wire S9390;
wire S9391;
wire S9392;
wire S9393;
wire S9394;
wire S9395;
wire S9396;
wire S9397;
wire S9398;
wire S9399;
wire S9400;
wire S9401;
wire S9402;
wire S9403;
wire S9404;
wire S9405;
wire S9406;
wire S9407;
wire S9408;
wire S9409;
wire S9410;
wire S9411;
wire S9412;
wire S9413;
wire S9414;
wire S9415;
wire S9416;
wire S9417;
wire S9418;
wire S9419;
wire S9420;
wire S9421;
wire S9422;
wire S9423;
wire S9424;
wire S9425;
wire S9426;
wire S9427;
wire S9428;
wire S9429;
wire S9430;
wire S9431;
wire S9432;
wire S9433;
wire S9434;
wire S9435;
wire S9436;
wire S9437;
wire S9438;
wire S9439;
wire S9440;
wire S9441;
wire S9442;
wire S9443;
wire S9444;
wire S9445;
wire S9446;
wire S9447;
wire S9448;
wire S9449;
wire S9450;
wire S9451;
wire S9452;
wire S9453;
wire S9454;
wire S9455;
wire S9456;
wire S9457;
wire S9458;
wire S9459;
wire S9460;
wire S9461;
wire S9462;
wire S9463;
wire S9464;
wire S9465;
wire S9466;
wire S9467;
wire S9468;
wire S9469;
wire S9470;
wire S9471;
wire S9472;
wire S9473;
wire S9474;
wire S9475;
wire S9476;
wire S9477;
wire S9478;
wire S9479;
wire S9480;
wire S9481;
wire S9482;
wire S9483;
wire S9484;
wire S9485;
wire S9486;
wire S9487;
wire S9488;
wire S9489;
wire S9490;
wire S9491;
wire S9492;
wire S9493;
wire S9494;
wire S9495;
wire S9496;
wire S9497;
wire S9498;
wire S9499;
wire S9500;
wire S9501;
wire S9502;
wire S9503;
wire S9504;
wire S9505;
wire S9506;
wire S9507;
wire S9508;
wire S9509;
wire S9510;
wire S9511;
wire S9512;
wire S9513;
wire S9514;
wire S9515;
wire S9516;
wire S9517;
wire S9518;
wire S9519;
wire S9520;
wire S9521;
wire S9522;
wire S9523;
wire S9524;
wire S9525;
wire S9526;
wire S9527;
wire S9528;
wire S9529;
wire S9530;
wire S9531;
wire S9532;
wire S9533;
wire S9534;
wire S9535;
wire S9536;
wire S9537;
wire S9538;
wire S9539;
wire S9540;
wire S9541;
wire S9542;
wire S9543;
wire S9544;
wire S9545;
wire S9546;
wire S9547;
wire S9548;
wire S9549;
wire S9550;
wire S9551;
wire S9552;
wire S9553;
wire S9554;
wire S9555;
wire S9556;
wire S9557;
wire S9558;
wire S9559;
wire S9560;
wire S9561;
wire S9562;
wire S9563;
wire S9564;
wire S9565;
wire S9566;
wire S9567;
wire S9568;
wire S9569;
wire S9570;
wire S9571;
wire S9572;
wire S9573;
wire S9574;
wire S9575;
wire S9576;
wire S9577;
wire S9578;
wire S9579;
wire S9580;
wire S9581;
wire S9582;
wire S9583;
wire S9584;
wire S9585;
wire S9586;
wire S9587;
wire S9588;
wire S9589;
wire S9590;
wire S9591;
wire S9592;
wire S9593;
wire S9594;
wire S9595;
wire S9596;
wire S9597;
wire S9598;
wire S9599;
wire S9600;
wire S9601;
wire S9602;
wire S9603;
wire S9604;
wire S9605;
wire S9606;
wire S9607;
wire S9608;
wire S9609;
wire S9610;
wire S9611;
wire S9612;
wire S9613;
wire S9614;
wire S9615;
wire S9616;
wire S9617;
wire S9618;
wire S9619;
wire S9620;
wire S9621;
wire S9622;
wire S9623;
wire S9624;
wire S9625;
wire S9626;
wire S9627;
wire S9628;
wire S9629;
wire S9630;
wire S9631;
wire S9632;
wire S9633;
wire S9634;
wire S9635;
wire S9636;
wire S9637;
wire S9638;
wire S9639;
wire S9640;
wire S9641;
wire S9642;
wire S9643;
wire S9644;
wire S9645;
wire S9646;
wire S9647;
wire S9648;
wire S9649;
wire S9650;
wire S9651;
wire S9652;
wire S9653;
wire S9654;
wire S9655;
wire S9656;
wire S9657;
wire S9658;
wire S9659;
wire S9660;
wire S9661;
wire S9662;
wire S9663;
wire S9664;
wire S9665;
wire S9666;
wire S9667;
wire S9668;
wire S9669;
wire S9670;
wire S9671;
wire S9672;
wire S9673;
wire S9674;
wire S9675;
wire S9676;
wire S9677;
wire S9678;
wire S9679;
wire S9680;
wire S9681;
wire S9682;
wire S9683;
wire S9684;
wire S9685;
wire S9686;
wire S9687;
wire S9688;
wire S9689;
wire S9690;
wire S9691;
wire S9692;
wire S9693;
wire S9694;
wire S9695;
wire S9696;
wire S9697;
wire S9698;
wire S9699;
wire S9700;
wire S9701;
wire S9702;
wire S9703;
wire S9704;
wire S9705;
wire S9706;
wire S9707;
wire S9708;
wire S9709;
wire S9710;
wire S9711;
wire S9712;
wire S9713;
wire S9714;
wire S9715;
wire S9716;
wire S9717;
wire S9718;
wire S9719;
wire S9720;
wire S9721;
wire S9722;
wire S9723;
wire S9724;
wire S9725;
wire S9726;
wire S9727;
wire S9728;
wire S9729;
wire S9730;
wire S9731;
wire S9732;
wire S9733;
wire S9734;
wire S9735;
wire S9736;
wire S9737;
wire S9738;
wire S9739;
wire S9740;
wire S9741;
wire S9742;
wire S9743;
wire S9744;
wire S9745;
wire S9746;
wire S9747;
wire S9748;
wire S9749;
wire S9750;
wire S9751;
wire S9752;
wire S9753;
wire S9754;
wire S9755;
wire S9756;
wire S9757;
wire S9758;
wire S9759;
wire S9760;
wire S9761;
wire S9762;
wire S9763;
wire S9764;
wire S9765;
wire S9766;
wire S9767;
wire S9768;
wire S9769;
wire S9770;
wire S9771;
wire S9772;
wire S9773;
wire S9774;
wire S9775;
wire S9776;
wire S9777;
wire S9778;
wire S9779;
wire S9780;
wire S9781;
wire S9782;
wire S9783;
wire S9784;
wire S9785;
wire S9786;
wire S9787;
wire S9788;
wire S9789;
wire S9790;
wire S9791;
wire S9792;
wire S9793;
wire S9794;
wire S9795;
wire S9796;
wire S9797;
wire S9798;
wire S9799;
wire S9800;
wire S9801;
wire S9802;
wire S9803;
wire S9804;
wire S9805;
wire S9806;
wire S9807;
wire S9808;
wire S9809;
wire S9810;
wire S9811;
wire S9812;
wire S9813;
wire S9814;
wire S9815;
wire S9816;
wire S9817;
wire S9818;
wire S9819;
wire S9820;
wire S9821;
wire S9822;
wire S9823;
wire S9824;
wire S9825;
wire S9826;
wire S9827;
wire S9828;
wire S9829;
wire S9830;
wire S9831;
wire S9832;
wire S9833;
wire S9834;
wire S9835;
wire S9836;
wire S9837;
wire S9838;
wire S9839;
wire S9840;
wire S9841;
wire S9842;
wire S9843;
wire S9844;
wire S9845;
wire S9846;
wire S9847;
wire S9848;
wire S9849;
wire S9850;
wire S9851;
wire S9852;
wire S9853;
wire S9854;
wire S9855;
wire S9856;
wire S9857;
wire S9858;
wire S9859;
wire S9860;
wire S9861;
wire S9862;
wire S9863;
wire S9864;
wire S9865;
wire S9866;
wire S9867;
wire S9868;
wire S9869;
wire S9870;
wire S9871;
wire S9872;
wire S9873;
wire S9874;
wire S9875;
wire S9876;
wire S9877;
wire S9878;
wire S9879;
wire S9880;
wire S9881;
wire S9882;
wire S9883;
wire S9884;
wire S9885;
wire S9886;
wire S9887;
wire S9888;
wire S9889;
wire S9890;
wire S9891;
wire S9892;
wire S9893;
wire S9894;
wire S9895;
wire S9896;
wire S9897;
wire S9898;
wire S9899;
wire S9900;
wire S9901;
wire S9902;
wire S9903;
wire S9904;
wire S9905;
wire S9906;
wire S9907;
wire S9908;
wire S9909;
wire S9910;
wire S9911;
wire S9912;
wire S9913;
wire S9914;
wire S9915;
wire S9916;
wire S9917;
wire S9918;
wire S9919;
wire S9920;
wire S9921;
wire S9922;
wire S9923;
wire S9924;
wire S9925;
wire S9926;
wire S9927;
wire S9928;
wire S9929;
wire S9930;
wire S9931;
wire S9932;
wire S9933;
wire S9934;
wire S9935;
wire S9936;
wire S9937;
wire S9938;
wire S9939;
wire S9940;
wire S9941;
wire S9942;
wire S9943;
wire S9944;
wire S9945;
wire S9946;
wire S9947;
wire S9948;
wire S9949;
wire S9950;
wire S9951;
wire S9952;
wire S9953;
wire S9954;
wire S9955;
wire S9956;
wire S9957;
wire S9958;
wire S9959;
wire S9960;
wire S9961;
wire S9962;
wire S9963;
wire S9964;
wire S9965;
wire S9966;
wire S9967;
wire S9968;
wire S9969;
wire S9970;
wire S9971;
wire S9972;
wire S9973;
wire S9974;
wire S9975;
wire S9976;
wire S9977;
wire S9978;
wire S9979;
wire S9980;
wire S9981;
wire S9982;
wire S9983;
wire S9984;
wire S9985;
wire S9986;
wire S9987;
wire S9988;
wire S9989;
wire S9990;
wire S9991;
wire S9992;
wire S9993;
wire S9994;
wire S9995;
wire S9996;
wire S9997;
wire S9998;
wire S9999;
wire S10000;
wire S10001;
wire S10002;
wire S10003;
wire S10004;
wire S10005;
wire S10006;
wire S10007;
wire S10008;
wire S10009;
wire S10010;
wire S10011;
wire S10012;
wire S10013;
wire S10014;
wire S10015;
wire S10016;
wire S10017;
wire S10018;
wire S10019;
wire S10020;
wire S10021;
wire S10022;
wire S10023;
wire S10024;
wire S10025;
wire S10026;
wire S10027;
wire S10028;
wire S10029;
wire S10030;
wire S10031;
wire S10032;
wire S10033;
wire S10034;
wire S10035;
wire S10036;
wire S10037;
wire S10038;
wire S10039;
wire S10040;
wire S10041;
wire S10042;
wire S10043;
wire S10044;
wire S10045;
wire S10046;
wire S10047;
wire S10048;
wire S10049;
wire S10050;
wire S10051;
wire S10052;
wire S10053;
wire S10054;
wire S10055;
wire S10056;
wire S10057;
wire S10058;
wire S10059;
wire S10060;
wire S10061;
wire S10062;
wire S10063;
wire S10064;
wire S10065;
wire S10066;
wire S10067;
wire S10068;
wire S10069;
wire S10070;
wire S10071;
wire S10072;
wire S10073;
wire S10074;
wire S10075;
wire S10076;
wire S10077;
wire S10078;
wire S10079;
wire S10080;
wire S10081;
wire S10082;
wire S10083;
wire S10084;
wire S10085;
wire S10086;
wire S10087;
wire S10088;
wire S10089;
wire S10090;
wire S10091;
wire S10092;
wire S10093;
wire S10094;
wire S10095;
wire S10096;
wire S10097;
wire S10098;
wire S10099;
wire S10100;
wire S10101;
wire S10102;
wire S10103;
wire S10104;
wire S10105;
wire S10106;
wire S10107;
wire S10108;
wire S10109;
wire S10110;
wire S10111;
wire S10112;
wire S10113;
wire S10114;
wire S10115;
wire S10116;
wire S10117;
wire S10118;
wire S10119;
wire S10120;
wire S10121;
wire S10122;
wire S10123;
wire S10124;
wire S10125;
wire S10126;
wire S10127;
wire S10128;
wire S10129;
wire S10130;
wire S10131;
wire S10132;
wire S10133;
wire S10134;
wire S10135;
wire S10136;
wire S10137;
wire S10138;
wire S10139;
wire S10140;
wire S10141;
wire S10142;
wire S10143;
wire S10144;
wire S10145;
wire S10146;
wire S10147;
wire S10148;
wire S10149;
wire S10150;
wire S10151;
wire S10152;
wire S10153;
wire S10154;
wire S10155;
wire S10156;
wire S10157;
wire S10158;
wire S10159;
wire S10160;
wire S10161;
wire S10162;
wire S10163;
wire S10164;
wire S10165;
wire S10166;
wire S10167;
wire S10168;
wire S10169;
wire S10170;
wire S10171;
wire S10172;
wire S10173;
wire S10174;
wire S10175;
wire S10176;
wire S10177;
wire S10178;
wire S10179;
wire S10180;
wire S10181;
wire S10182;
wire S10183;
wire S10184;
wire S10185;
wire S10186;
wire S10187;
wire S10188;
wire S10189;
wire S10190;
wire S10191;
wire S10192;
wire S10193;
wire S10194;
wire S10195;
wire S10196;
wire S10197;
wire S10198;
wire S10199;
wire S10200;
wire S10201;
wire S10202;
wire S10203;
wire S10204;
wire S10205;
wire S10206;
wire S10207;
wire S10208;
wire S10209;
wire S10210;
wire S10211;
wire S10212;
wire S10213;
wire S10214;
wire S10215;
wire S10216;
wire S10217;
wire S10218;
wire S10219;
wire S10220;
wire S10221;
wire S10222;
wire S10223;
wire S10224;
wire S10225;
wire S10226;
wire S10227;
wire S10228;
wire S10229;
wire S10230;
wire S10231;
wire S10232;
wire S10233;
wire S10234;
wire S10235;
wire S10236;
wire S10237;
wire S10238;
wire S10239;
wire S10240;
wire S10241;
wire S10242;
wire S10243;
wire S10244;
wire S10245;
wire S10246;
wire S10247;
wire S10248;
wire S10249;
wire S10250;
wire S10251;
wire S10252;
wire S10253;
wire S10254;
wire S10255;
wire S10256;
wire S10257;
wire S10258;
wire S10259;
wire S10260;
wire S10261;
wire S10262;
wire S10263;
wire S10264;
wire S10265;
wire S10266;
wire S10267;
wire S10268;
wire S10269;
wire S10270;
wire S10271;
wire S10272;
wire S10273;
wire S10274;
wire S10275;
wire S10276;
wire S10277;
wire S10278;
wire S10279;
wire S10280;
wire S10281;
wire S10282;
wire S10283;
wire S10284;
wire S10285;
wire S10286;
wire S10287;
wire S10288;
wire S10289;
wire S10290;
wire S10291;
wire S10292;
wire S10293;
wire S10294;
wire S10295;
wire S10296;
wire S10297;
wire S10298;
wire S10299;
wire S10300;
wire S10301;
wire S10302;
wire S10303;
wire S10304;
wire S10305;
wire S10306;
wire S10307;
wire S10308;
wire S10309;
wire S10310;
wire S10311;
wire S10312;
wire S10313;
wire S10314;
wire S10315;
wire S10316;
wire S10317;
wire S10318;
wire S10319;
wire S10320;
wire S10321;
wire S10322;
wire S10323;
wire S10324;
wire S10325;
wire S10326;
wire S10327;
wire S10328;
wire S10329;
wire S10330;
wire S10331;
wire S10332;
wire S10333;
wire S10334;
wire S10335;
wire S10336;
wire S10337;
wire S10338;
wire S10339;
wire S10340;
wire S10341;
wire S10342;
wire S10343;
wire S10344;
wire S10345;
wire S10346;
wire S10347;
wire S10348;
wire S10349;
wire S10350;
wire S10351;
wire S10352;
wire S10353;
wire S10354;
wire S10355;
wire S10356;
wire S10357;
wire S10358;
wire S10359;
wire S10360;
wire S10361;
wire S10362;
wire S10363;
wire S10364;
wire S10365;
wire S10366;
wire S10367;
wire S10368;
wire S10369;
wire S10370;
wire S10371;
wire S10372;
wire S10373;
wire S10374;
wire S10375;
wire S10376;
wire S10377;
wire S10378;
wire S10379;
wire S10380;
wire S10381;
wire S10382;
wire S10383;
wire S10384;
wire S10385;
wire S10386;
wire S10387;
wire S10388;
wire S10389;
wire S10390;
wire S10391;
wire S10392;
wire S10393;
wire S10394;
wire S10395;
wire S10396;
wire S10397;
wire S10398;
wire S10399;
wire S10400;
wire S10401;
wire S10402;
wire S10403;
wire S10404;
wire S10405;
wire S10406;
wire S10407;
wire S10408;
wire S10409;
wire S10410;
wire S10411;
wire S10412;
wire S10413;
wire S10414;
wire S10415;
wire S10416;
wire S10417;
wire S10418;
wire S10419;
wire S10420;
wire S10421;
wire S10422;
wire S10423;
wire S10424;
wire S10425;
wire S10426;
wire S10427;
wire S10428;
wire S10429;
wire S10430;
wire S10431;
wire S10432;
wire S10433;
wire S10434;
wire S10435;
wire S10436;
wire S10437;
wire S10438;
wire S10439;
wire S10440;
wire S10441;
wire S10442;
wire S10443;
wire S10444;
wire S10445;
wire S10446;
wire S10447;
wire S10448;
wire S10449;
wire S10450;
wire S10451;
wire S10452;
wire S10453;
wire S10454;
wire S10455;
wire S10456;
wire S10457;
wire S10458;
wire S10459;
wire S10460;
wire S10461;
wire S10462;
wire S10463;
wire S10464;
wire S10465;
wire S10466;
wire S10467;
wire S10468;
wire S10469;
wire S10470;
wire S10471;
wire S10472;
wire S10473;
wire S10474;
wire S10475;
wire S10476;
wire S10477;
wire S10478;
wire S10479;
wire S10480;
wire S10481;
wire S10482;
wire S10483;
wire S10484;
wire S10485;
wire S10486;
wire S10487;
wire S10488;
wire S10489;
wire S10490;
wire S10491;
wire S10492;
wire S10493;
wire S10494;
wire S10495;
wire S10496;
wire S10497;
wire S10498;
wire S10499;
wire S10500;
wire S10501;
wire S10502;
wire S10503;
wire S10504;
wire S10505;
wire S10506;
wire S10507;
wire S10508;
wire S10509;
wire S10510;
wire S10511;
wire S10512;
wire S10513;
wire S10514;
wire S10515;
wire S10516;
wire S10517;
wire S10518;
wire S10519;
wire S10520;
wire S10521;
wire S10522;
wire S10523;
wire S10524;
wire S10525;
wire S10526;
wire S10527;
wire S10528;
wire S10529;
wire S10530;
wire S10531;
wire S10532;
wire S10533;
wire S10534;
wire S10535;
wire S10536;
wire S10537;
wire S10538;
wire S10539;
wire S10540;
wire S10541;
wire S10542;
wire S10543;
wire S10544;
wire S10545;
wire S10546;
wire S10547;
wire S10548;
wire S10549;
wire S10550;
wire S10551;
wire S10552;
wire S10553;
wire S10554;
wire S10555;
wire S10556;
wire S10557;
wire S10558;
wire S10559;
wire S10560;
wire S10561;
wire S10562;
wire S10563;
wire S10564;
wire S10565;
wire S10566;
wire S10567;
wire S10568;
wire S10569;
wire S10570;
wire S10571;
wire S10572;
wire S10573;
wire S10574;
wire S10575;
wire S10576;
wire S10577;
wire S10578;
wire S10579;
wire S10580;
wire S10581;
wire S10582;
wire S10583;
wire S10584;
wire S10585;
wire S10586;
wire S10587;
wire S10588;
wire S10589;
wire S10590;
wire S10591;
wire S10592;
wire S10593;
wire S10594;
wire S10595;
wire S10596;
wire S10597;
wire S10598;
wire S10599;
wire S10600;
wire S10601;
wire S10602;
wire S10603;
wire S10604;
wire S10605;
wire S10606;
wire S10607;
wire S10608;
wire S10609;
wire S10610;
wire S10611;
wire S10612;
wire S10613;
wire S10614;
wire S10615;
wire S10616;
wire S10617;
wire S10618;
wire S10619;
wire S10620;
wire S10621;
wire S10622;
wire S10623;
wire S10624;
wire S10625;
wire S10626;
wire S10627;
wire S10628;
wire S10629;
wire S10630;
wire S10631;
wire S10632;
wire S10633;
wire S10634;
wire S10635;
wire S10636;
wire S10637;
wire S10638;
wire S10639;
wire S10640;
wire S10641;
wire S10642;
wire S10643;
wire S10644;
wire S10645;
wire S10646;
wire S10647;
wire S10648;
wire S10649;
wire S10650;
wire S10651;
wire S10652;
wire S10653;
wire S10654;
wire S10655;
wire S10656;
wire S10657;
wire S10658;
wire S10659;
wire S10660;
wire S10661;
wire S10662;
wire S10663;
wire S10664;
wire S10665;
wire S10666;
wire S10667;
wire S10668;
wire S10669;
wire S10670;
wire S10671;
wire S10672;
wire S10673;
wire S10674;
wire S10675;
wire S10676;
wire S10677;
wire S10678;
wire S10679;
wire S10680;
wire S10681;
wire S10682;
wire S10683;
wire S10684;
wire S10685;
wire S10686;
wire S10687;
wire S10688;
wire S10689;
wire S10690;
wire S10691;
wire S10692;
wire S10693;
wire S10694;
wire S10695;
wire S10696;
wire S10697;
wire S10698;
wire S10699;
wire S10700;
wire S10701;
wire S10702;
wire S10703;
wire S10704;
wire S10705;
wire S10706;
wire S10707;
wire S10708;
wire S10709;
wire S10710;
wire S10711;
wire S10712;
wire S10713;
wire S10714;
wire S10715;
wire S10716;
wire S10717;
wire S10718;
wire S10719;
wire S10720;
wire S10721;
wire S10722;
wire S10723;
wire S10724;
wire S10725;
wire S10726;
wire S10727;
wire S10728;
wire S10729;
wire S10730;
wire S10731;
wire S10732;
wire S10733;
wire S10734;
wire S10735;
wire S10736;
wire S10737;
wire S10738;
wire S10739;
wire S10740;
wire S10741;
wire S10742;
wire S10743;
wire S10744;
wire S10745;
wire S10746;
wire S10747;
wire S10748;
wire S10749;
wire S10750;
wire S10751;
wire S10752;
wire S10753;
wire S10754;
wire S10755;
wire S10756;
wire S10757;
wire S10758;
wire S10759;
wire S10760;
wire S10761;
wire S10762;
wire S10763;
wire S10764;
wire S10765;
wire S10766;
wire S10767;
wire S10768;
wire S10769;
wire S10770;
wire S10771;
wire S10772;
wire S10773;
wire S10774;
wire S10775;
wire S10776;
wire S10777;
wire S10778;
wire S10779;
wire S10780;
wire S10781;
wire S10782;
wire S10783;
wire S10784;
wire S10785;
wire S10786;
wire S10787;
wire S10788;
wire S10789;
wire S10790;
wire S10791;
wire S10792;
wire S10793;
wire S10794;
wire S10795;
wire S10796;
wire S10797;
wire S10798;
wire S10799;
wire S10800;
wire S10801;
wire S10802;
wire S10803;
wire S10804;
wire S10805;
wire S10806;
wire S10807;
wire S10808;
wire S10809;
wire S10810;
wire S10811;
wire S10812;
wire S10813;
wire S10814;
wire S10815;
wire S10816;
wire S10817;
wire S10818;
wire S10819;
wire S10820;
wire S10821;
wire S10822;
wire S10823;
wire S10824;
wire S10825;
wire S10826;
wire S10827;
wire S10828;
wire S10829;
wire S10830;
wire S10831;
wire S10832;
wire S10833;
wire S10834;
wire S10835;
wire S10836;
wire S10837;
wire S10838;
wire S10839;
wire S10840;
wire S10841;
wire S10842;
wire S10843;
wire S10844;
wire S10845;
wire S10846;
wire S10847;
wire S10848;
wire S10849;
wire S10850;
wire S10851;
wire S10852;
wire S10853;
wire S10854;
wire S10855;
wire S10856;
wire S10857;
wire S10858;
wire S10859;
wire S10860;
wire S10861;
wire S10862;
wire S10863;
wire S10864;
wire S10865;
wire S10866;
wire S10867;
wire S10868;
wire S10869;
wire S10870;
wire S10871;
wire S10872;
wire S10873;
wire S10874;
wire S10875;
wire S10876;
wire S10877;
wire S10878;
wire S10879;
wire S10880;
wire S10881;
wire S10882;
wire S10883;
wire S10884;
wire S10885;
wire S10886;
wire S10887;
wire S10888;
wire S10889;
wire S10890;
wire S10891;
wire S10892;
wire S10893;
wire S10894;
wire S10895;
wire S10896;
wire S10897;
wire S10898;
wire S10899;
wire S10900;
wire S10901;
wire S10902;
wire S10903;
wire S10904;
wire S10905;
wire S10906;
wire S10907;
wire S10908;
wire S10909;
wire S10910;
wire S10911;
wire S10912;
wire S10913;
wire S10914;
wire S10915;
wire S10916;
wire S10917;
wire S10918;
wire S10919;
wire S10920;
wire S10921;
wire S10922;
wire S10923;
wire S10924;
wire S10925;
wire S10926;
wire S10927;
wire S10928;
wire S10929;
wire S10930;
wire S10931;
wire S10932;
wire S10933;
wire S10934;
wire S10935;
wire S10936;
wire S10937;
wire S10938;
wire S10939;
wire S10940;
wire S10941;
wire S10942;
wire S10943;
wire S10944;
wire S10945;
wire S10946;
wire S10947;
wire S10948;
wire S10949;
wire S10950;
wire S10951;
wire S10952;
wire S10953;
wire S10954;
wire S10955;
wire S10956;
wire S10957;
wire S10958;
wire S10959;
wire S10960;
wire S10961;
wire S10962;
wire S10963;
wire S10964;
wire S10965;
wire S10966;
wire S10967;
wire S10968;
wire S10969;
wire S10970;
wire S10971;
wire S10972;
wire S10973;
wire S10974;
wire S10975;
wire S10976;
wire S10977;
wire S10978;
wire S10979;
wire S10980;
wire S10981;
wire S10982;
wire S10983;
wire S10984;
wire S10985;
wire S10986;
wire S10987;
wire S10988;
wire S10989;
wire S10990;
wire S10991;
wire S10992;
wire S10993;
wire S10994;
wire S10995;
wire S10996;
wire S10997;
wire S10998;
wire S10999;
wire S11000;
wire S11001;
wire S11002;
wire S11003;
wire S11004;
wire S11005;
wire S11006;
wire S11007;
wire S11008;
wire S11009;
wire S11010;
wire S11011;
wire S11012;
wire S11013;
wire S11014;
wire S11015;
wire S11016;
wire S11017;
wire S11018;
wire S11019;
wire S11020;
wire S11021;
wire S11022;
wire S11023;
wire S11024;
wire S11025;
wire S11026;
wire S11027;
wire S11028;
wire S11029;
wire S11030;
wire S11031;
wire S11032;
wire S11033;
wire S11034;
wire S11035;
wire S11036;
wire S11037;
wire S11038;
wire S11039;
wire S11040;
wire S11041;
wire S11042;
wire S11043;
wire S11044;
wire S11045;
wire S11046;
wire S11047;
wire S11048;
wire S11049;
wire S11050;
wire S11051;
wire S11052;
wire S11053;
wire S11054;
wire S11055;
wire S11056;
wire S11057;
wire S11058;
wire S11059;
wire S11060;
wire S11061;
wire S11062;
wire S11063;
wire S11064;
wire S11065;
wire S11066;
wire S11067;
wire S11068;
wire S11069;
wire S11070;
wire S11071;
wire S11072;
wire S11073;
wire S11074;
wire S11075;
wire S11076;
wire S11077;
wire S11078;
wire S11079;
wire S11080;
wire S11081;
wire S11082;
wire S11083;
wire S11084;
wire S11085;
wire S11086;
wire S11087;
wire S11088;
wire S11089;
wire S11090;
wire S11091;
wire S11092;
wire S11093;
wire S11094;
wire S11095;
wire S11096;
wire S11097;
wire S11098;
wire S11099;
wire S11100;
wire S11101;
wire S11102;
wire S11103;
wire S11104;
wire S11105;
wire S11106;
wire S11107;
wire S11108;
wire S11109;
wire S11110;
wire S11111;
wire S11112;
wire S11113;
wire S11114;
wire S11115;
wire S11116;
wire S11117;
wire S11118;
wire S11119;
wire S11120;
wire S11121;
wire S11122;
wire S11123;
wire S11124;
wire S11125;
wire S11126;
wire S11127;
wire S11128;
wire S11129;
wire S11130;
wire S11131;
wire S11132;
wire S11133;
wire S11134;
wire S11135;
wire S11136;
wire S11137;
wire S11138;
wire S11139;
wire S11140;
wire S11141;
wire S11142;
wire S11143;
wire S11144;
wire S11145;
wire S11146;
wire S11147;
wire S11148;
wire S11149;
wire S11150;
wire S11151;
wire S11152;
wire S11153;
wire S11154;
wire S11155;
wire S11156;
wire S11157;
wire S11158;
wire S11159;
wire S11160;
wire S11161;
wire S11162;
wire S11163;
wire S11164;
wire S11165;
wire S11166;
wire S11167;
wire S11168;
wire S11169;
wire S11170;
wire S11171;
wire S11172;
wire S11173;
wire S11174;
wire S11175;
wire S11176;
wire S11177;
wire S11178;
wire S11179;
wire S11180;
wire S11181;
wire S11182;
wire S11183;
wire S11184;
wire S11185;
wire S11186;
wire S11187;
wire S11188;
wire S11189;
wire S11190;
wire S11191;
wire S11192;
wire S11193;
wire S11194;
wire S11195;
wire S11196;
wire S11197;
wire S11198;
wire S11199;
wire S11200;
wire S11201;
wire S11202;
wire S11203;
wire S11204;
wire S11205;
wire S11206;
wire S11207;
wire S11208;
wire S11209;
wire S11210;
wire S11211;
wire S11212;
wire S11213;
wire S11214;
wire S11215;
wire S11216;
wire S11217;
wire S11218;
wire S11219;
wire S11220;
wire S11221;
wire S11222;
wire S11223;
wire S11224;
wire S11225;
wire S11226;
wire S11227;
wire S11228;
wire S11229;
wire S11230;
wire S11231;
wire S11232;
wire S11233;
wire S11234;
wire S11235;
wire S11236;
wire S11237;
wire S11238;
wire S11239;
wire S11240;
wire S11241;
wire S11242;
wire S11243;
wire S11244;
wire S11245;
wire S11246;
wire S11247;
wire S11248;
wire S11249;
wire S11250;
wire S11251;
wire S11252;
wire S11253;
wire S11254;
wire S11255;
wire S11256;
wire S11257;
wire S11258;
wire S11259;
wire S11260;
wire S11261;
wire S11262;
wire S11263;
wire S11264;
wire S11265;
wire S11266;
wire S11267;
wire S11268;
wire S11269;
wire S11270;
wire S11271;
wire S11272;
wire S11273;
wire S11274;
wire S11275;
wire S11276;
wire S11277;
wire S11278;
wire S11279;
wire S11280;
wire S11281;
wire S11282;
wire S11283;
wire S11284;
wire S11285;
wire S11286;
wire S11287;
wire S11288;
wire S11289;
wire S11290;
wire S11291;
wire S11292;
wire S11293;
wire S11294;
wire S11295;
wire S11296;
wire S11297;
wire S11298;
wire S11299;
wire S11300;
wire S11301;
wire S11302;
wire S11303;
wire S11304;
wire S11305;
wire S11306;
wire S11307;
wire S11308;
wire S11309;
wire S11310;
wire S11311;
wire S11312;
wire S11313;
wire S11314;
wire S11315;
wire S11316;
wire S11317;
wire S11318;
wire S11319;
wire S11320;
wire S11321;
wire S11322;
wire S11323;
wire S11324;
wire S11325;
wire S11326;
wire S11327;
wire S11328;
wire S11329;
wire S11330;
wire S11331;
wire S11332;
wire S11333;
wire S11334;
wire S11335;
wire S11336;
wire S11337;
wire S11338;
wire S11339;
wire S11340;
wire S11341;
wire S11342;
wire S11343;
wire S11344;
wire S11345;
wire S11346;
wire S11347;
wire S11348;
wire S11349;
wire S11350;
wire S11351;
wire S11352;
wire S11353;
wire S11354;
wire S11355;
wire S11356;
wire S11357;
wire S11358;
wire S11359;
wire S11360;
wire S11361;
wire S11362;
wire S11363;
wire S11364;
wire S11365;
wire S11366;
wire S11367;
wire S11368;
wire S11369;
wire S11370;
wire S11371;
wire S11372;
wire S11373;
wire S11374;
wire S11375;
wire S11376;
wire S11377;
wire S11378;
wire S11379;
wire S11380;
wire S11381;
wire S11382;
wire S11383;
wire S11384;
wire S11385;
wire S11386;
wire S11387;
wire S11388;
wire S11389;
wire S11390;
wire S11391;
wire S11392;
wire S11393;
wire S11394;
wire S11395;
wire S11396;
wire S11397;
wire S11398;
wire S11399;
wire S11400;
wire S11401;
wire S11402;
wire S11403;
wire S11404;
wire S11405;
wire S11406;
wire S11407;
wire S11408;
wire S11409;
wire S11410;
wire S11411;
wire S11412;
wire S11413;
wire S11414;
wire S11415;
wire S11416;
wire S11417;
wire S11418;
wire S11419;
wire S11420;
wire S11421;
wire S11422;
wire S11423;
wire S11424;
wire S11425;
wire S11426;
wire S11427;
wire S11428;
wire S11429;
wire S11430;
wire S11431;
wire S11432;
wire S11433;
wire S11434;
wire S11435;
wire S11436;
wire S11437;
wire S11438;
wire S11439;
wire S11440;
wire S11441;
wire S11442;
wire S11443;
wire S11444;
wire S11445;
wire S11446;
wire S11447;
wire S11448;
wire S11449;
wire S11450;
wire S11451;
wire S11452;
wire S11453;
wire S11454;
wire S11455;
wire S11456;
wire S11457;
wire S11458;
wire S11459;
wire S11460;
wire S11461;
wire S11462;
wire S11463;
wire S11464;
wire S11465;
wire S11466;
wire S11467;
wire S11468;
wire S11469;
wire S11470;
wire S11471;
wire S11472;
wire S11473;
wire S11474;
wire S11475;
wire S11476;
wire S11477;
wire S11478;
wire S11479;
wire S11480;
wire S11481;
wire S11482;
wire S11483;
wire S11484;
wire S11485;
wire S11486;
wire S11487;
wire S11488;
wire S11489;
wire S11490;
wire S11491;
wire S11492;
wire S11493;
wire S11494;
wire S11495;
wire S11496;
wire S11497;
wire S11498;
wire S11499;
wire S11500;
wire S11501;
wire S11502;
wire S11503;
wire S11504;
wire S11505;
wire S11506;
wire S11507;
wire S11508;
wire S11509;
wire S11510;
wire S11511;
wire S11512;
wire S11513;
wire S11514;
wire S11515;
wire S11516;
wire S11517;
wire S11518;
wire S11519;
wire S11520;
wire S11521;
wire S11522;
wire S11523;
wire S11524;
wire S11525;
wire S11526;
wire S11527;
wire S11528;
wire S11529;
wire S11530;
wire S11531;
wire S11532;
wire S11533;
wire S11534;
wire S11535;
wire S11536;
wire S11537;
wire S11538;
wire S11539;
wire S11540;
wire S11541;
wire S11542;
wire S11543;
wire S11544;
wire S11545;
wire S11546;
wire S11547;
wire S11548;
wire S11549;
wire S11550;
wire S11551;
wire S11552;
wire S11553;
wire S11554;
wire S11555;
wire S11556;
wire S11557;
wire S11558;
wire S11559;
wire S11560;
wire S11561;
wire S11562;
wire S11563;
wire S11564;
wire S11565;
wire S11566;
wire S11567;
wire S11568;
wire S11569;
wire S11570;
wire S11571;
wire S11572;
wire S11573;
wire S11574;
wire S11575;
wire S11576;
wire S11577;
wire S11578;
wire S11579;
wire S11580;
wire S11581;
wire S11582;
wire S11583;
wire S11584;
wire S11585;
wire S11586;
wire S11587;
wire S11588;
wire S11589;
wire S11590;
wire S11591;
wire S11592;
wire S11593;
wire S11594;
wire S11595;
wire S11596;
wire S11597;
wire S11598;
wire S11599;
wire S11600;
wire S11601;
wire S11602;
wire S11603;
wire S11604;
wire S11605;
wire S11606;
wire S11607;
wire S11608;
wire S11609;
wire S11610;
wire S11611;
wire S11612;
wire S11613;
wire S11614;
wire S11615;
wire S11616;
wire S11617;
wire S11618;
wire S11619;
wire S11620;
wire S11621;
wire S11622;
wire S11623;
wire S11624;
wire S11625;
wire S11626;
wire S11627;
wire S11628;
wire S11629;
wire S11630;
wire S11631;
wire S11632;
wire S11633;
wire S11634;
wire S11635;
wire S11636;
wire S11637;
wire S11638;
wire S11639;
wire S11640;
wire S11641;
wire S11642;
wire S11643;
wire S11644;
wire S11645;
wire S11646;
wire S11647;
wire S11648;
wire S11649;
wire S11650;
wire S11651;
wire S11652;
wire S11653;
wire S11654;
wire S11655;
wire S11656;
wire S11657;
wire S11658;
wire S11659;
wire S11660;
wire S11661;
wire S11662;
wire S11663;
wire S11664;
wire S11665;
wire S11666;
wire S11667;
wire S11668;
wire S11669;
wire S11670;
wire S11671;
wire S11672;
wire S11673;
wire S11674;
wire S11675;
wire S11676;
wire S11677;
wire S11678;
wire S11679;
wire S11680;
wire S11681;
wire S11682;
wire S11683;
wire S11684;
wire S11685;
wire S11686;
wire S11687;
wire S11688;
wire S11689;
wire S11690;
wire S11691;
wire S11692;
wire S11693;
wire S11694;
wire S11695;
wire S11696;
wire S11697;
wire S11698;
wire S11699;
wire S11700;
wire S11701;
wire S11702;
wire S11703;
wire S11704;
wire S11705;
wire S11706;
wire S11707;
wire S11708;
wire S11709;
wire S11710;
wire S11711;
wire S11712;
wire S11713;
wire S11714;
wire S11715;
wire S11716;
wire S11717;
wire S11718;
wire S11719;
wire S11720;
wire S11721;
wire S11722;
wire S11723;
wire S11724;
wire S11725;
wire S11726;
wire S11727;
wire S11728;
wire S11729;
wire S11730;
wire S11731;
wire S11732;
wire S11733;
wire S11734;
wire S11735;
wire S11736;
wire S11737;
wire S11738;
wire S11739;
wire S11740;
wire S11741;
wire S11742;
wire S11743;
wire S11744;
wire S11745;
wire S11746;
wire S11747;
wire S11748;
wire S11749;
wire S11750;
wire S11751;
wire S11752;
wire S11753;
wire S11754;
wire S11755;
wire S11756;
wire S11757;
wire S11758;
wire S11759;
wire S11760;
wire S11761;
wire S11762;
wire S11763;
wire S11764;
wire S11765;
wire S11766;
wire S11767;
wire S11768;
wire S11769;
wire S11770;
wire S11771;
wire S11772;
wire S11773;
wire S11774;
wire S11775;
wire S11776;
wire S11777;
wire S11778;
wire S11779;
wire S11780;
wire S11781;
wire S11782;
wire S11783;
wire S11784;
wire S11785;
wire S11786;
wire S11787;
wire S11788;
wire S11789;
wire S11790;
wire S11791;
wire S11792;
wire S11793;
wire S11794;
wire S11795;
wire S11796;
wire S11797;
wire S11798;
wire S11799;
wire S11800;
wire S11801;
wire S11802;
wire S11803;
wire S11804;
wire S11805;
wire S11806;
wire S11807;
wire S11808;
wire S11809;
wire S11810;
wire S11811;
wire S11812;
wire S11813;
wire S11814;
wire S11815;
wire S11816;
wire S11817;
wire S11818;
wire S11819;
wire S11820;
wire S11821;
wire S11822;
wire S11823;
wire S11824;
wire S11825;
wire S11826;
wire S11827;
wire S11828;
wire S11829;
wire S11830;
wire S11831;
wire S11832;
wire S11833;
wire S11834;
wire S11835;
wire S11836;
wire S11837;
wire S11838;
wire S11839;
wire S11840;
wire S11841;
wire S11842;
wire S11843;
wire S11844;
wire S11845;
wire S11846;
wire S11847;
wire S11848;
wire S11849;
wire S11850;
wire S11851;
wire S11852;
wire S11853;
wire S11854;
wire S11855;
wire S11856;
wire S11857;
wire S11858;
wire S11859;
wire S11860;
wire S11861;
wire S11862;
wire S11863;
wire S11864;
wire S11865;
wire S11866;
wire S11867;
wire S11868;
wire S11869;
wire S11870;
wire S11871;
wire S11872;
wire S11873;
wire S11874;
wire S11875;
wire S11876;
wire S11877;
wire S11878;
wire S11879;
wire S11880;
wire S11881;
wire S11882;
wire S11883;
wire S11884;
wire S11885;
wire S11886;
wire S11887;
wire S11888;
wire S11889;
wire S11890;
wire S11891;
wire S11892;
wire S11893;
wire S11894;
wire S11895;
wire S11896;
wire S11897;
wire S11898;
wire S11899;
wire S11900;
wire S11901;
wire S11902;
wire S11903;
wire S11904;
wire S11905;
wire S11906;
wire S11907;
wire S11908;
wire S11909;
wire S11910;
wire S11911;
wire S11912;
wire S11913;
wire S11914;
wire S11915;
wire S11916;
wire S11917;
wire S11918;
wire S11919;
wire S11920;
wire S11921;
wire S11922;
wire S11923;
wire S11924;
wire S11925;
wire S11926;
wire S11927;
wire S11928;
wire S11929;
wire S11930;
wire S11931;
wire S11932;
wire S11933;
wire S11934;
wire S11935;
wire S11936;
wire S11937;
wire S11938;
wire S11939;
wire S11940;
wire S11941;
wire S11942;
wire S11943;
wire S11944;
wire S11945;
wire S11946;
wire S11947;
wire S11948;
wire S11949;
wire S11950;
wire S11951;
wire S11952;
wire S11953;
wire S11954;
wire S11955;
wire S11956;
wire S11957;
wire S11958;
wire S11959;
wire S11960;
wire S11961;
wire S11962;
wire S11963;
wire S11964;
wire S11965;
wire S11966;
wire S11967;
wire S11968;
wire S11969;
wire S11970;
wire S11971;
wire S11972;
wire S11973;
wire S11974;
wire S11975;
wire S11976;
wire S11977;
wire S11978;
wire S11979;
wire S11980;
wire S11981;
wire S11982;
wire S11983;
wire S11984;
wire S11985;
wire S11986;
wire S11987;
wire S11988;
wire S11989;
wire S11990;
wire S11991;
wire S11992;
wire S11993;
wire S11994;
wire S11995;
wire S11996;
wire S11997;
wire S11998;
wire S11999;
wire S12000;
wire S12001;
wire S12002;
wire S12003;
wire S12004;
wire S12005;
wire S12006;
wire S12007;
wire S12008;
wire S12009;
wire S12010;
wire S12011;
wire S12012;
wire S12013;
wire S12014;
wire S12015;
wire S12016;
wire S12017;
wire S12018;
wire S12019;
wire S12020;
wire S12021;
wire S12022;
wire S12023;
wire S12024;
wire S12025;
wire S12026;
wire S12027;
wire S12028;
wire S12029;
wire S12030;
wire S12031;
wire S12032;
wire S12033;
wire S12034;
wire S12035;
wire S12036;
wire S12037;
wire S12038;
wire S12039;
wire S12040;
wire S12041;
wire S12042;
wire S12043;
wire S12044;
wire S12045;
wire S12046;
wire S12047;
wire S12048;
wire S12049;
wire S12050;
wire S12051;
wire S12052;
wire S12053;
wire S12054;
wire S12055;
wire S12056;
wire S12057;
wire S12058;
wire S12059;
wire S12060;
wire S12061;
wire S12062;
wire S12063;
wire S12064;
wire S12065;
wire S12066;
wire S12067;
wire S12068;
wire S12069;
wire S12070;
wire S12071;
wire S12072;
wire S12073;
wire S12074;
wire S12075;
wire S12076;
wire S12077;
wire S12078;
wire S12079;
wire S12080;
wire S12081;
wire S12082;
wire S12083;
wire S12084;
wire S12085;
wire S12086;
wire S12087;
wire S12088;
wire S12089;
wire S12090;
wire S12091;
wire S12092;
wire S12093;
wire S12094;
wire S12095;
wire S12096;
wire S12097;
wire S12098;
wire S12099;
wire S12100;
wire S12101;
wire S12102;
wire S12103;
wire S12104;
wire S12105;
wire S12106;
wire S12107;
wire S12108;
wire S12109;
wire S12110;
wire S12111;
wire S12112;
wire S12113;
wire S12114;
wire S12115;
wire S12116;
wire S12117;
wire S12118;
wire S12119;
wire S12120;
wire S12121;
wire S12122;
wire S12123;
wire S12124;
wire S12125;
wire S12126;
wire S12127;
wire S12128;
wire S12129;
wire S12130;
wire S12131;
wire S12132;
wire S12133;
wire S12134;
wire S12135;
wire S12136;
wire S12137;
wire S12138;
wire S12139;
wire S12140;
wire S12141;
wire S12142;
wire S12143;
wire S12144;
wire S12145;
wire S12146;
wire S12147;
wire S12148;
wire S12149;
wire S12150;
wire S12151;
wire S12152;
wire S12153;
wire S12154;
wire S12155;
wire S12156;
wire S12157;
wire S12158;
wire S12159;
wire S12160;
wire S12161;
wire S12162;
wire S12163;
wire S12164;
wire S12165;
wire S12166;
wire S12167;
wire S12168;
wire S12169;
wire S12170;
wire S12171;
wire S12172;
wire S12173;
wire S12174;
wire S12175;
wire S12176;
wire S12177;
wire S12178;
wire S12179;
wire S12180;
wire S12181;
wire S12182;
wire S12183;
wire S12184;
wire S12185;
wire S12186;
wire S12187;
wire S12188;
wire S12189;
wire S12190;
wire S12191;
wire S12192;
wire S12193;
wire S12194;
wire S12195;
wire S12196;
wire S12197;
wire S12198;
wire S12199;
wire S12200;
wire S12201;
wire S12202;
wire S12203;
wire S12204;
wire S12205;
wire S12206;
wire S12207;
wire S12208;
wire S12209;
wire S12210;
wire S12211;
wire S12212;
wire S12213;
wire S12214;
wire S12215;
wire S12216;
wire S12217;
wire S12218;
wire S12219;
wire S12220;
wire S12221;
wire S12222;
wire S12223;
wire S12224;
wire S12225;
wire S12226;
wire S12227;
wire S12228;
wire S12229;
wire S12230;
wire S12231;
wire S12232;
wire S12233;
wire S12234;
wire S12235;
wire S12236;
wire S12237;
wire S12238;
wire S12239;
wire S12240;
wire S12241;
wire S12242;
wire S12243;
wire S12244;
wire S12245;
wire S12246;
wire S12247;
wire S12248;
wire S12249;
wire S12250;
wire S12251;
wire S12252;
wire S12253;
wire S12254;
wire S12255;
wire S12256;
wire S12257;
wire S12258;
wire S12259;
wire S12260;
wire S12261;
wire S12262;
wire S12263;
wire S12264;
wire S12265;
wire S12266;
wire S12267;
wire S12268;
wire S12269;
wire S12270;
wire S12271;
wire S12272;
wire S12273;
wire S12274;
wire S12275;
wire S12276;
wire S12277;
wire S12278;
wire S12279;
wire S12280;
wire S12281;
wire S12282;
wire S12283;
wire S12284;
wire S12285;
wire S12286;
wire S12287;
wire S12288;
wire S12289;
wire S12290;
wire S12291;
wire S12292;
wire S12293;
wire S12294;
wire S12295;
wire S12296;
wire S12297;
wire S12298;
wire S12299;
wire S12300;
wire S12301;
wire S12302;
wire S12303;
wire S12304;
wire S12305;
wire S12306;
wire S12307;
wire S12308;
wire S12309;
wire S12310;
wire S12311;
wire S12312;
wire S12313;
wire S12314;
wire S12315;
wire S12316;
wire S12317;
wire S12318;
wire S12319;
wire S12320;
wire S12321;
wire S12322;
wire S12323;
wire S12324;
wire S12325;
wire S12326;
wire S12327;
wire S12328;
wire S12329;
wire S12330;
wire S12331;
wire S12332;
wire S12333;
wire S12334;
wire S12335;
wire S12336;
wire S12337;
wire S12338;
wire S12339;
wire S12340;
wire S12341;
wire S12342;
wire S12343;
wire S12344;
wire S12345;
wire S12346;
wire S12347;
wire S12348;
wire S12349;
wire S12350;
wire S12351;
wire S12352;
wire S12353;
wire S12354;
wire S12355;
wire S12356;
wire S12357;
wire S12358;
wire S12359;
wire S12360;
wire S12361;
wire S12362;
wire S12363;
wire S12364;
wire S12365;
wire S12366;
wire S12367;
wire S12368;
wire S12369;
wire S12370;
wire S12371;
wire S12372;
wire S12373;
wire S12374;
wire S12375;
wire S12376;
wire S12377;
wire S12378;
wire S12379;
wire S12380;
wire S12381;
wire S12382;
wire S12383;
wire S12384;
wire S12385;
wire S12386;
wire S12387;
wire S12388;
wire S12389;
wire S12390;
wire S12391;
wire S12392;
wire S12393;
wire S12394;
wire S12395;
wire S12396;
wire S12397;
wire S12398;
wire S12399;
wire S12400;
wire S12401;
wire S12402;
wire S12403;
wire S12404;
wire S12405;
wire S12406;
wire S12407;
wire S12408;
wire S12409;
wire S12410;
wire S12411;
wire S12412;
wire S12413;
wire S12414;
wire S12415;
wire S12416;
wire S12417;
wire S12418;
wire S12419;
wire S12420;
wire S12421;
wire S12422;
wire S12423;
wire S12424;
wire S12425;
wire S12426;
wire S12427;
wire S12428;
wire S12429;
wire S12430;
wire S12431;
wire S12432;
wire S12433;
wire S12434;
wire S12435;
wire S12436;
wire S12437;
wire S12438;
wire S12439;
wire S12440;
wire S12441;
wire S12442;
wire S12443;
wire S12444;
wire S12445;
wire S12446;
wire S12447;
wire S12448;
wire S12449;
wire S12450;
wire S12451;
wire S12452;
wire S12453;
wire S12454;
wire S12455;
wire S12456;
wire S12457;
wire S12458;
wire S12459;
wire S12460;
wire S12461;
wire S12462;
wire S12463;
wire S12464;
wire S12465;
wire S12466;
wire S12467;
wire S12468;
wire S12469;
wire S12470;
wire S12471;
wire S12472;
wire S12473;
wire S12474;
wire S12475;
wire S12476;
wire S12477;
wire S12478;
wire S12479;
wire S12480;
wire S12481;
wire S12482;
wire S12483;
wire S12484;
wire S12485;
wire S12486;
wire S12487;
wire S12488;
wire S12489;
wire S12490;
wire S12491;
wire S12492;
wire S12493;
wire S12494;
wire S12495;
wire S12496;
wire S12497;
wire S12498;
wire S12499;
wire S12500;
wire S12501;
wire S12502;
wire S12503;
wire S12504;
wire S12505;
wire S12506;
wire S12507;
wire S12508;
wire S12509;
wire S12510;
wire S12511;
wire S12512;
wire S12513;
wire S12514;
wire S12515;
wire S12516;
wire S12517;
wire S12518;
wire S12519;
wire S12520;
wire S12521;
wire S12522;
wire S12523;
wire S12524;
wire S12525;
wire S12526;
wire S12527;
wire S12528;
wire S12529;
wire S12530;
wire S12531;
wire S12532;
wire S12533;
wire S12534;
wire S12535;
wire S12536;
wire S12537;
wire S12538;
wire S12539;
wire S12540;
wire S12541;
wire S12542;
wire S12543;
wire S12544;
wire S12545;
wire S12546;
wire S12547;
wire S12548;
wire S12549;
wire S12550;
wire S12551;
wire S12552;
wire S12553;
wire S12554;
wire S12555;
wire S12556;
wire S12557;
wire S12558;
wire S12559;
wire S12560;
wire S12561;
wire S12562;
wire S12563;
wire S12564;
wire S12565;
wire S12566;
wire S12567;
wire S12568;
wire S12569;
wire S12570;
wire S12571;
wire S12572;
wire S12573;
wire S12574;
wire S12575;
wire S12576;
wire S12577;
wire S12578;
wire S12579;
wire S12580;
wire S12581;
wire S12582;
wire S12583;
wire S12584;
wire S12585;
wire S12586;
wire S12587;
wire S12588;
wire S12589;
wire S12590;
wire S12591;
wire S12592;
wire S12593;
wire S12594;
wire S12595;
wire S12596;
wire S12597;
wire S12598;
wire S12599;
wire S12600;
wire S12601;
wire S12602;
wire S12603;
wire S12604;
wire S12605;
wire S12606;
wire S12607;
wire S12608;
wire S12609;
wire S12610;
wire S12611;
wire S12612;
wire S12613;
wire S12614;
wire S12615;
wire S12616;
wire S12617;
wire S12618;
wire S12619;
wire S12620;
wire S12621;
wire S12622;
wire S12623;
wire S12624;
wire S12625;
wire S12626;
wire S12627;
wire S12628;
wire S12629;
wire S12630;
wire S12631;
wire S12632;
wire S12633;
wire S12634;
wire S12635;
wire S12636;
wire S12637;
wire S12638;
wire S12639;
wire S12640;
wire S12641;
wire S12642;
wire S12643;
wire S12644;
wire S12645;
wire S12646;
wire S12647;
wire S12648;
wire S12649;
wire S12650;
wire S12651;
wire S12652;
wire S12653;
wire S12654;
wire S12655;
wire S12656;
wire S12657;
wire S12658;
wire S12659;
wire S12660;
wire S12661;
wire S12662;
wire S12663;
wire S12664;
wire S12665;
wire S12666;
wire S12667;
wire S12668;
wire S12669;
wire S12670;
wire S12671;
wire S12672;
wire S12673;
wire S12674;
wire S12675;
wire S12676;
wire S12677;
wire S12678;
wire S12679;
wire S12680;
wire S12681;
wire S12682;
wire S12683;
wire S12684;
wire S12685;
wire S12686;
wire S12687;
wire S12688;
wire S12689;
wire S12690;
wire S12691;
wire S12692;
wire S12693;
wire S12694;
wire S12695;
wire S12696;
wire S12697;
wire S12698;
wire S12699;
wire S12700;
wire S12701;
wire S12702;
wire S12703;
wire S12704;
wire S12705;
wire S12706;
wire S12707;
wire S12708;
wire S12709;
wire S12710;
wire S12711;
wire S12712;
wire S12713;
wire S12714;
wire S12715;
wire S12716;
wire S12717;
wire S12718;
wire S12719;
wire S12720;
wire S12721;
wire S12722;
wire S12723;
wire S12724;
wire S12725;
wire S12726;
wire S12727;
wire S12728;
wire S12729;
wire S12730;
wire S12731;
wire S12732;
wire S12733;
wire S12734;
wire S12735;
wire S12736;
wire S12737;
wire S12738;
wire S12739;
wire S12740;
wire S12741;
wire S12742;
wire S12743;
wire S12744;
wire S12745;
wire S12746;
wire S12747;
wire S12748;
wire S12749;
wire S12750;
wire S12751;
wire S12752;
wire S12753;
wire S12754;
wire S12755;
wire S12756;
wire S12757;
wire S12758;
wire S12759;
wire S12760;
wire S12761;
wire S12762;
wire S12763;
wire S12764;
wire S12765;
wire S12766;
wire S12767;
wire S12768;
wire S12769;
wire S12770;
wire S12771;
wire S12772;
wire S12773;
wire S12774;
wire S12775;
wire S12776;
wire S12777;
wire S12778;
wire S12779;
wire S12780;
wire S12781;
wire S12782;
wire S12783;
wire S12784;
wire S12785;
wire S12786;
wire S12787;
wire S12788;
wire S12789;
wire S12790;
wire S12791;
wire S12792;
wire S12793;
wire S12794;
wire S12795;
wire S12796;
wire S12797;
wire S12798;
wire S12799;
wire S12800;
wire S12801;
wire S12802;
wire S12803;
wire S12804;
wire S12805;
wire S12806;
wire S12807;
wire S12808;
wire S12809;
wire S12810;
wire S12811;
wire S12812;
wire S12813;
wire S12814;
wire S12815;
wire S12816;
wire S12817;
wire S12818;
wire S12819;
wire S12820;
wire S12821;
wire S12822;
wire S12823;
wire S12824;
wire S12825;
wire S12826;
wire S12827;
wire S12828;
wire S12829;
wire S12830;
wire S12831;
wire S12832;
wire S12833;
wire S12834;
wire S12835;
wire S12836;
wire S12837;
wire S12838;
wire S12839;
wire S12840;
wire S12841;
wire S12842;
wire S12843;
wire S12844;
wire S12845;
wire S12846;
wire S12847;
wire S12848;
wire S12849;
wire S12850;
wire S12851;
wire S12852;
wire S12853;
wire S12854;
wire S12855;
wire S12856;
wire S12857;
wire S12858;
wire S12859;
wire S12860;
wire S12861;
wire S12862;
wire S12863;
wire S12864;
wire S12865;
wire S12866;
wire S12867;
wire S12868;
wire S12869;
wire S12870;
wire S12871;
wire S12872;
wire S12873;
wire S12874;
wire S12875;
wire S12876;
wire S12877;
wire S12878;
wire S12879;
wire S12880;
wire S12881;
wire S12882;
wire S12883;
wire S12884;
wire S12885;
wire S12886;
wire S12887;
wire S12888;
wire S12889;
wire S12890;
wire S12891;
wire S12892;
wire S12893;
wire S12894;
wire S12895;
wire S12896;
wire S12897;
wire S12898;
wire S12899;
wire S12900;
wire S12901;
wire S12902;
wire S12903;
wire S12904;
wire S12905;
wire S12906;
wire S12907;
wire S12908;
wire S12909;
wire S12910;
wire S12911;
wire S12912;
wire S12913;
wire S12914;
wire S12915;
wire S12916;
wire S12917;
wire S12918;
wire S12919;
wire S12920;
wire S12921;
wire S12922;
wire S12923;
wire S12924;
wire S12925;
wire S12926;
wire S12927;
wire S12928;
wire S12929;
wire S12930;
wire S12931;
wire S12932;
wire S12933;
wire S12934;
wire S12935;
wire S12936;
wire S12937;
wire S12938;
wire S12939;
wire S12940;
wire S12941;
wire S12942;
wire S12943;
wire S12944;
wire S12945;
wire S12946;
wire S12947;
wire S12948;
wire S12949;
wire S12950;
wire S12951;
wire S12952;
wire S12953;
wire S12954;
wire S12955;
wire S12956;
wire S12957;
wire S12958;
wire S12959;
wire S12960;
wire S12961;
wire S12962;
wire S12963;
wire S12964;
wire S12965;
wire S12966;
wire S12967;
wire S12968;
wire S12969;
wire S12970;
wire S12971;
wire S12972;
wire S12973;
wire S12974;
wire S12975;
wire S12976;
wire S12977;
wire S12978;
wire S12979;
wire S12980;
wire S12981;
wire S12982;
wire S12983;
wire S12984;
wire S12985;
wire S12986;
wire S12987;
wire S12988;
wire S12989;
wire S12990;
wire S12991;
wire S12992;
wire S12993;
wire S12994;
wire S12995;
wire S12996;
wire S12997;
wire S12998;
wire S12999;
wire S13000;
wire S13001;
wire S13002;
wire S13003;
wire S13004;
wire S13005;
wire S13006;
wire S13007;
wire S13008;
wire S13009;
wire S13010;
wire S13011;
wire S13012;
wire S13013;
wire S13014;
wire S13015;
wire S13016;
wire S13017;
wire S13018;
wire S13019;
wire S13020;
wire S13021;
wire S13022;
wire S13023;
wire S13024;
wire S13025;
wire S13026;
wire S13027;
wire S13028;
wire S13029;
wire S13030;
wire S13031;
wire S13032;
wire S13033;
wire S13034;
wire S13035;
wire S13036;
wire S13037;
wire S13038;
wire S13039;
wire S13040;
wire S13041;
wire S13042;
wire S13043;
wire S13044;
wire S13045;
wire S13046;
wire S13047;
wire S13048;
wire S13049;
wire S13050;
wire S13051;
wire S13052;
wire S13053;
wire S13054;
wire S13055;
wire S13056;
wire S13057;
wire S13058;
wire S13059;
wire S13060;
wire S13061;
wire S13062;
wire S13063;
wire S13064;
wire S13065;
wire S13066;
wire S13067;
wire S13068;
wire S13069;
wire S13070;
wire S13071;
wire S13072;
wire S13073;
wire S13074;
wire S13075;
wire S13076;
wire S13077;
wire S13078;
wire S13079;
wire S13080;
wire S13081;
wire S13082;
wire S13083;
wire S13084;
wire S13085;
wire S13086;
wire S13087;
wire S13088;
wire S13089;
wire S13090;
wire S13091;
wire S13092;
wire S13093;
wire S13094;
wire S13095;
wire S13096;
wire S13097;
wire S13098;
wire S13099;
wire S13100;
wire S13101;
wire S13102;
wire S13103;
wire S13104;
wire S13105;
wire S13106;
wire S13107;
wire S13108;
wire S13109;
wire S13110;
wire S13111;
wire S13112;
wire S13113;
wire S13114;
wire S13115;
wire S13116;
wire S13117;
wire S13118;
wire S13119;
wire S13120;
wire S13121;
wire S13122;
wire S13123;
wire S13124;
wire S13125;
wire S13126;
wire S13127;
wire S13128;
wire S13129;
wire S13130;
wire S13131;
wire S13132;
wire S13133;
wire S13134;
wire S13135;
wire S13136;
wire S13137;
wire S13138;
wire S13139;
wire S13140;
wire S13141;
wire S13142;
wire S13143;
wire S13144;
wire S13145;
wire S13146;
wire S13147;
wire S13148;
wire S13149;
wire S13150;
wire S13151;
wire S13152;
wire S13153;
wire S13154;
wire S13155;
wire S13156;
wire S13157;
wire S13158;
wire S13159;
wire S13160;
wire S13161;
wire S13162;
wire S13163;
wire S13164;
wire S13165;
wire S13166;
wire S13167;
wire S13168;
wire S13169;
wire S13170;
wire S13171;
wire S13172;
wire S13173;
wire S13174;
wire S13175;
wire S13176;
wire S13177;
wire S13178;
wire S13179;
wire S13180;
wire S13181;
wire S13182;
wire S13183;
wire S13184;
wire S13185;
wire S13186;
wire S13187;
wire S13188;
wire S13189;
wire S13190;
wire S13191;
wire S13192;
wire S13193;
wire S13194;
wire S13195;
wire S13196;
wire S13197;
wire S13198;
wire S13199;
wire S13200;
wire S13201;
wire S13202;
wire S13203;
wire S13204;
wire S13205;
wire S13206;
wire S13207;
wire S13208;
wire S13209;
wire S13210;
wire S13211;
wire S13212;
wire S13213;
wire S13214;
wire S13215;
wire S13216;
wire S13217;
wire S13218;
wire S13219;
wire S13220;
wire S13221;
wire S13222;
wire S13223;
wire S13224;
wire S13225;
wire S13226;
wire S13227;
wire S13228;
wire S13229;
wire S13230;
wire S13231;
wire S13232;
wire S13233;
wire S13234;
wire S13235;
wire S13236;
wire S13237;
wire S13238;
wire S13239;
wire S13240;
wire S13241;
wire S13242;
wire S13243;
wire S13244;
wire S13245;
wire S13246;
wire S13247;
wire S13248;
wire S13249;
wire S13250;
wire S13251;
wire S13252;
wire S13253;
wire S13254;
wire S13255;
wire S13256;
wire S13257;
wire S13258;
wire S13259;
wire S13260;
wire S13261;
wire S13262;
wire S13263;
wire S13264;
wire S13265;
wire S13266;
wire S13267;
wire S13268;
wire S13269;
wire S13270;
wire S13271;
wire S13272;
wire S13273;
wire S13274;
wire S13275;
wire S13276;
wire S13277;
wire S13278;
wire S13279;
wire S13280;
wire S13281;
wire S13282;
wire S13283;
wire S13284;
wire S13285;
wire S13286;
wire S13287;
wire S13288;
wire S13289;
wire S13290;
wire S13291;
wire S13292;
wire S13293;
wire S13294;
wire S13295;
wire S13296;
wire S13297;
wire S13298;
wire S13299;
wire S13300;
wire S13301;
wire S13302;
wire S13303;
wire S13304;
wire S13305;
wire S13306;
wire S13307;
wire S13308;
wire S13309;
wire S13310;
wire S13311;
wire S13312;
wire S13313;
wire S13314;
wire S13315;
wire S13316;
wire S13317;
wire S13318;
wire S13319;
wire S13320;
wire S13321;
wire S13322;
wire S13323;
wire S13324;
wire S13325;
wire S13326;
wire S13327;
wire S13328;
wire S13329;
wire S13330;
wire S13331;
wire S13332;
wire S13333;
wire S13334;
wire S13335;
wire S13336;
wire S13337;
wire S13338;
wire S13339;
wire S13340;
wire S13341;
wire S13342;
wire S13343;
wire S13344;
wire S13345;
wire S13346;
wire S13347;
wire S13348;
wire S13349;
wire S13350;
wire S13351;
wire S13352;
wire S13353;
wire S13354;
wire S13355;
wire S13356;
wire S13357;
wire S13358;
wire S13359;
wire S13360;
wire S13361;
wire S13362;
wire S13363;
wire S13364;
wire S13365;
wire S13366;
wire S13367;
wire S13368;
wire S13369;
wire S13370;
wire S13371;
wire S13372;
wire S13373;
wire S13374;
wire S13375;
wire S13376;
wire S13377;
wire S13378;
wire S13379;
wire S13380;
wire S13381;
wire S13382;
wire S13383;
wire S13384;
wire S13385;
wire S13386;
wire S13387;
wire S13388;
wire S13389;
wire S13390;
wire S13391;
wire S13392;
wire S13393;
wire S13394;
wire S13395;
wire S13396;
wire S13397;
wire S13398;
wire S13399;
wire S13400;
wire S13401;
wire S13402;
wire S13403;
wire S13404;
wire S13405;
wire S13406;
wire S13407;
wire S13408;
wire S13409;
wire S13410;
wire S13411;
wire S13412;
wire S13413;
wire S13414;
wire S13415;
wire S13416;
wire S13417;
wire S13418;
wire S13419;
wire S13420;
wire S13421;
wire S13422;
wire S13423;
wire S13424;
wire S13425;
wire S13426;
wire S13427;
wire S13428;
wire S13429;
wire S13430;
wire S13431;
wire S13432;
wire S13433;
wire S13434;
wire S13435;
wire S13436;
wire S13437;
wire S13438;
wire S13439;
wire S13440;
wire S13441;
wire S13442;
wire S13443;
wire S13444;
wire S13445;
wire S13446;
wire S13447;
wire S13448;
wire S13449;
wire S13450;
wire S13451;
wire S13452;
wire S13453;
wire S13454;
wire S13455;
wire S13456;
wire S13457;
wire S13458;
wire S13459;
wire S13460;
wire S13461;
wire S13462;
wire S13463;
wire S13464;
wire S13465;
wire S13466;
wire S13467;
wire S13468;
wire S13469;
wire S13470;
wire S13471;
wire S13472;
wire S13473;
wire S13474;
wire S13475;
wire S13476;
wire S13477;
wire S13478;
wire S13479;
wire S13480;
wire S13481;
wire S13482;
wire S13483;
wire S13484;
wire S13485;
wire S13486;
wire S13487;
wire S13488;
wire S13489;
wire S13490;
wire S13491;
wire S13492;
wire S13493;
wire S13494;
wire S13495;
wire S13496;
wire S13497;
wire S13498;
wire S13499;
wire S13500;
wire S13501;
wire S13502;
wire S13503;
wire S13504;
wire S13505;
wire S13506;
wire S13507;
wire S13508;
wire S13509;
wire S13510;
wire S13511;
wire S13512;
wire S13513;
wire S13514;
wire S13515;
wire S13516;
wire S13517;
wire S13518;
wire S13519;
wire S13520;
wire S13521;
wire S13522;
wire S13523;
wire S13524;
wire S13525;
wire S13526;
wire S13527;
wire S13528;
wire S13529;
wire S13530;
wire S13531;
wire S13532;
wire S13533;
wire S13534;
wire S13535;
wire S13536;
wire S13537;
wire S13538;
wire S13539;
wire S13540;
wire S13541;
wire S13542;
wire S13543;
wire S13544;
wire S13545;
wire S13546;
wire S13547;
wire S13548;
wire S13549;
wire S13550;
wire S13551;
wire S13552;
wire S13553;
wire S13554;
wire S13555;
wire S13556;
wire S13557;
wire S13558;
wire S13559;
wire S13560;
wire S13561;
wire S13562;
wire S13563;
wire S13564;
wire S13565;
wire S13566;
wire S13567;
wire S13568;
wire S13569;
wire S13570;
wire S13571;
wire S13572;
wire S13573;
wire S13574;
wire S13575;
wire S13576;
wire S13577;
wire S13578;
wire S13579;
wire S13580;
wire S13581;
wire S13582;
wire S13583;
wire S13584;
wire S13585;
wire S13586;
wire S13587;
wire S13588;
wire S13589;
wire S13590;
wire S13591;
wire S13592;
wire S13593;
wire S13594;
wire S13595;
wire S13596;
wire S13597;
wire S13598;
wire S13599;
wire S13600;
wire S13601;
wire S13602;
wire S13603;
wire S13604;
wire S13605;
wire S13606;
wire S13607;
wire S13608;
wire S13609;
wire S13610;
wire S13611;
wire S13612;
wire S13613;
wire S13614;
wire S13615;
wire S13616;
wire S13617;
wire S13618;
wire S13619;
wire S13620;
wire S13621;
wire S13622;
wire S13623;
wire S13624;
wire S13625;
wire S13626;
wire S13627;
wire S13628;
wire S13629;
wire S13630;
wire S13631;
wire S13632;
wire S13633;
wire S13634;
wire S13635;
wire S13636;
wire S13637;
wire S13638;
wire S13639;
wire S13640;
wire S13641;
wire S13642;
wire S13643;
wire S13644;
wire S13645;
wire S13646;
wire S13647;
wire S13648;
wire S13649;
wire S13650;
wire S13651;
wire S13652;
wire S13653;
wire S13654;
wire S13655;
wire S13656;
wire S13657;
wire S13658;
wire S13659;
wire S13660;
wire S13661;
wire S13662;
wire S13663;
wire S13664;
wire S13665;
wire S13666;
wire S13667;
wire S13668;
wire S13669;
wire S13670;
wire S13671;
wire S13672;
wire S13673;
wire S13674;
wire S13675;
wire S13676;
wire S13677;
wire S13678;
wire S13679;
wire S13680;
wire S13681;
wire S13682;
wire S13683;
wire S13684;
wire S13685;
wire S13686;
wire S13687;
wire S13688;
wire S13689;
wire S13690;
wire S13691;
wire S13692;
wire S13693;
wire S13694;
wire S13695;
wire S13696;
wire S13697;
wire S13698;
wire S13699;
wire S13700;
wire S13701;
wire S13702;
wire S13703;
wire S13704;
wire S13705;
wire S13706;
wire S13707;
wire S13708;
wire S13709;
wire S13710;
wire S13711;
wire S13712;
wire S13713;
wire S13714;
wire S13715;
wire S13716;
wire S13717;
wire S13718;
wire S13719;
wire S13720;
wire S13721;
wire S13722;
wire S13723;
wire S13724;
wire S13725;
wire S13726;
wire S13727;
wire S13728;
wire S13729;
wire S13730;
wire S13731;
wire S13732;
wire S13733;
wire S13734;
wire S13735;
wire S13736;
wire S13737;
wire S13738;
wire S13739;
wire S13740;
wire S13741;
wire S13742;
wire S13743;
wire S13744;
wire S13745;
wire S13746;
wire S13747;
wire S13748;
wire S13749;
wire S13750;
wire S13751;
wire S13752;
wire S13753;
wire S13754;
wire S13755;
wire S13756;
wire S13757;
wire S13758;
wire S13759;
wire S13760;
wire S13761;
wire S13762;
wire S13763;
wire S13764;
wire S13765;
wire S13766;
wire S13767;
wire S13768;
wire S13769;
wire S13770;
wire S13771;
wire S13772;
wire S13773;
wire S13774;
wire S13775;
wire S13776;
wire S13777;
wire S13778;
wire S13779;
wire S13780;
wire S13781;
wire S13782;
wire S13783;
wire S13784;
wire S13785;
wire S13786;
wire S13787;
wire S13788;
wire S13789;
wire S13790;
wire S13791;
wire S13792;
wire S13793;
wire S13794;
wire S13795;
wire S13796;
wire S13797;
wire S13798;
wire S13799;
wire S13800;
wire S13801;
wire S13802;
wire S13803;
wire S13804;
wire S13805;
wire S13806;
wire S13807;
wire S13808;
wire S13809;
wire S13810;
wire S13811;
wire S13812;
wire S13813;
wire S13814;
wire S13815;
wire S13816;
wire S13817;
wire S13818;
wire S13819;
wire S13820;
wire S13821;
wire S13822;
wire S13823;
wire S13824;
wire S13825;
wire S13826;
wire S13827;
wire S13828;
wire S13829;
wire S13830;
wire S13831;
wire S13832;
wire S13833;
wire S13834;
wire S13835;
wire S13836;
wire S13837;
wire S13838;
wire S13839;
wire S13840;
wire S13841;
wire S13842;
wire S13843;
wire S13844;
wire S13845;
wire S13846;
wire S13847;
wire S13848;
wire S13849;
wire S13850;
wire S13851;
wire S13852;
wire S13853;
wire S13854;
wire S13855;
wire S13856;
wire S13857;
wire S13858;
wire S13859;
wire S13860;
wire S13861;
wire S13862;
wire S13863;
wire S13864;
wire S13865;
wire S13866;
wire S13867;
wire S13868;
wire S13869;
wire S13870;
wire S13871;
wire S13872;
wire S13873;
wire S13874;
wire S13875;
wire S13876;
wire S13877;
wire S13878;
wire S13879;
wire S13880;
wire S13881;
wire S13882;
wire S13883;
wire S13884;
wire S13885;
wire S13886;
wire S13887;
wire S13888;
wire S13889;
wire S13890;
wire S13891;
wire S13892;
wire S13893;
wire S13894;
wire S13895;
wire S13896;
wire S13897;
wire S13898;
wire S13899;
wire S13900;
wire S13901;
wire S13902;
wire S13903;
wire S13904;
wire S13905;
wire S13906;
wire S13907;
wire S13908;
wire S13909;
wire S13910;
wire S13911;
wire S13912;
wire S13913;
wire S13914;
wire S13915;
wire S13916;
wire S13917;
wire S13918;
wire S13919;
wire S13920;
wire S13921;
wire S13922;
wire S13923;
wire S13924;
wire S13925;
wire S13926;
wire S13927;
wire S13928;
wire S13929;
wire S13930;
wire S13931;
wire S13932;
wire S13933;
wire S13934;
wire S13935;
wire S13936;
wire S13937;
wire S13938;
wire S13939;
wire S13940;
wire S13941;
wire S13942;
wire S13943;
wire S13944;
wire S13945;
wire S13946;
wire S13947;
wire S13948;
wire S13949;
wire S13950;
wire S13951;
wire S13952;
wire S13953;
wire S13954;
wire S13955;
wire S13956;
wire S13957;
wire S13958;
wire S13959;
wire S13960;
wire S13961;
wire S13962;
wire S13963;
wire S13964;
wire S13965;
wire S13966;
wire S13967;
wire S13968;
wire S13969;
wire S13970;
wire S13971;
wire S13972;
wire S13973;
wire S13974;
wire S13975;
wire S13976;
wire S13977;
wire S13978;
wire S13979;
wire S13980;
wire S13981;
wire S13982;
wire S13983;
wire S13984;
wire S13985;
wire S13986;
wire S13987;
wire S13988;
wire S13989;
wire S13990;
wire S13991;
wire S13992;
wire S13993;
wire S13994;
wire S13995;
wire S13996;
wire S13997;
wire S13998;
wire S13999;
wire S14000;
wire S14001;
wire S14002;
wire S14003;
wire S14004;
wire S14005;
wire S14006;
wire S14007;
wire S14008;
wire S14009;
wire S14010;
wire S14011;
wire S14012;
wire S14013;
wire S14014;
wire S14015;
wire S14016;
wire S14017;
wire S14018;
wire S14019;
wire S14020;
wire S14021;
wire S14022;
wire S14023;
wire S14024;
wire S14025;
wire S14026;
wire S14027;
wire S14028;
wire S14029;
wire S14030;
wire S14031;
wire S14032;
wire S14033;
wire S14034;
wire S14035;
wire S14036;
wire S14037;
wire S14038;
wire S14039;
wire S14040;
wire S14041;
wire S14042;
wire S14043;
wire S14044;
wire S14045;
wire S14046;
wire S14047;
wire S14048;
wire S14049;
wire S14050;
wire S14051;
wire S14052;
wire S14053;
wire S14054;
wire S14055;
wire S14056;
wire S14057;
wire S14058;
wire S14059;
wire S14060;
wire S14061;
wire S14062;
wire S14063;
wire S14064;
wire S14065;
wire S14066;
wire S14067;
wire S14068;
wire S14069;
wire S14070;
wire S14071;
wire S14072;
wire S14073;
wire S14074;
wire S14075;
wire S14076;
wire S14077;
wire S14078;
wire S14079;
wire S14080;
wire S14081;
wire S14082;
wire S14083;
wire S14084;
wire S14085;
wire S14086;
wire S14087;
wire S14088;
wire S14089;
wire S14090;
wire S14091;
wire S14092;
wire S14093;
wire S14094;
wire S14095;
wire S14096;
wire S14097;
wire S14098;
wire S14099;
wire S14100;
wire S14101;
wire S14102;
wire S14103;
wire S14104;
wire S14105;
wire S14106;
wire S14107;
wire S14108;
wire S14109;
wire S14110;
wire S14111;
wire S14112;
wire S14113;
wire S14114;
wire S14115;
wire S14116;
wire S14117;
wire S14118;
wire S14119;
wire S14120;
wire S14121;
wire S14122;
wire S14123;
wire S14124;
wire S14125;
wire S14126;
wire S14127;
wire S14128;
wire S14129;
wire S14130;
wire S14131;
wire S14132;
wire S14133;
wire S14134;
wire S14135;
wire S14136;
wire S14137;
wire S14138;
wire S14139;
wire S14140;
wire S14141;
wire S14142;
wire S14143;
wire S14144;
wire S14145;
wire S14146;
wire S14147;
wire S14148;
wire S14149;
wire S14150;
wire S14151;
wire S14152;
wire S14153;
wire S14154;
wire S14155;
wire S14156;
wire S14157;
wire S14158;
wire S14159;
wire S14160;
wire S14161;
wire S14162;
wire S14163;
wire S14164;
wire S14165;
wire S14166;
wire S14167;
wire S14168;
wire S14169;
wire S14170;
wire S14171;
wire S14172;
wire S14173;
wire S14174;
wire S14175;
wire S14176;
wire S14177;
wire S14178;
wire S14179;
wire S14180;
wire S14181;
wire S14182;
wire S14183;
wire S14184;
wire S14185;
wire S14186;
wire S14187;
wire S14188;
wire S14189;
wire S14190;
wire S14191;
wire S14192;
wire S14193;
wire S14194;
wire S14195;
wire S14196;
wire S14197;
wire S14198;
wire S14199;
wire S14200;
wire S14201;
wire S14202;
wire S14203;
wire S14204;
wire S14205;
wire S14206;
wire S14207;
wire S14208;
wire S14209;
wire S14210;
wire S14211;
wire S14212;
wire S14213;
wire S14214;
wire S14215;
wire S14216;
wire S14217;
wire S14218;
wire S14219;
wire S14220;
wire S14221;
wire S14222;
wire S14223;
wire S14224;
wire S14225;
wire S14226;
wire S14227;
wire S14228;
wire S14229;
wire S14230;
wire S14231;
wire S14232;
wire S14233;
wire S14234;
wire S14235;
wire S14236;
wire S14237;
wire S14238;
wire S14239;
wire S14240;
wire S14241;
wire S14242;
wire S14243;
wire S14244;
wire S14245;
wire S14246;
wire S14247;
wire S14248;
wire S14249;
wire S14250;
wire S14251;
wire S14252;
wire S14253;
wire S14254;
wire S14255;
wire S14256;
wire S14257;
wire S14258;
wire S14259;
wire S14260;
wire S14261;
wire S14262;
wire S14263;
wire S14264;
wire S14265;
wire S14266;
wire S14267;
wire S14268;
wire S14269;
wire S14270;
wire S14271;
wire S14272;
wire S14273;
wire S14274;
wire S14275;
wire S14276;
wire S14277;
wire S14278;
wire S14279;
wire S14280;
wire S14281;
wire S14282;
wire S14283;
wire S14284;
wire S14285;
wire S14286;
wire S14287;
wire S14288;
wire S14289;
wire S14290;
wire S14291;
wire S14292;
wire S14293;
wire S14294;
wire S14295;
wire S14296;
wire S14297;
wire S14298;
wire S14299;
wire S14300;
wire S14301;
wire S14302;
wire S14303;
wire S14304;
wire S14305;
wire S14306;
wire S14307;
wire S14308;
wire S14309;
wire S14310;
wire S14311;
wire S14312;
wire S14313;
wire S14314;
wire S14315;
wire S14316;
wire S14317;
wire S14318;
wire S14319;
wire S14320;
wire S14321;
wire S14322;
wire S14323;
wire S14324;
wire S14325;
wire S14326;
wire S14327;
wire S14328;
wire S14329;
wire S14330;
wire S14331;
wire S14332;
wire S14333;
wire S14334;
wire S14335;
wire S14336;
wire S14337;
wire S14338;
wire S14339;
wire S14340;
wire S14341;
wire S14342;
wire S14343;
wire S14344;
wire S14345;
wire S14346;
wire S14347;
wire S14348;
wire S14349;
wire S14350;
wire S14351;
wire S14352;
wire S14353;
wire S14354;
wire S14355;
wire S14356;
wire S14357;
wire S14358;
wire S14359;
wire S14360;
wire S14361;
wire S14362;
wire S14363;
wire S14364;
wire S14365;
wire S14366;
wire S14367;
wire S14368;
wire S14369;
wire S14370;
wire S14371;
wire S14372;
wire S14373;
wire S14374;
wire S14375;
wire S14376;
wire S14377;
wire S14378;
wire S14379;
wire S14380;
wire S14381;
wire S14382;
wire S14383;
wire S14384;
wire S14385;
wire S14386;
wire S14387;
wire S14388;
wire S14389;
wire S14390;
wire S14391;
wire S14392;
wire S14393;
wire S14394;
wire S14395;
wire S14396;
wire S14397;
wire S14398;
wire S14399;
wire S14400;
wire S14401;
wire S14402;
wire S14403;
wire S14404;
wire S14405;
wire S14406;
wire S14407;
wire S14408;
wire S14409;
wire S14410;
wire S14411;
wire S14412;
wire S14413;
wire S14414;
wire S14415;
wire S14416;
wire S14417;
wire S14418;
wire S14419;
wire S14420;
wire S14421;
wire S14422;
wire S14423;
wire S14424;
wire S14425;
wire S14426;
wire S14427;
wire S14428;
wire S14429;
wire S14430;
wire S14431;
wire S14432;
wire S14433;
wire S14434;
wire S14435;
wire S14436;
wire S14437;
wire S14438;
wire S14439;
wire S14440;
wire S14441;
wire S14442;
wire S14443;
wire S14444;
wire S14445;
wire S14446;
wire S14447;
wire S14448;
wire S14449;
wire S14450;
wire S14451;
wire S14452;
wire S14453;
wire S14454;
wire S14455;
wire S14456;
wire S14457;
wire S14458;
wire S14459;
wire S14460;
wire S14461;
wire S14462;
wire S14463;
wire S14464;
wire S14465;
wire S14466;
wire S14467;
wire S14468;
wire S14469;
wire S14470;
wire S14471;
wire S14472;
wire S14473;
wire S14474;
wire S14475;
wire S14476;
wire S14477;
wire S14478;
wire S14479;
wire S14480;
wire S14481;
wire S14482;
wire S14483;
wire S14484;
wire S14485;
wire S14486;
wire S14487;
wire S14488;
wire S14489;
wire S14490;
wire S14491;
wire S14492;
wire S14493;
wire S14494;
wire S14495;
wire S14496;
wire S14497;
wire S14498;
wire S14499;
wire S14500;
wire S14501;
wire S14502;
wire S14503;
wire S14504;
wire S14505;
wire S14506;
wire S14507;
wire S14508;
wire S14509;
wire S14510;
wire S14511;
wire S14512;
wire S14513;
wire S14514;
wire S14515;
wire S14516;
wire S14517;
wire S14518;
wire S14519;
wire S14520;
wire S14521;
wire S14522;
wire S14523;
wire S14524;
wire S14525;
wire S14526;
wire S14527;
wire S14528;
wire S14529;
wire S14530;
wire S14531;
wire S14532;
wire S14533;
wire S14534;
wire S14535;
wire S14536;
wire S14537;
wire S14538;
wire S14539;
wire S14540;
wire S14541;
wire S14542;
wire S14543;
wire S14544;
wire S14545;
wire S14546;
wire S14547;
wire S14548;
wire S14549;
wire S14550;
wire S14551;
wire S14552;
wire S14553;
wire S14554;
wire S14555;
wire S14556;
wire S14557;
wire S14558;
wire S14559;
wire S14560;
wire S14561;
wire S14562;
wire S14563;
wire S14564;
wire S14565;
wire S14566;
wire S14567;
wire S14568;
wire S14569;
wire S14570;
wire S14571;
wire S14572;
wire S14573;
wire S14574;
wire S14575;
wire S14576;
wire S14577;
wire S14578;
wire S14579;
wire S14580;
wire S14581;
wire S14582;
wire S14583;
wire S14584;
wire S14585;
wire S14586;
wire S14587;
wire S14588;
wire S14589;
wire S14590;
wire S14591;
wire S14592;
wire S14593;
wire S14594;
wire S14595;
wire S14596;
wire S14597;
wire S14598;
wire S14599;
wire S14600;
wire S14601;
wire S14602;
wire S14603;
wire S14604;
wire S14605;
wire S14606;
wire S14607;
wire S14608;
wire S14609;
wire S14610;
wire S14611;
wire S14612;
wire S14613;
wire S14614;
wire S14615;
wire S14616;
wire S14617;
wire S14618;
wire S14619;
wire S14620;
wire S14621;
wire S14622;
wire S14623;
wire S14624;
wire S14625;
wire S14626;
wire S14627;
wire S14628;
wire S14629;
wire S14630;
wire S14631;
wire S14632;
wire S14633;
wire S14634;
wire S14635;
wire S14636;
wire S14637;
wire S14638;
wire S14639;
wire S14640;
wire S14641;
wire S14642;
wire S14643;
wire S14644;
wire S14645;
wire S14646;
wire S14647;
wire S14648;
wire S14649;
wire S14650;
wire S14651;
wire S14652;
wire S14653;
wire S14654;
wire S14655;
wire S14656;
wire S14657;
wire S14658;
wire S14659;
wire S14660;
wire S14661;
wire S14662;
wire S14663;
wire S14664;
wire S14665;
wire S14666;
wire S14667;
wire S14668;
wire S14669;
wire S14670;
wire S14671;
wire S14672;
wire S14673;
wire S14674;
wire S14675;
wire S14676;
wire S14677;
wire S14678;
wire S14679;
wire S14680;
wire S14681;
wire S14682;
wire S14683;
wire S14684;
wire S14685;
wire S14686;
wire S14687;
wire S14688;
wire S14689;
wire S14690;
wire S14691;
wire S14692;
wire S14693;
wire S14694;
wire S14695;
wire S14696;
wire S14697;
wire S14698;
wire S14699;
wire S14700;
wire S14701;
wire S14702;
wire S14703;
wire S14704;
wire S14705;
wire S14706;
wire S14707;
wire S14708;
wire S14709;
wire S14710;
wire S14711;
wire S14712;
wire S14713;
wire S14714;
wire S14715;
wire S14716;
wire S14717;
wire S14718;
wire S14719;
wire S14720;
wire S14721;
wire S14722;
wire S14723;
wire S14724;
wire S14725;
wire S14726;
wire S14727;
wire S14728;
wire S14729;
wire S14730;
wire S14731;
wire S14732;
wire S14733;
wire S14734;
wire S14735;
wire S14736;
wire S14737;
wire S14738;
wire S14739;
wire S14740;
wire S14741;
wire S14742;
wire S14743;
wire S14744;
wire S14745;
wire S14746;
wire S14747;
wire S14748;
wire S14749;
wire S14750;
wire S14751;
wire S14752;
wire S14753;
wire S14754;
wire S14755;
wire S14756;
wire S14757;
wire S14758;
wire S14759;
wire S14760;
wire S14761;
wire S14762;
wire S14763;
wire S14764;
wire S14765;
wire S14766;
wire S14767;
wire S14768;
wire S14769;
wire S14770;
wire S14771;
wire S14772;
wire S14773;
wire S14774;
wire S14775;
wire S14776;
wire S14777;
wire S14778;
wire S14779;
wire S14780;
wire S14781;
wire S14782;
wire S14783;
wire S14784;
wire S14785;
wire S14786;
wire S14787;
wire S14788;
wire S14789;
wire S14790;
wire S14791;
wire S14792;
wire S14793;
wire S14794;
wire S14795;
wire S14796;
wire S14797;
wire S14798;
wire S14799;
wire S14800;
wire S14801;
wire S14802;
wire S14803;
wire S14804;
wire S14805;
wire S14806;
wire S14807;
wire S14808;
wire S14809;
wire S14810;
wire S14811;
wire S14812;
wire S14813;
wire S14814;
wire S14815;
wire S14816;
wire S14817;
wire S14818;
wire S14819;
wire S14820;
wire S14821;
wire S14822;
wire S14823;
wire S14824;
wire S14825;
wire S14826;
wire S14827;
wire S14828;
wire S14829;
wire S14830;
wire S14831;
wire S14832;
wire S14833;
wire S14834;
wire S14835;
wire S14836;
wire S14837;
wire S14838;
wire S14839;
wire S14840;
wire S14841;
wire S14842;
wire S14843;
wire S14844;
wire S14845;
wire S14846;
wire S14847;
wire S14848;
wire S14849;
wire S14850;
wire S14851;
wire S14852;
wire S14853;
wire S14854;
wire S14855;
wire S14856;
wire S14857;
wire S14858;
wire S14859;
wire S14860;
wire S14861;
wire S14862;
wire S14863;
wire S14864;
wire S14865;
wire S14866;
wire S14867;
wire S14868;
wire S14869;
wire S14870;
wire S14871;
wire S14872;
wire S14873;
wire S14874;
wire S14875;
wire S14876;
wire S14877;
wire S14878;
wire S14879;
wire S14880;
wire S14881;
wire S14882;
wire S14883;
wire S14884;
wire S14885;
wire S14886;
wire S14887;
wire S14888;
wire S14889;
wire S14890;
wire S14891;
wire S14892;
wire S14893;
wire S14894;
wire S14895;
wire S14896;
wire S14897;
wire S14898;
wire S14899;
wire S14900;
wire S14901;
wire S14902;
wire S14903;
wire S14904;
wire S14905;
wire S14906;
wire S14907;
wire S14908;
wire S14909;
wire S14910;
wire S14911;
wire S14912;
wire S14913;
wire S14914;
wire S14915;
wire S14916;
wire S14917;
wire S14918;
wire S14919;
wire S14920;
wire S14921;
wire S14922;
wire S14923;
wire S14924;
wire S14925;
wire S14926;
wire S14927;
wire S14928;
wire S14929;
wire S14930;
wire S14931;
wire S14932;
wire S14933;
wire S14934;
wire S14935;
wire S14936;
wire S14937;
wire S14938;
wire S14939;
wire S14940;
wire S14941;
wire S14942;
wire S14943;
wire S14944;
wire S14945;
wire S14946;
wire S14947;
wire S14948;
wire S14949;
wire S14950;
wire S14951;
wire S14952;
wire S14953;
wire S14954;
wire S14955;
wire S14956;
wire S14957;
wire S14958;
wire S14959;
wire S14960;
wire S14961;
wire S14962;
wire S14963;
wire S14964;
wire S14965;
wire S14966;
wire S14967;
wire S14968;
wire S14969;
wire S14970;
wire S14971;
wire S14972;
wire S14973;
wire S14974;
wire S14975;
wire S14976;
wire S14977;
wire S14978;
wire S14979;
wire S14980;
wire S14981;
wire S14982;
wire S14983;
wire S14984;
wire S14985;
wire S14986;
wire S14987;
wire S14988;
wire S14989;
wire S14990;
wire S14991;
wire S14992;
wire S14993;
wire S14994;
wire S14995;
wire S14996;
wire S14997;
wire S14998;
wire S14999;
wire S15000;
wire S15001;
wire S15002;
wire S15003;
wire S15004;
wire S15005;
wire S15006;
wire S15007;
wire S15008;
wire S15009;
wire S15010;
wire S15011;
wire S15012;
wire S15013;
wire S15014;
wire S15015;
wire S15016;
wire S15017;
wire S15018;
wire S15019;
wire S15020;
wire S15021;
wire S15022;
wire S15023;
wire S15024;
wire S15025;
wire S15026;
wire S15027;
wire S15028;
wire S15029;
wire S15030;
wire S15031;
wire S15032;
wire S15033;
wire S15034;
wire S15035;
wire S15036;
wire S15037;
wire S15038;
wire S15039;
wire S15040;
wire S15041;
wire S15042;
wire S15043;
wire S15044;
wire S15045;
wire S15046;
wire S15047;
wire S15048;
wire S15049;
wire S15050;
wire S15051;
wire S15052;
wire S15053;
wire S15054;
wire S15055;
wire S15056;
wire S15057;
wire S15058;
wire S15059;
wire S15060;
wire S15061;
wire S15062;
wire S15063;
wire S15064;
wire S15065;
wire S15066;
wire S15067;
wire S15068;
wire S15069;
wire S15070;
wire S15071;
wire S15072;
wire S15073;
wire S15074;
wire S15075;
wire S15076;
wire S15077;
wire S15078;
wire S15079;
wire S15080;
wire S15081;
wire S15082;
wire S15083;
wire S15084;
wire S15085;
wire S15086;
wire S15087;
wire S15088;
wire S15089;
wire S15090;
wire S15091;
wire S15092;
wire S15093;
wire S15094;
wire S15095;
wire S15096;
wire S15097;
wire S15098;
wire S15099;
wire S15100;
wire S15101;
wire S15102;
wire S15103;
wire S15104;
wire S15105;
wire S15106;
wire S15107;
wire S15108;
wire S15109;
wire S15110;
wire S15111;
wire S15112;
wire S15113;
wire S15114;
wire S15115;
wire S15116;
wire S15117;
wire S15118;
wire S15119;
wire S15120;
wire S15121;
wire S15122;
wire S15123;
wire S15124;
wire S15125;
wire S15126;
wire S15127;
wire S15128;
wire S15129;
wire S15130;
wire S15131;
wire S15132;
wire S15133;
wire S15134;
wire S15135;
wire S15136;
wire S15137;
wire S15138;
wire S15139;
wire S15140;
wire S15141;
wire S15142;
wire S15143;
wire S15144;
wire S15145;
wire S15146;
wire S15147;
wire S15148;
wire S15149;
wire S15150;
wire S15151;
wire S15152;
wire S15153;
wire S15154;
wire S15155;
wire S15156;
wire S15157;
wire S15158;
wire S15159;
wire S15160;
wire S15161;
wire S15162;
wire S15163;
wire S15164;
wire S15165;
wire S15166;
wire S15167;
wire S15168;
wire S15169;
wire S15170;
wire S15171;
wire S15172;
wire S15173;
wire S15174;
wire S15175;
wire S15176;
wire S15177;
wire S15178;
wire S15179;
wire S15180;
wire S15181;
wire S15182;
wire S15183;
wire S15184;
wire S15185;
wire S15186;
wire S15187;
wire S15188;
wire S15189;
wire S15190;
wire S15191;
wire S15192;
wire S15193;
wire S15194;
wire S15195;
wire S15196;
wire S15197;
wire S15198;
wire S15199;
wire S15200;
wire S15201;
wire S15202;
wire S15203;
wire S15204;
wire S15205;
wire S15206;
wire S15207;
wire S15208;
wire S15209;
wire S15210;
wire S15211;
wire S15212;
wire S15213;
wire S15214;
wire S15215;
wire S15216;
wire S15217;
wire S15218;
wire S15219;
wire S15220;
wire S15221;
wire S15222;
wire S15223;
wire S15224;
wire S15225;
wire S15226;
wire S15227;
wire S15228;
wire S15229;
wire S15230;
wire S15231;
wire S15232;
wire S15233;
wire S15234;
wire S15235;
wire S15236;
wire S15237;
wire S15238;
wire S15239;
wire S15240;
wire S15241;
wire S15242;
wire S15243;
wire S15244;
wire S15245;
wire S15246;
wire S15247;
wire S15248;
wire S15249;
wire S15250;
wire S15251;
wire S15252;
wire S15253;
wire S15254;
wire S15255;
wire S15256;
wire S15257;
wire S15258;
wire S15259;
wire S15260;
wire S15261;
wire S15262;
wire S15263;
wire S15264;
wire S15265;
wire S15266;
wire S15267;
wire S15268;
wire S15269;
wire S15270;
wire S15271;
wire S15272;
wire S15273;
wire S15274;
wire S15275;
wire S15276;
wire S15277;
wire S15278;
wire S15279;
wire S15280;
wire S15281;
wire S15282;
wire S15283;
wire S15284;
wire S15285;
wire S15286;
wire S15287;
wire S15288;
wire S15289;
wire S15290;
wire S15291;
wire S15292;
wire S15293;
wire S15294;
wire S15295;
wire S15296;
wire S15297;
wire S15298;
wire S15299;
wire S15300;
wire S15301;
wire S15302;
wire S15303;
wire S15304;
wire S15305;
wire S15306;
wire S15307;
wire S15308;
wire S15309;
wire S15310;
wire S15311;
wire S15312;
wire S15313;
wire S15314;
wire S15315;
wire S15316;
wire S15317;
wire S15318;
wire S15319;
wire S15320;
wire S15321;
wire S15322;
wire S15323;
wire S15324;
wire S15325;
wire S15326;
wire S15327;
wire S15328;
wire S15329;
wire S15330;
wire S15331;
wire S15332;
wire S15333;
wire S15334;
wire S15335;
wire S15336;
wire S15337;
wire S15338;
wire S15339;
wire S15340;
wire S15341;
wire S15342;
wire S15343;
wire S15344;
wire S15345;
wire S15346;
wire S15347;
wire S15348;
wire S15349;
wire S15350;
wire S15351;
wire S15352;
wire S15353;
wire S15354;
wire S15355;
wire S15356;
wire S15357;
wire S15358;
wire S15359;
wire S15360;
wire S15361;
wire S15362;
wire S15363;
wire S15364;
wire S15365;
wire S15366;
wire S15367;
wire S15368;
wire S15369;
wire S15370;
wire S15371;
wire S15372;
wire S15373;
wire S15374;
wire S15375;
wire S15376;
wire S15377;
wire S15378;
wire S15379;
wire S15380;
wire S15381;
wire S15382;
wire S15383;
wire S15384;
wire S15385;
wire S15386;
wire S15387;
wire S15388;
wire S15389;
wire S15390;
wire S15391;
wire S15392;
wire S15393;
wire S15394;
wire S15395;
wire S15396;
wire S15397;
wire S15398;
wire S15399;
wire S15400;
wire S15401;
wire S15402;
wire S15403;
wire S15404;
wire S15405;
wire S15406;
wire S15407;
wire S15408;
wire S15409;
wire S15410;
wire S15411;
wire S15412;
wire S15413;
wire S15414;
wire S15415;
wire S15416;
wire S15417;
wire S15418;
wire S15419;
wire S15420;
wire S15421;
wire S15422;
wire S15423;
wire S15424;
wire S15425;
wire S15426;
wire S15427;
wire S15428;
wire S15429;
wire S15430;
wire S15431;
wire S15432;
wire S15433;
wire S15434;
wire S15435;
wire S15436;
wire S15437;
wire S15438;
wire S15439;
wire S15440;
wire S15441;
wire S15442;
wire S15443;
wire S15444;
wire S15445;
wire S15446;
wire S15447;
wire S15448;
wire S15449;
wire S15450;
wire S15451;
wire S15452;
wire S15453;
wire S15454;
wire S15455;
wire S15456;
wire S15457;
wire S15458;
wire S15459;
wire S15460;
wire S15461;
wire S15462;
wire S15463;
wire S15464;
wire S15465;
wire S15466;
wire S15467;
wire S15468;
wire S15469;
wire S15470;
wire S15471;
wire S15472;
wire S15473;
wire S15474;
wire S15475;
wire S15476;
wire S15477;
wire S15478;
wire S15479;
wire S15480;
wire S15481;
wire S15482;
wire S15483;
wire S15484;
wire S15485;
wire S15486;
wire S15487;
wire S15488;
wire S15489;
wire S15490;
wire S15491;
wire S15492;
wire S15493;
wire S15494;
wire S15495;
wire S15496;
wire S15497;
wire S15498;
wire S15499;
wire S15500;
wire S15501;
wire S15502;
wire S15503;
wire S15504;
wire S15505;
wire S15506;
wire S15507;
wire S15508;
wire S15509;
wire S15510;
wire S15511;
wire S15512;
wire S15513;
wire S15514;
wire S15515;
wire S15516;
wire S15517;
wire S15518;
wire S15519;
wire S15520;
wire S15521;
wire S15522;
wire S15523;
wire S15524;
wire S15525;
wire S15526;
wire S15527;
wire S15528;
wire S15529;
wire S15530;
wire S15531;
wire S15532;
wire S15533;
wire S15534;
wire S15535;
wire S15536;
wire S15537;
wire S15538;
wire S15539;
wire S15540;
wire S15541;
wire S15542;
wire S15543;
wire S15544;
wire S15545;
wire S15546;
wire S15547;
wire S15548;
wire S15549;
wire S15550;
wire S15551;
wire S15552;
wire S15553;
wire S15554;
wire S15555;
wire S15556;
wire S15557;
wire S15558;
wire S15559;
wire S15560;
wire S15561;
wire S15562;
wire S15563;
wire S15564;
wire S15565;
wire S15566;
wire S15567;
wire S15568;
wire S15569;
wire S15570;
wire S15571;
wire S15572;
wire S15573;
wire S15574;
wire S15575;
wire S15576;
wire S15577;
wire S15578;
wire S15579;
wire S15580;
wire S15581;
wire S15582;
wire S15583;
wire S15584;
wire S15585;
wire S15586;
wire S15587;
wire S15588;
wire S15589;
wire S15590;
wire S15591;
wire S15592;
wire S15593;
wire S15594;
wire S15595;
wire S15596;
wire S15597;
wire S15598;
wire S15599;
wire S15600;
wire S15601;
wire S15602;
wire S15603;
wire S15604;
wire S15605;
wire S15606;
wire S15607;
wire S15608;
wire S15609;
wire S15610;
wire S15611;
wire S15612;
wire S15613;
wire S15614;
wire S15615;
wire S15616;
wire S15617;
wire S15618;
wire S15619;
wire S15620;
wire S15621;
wire S15622;
wire S15623;
wire S15624;
wire S15625;
wire S15626;
wire S15627;
wire S15628;
wire S15629;
wire S15630;
wire S15631;
wire S15632;
wire S15633;
wire S15634;
wire S15635;
wire S15636;
wire S15637;
wire S15638;
wire S15639;
wire S15640;
wire S15641;
wire S15642;
wire S15643;
wire S15644;
wire S15645;
wire S15646;
wire S15647;
wire S15648;
wire S15649;
wire S15650;
wire S15651;
wire S15652;
wire S15653;
wire S15654;
wire S15655;
wire S15656;
wire S15657;
wire S15658;
wire S15659;
wire S15660;
wire S15661;
wire S15662;
wire S15663;
wire S15664;
wire S15665;
wire S15666;
wire S15667;
wire S15668;
wire S15669;
wire S15670;
wire S15671;
wire S15672;
wire S15673;
wire S15674;
wire S15675;
wire S15676;
wire S15677;
wire S15678;
wire S15679;
wire S15680;
wire S15681;
wire S15682;
wire S15683;
wire S15684;
wire S15685;
wire S15686;
wire S15687;
wire S15688;
wire S15689;
wire S15690;
wire S15691;
wire S15692;
wire S15693;
wire S15694;
wire S15695;
wire S15696;
wire S15697;
wire S15698;
wire S15699;
wire S15700;
wire S15701;
wire S15702;
wire S15703;
wire S15704;
wire S15705;
wire S15706;
wire S15707;
wire S15708;
wire S15709;
wire S15710;
wire S15711;
wire S15712;
wire S15713;
wire S15714;
wire S15715;
wire S15716;
wire S15717;
wire S15718;
wire S15719;
wire S15720;
wire S15721;
wire S15722;
wire S15723;
wire S15724;
wire S15725;
wire S15726;
wire S15727;
wire S15728;
wire S15729;
wire S15730;
wire S15731;
wire S15732;
wire S15733;
wire S15734;
wire S15735;
wire S15736;
wire S15737;
wire S15738;
wire S15739;
wire S15740;
wire S15741;
wire S15742;
wire S15743;
wire S15744;
wire S15745;
wire S15746;
wire S15747;
wire S15748;
wire S15749;
wire S15750;
wire S15751;
wire S15752;
wire S15753;
wire S15754;
wire S15755;
wire S15756;
wire S15757;
wire S15758;
wire S15759;
wire S15760;
wire S15761;
wire S15762;
wire S15763;
wire S15764;
wire S15765;
wire S15766;
wire S15767;
wire S15768;
wire S15769;
wire S15770;
wire S15771;
wire S15772;
wire S15773;
wire S15774;
wire S15775;
wire S15776;
wire S15777;
wire S15778;
wire S15779;
wire S15780;
wire S15781;
wire S15782;
wire S15783;
wire S15784;
wire S15785;
wire S15786;
wire S15787;
wire S15788;
wire S15789;
wire S15790;
wire S15791;
wire S15792;
wire S15793;
wire S15794;
wire S15795;
wire S15796;
wire S15797;
wire S15798;
wire S15799;
wire S15800;
wire S15801;
wire S15802;
wire S15803;
wire S15804;
wire S15805;
wire S15806;
wire S15807;
wire S15808;
wire S15809;
wire S15810;
wire S15811;
wire S15812;
wire S15813;
wire S15814;
wire S15815;
wire S15816;
wire S15817;
wire S15818;
wire S15819;
wire S15820;
wire S15821;
wire S15822;
wire S15823;
wire S15824;
wire S15825;
wire S15826;
wire S15827;
wire S15828;
wire S15829;
wire S15830;
wire S15831;
wire S15832;
wire S15833;
wire S15834;
wire S15835;
wire S15836;
wire S15837;
wire S15838;
wire S15839;
wire S15840;
wire S15841;
wire S15842;
wire S15843;
wire S15844;
wire S15845;
wire S15846;
wire S15847;
wire S15848;
wire S15849;
wire S15850;
wire S15851;
wire S15852;
wire S15853;
wire S15854;
wire S15855;
wire S15856;
wire S15857;
wire S15858;
wire S15859;
wire S15860;
wire S15861;
wire S15862;
wire S15863;
wire S15864;
wire S15865;
wire S15866;
wire S15867;
wire S15868;
wire S15869;
wire S15870;
wire S15871;
wire S15872;
wire S15873;
wire S15874;
wire S15875;
wire S15876;
wire S15877;
wire S15878;
wire S15879;
wire S15880;
wire S15881;
wire S15882;
wire S15883;
wire S15884;
wire S15885;
wire S15886;
wire S15887;
wire S15888;
wire S15889;
wire S15890;
wire S15891;
wire S15892;
wire S15893;
wire S15894;
wire S15895;
wire S15896;
wire S15897;
wire S15898;
wire S15899;
wire S15900;
wire S15901;
wire S15902;
wire S15903;
wire S15904;
wire S15905;
wire S15906;
wire S15907;
wire S15908;
wire S15909;
wire S15910;
wire S15911;
wire S15912;
wire S15913;
wire S15914;
wire S15915;
wire S15916;
wire S15917;
wire S15918;
wire S15919;
wire S15920;
wire S15921;
wire S15922;
wire S15923;
wire S15924;
wire S15925;
wire S15926;
wire S15927;
wire S15928;
wire S15929;
wire S15930;
wire S15931;
wire S15932;
wire S15933;
wire S15934;
wire S15935;
wire S15936;
wire S15937;
wire S15938;
wire S15939;
wire S15940;
wire S15941;
wire S15942;
wire S15943;
wire S15944;
wire S15945;
wire S15946;
wire S15947;
wire S15948;
wire S15949;
wire S15950;
wire S15951;
wire S15952;
wire S15953;
wire S15954;
wire S15955;
wire S15956;
wire S15957;
wire S15958;
wire S15959;
wire S15960;
wire S15961;
wire S15962;
wire S15963;
wire S15964;
wire S15965;
wire S15966;
wire S15967;
wire S15968;
wire S15969;
wire S15970;
wire S15971;
wire S15972;
wire S15973;
wire S15974;
wire S15975;
wire S15976;
wire S15977;
wire S15978;
wire S15979;
wire S15980;
wire S15981;
wire S15982;
wire S15983;
wire S15984;
wire S15985;
wire S15986;
wire S15987;
wire S15988;
wire S15989;
wire S15990;
wire S15991;
wire S15992;
wire S15993;
wire S15994;
wire S15995;
wire S15996;
wire S15997;
wire S15998;
wire S15999;
wire S16000;
wire S16001;
wire S16002;
wire S16003;
wire S16004;
wire S16005;
wire S16006;
wire S16007;
wire S16008;
wire S16009;
wire S16010;
wire S16011;
wire S16012;
wire S16013;
wire S16014;
wire S16015;
wire S16016;
wire S16017;
wire S16018;
wire S16019;
wire S16020;
wire S16021;
wire S16022;
wire S16023;
wire S16024;
wire S16025;
wire S16026;
wire S16027;
wire S16028;
wire S16029;
wire S16030;
wire S16031;
wire S16032;
wire S16033;
wire S16034;
wire S16035;
wire S16036;
wire S16037;
wire S16038;
wire S16039;
wire S16040;
wire S16041;
wire S16042;
wire S16043;
wire S16044;
wire S16045;
wire S16046;
wire S16047;
wire S16048;
wire S16049;
wire S16050;
wire S16051;
wire S16052;
wire S16053;
wire S16054;
wire S16055;
wire S16056;
wire S16057;
wire S16058;
wire S16059;
wire S16060;
wire S16061;
wire S16062;
wire S16063;
wire S16064;
wire S16065;
wire S16066;
wire S16067;
wire S16068;
wire S16069;
wire S16070;
wire S16071;
wire S16072;
wire S16073;
wire S16074;
wire S16075;
wire S16076;
wire S16077;
wire S16078;
wire S16079;
wire S16080;
wire S16081;
wire S16082;
wire S16083;
wire S16084;
wire S16085;
wire S16086;
wire S16087;
wire S16088;
wire S16089;
wire S16090;
wire S16091;
wire S16092;
wire S16093;
wire S16094;
wire S16095;
wire S16096;
wire S16097;
wire S16098;
wire S16099;
wire S16100;
wire S16101;
wire S16102;
wire S16103;
wire S16104;
wire S16105;
wire S16106;
wire S16107;
wire S16108;
wire S16109;
wire S16110;
wire S16111;
wire S16112;
wire S16113;
wire S16114;
wire S16115;
wire S16116;
wire S16117;
wire S16118;
wire S16119;
wire S16120;
wire S16121;
wire S16122;
wire S16123;
wire S16124;
wire S16125;
wire S16126;
wire S16127;
wire S16128;
wire S16129;
wire S16130;
wire S16131;
wire S16132;
wire S16133;
wire S16134;
wire S16135;
wire S16136;
wire S16137;
wire S16138;
wire S16139;
wire S16140;
wire S16141;
wire S16142;
wire S16143;
wire S16144;
wire S16145;
wire S16146;
wire S16147;
wire S16148;
wire S16149;
wire S16150;
wire S16151;
wire S16152;
wire S16153;
wire S16154;
wire S16155;
wire S16156;
wire S16157;
wire S16158;
wire S16159;
wire S16160;
wire S16161;
wire S16162;
wire S16163;
wire S16164;
wire S16165;
wire S16166;
wire S16167;
wire S16168;
wire S16169;
wire S16170;
wire S16171;
wire S16172;
wire S16173;
wire S16174;
wire S16175;
wire S16176;
wire S16177;
wire S16178;
wire S16179;
wire S16180;
wire S16181;
wire S16182;
wire S16183;
wire S16184;
wire S16185;
wire S16186;
wire S16187;
wire S16188;
wire S16189;
wire S16190;
wire S16191;
wire S16192;
wire S16193;
wire S16194;
wire S16195;
wire S16196;
wire S16197;
wire S16198;
wire S16199;
wire S16200;
wire S16201;
wire S16202;
wire S16203;
wire S16204;
wire S16205;
wire S16206;
wire S16207;
wire S16208;
wire S16209;
wire S16210;
wire S16211;
wire S16212;
wire S16213;
wire S16214;
wire S16215;
wire S16216;
wire S16217;
wire S16218;
wire S16219;
wire S16220;
wire S16221;
wire S16222;
wire S16223;
wire S16224;
wire S16225;
wire S16226;
wire S16227;
wire S16228;
wire S16229;
wire S16230;
wire S16231;
wire S16232;
wire S16233;
wire S16234;
wire S16235;
wire S16236;
wire S16237;
wire S16238;
wire S16239;
wire S16240;
wire S16241;
wire S16242;
wire S16243;
wire S16244;
wire S16245;
wire S16246;
wire S16247;
wire S16248;
wire S16249;
wire S16250;
wire S16251;
wire S16252;
wire S16253;
wire S16254;
wire S16255;
wire S16256;
wire S16257;
wire S16258;
wire S16259;
wire S16260;
wire S16261;
wire S16262;
wire S16263;
wire S16264;
wire S16265;
wire S16266;
wire S16267;
wire S16268;
wire S16269;
wire S16270;
wire S16271;
wire S16272;
wire S16273;
wire S16274;
wire S16275;
wire S16276;
wire S16277;
wire S16278;
wire S16279;
wire S16280;
wire S16281;
wire S16282;
wire S16283;
wire S16284;
wire S16285;
wire S16286;
wire S16287;
wire S16288;
wire S16289;
wire S16290;
wire S16291;
wire S16292;
wire S16293;
wire S16294;
wire S16295;
wire S16296;
wire S16297;
wire S16298;
wire S16299;
wire S16300;
wire S16301;
wire S16302;
wire S16303;
wire S16304;
wire S16305;
wire S16306;
wire S16307;
wire S16308;
wire S16309;
wire S16310;
wire S16311;
wire S16312;
wire S16313;
wire S16314;
wire S16315;
wire S16316;
wire S16317;
wire S16318;
wire S16319;
wire S16320;
wire S16321;
wire S16322;
wire S16323;
wire S16324;
wire S16325;
wire S16326;
wire S16327;
wire S16328;
wire S16329;
wire S16330;
wire S16331;
wire S16332;
wire S16333;
wire S16334;
wire S16335;
wire S16336;
wire S16337;
wire S16338;
wire S16339;
wire S16340;
wire S16341;
wire S16342;
wire S16343;
wire S16344;
wire S16345;
wire S16346;
wire S16347;
wire S16348;
wire S16349;
wire S16350;
wire S16351;
wire S16352;
wire S16353;
wire S16354;
wire S16355;
wire S16356;
wire S16357;
wire S16358;
wire S16359;
wire S16360;
wire S16361;
wire S16362;
wire S16363;
wire S16364;
wire S16365;
wire S16366;
wire S16367;
wire S16368;
wire S16369;
wire S16370;
wire S16371;
wire S16372;
wire S16373;
wire S16374;
wire S16375;
wire S16376;
wire S16377;
wire S16378;
wire S16379;
wire S16380;
wire S16381;
wire S16382;
wire S16383;
wire S16384;
wire S16385;
wire S16386;
wire S16387;
wire S16388;
wire S16389;
wire S16390;
wire S16391;
wire S16392;
wire S16393;
wire S16394;
wire S16395;
wire S16396;
wire S16397;
wire S16398;
wire S16399;
wire S16400;
wire S16401;
wire S16402;
wire S16403;
wire S16404;
wire S16405;
wire S16406;
wire S16407;
wire S16408;
wire S16409;
wire S16410;
wire S16411;
wire S16412;
wire S16413;
wire S16414;
wire S16415;
wire S16416;
wire S16417;
wire S16418;
wire S16419;
wire S16420;
wire S16421;
wire S16422;
wire S16423;
wire S16424;
wire S16425;
wire S16426;
wire S16427;
wire S16428;
wire S16429;
wire S16430;
wire S16431;
wire S16432;
wire S16433;
wire S16434;
wire S16435;
wire S16436;
wire S16437;
wire S16438;
wire S16439;
wire S16440;
wire S16441;
wire S16442;
wire S16443;
wire S16444;
wire S16445;
wire S16446;
wire S16447;
wire S16448;
wire S16449;
wire S16450;
wire S16451;
wire S16452;
wire S16453;
wire S16454;
wire S16455;
wire S16456;
wire S16457;
wire S16458;
wire S16459;
wire S16460;
wire S16461;
wire S16462;
wire S16463;
wire S16464;
wire S16465;
wire S16466;
wire S16467;
wire S16468;
wire S16469;
wire S16470;
wire S16471;
wire S16472;
wire S16473;
wire S16474;
wire S16475;
wire S16476;
wire S16477;
wire S16478;
wire S16479;
wire S16480;
wire S16481;
wire S16482;
wire S16483;
wire S16484;
wire S16485;
wire S16486;
wire S16487;
wire S16488;
wire S16489;
wire S16490;
wire S16491;
wire S16492;
wire S16493;
wire S16494;
wire S16495;
wire S16496;
wire S16497;
wire S16498;
wire S16499;
wire S16500;
wire S16501;
wire S16502;
wire S16503;
wire S16504;
wire S16505;
wire S16506;
wire S16507;
wire S16508;
wire S16509;
wire S16510;
wire S16511;
wire S16512;
wire S16513;
wire S16514;
wire S16515;
wire S16516;
wire S16517;
wire S16518;
wire S16519;
wire S16520;
wire S16521;
wire S16522;
wire S16523;
wire S16524;
wire S16525;
wire S16526;
wire S16527;
wire S16528;
wire S16529;
wire S16530;
wire S16531;
wire S16532;
wire S16533;
wire S16534;
wire S16535;
wire S16536;
wire S16537;
wire S16538;
wire S16539;
wire S16540;
wire S16541;
wire S16542;
wire S16543;
wire S16544;
wire S16545;
wire S16546;
wire S16547;
wire S16548;
wire S16549;
wire S16550;
wire S16551;
wire S16552;
wire S16553;
wire S16554;
wire S16555;
wire S16556;
wire S16557;
wire S16558;
wire S16559;
wire S16560;
wire S16561;
wire S16562;
wire S16563;
wire S16564;
wire S16565;
wire S16566;
wire S16567;
wire S16568;
wire S16569;
wire S16570;
wire S16571;
wire S16572;
wire S16573;
wire S16574;
wire S16575;
wire S16576;
wire S16577;
wire S16578;
wire S16579;
wire S16580;
wire S16581;
wire S16582;
wire S16583;
wire S16584;
wire S16585;
wire S16586;
wire S16587;
wire S16588;
wire S16589;
wire S16590;
wire S16591;
wire S16592;
wire S16593;
wire S16594;
wire S16595;
wire S16596;
wire S16597;
wire S16598;
wire S16599;
wire S16600;
wire S16601;
wire S16602;
wire S16603;
wire S16604;
wire S16605;
wire S16606;
wire S16607;
wire S16608;
wire S16609;
wire S16610;
wire S16611;
wire S16612;
wire S16613;
wire S16614;
wire S16615;
wire S16616;
wire S16617;
wire S16618;
wire S16619;
wire S16620;
wire S16621;
wire S16622;
wire S16623;
wire S16624;
wire S16625;
wire S16626;
wire S16627;
wire S16628;
wire S16629;
wire S16630;
wire S16631;
wire S16632;
wire S16633;
wire S16634;
wire S16635;
wire S16636;
wire S16637;
wire S16638;
wire S16639;
wire S16640;
wire S16641;
wire S16642;
wire S16643;
wire S16644;
wire S16645;
wire S16646;
wire S16647;
wire S16648;
wire S16649;
wire S16650;
wire S16651;
wire S16652;
wire S16653;
wire S16654;
wire S16655;
wire S16656;
wire S16657;
wire S16658;
wire S16659;
wire S16660;
wire S16661;
wire S16662;
wire S16663;
wire S16664;
wire S16665;
wire S16666;
wire S16667;
wire S16668;
wire S16669;
wire S16670;
wire S16671;
wire S16672;
wire S16673;
wire S16674;
wire S16675;
wire S16676;
wire S16677;
wire S16678;
wire S16679;
wire S16680;
wire S16681;
wire S16682;
wire S16683;
wire S16684;
wire S16685;
wire S16686;
wire S16687;
wire S16688;
wire S16689;
wire S16690;
wire S16691;
wire S16692;
wire S16693;
wire S16694;
wire S16695;
wire S16696;
wire S16697;
wire S16698;
wire S16699;
wire S16700;
wire S16701;
wire S16702;
wire S16703;
wire S16704;
wire S16705;
wire S16706;
wire S16707;
wire S16708;
wire S16709;
wire S16710;
wire S16711;
wire S16712;
wire S16713;
wire S16714;
wire S16715;
wire S16716;
wire S16717;
wire S16718;
wire S16719;
wire S16720;
wire S16721;
wire S16722;
wire S16723;
wire S16724;
wire S16725;
wire S16726;
wire S16727;
wire S16728;
wire S16729;
wire S16730;
wire S16731;
wire S16732;
wire S16733;
wire S16734;
wire S16735;
wire S16736;
wire S16737;
wire S16738;
wire S16739;
wire S16740;
wire S16741;
wire S16742;
wire S16743;
wire S16744;
wire S16745;
wire S16746;
wire S16747;
wire S16748;
wire S16749;
wire S16750;
wire S16751;
wire S16752;
wire S16753;
wire S16754;
wire S16755;
wire S16756;
wire S16757;
wire S16758;
wire S16759;
wire S16760;
wire S16761;
wire S16762;
wire S16763;
wire S16764;
wire S16765;
wire S16766;
wire S16767;
wire S16768;
wire S16769;
wire S16770;
wire S16771;
wire S16772;
wire S16773;
wire S16774;
wire S16775;
wire S16776;
wire S16777;
wire S16778;
wire S16779;
wire S16780;
wire S16781;
wire S16782;
wire S16783;
wire S16784;
wire S16785;
wire S16786;
wire S16787;
wire S16788;
wire S16789;
wire S16790;
wire S16791;
wire S16792;
wire S16793;
wire S16794;
wire S16795;
wire S16796;
wire S16797;
wire S16798;
wire S16799;
wire S16800;
wire S16801;
wire S16802;
wire S16803;
wire S16804;
wire S16805;
wire S16806;
wire S16807;
wire S16808;
wire S16809;
wire S16810;
wire S16811;
wire S16812;
wire S16813;
wire S16814;
wire S16815;
wire S16816;
wire S16817;
wire S16818;
wire S16819;
wire S16820;
wire S16821;
wire S16822;
wire S16823;
wire S16824;
wire S16825;
wire S16826;
wire S16827;
wire S16828;
wire S16829;
wire S16830;
wire S16831;
wire S16832;
wire S16833;
wire S16834;
wire S16835;
wire S16836;
wire S16837;
wire S16838;
wire S16839;
wire S16840;
wire S16841;
wire S16842;
wire S16843;
wire S16844;
wire S16845;
wire S16846;
wire S16847;
wire S16848;
wire S16849;
wire S16850;
wire S16851;
wire S16852;
wire S16853;
wire S16854;
wire S16855;
wire S16856;
wire S16857;
wire S16858;
wire S16859;
wire S16860;
wire S16861;
wire S16862;
wire S16863;
wire S16864;
wire S16865;
wire S16866;
wire S16867;
wire S16868;
wire S16869;
wire S16870;
wire S16871;
wire S16872;
wire S16873;
wire S16874;
wire S16875;
wire S16876;
wire S16877;
wire S16878;
wire S16879;
wire S16880;
wire S16881;
wire S16882;
wire S16883;
wire S16884;
wire S16885;
wire S16886;
wire S16887;
wire S16888;
wire S16889;
wire S16890;
wire S16891;
wire S16892;
wire S16893;
wire S16894;
wire S16895;
wire S16896;
wire S16897;
wire S16898;
wire S16899;
wire S16900;
wire S16901;
wire S16902;
wire S16903;
wire S16904;
wire S16905;
wire S16906;
wire S16907;
wire S16908;
wire S16909;
wire S16910;
wire S16911;
wire S16912;
wire S16913;
wire S16914;
wire S16915;
wire S16916;
wire S16917;
wire S16918;
wire S16919;
wire S16920;
wire S16921;
wire S16922;
wire S16923;
wire S16924;
wire S16925;
wire S16926;
wire S16927;
wire S16928;
wire S16929;
wire S16930;
wire S16931;
wire S16932;
wire S16933;
wire S16934;
wire S16935;
wire S16936;
wire S16937;
wire S16938;
wire S16939;
wire S16940;
wire S16941;
wire S16942;
wire S16943;
wire S16944;
wire S16945;
wire S16946;
wire S16947;
wire S16948;
wire S16949;
wire S16950;
wire S16951;
wire S16952;
wire S16953;
wire S16954;
wire S16955;
wire S16956;
wire S16957;
wire S16958;
wire S16959;
wire S16960;
wire S16961;
wire S16962;
wire S16963;
wire S16964;
wire S16965;
wire S16966;
wire S16967;
wire S16968;
wire S16969;
wire S16970;
wire S16971;
wire S16972;
wire S16973;
wire S16974;
wire S16975;
wire S16976;
wire S16977;
wire S16978;
wire S16979;
wire S16980;
wire S16981;
wire S16982;
wire S16983;
wire S16984;
wire S16985;
wire S16986;
wire S16987;
wire S16988;
wire S16989;
wire S16990;
wire S16991;
wire S16992;
wire S16993;
wire S16994;
wire S16995;
wire S16996;
wire S16997;
wire S16998;
wire S16999;
wire S17000;
wire S17001;
wire S17002;
wire S17003;
wire S17004;
wire S17005;
wire S17006;
wire S17007;
wire S17008;
wire S17009;
wire S17010;
wire S17011;
wire S17012;
wire S17013;
wire S17014;
wire S17015;
wire S17016;
wire S17017;
wire S17018;
wire S17019;
wire S17020;
wire S17021;
wire S17022;
wire S17023;
wire S17024;
wire S17025;
wire S17026;
wire S17027;
wire S17028;
wire S17029;
wire S17030;
wire S17031;
wire S17032;
wire S17033;
wire S17034;
wire S17035;
wire S17036;
wire S17037;
wire S17038;
wire S17039;
wire S17040;
wire S17041;
wire S17042;
wire S17043;
wire S17044;
wire S17045;
wire S17046;
wire S17047;
wire S17048;
wire S17049;
wire S17050;
wire S17051;
wire S17052;
wire S17053;
wire S17054;
wire S17055;
wire S17056;
wire S17057;
wire S17058;
wire S17059;
wire S17060;
wire S17061;
wire S17062;
wire S17063;
wire S17064;
wire S17065;
wire S17066;
wire S17067;
wire S17068;
wire S17069;
wire S17070;
wire S17071;
wire S17072;
wire S17073;
wire S17074;
wire S17075;
wire S17076;
wire S17077;
wire S17078;
wire S17079;
wire S17080;
wire S17081;
wire S17082;
wire S17083;
wire S17084;
wire S17085;
wire S17086;
wire S17087;
wire S17088;
wire S17089;
wire S17090;
wire S17091;
wire S17092;
wire S17093;
wire S17094;
wire S17095;
wire S17096;
wire S17097;
wire S17098;
wire S17099;
wire S17100;
wire S17101;
wire S17102;
wire S17103;
wire S17104;
wire S17105;
wire S17106;
wire S17107;
wire S17108;
wire S17109;
wire S17110;
wire S17111;
wire S17112;
wire S17113;
wire S17114;
wire S17115;
wire S17116;
wire S17117;
wire S17118;
wire S17119;
wire S17120;
wire S17121;
wire S17122;
wire S17123;
wire S17124;
wire S17125;
wire S17126;
wire S17127;
wire S17128;
wire S17129;
wire S17130;
wire S17131;
wire S17132;
wire S17133;
wire S17134;
wire S17135;
wire S17136;
wire S17137;
wire S17138;
wire S17139;
wire S17140;
wire S17141;
wire S17142;
wire S17143;
wire S17144;
wire S17145;
wire S17146;
wire S17147;
wire S17148;
wire S17149;
wire S17150;
wire S17151;
wire S17152;
wire S17153;
wire S17154;
wire S17155;
wire S17156;
wire S17157;
wire S17158;
wire S17159;
wire S17160;
wire S17161;
wire S17162;
wire S17163;
wire S17164;
wire S17165;
wire S17166;
wire S17167;
wire S17168;
wire S17169;
wire S17170;
wire S17171;
wire S17172;
wire S17173;
wire S17174;
wire S17175;
wire S17176;
wire S17177;
wire S17178;
wire S17179;
wire S17180;
wire S17181;
wire S17182;
wire S17183;
wire S17184;
wire S17185;
wire S17186;
wire S17187;
wire S17188;
wire S17189;
wire S17190;
wire S17191;
wire S17192;
wire S17193;
wire S17194;
wire S17195;
wire S17196;
wire S17197;
wire S17198;
wire S17199;
wire S17200;
wire S17201;
wire S17202;
wire S17203;
wire S17204;
wire S17205;
wire S17206;
wire S17207;
wire S17208;
wire S17209;
wire S17210;
wire S17211;
wire S17212;
wire S17213;
wire S17214;
wire S17215;
wire S17216;
wire S17217;
wire S17218;
wire S17219;
wire S17220;
wire S17221;
wire S17222;
wire S17223;
wire S17224;
wire S17225;
wire S17226;
wire S17227;
wire S17228;
wire S17229;
wire S17230;
wire S17231;
wire S17232;
wire S17233;
wire S17234;
wire S17235;
wire S17236;
wire S17237;
wire S17238;
wire S17239;
wire S17240;
wire S17241;
wire S17242;
wire S17243;
wire S17244;
wire S17245;
wire S17246;
wire S17247;
wire S17248;
wire S17249;
wire S17250;
wire S17251;
wire S17252;
wire S17253;
wire S17254;
wire S17255;
wire S17256;
wire S17257;
wire S17258;
wire S17259;
wire S17260;
wire S17261;
wire S17262;
wire S17263;
wire S17264;
wire S17265;
wire S17266;
wire S17267;
wire S17268;
wire S17269;
wire S17270;
wire S17271;
wire S17272;
wire S17273;
wire S17274;
wire S17275;
wire S17276;
wire S17277;
wire S17278;
wire S17279;
wire S17280;
wire S17281;
wire S17282;
wire S17283;
wire S17284;
wire S17285;
wire S17286;
wire S17287;
wire S17288;
wire S17289;
wire S17290;
wire S17291;
wire S17292;
wire S17293;
wire S17294;
wire S17295;
wire S17296;
wire S17297;
wire S17298;
wire S17299;
wire S17300;
wire S17301;
wire S17302;
wire S17303;
wire S17304;
wire S17305;
wire S17306;
wire S17307;
wire S17308;
wire S17309;
wire S17310;
wire S17311;
wire S17312;
wire S17313;
wire S17314;
wire S17315;
wire S17316;
wire S17317;
wire S17318;
wire S17319;
wire S17320;
wire S17321;
wire S17322;
wire S17323;
wire S17324;
wire S17325;
wire S17326;
wire S17327;
wire S17328;
wire S17329;
wire S17330;
wire S17331;
wire S17332;
wire S17333;
wire S17334;
wire S17335;
wire S17336;
wire S17337;
wire S17338;
wire S17339;
wire S17340;
wire S17341;
wire S17342;
wire S17343;
wire S17344;
wire S17345;
wire S17346;
wire S17347;
wire S17348;
wire S17349;
wire S17350;
wire S17351;
wire S17352;
wire S17353;
wire S17354;
wire S17355;
wire S17356;
wire S17357;
wire S17358;
wire S17359;
wire S17360;
wire S17361;
wire S17362;
wire S17363;
wire S17364;
wire S17365;
wire S17366;
wire S17367;
wire S17368;
wire S17369;
wire S17370;
wire S17371;
wire S17372;
wire S17373;
wire S17374;
wire S17375;
wire S17376;
wire S17377;
wire S17378;
wire S17379;
wire S17380;
wire S17381;
wire S17382;
wire S17383;
wire S17384;
wire S17385;
wire S17386;
wire S17387;
wire S17388;
wire S17389;
wire S17390;
wire S17391;
wire S17392;
wire S17393;
wire S17394;
wire S17395;
wire S17396;
wire S17397;
wire S17398;
wire S17399;
wire S17400;
wire S17401;
wire S17402;
wire S17403;
wire S17404;
wire S17405;
wire S17406;
wire S17407;
wire S17408;
wire S17409;
wire S17410;
wire S17411;
wire S17412;
wire S17413;
wire S17414;
wire S17415;
wire S17416;
wire S17417;
wire S17418;
wire S17419;
wire S17420;
wire S17421;
wire S17422;
wire S17423;
wire S17424;
wire S17425;
wire S17426;
wire S17427;
wire S17428;
wire S17429;
wire S17430;
wire S17431;
wire S17432;
wire S17433;
wire S17434;
wire S17435;
wire S17436;
wire S17437;
wire S17438;
wire S17439;
wire S17440;
wire S17441;
wire S17442;
wire S17443;
wire S17444;
wire S17445;
wire S17446;
wire S17447;
wire S17448;
wire S17449;
wire S17450;
wire S17451;
wire S17452;
wire S17453;
wire S17454;
wire S17455;
wire S17456;
wire S17457;
wire S17458;
wire S17459;
wire S17460;
wire S17461;
wire S17462;
wire S17463;
wire S17464;
wire S17465;
wire S17466;
wire S17467;
wire S17468;
wire S17469;
wire S17470;
wire S17471;
wire S17472;
wire S17473;
wire S17474;
wire S17475;
wire S17476;
wire S17477;
wire S17478;
wire S17479;
wire S17480;
wire S17481;
wire S17482;
wire S17483;
wire S17484;
wire S17485;
wire S17486;
wire S17487;
wire S17488;
wire S17489;
wire S17490;
wire S17491;
wire S17492;
wire S17493;
wire S17494;
wire S17495;
wire S17496;
wire S17497;
wire S17498;
wire S17499;
wire S17500;
wire S17501;
wire S17502;
wire S17503;
wire S17504;
wire S17505;
wire S17506;
wire S17507;
wire S17508;
wire S17509;
wire S17510;
wire S17511;
wire S17512;
wire S17513;
wire S17514;
wire S17515;
wire S17516;
wire S17517;
wire S17518;
wire S17519;
wire S17520;
wire S17521;
wire S17522;
wire S17523;
wire S17524;
wire S17525;
wire S17526;
wire S17527;
wire S17528;
wire S17529;
wire S17530;
wire S17531;
wire S17532;
wire S17533;
wire S17534;
wire S17535;
wire S17536;
wire S17537;
wire S17538;
wire S17539;
wire S17540;
wire S17541;
wire S17542;
wire S17543;
wire S17544;
wire S17545;
wire S17546;
wire S17547;
wire S17548;
wire S17549;
wire S17550;
wire S17551;
wire S17552;
wire S17553;
wire S17554;
wire S17555;
wire S17556;
wire S17557;
wire S17558;
wire S17559;
wire S17560;
wire S17561;
wire S17562;
wire S17563;
wire S17564;
wire S17565;
wire S17566;
wire S17567;
wire S17568;
wire S17569;
wire S17570;
wire S17571;
wire S17572;
wire S17573;
wire S17574;
wire S17575;
wire S17576;
wire S17577;
wire S17578;
wire S17579;
wire S17580;
wire S17581;
wire S17582;
wire S17583;
wire S17584;
wire S17585;
wire S17586;
wire S17587;
wire S17588;
wire S17589;
wire S17590;
wire S17591;
wire S17592;
wire S17593;
wire S17594;
wire S17595;
wire S17596;
wire S17597;
wire S17598;
wire S17599;
wire S17600;
wire S17601;
wire S17602;
wire S17603;
wire S17604;
wire S17605;
wire S17606;
wire S17607;
wire S17608;
wire S17609;
wire S17610;
wire S17611;
wire S17612;
wire S17613;
wire S17614;
wire S17615;
wire S17616;
wire S17617;
wire S17618;
wire S17619;
wire S17620;
wire S17621;
wire S17622;
wire S17623;
wire S17624;
wire S17625;
wire S17626;
wire S17627;
wire S17628;
wire S17629;
wire S17630;
wire S17631;
wire S17632;
wire S17633;
wire S17634;
wire S17635;
wire S17636;
wire S17637;
wire S17638;
wire S17639;
wire S17640;
wire S17641;
wire S17642;
wire S17643;
wire S17644;
wire S17645;
wire S17646;
wire S17647;
wire S17648;
wire S17649;
wire S17650;
wire S17651;
wire S17652;
wire S17653;
wire S17654;
wire S17655;
wire S17656;
wire S17657;
wire S17658;
wire S17659;
wire S17660;
wire S17661;
wire S17662;
wire S17663;
wire S17664;
wire S17665;
wire S17666;
wire S17667;
wire S17668;
wire S17669;
wire S17670;
wire S17671;
wire S17672;
wire S17673;
wire S17674;
wire S17675;
wire S17676;
wire S17677;
wire S17678;
wire S17679;
wire S17680;
wire S17681;
wire S17682;
wire S17683;
wire S17684;
wire S17685;
wire S17686;
wire S17687;
wire S17688;
wire S17689;
wire S17690;
wire S17691;
wire S17692;
wire S17693;
wire S17694;
wire S17695;
wire S17696;
wire S17697;
wire S17698;
wire S17699;
wire S17700;
wire S17701;
wire S17702;
wire S17703;
wire S17704;
wire S17705;
wire S17706;
wire S17707;
wire S17708;
wire S17709;
wire S17710;
wire S17711;
wire S17712;
wire S17713;
wire S17714;
wire S17715;
wire S17716;
wire S17717;
wire S17718;
wire S17719;
wire S17720;
wire S17721;
wire S17722;
wire S17723;
wire S17724;
wire S17725;
wire S17726;
wire S17727;
wire S17728;
wire S17729;
wire S17730;
wire S17731;
wire S17732;
wire S17733;
wire S17734;
wire S17735;
wire S17736;
wire S17737;
wire S17738;
wire S17739;
wire S17740;
wire S17741;
wire S17742;
wire S17743;
wire S17744;
wire S17745;
wire S17746;
wire S17747;
wire S17748;
wire S17749;
wire S17750;
wire S17751;
wire S17752;
wire S17753;
wire S17754;
wire S17755;
wire S17756;
wire S17757;
wire S17758;
wire S17759;
wire S17760;
wire S17761;
wire S17762;
wire S17763;
wire S17764;
wire S17765;
wire S17766;
wire S17767;
wire S17768;
wire S17769;
wire S17770;
wire S17771;
wire S17772;
wire S17773;
wire S17774;
wire S17775;
wire S17776;
wire S17777;
wire S17778;
wire S17779;
wire S17780;
wire S17781;
wire S17782;
wire S17783;
wire S17784;
wire S17785;
wire S17786;
wire S17787;
wire S17788;
wire S17789;
wire S17790;
wire S17791;
wire S17792;
wire S17793;
wire S17794;
wire S17795;
wire S17796;
wire S17797;
wire S17798;
wire S17799;
wire S17800;
wire S17801;
wire S17802;
wire S17803;
wire S17804;
wire S17805;
wire S17806;
wire S17807;
wire S17808;
wire S17809;
wire S17810;
wire S17811;
wire S17812;
wire S17813;
wire S17814;
wire S17815;
wire S17816;
wire S17817;
wire S17818;
wire S17819;
wire S17820;
wire S17821;
wire S17822;
wire S17823;
wire S17824;
wire S17825;
wire S17826;
wire S17827;
wire S17828;
wire S17829;
wire S17830;
wire S17831;
wire S17832;
wire S17833;
wire S17834;
wire S17835;
wire S17836;
wire S17837;
wire S17838;
wire S17839;
wire S17840;
wire S17841;
wire S17842;
wire S17843;
wire S17844;
wire S17845;
wire S17846;
wire S17847;
wire S17848;
wire S17849;
wire S17850;
wire S17851;
wire S17852;
wire S17853;
wire S17854;
wire S17855;
wire S17856;
wire S17857;
wire S17858;
wire S17859;
wire S17860;
wire S17861;
wire S17862;
wire S17863;
wire S17864;
wire S17865;
wire S17866;
wire S17867;
wire S17868;
wire S17869;
wire S17870;
wire S17871;
wire S17872;
wire S17873;
wire S17874;
wire S17875;
wire S17876;
wire S17877;
wire S17878;
wire S17879;
wire S17880;
wire S17881;
wire S17882;
wire S17883;
wire S17884;
wire S17885;
wire S17886;
wire S17887;
wire S17888;
wire S17889;
wire S17890;
wire S17891;
wire S17892;
wire S17893;
wire S17894;
wire S17895;
wire S17896;
wire S17897;
wire S17898;
wire S17899;
wire S17900;
wire S17901;
wire S17902;
wire S17903;
wire S17904;
wire S17905;
wire S17906;
wire S17907;
wire S17908;
wire S17909;
wire S17910;
wire S17911;
wire S17912;
wire S17913;
wire S17914;
wire S17915;
wire S17916;
wire S17917;
wire S17918;
wire S17919;
wire S17920;
wire S17921;
wire S17922;
wire S17923;
wire S17924;
wire S17925;
wire S17926;
wire S17927;
wire S17928;
wire S17929;
wire S17930;
wire S17931;
wire S17932;
wire S17933;
wire S17934;
wire S17935;
wire S17936;
wire S17937;
wire S17938;
wire S17939;
wire S17940;
wire S17941;
wire S17942;
wire S17943;
wire S17944;
wire S17945;
wire S17946;
wire S17947;
wire S17948;
wire S17949;
wire S17950;
wire S17951;
wire S17952;
wire S17953;
wire S17954;
wire S17955;
wire S17956;
wire S17957;
wire S17958;
wire S17959;
wire S17960;
wire S17961;
wire S17962;
wire S17963;
wire S17964;
wire S17965;
wire S17966;
wire S17967;
wire S17968;
wire S17969;
wire S17970;
wire S17971;
wire S17972;
wire S17973;
wire S17974;
wire S17975;
wire S17976;
wire S17977;
wire S17978;
wire S17979;
wire S17980;
wire S17981;
wire S17982;
wire S17983;
wire S17984;
wire S17985;
wire S17986;
wire S17987;
wire S17988;
wire S17989;
wire S17990;
wire S17991;
wire S17992;
wire S17993;
wire S17994;
wire S17995;
wire S17996;
wire S17997;
wire S17998;
wire S17999;
wire S18000;
wire S18001;
wire S18002;
wire S18003;
wire S18004;
wire S18005;
wire S18006;
wire S18007;
wire S18008;
wire S18009;
wire S18010;
wire S18011;
wire S18012;
wire S18013;
wire S18014;
wire S18015;
wire S18016;
wire S18017;
wire S18018;
wire S18019;
wire S18020;
wire S18021;
wire S18022;
wire S18023;
wire S18024;
wire S18025;
wire S18026;
wire S18027;
wire S18028;
wire S18029;
wire S18030;
wire S18031;
wire S18032;
wire S18033;
wire S18034;
wire S18035;
wire S18036;
wire S18037;
wire S18038;
wire S18039;
wire S18040;
wire S18041;
wire S18042;
wire S18043;
wire S18044;
wire S18045;
wire S18046;
wire S18047;
wire S18048;
wire S18049;
wire S18050;
wire S18051;
wire S18052;
wire S18053;
wire S18054;
wire S18055;
wire S18056;
wire S18057;
wire S18058;
wire S18059;
wire S18060;
wire S18061;
wire S18062;
wire S18063;
wire S18064;
wire S18065;
wire S18066;
wire S18067;
wire S18068;
wire S18069;
wire S18070;
wire S18071;
wire S18072;
wire S18073;
wire S18074;
wire S18075;
wire S18076;
wire S18077;
wire S18078;
wire S18079;
wire S18080;
wire S18081;
wire S18082;
wire S18083;
wire S18084;
wire S18085;
wire S18086;
wire S18087;
wire S18088;
wire S18089;
wire S18090;
wire S18091;
wire S18092;
wire S18093;
wire S18094;
wire S18095;
wire S18096;
wire S18097;
wire S18098;
wire S18099;
wire S18100;
wire S18101;
wire S18102;
wire S18103;
wire S18104;
wire S18105;
wire S18106;
wire S18107;
wire S18108;
wire S18109;
wire S18110;
wire S18111;
wire S18112;
wire S18113;
wire S18114;
wire S18115;
wire S18116;
wire S18117;
wire S18118;
wire S18119;
wire S18120;
wire S18121;
wire S18122;
wire S18123;
wire S18124;
wire S18125;
wire S18126;
wire S18127;
wire S18128;
wire S18129;
wire S18130;
wire S18131;
wire S18132;
wire S18133;
wire S18134;
wire S18135;
wire S18136;
wire S18137;
wire S18138;
wire S18139;
wire S18140;
wire S18141;
wire S18142;
wire S18143;
wire S18144;
wire S18145;
wire S18146;
wire S18147;
wire S18148;
wire S18149;
wire S18150;
wire S18151;
wire S18152;
wire S18153;
wire S18154;
wire S18155;
wire S18156;
wire S18157;
wire S18158;
wire S18159;
wire S18160;
wire S18161;
wire S18162;
wire S18163;
wire S18164;
wire S18165;
wire S18166;
wire S18167;
wire S18168;
wire S18169;
wire S18170;
wire S18171;
wire S18172;
wire S18173;
wire S18174;
wire S18175;
wire S18176;
wire S18177;
wire S18178;
wire S18179;
wire S18180;
wire S18181;
wire S18182;
wire S18183;
wire S18184;
wire S18185;
wire S18186;
wire S18187;
wire S18188;
wire S18189;
wire S18190;
wire S18191;
wire S18192;
wire S18193;
wire S18194;
wire S18195;
wire S18196;
wire S18197;
wire S18198;
wire S18199;
wire S18200;
wire S18201;
wire S18202;
wire S18203;
wire S18204;
wire S18205;
wire S18206;
wire S18207;
wire S18208;
wire S18209;
wire S18210;
wire S18211;
wire S18212;
wire S18213;
wire S18214;
wire S18215;
wire S18216;
wire S18217;
wire S18218;
wire S18219;
wire S18220;
wire S18221;
wire S18222;
wire S18223;
wire S18224;
wire S18225;
wire S18226;
wire S18227;
wire S18228;
wire S18229;
wire S18230;
wire S18231;
wire S18232;
wire S18233;
wire S18234;
wire S18235;
wire S18236;
wire S18237;
wire S18238;
wire S18239;
wire S18240;
wire S18241;
wire S18242;
wire S18243;
wire S18244;
wire S18245;
wire S18246;
wire S18247;
wire S18248;
wire S18249;
wire S18250;
wire S18251;
wire S18252;
wire S18253;
wire S18254;
wire S18255;
wire S18256;
wire S18257;
wire S18258;
wire S18259;
wire S18260;
wire S18261;
wire S18262;
wire S18263;
wire S18264;
wire S18265;
wire S18266;
wire S18267;
wire S18268;
wire S18269;
wire S18270;
wire S18271;
wire S18272;
wire S18273;
wire S18274;
wire S18275;
wire S18276;
wire S18277;
wire S18278;
wire S18279;
wire S18280;
wire S18281;
wire S18282;
wire S18283;
wire S18284;
wire S18285;
wire S18286;
wire S18287;
wire S18288;
wire S18289;
wire S18290;
wire S18291;
wire S18292;
wire S18293;
wire S18294;
wire S18295;
wire S18296;
wire S18297;
wire S18298;
wire S18299;
wire S18300;
wire S18301;
wire S18302;
wire S18303;
wire S18304;
wire S18305;
wire S18306;
wire S18307;
wire S18308;
wire S18309;
wire S18310;
wire S18311;
wire S18312;
wire S18313;
wire S18314;
wire S18315;
wire S18316;
wire S18317;
wire S18318;
wire S18319;
wire S18320;
wire S18321;
wire S18322;
wire S18323;
wire S18324;
wire S18325;
wire S18326;
wire S18327;
wire S18328;
wire S18329;
wire S18330;
wire S18331;
wire S18332;
wire S18333;
wire S18334;
wire S18335;
wire S18336;
wire S18337;
wire S18338;
wire S18339;
wire S18340;
wire S18341;
wire S18342;
wire S18343;
wire S18344;
wire S18345;
wire S18346;
wire S18347;
wire S18348;
wire S18349;
wire S18350;
wire S18351;
wire S18352;
wire S18353;
wire S18354;
wire S18355;
wire S18356;
wire S18357;
wire S18358;
wire S18359;
wire S18360;
wire S18361;
wire S18362;
wire S18363;
wire S18364;
wire S18365;
wire S18366;
wire S18367;
wire S18368;
wire S18369;
wire S18370;
wire S18371;
wire S18372;
wire S18373;
wire S18374;
wire S18375;
wire S18376;
wire S18377;
wire S18378;
wire S18379;
wire S18380;
wire S18381;
wire S18382;
wire S18383;
wire S18384;
wire S18385;
wire S18386;
wire S18387;
wire S18388;
wire S18389;
wire S18390;
wire S18391;
wire S18392;
wire S18393;
wire S18394;
wire S18395;
wire S18396;
wire S18397;
wire S18398;
wire S18399;
wire S18400;
wire S18401;
wire S18402;
wire S18403;
wire S18404;
wire S18405;
wire S18406;
wire S18407;
wire S18408;
wire S18409;
wire S18410;
wire S18411;
wire S18412;
wire S18413;
wire S18414;
wire S18415;
wire S18416;
wire S18417;
wire S18418;
wire S18419;
wire S18420;
wire S18421;
wire S18422;
wire S18423;
wire S18424;
wire S18425;
wire S18426;
wire S18427;
wire S18428;
wire S18429;
wire S18430;
wire S18431;
wire S18432;
wire S18433;
wire S18434;
wire S18435;
wire S18436;
wire S18437;
wire S18438;
wire S18439;
wire S18440;
wire S18441;
wire S18442;
wire S18443;
wire S18444;
wire S18445;
wire S18446;
wire S18447;
wire S18448;
wire S18449;
wire S18450;
wire S18451;
wire S18452;
wire S18453;
wire S18454;
wire S18455;
wire S18456;
wire S18457;
wire S18458;
wire S18459;
wire S18460;
wire S18461;
wire S18462;
wire S18463;
wire S18464;
wire S18465;
wire S18466;
wire S18467;
wire S18468;
wire S18469;
wire S18470;
wire S18471;
wire S18472;
wire S18473;
wire S18474;
wire S18475;
wire S18476;
wire S18477;
wire S18478;
wire S18479;
wire S18480;
wire S18481;
wire S18482;
wire S18483;
wire S18484;
wire S18485;
wire S18486;
wire S18487;
wire S18488;
wire S18489;
wire S18490;
wire S18491;
wire S18492;
wire S18493;
wire S18494;
wire S18495;
wire S18496;
wire S18497;
wire S18498;
wire S18499;
wire S18500;
wire S18501;
wire S18502;
wire S18503;
wire S18504;
wire S18505;
wire S18506;
wire S18507;
wire S18508;
wire S18509;
wire S18510;
wire S18511;
wire S18512;
wire S18513;
wire S18514;
wire S18515;
wire S18516;
wire S18517;
wire S18518;
wire S18519;
wire S18520;
wire S18521;
wire S18522;
wire S18523;
wire S18524;
wire S18525;
wire S18526;
wire S18527;
wire S18528;
wire S18529;
wire S18530;
wire S18531;
wire S18532;
wire S18533;
wire S18534;
wire S18535;
wire S18536;
wire S18537;
wire S18538;
wire S18539;
wire S18540;
wire S18541;
wire S18542;
wire S18543;
wire S18544;
wire S18545;
wire S18546;
wire S18547;
wire S18548;
wire S18549;
wire S18550;
wire S18551;
wire S18552;
wire S18553;
wire S18554;
wire S18555;
wire S18556;
wire S18557;
wire S18558;
wire S18559;
wire S18560;
wire S18561;
wire S18562;
wire S18563;
wire S18564;
wire S18565;
wire S18566;
wire S18567;
wire S18568;
wire S18569;
wire S18570;
wire S18571;
wire S18572;
wire S18573;
wire S18574;
wire S18575;
wire S18576;
wire S18577;
wire S18578;
wire S18579;
wire S18580;
wire S18581;
wire S18582;
wire S18583;
wire S18584;
wire S18585;
wire S18586;
wire S18587;
wire S18588;
wire S18589;
wire S18590;
wire S18591;
wire S18592;
wire S18593;
wire S18594;
wire S18595;
wire S18596;
wire S18597;
wire S18598;
wire S18599;
wire S18600;
wire S18601;
wire S18602;
wire S18603;
wire S18604;
wire S18605;
wire S18606;
wire S18607;
wire S18608;
wire S18609;
wire S18610;
wire S18611;
wire S18612;
wire S18613;
wire S18614;
wire S18615;
wire S18616;
wire S18617;
wire S18618;
wire S18619;
wire S18620;
wire S18621;
wire S18622;
wire S18623;
wire S18624;
wire S18625;
wire S18626;
wire S18627;
wire S18628;
wire S18629;
wire S18630;
wire S18631;
wire S18632;
wire S18633;
wire S18634;
wire S18635;
wire S18636;
wire S18637;
wire S18638;
wire S18639;
wire S18640;
wire S18641;
wire S18642;
wire S18643;
wire S18644;
wire S18645;
wire S18646;
wire S18647;
wire S18648;
wire S18649;
wire S18650;
wire S18651;
wire S18652;
wire S18653;
wire S18654;
wire S18655;
wire S18656;
wire S18657;
wire S18658;
wire S18659;
wire S18660;
wire S18661;
wire S18662;
wire S18663;
wire S18664;
wire S18665;
wire S18666;
wire S18667;
wire S18668;
wire S18669;
wire S18670;
wire S18671;
wire S18672;
wire S18673;
wire S18674;
wire S18675;
wire S18676;
wire S18677;
wire S18678;
wire S18679;
wire S18680;
wire S18681;
wire S18682;
wire S18683;
wire S18684;
wire S18685;
wire S18686;
wire S18687;
wire S18688;
wire S18689;
wire S18690;
wire S18691;
wire S18692;
wire S18693;
wire S18694;
wire S18695;
wire S18696;
wire S18697;
wire S18698;
wire S18699;
wire S18700;
wire S18701;
wire S18702;
wire S18703;
wire S18704;
wire S18705;
wire S18706;
wire S18707;
wire S18708;
wire S18709;
wire S18710;
wire S18711;
wire S18712;
wire S18713;
wire S18714;
wire S18715;
wire S18716;
wire S18717;
wire S18718;
wire S18719;
wire S18720;
wire S18721;
wire S18722;
wire S18723;
wire S18724;
wire S18725;
wire S18726;
wire S18727;
wire S18728;
wire S18729;
wire S18730;
wire S18731;
wire S18732;
wire S18733;
wire S18734;
wire S18735;
wire S18736;
wire S18737;
wire S18738;
wire S18739;
wire S18740;
wire S18741;
wire S18742;
wire S18743;
wire S18744;
wire S18745;
wire S18746;
wire S18747;
wire S18748;
wire S18749;
wire S18750;
wire S18751;
wire S18752;
wire S18753;
wire S18754;
wire S18755;
wire S18756;
wire S18757;
wire S18758;
wire S18759;
wire S18760;
wire S18761;
wire S18762;
wire S18763;
wire S18764;
wire S18765;
wire S18766;
wire S18767;
wire S18768;
wire S18769;
wire S18770;
wire S18771;
wire S18772;
wire S18773;
wire S18774;
wire S18775;
wire S18776;
wire S18777;
wire S18778;
wire S18779;
wire S18780;
wire S18781;
wire S18782;
wire S18783;
wire S18784;
wire S18785;
wire S18786;
wire S18787;
wire S18788;
wire S18789;
wire S18790;
wire S18791;
wire S18792;
wire S18793;
wire S18794;
wire S18795;
wire S18796;
wire S18797;
wire S18798;
wire S18799;
wire S18800;
wire S18801;
wire S18802;
wire S18803;
wire S18804;
wire S18805;
wire S18806;
wire S18807;
wire S18808;
wire S18809;
wire S18810;
wire S18811;
wire S18812;
wire S18813;
wire S18814;
wire S18815;
wire S18816;
wire S18817;
wire S18818;
wire S18819;
wire S18820;
wire S18821;
wire S18822;
wire S18823;
wire S18824;
wire S18825;
wire S18826;
wire S18827;
wire S18828;
wire S18829;
wire S18830;
wire S18831;
wire S18832;
wire S18833;
wire S18834;
wire S18835;
wire S18836;
wire S18837;
wire S18838;
wire S18839;
wire S18840;
wire S18841;
wire S18842;
wire S18843;
wire S18844;
wire S18845;
wire S18846;
wire S18847;
wire S18848;
wire S18849;
wire S18850;
wire S18851;
wire S18852;
wire S18853;
wire S18854;
wire S18855;
wire S18856;
wire S18857;
wire S18858;
wire S18859;
wire S18860;
wire S18861;
wire S18862;
wire S18863;
wire S18864;
wire S18865;
wire S18866;
wire S18867;
wire S18868;
wire S18869;
wire S18870;
wire S18871;
wire S18872;
wire S18873;
wire S18874;
wire S18875;
wire S18876;
wire S18877;
wire S18878;
wire S18879;
wire S18880;
wire S18881;
wire S18882;
wire S18883;
wire S18884;
wire S18885;
wire S18886;
wire S18887;
wire S18888;
wire S18889;
wire S18890;
wire S18891;
wire S18892;
wire S18893;
wire S18894;
wire S18895;
wire S18896;
wire S18897;
wire S18898;
wire S18899;
wire S18900;
wire S18901;
wire S18902;
wire S18903;
wire S18904;
wire S18905;
wire S18906;
wire S18907;
wire S18908;
wire S18909;
wire S18910;
wire S18911;
wire S18912;
wire S18913;
wire S18914;
wire S18915;
wire S18916;
wire S18917;
wire S18918;
wire S18919;
wire S18920;
wire S18921;
wire S18922;
wire S18923;
wire S18924;
wire S18925;
wire S18926;
wire S18927;
wire S18928;
wire S18929;
wire S18930;
wire S18931;
wire S18932;
wire S18933;
wire S18934;
wire S18935;
wire S18936;
wire S18937;
wire S18938;
wire S18939;
wire S18940;
wire S18941;
wire S18942;
wire S18943;
wire S18944;
wire S18945;
wire S18946;
wire S18947;
wire S18948;
wire S18949;
wire S18950;
wire S18951;
wire S18952;
wire S18953;
wire S18954;
wire S18955;
wire S18956;
wire S18957;
wire S18958;
wire S18959;
wire S18960;
wire S18961;
wire S18962;
wire S18963;
wire S18964;
wire S18965;
wire S18966;
wire S18967;
wire S18968;
wire S18969;
wire S18970;
wire S18971;
wire S18972;
wire S18973;
wire S18974;
wire S18975;
wire S18976;
wire S18977;
wire S18978;
wire S18979;
wire S18980;
wire S18981;
wire S18982;
wire S18983;
wire S18984;
wire S18985;
wire S18986;
wire S18987;
wire S18988;
wire S18989;
wire S18990;
wire S18991;
wire S18992;
wire S18993;
wire S18994;
wire S18995;
wire S18996;
wire S18997;
wire S18998;
wire S18999;
wire S19000;
wire S19001;
wire S19002;
wire S19003;
wire S19004;
wire S19005;
wire S19006;
wire S19007;
wire S19008;
wire S19009;
wire S19010;
wire S19011;
wire S19012;
wire S19013;
wire S19014;
wire S19015;
wire S19016;
wire S19017;
wire S19018;
wire S19019;
wire S19020;
wire S19021;
wire S19022;
wire S19023;
wire S19024;
wire S19025;
wire S19026;
wire S19027;
wire S19028;
wire S19029;
wire S19030;
wire S19031;
wire S19032;
wire S19033;
wire S19034;
wire S19035;
wire S19036;
wire S19037;
wire S19038;
wire S19039;
wire S19040;
wire S19041;
wire S19042;
wire S19043;
wire S19044;
wire S19045;
wire S19046;
wire S19047;
wire S19048;
wire S19049;
wire S19050;
wire S19051;
wire S19052;
wire S19053;
wire S19054;
wire S19055;
wire S19056;
wire S19057;
wire S19058;
wire S19059;
wire S19060;
wire S19061;
wire S19062;
wire S19063;
wire S19064;
wire S19065;
wire S19066;
wire S19067;
wire S19068;
wire S19069;
wire S19070;
wire S19071;
wire S19072;
wire S19073;
wire S19074;
wire S19075;
wire S19076;
wire S19077;
wire S19078;
wire S19079;
wire S19080;
wire S19081;
wire S19082;
wire S19083;
wire S19084;
wire S19085;
wire S19086;
wire S19087;
wire S19088;
wire S19089;
wire S19090;
wire S19091;
wire S19092;
wire S19093;
wire S19094;
wire S19095;
wire S19096;
wire S19097;
wire S19098;
wire S19099;
wire S19100;
wire S19101;
wire S19102;
wire S19103;
wire S19104;
wire S19105;
wire S19106;
wire S19107;
wire S19108;
wire S19109;
wire S19110;
wire S19111;
wire S19112;
wire S19113;
wire S19114;
wire S19115;
wire S19116;
wire S19117;
wire S19118;
wire S19119;
wire S19120;
wire S19121;
wire S19122;
wire S19123;
wire S19124;
wire S19125;
wire S19126;
wire S19127;
wire S19128;
wire S19129;
wire S19130;
wire S19131;
wire S19132;
wire S19133;
wire S19134;
wire S19135;
wire S19136;
wire S19137;
wire S19138;
wire S19139;
wire S19140;
wire S19141;
wire S19142;
wire S19143;
wire S19144;
wire S19145;
wire S19146;
wire S19147;
wire S19148;
wire S19149;
wire S19150;
wire S19151;
wire S19152;
wire S19153;
wire S19154;
wire S19155;
wire S19156;
wire S19157;
wire S19158;
wire S19159;
wire S19160;
wire S19161;
wire S19162;
wire S19163;
wire S19164;
wire S19165;
wire S19166;
wire S19167;
wire S19168;
wire S19169;
wire S19170;
wire S19171;
wire S19172;
wire S19173;
wire S19174;
wire S19175;
wire S19176;
wire S19177;
wire S19178;
wire S19179;
wire S19180;
wire S19181;
wire S19182;
wire S19183;
wire S19184;
wire S19185;
wire S19186;
wire S19187;
wire S19188;
wire S19189;
wire S19190;
wire S19191;
wire S19192;
wire S19193;
wire S19194;
wire S19195;
wire S19196;
wire S19197;
wire S19198;
wire S19199;
wire S19200;
wire S19201;
wire S19202;
wire S19203;
wire S19204;
wire S19205;
wire S19206;
wire S19207;
wire S19208;
wire S19209;
wire S19210;
wire S19211;
wire S19212;
wire S19213;
wire S19214;
wire S19215;
wire S19216;
wire S19217;
wire S19218;
wire S19219;
wire S19220;
wire S19221;
wire S19222;
wire S19223;
wire S19224;
wire S19225;
wire S19226;
wire S19227;
wire S19228;
wire S19229;
wire S19230;
wire S19231;
wire S19232;
wire S19233;
wire S19234;
wire S19235;
wire S19236;
wire S19237;
wire S19238;
wire S19239;
wire S19240;
wire S19241;
wire S19242;
wire S19243;
wire S19244;
wire S19245;
wire S19246;
wire S19247;
wire S19248;
wire S19249;
wire S19250;
wire S19251;
wire S19252;
wire S19253;
wire S19254;
wire S19255;
wire S19256;
wire S19257;
wire S19258;
wire S19259;
wire S19260;
wire S19261;
wire S19262;
wire S19263;
wire S19264;
wire S19265;
wire S19266;
wire S19267;
wire S19268;
wire S19269;
wire S19270;
wire S19271;
wire S19272;
wire S19273;
wire S19274;
wire S19275;
wire S19276;
wire S19277;
wire S19278;
wire S19279;
wire S19280;
wire S19281;
wire S19282;
wire S19283;
wire S19284;
wire S19285;
wire S19286;
wire S19287;
wire S19288;
wire S19289;
wire S19290;
wire S19291;
wire S19292;
wire S19293;
wire S19294;
wire S19295;
wire S19296;
wire S19297;
wire S19298;
wire S19299;
wire S19300;
wire S19301;
wire S19302;
wire S19303;
wire S19304;
wire S19305;
wire S19306;
wire S19307;
wire S19308;
wire S19309;
wire S19310;
wire S19311;
wire S19312;
wire S19313;
wire S19314;
wire S19315;
wire S19316;
wire S19317;
wire S19318;
wire S19319;
wire S19320;
wire S19321;
wire S19322;
wire S19323;
wire S19324;
wire S19325;
wire S19326;
wire S19327;
wire S19328;
wire S19329;
wire S19330;
wire S19331;
wire S19332;
wire S19333;
wire S19334;
wire S19335;
wire S19336;
wire S19337;
wire S19338;
wire S19339;
wire S19340;
wire S19341;
wire S19342;
wire S19343;
wire S19344;
wire S19345;
wire S19346;
wire S19347;
wire S19348;
wire S19349;
wire S19350;
wire S19351;
wire S19352;
wire S19353;
wire S19354;
wire S19355;
wire S19356;
wire S19357;
wire S19358;
wire S19359;
wire S19360;
wire S19361;
wire S19362;
wire S19363;
wire S19364;
wire S19365;
wire S19366;
wire S19367;
wire S19368;
wire S19369;
wire S19370;
wire S19371;
wire S19372;
wire S19373;
wire S19374;
wire S19375;
wire S19376;
wire S19377;
wire S19378;
wire S19379;
wire S19380;
wire S19381;
wire S19382;
wire S19383;
wire S19384;
wire S19385;
wire S19386;
wire S19387;
wire S19388;
wire S19389;
wire S19390;
wire S19391;
wire S19392;
wire S19393;
wire S19394;
wire S19395;
wire S19396;
wire S19397;
wire S19398;
wire S19399;
wire S19400;
wire S19401;
wire S19402;
wire S19403;
wire S19404;
wire S19405;
wire S19406;
wire S19407;
wire S19408;
wire S19409;
wire S19410;
wire S19411;
wire S19412;
wire S19413;
wire S19414;
wire S19415;
wire S19416;
wire S19417;
wire S19418;
wire S19419;
wire S19420;
wire S19421;
wire S19422;
wire S19423;
wire S19424;
wire S19425;
wire S19426;
wire S19427;
wire S19428;
wire S19429;
wire S19430;
wire S19431;
wire S19432;
wire S19433;
wire S19434;
wire S19435;
wire S19436;
wire S19437;
wire S19438;
wire S19439;
wire S19440;
wire S19441;
wire S19442;
wire S19443;
wire S19444;
wire S19445;
wire S19446;
wire S19447;
wire S19448;
wire S19449;
wire S19450;
wire S19451;
wire S19452;
wire S19453;
wire S19454;
wire S19455;
wire S19456;
wire S19457;
wire S19458;
wire S19459;
wire S19460;
wire S19461;
wire S19462;
wire S19463;
wire S19464;
wire S19465;
wire S19466;
wire S19467;
wire S19468;
wire S19469;
wire S19470;
wire S19471;
wire S19472;
wire S19473;
wire S19474;
wire S19475;
wire S19476;
wire S19477;
wire S19478;
wire S19479;
wire S19480;
wire S19481;
wire S19482;
wire S19483;
wire S19484;
wire S19485;
wire S19486;
wire S19487;
wire S19488;
wire S19489;
wire S19490;
wire S19491;
wire S19492;
wire S19493;
wire S19494;
wire S19495;
wire S19496;
wire S19497;
wire S19498;
wire S19499;
wire S19500;
wire S19501;
wire S19502;
wire S19503;
wire S19504;
wire S19505;
wire S19506;
wire S19507;
wire S19508;
wire S19509;
wire S19510;
wire S19511;
wire S19512;
wire S19513;
wire S19514;
wire S19515;
wire S19516;
wire S19517;
wire S19518;
wire S19519;
wire S19520;
wire S19521;
wire S19522;
wire S19523;
wire S19524;
wire S19525;
wire S19526;
wire S19527;
wire S19528;
wire S19529;
wire S19530;
wire S19531;
wire S19532;
wire S19533;
wire S19534;
wire S19535;
wire S19536;
wire S19537;
wire S19538;
wire S19539;
wire S19540;
wire S19541;
wire S19542;
wire S19543;
wire S19544;
wire S19545;
wire S19546;
wire S19547;
wire S19548;
wire S19549;
wire S19550;
wire S19551;
wire S19552;
wire S19553;
wire S19554;
wire S19555;
wire S19556;
wire S19557;
wire S19558;
wire S19559;
wire S19560;
wire S19561;
wire S19562;
wire S19563;
wire S19564;
wire S19565;
wire S19566;
wire S19567;
wire S19568;
wire S19569;
wire S19570;
wire S19571;
wire S19572;
wire S19573;
wire S19574;
wire S19575;
wire S19576;
wire S19577;
wire S19578;
wire S19579;
wire S19580;
wire S19581;
wire S19582;
wire S19583;
wire S19584;
wire S19585;
wire S19586;
wire S19587;
wire S19588;
wire S19589;
wire S19590;
wire S19591;
wire S19592;
wire S19593;
wire S19594;
wire S19595;
wire S19596;
wire S19597;
wire S19598;
wire S19599;
wire S19600;
wire S19601;
wire S19602;
wire S19603;
wire S19604;
wire S19605;
wire S19606;
wire S19607;
wire S19608;
wire S19609;
wire S19610;
wire S19611;
wire S19612;
wire S19613;
wire S19614;
wire S19615;
wire S19616;
wire S19617;
wire S19618;
wire S19619;
wire S19620;
wire S19621;
wire S19622;
wire S19623;
wire S19624;
wire S19625;
wire S19626;
wire S19627;
wire S19628;
wire S19629;
wire S19630;
wire S19631;
wire S19632;
wire S19633;
wire S19634;
wire S19635;
wire S19636;
wire S19637;
wire S19638;
wire S19639;
wire S19640;
wire S19641;
wire S19642;
wire S19643;
wire S19644;
wire S19645;
wire S19646;
wire S19647;
wire S19648;
wire S19649;
wire S19650;
wire S19651;
wire S19652;
wire S19653;
wire S19654;
wire S19655;
wire S19656;
wire S19657;
wire S19658;
wire S19659;
wire S19660;
wire S19661;
wire S19662;
wire S19663;
wire S19664;
wire S19665;
wire S19666;
wire S19667;
wire S19668;
wire S19669;
wire S19670;
wire S19671;
wire S19672;
wire S19673;
wire S19674;
wire S19675;
wire S19676;
wire S19677;
wire S19678;
wire S19679;
wire S19680;
wire S19681;
wire S19682;
wire S19683;
wire S19684;
wire S19685;
wire S19686;
wire S19687;
wire S19688;
wire S19689;
wire S19690;
wire S19691;
wire S19692;
wire S19693;
wire S19694;
wire S19695;
wire S19696;
wire S19697;
wire S19698;
wire S19699;
wire S19700;
wire S19701;
wire S19702;
wire S19703;
wire S19704;
wire S19705;
wire S19706;
wire S19707;
wire S19708;
wire S19709;
wire S19710;
wire S19711;
wire S19712;
wire S19713;
wire S19714;
wire S19715;
wire S19716;
wire S19717;
wire S19718;
wire S19719;
wire S19720;
wire S19721;
wire S19722;
wire S19723;
wire S19724;
wire S19725;
wire S19726;
wire S19727;
wire S19728;
wire S19729;
wire S19730;
wire S19731;
wire S19732;
wire S19733;
wire S19734;
wire S19735;
wire S19736;
wire S19737;
wire S19738;
wire S19739;
wire S19740;
wire S19741;
wire S19742;
wire S19743;
wire S19744;
wire S19745;
wire S19746;
wire S19747;
wire S19748;
wire S19749;
wire S19750;
wire S19751;
wire S19752;
wire S19753;
wire S19754;
wire S19755;
wire S19756;
wire S19757;
wire S19758;
wire S19759;
wire S19760;
wire S19761;
wire S19762;
wire S19763;
wire S19764;
wire S19765;
wire S19766;
wire S19767;
wire S19768;
wire S19769;
wire S19770;
wire S19771;
wire S19772;
wire S19773;
wire S19774;
wire S19775;
wire S19776;
wire S19777;
wire S19778;
wire S19779;
wire S19780;
wire S19781;
wire S19782;
wire S19783;
wire S19784;
wire S19785;
wire S19786;
wire S19787;
wire S19788;
wire S19789;
wire S19790;
wire S19791;
wire S19792;
wire S19793;
wire S19794;
wire S19795;
wire S19796;
wire S19797;
wire S19798;
wire S19799;
wire S19800;
wire S19801;
wire S19802;
wire S19803;
wire S19804;
wire S19805;
wire S19806;
wire S19807;
wire S19808;
wire S19809;
wire S19810;
wire S19811;
wire S19812;
wire S19813;
wire S19814;
wire S19815;
wire S19816;
wire S19817;
wire S19818;
wire S19819;
wire S19820;
wire S19821;
wire S19822;
wire S19823;
wire S19824;
wire S19825;
wire S19826;
wire S19827;
wire S19828;
wire S19829;
wire S19830;
wire S19831;
wire S19832;
wire S19833;
wire S19834;
wire S19835;
wire S19836;
wire S19837;
wire S19838;
wire S19839;
wire S19840;
wire S19841;
wire S19842;
wire S19843;
wire S19844;
wire S19845;
wire S19846;
wire S19847;
wire S19848;
wire S19849;
wire S19850;
wire S19851;
wire S19852;
wire S19853;
wire S19854;
wire S19855;
wire S19856;
wire S19857;
wire S19858;
wire S19859;
wire S19860;
wire S19861;
wire S19862;
wire S19863;
wire S19864;
wire S19865;
wire S19866;
wire S19867;
wire S19868;
wire S19869;
wire S19870;
wire S19871;
wire S19872;
wire S19873;
wire S19874;
wire S19875;
wire S19876;
wire S19877;
wire S19878;
wire S19879;
wire S19880;
wire S19881;
wire S19882;
wire S19883;
wire S19884;
wire S19885;
wire S19886;
wire S19887;
wire S19888;
wire S19889;
wire S19890;
wire S19891;
wire S19892;
wire S19893;
wire S19894;
wire S19895;
wire S19896;
wire S19897;
wire S19898;
wire S19899;
wire S19900;
wire S19901;
wire S19902;
wire S19903;
wire S19904;
wire S19905;
wire S19906;
wire S19907;
wire S19908;
wire S19909;
wire S19910;
wire S19911;
wire S19912;
wire S19913;
wire S19914;
wire S19915;
wire S19916;
wire S19917;
wire S19918;
wire S19919;
wire S19920;
wire S19921;
wire S19922;
wire S19923;
wire S19924;
wire S19925;
wire S19926;
wire S19927;
wire S19928;
wire S19929;
wire S19930;
wire S19931;
wire S19932;
wire S19933;
wire S19934;
wire S19935;
wire S19936;
wire S19937;
wire S19938;
wire S19939;
wire S19940;
wire S19941;
wire S19942;
wire S19943;
wire S19944;
wire S19945;
wire S19946;
wire S19947;
wire S19948;
wire S19949;
wire S19950;
wire S19951;
wire S19952;
wire S19953;
wire S19954;
wire S19955;
wire S19956;
wire S19957;
wire S19958;
wire S19959;
wire S19960;
wire S19961;
wire S19962;
wire S19963;
wire S19964;
wire S19965;
wire S19966;
wire S19967;
wire S19968;
wire S19969;
wire S19970;
wire S19971;
wire S19972;
wire S19973;
wire S19974;
wire S19975;
wire S19976;
wire S19977;
wire S19978;
wire S19979;
wire S19980;
wire S19981;
wire S19982;
wire S19983;
wire S19984;
wire S19985;
wire S19986;
wire S19987;
wire S19988;
wire S19989;
wire S19990;
wire S19991;
wire S19992;
wire S19993;
wire S19994;
wire S19995;
wire S19996;
wire S19997;
wire S19998;
wire S19999;
wire S20000;
wire S20001;
wire S20002;
wire S20003;
wire S20004;
wire S20005;
wire S20006;
wire S20007;
wire S20008;
wire S20009;
wire S20010;
wire S20011;
wire S20012;
wire S20013;
wire S20014;
wire S20015;
wire S20016;
wire S20017;
wire S20018;
wire S20019;
wire S20020;
wire S20021;
wire S20022;
wire S20023;
wire S20024;
wire S20025;
wire S20026;
wire S20027;
wire S20028;
wire S20029;
wire S20030;
wire S20031;
wire S20032;
wire S20033;
wire S20034;
wire S20035;
wire S20036;
wire S20037;
wire S20038;
wire S20039;
wire S20040;
wire S20041;
wire S20042;
wire S20043;
wire S20044;
wire S20045;
wire S20046;
wire S20047;
wire S20048;
wire S20049;
wire S20050;
wire S20051;
wire S20052;
wire S20053;
wire S20054;
wire S20055;
wire S20056;
wire S20057;
wire S20058;
wire S20059;
wire S20060;
wire S20061;
wire S20062;
wire S20063;
wire S20064;
wire S20065;
wire S20066;
wire S20067;
wire S20068;
wire S20069;
wire S20070;
wire S20071;
wire S20072;
wire S20073;
wire S20074;
wire S20075;
wire S20076;
wire S20077;
wire S20078;
wire S20079;
wire S20080;
wire S20081;
wire S20082;
wire S20083;
wire S20084;
wire S20085;
wire S20086;
wire S20087;
wire S20088;
wire S20089;
wire S20090;
wire S20091;
wire S20092;
wire S20093;
wire S20094;
wire S20095;
wire S20096;
wire S20097;
wire S20098;
wire S20099;
wire S20100;
wire S20101;
wire S20102;
wire S20103;
wire S20104;
wire S20105;
wire S20106;
wire S20107;
wire S20108;
wire S20109;
wire S20110;
wire S20111;
wire S20112;
wire S20113;
wire S20114;
wire S20115;
wire S20116;
wire S20117;
wire S20118;
wire S20119;
wire S20120;
wire S20121;
wire S20122;
wire S20123;
wire S20124;
wire S20125;
wire S20126;
wire S20127;
wire S20128;
wire S20129;
wire S20130;
wire S20131;
wire S20132;
wire S20133;
wire S20134;
wire S20135;
wire S20136;
wire S20137;
wire S20138;
wire S20139;
wire S20140;
wire S20141;
wire S20142;
wire S20143;
wire S20144;
wire S20145;
wire S20146;
wire S20147;
wire S20148;
wire S20149;
wire S20150;
wire S20151;
wire S20152;
wire S20153;
wire S20154;
wire S20155;
wire S20156;
wire S20157;
wire S20158;
wire S20159;
wire S20160;
wire S20161;
wire S20162;
wire S20163;
wire S20164;
wire S20165;
wire S20166;
wire S20167;
wire S20168;
wire S20169;
wire S20170;
wire S20171;
wire S20172;
wire S20173;
wire S20174;
wire S20175;
wire S20176;
wire S20177;
wire S20178;
wire S20179;
wire S20180;
wire S20181;
wire S20182;
wire S20183;
wire S20184;
wire S20185;
wire S20186;
wire S20187;
wire S20188;
wire S20189;
wire S20190;
wire S20191;
wire S20192;
wire S20193;
wire S20194;
wire S20195;
wire S20196;
wire S20197;
wire S20198;
wire S20199;
wire S20200;
wire S20201;
wire S20202;
wire S20203;
wire S20204;
wire S20205;
wire S20206;
wire S20207;
wire S20208;
wire S20209;
wire S20210;
wire S20211;
wire S20212;
wire S20213;
wire S20214;
wire S20215;
wire S20216;
wire S20217;
wire S20218;
wire S20219;
wire S20220;
wire S20221;
wire S20222;
wire S20223;
wire S20224;
wire S20225;
wire S20226;
wire S20227;
wire S20228;
wire S20229;
wire S20230;
wire S20231;
wire S20232;
wire S20233;
wire S20234;
wire S20235;
wire S20236;
wire S20237;
wire S20238;
wire S20239;
wire S20240;
wire S20241;
wire S20242;
wire S20243;
wire S20244;
wire S20245;
wire S20246;
wire S20247;
wire S20248;
wire S20249;
wire S20250;
wire S20251;
wire S20252;
wire S20253;
wire S20254;
wire S20255;
wire S20256;
wire S20257;
wire S20258;
wire S20259;
wire S20260;
wire S20261;
wire S20262;
wire S20263;
wire S20264;
wire S20265;
wire S20266;
wire S20267;
wire S20268;
wire S20269;
wire S20270;
wire S20271;
wire S20272;
wire S20273;
wire S20274;
wire S20275;
wire S20276;
wire S20277;
wire S20278;
wire S20279;
wire S20280;
wire S20281;
wire S20282;
wire S20283;
wire S20284;
wire S20285;
wire S20286;
wire S20287;
wire S20288;
wire S20289;
wire S20290;
wire S20291;
wire S20292;
wire S20293;
wire S20294;
wire S20295;
wire S20296;
wire S20297;
wire S20298;
wire S20299;
wire S20300;
wire S20301;
wire S20302;
wire S20303;
wire S20304;
wire S20305;
wire S20306;
wire S20307;
wire S20308;
wire S20309;
wire S20310;
wire S20311;
wire S20312;
wire S20313;
wire S20314;
wire S20315;
wire S20316;
wire S20317;
wire S20318;
wire S20319;
wire S20320;
wire S20321;
wire S20322;
wire S20323;
wire S20324;
wire S20325;
wire S20326;
wire S20327;
wire S20328;
wire S20329;
wire S20330;
wire S20331;
wire S20332;
wire S20333;
wire S20334;
wire S20335;
wire S20336;
wire S20337;
wire S20338;
wire S20339;
wire S20340;
wire S20341;
wire S20342;
wire S20343;
wire S20344;
wire S20345;
wire S20346;
wire S20347;
wire S20348;
wire S20349;
wire S20350;
wire S20351;
wire S20352;
wire S20353;
wire S20354;
wire S20355;
wire S20356;
wire S20357;
wire S20358;
wire S20359;
wire S20360;
wire S20361;
wire S20362;
wire S20363;
wire S20364;
wire S20365;
wire S20366;
wire S20367;
wire S20368;
wire S20369;
wire S20370;
wire S20371;
wire S20372;
wire S20373;
wire S20374;
wire S20375;
wire S20376;
wire S20377;
wire S20378;
wire S20379;
wire S20380;
wire S20381;
wire S20382;
wire S20383;
wire S20384;
wire S20385;
wire S20386;
wire S20387;
wire S20388;
wire S20389;
wire S20390;
wire S20391;
wire S20392;
wire S20393;
wire S20394;
wire S20395;
wire S20396;
wire S20397;
wire S20398;
wire S20399;
wire S20400;
wire S20401;
wire S20402;
wire S20403;
wire S20404;
wire S20405;
wire S20406;
wire S20407;
wire S20408;
wire S20409;
wire S20410;
wire S20411;
wire S20412;
wire S20413;
wire S20414;
wire S20415;
wire S20416;
wire S20417;
wire S20418;
wire S20419;
wire S20420;
wire S20421;
wire S20422;
wire S20423;
wire S20424;
wire S20425;
wire S20426;
wire S20427;
wire S20428;
wire S20429;
wire S20430;
wire S20431;
wire S20432;
wire S20433;
wire S20434;
wire S20435;
wire S20436;
wire S20437;
wire S20438;
wire S20439;
wire S20440;
wire S20441;
wire S20442;
wire S20443;
wire S20444;
wire S20445;
wire S20446;
wire S20447;
wire S20448;
wire S20449;
wire S20450;
wire S20451;
wire S20452;
wire S20453;
wire S20454;
wire S20455;
wire S20456;
wire S20457;
wire S20458;
wire S20459;
wire S20460;
wire S20461;
wire S20462;
wire S20463;
wire S20464;
wire S20465;
wire S20466;
wire S20467;
wire S20468;
wire S20469;
wire S20470;
wire S20471;
wire S20472;
wire S20473;
wire S20474;
wire S20475;
wire S20476;
wire S20477;
wire S20478;
wire S20479;
wire S20480;
wire S20481;
wire S20482;
wire S20483;
wire S20484;
wire S20485;
wire S20486;
wire S20487;
wire S20488;
wire S20489;
wire S20490;
wire S20491;
wire S20492;
wire S20493;
wire S20494;
wire S20495;
wire S20496;
wire S20497;
wire S20498;
wire S20499;
wire S20500;
wire S20501;
wire S20502;
wire S20503;
wire S20504;
wire S20505;
wire S20506;
wire S20507;
wire S20508;
wire S20509;
wire S20510;
wire S20511;
wire S20512;
wire S20513;
wire S20514;
wire S20515;
wire S20516;
wire S20517;
wire S20518;
wire S20519;
wire S20520;
wire S20521;
wire S20522;
wire S20523;
wire S20524;
wire S20525;
wire S20526;
wire S20527;
wire S20528;
wire S20529;
wire S20530;
wire S20531;
wire S20532;
wire S20533;
wire S20534;
wire S20535;
wire S20536;
wire S20537;
wire S20538;
wire S20539;
wire S20540;
wire S20541;
wire S20542;
wire S20543;
wire S20544;
wire S20545;
wire S20546;
wire S20547;
wire S20548;
wire S20549;
wire S20550;
wire S20551;
wire S20552;
wire S20553;
wire S20554;
wire S20555;
wire S20556;
wire S20557;
wire S20558;
wire S20559;
wire S20560;
wire S20561;
wire S20562;
wire S20563;
wire S20564;
wire S20565;
wire S20566;
wire S20567;
wire S20568;
wire S20569;
wire S20570;
wire S20571;
wire S20572;
wire S20573;
wire S20574;
wire S20575;
wire S20576;
wire S20577;
wire S20578;
wire S20579;
wire S20580;
wire S20581;
wire S20582;
wire S20583;
wire S20584;
wire S20585;
wire S20586;
wire S20587;
wire S20588;
wire S20589;
wire S20590;
wire S20591;
wire S20592;
wire S20593;
wire S20594;
wire S20595;
wire S20596;
wire S20597;
wire S20598;
wire S20599;
wire S20600;
wire S20601;
wire S20602;
wire S20603;
wire S20604;
wire S20605;
wire S20606;
wire S20607;
wire S20608;
wire S20609;
wire S20610;
wire S20611;
wire S20612;
wire S20613;
wire S20614;
wire S20615;
wire S20616;
wire S20617;
wire S20618;
wire S20619;
wire S20620;
wire S20621;
wire S20622;
wire S20623;
wire S20624;
wire S20625;
wire S20626;
wire S20627;
wire S20628;
wire S20629;
wire S20630;
wire S20631;
wire S20632;
wire S20633;
wire S20634;
wire S20635;
wire S20636;
wire S20637;
wire S20638;
wire S20639;
wire S20640;
wire S20641;
wire S20642;
wire S20643;
wire S20644;
wire S20645;
wire S20646;
wire S20647;
wire S20648;
wire S20649;
wire S20650;
wire S20651;
wire S20652;
wire S20653;
wire S20654;
wire S20655;
wire S20656;
wire S20657;
wire S20658;
wire S20659;
wire S20660;
wire S20661;
wire S20662;
wire S20663;
wire S20664;
wire S20665;
wire S20666;
wire S20667;
wire S20668;
wire S20669;
wire S20670;
wire S20671;
wire S20672;
wire S20673;
wire S20674;
wire S20675;
wire S20676;
wire S20677;
wire S20678;
wire S20679;
wire S20680;
wire S20681;
wire S20682;
wire S20683;
wire S20684;
wire S20685;
wire S20686;
wire S20687;
wire S20688;
wire S20689;
wire S20690;
wire S20691;
wire S20692;
wire S20693;
wire S20694;
wire S20695;
wire S20696;
wire S20697;
wire S20698;
wire S20699;
wire S20700;
wire S20701;
wire S20702;
wire S20703;
wire S20704;
wire S20705;
wire S20706;
wire S20707;
wire S20708;
wire S20709;
wire S20710;
wire S20711;
wire S20712;
wire S20713;
wire S20714;
wire S20715;
wire S20716;
wire S20717;
wire S20718;
wire S20719;
wire S20720;
wire S20721;
wire S20722;
wire S20723;
wire S20724;
wire S20725;
wire S20726;
wire S20727;
wire S20728;
wire S20729;
wire S20730;
wire S20731;
wire S20732;
wire S20733;
wire S20734;
wire S20735;
wire S20736;
wire S20737;
wire S20738;
wire S20739;
wire S20740;
wire S20741;
wire S20742;
wire S20743;
wire S20744;
wire S20745;
wire S20746;
wire S20747;
wire S20748;
wire S20749;
wire S20750;
wire S20751;
wire S20752;
wire S20753;
wire S20754;
wire S20755;
wire S20756;
wire S20757;
wire S20758;
wire S20759;
wire S20760;
wire S20761;
wire S20762;
wire S20763;
wire S20764;
wire S20765;
wire S20766;
wire S20767;
wire S20768;
wire S20769;
wire S20770;
wire S20771;
wire S20772;
wire S20773;
wire S20774;
wire S20775;
wire S20776;
wire S20777;
wire S20778;
wire S20779;
wire S20780;
wire S20781;
wire S20782;
wire S20783;
wire S20784;
wire S20785;
wire S20786;
wire S20787;
wire S20788;
wire S20789;
wire S20790;
wire S20791;
wire S20792;
wire S20793;
wire S20794;
wire S20795;
wire S20796;
wire S20797;
wire S20798;
wire S20799;
wire S20800;
wire S20801;
wire S20802;
wire S20803;
wire S20804;
wire S20805;
wire S20806;
wire S20807;
wire S20808;
wire S20809;
wire S20810;
wire S20811;
wire S20812;
wire S20813;
wire S20814;
wire S20815;
wire S20816;
wire S20817;
wire S20818;
wire S20819;
wire S20820;
wire S20821;
wire S20822;
wire S20823;
wire S20824;
wire S20825;
wire S20826;
wire S20827;
wire S20828;
wire S20829;
wire S20830;
wire S20831;
wire S20832;
wire S20833;
wire S20834;
wire S20835;
wire S20836;
wire S20837;
wire S20838;
wire S20839;
wire S20840;
wire S20841;
wire S20842;
wire S20843;
wire S20844;
wire S20845;
wire S20846;
wire S20847;
wire S20848;
wire S20849;
wire S20850;
wire S20851;
wire S20852;
wire S20853;
wire S20854;
wire S20855;
wire S20856;
wire S20857;
wire S20858;
wire S20859;
wire S20860;
wire S20861;
wire S20862;
wire S20863;
wire S20864;
wire S20865;
wire S20866;
wire S20867;
wire S20868;
wire S20869;
wire S20870;
wire S20871;
wire S20872;
wire S20873;
wire S20874;
wire S20875;
wire S20876;
wire S20877;
wire S20878;
wire S20879;
wire S20880;
wire S20881;
wire S20882;
wire S20883;
wire S20884;
wire S20885;
wire S20886;
wire S20887;
wire S20888;
wire S20889;
wire S20890;
wire S20891;
wire S20892;
wire S20893;
wire S20894;
wire S20895;
wire S20896;
wire S20897;
wire S20898;
wire S20899;
wire S20900;
wire S20901;
wire S20902;
wire S20903;
wire S20904;
wire S20905;
wire S20906;
wire S20907;
wire S20908;
wire S20909;
wire S20910;
wire S20911;
wire S20912;
wire S20913;
wire S20914;
wire S20915;
wire S20916;
wire S20917;
wire S20918;
wire S20919;
wire S20920;
wire S20921;
wire S20922;
wire S20923;
wire S20924;
wire S20925;
wire S20926;
wire S20927;
wire S20928;
wire S20929;
wire S20930;
wire S20931;
wire S20932;
wire S20933;
wire S20934;
wire S20935;
wire S20936;
wire S20937;
wire S20938;
wire S20939;
wire S20940;
wire S20941;
wire S20942;
wire S20943;
wire S20944;
wire S20945;
wire S20946;
wire S20947;
wire S20948;
wire S20949;
wire S20950;
wire S20951;
wire S20952;
wire S20953;
wire S20954;
wire S20955;
wire S20956;
wire S20957;
wire S20958;
wire S20959;
wire S20960;
wire S20961;
wire S20962;
wire S20963;
wire S20964;
wire S20965;
wire S20966;
wire S20967;
wire S20968;
wire S20969;
wire S20970;
wire S20971;
wire S20972;
wire S20973;
wire S20974;
wire S20975;
wire S20976;
wire S20977;
wire S20978;
wire S20979;
wire S20980;
wire S20981;
wire S20982;
wire S20983;
wire S20984;
wire S20985;
wire S20986;
wire S20987;
wire S20988;
wire S20989;
wire S20990;
wire S20991;
wire S20992;
wire S20993;
wire S20994;
wire S20995;
wire S20996;
wire S20997;
wire S20998;
wire S20999;
wire S21000;
wire S21001;
wire S21002;
wire S21003;
wire S21004;
wire S21005;
wire S21006;
wire S21007;
wire S21008;
wire S21009;
wire S21010;
wire S21011;
wire S21012;
wire S21013;
wire S21014;
wire S21015;
wire S21016;
wire S21017;
wire S21018;
wire S21019;
wire S21020;
wire S21021;
wire S21022;
wire S21023;
wire S21024;
wire S21025;
wire S21026;
wire S21027;
wire S21028;
wire S21029;
wire S21030;
wire S21031;
wire S21032;
wire S21033;
wire S21034;
wire S21035;
wire S21036;
wire S21037;
wire S21038;
wire S21039;
wire S21040;
wire S21041;
wire S21042;
wire S21043;
wire S21044;
wire S21045;
wire S21046;
wire S21047;
wire S21048;
wire S21049;
wire S21050;
wire S21051;
wire S21052;
wire S21053;
wire S21054;
wire S21055;
wire S21056;
wire S21057;
wire S21058;
wire S21059;
wire S21060;
wire S21061;
wire S21062;
wire S21063;
wire S21064;
wire S21065;
wire S21066;
wire S21067;
wire S21068;
wire S21069;
wire S21070;
wire S21071;
wire S21072;
wire S21073;
wire S21074;
wire S21075;
wire S21076;
wire S21077;
wire S21078;
wire S21079;
wire S21080;
wire S21081;
wire S21082;
wire S21083;
wire S21084;
wire S21085;
wire S21086;
wire S21087;
wire S21088;
wire S21089;
wire S21090;
wire S21091;
wire S21092;
wire S21093;
wire S21094;
wire S21095;
wire S21096;
wire S21097;
wire S21098;
wire S21099;
wire S21100;
wire S21101;
wire S21102;
wire S21103;
wire S21104;
wire S21105;
wire S21106;
wire S21107;
wire S21108;
wire S21109;
wire S21110;
wire S21111;
wire S21112;
wire S21113;
wire S21114;
wire S21115;
wire S21116;
wire S21117;
wire S21118;
wire S21119;
wire S21120;
wire S21121;
wire S21122;
wire S21123;
wire S21124;
wire S21125;
wire S21126;
wire S21127;
wire S21128;
wire S21129;
wire S21130;
wire S21131;
wire S21132;
wire S21133;
wire S21134;
wire S21135;
wire S21136;
wire S21137;
wire S21138;
wire S21139;
wire S21140;
wire S21141;
wire S21142;
wire S21143;
wire S21144;
wire S21145;
wire S21146;
wire S21147;
wire S21148;
wire S21149;
wire S21150;
wire S21151;
wire S21152;
wire S21153;
wire S21154;
wire S21155;
wire S21156;
wire S21157;
wire S21158;
wire S21159;
wire S21160;
wire S21161;
wire S21162;
wire S21163;
wire S21164;
wire S21165;
wire S21166;
wire S21167;
wire S21168;
wire S21169;
wire S21170;
wire S21171;
wire S21172;
wire S21173;
wire S21174;
wire S21175;
wire S21176;
wire S21177;
wire S21178;
wire S21179;
wire S21180;
wire S21181;
wire S21182;
wire S21183;
wire S21184;
wire S21185;
wire S21186;
wire S21187;
wire S21188;
wire S21189;
wire S21190;
wire S21191;
wire S21192;
wire S21193;
wire S21194;
wire S21195;
wire S21196;
wire S21197;
wire S21198;
wire S21199;
wire S21200;
wire S21201;
wire S21202;
wire S21203;
wire S21204;
wire S21205;
wire S21206;
wire S21207;
wire S21208;
wire S21209;
wire S21210;
wire S21211;
wire S21212;
wire S21213;
wire S21214;
wire S21215;
wire S21216;
wire S21217;
wire S21218;
wire S21219;
wire S21220;
wire S21221;
wire S21222;
wire S21223;
wire S21224;
wire S21225;
wire S21226;
wire S21227;
wire S21228;
wire S21229;
wire S21230;
wire S21231;
wire S21232;
wire S21233;
wire S21234;
wire S21235;
wire S21236;
wire S21237;
wire S21238;
wire S21239;
wire S21240;
wire S21241;
wire S21242;
wire S21243;
wire S21244;
wire S21245;
wire S21246;
wire S21247;
wire S21248;
wire S21249;
wire S21250;
wire S21251;
wire S21252;
wire S21253;
wire S21254;
wire S21255;
wire S21256;
wire S21257;
wire S21258;
wire S21259;
wire S21260;
wire S21261;
wire S21262;
wire S21263;
wire S21264;
wire S21265;
wire S21266;
wire S21267;
wire S21268;
wire S21269;
wire S21270;
wire S21271;
wire S21272;
wire S21273;
wire S21274;
wire S21275;
wire S21276;
wire S21277;
wire S21278;
wire S21279;
wire S21280;
wire S21281;
wire S21282;
wire S21283;
wire S21284;
wire S21285;
wire S21286;
wire S21287;
wire S21288;
wire S21289;
wire S21290;
wire S21291;
wire S21292;
wire S21293;
wire S21294;
wire S21295;
wire S21296;
wire S21297;
wire S21298;
wire S21299;
wire S21300;
wire S21301;
wire S21302;
wire S21303;
wire S21304;
wire S21305;
wire S21306;
wire S21307;
wire S21308;
wire S21309;
wire S21310;
wire S21311;
wire S21312;
wire S21313;
wire S21314;
wire S21315;
wire S21316;
wire S21317;
wire S21318;
wire S21319;
wire S21320;
wire S21321;
wire S21322;
wire S21323;
wire S21324;
wire S21325;
wire S21326;
wire S21327;
wire S21328;
wire S21329;
wire S21330;
wire S21331;
wire S21332;
wire S21333;
wire S21334;
wire S21335;
wire S21336;
wire S21337;
wire S21338;
wire S21339;
wire S21340;
wire S21341;
wire S21342;
wire S21343;
wire S21344;
wire S21345;
wire S21346;
wire S21347;
wire S21348;
wire S21349;
wire S21350;
wire S21351;
wire S21352;
wire S21353;
wire S21354;
wire S21355;
wire S21356;
wire S21357;
wire S21358;
wire S21359;
wire S21360;
wire S21361;
wire S21362;
wire S21363;
wire S21364;
wire S21365;
wire S21366;
wire S21367;
wire S21368;
wire S21369;
wire S21370;
wire S21371;
wire S21372;
wire S21373;
wire S21374;
wire S21375;
wire S21376;
wire S21377;
wire S21378;
wire S21379;
wire S21380;
wire S21381;
wire S21382;
wire S21383;
wire S21384;
wire S21385;
wire S21386;
wire S21387;
wire S21388;
wire S21389;
wire S21390;
wire S21391;
wire S21392;
wire S21393;
wire S21394;
wire S21395;
wire S21396;
wire S21397;
wire S21398;
wire S21399;
wire S21400;
wire S21401;
wire S21402;
wire S21403;
wire S21404;
wire S21405;
wire S21406;
wire S21407;
wire S21408;
wire S21409;
wire S21410;
wire S21411;
wire S21412;
wire S21413;
wire S21414;
wire S21415;
wire S21416;
wire S21417;
wire S21418;
wire S21419;
wire S21420;
wire S21421;
wire S21422;
wire S21423;
wire S21424;
wire S21425;
wire S21426;
wire S21427;
wire S21428;
wire S21429;
wire S21430;
wire S21431;
wire S21432;
wire S21433;
wire S21434;
wire S21435;
wire S21436;
wire S21437;
wire S21438;
wire S21439;
wire S21440;
wire S21441;
wire S21442;
wire S21443;
wire S21444;
wire S21445;
wire S21446;
wire S21447;
wire S21448;
wire S21449;
wire S21450;
wire S21451;
wire S21452;
wire S21453;
wire S21454;
wire S21455;
wire S21456;
wire S21457;
wire S21458;
wire S21459;
wire S21460;
wire S21461;
wire S21462;
wire S21463;
wire S21464;
wire S21465;
wire S21466;
wire S21467;
wire S21468;
wire S21469;
wire S21470;
wire S21471;
wire S21472;
wire S21473;
wire S21474;
wire S21475;
wire S21476;
wire S21477;
wire S21478;
wire S21479;
wire S21480;
wire S21481;
wire S21482;
wire S21483;
wire S21484;
wire S21485;
wire S21486;
wire S21487;
wire S21488;
wire S21489;
wire S21490;
wire S21491;
wire S21492;
wire S21493;
wire S21494;
wire S21495;
wire S21496;
wire S21497;
wire S21498;
wire S21499;
wire S21500;
wire S21501;
wire S21502;
wire S21503;
wire S21504;
wire S21505;
wire S21506;
wire S21507;
wire S21508;
wire S21509;
wire S21510;
wire S21511;
wire S21512;
wire S21513;
wire S21514;
wire S21515;
wire S21516;
wire S21517;
wire S21518;
wire S21519;
wire S21520;
wire S21521;
wire S21522;
wire S21523;
wire S21524;
wire S21525;
wire S21526;
wire S21527;
wire S21528;
wire S21529;
wire S21530;
wire S21531;
wire S21532;
wire S21533;
wire S21534;
wire S21535;
wire S21536;
wire S21537;
wire S21538;
wire S21539;
wire S21540;
wire S21541;
wire S21542;
wire S21543;
wire S21544;
wire S21545;
wire S21546;
wire S21547;
wire S21548;
wire S21549;
wire S21550;
wire S21551;
wire S21552;
wire S21553;
wire S21554;
wire S21555;
wire S21556;
wire S21557;
wire S21558;
wire S21559;
wire S21560;
wire S21561;
wire S21562;
wire S21563;
wire S21564;
wire S21565;
wire S21566;
wire S21567;
wire S21568;
wire S21569;
wire S21570;
wire S21571;
wire S21572;
wire S21573;
wire S21574;
wire S21575;
wire S21576;
wire S21577;
wire S21578;
wire S21579;
wire S21580;
wire S21581;
wire S21582;
wire S21583;
wire S21584;
wire S21585;
wire S21586;
wire S21587;
wire S21588;
wire S21589;
wire S21590;
wire S21591;
wire S21592;
wire S21593;
wire S21594;
wire S21595;
wire S21596;
wire S21597;
wire S21598;
wire S21599;
wire S21600;
wire S21601;
wire S21602;
wire S21603;
wire S21604;
wire S21605;
wire S21606;
wire S21607;
wire S21608;
wire S21609;
wire S21610;
wire S21611;
wire S21612;
wire S21613;
wire S21614;
wire S21615;
wire S21616;
wire S21617;
wire S21618;
wire S21619;
wire S21620;
wire S21621;
wire S21622;
wire S21623;
wire S21624;
wire S21625;
wire S21626;
wire S21627;
wire S21628;
wire S21629;
wire S21630;
wire S21631;
wire S21632;
wire S21633;
wire S21634;
wire S21635;
wire S21636;
wire S21637;
wire S21638;
wire S21639;
wire S21640;
wire S21641;
wire S21642;
wire S21643;
wire S21644;
wire S21645;
wire S21646;
wire S21647;
wire S21648;
wire S21649;
wire S21650;
wire S21651;
wire S21652;
wire S21653;
wire S21654;
wire S21655;
wire S21656;
wire S21657;
wire S21658;
wire S21659;
wire S21660;
wire S21661;
wire S21662;
wire S21663;
wire S21664;
wire S21665;
wire S21666;
wire S21667;
wire S21668;
wire S21669;
wire S21670;
wire S21671;
wire S21672;
wire S21673;
wire S21674;
wire S21675;
wire S21676;
wire S21677;
wire S21678;
wire S21679;
wire S21680;
wire S21681;
wire S21682;
wire S21683;
wire S21684;
wire S21685;
wire S21686;
wire S21687;
wire S21688;
wire S21689;
wire S21690;
wire S21691;
wire S21692;
wire S21693;
wire S21694;
wire S21695;
wire S21696;
wire S21697;
wire S21698;
wire S21699;
wire S21700;
wire S21701;
wire S21702;
wire S21703;
wire S21704;
wire S21705;
wire S21706;
wire S21707;
wire S21708;
wire S21709;
wire S21710;
wire S21711;
wire S21712;
wire S21713;
wire S21714;
wire S21715;
wire S21716;
wire S21717;
wire S21718;
wire S21719;
wire S21720;
wire S21721;
wire S21722;
wire S21723;
wire S21724;
wire S21725;
wire S21726;
wire S21727;
wire S21728;
wire S21729;
wire S21730;
wire S21731;
wire S21732;
wire S21733;
wire S21734;
wire S21735;
wire S21736;
wire S21737;
wire S21738;
wire S21739;
wire S21740;
wire S21741;
wire S21742;
wire S21743;
wire S21744;
wire S21745;
wire S21746;
wire S21747;
wire S21748;
wire S21749;
wire S21750;
wire S21751;
wire S21752;
wire S21753;
wire S21754;
wire S21755;
wire S21756;
wire S21757;
wire S21758;
wire S21759;
wire S21760;
wire S21761;
wire S21762;
wire S21763;
wire S21764;
wire S21765;
wire S21766;
wire S21767;
wire S21768;
wire S21769;
wire S21770;
wire S21771;
wire S21772;
wire S21773;
wire S21774;
wire S21775;
wire S21776;
wire S21777;
wire S21778;
wire S21779;
wire S21780;
wire S21781;
wire S21782;
wire S21783;
wire S21784;
wire S21785;
wire S21786;
wire S21787;
wire S21788;
wire S21789;
wire S21790;
wire S21791;
wire S21792;
wire S21793;
wire S21794;
wire S21795;
wire S21796;
wire S21797;
wire S21798;
wire S21799;
wire S21800;
wire S21801;
wire S21802;
wire S21803;
wire S21804;
wire S21805;
wire S21806;
wire S21807;
wire S21808;
wire S21809;
wire S21810;
wire S21811;
wire S21812;
wire S21813;
wire S21814;
wire S21815;
wire S21816;
wire S21817;
wire S21818;
wire S21819;
wire S21820;
wire S21821;
wire S21822;
wire S21823;
wire S21824;
wire S21825;
wire S21826;
wire S21827;
wire S21828;
wire S21829;
wire S21830;
wire S21831;
wire S21832;
wire S21833;
wire S21834;
wire S21835;
wire S21836;
wire S21837;
wire S21838;
wire S21839;
wire S21840;
wire S21841;
wire S21842;
wire S21843;
wire S21844;
wire S21845;
wire S21846;
wire S21847;
wire S21848;
wire S21849;
wire S21850;
wire S21851;
wire S21852;
wire S21853;
wire S21854;
wire S21855;
wire S21856;
wire S21857;
wire S21858;
wire S21859;
wire S21860;
wire S21861;
wire S21862;
wire S21863;
wire S21864;
wire S21865;
wire S21866;
wire S21867;
wire S21868;
wire S21869;
wire S21870;
wire S21871;
wire S21872;
wire S21873;
wire S21874;
wire S21875;
wire S21876;
wire S21877;
wire S21878;
wire S21879;
wire S21880;
wire S21881;
wire S21882;
wire S21883;
wire S21884;
wire S21885;
wire S21886;
wire S21887;
wire S21888;
wire S21889;
wire S21890;
wire S21891;
wire S21892;
wire S21893;
wire S21894;
wire S21895;
wire S21896;
wire S21897;
wire S21898;
wire S21899;
wire S21900;
wire S21901;
wire S21902;
wire S21903;
wire S21904;
wire S21905;
wire S21906;
wire S21907;
wire S21908;
wire S21909;
wire S21910;
wire S21911;
wire S21912;
wire S21913;
wire S21914;
wire S21915;
wire S21916;
wire S21917;
wire S21918;
wire S21919;
wire S21920;
wire S21921;
wire S21922;
wire S21923;
wire S21924;
wire S21925;
wire S21926;
wire S21927;
wire S21928;
wire S21929;
wire S21930;
wire S21931;
wire S21932;
wire S21933;
wire S21934;
wire S21935;
wire S21936;
wire S21937;
wire S21938;
wire S21939;
wire S21940;
wire S21941;
wire S21942;
wire S21943;
wire S21944;
wire S21945;
wire S21946;
wire S21947;
wire S21948;
wire S21949;
wire S21950;
wire S21951;
wire S21952;
wire S21953;
wire S21954;
wire S21955;
wire S21956;
wire S21957;
wire S21958;
wire S21959;
wire S21960;
wire S21961;
wire S21962;
wire S21963;
wire S21964;
wire S21965;
wire S21966;
wire S21967;
wire S21968;
wire S21969;
wire S21970;
wire S21971;
wire S21972;
wire S21973;
wire S21974;
wire S21975;
wire S21976;
wire S21977;
wire S21978;
wire S21979;
wire S21980;
wire S21981;
wire S21982;
wire S21983;
wire S21984;
wire S21985;
wire S21986;
wire S21987;
wire S21988;
wire S21989;
wire S21990;
wire S21991;
wire S21992;
wire S21993;
wire S21994;
wire S21995;
wire S21996;
wire S21997;
wire S21998;
wire S21999;
wire S22000;
wire S22001;
wire S22002;
wire S22003;
wire S22004;
wire S22005;
wire S22006;
wire S22007;
wire S22008;
wire S22009;
wire S22010;
wire S22011;
wire S22012;
wire S22013;
wire S22014;
wire S22015;
wire S22016;
wire S22017;
wire S22018;
wire S22019;
wire S22020;
wire S22021;
wire S22022;
wire S22023;
wire S22024;
wire S22025;
wire S22026;
wire S22027;
wire S22028;
wire S22029;
wire S22030;
wire S22031;
wire S22032;
wire S22033;
wire S22034;
wire S22035;
wire S22036;
wire S22037;
wire S22038;
wire S22039;
wire S22040;
wire S22041;
wire S22042;
wire S22043;
wire S22044;
wire S22045;
wire S22046;
wire S22047;
wire S22048;
wire S22049;
wire S22050;
wire S22051;
wire S22052;
wire S22053;
wire S22054;
wire S22055;
wire S22056;
wire S22057;
wire S22058;
wire S22059;
wire S22060;
wire S22061;
wire S22062;
wire S22063;
wire S22064;
wire S22065;
wire S22066;
wire S22067;
wire S22068;
wire S22069;
wire S22070;
wire S22071;
wire S22072;
wire S22073;
wire S22074;
wire S22075;
wire S22076;
wire S22077;
wire S22078;
wire S22079;
wire S22080;
wire S22081;
wire S22082;
wire S22083;
wire S22084;
wire S22085;
wire S22086;
wire S22087;
wire S22088;
wire S22089;
wire S22090;
wire S22091;
wire S22092;
wire S22093;
wire S22094;
wire S22095;
wire S22096;
wire S22097;
wire S22098;
wire S22099;
wire S22100;
wire S22101;
wire S22102;
wire S22103;
wire S22104;
wire S22105;
wire S22106;
wire S22107;
wire S22108;
wire S22109;
wire S22110;
wire S22111;
wire S22112;
wire S22113;
wire S22114;
wire S22115;
wire S22116;
wire S22117;
wire S22118;
wire S22119;
wire S22120;
wire S22121;
wire S22122;
wire S22123;
wire S22124;
wire S22125;
wire S22126;
wire S22127;
wire S22128;
wire S22129;
wire S22130;
wire S22131;
wire S22132;
wire S22133;
wire S22134;
wire S22135;
wire S22136;
wire S22137;
wire S22138;
wire S22139;
wire S22140;
wire S22141;
wire S22142;
wire S22143;
wire S22144;
wire S22145;
wire S22146;
wire S22147;
wire S22148;
wire S22149;
wire S22150;
wire S22151;
wire S22152;
wire S22153;
wire S22154;
wire S22155;
wire S22156;
wire S22157;
wire S22158;
wire S22159;
wire S22160;
wire S22161;
wire S22162;
wire S22163;
wire S22164;
wire S22165;
wire S22166;
wire S22167;
wire S22168;
wire S22169;
wire S22170;
wire S22171;
wire S22172;
wire S22173;
wire S22174;
wire S22175;
wire S22176;
wire S22177;
wire S22178;
wire S22179;
wire S22180;
wire S22181;
wire S22182;
wire S22183;
wire S22184;
wire S22185;
wire S22186;
wire S22187;
wire S22188;
wire S22189;
wire S22190;
wire S22191;
wire S22192;
wire S22193;
wire S22194;
wire S22195;
wire S22196;
wire S22197;
wire S22198;
wire S22199;
wire S22200;
wire S22201;
wire S22202;
wire S22203;
wire S22204;
wire S22205;
wire S22206;
wire S22207;
wire S22208;
wire S22209;
wire S22210;
wire S22211;
wire S22212;
wire S22213;
wire S22214;
wire S22215;
wire S22216;
wire S22217;
wire S22218;
wire S22219;
wire S22220;
wire S22221;
wire S22222;
wire S22223;
wire S22224;
wire S22225;
wire S22226;
wire S22227;
wire S22228;
wire S22229;
wire S22230;
wire S22231;
wire S22232;
wire S22233;
wire S22234;
wire S22235;
wire S22236;
wire S22237;
wire S22238;
wire S22239;
wire S22240;
wire S22241;
wire S22242;
wire S22243;
wire S22244;
wire S22245;
wire S22246;
wire S22247;
wire S22248;
wire S22249;
wire S22250;
wire S22251;
wire S22252;
wire S22253;
wire S22254;
wire S22255;
wire S22256;
wire S22257;
wire S22258;
wire S22259;
wire S22260;
wire S22261;
wire S22262;
wire S22263;
wire S22264;
wire S22265;
wire S22266;
wire S22267;
wire S22268;
wire S22269;
wire S22270;
wire S22271;
wire S22272;
wire S22273;
wire S22274;
wire S22275;
wire S22276;
wire S22277;
wire S22278;
wire S22279;
wire S22280;
wire S22281;
wire S22282;
wire S22283;
wire S22284;
wire S22285;
wire S22286;
wire S22287;
wire S22288;
wire S22289;
wire S22290;
wire S22291;
wire S22292;
wire S22293;
wire S22294;
wire S22295;
wire S22296;
wire S22297;
wire S22298;
wire S22299;
wire S22300;
wire S22301;
wire S22302;
wire S22303;
wire S22304;
wire S22305;
wire S22306;
wire S22307;
wire S22308;
wire S22309;
wire S22310;
wire S22311;
wire S22312;
wire S22313;
wire S22314;
wire S22315;
wire S22316;
wire S22317;
wire S22318;
wire S22319;
wire S22320;
wire S22321;
wire S22322;
wire S22323;
wire S22324;
wire S22325;
wire S22326;
wire S22327;
wire S22328;
wire S22329;
wire S22330;
wire S22331;
wire S22332;
wire S22333;
wire S22334;
wire S22335;
wire S22336;
wire S22337;
wire S22338;
wire S22339;
wire S22340;
wire S22341;
wire S22342;
wire S22343;
wire S22344;
wire S22345;
wire S22346;
wire S22347;
wire S22348;
wire S22349;
wire S22350;
wire S22351;
wire S22352;
wire S22353;
wire S22354;
wire S22355;
wire S22356;
wire S22357;
wire S22358;
wire S22359;
wire S22360;
wire S22361;
wire S22362;
wire S22363;
wire S22364;
wire S22365;
wire S22366;
wire S22367;
wire S22368;
wire S22369;
wire S22370;
wire S22371;
wire S22372;
wire S22373;
wire S22374;
wire S22375;
wire S22376;
wire S22377;
wire S22378;
wire S22379;
wire S22380;
wire S22381;
wire S22382;
wire S22383;
wire S22384;
wire S22385;
wire S22386;
wire S22387;
wire S22388;
wire S22389;
wire S22390;
wire S22391;
wire S22392;
wire S22393;
wire S22394;
wire S22395;
wire S22396;
wire S22397;
wire S22398;
wire S22399;
wire S22400;
wire S22401;
wire S22402;
wire S22403;
wire S22404;
wire S22405;
wire S22406;
wire S22407;
wire S22408;
wire S22409;
wire S22410;
wire S22411;
wire S22412;
wire S22413;
wire S22414;
wire S22415;
wire S22416;
wire S22417;
wire S22418;
wire S22419;
wire S22420;
wire S22421;
wire S22422;
wire S22423;
wire S22424;
wire S22425;
wire S22426;
wire S22427;
wire S22428;
wire S22429;
wire S22430;
wire S22431;
wire S22432;
wire S22433;
wire S22434;
wire S22435;
wire S22436;
wire S22437;
wire S22438;
wire S22439;
wire S22440;
wire S22441;
wire S22442;
wire S22443;
wire S22444;
wire S22445;
wire S22446;
wire S22447;
wire S22448;
wire S22449;
wire S22450;
wire S22451;
wire S22452;
wire S22453;
wire S22454;
wire S22455;
wire S22456;
wire S22457;
wire S22458;
wire S22459;
wire S22460;
wire S22461;
wire S22462;
wire S22463;
wire S22464;
wire S22465;
wire S22466;
wire S22467;
wire S22468;
wire S22469;
wire S22470;
wire S22471;
wire S22472;
wire S22473;
wire S22474;
wire S22475;
wire S22476;
wire S22477;
wire S22478;
wire S22479;
wire S22480;
wire S22481;
wire S22482;
wire S22483;
wire S22484;
wire S22485;
wire S22486;
wire S22487;
wire S22488;
wire S22489;
wire S22490;
wire S22491;
wire S22492;
wire S22493;
wire S22494;
wire S22495;
wire S22496;
wire S22497;
wire S22498;
wire S22499;
wire S22500;
wire S22501;
wire S22502;
wire S22503;
wire S22504;
wire S22505;
wire S22506;
wire S22507;
wire S22508;
wire S22509;
wire S22510;
wire S22511;
wire S22512;
wire S22513;
wire S22514;
wire S22515;
wire S22516;
wire S22517;
wire S22518;
wire S22519;
wire S22520;
wire S22521;
wire S22522;
wire S22523;
wire S22524;
wire S22525;
wire S22526;
wire S22527;
wire S22528;
wire S22529;
wire S22530;
wire S22531;
wire S22532;
wire S22533;
wire S22534;
wire S22535;
wire S22536;
wire S22537;
wire S22538;
wire S22539;
wire S22540;
wire S22541;
wire S22542;
wire S22543;
wire S22544;
wire S22545;
wire S22546;
wire S22547;
wire S22548;
wire S22549;
wire S22550;
wire S22551;
wire S22552;
wire S22553;
wire S22554;
wire S22555;
wire S22556;
wire S22557;
wire S22558;
wire S22559;
wire S22560;
wire S22561;
wire S22562;
wire S22563;
wire S22564;
wire S22565;
wire S22566;
wire S22567;
wire S22568;
wire S22569;
wire S22570;
wire S22571;
wire S22572;
wire S22573;
wire S22574;
wire S22575;
wire S22576;
wire S22577;
wire S22578;
wire S22579;
wire S22580;
wire S22581;
wire S22582;
wire S22583;
wire S22584;
wire S22585;
wire S22586;
wire S22587;
wire S22588;
wire S22589;
wire S22590;
wire S22591;
wire S22592;
wire S22593;
wire S22594;
wire S22595;
wire S22596;
wire S22597;
wire S22598;
wire S22599;
wire S22600;
wire S22601;
wire S22602;
wire S22603;
wire S22604;
wire S22605;
wire S22606;
wire S22607;
wire S22608;
wire S22609;
wire S22610;
wire S22611;
wire S22612;
wire S22613;
wire S22614;
wire S22615;
wire S22616;
wire S22617;
wire S22618;
wire S22619;
wire S22620;
wire S22621;
wire S22622;
wire S22623;
wire S22624;
wire S22625;
wire S22626;
wire S22627;
wire S22628;
wire S22629;
wire S22630;
wire S22631;
wire S22632;
wire S22633;
wire S22634;
wire S22635;
wire S22636;
wire S22637;
wire S22638;
wire S22639;
wire S22640;
wire S22641;
wire S22642;
wire S22643;
wire S22644;
wire S22645;
wire S22646;
wire S22647;
wire S22648;
wire S22649;
wire S22650;
wire S22651;
wire S22652;
wire S22653;
wire S22654;
wire S22655;
wire S22656;
wire S22657;
wire S22658;
wire S22659;
wire S22660;
wire S22661;
wire S22662;
wire S22663;
wire S22664;
wire S22665;
wire S22666;
wire S22667;
wire S22668;
wire S22669;
wire S22670;
wire S22671;
wire S22672;
wire S22673;
wire S22674;
wire S22675;
wire S22676;
wire S22677;
wire S22678;
wire S22679;
wire S22680;
wire S22681;
wire S22682;
wire S22683;
wire S22684;
wire S22685;
wire S22686;
wire S22687;
wire S22688;
wire S22689;
wire S22690;
wire S22691;
wire S22692;
wire S22693;
wire S22694;
wire S22695;
wire S22696;
wire S22697;
wire S22698;
wire S22699;
wire S22700;
wire S22701;
wire S22702;
wire S22703;
wire S22704;
wire S22705;
wire S22706;
wire S22707;
wire S22708;
wire S22709;
wire S22710;
wire S22711;
wire S22712;
wire S22713;
wire S22714;
wire S22715;
wire S22716;
wire S22717;
wire S22718;
wire S22719;
wire S22720;
wire S22721;
wire S22722;
wire S22723;
wire S22724;
wire S22725;
wire S22726;
wire S22727;
wire S22728;
wire S22729;
wire S22730;
wire S22731;
wire S22732;
wire S22733;
wire S22734;
wire S22735;
wire S22736;
wire S22737;
wire S22738;
wire S22739;
wire S22740;
wire S22741;
wire S22742;
wire S22743;
wire S22744;
wire S22745;
wire S22746;
wire S22747;
wire S22748;
wire S22749;
wire S22750;
wire S22751;
wire S22752;
wire S22753;
wire S22754;
wire S22755;
wire S22756;
wire S22757;
wire S22758;
wire S22759;
wire S22760;
wire S22761;
wire S22762;
wire S22763;
wire S22764;
wire S22765;
wire S22766;
wire S22767;
wire S22768;
wire S22769;
wire S22770;
wire S22771;
wire S22772;
wire S22773;
wire S22774;
wire S22775;
wire S22776;
wire S22777;
wire S22778;
wire S22779;
wire S22780;
wire S22781;
wire S22782;
wire S22783;
wire S22784;
wire S22785;
wire S22786;
wire S22787;
wire S22788;
wire S22789;
wire S22790;
wire S22791;
wire S22792;
wire S22793;
wire S22794;
wire S22795;
wire S22796;
wire S22797;
wire S22798;
wire S22799;
wire S22800;
wire S22801;
wire S22802;
wire S22803;
wire S22804;
wire S22805;
wire S22806;
wire S22807;
wire S22808;
wire S22809;
wire S22810;
wire S22811;
wire S22812;
wire S22813;
wire S22814;
wire S22815;
wire S22816;
wire S22817;
wire S22818;
wire S22819;
wire S22820;
wire S22821;
wire S22822;
wire S22823;
wire S22824;
wire S22825;
wire S22826;
wire S22827;
wire S22828;
wire S22829;
wire S22830;
wire S22831;
wire S22832;
wire S22833;
wire S22834;
wire S22835;
wire S22836;
wire S22837;
wire S22838;
wire S22839;
wire S22840;
wire S22841;
wire S22842;
wire S22843;
wire S22844;
wire S22845;
wire S22846;
wire S22847;
wire S22848;
wire S22849;
wire S22850;
wire S22851;
wire S22852;
wire S22853;
wire S22854;
wire S22855;
wire S22856;
wire S22857;
wire S22858;
wire S22859;
wire S22860;
wire S22861;
wire S22862;
wire S22863;
wire S22864;
wire S22865;
wire S22866;
wire S22867;
wire S22868;
wire S22869;
wire S22870;
wire S22871;
wire S22872;
wire S22873;
wire S22874;
wire S22875;
wire S22876;
wire S22877;
wire S22878;
wire S22879;
wire S22880;
wire S22881;
wire S22882;
wire S22883;
wire S22884;
wire S22885;
wire S22886;
wire S22887;
wire S22888;
wire S22889;
wire S22890;
wire S22891;
wire S22892;
wire S22893;
wire S22894;
wire S22895;
wire S22896;
wire S22897;
wire S22898;
wire S22899;
wire S22900;
wire S22901;
wire S22902;
wire S22903;
wire S22904;
wire S22905;
wire S22906;
wire S22907;
wire S22908;
wire S22909;
wire S22910;
wire S22911;
wire S22912;
wire S22913;
wire S22914;
wire S22915;
wire S22916;
wire S22917;
wire S22918;
wire S22919;
wire S22920;
wire S22921;
wire S22922;
wire S22923;
wire S22924;
wire S22925;
wire S22926;
wire S22927;
wire S22928;
wire S22929;
wire S22930;
wire S22931;
wire S22932;
wire S22933;
wire S22934;
wire S22935;
wire S22936;
wire S22937;
wire S22938;
wire S22939;
wire S22940;
wire S22941;
wire S22942;
wire S22943;
wire S22944;
wire S22945;
wire S22946;
wire S22947;
wire S22948;
wire S22949;
wire S22950;
wire S22951;
wire S22952;
wire S22953;
wire S22954;
wire S22955;
wire S22956;
wire S22957;
wire S22958;
wire S22959;
wire S22960;
wire S22961;
wire S22962;
wire S22963;
wire S22964;
wire S22965;
wire S22966;
wire S22967;
wire S22968;
wire S22969;
wire S22970;
wire S22971;
wire S22972;
wire S22973;
wire S22974;
wire S22975;
wire S22976;
wire S22977;
wire S22978;
wire S22979;
wire S22980;
wire S22981;
wire S22982;
wire S22983;
wire S22984;
wire S22985;
wire S22986;
wire S22987;
wire S22988;
wire S22989;
wire S22990;
wire S22991;
wire S22992;
wire S22993;
wire S22994;
wire S22995;
wire S22996;
wire S22997;
wire S22998;
wire S22999;
wire S23000;
wire S23001;
wire S23002;
wire S23003;
wire S23004;
wire S23005;
wire S23006;
wire S23007;
wire S23008;
wire S23009;
wire S23010;
wire S23011;
wire S23012;
wire S23013;
wire S23014;
wire S23015;
wire S23016;
wire S23017;
wire S23018;
wire S23019;
wire S23020;
wire S23021;
wire S23022;
wire S23023;
wire S23024;
wire S23025;
wire S23026;
wire S23027;
wire S23028;
wire S23029;
wire S23030;
wire S23031;
wire S23032;
wire S23033;
wire S23034;
wire S23035;
wire S23036;
wire S23037;
wire S23038;
wire S23039;
wire S23040;
wire S23041;
wire S23042;
wire S23043;
wire S23044;
wire S23045;
wire S23046;
wire S23047;
wire S23048;
wire S23049;
wire S23050;
wire S23051;
wire S23052;
wire S23053;
wire S23054;
wire S23055;
wire S23056;
wire S23057;
wire S23058;
wire S23059;
wire S23060;
wire S23061;
wire S23062;
wire S23063;
wire S23064;
wire S23065;
wire S23066;
wire S23067;
wire S23068;
wire S23069;
wire S23070;
wire S23071;
wire S23072;
wire S23073;
wire S23074;
wire S23075;
wire S23076;
wire S23077;
wire S23078;
wire S23079;
wire S23080;
wire S23081;
wire S23082;
wire S23083;
wire S23084;
wire S23085;
wire S23086;
wire S23087;
wire S23088;
wire S23089;
wire S23090;
wire S23091;
wire S23092;
wire S23093;
wire S23094;
wire S23095;
wire S23096;
wire S23097;
wire S23098;
wire S23099;
wire S23100;
wire S23101;
wire S23102;
wire S23103;
wire S23104;
wire S23105;
wire S23106;
wire S23107;
wire S23108;
wire S23109;
wire S23110;
wire S23111;
wire S23112;
wire S23113;
wire S23114;
wire S23115;
wire S23116;
wire S23117;
wire S23118;
wire S23119;
wire S23120;
wire S23121;
wire S23122;
wire S23123;
wire S23124;
wire S23125;
wire S23126;
wire S23127;
wire S23128;
wire S23129;
wire S23130;
wire S23131;
wire S23132;
wire S23133;
wire S23134;
wire S23135;
wire S23136;
wire S23137;
wire S23138;
wire S23139;
wire S23140;
wire S23141;
wire S23142;
wire S23143;
wire S23144;
wire S23145;
wire S23146;
wire S23147;
wire S23148;
wire S23149;
wire S23150;
wire S23151;
wire S23152;
wire S23153;
wire S23154;
wire S23155;
wire S23156;
wire S23157;
wire S23158;
wire S23159;
wire S23160;
wire S23161;
wire S23162;
wire S23163;
wire S23164;
wire S23165;
wire S23166;
wire S23167;
wire S23168;
wire S23169;
wire S23170;
wire S23171;
wire S23172;
wire S23173;
wire S23174;
wire S23175;
wire S23176;
wire S23177;
wire S23178;
wire S23179;
wire S23180;
wire S23181;
wire S23182;
wire S23183;
wire S23184;
wire S23185;
wire S23186;
wire S23187;
wire S23188;
wire S23189;
wire S23190;
wire S23191;
wire S23192;
wire S23193;
wire S23194;
wire S23195;
wire S23196;
wire S23197;
wire S23198;
wire S23199;
wire S23200;
wire S23201;
wire S23202;
wire S23203;
wire S23204;
wire S23205;
wire S23206;
wire S23207;
wire S23208;
wire S23209;
wire S23210;
wire S23211;
wire S23212;
wire S23213;
wire S23214;
wire S23215;
wire S23216;
wire S23217;
wire S23218;
wire S23219;
wire S23220;
wire S23221;
wire S23222;
wire S23223;
wire S23224;
wire S23225;
wire S23226;
wire S23227;
wire S23228;
wire S23229;
wire S23230;
wire S23231;
wire S23232;
wire S23233;
wire S23234;
wire S23235;
wire S23236;
wire S23237;
wire S23238;
wire S23239;
wire S23240;
wire S23241;
wire S23242;
wire S23243;
wire S23244;
wire S23245;
wire S23246;
wire S23247;
wire S23248;
wire S23249;
wire S23250;
wire S23251;
wire S23252;
wire S23253;
wire S23254;
wire S23255;
wire S23256;
wire S23257;
wire S23258;
wire S23259;
wire S23260;
wire S23261;
wire S23262;
wire S23263;
wire S23264;
wire S23265;
wire S23266;
wire S23267;
wire S23268;
wire S23269;
wire S23270;
wire S23271;
wire S23272;
wire S23273;
wire S23274;
wire S23275;
wire S23276;
wire S23277;
wire S23278;
wire S23279;
wire S23280;
wire S23281;
wire S23282;
wire S23283;
wire S23284;
wire S23285;
wire S23286;
wire S23287;
wire S23288;
wire S23289;
wire S23290;
wire S23291;
wire S23292;
wire S23293;
wire S23294;
wire S23295;
wire S23296;
wire S23297;
wire S23298;
wire S23299;
wire S23300;
wire S23301;
wire S23302;
wire S23303;
wire S23304;
wire S23305;
wire S23306;
wire S23307;
wire S23308;
wire S23309;
wire S23310;
wire S23311;
wire S23312;
wire S23313;
wire S23314;
wire S23315;
wire S23316;
wire S23317;
wire S23318;
wire S23319;
wire S23320;
wire S23321;
wire S23322;
wire S23323;
wire S23324;
wire S23325;
wire S23326;
wire S23327;
wire S23328;
wire S23329;
wire S23330;
wire S23331;
wire S23332;
wire S23333;
wire S23334;
wire S23335;
wire S23336;
wire S23337;
wire S23338;
wire S23339;
wire S23340;
wire S23341;
wire S23342;
wire S23343;
wire S23344;
wire S23345;
wire S23346;
wire S23347;
wire S23348;
wire S23349;
wire S23350;
wire S23351;
wire S23352;
wire S23353;
wire S23354;
wire S23355;
wire S23356;
wire S23357;
wire S23358;
wire S23359;
wire S23360;
wire S23361;
wire S23362;
wire S23363;
wire S23364;
wire S23365;
wire S23366;
wire S23367;
wire S23368;
wire S23369;
wire S23370;
wire S23371;
wire S23372;
wire S23373;
wire S23374;
wire S23375;
wire S23376;
wire S23377;
wire S23378;
wire S23379;
wire S23380;
wire S23381;
wire S23382;
wire S23383;
wire S23384;
wire S23385;
wire S23386;
wire S23387;
wire S23388;
wire S23389;
wire S23390;
wire S23391;
wire S23392;
wire S23393;
wire S23394;
wire S23395;
wire S23396;
wire S23397;
wire S23398;
wire S23399;
wire S23400;
wire S23401;
wire S23402;
wire S23403;
wire S23404;
wire S23405;
wire S23406;
wire S23407;
wire S23408;
wire S23409;
wire S23410;
wire S23411;
wire S23412;
wire S23413;
wire S23414;
wire S23415;
wire S23416;
wire S23417;
wire S23418;
wire S23419;
wire S23420;
wire S23421;
wire S23422;
wire S23423;
wire S23424;
wire S23425;
wire S23426;
wire S23427;
wire S23428;
wire S23429;
wire S23430;
wire S23431;
wire S23432;
wire S23433;
wire S23434;
wire S23435;
wire S23436;
wire S23437;
wire S23438;
wire S23439;
wire S23440;
wire S23441;
wire S23442;
wire S23443;
wire S23444;
wire S23445;
wire S23446;
wire S23447;
wire S23448;
wire S23449;
wire S23450;
wire S23451;
wire S23452;
wire S23453;
wire S23454;
wire S23455;
wire S23456;
wire S23457;
wire S23458;
wire S23459;
wire S23460;
wire S23461;
wire S23462;
wire S23463;
wire S23464;
wire S23465;
wire S23466;
wire S23467;
wire S23468;
wire S23469;
wire S23470;
wire S23471;
wire S23472;
wire S23473;
wire S23474;
wire S23475;
wire S23476;
wire S23477;
wire S23478;
wire S23479;
wire S23480;
wire S23481;
wire S23482;
wire S23483;
wire S23484;
wire S23485;
wire S23486;
wire S23487;
wire S23488;
wire S23489;
wire S23490;
wire S23491;
wire S23492;
wire S23493;
wire S23494;
wire S23495;
wire S23496;
wire S23497;
wire S23498;
wire S23499;
wire S23500;
wire S23501;
wire S23502;
wire S23503;
wire S23504;
wire S23505;
wire S23506;
wire S23507;
wire S23508;
wire S23509;
wire S23510;
wire S23511;
wire S23512;
wire S23513;
wire S23514;
wire S23515;
wire S23516;
wire S23517;
wire S23518;
wire S23519;
wire S23520;
wire S23521;
wire S23522;
wire S23523;
wire S23524;
wire S23525;
wire S23526;
wire S23527;
wire S23528;
wire S23529;
wire S23530;
wire S23531;
wire S23532;
wire S23533;
wire S23534;
wire S23535;
wire S23536;
wire S23537;
wire S23538;
wire S23539;
wire S23540;
wire S23541;
wire S23542;
wire S23543;
wire S23544;
wire S23545;
wire S23546;
wire S23547;
wire S23548;
wire S23549;
wire S23550;
wire S23551;
wire S23552;
wire S23553;
wire S23554;
wire S23555;
wire S23556;
wire S23557;
wire S23558;
wire S23559;
wire S23560;
wire S23561;
wire S23562;
wire S23563;
wire S23564;
wire S23565;
wire S23566;
wire S23567;
wire S23568;
wire S23569;
wire S23570;
wire S23571;
wire S23572;
wire S23573;
wire S23574;
wire S23575;
wire S23576;
wire S23577;
wire S23578;
wire S23579;
wire S23580;
wire S23581;
wire S23582;
wire S23583;
wire S23584;
wire S23585;
wire S23586;
wire S23587;
wire S23588;
wire S23589;
wire S23590;
wire S23591;
wire S23592;
wire S23593;
wire S23594;
wire S23595;
wire S23596;
wire S23597;
wire S23598;
wire S23599;
wire S23600;
wire S23601;
wire S23602;
wire S23603;
wire S23604;
wire S23605;
wire S23606;
wire S23607;
wire S23608;
wire S23609;
wire S23610;
wire S23611;
wire S23612;
wire S23613;
wire S23614;
wire S23615;
wire S23616;
wire S23617;
wire S23618;
wire S23619;
wire S23620;
wire S23621;
wire S23622;
wire S23623;
wire S23624;
wire S23625;
wire S23626;
wire S23627;
wire S23628;
wire S23629;
wire S23630;
wire S23631;
wire S23632;
wire S23633;
wire S23634;
wire S23635;
wire S23636;
wire S23637;
wire S23638;
wire S23639;
wire S23640;
wire S23641;
wire S23642;
wire S23643;
wire S23644;
wire S23645;
wire S23646;
wire S23647;
wire S23648;
wire S23649;
wire S23650;
wire S23651;
wire S23652;
wire S23653;
wire S23654;
wire S23655;
wire S23656;
wire S23657;
wire S23658;
wire S23659;
wire S23660;
wire S23661;
wire S23662;
wire S23663;
wire S23664;
wire S23665;
wire S23666;
wire S23667;
wire S23668;
wire S23669;
wire S23670;
wire S23671;
wire S23672;
wire S23673;
wire S23674;
wire S23675;
wire S23676;
wire S23677;
wire S23678;
wire S23679;
wire S23680;
wire S23681;
wire S23682;
wire S23683;
wire S23684;
wire S23685;
wire S23686;
wire S23687;
wire S23688;
wire S23689;
wire S23690;
wire S23691;
wire S23692;
wire S23693;
wire S23694;
wire S23695;
wire S23696;
wire S23697;
wire S23698;
wire S23699;
wire S23700;
wire S23701;
wire S23702;
wire S23703;
wire S23704;
wire S23705;
wire S23706;
wire S23707;
wire S23708;
wire S23709;
wire S23710;
wire S23711;
wire S23712;
wire S23713;
wire S23714;
wire S23715;
wire S23716;
wire S23717;
wire S23718;
wire S23719;
wire S23720;
wire S23721;
wire S23722;
wire S23723;
wire S23724;
wire S23725;
wire S23726;
wire S23727;
wire S23728;
wire S23729;
wire S23730;
wire S23731;
wire S23732;
wire S23733;
wire S23734;
wire S23735;
wire S23736;
wire S23737;
wire S23738;
wire S23739;
wire S23740;
wire S23741;
wire S23742;
wire S23743;
wire S23744;
wire S23745;
wire S23746;
wire S23747;
wire S23748;
wire S23749;
wire S23750;
wire S23751;
wire S23752;
wire S23753;
wire S23754;
wire S23755;
wire S23756;
wire S23757;
wire S23758;
wire S23759;
wire S23760;
wire S23761;
wire S23762;
wire S23763;
wire S23764;
wire S23765;
wire S23766;
wire S23767;
wire S23768;
wire S23769;
wire S23770;
wire S23771;
wire S23772;
wire S23773;
wire S23774;
wire S23775;
wire S23776;
wire S23777;
wire S23778;
wire S23779;
wire S23780;
wire S23781;
wire S23782;
wire S23783;
wire S23784;
wire S23785;
wire S23786;
wire S23787;
wire S23788;
wire S23789;
wire S23790;
wire S23791;
wire S23792;
wire S23793;
wire S23794;
wire S23795;
wire S23796;
wire S23797;
wire S23798;
wire S23799;
wire S23800;
wire S23801;
wire S23802;
wire S23803;
wire S23804;
wire S23805;
wire S23806;
wire S23807;
wire S23808;
wire S23809;
wire S23810;
wire S23811;
wire S23812;
wire S23813;
wire S23814;
wire S23815;
wire S23816;
wire S23817;
wire S23818;
wire S23819;
wire S23820;
wire S23821;
wire S23822;
wire S23823;
wire S23824;
wire S23825;
wire S23826;
wire S23827;
wire S23828;
wire S23829;
wire S23830;
wire S23831;
wire S23832;
wire S23833;
wire S23834;
wire S23835;
wire S23836;
wire S23837;
wire S23838;
wire S23839;
wire S23840;
wire S23841;
wire S23842;
wire S23843;
wire S23844;
wire S23845;
wire S23846;
wire S23847;
wire S23848;
wire S23849;
wire S23850;
wire S23851;
wire S23852;
wire S23853;
wire S23854;
wire S23855;
wire S23856;
wire S23857;
wire S23858;
wire S23859;
wire S23860;
wire S23861;
wire S23862;
wire S23863;
wire S23864;
wire S23865;
wire S23866;
wire S23867;
wire S23868;
wire S23869;
wire S23870;
wire S23871;
wire S23872;
wire S23873;
wire S23874;
wire S23875;
wire S23876;
wire S23877;
wire S23878;
wire S23879;
wire S23880;
wire S23881;
wire S23882;
wire S23883;
wire S23884;
wire S23885;
wire S23886;
wire S23887;
wire S23888;
wire S23889;
wire S23890;
wire S23891;
wire S23892;
wire S23893;
wire S23894;
wire S23895;
wire S23896;
wire S23897;
wire S23898;
wire S23899;
wire S23900;
wire S23901;
wire S23902;
wire S23903;
wire S23904;
wire S23905;
wire S23906;
wire S23907;
wire S23908;
wire S23909;
wire S23910;
wire S23911;
wire S23912;
wire S23913;
wire S23914;
wire S23915;
wire S23916;
wire S23917;
wire S23918;
wire S23919;
wire S23920;
wire S23921;
wire S23922;
wire S23923;
wire S23924;
wire S23925;
wire S23926;
wire S23927;
wire S23928;
wire S23929;
wire S23930;
wire S23931;
wire S23932;
wire S23933;
wire S23934;
wire S23935;
wire S23936;
wire S23937;
wire S23938;
wire S23939;
wire S23940;
wire S23941;
wire S23942;
wire S23943;
wire S23944;
wire S23945;
wire S23946;
wire S23947;
wire S23948;
wire S23949;
wire S23950;
wire S23951;
wire S23952;
wire S23953;
wire S23954;
wire S23955;
wire S23956;
wire S23957;
wire S23958;
wire S23959;
wire S23960;
wire S23961;
wire S23962;
wire S23963;
wire S23964;
wire S23965;
wire S23966;
wire S23967;
wire S23968;
wire S23969;
wire S23970;
wire S23971;
wire S23972;
wire S23973;
wire S23974;
wire S23975;
wire S23976;
wire S23977;
wire S23978;
wire S23979;
wire S23980;
wire S23981;
wire S23982;
wire S23983;
wire S23984;
wire S23985;
wire S23986;
wire S23987;
wire S23988;
wire S23989;
wire S23990;
wire S23991;
wire S23992;
wire S23993;
wire S23994;
wire S23995;
wire S23996;
wire S23997;
wire S23998;
wire S23999;
wire S24000;
wire S24001;
wire S24002;
wire S24003;
wire S24004;
wire S24005;
wire S24006;
wire S24007;
wire S24008;
wire S24009;
wire S24010;
wire S24011;
wire S24012;
wire S24013;
wire S24014;
wire S24015;
wire S24016;
wire S24017;
wire S24018;
wire S24019;
wire S24020;
wire S24021;
wire S24022;
wire S24023;
wire S24024;
wire S24025;
wire S24026;
wire S24027;
wire S24028;
wire S24029;
wire S24030;
wire S24031;
wire S24032;
wire S24033;
wire S24034;
wire S24035;
wire S24036;
wire S24037;
wire S24038;
wire S24039;
wire S24040;
wire S24041;
wire S24042;
wire S24043;
wire S24044;
wire S24045;
wire S24046;
wire S24047;
wire S24048;
wire S24049;
wire S24050;
wire S24051;
wire S24052;
wire S24053;
wire S24054;
wire S24055;
wire S24056;
wire S24057;
wire S24058;
wire S24059;
wire S24060;
wire S24061;
wire S24062;
wire S24063;
wire S24064;
wire S24065;
wire S24066;
wire S24067;
wire S24068;
wire S24069;
wire S24070;
wire S24071;
wire S24072;
wire S24073;
wire S24074;
wire S24075;
wire S24076;
wire S24077;
wire S24078;
wire S24079;
wire S24080;
wire S24081;
wire S24082;
wire S24083;
wire S24084;
wire S24085;
wire S24086;
wire S24087;
wire S24088;
wire S24089;
wire S24090;
wire S24091;
wire S24092;
wire S24093;
wire S24094;
wire S24095;
wire S24096;
wire S24097;
wire S24098;
wire S24099;
wire S24100;
wire S24101;
wire S24102;
wire S24103;
wire S24104;
wire S24105;
wire S24106;
wire S24107;
wire S24108;
wire S24109;
wire S24110;
wire S24111;
wire S24112;
wire S24113;
wire S24114;
wire S24115;
wire S24116;
wire S24117;
wire S24118;
wire S24119;
wire S24120;
wire S24121;
wire S24122;
wire S24123;
wire S24124;
wire S24125;
wire S24126;
wire S24127;
wire S24128;
wire S24129;
wire S24130;
wire S24131;
wire S24132;
wire S24133;
wire S24134;
wire S24135;
wire S24136;
wire S24137;
wire S24138;
wire S24139;
wire S24140;
wire S24141;
wire S24142;
wire S24143;
wire S24144;
wire S24145;
wire S24146;
wire S24147;
wire S24148;
wire S24149;
wire S24150;
wire S24151;
wire S24152;
wire S24153;
wire S24154;
wire S24155;
wire S24156;
wire S24157;
wire S24158;
wire S24159;
wire S24160;
wire S24161;
wire S24162;
wire S24163;
wire S24164;
wire S24165;
wire S24166;
wire S24167;
wire S24168;
wire S24169;
wire S24170;
wire S24171;
wire S24172;
wire S24173;
wire S24174;
wire S24175;
wire S24176;
wire S24177;
wire S24178;
wire S24179;
wire S24180;
wire S24181;
wire S24182;
wire S24183;
wire S24184;
wire S24185;
wire S24186;
wire S24187;
wire S24188;
wire S24189;
wire S24190;
wire S24191;
wire S24192;
wire S24193;
wire S24194;
wire S24195;
wire S24196;
wire S24197;
wire S24198;
wire S24199;
wire S24200;
wire S24201;
wire S24202;
wire S24203;
wire S24204;
wire S24205;
wire S24206;
wire S24207;
wire S24208;
wire S24209;
wire S24210;
wire S24211;
wire S24212;
wire S24213;
wire S24214;
wire S24215;
wire S24216;
wire S24217;
wire S24218;
wire S24219;
wire S24220;
wire S24221;
wire S24222;
wire S24223;
wire S24224;
wire S24225;
wire S24226;
wire S24227;
wire S24228;
wire S24229;
wire S24230;
wire S24231;
wire S24232;
wire S24233;
wire S24234;
wire S24235;
wire S24236;
wire S24237;
wire S24238;
wire S24239;
wire S24240;
wire S24241;
wire S24242;
wire S24243;
wire S24244;
wire S24245;
wire S24246;
wire S24247;
wire S24248;
wire S24249;
wire S24250;
wire S24251;
wire S24252;
wire S24253;
wire S24254;
wire S24255;
wire S24256;
wire S24257;
wire S24258;
wire S24259;
wire S24260;
wire S24261;
wire S24262;
wire S24263;
wire S24264;
wire S24265;
wire S24266;
wire S24267;
wire S24268;
wire S24269;
wire S24270;
wire S24271;
wire S24272;
wire S24273;
wire S24274;
wire S24275;
wire S24276;
wire S24277;
wire S24278;
wire S24279;
wire S24280;
wire S24281;
wire S24282;
wire S24283;
wire S24284;
wire S24285;
wire S24286;
wire S24287;
wire S24288;
wire S24289;
wire S24290;
wire S24291;
wire S24292;
wire S24293;
wire S24294;
wire S24295;
wire S24296;
wire S24297;
wire S24298;
wire S24299;
wire S24300;
wire S24301;
wire S24302;
wire S24303;
wire S24304;
wire S24305;
wire S24306;
wire S24307;
wire S24308;
wire S24309;
wire S24310;
wire S24311;
wire S24312;
wire S24313;
wire S24314;
wire S24315;
wire S24316;
wire S24317;
wire S24318;
wire S24319;
wire S24320;
wire S24321;
wire S24322;
wire S24323;
wire S24324;
wire S24325;
wire S24326;
wire S24327;
wire S24328;
wire S24329;
wire S24330;
wire S24331;
wire S24332;
wire S24333;
wire S24334;
wire S24335;
wire S24336;
wire S24337;
wire S24338;
wire S24339;
wire S24340;
wire S24341;
wire S24342;
wire S24343;
wire S24344;
wire S24345;
wire S24346;
wire S24347;
wire S24348;
wire S24349;
wire S24350;
wire S24351;
wire S24352;
wire S24353;
wire S24354;
wire S24355;
wire S24356;
wire S24357;
wire S24358;
wire S24359;
wire S24360;
wire S24361;
wire S24362;
wire S24363;
wire S24364;
wire S24365;
wire S24366;
wire S24367;
wire S24368;
wire S24369;
wire S24370;
wire S24371;
wire S24372;
wire S24373;
wire S24374;
wire S24375;
wire S24376;
wire S24377;
wire S24378;
wire S24379;
wire S24380;
wire S24381;
wire S24382;
wire S24383;
wire S24384;
wire S24385;
wire S24386;
wire S24387;
wire S24388;
wire S24389;
wire S24390;
wire S24391;
wire S24392;
wire S24393;
wire S24394;
wire S24395;
wire S24396;
wire S24397;
wire S24398;
wire S24399;
wire S24400;
wire S24401;
wire S24402;
wire S24403;
wire S24404;
wire S24405;
wire S24406;
wire S24407;
wire S24408;
wire S24409;
wire S24410;
wire S24411;
wire S24412;
wire S24413;
wire S24414;
wire S24415;
wire S24416;
wire S24417;
wire S24418;
wire S24419;
wire S24420;
wire S24421;
wire S24422;
wire S24423;
wire S24424;
wire S24425;
wire S24426;
wire S24427;
wire S24428;
wire S24429;
wire S24430;
wire S24431;
wire S24432;
wire S24433;
wire S24434;
wire S24435;
wire S24436;
wire S24437;
wire S24438;
wire S24439;
wire S24440;
wire S24441;
wire S24442;
wire S24443;
wire S24444;
wire S24445;
wire S24446;
wire S24447;
wire S24448;
wire S24449;
wire S24450;
wire S24451;
wire S24452;
wire S24453;
wire S24454;
wire S24455;
wire S24456;
wire S24457;
wire S24458;
wire S24459;
wire S24460;
wire S24461;
wire S24462;
wire S24463;
wire S24464;
wire S24465;
wire S24466;
wire S24467;
wire S24468;
wire S24469;
wire S24470;
wire S24471;
wire S24472;
wire S24473;
wire S24474;
wire S24475;
wire S24476;
wire S24477;
wire S24478;
wire S24479;
wire S24480;
wire S24481;
wire S24482;
wire S24483;
wire S24484;
wire S24485;
wire S24486;
wire S24487;
wire S24488;
wire S24489;
wire S24490;
wire S24491;
wire S24492;
wire S24493;
wire S24494;
wire S24495;
wire S24496;
wire S24497;
wire S24498;
wire S24499;
wire S24500;
wire S24501;
wire S24502;
wire S24503;
wire S24504;
wire S24505;
wire S24506;
wire S24507;
wire S24508;
wire S24509;
wire S24510;
wire S24511;
wire S24512;
wire S24513;
wire S24514;
wire S24515;
wire S24516;
wire S24517;
wire S24518;
wire S24519;
wire S24520;
wire S24521;
wire S24522;
wire S24523;
wire S24524;
wire S24525;
wire S24526;
wire S24527;
wire S24528;
wire S24529;
wire S24530;
wire S24531;
wire S24532;
wire S24533;
wire S24534;
wire S24535;
wire S24536;
wire S24537;
wire S24538;
wire S24539;
wire S24540;
wire S24541;
wire S24542;
wire S24543;
wire S24544;
wire S24545;
wire S24546;
wire S24547;
wire S24548;
wire S24549;
wire S24550;
wire S24551;
wire S24552;
wire S24553;
wire S24554;
wire S24555;
wire S24556;
wire S24557;
wire S24558;
wire S24559;
wire S24560;
wire S24561;
wire S24562;
wire S24563;
wire S24564;
wire S24565;
wire S24566;
wire S24567;
wire S24568;
wire S24569;
wire S24570;
wire S24571;
wire S24572;
wire S24573;
wire S24574;
wire S24575;
wire S24576;
wire S24577;
wire S24578;
wire S24579;
wire S24580;
wire S24581;
wire S24582;
wire S24583;
wire S24584;
wire S24585;
wire S24586;
wire S24587;
wire S24588;
wire S24589;
wire S24590;
wire S24591;
wire S24592;
wire S24593;
wire S24594;
wire S24595;
wire S24596;
wire S24597;
wire S24598;
wire S24599;
wire S24600;
wire S24601;
wire S24602;
wire S24603;
wire S24604;
wire S24605;
wire S24606;
wire S24607;
wire S24608;
wire S24609;
wire S24610;
wire S24611;
wire S24612;
wire S24613;
wire S24614;
wire S24615;
wire S24616;
wire S24617;
wire S24618;
wire S24619;
wire S24620;
wire S24621;
wire S24622;
wire S24623;
wire S24624;
wire S24625;
wire S24626;
wire S24627;
wire S24628;
wire S24629;
wire S24630;
wire S24631;
wire S24632;
wire S24633;
wire S24634;
wire S24635;
wire S24636;
wire S24637;
wire S24638;
wire S24639;
wire S24640;
wire S24641;
wire S24642;
wire S24643;
wire S24644;
wire S24645;
wire S24646;
wire S24647;
wire S24648;
wire S24649;
wire S24650;
wire S24651;
wire S24652;
wire S24653;
wire S24654;
wire S24655;
wire S24656;
wire S24657;
wire S24658;
wire S24659;
wire S24660;
wire S24661;
wire S24662;
wire S24663;
wire S24664;
wire S24665;
wire S24666;
wire S24667;
wire S24668;
wire S24669;
wire S24670;
wire S24671;
wire S24672;
wire S24673;
wire S24674;
wire S24675;
wire S24676;
wire S24677;
wire S24678;
wire S24679;
wire S24680;
wire S24681;
wire S24682;
wire S24683;
wire S24684;
wire S24685;
wire S24686;
wire S24687;
wire S24688;
wire S24689;
wire S24690;
wire S24691;
wire S24692;
wire S24693;
wire S24694;
wire S24695;
wire S24696;
wire S24697;
wire S24698;
wire S24699;
wire S24700;
wire S24701;
wire S24702;
wire S24703;
wire S24704;
wire S24705;
wire S24706;
wire S24707;
wire S24708;
wire S24709;
wire S24710;
wire S24711;
wire S24712;
wire S24713;
wire S24714;
wire S24715;
wire S24716;
wire S24717;
wire S24718;
wire S24719;
wire S24720;
wire S24721;
wire S24722;
wire S24723;
wire S24724;
wire S24725;
wire S24726;
wire S24727;
wire S24728;
wire S24729;
wire S24730;
wire S24731;
wire S24732;
wire S24733;
wire S24734;
wire S24735;
wire S24736;
wire S24737;
wire S24738;
wire S24739;
wire S24740;
wire S24741;
wire S24742;
wire S24743;
wire S24744;
wire S24745;
wire S24746;
wire S24747;
wire S24748;
wire S24749;
wire S24750;
wire S24751;
wire S24752;
wire S24753;
wire S24754;
wire S24755;
wire S24756;
wire S24757;
wire S24758;
wire S24759;
wire S24760;
wire S24761;
wire S24762;
wire S24763;
wire S24764;
wire S24765;
wire S24766;
wire S24767;
wire S24768;
wire S24769;
wire S24770;
wire S24771;
wire S24772;
wire S24773;
wire S24774;
wire S24775;
wire S24776;
wire S24777;
wire S24778;
wire S24779;
wire S24780;
wire S24781;
wire S24782;
wire S24783;
wire S24784;
wire S24785;
wire S24786;
wire S24787;
wire S24788;
wire S24789;
wire S24790;
wire S24791;
wire S24792;
wire S24793;
wire S24794;
wire S24795;
wire S24796;
wire S24797;
wire S24798;
wire S24799;
wire S24800;
wire S24801;
wire S24802;
wire S24803;
wire S24804;
wire S24805;
wire S24806;
wire S24807;
wire S24808;
wire S24809;
wire S24810;
wire S24811;
wire S24812;
wire S24813;
wire S24814;
wire S24815;
wire S24816;
wire S24817;
wire S24818;
wire S24819;
wire S24820;
wire S24821;
wire S24822;
wire S24823;
wire S24824;
wire S24825;
wire S24826;
wire S24827;
wire S24828;
wire S24829;
wire S24830;
wire S24831;
wire S24832;
wire S24833;
wire S24834;
wire S24835;
wire S24836;
wire S24837;
wire S24838;
wire S24839;
wire S24840;
wire S24841;
wire S24842;
wire S24843;
wire S24844;
wire S24845;
wire S24846;
wire S24847;
wire S24848;
wire S24849;
wire S24850;
wire S24851;
wire S24852;
wire S24853;
wire S24854;
wire S24855;
wire S24856;
wire S24857;
wire S24858;
wire S24859;
wire S24860;
wire S24861;
wire S24862;
wire S24863;
wire S24864;
wire S24865;
wire S24866;
wire S24867;
wire S24868;
wire S24869;
wire S24870;
wire S24871;
wire S24872;
wire S24873;
wire S24874;
wire S24875;
wire S24876;
wire S24877;
wire S24878;
wire S24879;
wire S24880;
wire S24881;
wire S24882;
wire S24883;
wire S24884;
wire S24885;
wire S24886;
wire S24887;
wire S24888;
wire S24889;
wire S24890;
wire S24891;
wire S24892;
wire S24893;
wire S24894;
wire S24895;
wire S24896;
wire S24897;
wire S24898;
wire S24899;
wire S24900;
wire S24901;
wire S24902;
wire S24903;
wire S24904;
wire S24905;
wire S24906;
wire S24907;
wire S24908;
wire S24909;
wire S24910;
wire S24911;
wire S24912;
wire S24913;
wire S24914;
wire S24915;
wire S24916;
wire S24917;
wire S24918;
wire S24919;
wire S24920;
wire S24921;
wire S24922;
wire S24923;
wire S24924;
wire S24925;
wire S24926;
wire S24927;
wire S24928;
wire S24929;
wire S24930;
wire S24931;
wire S24932;
wire S24933;
wire S24934;
wire S24935;
wire S24936;
wire S24937;
wire S24938;
wire S24939;
wire S24940;
wire S24941;
wire S24942;
wire S24943;
wire S24944;
wire S24945;
wire S24946;
wire S24947;
wire S24948;
wire S24949;
wire S24950;
wire S24951;
wire S24952;
wire S24953;
wire S24954;
wire S24955;
wire S24956;
wire S24957;
wire S24958;
wire S24959;
wire S24960;
wire S24961;
wire S24962;
wire S24963;
wire S24964;
wire S24965;
wire S24966;
wire S24967;
wire S24968;
wire S24969;
wire S24970;
wire S24971;
wire S24972;
wire S24973;
wire S24974;
wire S24975;
wire S24976;
wire S24977;
wire S24978;
wire S24979;
wire S24980;
wire S24981;
wire S24982;
wire S24983;
wire S24984;
wire S24985;
wire S24986;
wire S24987;
wire S24988;
wire S24989;
wire S24990;
wire S24991;
wire S24992;
wire S24993;
wire S24994;
wire S24995;
wire S24996;
wire S24997;
wire S24998;
wire S24999;
wire S25000;
wire S25001;
wire S25002;
wire S25003;
wire S25004;
wire S25005;
wire S25006;
wire S25007;
wire S25008;
wire S25009;
wire S25010;
wire S25011;
wire S25012;
wire S25013;
wire S25014;
wire S25015;
wire S25016;
wire S25017;
wire S25018;
wire S25019;
wire S25020;
wire S25021;
wire S25022;
wire S25023;
wire S25024;
wire S25025;
wire S25026;
wire S25027;
wire S25028;
wire S25029;
wire S25030;
wire S25031;
wire S25032;
wire S25033;
wire S25034;
wire S25035;
wire S25036;
wire S25037;
wire S25038;
wire S25039;
wire S25040;
wire S25041;
wire S25042;
wire S25043;
wire S25044;
wire S25045;
wire S25046;
wire S25047;
wire S25048;
wire S25049;
wire S25050;
wire S25051;
wire S25052;
wire S25053;
wire S25054;
wire S25055;
wire S25056;
wire S25057;
wire S25058;
wire S25059;
wire S25060;
wire S25061;
wire S25062;
wire S25063;
wire S25064;
wire S25065;
wire S25066;
wire S25067;
wire S25068;
wire S25069;
wire S25070;
wire S25071;
wire S25072;
wire S25073;
wire S25074;
wire S25075;
wire S25076;
wire S25077;
wire S25078;
wire S25079;
wire S25080;
wire S25081;
wire S25082;
wire S25083;
wire S25084;
wire S25085;
wire S25086;
wire S25087;
wire S25088;
wire S25089;
wire S25090;
wire S25091;
wire S25092;
wire S25093;
wire S25094;
wire S25095;
wire S25096;
wire S25097;
wire S25098;
wire S25099;
wire S25100;
wire S25101;
wire S25102;
wire S25103;
wire S25104;
wire S25105;
wire S25106;
wire S25107;
wire S25108;
wire S25109;
wire S25110;
wire S25111;
wire S25112;
wire S25113;
wire S25114;
wire S25115;
wire S25116;
wire S25117;
wire S25118;
wire S25119;
wire S25120;
wire S25121;
wire S25122;
wire S25123;
wire S25124;
wire S25125;
wire S25126;
wire S25127;
wire S25128;
wire S25129;
wire S25130;
wire S25131;
wire S25132;
wire S25133;
wire S25134;
wire S25135;
wire S25136;
wire S25137;
wire S25138;
wire S25139;
wire S25140;
wire S25141;
wire S25142;
wire S25143;
wire S25144;
wire S25145;
wire S25146;
wire S25147;
wire S25148;
wire S25149;
wire S25150;
wire S25151;
wire S25152;
wire S25153;
wire S25154;
wire S25155;
wire S25156;
wire S25157;
wire S25158;
wire S25159;
wire S25160;
wire S25161;
wire S25162;
wire S25163;
wire S25164;
wire S25165;
wire S25166;
wire S25167;
wire S25168;
wire S25169;
wire S25170;
wire S25171;
wire S25172;
wire S25173;
wire S25174;
wire S25175;
wire S25176;
wire S25177;
wire S25178;
wire S25179;
wire S25180;
wire S25181;
wire S25182;
wire S25183;
wire S25184;
wire S25185;
wire S25186;
wire S25187;
wire S25188;
wire S25189;
wire S25190;
wire S25191;
wire S25192;
wire S25193;
wire S25194;
wire S25195;
wire S25196;
wire S25197;
wire S25198;
wire S25199;
wire S25200;
wire S25201;
wire S25202;
wire S25203;
wire S25204;
wire S25205;
wire S25206;
wire S25207;
wire S25208;
wire S25209;
wire S25210;
wire S25211;
wire S25212;
wire S25213;
wire S25214;
wire S25215;
wire S25216;
wire S25217;
wire S25218;
wire S25219;
wire S25220;
wire S25221;
wire S25222;
wire S25223;
wire S25224;
wire S25225;
wire S25226;
wire S25227;
wire S25228;
wire S25229;
wire S25230;
wire S25231;
wire S25232;
wire S25233;
wire S25234;
wire S25235;
wire S25236;
wire S25237;
wire S25238;
wire S25239;
wire S25240;
wire S25241;
wire S25242;
wire S25243;
wire S25244;
wire S25245;
wire S25246;
wire S25247;
wire S25248;
wire S25249;
wire S25250;
wire S25251;
wire S25252;
wire S25253;
wire S25254;
wire S25255;
wire S25256;
wire S25257;
wire S25258;
wire S25259;
wire S25260;
wire S25261;
wire S25262;
wire S25263;
wire S25264;
wire S25265;
wire S25266;
wire S25267;
wire S25268;
wire S25269;
wire S25270;
wire S25271;
wire S25272;
wire S25273;
wire S25274;
wire S25275;
wire S25276;
wire S25277;
wire S25278;
wire S25279;
wire S25280;
wire S25281;
wire S25282;
wire S25283;
wire S25284;
wire S25285;
wire S25286;
wire S25287;
wire S25288;
wire S25289;
wire S25290;
wire S25291;
wire S25292;
wire S25293;
wire S25294;
wire S25295;
wire S25296;
wire S25297;
wire S25298;
wire S25299;
wire S25300;
wire S25301;
wire S25302;
wire S25303;
wire S25304;
wire S25305;
wire S25306;
wire S25307;
wire S25308;
wire S25309;
wire S25310;
wire S25311;
wire S25312;
wire S25313;
wire S25314;
wire S25315;
wire S25316;
wire S25317;
wire S25318;
wire S25319;
wire S25320;
wire S25321;
wire S25322;
wire S25323;
wire S25324;
wire S25325;
wire S25326;
wire S25327;
wire S25328;
wire S25329;
wire S25330;
wire S25331;
wire S25332;
wire S25333;
wire S25334;
wire S25335;
wire S25336;
wire S25337;
wire S25338;
wire S25339;
wire S25340;
wire S25341;
wire S25342;
wire S25343;
wire S25344;
wire S25345;
wire S25346;
wire S25347;
wire S25348;
wire S25349;
wire S25350;
wire S25351;
wire S25352;
wire S25353;
wire S25354;
wire S25355;
wire S25356;
wire S25357;
wire S25358;
wire S25359;
wire S25360;
wire S25361;
wire S25362;
wire S25363;
wire S25364;
wire S25365;
wire S25366;
wire S25367;
wire S25368;
wire S25369;
wire S25370;
wire S25371;
wire S25372;
wire S25373;
wire S25374;
wire S25375;
wire S25376;
wire S25377;
wire S25378;
wire S25379;
wire S25380;
wire S25381;
wire S25382;
wire S25383;
wire S25384;
wire S25385;
wire S25386;
wire S25387;
wire S25388;
wire S25389;
wire S25390;
wire S25391;
wire S25392;
wire S25393;
wire S25394;
wire S25395;
wire S25396;
wire S25397;
wire S25398;
wire S25399;
wire S25400;
wire S25401;
wire S25402;
wire S25403;
wire S25404;
wire S25405;
wire S25406;
wire S25407;
wire S25408;
wire S25409;
wire S25410;
wire S25411;
wire S25412;
wire S25413;
wire S25414;
wire S25415;
wire S25416;
wire S25417;
wire S25418;
wire S25419;
wire S25420;
wire S25421;
wire S25422;
wire S25423;
wire S25424;
wire S25425;
wire S25426;
wire S25427;
wire S25428;
wire S25429;
wire S25430;
wire S25431;
wire S25432;
wire S25433;
wire S25434;
wire S25435;
wire S25436;
wire S25437;
wire S25438;
wire S25439;
wire S25440;
wire S25441;
wire S25442;
wire S25443;
wire S25444;
wire S25445;
wire S25446;
wire S25447;
wire S25448;
wire S25449;
wire S25450;
wire S25451;
wire S25452;
wire S25453;
wire S25454;
wire S25455;
wire S25456;
wire S25457;
wire S25458;
wire S25459;
wire S25460;
wire S25461;
wire S25462;
wire S25463;
wire S25464;
wire S25465;
wire S25466;
wire S25467;
wire S25468;
wire S25469;
wire S25470;
wire S25471;
wire S25472;
wire S25473;
wire S25474;
wire S25475;
wire S25476;
wire S25477;
wire S25478;
wire S25479;
wire S25480;
wire S25481;
wire S25482;
wire S25483;
wire S25484;
wire S25485;
wire S25486;
wire S25487;
wire S25488;
wire S25489;
wire S25490;
wire S25491;
wire S25492;
wire S25493;
wire S25494;
wire S25495;
wire S25496;
wire S25497;
wire S25498;
wire S25499;
wire S25500;
wire S25501;
wire S25502;
wire S25503;
wire S25504;
wire S25505;
wire S25506;
wire S25507;
wire S25508;
wire S25509;
wire S25510;
wire S25511;
wire S25512;
wire S25513;
wire S25514;
wire S25515;
wire S25516;
wire S25517;
wire S25518;
wire S25519;
wire S25520;
wire S25521;
wire S25522;
wire S25523;
wire S25524;
wire S25525;
wire S25526;
wire S25527;
wire S25528;
wire S25529;
wire S25530;
wire S25531;
wire S25532;
wire S25533;
wire S25534;
wire S25535;
wire S25536;
wire S25537;
wire S25538;
wire S25539;
wire S25540;
wire S25541;
wire S25542;
wire S25543;
wire S25544;
wire S25545;
wire S25546;
wire S25547;
wire S25548;
wire S25549;
wire S25550;
wire S25551;
wire S25552;
wire S25553;
wire S25554;
wire S25555;
wire S25556;
wire S25557;
wire S25558;
wire S25559;
wire S25560;
wire S25561;
wire S25562;
wire S25563;
wire S25564;
wire S25565;
wire S25566;
wire S25567;
wire S25568;
wire S25569;
wire S25570;
wire S25571;
wire S25572;
wire S25573;
wire S25574;
wire S25575;
wire S25576;
wire S25577;
wire S25578;
wire S25579;
wire S25580;
wire S25581;
wire S25582;
wire S25583;
wire S25584;
wire S25585;
wire S25586;
wire S25587;
wire S25588;
wire S25589;
wire S25590;
wire S25591;
wire S25592;
wire S25593;
wire S25594;
wire S25595;
wire S25596;
wire S25597;
wire S25598;
wire S25599;
wire S25600;
wire S25601;
wire S25602;
wire S25603;
wire S25604;
wire S25605;
wire S25606;
wire S25607;
wire S25608;
wire S25609;
wire S25610;
wire S25611;
wire S25612;
wire S25613;
wire S25614;
wire S25615;
wire S25616;
wire S25617;
wire S25618;
wire S25619;
wire S25620;
wire S25621;
wire S25622;
wire S25623;
wire S25624;
wire S25625;
wire S25626;
wire S25627;
wire S25628;
wire S25629;
wire S25630;
wire S25631;
wire S25632;
wire S25633;
wire S25634;
wire S25635;
wire S25636;
wire S25637;
wire S25638;
wire S25639;
wire S25640;
wire S25641;
wire S25642;
wire S25643;
wire S25644;
wire S25645;
wire S25646;
wire S25647;
wire S25648;
wire S25649;
wire S25650;
wire S25651;
wire S25652;
wire S25653;
wire S25654;
wire S25655;
wire S25656;
wire S25657;
wire S25658;
wire S25659;
wire S25660;
wire S25661;
wire S25662;
wire S25663;
wire S25664;
wire S25665;
wire S25666;
wire S25667;
wire S25668;
wire S25669;
wire S25670;
wire S25671;
wire S25672;
wire S25673;
wire S25674;
wire S25675;
wire S25676;
wire S25677;
wire S25678;
wire S25679;
wire S25680;
wire S25681;
wire S25682;
wire S25683;
wire S25684;
wire S25685;
wire S25686;
wire S25687;
wire S25688;
wire S25689;
wire S25690;
wire S25691;
wire S25692;
wire S25693;
wire S25694;
wire S25695;
wire S25696;
wire S25697;
wire S25698;
wire S25699;
wire S25700;
wire S25701;
wire S25702;
wire S25703;
wire S25704;
wire S25705;
wire S25706;
wire S25707;
wire S25708;
wire S25709;
wire S25710;
wire S25711;
wire S25712;
wire S25713;
wire S25714;
wire S25715;
wire S25716;
wire S25717;
wire S25718;
wire S25719;
wire S25720;
wire S25721;
wire S25722;
wire S25723;
wire S25724;
wire S25725;
wire S25726;
wire S25727;
wire S25728;
wire S25729;
wire S25730;
wire S25731;
wire S25732;
wire S25733;
wire S25734;
wire S25735;
wire S25736;
wire S25737;
wire S25738;
wire S25739;
wire S25740;
wire S25741;
wire S25742;
wire S25743;
wire S25744;
wire S25745;
wire S25746;
wire S25747;
wire S25748;
wire S25749;
wire S25750;
wire S25751;
wire S25752;
wire S25753;
wire S25754;
wire S25755;
wire S25756;
wire S25757;
wire S25758;
wire S25759;
wire S25760;
wire S25761;
wire S25762;
wire S25763;
wire S25764;
wire S25765;
wire S25766;
wire S25767;
wire S25768;
wire S25769;
wire S25770;
wire S25771;
wire S25772;
wire S25773;
wire S25774;
wire S25775;
wire S25776;
wire S25777;
wire S25778;
wire S25779;
wire S25780;
wire S25781;
wire S25782;
wire S25783;
wire S25784;
wire S25785;
wire S25786;
wire S25787;
wire S25788;
wire S25789;
wire S25790;
wire S25791;
wire S25792;
wire S25793;
wire S25794;
wire S25795;
wire S25796;
wire S25797;
wire S25798;
wire S25799;
wire S25800;
wire S25801;
wire S25802;
wire S25803;
wire S25804;
wire S25805;
wire S25806;
wire S25807;
wire S25808;
wire S25809;
wire S25810;
wire S25811;
wire S25812;
wire S25813;
wire S25814;
wire S25815;
wire S25816;
wire S25817;
wire S25818;
wire S25819;
wire S25820;
wire S25821;
wire S25822;
wire S25823;
wire S25824;
wire S25825;
wire S25826;
wire S25827;
wire S25828;
wire S25829;
wire S25830;
wire S25831;
wire S25832;
wire S25833;
wire S25834;
wire S25835;
wire S25836;
wire S25837;
wire S25838;
wire S25839;
wire S25840;
wire S25841;
wire S25842;
wire S25843;
wire S25844;
wire S25845;
wire S25846;
wire S25847;
wire S25848;
wire S25849;
wire S25850;
wire S25851;
wire S25852;
wire S25853;
wire S25854;
wire S25855;
wire S25856;
wire S25857;
wire S25858;
wire S25859;
wire S25860;
wire S25861;
wire S25862;
wire S25863;
wire S25864;
wire S25865;
wire S25866;
wire S25867;
wire S25868;
wire S25869;
wire S25870;
wire S25871;
wire S25872;
wire S25873;
wire S25874;
wire S25875;
wire S25876;
wire S25877;
wire S25878;
wire S25879;
wire S25880;
wire S25881;
wire S25882;
wire S25883;
wire S25884;
wire S25885;
wire S25886;
wire S25887;
wire S25888;
wire S25889;
wire S25890;
wire S25891;
wire S25892;
wire S25893;
wire S25894;
wire S25895;
wire S25896;
wire S25897;
wire S25898;
wire S25899;
wire S25900;
wire S25901;
wire S25902;
wire S25903;
wire S25904;
wire S25905;
wire S25906;
wire S25907;
wire S25908;
wire S25909;
wire S25910;
wire S25911;
wire S25912;
wire S25913;
wire S25914;
wire S25915;
wire S25916;
wire S25917;
wire S25918;
wire S25919;
wire S25920;
wire S25921;
wire S25922;
wire S25923;
wire S25924;
wire S25925;
wire S25926;
wire S25927;
wire S25928;
wire S25929;
wire S25930;
wire S25931;
wire S25932;
wire S25933;
wire S25934;
wire S25935;
wire S25936;
wire S25937;
wire S25938;
wire S25939;
wire S25940;
wire S25941;
wire S25942;
wire S25943;
wire S25944;
wire S25945;
wire S25946;
wire S25947;
wire S25948;
wire S25949;
wire S25950;
wire S25951;
wire S25952;
wire S25953;
wire S25954;
wire S25955;
wire S25956;
wire S25957;
wire new_0;
wire new_10;
wire new_11;
wire new_12;
wire new_13;
wire new_14;
wire new_15;
wire new_16;
wire new_17;
wire new_18;
wire new_19;
wire new_1;
wire new_20;
wire new_21;
wire new_22;
wire new_23;
wire new_24;
wire new_25;
wire new_26;
wire new_27;
wire new_28;
wire new_29;
wire new_2;
wire new_30;
wire new_31;
wire new_3;
wire new_4;
wire new_5;
wire new_6;
wire new_7;
wire new_8;
wire new_9;
wire rot_0;
wire rot_10;
wire rot_11;
wire rot_12;
wire rot_13;
wire rot_14;
wire rot_15;
wire rot_16;
wire rot_17;
wire rot_18;
wire rot_19;
wire rot_1;
wire rot_20;
wire rot_21;
wire rot_22;
wire rot_23;
wire rot_24;
wire rot_25;
wire rot_26;
wire rot_27;
wire rot_28;
wire rot_29;
wire rot_2;
wire rot_30;
wire rot_31;
wire rot_3;
wire rot_4;
wire rot_5;
wire rot_6;
wire rot_7;
wire rot_8;
wire rot_9;
wire temp_0;
wire temp_10;
wire temp_11;
wire temp_12;
wire temp_13;
wire temp_14;
wire temp_15;
wire temp_16;
wire temp_17;
wire temp_18;
wire temp_19;
wire temp_1;
wire temp_20;
wire temp_21;
wire temp_22;
wire temp_23;
wire temp_24;
wire temp_25;
wire temp_26;
wire temp_27;
wire temp_28;
wire temp_29;
wire temp_2;
wire temp_30;
wire temp_31;
wire temp_3;
wire temp_4;
wire temp_5;
wire temp_6;
wire temp_7;
wire temp_8;
wire temp_9;
input [127:0] key;output [1407:0] w;
INV_X1 #() 
INV_X1_1_ (
  .A({ S27 }),
  .ZN({ S156 })
);
NAND2_X1 #() 
NAND2_X1_1_ (
  .A1({ S29 }),
  .A2({ S25956[11] }),
  .ZN({ S157 })
);
OAI21_X1 #() 
OAI21_X1_1_ (
  .A({ S157 }),
  .B1({ S156 }),
  .B2({ S25956[11] }),
  .ZN({ S116 })
);
INV_X1 #() 
INV_X1_2_ (
  .A({ S56 }),
  .ZN({ S158 })
);
NAND2_X1 #() 
NAND2_X1_2_ (
  .A1({ S58 }),
  .A2({ S25956[3] }),
  .ZN({ S159 })
);
OAI21_X1 #() 
OAI21_X1_2_ (
  .A({ S159 }),
  .B1({ S158 }),
  .B2({ S25956[3] }),
  .ZN({ S117 })
);
INV_X1 #() 
INV_X1_3_ (
  .A({ S66 }),
  .ZN({ S160 })
);
NAND2_X1 #() 
NAND2_X1_3_ (
  .A1({ S67 }),
  .A2({ S25956[27] }),
  .ZN({ S161 })
);
OAI21_X1 #() 
OAI21_X1_3_ (
  .A({ S161 }),
  .B1({ S160 }),
  .B2({ S25956[27] }),
  .ZN({ S118 })
);
INV_X1 #() 
INV_X1_4_ (
  .A({ S69 }),
  .ZN({ S162 })
);
NAND2_X1 #() 
NAND2_X1_4_ (
  .A1({ S70 }),
  .A2({ S25956[19] }),
  .ZN({ S163 })
);
OAI21_X1 #() 
OAI21_X1_4_ (
  .A({ S163 }),
  .B1({ S162 }),
  .B2({ S25956[19] }),
  .ZN({ S119 })
);
INV_X1 #() 
INV_X1_5_ (
  .A({ S72 }),
  .ZN({ S164 })
);
NAND2_X1 #() 
NAND2_X1_5_ (
  .A1({ S73 }),
  .A2({ S65 }),
  .ZN({ S165 })
);
OAI21_X1 #() 
OAI21_X1_5_ (
  .A({ S165 }),
  .B1({ S164 }),
  .B2({ S65 }),
  .ZN({ S120 })
);
INV_X1 #() 
INV_X1_6_ (
  .A({ S75 }),
  .ZN({ S166 })
);
NAND2_X1 #() 
NAND2_X1_6_ (
  .A1({ S76 }),
  .A2({ S68 }),
  .ZN({ S167 })
);
OAI21_X1 #() 
OAI21_X1_6_ (
  .A({ S167 }),
  .B1({ S166 }),
  .B2({ S68 }),
  .ZN({ S121 })
);
INV_X1 #() 
INV_X1_7_ (
  .A({ S78 }),
  .ZN({ S168 })
);
NAND2_X1 #() 
NAND2_X1_7_ (
  .A1({ S79 }),
  .A2({ S71 }),
  .ZN({ S169 })
);
OAI21_X1 #() 
OAI21_X1_7_ (
  .A({ S169 }),
  .B1({ S168 }),
  .B2({ S71 }),
  .ZN({ S122 })
);
INV_X1 #() 
INV_X1_8_ (
  .A({ S81 }),
  .ZN({ S170 })
);
NAND2_X1 #() 
NAND2_X1_8_ (
  .A1({ S82 }),
  .A2({ S50 }),
  .ZN({ S171 })
);
OAI21_X1 #() 
OAI21_X1_8_ (
  .A({ S171 }),
  .B1({ S170 }),
  .B2({ S50 }),
  .ZN({ S123 })
);
INV_X1 #() 
INV_X1_9_ (
  .A({ S84 }),
  .ZN({ S172 })
);
NAND2_X1 #() 
NAND2_X1_9_ (
  .A1({ S85 }),
  .A2({ S77 }),
  .ZN({ S173 })
);
OAI21_X1 #() 
OAI21_X1_9_ (
  .A({ S173 }),
  .B1({ S172 }),
  .B2({ S77 }),
  .ZN({ S124 })
);
INV_X1 #() 
INV_X1_10_ (
  .A({ S87 }),
  .ZN({ S174 })
);
NAND2_X1 #() 
NAND2_X1_10_ (
  .A1({ S88 }),
  .A2({ S80 }),
  .ZN({ S175 })
);
OAI21_X1 #() 
OAI21_X1_10_ (
  .A({ S175 }),
  .B1({ S174 }),
  .B2({ S80 }),
  .ZN({ S125 })
);
INV_X1 #() 
INV_X1_11_ (
  .A({ S90 }),
  .ZN({ S176 })
);
NAND2_X1 #() 
NAND2_X1_11_ (
  .A1({ S91 }),
  .A2({ S83 }),
  .ZN({ S177 })
);
OAI21_X1 #() 
OAI21_X1_11_ (
  .A({ S177 }),
  .B1({ S176 }),
  .B2({ S83 }),
  .ZN({ S126 })
);
INV_X1 #() 
INV_X1_12_ (
  .A({ S93 }),
  .ZN({ S178 })
);
NAND2_X1 #() 
NAND2_X1_12_ (
  .A1({ S94 }),
  .A2({ S74 }),
  .ZN({ S179 })
);
OAI21_X1 #() 
OAI21_X1_12_ (
  .A({ S179 }),
  .B1({ S178 }),
  .B2({ S74 }),
  .ZN({ S127 })
);
INV_X1 #() 
INV_X1_13_ (
  .A({ S96 }),
  .ZN({ S180 })
);
NAND2_X1 #() 
NAND2_X1_13_ (
  .A1({ S97 }),
  .A2({ S89 }),
  .ZN({ S181 })
);
OAI21_X1 #() 
OAI21_X1_13_ (
  .A({ S181 }),
  .B1({ S180 }),
  .B2({ S89 }),
  .ZN({ S128 })
);
INV_X1 #() 
INV_X1_14_ (
  .A({ S99 }),
  .ZN({ S182 })
);
NAND2_X1 #() 
NAND2_X1_14_ (
  .A1({ S100 }),
  .A2({ S92 }),
  .ZN({ S183 })
);
OAI21_X1 #() 
OAI21_X1_14_ (
  .A({ S183 }),
  .B1({ S182 }),
  .B2({ S92 }),
  .ZN({ S129 })
);
INV_X1 #() 
INV_X1_15_ (
  .A({ S102 }),
  .ZN({ S184 })
);
NAND2_X1 #() 
NAND2_X1_15_ (
  .A1({ S103 }),
  .A2({ S95 }),
  .ZN({ S185 })
);
OAI21_X1 #() 
OAI21_X1_15_ (
  .A({ S185 }),
  .B1({ S184 }),
  .B2({ S95 }),
  .ZN({ S130 })
);
INV_X1 #() 
INV_X1_16_ (
  .A({ S105 }),
  .ZN({ S186 })
);
NAND2_X1 #() 
NAND2_X1_16_ (
  .A1({ S106 }),
  .A2({ S86 }),
  .ZN({ S187 })
);
OAI21_X1 #() 
OAI21_X1_16_ (
  .A({ S187 }),
  .B1({ S186 }),
  .B2({ S86 }),
  .ZN({ S131 })
);
INV_X1 #() 
INV_X1_17_ (
  .A({ S108 }),
  .ZN({ S188 })
);
NAND2_X1 #() 
NAND2_X1_17_ (
  .A1({ S109 }),
  .A2({ S101 }),
  .ZN({ S189 })
);
OAI21_X1 #() 
OAI21_X1_17_ (
  .A({ S189 }),
  .B1({ S188 }),
  .B2({ S101 }),
  .ZN({ S132 })
);
INV_X1 #() 
INV_X1_18_ (
  .A({ S111 }),
  .ZN({ S190 })
);
NAND2_X1 #() 
NAND2_X1_18_ (
  .A1({ S112 }),
  .A2({ S104 }),
  .ZN({ S191 })
);
OAI21_X1 #() 
OAI21_X1_18_ (
  .A({ S191 }),
  .B1({ S190 }),
  .B2({ S104 }),
  .ZN({ S133 })
);
INV_X1 #() 
INV_X1_19_ (
  .A({ S114 }),
  .ZN({ S192 })
);
NAND2_X1 #() 
NAND2_X1_19_ (
  .A1({ S115 }),
  .A2({ S107 }),
  .ZN({ S193 })
);
OAI21_X1 #() 
OAI21_X1_19_ (
  .A({ S193 }),
  .B1({ S192 }),
  .B2({ S107 }),
  .ZN({ S134 })
);
INV_X1 #() 
INV_X1_20_ (
  .A({ S1 }),
  .ZN({ S194 })
);
NAND2_X1 #() 
NAND2_X1_20_ (
  .A1({ S2 }),
  .A2({ S98 }),
  .ZN({ S195 })
);
OAI21_X1 #() 
OAI21_X1_20_ (
  .A({ S195 }),
  .B1({ S194 }),
  .B2({ S98 }),
  .ZN({ S135 })
);
INV_X1 #() 
INV_X1_21_ (
  .A({ S4 }),
  .ZN({ S196 })
);
NAND2_X1 #() 
NAND2_X1_21_ (
  .A1({ S5 }),
  .A2({ S113 }),
  .ZN({ S197 })
);
OAI21_X1 #() 
OAI21_X1_21_ (
  .A({ S197 }),
  .B1({ S196 }),
  .B2({ S113 }),
  .ZN({ S136 })
);
INV_X1 #() 
INV_X1_22_ (
  .A({ S7 }),
  .ZN({ S198 })
);
NAND2_X1 #() 
NAND2_X1_22_ (
  .A1({ S8 }),
  .A2({ S0 }),
  .ZN({ S199 })
);
OAI21_X1 #() 
OAI21_X1_22_ (
  .A({ S199 }),
  .B1({ S198 }),
  .B2({ S0 }),
  .ZN({ S137 })
);
INV_X1 #() 
INV_X1_23_ (
  .A({ S10 }),
  .ZN({ S200 })
);
NAND2_X1 #() 
NAND2_X1_23_ (
  .A1({ S11 }),
  .A2({ S3 }),
  .ZN({ S201 })
);
OAI21_X1 #() 
OAI21_X1_23_ (
  .A({ S201 }),
  .B1({ S200 }),
  .B2({ S3 }),
  .ZN({ S138 })
);
INV_X1 #() 
INV_X1_24_ (
  .A({ S13 }),
  .ZN({ S202 })
);
NAND2_X1 #() 
NAND2_X1_24_ (
  .A1({ S14 }),
  .A2({ S110 }),
  .ZN({ S203 })
);
OAI21_X1 #() 
OAI21_X1_24_ (
  .A({ S203 }),
  .B1({ S202 }),
  .B2({ S110 }),
  .ZN({ S139 })
);
INV_X1 #() 
INV_X1_25_ (
  .A({ S16 }),
  .ZN({ S204 })
);
NAND2_X1 #() 
NAND2_X1_25_ (
  .A1({ S17 }),
  .A2({ S9 }),
  .ZN({ S205 })
);
OAI21_X1 #() 
OAI21_X1_25_ (
  .A({ S205 }),
  .B1({ S204 }),
  .B2({ S9 }),
  .ZN({ S140 })
);
INV_X1 #() 
INV_X1_26_ (
  .A({ S19 }),
  .ZN({ S206 })
);
NAND2_X1 #() 
NAND2_X1_26_ (
  .A1({ S20 }),
  .A2({ S12 }),
  .ZN({ S207 })
);
OAI21_X1 #() 
OAI21_X1_26_ (
  .A({ S207 }),
  .B1({ S206 }),
  .B2({ S12 }),
  .ZN({ S141 })
);
INV_X1 #() 
INV_X1_27_ (
  .A({ S22 }),
  .ZN({ S208 })
);
NAND2_X1 #() 
NAND2_X1_27_ (
  .A1({ S23 }),
  .A2({ S15 }),
  .ZN({ S209 })
);
OAI21_X1 #() 
OAI21_X1_27_ (
  .A({ S209 }),
  .B1({ S208 }),
  .B2({ S15 }),
  .ZN({ S142 })
);
INV_X1 #() 
INV_X1_28_ (
  .A({ S25 }),
  .ZN({ S210 })
);
NAND2_X1 #() 
NAND2_X1_28_ (
  .A1({ S26 }),
  .A2({ S6 }),
  .ZN({ S211 })
);
OAI21_X1 #() 
OAI21_X1_28_ (
  .A({ S211 }),
  .B1({ S210 }),
  .B2({ S6 }),
  .ZN({ S143 })
);
INV_X1 #() 
INV_X1_29_ (
  .A({ S30 }),
  .ZN({ S212 })
);
NAND2_X1 #() 
NAND2_X1_29_ (
  .A1({ S31 }),
  .A2({ S21 }),
  .ZN({ S213 })
);
OAI21_X1 #() 
OAI21_X1_29_ (
  .A({ S213 }),
  .B1({ S212 }),
  .B2({ S21 }),
  .ZN({ S144 })
);
INV_X1 #() 
INV_X1_30_ (
  .A({ S33 }),
  .ZN({ S214 })
);
NAND2_X1 #() 
NAND2_X1_30_ (
  .A1({ S34 }),
  .A2({ S24 }),
  .ZN({ S215 })
);
OAI21_X1 #() 
OAI21_X1_30_ (
  .A({ S215 }),
  .B1({ S214 }),
  .B2({ S24 }),
  .ZN({ S145 })
);
INV_X1 #() 
INV_X1_31_ (
  .A({ S36 }),
  .ZN({ S216 })
);
NAND2_X1 #() 
NAND2_X1_31_ (
  .A1({ S37 }),
  .A2({ S28 }),
  .ZN({ S217 })
);
OAI21_X1 #() 
OAI21_X1_31_ (
  .A({ S217 }),
  .B1({ S216 }),
  .B2({ S28 }),
  .ZN({ S146 })
);
INV_X1 #() 
INV_X1_32_ (
  .A({ S39 }),
  .ZN({ S218 })
);
NAND2_X1 #() 
NAND2_X1_32_ (
  .A1({ S40 }),
  .A2({ S18 }),
  .ZN({ S219 })
);
OAI21_X1 #() 
OAI21_X1_32_ (
  .A({ S219 }),
  .B1({ S218 }),
  .B2({ S18 }),
  .ZN({ S147 })
);
INV_X1 #() 
INV_X1_33_ (
  .A({ S42 }),
  .ZN({ S220 })
);
NAND2_X1 #() 
NAND2_X1_33_ (
  .A1({ S43 }),
  .A2({ S35 }),
  .ZN({ S221 })
);
OAI21_X1 #() 
OAI21_X1_33_ (
  .A({ S221 }),
  .B1({ S220 }),
  .B2({ S35 }),
  .ZN({ S148 })
);
INV_X1 #() 
INV_X1_34_ (
  .A({ S45 }),
  .ZN({ S222 })
);
NAND2_X1 #() 
NAND2_X1_34_ (
  .A1({ S46 }),
  .A2({ S38 }),
  .ZN({ S223 })
);
OAI21_X1 #() 
OAI21_X1_34_ (
  .A({ S223 }),
  .B1({ S222 }),
  .B2({ S38 }),
  .ZN({ S149 })
);
INV_X1 #() 
INV_X1_35_ (
  .A({ S48 }),
  .ZN({ S224 })
);
NAND2_X1 #() 
NAND2_X1_35_ (
  .A1({ S49 }),
  .A2({ S41 }),
  .ZN({ S225 })
);
OAI21_X1 #() 
OAI21_X1_35_ (
  .A({ S225 }),
  .B1({ S224 }),
  .B2({ S41 }),
  .ZN({ S150 })
);
INV_X1 #() 
INV_X1_36_ (
  .A({ S52 }),
  .ZN({ S226 })
);
NAND2_X1 #() 
NAND2_X1_36_ (
  .A1({ S53 }),
  .A2({ S32 }),
  .ZN({ S227 })
);
OAI21_X1 #() 
OAI21_X1_36_ (
  .A({ S227 }),
  .B1({ S226 }),
  .B2({ S32 }),
  .ZN({ S151 })
);
INV_X1 #() 
INV_X1_37_ (
  .A({ S55 }),
  .ZN({ S228 })
);
NAND2_X1 #() 
NAND2_X1_37_ (
  .A1({ S57 }),
  .A2({ S54 }),
  .ZN({ S229 })
);
OAI21_X1 #() 
OAI21_X1_37_ (
  .A({ S229 }),
  .B1({ S228 }),
  .B2({ S54 }),
  .ZN({ S152 })
);
INV_X1 #() 
INV_X1_38_ (
  .A({ S59 }),
  .ZN({ S230 })
);
NAND2_X1 #() 
NAND2_X1_38_ (
  .A1({ S60 }),
  .A2({ S51 }),
  .ZN({ S231 })
);
OAI21_X1 #() 
OAI21_X1_38_ (
  .A({ S231 }),
  .B1({ S230 }),
  .B2({ S51 }),
  .ZN({ S153 })
);
INV_X1 #() 
INV_X1_39_ (
  .A({ S61 }),
  .ZN({ S232 })
);
NAND2_X1 #() 
NAND2_X1_39_ (
  .A1({ S62 }),
  .A2({ S47 }),
  .ZN({ S233 })
);
OAI21_X1 #() 
OAI21_X1_39_ (
  .A({ S233 }),
  .B1({ S232 }),
  .B2({ S47 }),
  .ZN({ S154 })
);
INV_X1 #() 
INV_X1_40_ (
  .A({ S63 }),
  .ZN({ S234 })
);
NAND2_X1 #() 
NAND2_X1_40_ (
  .A1({ S64 }),
  .A2({ S44 }),
  .ZN({ S235 })
);
OAI21_X1 #() 
OAI21_X1_40_ (
  .A({ S235 }),
  .B1({ S234 }),
  .B2({ S44 }),
  .ZN({ S155 })
);
AOI21_X1 #() 
AOI21_X1_1_ (
  .A({ S5495 }),
  .B1({ S6076 }),
  .B2({ S25957[645] }),
  .ZN({ S6077 })
);
NAND2_X1 #() 
NAND2_X1_41_ (
  .A1({ S6077 }),
  .A2({ S6075 }),
  .ZN({ S6078 })
);
NAND3_X1 #() 
NAND3_X1_1_ (
  .A1({ S6074 }),
  .A2({ S6078 }),
  .A3({ S25957[646] }),
  .ZN({ S6079 })
);
OAI21_X1 #() 
OAI21_X1_41_ (
  .A({ S6027 }),
  .B1({ S6025 }),
  .B2({ S5533 }),
  .ZN({ S6080 })
);
NAND2_X1 #() 
NAND2_X1_42_ (
  .A1({ S6080 }),
  .A2({ S25957[645] }),
  .ZN({ S6082 })
);
OAI21_X1 #() 
OAI21_X1_42_ (
  .A({ S6029 }),
  .B1({ S6030 }),
  .B2({ S25957[643] }),
  .ZN({ S6083 })
);
NAND2_X1 #() 
NAND2_X1_43_ (
  .A1({ S6083 }),
  .A2({ S25957[644] }),
  .ZN({ S6084 })
);
AOI21_X1 #() 
AOI21_X1_2_ (
  .A({ S25957[643] }),
  .B1({ S5604 }),
  .B2({ S5512 }),
  .ZN({ S6085 })
);
AOI21_X1 #() 
AOI21_X1_3_ (
  .A({ S6085 }),
  .B1({ S5748 }),
  .B2({ S25957[643] }),
  .ZN({ S6086 })
);
OAI211_X1 #() 
OAI211_X1_1_ (
  .A({ S5494 }),
  .B({ S6084 }),
  .C1({ S6086 }),
  .C2({ S25957[644] }),
  .ZN({ S6087 })
);
NAND3_X1 #() 
NAND3_X1_2_ (
  .A1({ S6087 }),
  .A2({ S6082 }),
  .A3({ S5465 }),
  .ZN({ S6088 })
);
NAND3_X1 #() 
NAND3_X1_3_ (
  .A1({ S6088 }),
  .A2({ S25957[647] }),
  .A3({ S6079 }),
  .ZN({ S6089 })
);
NAND3_X1 #() 
NAND3_X1_4_ (
  .A1({ S6089 }),
  .A2({ S25957[745] }),
  .A3({ S6069 }),
  .ZN({ S6090 })
);
NAND3_X1 #() 
NAND3_X1_5_ (
  .A1({ S6090 }),
  .A2({ S3355 }),
  .A3({ S6054 }),
  .ZN({ S6091 })
);
NAND3_X1 #() 
NAND3_X1_6_ (
  .A1({ S6035 }),
  .A2({ S6053 }),
  .A3({ S25957[745] }),
  .ZN({ S6093 })
);
NAND3_X1 #() 
NAND3_X1_7_ (
  .A1({ S6089 }),
  .A2({ S6013 }),
  .A3({ S6069 }),
  .ZN({ S6094 })
);
NAND3_X1 #() 
NAND3_X1_8_ (
  .A1({ S6094 }),
  .A2({ S25957[809] }),
  .A3({ S6093 }),
  .ZN({ S6095 })
);
NAND3_X1 #() 
NAND3_X1_9_ (
  .A1({ S6091 }),
  .A2({ S6095 }),
  .A3({ S4806 }),
  .ZN({ S6096 })
);
NAND3_X1 #() 
NAND3_X1_10_ (
  .A1({ S6094 }),
  .A2({ S3355 }),
  .A3({ S6093 }),
  .ZN({ S6097 })
);
NAND3_X1 #() 
NAND3_X1_11_ (
  .A1({ S6090 }),
  .A2({ S25957[809] }),
  .A3({ S6054 }),
  .ZN({ S6098 })
);
NAND3_X1 #() 
NAND3_X1_12_ (
  .A1({ S6097 }),
  .A2({ S6098 }),
  .A3({ S25957[649] }),
  .ZN({ S6099 })
);
NAND2_X1 #() 
NAND2_X1_44_ (
  .A1({ S6096 }),
  .A2({ S6099 }),
  .ZN({ S25957[521] })
);
NAND2_X1 #() 
NAND2_X1_45_ (
  .A1({ S3473 }),
  .A2({ S3476 }),
  .ZN({ S6100 })
);
INV_X1 #() 
INV_X1_41_ (
  .A({ S6100 }),
  .ZN({ S25957[682] })
);
NAND2_X1 #() 
NAND2_X1_46_ (
  .A1({ S1007 }),
  .A2({ S1008 }),
  .ZN({ S25957[874] })
);
XNOR2_X1 #() 
XNOR2_X1_1_ (
  .A({ S25957[874] }),
  .B({ S3412 }),
  .ZN({ S25957[842] })
);
INV_X1 #() 
INV_X1_42_ (
  .A({ S25957[842] }),
  .ZN({ S6102 })
);
NAND3_X1 #() 
NAND3_X1_13_ (
  .A1({ S5565 }),
  .A2({ S5714 }),
  .A3({ S25957[643] }),
  .ZN({ S6103 })
);
OAI211_X1 #() 
OAI211_X1_2_ (
  .A({ S6103 }),
  .B({ S25957[644] }),
  .C1({ S5627 }),
  .C2({ S5773 }),
  .ZN({ S6104 })
);
NAND4_X1 #() 
NAND4_X1_1_ (
  .A1({ S5501 }),
  .A2({ S25957[643] }),
  .A3({ S5475 }),
  .A4({ S5508 }),
  .ZN({ S6105 })
);
AOI22_X1 #() 
AOI22_X1_1_ (
  .A1({ S5608 }),
  .A2({ S0 }),
  .B1({ S3849 }),
  .B2({ S3846 }),
  .ZN({ S6106 })
);
AOI21_X1 #() 
AOI21_X1_4_ (
  .A({ S5494 }),
  .B1({ S6106 }),
  .B2({ S6105 }),
  .ZN({ S6107 })
);
NAND2_X1 #() 
NAND2_X1_47_ (
  .A1({ S6107 }),
  .A2({ S6104 }),
  .ZN({ S6108 })
);
NAND2_X1 #() 
NAND2_X1_48_ (
  .A1({ S5623 }),
  .A2({ S25957[643] }),
  .ZN({ S6109 })
);
NAND3_X1 #() 
NAND3_X1_14_ (
  .A1({ S5756 }),
  .A2({ S25957[644] }),
  .A3({ S6109 }),
  .ZN({ S6111 })
);
NAND3_X1 #() 
NAND3_X1_15_ (
  .A1({ S5642 }),
  .A2({ S5495 }),
  .A3({ S5931 }),
  .ZN({ S6112 })
);
NAND3_X1 #() 
NAND3_X1_16_ (
  .A1({ S6112 }),
  .A2({ S5494 }),
  .A3({ S6111 }),
  .ZN({ S6113 })
);
NAND3_X1 #() 
NAND3_X1_17_ (
  .A1({ S6113 }),
  .A2({ S5530 }),
  .A3({ S6108 }),
  .ZN({ S6114 })
);
OAI211_X1 #() 
OAI211_X1_3_ (
  .A({ S25957[643] }),
  .B({ S5497 }),
  .C1({ S5498 }),
  .C2({ S5471 }),
  .ZN({ S6115 })
);
AND3_X1 #() 
AND3_X1_1_ (
  .A1({ S6115 }),
  .A2({ S5590 }),
  .A3({ S5495 }),
  .ZN({ S6116 })
);
AOI21_X1 #() 
AOI21_X1_5_ (
  .A({ S0 }),
  .B1({ S5565 }),
  .B2({ S5488 }),
  .ZN({ S6117 })
);
OAI21_X1 #() 
OAI21_X1_43_ (
  .A({ S25957[644] }),
  .B1({ S5554 }),
  .B2({ S25957[643] }),
  .ZN({ S6118 })
);
OAI21_X1 #() 
OAI21_X1_44_ (
  .A({ S25957[645] }),
  .B1({ S6118 }),
  .B2({ S6117 }),
  .ZN({ S6119 })
);
INV_X1 #() 
INV_X1_43_ (
  .A({ S6109 }),
  .ZN({ S6120 })
);
NAND3_X1 #() 
NAND3_X1_18_ (
  .A1({ S5609 }),
  .A2({ S5495 }),
  .A3({ S5607 }),
  .ZN({ S6122 })
);
OAI21_X1 #() 
OAI21_X1_45_ (
  .A({ S25957[644] }),
  .B1({ S25957[643] }),
  .B2({ S5551 }),
  .ZN({ S6123 })
);
OAI211_X1 #() 
OAI211_X1_4_ (
  .A({ S6122 }),
  .B({ S5494 }),
  .C1({ S6123 }),
  .C2({ S6120 }),
  .ZN({ S6124 })
);
OAI211_X1 #() 
OAI211_X1_5_ (
  .A({ S6124 }),
  .B({ S25957[647] }),
  .C1({ S6116 }),
  .C2({ S6119 }),
  .ZN({ S6125 })
);
NAND2_X1 #() 
NAND2_X1_49_ (
  .A1({ S6114 }),
  .A2({ S6125 }),
  .ZN({ S6126 })
);
NAND2_X1 #() 
NAND2_X1_50_ (
  .A1({ S6126 }),
  .A2({ S5465 }),
  .ZN({ S6127 })
);
OAI21_X1 #() 
OAI21_X1_46_ (
  .A({ S0 }),
  .B1({ S5942 }),
  .B2({ S5623 }),
  .ZN({ S6128 })
);
AOI21_X1 #() 
AOI21_X1_6_ (
  .A({ S5495 }),
  .B1({ S6062 }),
  .B2({ S25957[643] }),
  .ZN({ S6129 })
);
NAND2_X1 #() 
NAND2_X1_51_ (
  .A1({ S6128 }),
  .A2({ S6129 }),
  .ZN({ S6130 })
);
NAND3_X1 #() 
NAND3_X1_19_ (
  .A1({ S5489 }),
  .A2({ S25957[643] }),
  .A3({ S5704 }),
  .ZN({ S6131 })
);
NOR2_X1 #() 
NOR2_X1_1_ (
  .A1({ S5559 }),
  .A2({ S25957[644] }),
  .ZN({ S6133 })
);
NAND2_X1 #() 
NAND2_X1_52_ (
  .A1({ S6131 }),
  .A2({ S6133 }),
  .ZN({ S6134 })
);
NAND3_X1 #() 
NAND3_X1_20_ (
  .A1({ S6134 }),
  .A2({ S6130 }),
  .A3({ S25957[645] }),
  .ZN({ S6135 })
);
OAI21_X1 #() 
OAI21_X1_47_ (
  .A({ S25957[644] }),
  .B1({ S5504 }),
  .B2({ S25957[641] }),
  .ZN({ S6136 })
);
NAND3_X1 #() 
NAND3_X1_21_ (
  .A1({ S5561 }),
  .A2({ S5495 }),
  .A3({ S5920 }),
  .ZN({ S6137 })
);
OAI21_X1 #() 
OAI21_X1_48_ (
  .A({ S5484 }),
  .B1({ S5479 }),
  .B2({ S5508 }),
  .ZN({ S6138 })
);
NOR3_X1 #() 
NOR3_X1_1_ (
  .A1({ S6138 }),
  .A2({ S5623 }),
  .A3({ S0 }),
  .ZN({ S6139 })
);
OAI211_X1 #() 
OAI211_X1_6_ (
  .A({ S5494 }),
  .B({ S6137 }),
  .C1({ S6139 }),
  .C2({ S6136 }),
  .ZN({ S6140 })
);
AND3_X1 #() 
AND3_X1_2_ (
  .A1({ S6135 }),
  .A2({ S25957[647] }),
  .A3({ S6140 }),
  .ZN({ S6141 })
);
NAND3_X1 #() 
NAND3_X1_22_ (
  .A1({ S0 }),
  .A2({ S25957[640] }),
  .A3({ S5544 }),
  .ZN({ S6142 })
);
OAI211_X1 #() 
OAI211_X1_7_ (
  .A({ S25957[645] }),
  .B({ S6142 }),
  .C1({ S5499 }),
  .C2({ S5502 }),
  .ZN({ S6144 })
);
NAND4_X1 #() 
NAND4_X1_2_ (
  .A1({ S5604 }),
  .A2({ S5485 }),
  .A3({ S5484 }),
  .A4({ S0 }),
  .ZN({ S6145 })
);
NAND3_X1 #() 
NAND3_X1_23_ (
  .A1({ S6145 }),
  .A2({ S5494 }),
  .A3({ S6109 }),
  .ZN({ S6146 })
);
AOI21_X1 #() 
AOI21_X1_7_ (
  .A({ S25957[644] }),
  .B1({ S6144 }),
  .B2({ S6146 }),
  .ZN({ S6147 })
);
OAI21_X1 #() 
OAI21_X1_49_ (
  .A({ S5543 }),
  .B1({ S5722 }),
  .B2({ S5759 }),
  .ZN({ S6148 })
);
NAND2_X1 #() 
NAND2_X1_53_ (
  .A1({ S6148 }),
  .A2({ S25957[645] }),
  .ZN({ S6149 })
);
NAND3_X1 #() 
NAND3_X1_24_ (
  .A1({ S5604 }),
  .A2({ S25957[643] }),
  .A3({ S5484 }),
  .ZN({ S6150 })
);
NAND3_X1 #() 
NAND3_X1_25_ (
  .A1({ S5635 }),
  .A2({ S0 }),
  .A3({ S25957[640] }),
  .ZN({ S6151 })
);
NAND3_X1 #() 
NAND3_X1_26_ (
  .A1({ S6150 }),
  .A2({ S6151 }),
  .A3({ S5494 }),
  .ZN({ S6152 })
);
AOI21_X1 #() 
AOI21_X1_8_ (
  .A({ S5495 }),
  .B1({ S6149 }),
  .B2({ S6152 }),
  .ZN({ S6153 })
);
NOR3_X1 #() 
NOR3_X1_2_ (
  .A1({ S6147 }),
  .A2({ S6153 }),
  .A3({ S25957[647] }),
  .ZN({ S6155 })
);
OAI21_X1 #() 
OAI21_X1_50_ (
  .A({ S25957[646] }),
  .B1({ S6155 }),
  .B2({ S6141 }),
  .ZN({ S6156 })
);
AOI21_X1 #() 
AOI21_X1_9_ (
  .A({ S6102 }),
  .B1({ S6156 }),
  .B2({ S6127 }),
  .ZN({ S6157 })
);
NAND2_X1 #() 
NAND2_X1_54_ (
  .A1({ S6148 }),
  .A2({ S25957[644] }),
  .ZN({ S6158 })
);
OAI211_X1 #() 
OAI211_X1_8_ (
  .A({ S5495 }),
  .B({ S6142 }),
  .C1({ S5499 }),
  .C2({ S5502 }),
  .ZN({ S6159 })
);
NAND3_X1 #() 
NAND3_X1_27_ (
  .A1({ S6159 }),
  .A2({ S6158 }),
  .A3({ S25957[645] }),
  .ZN({ S6160 })
);
NAND3_X1 #() 
NAND3_X1_28_ (
  .A1({ S6150 }),
  .A2({ S6151 }),
  .A3({ S25957[644] }),
  .ZN({ S6161 })
);
NAND3_X1 #() 
NAND3_X1_29_ (
  .A1({ S6145 }),
  .A2({ S5495 }),
  .A3({ S6109 }),
  .ZN({ S6162 })
);
NAND3_X1 #() 
NAND3_X1_30_ (
  .A1({ S6162 }),
  .A2({ S6161 }),
  .A3({ S5494 }),
  .ZN({ S6163 })
);
AND3_X1 #() 
AND3_X1_3_ (
  .A1({ S6160 }),
  .A2({ S25957[646] }),
  .A3({ S6163 }),
  .ZN({ S6164 })
);
AOI21_X1 #() 
AOI21_X1_10_ (
  .A({ S25957[646] }),
  .B1({ S6113 }),
  .B2({ S6108 }),
  .ZN({ S6166 })
);
OAI21_X1 #() 
OAI21_X1_51_ (
  .A({ S5530 }),
  .B1({ S6164 }),
  .B2({ S6166 }),
  .ZN({ S6167 })
);
OAI211_X1 #() 
OAI211_X1_9_ (
  .A({ S5465 }),
  .B({ S6124 }),
  .C1({ S6116 }),
  .C2({ S6119 }),
  .ZN({ S6168 })
);
NAND3_X1 #() 
NAND3_X1_31_ (
  .A1({ S6135 }),
  .A2({ S25957[646] }),
  .A3({ S6140 }),
  .ZN({ S6169 })
);
NAND3_X1 #() 
NAND3_X1_32_ (
  .A1({ S6168 }),
  .A2({ S6169 }),
  .A3({ S25957[647] }),
  .ZN({ S6170 })
);
AOI21_X1 #() 
AOI21_X1_11_ (
  .A({ S25957[842] }),
  .B1({ S6167 }),
  .B2({ S6170 }),
  .ZN({ S6171 })
);
OAI21_X1 #() 
OAI21_X1_52_ (
  .A({ S25957[682] }),
  .B1({ S6157 }),
  .B2({ S6171 }),
  .ZN({ S6172 })
);
NAND3_X1 #() 
NAND3_X1_33_ (
  .A1({ S6167 }),
  .A2({ S25957[842] }),
  .A3({ S6170 }),
  .ZN({ S6173 })
);
NAND3_X1 #() 
NAND3_X1_34_ (
  .A1({ S6156 }),
  .A2({ S6127 }),
  .A3({ S6102 }),
  .ZN({ S6174 })
);
NAND3_X1 #() 
NAND3_X1_35_ (
  .A1({ S6174 }),
  .A2({ S6100 }),
  .A3({ S6173 }),
  .ZN({ S6175 })
);
NAND3_X1 #() 
NAND3_X1_36_ (
  .A1({ S6172 }),
  .A2({ S25957[650] }),
  .A3({ S6175 }),
  .ZN({ S6177 })
);
NAND3_X1 #() 
NAND3_X1_37_ (
  .A1({ S6174 }),
  .A2({ S25957[682] }),
  .A3({ S6173 }),
  .ZN({ S6178 })
);
OAI21_X1 #() 
OAI21_X1_53_ (
  .A({ S6100 }),
  .B1({ S6157 }),
  .B2({ S6171 }),
  .ZN({ S6179 })
);
NAND3_X1 #() 
NAND3_X1_38_ (
  .A1({ S6179 }),
  .A2({ S4816 }),
  .A3({ S6178 }),
  .ZN({ S6180 })
);
NAND2_X1 #() 
NAND2_X1_55_ (
  .A1({ S6177 }),
  .A2({ S6180 }),
  .ZN({ S25957[522] })
);
NAND3_X1 #() 
NAND3_X1_39_ (
  .A1({ S4735 }),
  .A2({ S4736 }),
  .A3({ S25957[793] }),
  .ZN({ S6181 })
);
NAND3_X1 #() 
NAND3_X1_40_ (
  .A1({ S4729 }),
  .A2({ S4733 }),
  .A3({ S3527 }),
  .ZN({ S6182 })
);
NAND3_X1 #() 
NAND3_X1_41_ (
  .A1({ S25957[664] }),
  .A2({ S6181 }),
  .A3({ S6182 }),
  .ZN({ S6183 })
);
INV_X1 #() 
INV_X1_44_ (
  .A({ S6183 }),
  .ZN({ S10 })
);
NAND2_X1 #() 
NAND2_X1_56_ (
  .A1({ S2065 }),
  .A2({ S2044 }),
  .ZN({ S25957[856] })
);
NAND3_X1 #() 
NAND3_X1_42_ (
  .A1({ S4671 }),
  .A2({ S4645 }),
  .A3({ S25957[856] }),
  .ZN({ S6185 })
);
INV_X1 #() 
INV_X1_45_ (
  .A({ S25957[856] }),
  .ZN({ S6186 })
);
NAND3_X1 #() 
NAND3_X1_43_ (
  .A1({ S4674 }),
  .A2({ S4673 }),
  .A3({ S6186 }),
  .ZN({ S6187 })
);
NAND3_X1 #() 
NAND3_X1_44_ (
  .A1({ S6185 }),
  .A2({ S6187 }),
  .A3({ S1088 }),
  .ZN({ S6188 })
);
NAND3_X1 #() 
NAND3_X1_45_ (
  .A1({ S4674 }),
  .A2({ S4673 }),
  .A3({ S25957[856] }),
  .ZN({ S6189 })
);
NAND3_X1 #() 
NAND3_X1_46_ (
  .A1({ S4671 }),
  .A2({ S4645 }),
  .A3({ S6186 }),
  .ZN({ S6190 })
);
NAND3_X1 #() 
NAND3_X1_47_ (
  .A1({ S6189 }),
  .A2({ S6190 }),
  .A3({ S25957[920] }),
  .ZN({ S6191 })
);
NAND2_X1 #() 
NAND2_X1_57_ (
  .A1({ S6188 }),
  .A2({ S6191 }),
  .ZN({ S6192 })
);
NAND3_X1 #() 
NAND3_X1_48_ (
  .A1({ S4734 }),
  .A2({ S4737 }),
  .A3({ S6192 }),
  .ZN({ S11 })
);
NAND2_X1 #() 
NAND2_X1_58_ (
  .A1({ S3597 }),
  .A2({ S3600 }),
  .ZN({ S6193 })
);
INV_X1 #() 
INV_X1_46_ (
  .A({ S6193 }),
  .ZN({ S25957[679] })
);
NAND3_X1 #() 
NAND3_X1_49_ (
  .A1({ S4493 }),
  .A2({ S4489 }),
  .A3({ S25957[956] }),
  .ZN({ S6195 })
);
NAND3_X1 #() 
NAND3_X1_50_ (
  .A1({ S4499 }),
  .A2({ S4498 }),
  .A3({ S1942 }),
  .ZN({ S6196 })
);
NAND3_X1 #() 
NAND3_X1_51_ (
  .A1({ S6195 }),
  .A2({ S6196 }),
  .A3({ S3483 }),
  .ZN({ S6197 })
);
AOI21_X1 #() 
AOI21_X1_12_ (
  .A({ S1942 }),
  .B1({ S4499 }),
  .B2({ S4498 }),
  .ZN({ S6198 })
);
AOI21_X1 #() 
AOI21_X1_13_ (
  .A({ S25957[956] }),
  .B1({ S4493 }),
  .B2({ S4489 }),
  .ZN({ S6199 })
);
OAI21_X1 #() 
OAI21_X1_54_ (
  .A({ S25957[796] }),
  .B1({ S6198 }),
  .B2({ S6199 }),
  .ZN({ S6200 })
);
NAND2_X1 #() 
NAND2_X1_59_ (
  .A1({ S6200 }),
  .A2({ S6197 }),
  .ZN({ S6201 })
);
NAND3_X1 #() 
NAND3_X1_52_ (
  .A1({ S6181 }),
  .A2({ S6182 }),
  .A3({ S25957[666] }),
  .ZN({ S6202 })
);
NAND3_X1 #() 
NAND3_X1_53_ (
  .A1({ S6183 }),
  .A2({ S11 }),
  .A3({ S25957[666] }),
  .ZN({ S6203 })
);
OAI21_X1 #() 
OAI21_X1_55_ (
  .A({ S25957[922] }),
  .B1({ S4784 }),
  .B2({ S4787 }),
  .ZN({ S6205 })
);
NAND3_X1 #() 
NAND3_X1_54_ (
  .A1({ S4790 }),
  .A2({ S1033 }),
  .A3({ S4789 }),
  .ZN({ S6206 })
);
NAND2_X1 #() 
NAND2_X1_60_ (
  .A1({ S6205 }),
  .A2({ S6206 }),
  .ZN({ S6207 })
);
NAND3_X1 #() 
NAND3_X1_55_ (
  .A1({ S6207 }),
  .A2({ S6188 }),
  .A3({ S6191 }),
  .ZN({ S6208 })
);
NAND3_X1 #() 
NAND3_X1_56_ (
  .A1({ S6208 }),
  .A2({ S6181 }),
  .A3({ S6182 }),
  .ZN({ S6209 })
);
NAND3_X1 #() 
NAND3_X1_57_ (
  .A1({ S4676 }),
  .A2({ S6207 }),
  .A3({ S4679 }),
  .ZN({ S6210 })
);
NAND3_X1 #() 
NAND3_X1_58_ (
  .A1({ S6210 }),
  .A2({ S4734 }),
  .A3({ S4737 }),
  .ZN({ S6211 })
);
NAND2_X1 #() 
NAND2_X1_61_ (
  .A1({ S6211 }),
  .A2({ S6209 }),
  .ZN({ S6212 })
);
AOI21_X1 #() 
AOI21_X1_14_ (
  .A({ S3 }),
  .B1({ S6203 }),
  .B2({ S6212 }),
  .ZN({ S6213 })
);
NAND2_X1 #() 
NAND2_X1_62_ (
  .A1({ S6208 }),
  .A2({ S3 }),
  .ZN({ S6214 })
);
INV_X1 #() 
INV_X1_47_ (
  .A({ S6214 }),
  .ZN({ S6216 })
);
AOI21_X1 #() 
AOI21_X1_15_ (
  .A({ S6213 }),
  .B1({ S6202 }),
  .B2({ S6216 }),
  .ZN({ S6217 })
);
NOR2_X1 #() 
NOR2_X1_2_ (
  .A1({ S6217 }),
  .A2({ S6201 }),
  .ZN({ S6218 })
);
NAND3_X1 #() 
NAND3_X1_59_ (
  .A1({ S6183 }),
  .A2({ S11 }),
  .A3({ S6207 }),
  .ZN({ S6219 })
);
NAND3_X1 #() 
NAND3_X1_60_ (
  .A1({ S25957[664] }),
  .A2({ S4734 }),
  .A3({ S4737 }),
  .ZN({ S6220 })
);
NAND2_X1 #() 
NAND2_X1_63_ (
  .A1({ S6220 }),
  .A2({ S25957[666] }),
  .ZN({ S6221 })
);
NAND3_X1 #() 
NAND3_X1_61_ (
  .A1({ S6219 }),
  .A2({ S3 }),
  .A3({ S6221 }),
  .ZN({ S6222 })
);
NAND3_X1 #() 
NAND3_X1_62_ (
  .A1({ S4734 }),
  .A2({ S4737 }),
  .A3({ S6207 }),
  .ZN({ S6223 })
);
INV_X1 #() 
INV_X1_48_ (
  .A({ S6223 }),
  .ZN({ S6224 })
);
AOI21_X1 #() 
AOI21_X1_16_ (
  .A({ S25957[668] }),
  .B1({ S6224 }),
  .B2({ S25957[667] }),
  .ZN({ S6225 })
);
AOI21_X1 #() 
AOI21_X1_17_ (
  .A({ S6218 }),
  .B1({ S6222 }),
  .B2({ S6225 }),
  .ZN({ S6227 })
);
NAND3_X1 #() 
NAND3_X1_63_ (
  .A1({ S25957[666] }),
  .A2({ S6188 }),
  .A3({ S6191 }),
  .ZN({ S6228 })
);
INV_X1 #() 
INV_X1_49_ (
  .A({ S6228 }),
  .ZN({ S6229 })
);
NAND3_X1 #() 
NAND3_X1_64_ (
  .A1({ S3 }),
  .A2({ S6181 }),
  .A3({ S6182 }),
  .ZN({ S6230 })
);
NOR2_X1 #() 
NOR2_X1_3_ (
  .A1({ S6230 }),
  .A2({ S6229 }),
  .ZN({ S6231 })
);
NAND2_X1 #() 
NAND2_X1_64_ (
  .A1({ S6181 }),
  .A2({ S6182 }),
  .ZN({ S6232 })
);
OAI21_X1 #() 
OAI21_X1_56_ (
  .A({ S25957[667] }),
  .B1({ S6232 }),
  .B2({ S6229 }),
  .ZN({ S6233 })
);
NAND2_X1 #() 
NAND2_X1_65_ (
  .A1({ S6233 }),
  .A2({ S25957[668] }),
  .ZN({ S6234 })
);
NAND2_X1 #() 
NAND2_X1_66_ (
  .A1({ S6210 }),
  .A2({ S3 }),
  .ZN({ S6235 })
);
NAND2_X1 #() 
NAND2_X1_67_ (
  .A1({ S6230 }),
  .A2({ S6235 }),
  .ZN({ S6236 })
);
NAND2_X1 #() 
NAND2_X1_68_ (
  .A1({ S6183 }),
  .A2({ S6201 }),
  .ZN({ S6238 })
);
OAI221_X1 #() 
OAI221_X1_1_ (
  .A({ S25957[669] }),
  .B1({ S6236 }),
  .B2({ S6238 }),
  .C1({ S6234 }),
  .C2({ S6231 }),
  .ZN({ S6239 })
);
OAI21_X1 #() 
OAI21_X1_57_ (
  .A({ S6239 }),
  .B1({ S6227 }),
  .B2({ S25957[669] }),
  .ZN({ S6240 })
);
NAND3_X1 #() 
NAND3_X1_65_ (
  .A1({ S4734 }),
  .A2({ S4737 }),
  .A3({ S25957[666] }),
  .ZN({ S6241 })
);
NAND2_X1 #() 
NAND2_X1_69_ (
  .A1({ S6241 }),
  .A2({ S25957[667] }),
  .ZN({ S6242 })
);
NOR2_X1 #() 
NOR2_X1_4_ (
  .A1({ S6242 }),
  .A2({ S10 }),
  .ZN({ S6243 })
);
INV_X1 #() 
INV_X1_50_ (
  .A({ S6243 }),
  .ZN({ S6244 })
);
NAND3_X1 #() 
NAND3_X1_66_ (
  .A1({ S6181 }),
  .A2({ S6182 }),
  .A3({ S6192 }),
  .ZN({ S6245 })
);
NAND2_X1 #() 
NAND2_X1_70_ (
  .A1({ S6245 }),
  .A2({ S3 }),
  .ZN({ S6246 })
);
AOI21_X1 #() 
AOI21_X1_18_ (
  .A({ S6201 }),
  .B1({ S6244 }),
  .B2({ S6246 }),
  .ZN({ S6247 })
);
OAI211_X1 #() 
OAI211_X1_10_ (
  .A({ S6202 }),
  .B({ S6228 }),
  .C1({ S25957[665] }),
  .C2({ S6210 }),
  .ZN({ S6249 })
);
OAI21_X1 #() 
OAI21_X1_58_ (
  .A({ S6201 }),
  .B1({ S6220 }),
  .B2({ S3 }),
  .ZN({ S6250 })
);
NOR2_X1 #() 
NOR2_X1_5_ (
  .A1({ S6249 }),
  .A2({ S6250 }),
  .ZN({ S6251 })
);
NOR3_X1 #() 
NOR3_X1_3_ (
  .A1({ S6247 }),
  .A2({ S6251 }),
  .A3({ S25957[669] }),
  .ZN({ S6252 })
);
NAND2_X1 #() 
NAND2_X1_71_ (
  .A1({ S6192 }),
  .A2({ S25957[666] }),
  .ZN({ S6253 })
);
NAND4_X1 #() 
NAND4_X1_3_ (
  .A1({ S25957[664] }),
  .A2({ S4734 }),
  .A3({ S4737 }),
  .A4({ S6207 }),
  .ZN({ S6254 })
);
NAND3_X1 #() 
NAND3_X1_67_ (
  .A1({ S6254 }),
  .A2({ S25957[667] }),
  .A3({ S6253 }),
  .ZN({ S6255 })
);
NAND2_X1 #() 
NAND2_X1_72_ (
  .A1({ S25957[665] }),
  .A2({ S6210 }),
  .ZN({ S6256 })
);
OAI21_X1 #() 
OAI21_X1_59_ (
  .A({ S6255 }),
  .B1({ S25957[667] }),
  .B2({ S6256 }),
  .ZN({ S6257 })
);
NAND4_X1 #() 
NAND4_X1_4_ (
  .A1({ S6181 }),
  .A2({ S6182 }),
  .A3({ S6192 }),
  .A4({ S25957[666] }),
  .ZN({ S6258 })
);
NAND2_X1 #() 
NAND2_X1_73_ (
  .A1({ S6258 }),
  .A2({ S6220 }),
  .ZN({ S6260 })
);
NAND2_X1 #() 
NAND2_X1_74_ (
  .A1({ S6183 }),
  .A2({ S6253 }),
  .ZN({ S6261 })
);
NAND2_X1 #() 
NAND2_X1_75_ (
  .A1({ S6202 }),
  .A2({ S3 }),
  .ZN({ S6262 })
);
INV_X1 #() 
INV_X1_51_ (
  .A({ S6262 }),
  .ZN({ S6263 })
);
AOI22_X1 #() 
AOI22_X1_2_ (
  .A1({ S6263 }),
  .A2({ S6261 }),
  .B1({ S6260 }),
  .B2({ S25957[667] }),
  .ZN({ S6264 })
);
OAI21_X1 #() 
OAI21_X1_60_ (
  .A({ S25957[669] }),
  .B1({ S6264 }),
  .B2({ S25957[668] }),
  .ZN({ S6265 })
);
AOI21_X1 #() 
AOI21_X1_19_ (
  .A({ S6265 }),
  .B1({ S6257 }),
  .B2({ S25957[668] }),
  .ZN({ S6266 })
);
NOR3_X1 #() 
NOR3_X1_4_ (
  .A1({ S6252 }),
  .A2({ S6266 }),
  .A3({ S4354 }),
  .ZN({ S6267 })
);
AOI21_X1 #() 
AOI21_X1_20_ (
  .A({ S6267 }),
  .B1({ S6240 }),
  .B2({ S4354 }),
  .ZN({ S6268 })
);
NAND2_X1 #() 
NAND2_X1_76_ (
  .A1({ S6268 }),
  .A2({ S25957[671] }),
  .ZN({ S6269 })
);
INV_X1 #() 
INV_X1_52_ (
  .A({ S6241 }),
  .ZN({ S6271 })
);
AOI21_X1 #() 
AOI21_X1_21_ (
  .A({ S25957[667] }),
  .B1({ S6192 }),
  .B2({ S25957[666] }),
  .ZN({ S6272 })
);
INV_X1 #() 
INV_X1_53_ (
  .A({ S6272 }),
  .ZN({ S6273 })
);
NOR2_X1 #() 
NOR2_X1_6_ (
  .A1({ S6271 }),
  .A2({ S6273 }),
  .ZN({ S6274 })
);
NAND2_X1 #() 
NAND2_X1_77_ (
  .A1({ S6254 }),
  .A2({ S6202 }),
  .ZN({ S6275 })
);
NAND2_X1 #() 
NAND2_X1_78_ (
  .A1({ S6275 }),
  .A2({ S25957[667] }),
  .ZN({ S6276 })
);
NAND2_X1 #() 
NAND2_X1_79_ (
  .A1({ S6276 }),
  .A2({ S6201 }),
  .ZN({ S6277 })
);
AOI21_X1 #() 
AOI21_X1_22_ (
  .A({ S6207 }),
  .B1({ S4596 }),
  .B2({ S4593 }),
  .ZN({ S6278 })
);
AOI21_X1 #() 
AOI21_X1_23_ (
  .A({ S6201 }),
  .B1({ S25957[665] }),
  .B2({ S6278 }),
  .ZN({ S6279 })
);
AOI21_X1 #() 
AOI21_X1_24_ (
  .A({ S25957[667] }),
  .B1({ S6192 }),
  .B2({ S6207 }),
  .ZN({ S6280 })
);
NAND2_X1 #() 
NAND2_X1_80_ (
  .A1({ S6258 }),
  .A2({ S6280 }),
  .ZN({ S6282 })
);
NAND3_X1 #() 
NAND3_X1_68_ (
  .A1({ S6183 }),
  .A2({ S25957[667] }),
  .A3({ S6253 }),
  .ZN({ S6283 })
);
NAND3_X1 #() 
NAND3_X1_69_ (
  .A1({ S6279 }),
  .A2({ S6282 }),
  .A3({ S6283 }),
  .ZN({ S6284 })
);
OAI211_X1 #() 
OAI211_X1_11_ (
  .A({ S25957[669] }),
  .B({ S6284 }),
  .C1({ S6277 }),
  .C2({ S6274 }),
  .ZN({ S6285 })
);
NAND3_X1 #() 
NAND3_X1_70_ (
  .A1({ S6181 }),
  .A2({ S6182 }),
  .A3({ S6207 }),
  .ZN({ S6286 })
);
AND2_X1 #() 
AND2_X1_1_ (
  .A1({ S6228 }),
  .A2({ S25957[667] }),
  .ZN({ S6287 })
);
NAND2_X1 #() 
NAND2_X1_81_ (
  .A1({ S6287 }),
  .A2({ S6286 }),
  .ZN({ S6288 })
);
NAND4_X1 #() 
NAND4_X1_5_ (
  .A1({ S6286 }),
  .A2({ S6241 }),
  .A3({ S6253 }),
  .A4({ S6210 }),
  .ZN({ S6289 })
);
AOI21_X1 #() 
AOI21_X1_25_ (
  .A({ S25957[668] }),
  .B1({ S6289 }),
  .B2({ S3 }),
  .ZN({ S6290 })
);
NAND2_X1 #() 
NAND2_X1_82_ (
  .A1({ S6183 }),
  .A2({ S25957[666] }),
  .ZN({ S6291 })
);
AOI21_X1 #() 
AOI21_X1_26_ (
  .A({ S3 }),
  .B1({ S6212 }),
  .B2({ S6291 }),
  .ZN({ S6293 })
);
NAND3_X1 #() 
NAND3_X1_71_ (
  .A1({ S6220 }),
  .A2({ S6245 }),
  .A3({ S25957[666] }),
  .ZN({ S6294 })
);
AOI21_X1 #() 
AOI21_X1_27_ (
  .A({ S25957[667] }),
  .B1({ S6294 }),
  .B2({ S6210 }),
  .ZN({ S6295 })
);
NOR3_X1 #() 
NOR3_X1_5_ (
  .A1({ S6295 }),
  .A2({ S6293 }),
  .A3({ S6201 }),
  .ZN({ S6296 })
);
AOI21_X1 #() 
AOI21_X1_28_ (
  .A({ S6296 }),
  .B1({ S6290 }),
  .B2({ S6288 }),
  .ZN({ S6297 })
);
OAI21_X1 #() 
OAI21_X1_61_ (
  .A({ S6285 }),
  .B1({ S6297 }),
  .B2({ S25957[669] }),
  .ZN({ S6298 })
);
AOI21_X1 #() 
AOI21_X1_29_ (
  .A({ S6207 }),
  .B1({ S6220 }),
  .B2({ S6245 }),
  .ZN({ S6299 })
);
NOR2_X1 #() 
NOR2_X1_7_ (
  .A1({ S6192 }),
  .A2({ S25957[666] }),
  .ZN({ S6300 })
);
NAND2_X1 #() 
NAND2_X1_83_ (
  .A1({ S25957[665] }),
  .A2({ S6300 }),
  .ZN({ S6301 })
);
NAND2_X1 #() 
NAND2_X1_84_ (
  .A1({ S6301 }),
  .A2({ S3 }),
  .ZN({ S6302 })
);
OAI21_X1 #() 
OAI21_X1_62_ (
  .A({ S25957[668] }),
  .B1({ S6302 }),
  .B2({ S6299 }),
  .ZN({ S6304 })
);
AOI21_X1 #() 
AOI21_X1_30_ (
  .A({ S6304 }),
  .B1({ S6258 }),
  .B2({ S25957[667] }),
  .ZN({ S6305 })
);
INV_X1 #() 
INV_X1_54_ (
  .A({ S25957[669] }),
  .ZN({ S6306 })
);
INV_X1 #() 
INV_X1_55_ (
  .A({ S6278 }),
  .ZN({ S6307 })
);
NOR2_X1 #() 
NOR2_X1_8_ (
  .A1({ S10 }),
  .A2({ S6307 }),
  .ZN({ S6308 })
);
NAND2_X1 #() 
NAND2_X1_85_ (
  .A1({ S6202 }),
  .A2({ S6253 }),
  .ZN({ S6309 })
);
NAND3_X1 #() 
NAND3_X1_72_ (
  .A1({ S6309 }),
  .A2({ S3 }),
  .A3({ S6245 }),
  .ZN({ S6310 })
);
NAND2_X1 #() 
NAND2_X1_86_ (
  .A1({ S6310 }),
  .A2({ S6201 }),
  .ZN({ S6311 })
);
OAI21_X1 #() 
OAI21_X1_63_ (
  .A({ S6306 }),
  .B1({ S6311 }),
  .B2({ S6308 }),
  .ZN({ S6312 })
);
NOR2_X1 #() 
NOR2_X1_9_ (
  .A1({ S6305 }),
  .A2({ S6312 }),
  .ZN({ S6313 })
);
NAND3_X1 #() 
NAND3_X1_73_ (
  .A1({ S6220 }),
  .A2({ S6286 }),
  .A3({ S25957[667] }),
  .ZN({ S6315 })
);
NAND2_X1 #() 
NAND2_X1_87_ (
  .A1({ S6223 }),
  .A2({ S6210 }),
  .ZN({ S6316 })
);
OR2_X1 #() 
OR2_X1_1_ (
  .A1({ S6316 }),
  .A2({ S6262 }),
  .ZN({ S6317 })
);
AOI21_X1 #() 
AOI21_X1_31_ (
  .A({ S25957[668] }),
  .B1({ S6317 }),
  .B2({ S6315 }),
  .ZN({ S6318 })
);
NAND2_X1 #() 
NAND2_X1_88_ (
  .A1({ S6228 }),
  .A2({ S25957[667] }),
  .ZN({ S6319 })
);
NOR2_X1 #() 
NOR2_X1_10_ (
  .A1({ S6224 }),
  .A2({ S6319 }),
  .ZN({ S6320 })
);
OAI21_X1 #() 
OAI21_X1_64_ (
  .A({ S25957[668] }),
  .B1({ S25957[667] }),
  .B2({ S6192 }),
  .ZN({ S6321 })
);
OAI21_X1 #() 
OAI21_X1_65_ (
  .A({ S25957[669] }),
  .B1({ S6320 }),
  .B2({ S6321 }),
  .ZN({ S6322 })
);
OAI21_X1 #() 
OAI21_X1_66_ (
  .A({ S4354 }),
  .B1({ S6318 }),
  .B2({ S6322 }),
  .ZN({ S6323 })
);
OAI22_X1 #() 
OAI22_X1_1_ (
  .A1({ S6298 }),
  .A2({ S4354 }),
  .B1({ S6313 }),
  .B2({ S6323 }),
  .ZN({ S6324 })
);
OAI21_X1 #() 
OAI21_X1_67_ (
  .A({ S6269 }),
  .B1({ S6324 }),
  .B2({ S25957[671] }),
  .ZN({ S6326 })
);
NAND2_X1 #() 
NAND2_X1_89_ (
  .A1({ S6326 }),
  .A2({ S3595 }),
  .ZN({ S6327 })
);
NOR2_X1 #() 
NOR2_X1_11_ (
  .A1({ S6326 }),
  .A2({ S3595 }),
  .ZN({ S6328 })
);
INV_X1 #() 
INV_X1_56_ (
  .A({ S6328 }),
  .ZN({ S6329 })
);
NAND2_X1 #() 
NAND2_X1_90_ (
  .A1({ S6329 }),
  .A2({ S6327 }),
  .ZN({ S25957[583] })
);
NAND2_X1 #() 
NAND2_X1_91_ (
  .A1({ S25957[583] }),
  .A2({ S25957[679] }),
  .ZN({ S6330 })
);
NAND3_X1 #() 
NAND3_X1_74_ (
  .A1({ S6329 }),
  .A2({ S6193 }),
  .A3({ S6327 }),
  .ZN({ S6331 })
);
NAND2_X1 #() 
NAND2_X1_92_ (
  .A1({ S6330 }),
  .A2({ S6331 }),
  .ZN({ S6332 })
);
NAND2_X1 #() 
NAND2_X1_93_ (
  .A1({ S6332 }),
  .A2({ S5530 }),
  .ZN({ S6333 })
);
INV_X1 #() 
INV_X1_57_ (
  .A({ S6332 }),
  .ZN({ S25957[551] })
);
NAND2_X1 #() 
NAND2_X1_94_ (
  .A1({ S25957[551] }),
  .A2({ S25957[647] }),
  .ZN({ S6335 })
);
AND2_X1 #() 
AND2_X1_2_ (
  .A1({ S6335 }),
  .A2({ S6333 }),
  .ZN({ S25957[519] })
);
NAND2_X1 #() 
NAND2_X1_95_ (
  .A1({ S1213 }),
  .A2({ S1210 }),
  .ZN({ S6336 })
);
XNOR2_X1 #() 
XNOR2_X1_2_ (
  .A({ S6336 }),
  .B({ S25957[966] }),
  .ZN({ S25957[838] })
);
NAND2_X1 #() 
NAND2_X1_96_ (
  .A1({ S6203 }),
  .A2({ S3 }),
  .ZN({ S6337 })
);
AOI21_X1 #() 
AOI21_X1_32_ (
  .A({ S3 }),
  .B1({ S6221 }),
  .B2({ S6208 }),
  .ZN({ S6338 })
);
NOR2_X1 #() 
NOR2_X1_12_ (
  .A1({ S6338 }),
  .A2({ S25957[669] }),
  .ZN({ S6339 })
);
NAND2_X1 #() 
NAND2_X1_97_ (
  .A1({ S6339 }),
  .A2({ S6337 }),
  .ZN({ S6340 })
);
NOR2_X1 #() 
NOR2_X1_13_ (
  .A1({ S6228 }),
  .A2({ S3 }),
  .ZN({ S6341 })
);
INV_X1 #() 
INV_X1_58_ (
  .A({ S6341 }),
  .ZN({ S6342 })
);
NAND3_X1 #() 
NAND3_X1_75_ (
  .A1({ S6342 }),
  .A2({ S25957[669] }),
  .A3({ S6209 }),
  .ZN({ S6344 })
);
AOI21_X1 #() 
AOI21_X1_33_ (
  .A({ S25957[668] }),
  .B1({ S6340 }),
  .B2({ S6344 }),
  .ZN({ S6345 })
);
NAND3_X1 #() 
NAND3_X1_76_ (
  .A1({ S6223 }),
  .A2({ S3 }),
  .A3({ S6192 }),
  .ZN({ S6346 })
);
OAI211_X1 #() 
OAI211_X1_12_ (
  .A({ S6346 }),
  .B({ S6306 }),
  .C1({ S3 }),
  .C2({ S6286 }),
  .ZN({ S6347 })
);
NAND4_X1 #() 
NAND4_X1_6_ (
  .A1({ S25957[664] }),
  .A2({ S6181 }),
  .A3({ S6182 }),
  .A4({ S25957[666] }),
  .ZN({ S6348 })
);
NAND2_X1 #() 
NAND2_X1_98_ (
  .A1({ S6348 }),
  .A2({ S6210 }),
  .ZN({ S6349 })
);
NAND2_X1 #() 
NAND2_X1_99_ (
  .A1({ S11 }),
  .A2({ S6208 }),
  .ZN({ S6350 })
);
NAND2_X1 #() 
NAND2_X1_100_ (
  .A1({ S6350 }),
  .A2({ S25957[667] }),
  .ZN({ S6351 })
);
OAI21_X1 #() 
OAI21_X1_68_ (
  .A({ S6351 }),
  .B1({ S25957[667] }),
  .B2({ S6349 }),
  .ZN({ S6352 })
);
OAI21_X1 #() 
OAI21_X1_69_ (
  .A({ S6347 }),
  .B1({ S6352 }),
  .B2({ S6306 }),
  .ZN({ S6353 })
);
AOI21_X1 #() 
AOI21_X1_34_ (
  .A({ S6345 }),
  .B1({ S25957[668] }),
  .B2({ S6353 }),
  .ZN({ S6355 })
);
NAND3_X1 #() 
NAND3_X1_77_ (
  .A1({ S6232 }),
  .A2({ S6192 }),
  .A3({ S25957[666] }),
  .ZN({ S6356 })
);
NAND3_X1 #() 
NAND3_X1_78_ (
  .A1({ S6356 }),
  .A2({ S25957[667] }),
  .A3({ S6183 }),
  .ZN({ S6357 })
);
NAND3_X1 #() 
NAND3_X1_79_ (
  .A1({ S6357 }),
  .A2({ S25957[668] }),
  .A3({ S6214 }),
  .ZN({ S6358 })
);
INV_X1 #() 
INV_X1_59_ (
  .A({ S6286 }),
  .ZN({ S6359 })
);
OAI221_X1 #() 
OAI221_X1_2_ (
  .A({ S6201 }),
  .B1({ S6242 }),
  .B2({ S6359 }),
  .C1({ S6275 }),
  .C2({ S25957[667] }),
  .ZN({ S6360 })
);
NAND3_X1 #() 
NAND3_X1_80_ (
  .A1({ S6360 }),
  .A2({ S25957[669] }),
  .A3({ S6358 }),
  .ZN({ S6361 })
);
NAND4_X1 #() 
NAND4_X1_7_ (
  .A1({ S3 }),
  .A2({ S4734 }),
  .A3({ S4737 }),
  .A4({ S6207 }),
  .ZN({ S6362 })
);
OAI22_X1 #() 
OAI22_X1_2_ (
  .A1({ S6275 }),
  .A2({ S3 }),
  .B1({ S6192 }),
  .B2({ S6362 }),
  .ZN({ S6363 })
);
NAND3_X1 #() 
NAND3_X1_81_ (
  .A1({ S6258 }),
  .A2({ S6223 }),
  .A3({ S6208 }),
  .ZN({ S6364 })
);
NAND2_X1 #() 
NAND2_X1_101_ (
  .A1({ S6364 }),
  .A2({ S25957[667] }),
  .ZN({ S6366 })
);
AOI21_X1 #() 
AOI21_X1_35_ (
  .A({ S25957[669] }),
  .B1({ S6366 }),
  .B2({ S6201 }),
  .ZN({ S6367 })
);
OAI21_X1 #() 
OAI21_X1_70_ (
  .A({ S6367 }),
  .B1({ S6201 }),
  .B2({ S6363 }),
  .ZN({ S6368 })
);
NAND3_X1 #() 
NAND3_X1_82_ (
  .A1({ S6368 }),
  .A2({ S4354 }),
  .A3({ S6361 }),
  .ZN({ S6369 })
);
OAI21_X1 #() 
OAI21_X1_71_ (
  .A({ S6369 }),
  .B1({ S6355 }),
  .B2({ S4354 }),
  .ZN({ S6370 })
);
NAND2_X1 #() 
NAND2_X1_102_ (
  .A1({ S25957[665] }),
  .A2({ S6278 }),
  .ZN({ S6371 })
);
AOI21_X1 #() 
AOI21_X1_36_ (
  .A({ S25957[666] }),
  .B1({ S6191 }),
  .B2({ S6188 }),
  .ZN({ S6372 })
);
INV_X1 #() 
INV_X1_60_ (
  .A({ S6230 }),
  .ZN({ S6373 })
);
NAND2_X1 #() 
NAND2_X1_103_ (
  .A1({ S6373 }),
  .A2({ S6372 }),
  .ZN({ S6374 })
);
AND2_X1 #() 
AND2_X1_3_ (
  .A1({ S6374 }),
  .A2({ S6371 }),
  .ZN({ S6375 })
);
AOI21_X1 #() 
AOI21_X1_37_ (
  .A({ S6201 }),
  .B1({ S6375 }),
  .B2({ S6310 }),
  .ZN({ S6377 })
);
NAND2_X1 #() 
NAND2_X1_104_ (
  .A1({ S25957[665] }),
  .A2({ S6372 }),
  .ZN({ S6378 })
);
NAND2_X1 #() 
NAND2_X1_105_ (
  .A1({ S6378 }),
  .A2({ S25957[667] }),
  .ZN({ S6379 })
);
INV_X1 #() 
INV_X1_61_ (
  .A({ S6379 }),
  .ZN({ S6380 })
);
AOI21_X1 #() 
AOI21_X1_38_ (
  .A({ S25957[667] }),
  .B1({ S6348 }),
  .B2({ S11 }),
  .ZN({ S6381 })
);
AOI211_X1 #() 
AOI211_X1_1_ (
  .A({ S25957[668] }),
  .B({ S6381 }),
  .C1({ S6241 }),
  .C2({ S6380 }),
  .ZN({ S6382 })
);
OAI21_X1 #() 
OAI21_X1_72_ (
  .A({ S25957[669] }),
  .B1({ S6382 }),
  .B2({ S6377 }),
  .ZN({ S6383 })
);
NAND2_X1 #() 
NAND2_X1_106_ (
  .A1({ S6220 }),
  .A2({ S6207 }),
  .ZN({ S6384 })
);
OAI21_X1 #() 
OAI21_X1_73_ (
  .A({ S6233 }),
  .B1({ S6384 }),
  .B2({ S25957[667] }),
  .ZN({ S6385 })
);
INV_X1 #() 
INV_X1_62_ (
  .A({ S6212 }),
  .ZN({ S6386 })
);
NOR2_X1 #() 
NOR2_X1_14_ (
  .A1({ S6386 }),
  .A2({ S6273 }),
  .ZN({ S6388 })
);
AOI21_X1 #() 
AOI21_X1_39_ (
  .A({ S3 }),
  .B1({ S6258 }),
  .B2({ S6208 }),
  .ZN({ S6389 })
);
OAI21_X1 #() 
OAI21_X1_74_ (
  .A({ S6201 }),
  .B1({ S6388 }),
  .B2({ S6389 }),
  .ZN({ S6390 })
);
OAI21_X1 #() 
OAI21_X1_75_ (
  .A({ S6390 }),
  .B1({ S6201 }),
  .B2({ S6385 }),
  .ZN({ S6391 })
);
AOI21_X1 #() 
AOI21_X1_40_ (
  .A({ S25957[670] }),
  .B1({ S6391 }),
  .B2({ S6306 }),
  .ZN({ S6392 })
);
OAI21_X1 #() 
OAI21_X1_76_ (
  .A({ S25957[668] }),
  .B1({ S6388 }),
  .B2({ S6338 }),
  .ZN({ S6393 })
);
NAND4_X1 #() 
NAND4_X1_8_ (
  .A1({ S6241 }),
  .A2({ S6286 }),
  .A3({ S6272 }),
  .A4({ S6210 }),
  .ZN({ S6394 })
);
INV_X1 #() 
INV_X1_63_ (
  .A({ S6394 }),
  .ZN({ S6395 })
);
OAI21_X1 #() 
OAI21_X1_77_ (
  .A({ S25957[667] }),
  .B1({ S6232 }),
  .B2({ S6372 }),
  .ZN({ S6396 })
);
OAI21_X1 #() 
OAI21_X1_78_ (
  .A({ S6201 }),
  .B1({ S6396 }),
  .B2({ S6229 }),
  .ZN({ S6397 })
);
OAI21_X1 #() 
OAI21_X1_79_ (
  .A({ S6393 }),
  .B1({ S6395 }),
  .B2({ S6397 }),
  .ZN({ S6399 })
);
NAND2_X1 #() 
NAND2_X1_107_ (
  .A1({ S6399 }),
  .A2({ S6306 }),
  .ZN({ S6400 })
);
NAND2_X1 #() 
NAND2_X1_108_ (
  .A1({ S11 }),
  .A2({ S6207 }),
  .ZN({ S6401 })
);
AND2_X1 #() 
AND2_X1_4_ (
  .A1({ S6221 }),
  .A2({ S6401 }),
  .ZN({ S6402 })
);
NAND3_X1 #() 
NAND3_X1_83_ (
  .A1({ S6202 }),
  .A2({ S3 }),
  .A3({ S6228 }),
  .ZN({ S6403 })
);
OAI21_X1 #() 
OAI21_X1_80_ (
  .A({ S6403 }),
  .B1({ S6402 }),
  .B2({ S3 }),
  .ZN({ S6404 })
);
NAND2_X1 #() 
NAND2_X1_109_ (
  .A1({ S6244 }),
  .A2({ S6230 }),
  .ZN({ S6405 })
);
MUX2_X1 #() 
MUX2_X1_1_ (
  .A({ S6405 }),
  .B({ S6404 }),
  .S({ S25957[668] }),
  .Z({ S6406 })
);
AOI21_X1 #() 
AOI21_X1_41_ (
  .A({ S4354 }),
  .B1({ S6406 }),
  .B2({ S25957[669] }),
  .ZN({ S6407 })
);
AOI22_X1 #() 
AOI22_X1_3_ (
  .A1({ S6407 }),
  .A2({ S6400 }),
  .B1({ S6392 }),
  .B2({ S6383 }),
  .ZN({ S6408 })
);
NAND2_X1 #() 
NAND2_X1_110_ (
  .A1({ S6408 }),
  .A2({ S25957[671] }),
  .ZN({ S6410 })
);
OAI21_X1 #() 
OAI21_X1_81_ (
  .A({ S6410 }),
  .B1({ S25957[671] }),
  .B2({ S6370 }),
  .ZN({ S6411 })
);
OR2_X1 #() 
OR2_X1_2_ (
  .A1({ S6411 }),
  .A2({ S25957[838] }),
  .ZN({ S6412 })
);
NAND2_X1 #() 
NAND2_X1_111_ (
  .A1({ S6411 }),
  .A2({ S25957[838] }),
  .ZN({ S6413 })
);
AOI21_X1 #() 
AOI21_X1_42_ (
  .A({ S25957[774] }),
  .B1({ S6412 }),
  .B2({ S6413 }),
  .ZN({ S6414 })
);
NAND2_X1 #() 
NAND2_X1_112_ (
  .A1({ S6412 }),
  .A2({ S6413 }),
  .ZN({ S25957[582] })
);
NOR2_X1 #() 
NOR2_X1_15_ (
  .A1({ S25957[582] }),
  .A2({ S2900 }),
  .ZN({ S6415 })
);
NOR2_X1 #() 
NOR2_X1_16_ (
  .A1({ S6415 }),
  .A2({ S6414 }),
  .ZN({ S6416 })
);
INV_X1 #() 
INV_X1_64_ (
  .A({ S6416 }),
  .ZN({ S25957[518] })
);
NAND2_X1 #() 
NAND2_X1_113_ (
  .A1({ S24295 }),
  .A2({ S24296 }),
  .ZN({ S25957[933] })
);
XNOR2_X1 #() 
XNOR2_X1_3_ (
  .A({ S3682 }),
  .B({ S25957[933] }),
  .ZN({ S25957[805] })
);
NAND2_X1 #() 
NAND2_X1_114_ (
  .A1({ S3749 }),
  .A2({ S3750 }),
  .ZN({ S25957[709] })
);
XOR2_X1 #() 
XOR2_X1_1_ (
  .A({ S25957[709] }),
  .B({ S25957[805] }),
  .Z({ S25957[677] })
);
INV_X1 #() 
INV_X1_65_ (
  .A({ S25957[709] }),
  .ZN({ S6418 })
);
NAND2_X1 #() 
NAND2_X1_115_ (
  .A1({ S6349 }),
  .A2({ S25957[667] }),
  .ZN({ S6419 })
);
NAND3_X1 #() 
NAND3_X1_84_ (
  .A1({ S6378 }),
  .A2({ S3 }),
  .A3({ S6228 }),
  .ZN({ S6420 })
);
NAND2_X1 #() 
NAND2_X1_116_ (
  .A1({ S6419 }),
  .A2({ S6420 }),
  .ZN({ S6421 })
);
INV_X1 #() 
INV_X1_66_ (
  .A({ S6384 }),
  .ZN({ S6422 })
);
AOI21_X1 #() 
AOI21_X1_43_ (
  .A({ S6201 }),
  .B1({ S6422 }),
  .B2({ S25957[667] }),
  .ZN({ S6423 })
);
INV_X1 #() 
INV_X1_67_ (
  .A({ S6209 }),
  .ZN({ S6424 })
);
NAND2_X1 #() 
NAND2_X1_117_ (
  .A1({ S6424 }),
  .A2({ S6253 }),
  .ZN({ S6426 })
);
NAND3_X1 #() 
NAND3_X1_85_ (
  .A1({ S6426 }),
  .A2({ S3 }),
  .A3({ S6223 }),
  .ZN({ S6427 })
);
AOI22_X1 #() 
AOI22_X1_4_ (
  .A1({ S6421 }),
  .A2({ S6201 }),
  .B1({ S6423 }),
  .B2({ S6427 }),
  .ZN({ S6428 })
);
AOI21_X1 #() 
AOI21_X1_44_ (
  .A({ S4354 }),
  .B1({ S6428 }),
  .B2({ S6306 }),
  .ZN({ S6429 })
);
INV_X1 #() 
INV_X1_68_ (
  .A({ S6294 }),
  .ZN({ S6430 })
);
OAI211_X1 #() 
OAI211_X1_13_ (
  .A({ S6286 }),
  .B({ S3 }),
  .C1({ S25957[665] }),
  .C2({ S6300 }),
  .ZN({ S6431 })
);
OAI211_X1 #() 
OAI211_X1_14_ (
  .A({ S25957[668] }),
  .B({ S6431 }),
  .C1({ S6430 }),
  .C2({ S6379 }),
  .ZN({ S6432 })
);
NOR2_X1 #() 
NOR2_X1_17_ (
  .A1({ S25957[664] }),
  .A2({ S3 }),
  .ZN({ S6433 })
);
NAND3_X1 #() 
NAND3_X1_86_ (
  .A1({ S6245 }),
  .A2({ S3 }),
  .A3({ S6208 }),
  .ZN({ S6434 })
);
INV_X1 #() 
INV_X1_69_ (
  .A({ S6434 }),
  .ZN({ S6435 })
);
OAI21_X1 #() 
OAI21_X1_82_ (
  .A({ S6201 }),
  .B1({ S6435 }),
  .B2({ S6433 }),
  .ZN({ S6437 })
);
NAND3_X1 #() 
NAND3_X1_87_ (
  .A1({ S6432 }),
  .A2({ S25957[669] }),
  .A3({ S6437 }),
  .ZN({ S6438 })
);
NAND4_X1 #() 
NAND4_X1_9_ (
  .A1({ S6220 }),
  .A2({ S6245 }),
  .A3({ S6210 }),
  .A4({ S3 }),
  .ZN({ S6439 })
);
NAND3_X1 #() 
NAND3_X1_88_ (
  .A1({ S6294 }),
  .A2({ S25957[667] }),
  .A3({ S6254 }),
  .ZN({ S6440 })
);
AOI21_X1 #() 
AOI21_X1_45_ (
  .A({ S6201 }),
  .B1({ S6440 }),
  .B2({ S6439 }),
  .ZN({ S6441 })
);
NAND2_X1 #() 
NAND2_X1_118_ (
  .A1({ S6316 }),
  .A2({ S6230 }),
  .ZN({ S6442 })
);
AOI21_X1 #() 
AOI21_X1_46_ (
  .A({ S6201 }),
  .B1({ S6442 }),
  .B2({ S6235 }),
  .ZN({ S6443 })
);
NAND2_X1 #() 
NAND2_X1_119_ (
  .A1({ S6201 }),
  .A2({ S6319 }),
  .ZN({ S6444 })
);
AOI21_X1 #() 
AOI21_X1_47_ (
  .A({ S6444 }),
  .B1({ S6426 }),
  .B2({ S3 }),
  .ZN({ S6445 })
);
OAI21_X1 #() 
OAI21_X1_83_ (
  .A({ S25957[669] }),
  .B1({ S6443 }),
  .B2({ S6445 }),
  .ZN({ S6446 })
);
NOR2_X1 #() 
NOR2_X1_18_ (
  .A1({ S6348 }),
  .A2({ S25957[667] }),
  .ZN({ S6448 })
);
OAI21_X1 #() 
OAI21_X1_84_ (
  .A({ S6306 }),
  .B1({ S6448 }),
  .B2({ S6250 }),
  .ZN({ S6449 })
);
OAI21_X1 #() 
OAI21_X1_85_ (
  .A({ S6446 }),
  .B1({ S6449 }),
  .B2({ S6441 }),
  .ZN({ S6450 })
);
AOI22_X1 #() 
AOI22_X1_5_ (
  .A1({ S6429 }),
  .A2({ S6438 }),
  .B1({ S6450 }),
  .B2({ S4354 }),
  .ZN({ S6451 })
);
NOR2_X1 #() 
NOR2_X1_19_ (
  .A1({ S6311 }),
  .A2({ S6338 }),
  .ZN({ S6452 })
);
NAND3_X1 #() 
NAND3_X1_89_ (
  .A1({ S6384 }),
  .A2({ S3 }),
  .A3({ S6258 }),
  .ZN({ S6453 })
);
NAND2_X1 #() 
NAND2_X1_120_ (
  .A1({ S6433 }),
  .A2({ S6223 }),
  .ZN({ S6454 })
);
AOI21_X1 #() 
AOI21_X1_48_ (
  .A({ S6201 }),
  .B1({ S6453 }),
  .B2({ S6454 }),
  .ZN({ S6455 })
);
NAND3_X1 #() 
NAND3_X1_90_ (
  .A1({ S6228 }),
  .A2({ S4734 }),
  .A3({ S4737 }),
  .ZN({ S6456 })
);
NAND2_X1 #() 
NAND2_X1_121_ (
  .A1({ S6456 }),
  .A2({ S3 }),
  .ZN({ S6457 })
);
INV_X1 #() 
INV_X1_70_ (
  .A({ S6457 }),
  .ZN({ S6459 })
);
NAND3_X1 #() 
NAND3_X1_91_ (
  .A1({ S6396 }),
  .A2({ S6201 }),
  .A3({ S6342 }),
  .ZN({ S6460 })
);
OAI21_X1 #() 
OAI21_X1_86_ (
  .A({ S25957[669] }),
  .B1({ S6460 }),
  .B2({ S6459 }),
  .ZN({ S6461 })
);
NAND3_X1 #() 
NAND3_X1_92_ (
  .A1({ S6223 }),
  .A2({ S25957[667] }),
  .A3({ S6208 }),
  .ZN({ S6462 })
);
NAND3_X1 #() 
NAND3_X1_93_ (
  .A1({ S6245 }),
  .A2({ S3 }),
  .A3({ S25957[666] }),
  .ZN({ S6463 })
);
NAND3_X1 #() 
NAND3_X1_94_ (
  .A1({ S6462 }),
  .A2({ S6463 }),
  .A3({ S25957[668] }),
  .ZN({ S6464 })
);
NAND2_X1 #() 
NAND2_X1_122_ (
  .A1({ S6464 }),
  .A2({ S6306 }),
  .ZN({ S6465 })
);
OAI221_X1 #() 
OAI221_X1_3_ (
  .A({ S25957[670] }),
  .B1({ S6461 }),
  .B2({ S6455 }),
  .C1({ S6452 }),
  .C2({ S6465 }),
  .ZN({ S6466 })
);
AOI21_X1 #() 
AOI21_X1_49_ (
  .A({ S6278 }),
  .B1({ S6183 }),
  .B2({ S6210 }),
  .ZN({ S6467 })
);
OAI21_X1 #() 
OAI21_X1_87_ (
  .A({ S25957[668] }),
  .B1({ S6308 }),
  .B2({ S6467 }),
  .ZN({ S6468 })
);
NAND3_X1 #() 
NAND3_X1_95_ (
  .A1({ S6223 }),
  .A2({ S6245 }),
  .A3({ S3 }),
  .ZN({ S6470 })
);
AOI21_X1 #() 
AOI21_X1_50_ (
  .A({ S25957[668] }),
  .B1({ S6232 }),
  .B2({ S25957[667] }),
  .ZN({ S6471 })
);
AOI21_X1 #() 
AOI21_X1_51_ (
  .A({ S6306 }),
  .B1({ S6471 }),
  .B2({ S6470 }),
  .ZN({ S6472 })
);
NOR2_X1 #() 
NOR2_X1_20_ (
  .A1({ S25957[665] }),
  .A2({ S6210 }),
  .ZN({ S6473 })
);
OAI21_X1 #() 
OAI21_X1_88_ (
  .A({ S25957[667] }),
  .B1({ S6299 }),
  .B2({ S6473 }),
  .ZN({ S6474 })
);
NAND3_X1 #() 
NAND3_X1_96_ (
  .A1({ S6474 }),
  .A2({ S6201 }),
  .A3({ S6302 }),
  .ZN({ S6475 })
);
NAND2_X1 #() 
NAND2_X1_123_ (
  .A1({ S6216 }),
  .A2({ S6232 }),
  .ZN({ S6476 })
);
OAI21_X1 #() 
OAI21_X1_89_ (
  .A({ S6476 }),
  .B1({ S6219 }),
  .B2({ S3 }),
  .ZN({ S6477 })
);
AOI21_X1 #() 
AOI21_X1_52_ (
  .A({ S25957[669] }),
  .B1({ S6477 }),
  .B2({ S25957[668] }),
  .ZN({ S6478 })
);
AOI22_X1 #() 
AOI22_X1_6_ (
  .A1({ S6478 }),
  .A2({ S6475 }),
  .B1({ S6472 }),
  .B2({ S6468 }),
  .ZN({ S6479 })
);
NAND2_X1 #() 
NAND2_X1_124_ (
  .A1({ S6479 }),
  .A2({ S4354 }),
  .ZN({ S6481 })
);
NAND3_X1 #() 
NAND3_X1_97_ (
  .A1({ S6481 }),
  .A2({ S6466 }),
  .A3({ S25957[671] }),
  .ZN({ S6482 })
);
OAI211_X1 #() 
OAI211_X1_15_ (
  .A({ S6482 }),
  .B({ S25957[741] }),
  .C1({ S6451 }),
  .C2({ S25957[671] }),
  .ZN({ S6483 })
);
OAI22_X1 #() 
OAI22_X1_3_ (
  .A1({ S6452 }),
  .A2({ S6465 }),
  .B1({ S6461 }),
  .B2({ S6455 }),
  .ZN({ S6484 })
);
NAND2_X1 #() 
NAND2_X1_125_ (
  .A1({ S6484 }),
  .A2({ S25957[670] }),
  .ZN({ S6485 })
);
OAI211_X1 #() 
OAI211_X1_16_ (
  .A({ S6485 }),
  .B({ S25957[671] }),
  .C1({ S25957[670] }),
  .C2({ S6479 }),
  .ZN({ S6486 })
);
NAND2_X1 #() 
NAND2_X1_126_ (
  .A1({ S6421 }),
  .A2({ S6201 }),
  .ZN({ S6487 })
);
NAND2_X1 #() 
NAND2_X1_127_ (
  .A1({ S6423 }),
  .A2({ S6427 }),
  .ZN({ S6488 })
);
NAND3_X1 #() 
NAND3_X1_98_ (
  .A1({ S6487 }),
  .A2({ S6488 }),
  .A3({ S6306 }),
  .ZN({ S6489 })
);
NAND3_X1 #() 
NAND3_X1_99_ (
  .A1({ S6489 }),
  .A2({ S25957[670] }),
  .A3({ S6438 }),
  .ZN({ S6490 })
);
NAND2_X1 #() 
NAND2_X1_128_ (
  .A1({ S6450 }),
  .A2({ S4354 }),
  .ZN({ S6492 })
);
NAND3_X1 #() 
NAND3_X1_100_ (
  .A1({ S6492 }),
  .A2({ S4284 }),
  .A3({ S6490 }),
  .ZN({ S6493 })
);
NAND3_X1 #() 
NAND3_X1_101_ (
  .A1({ S6486 }),
  .A2({ S6493 }),
  .A3({ S3748 }),
  .ZN({ S6494 })
);
NAND3_X1 #() 
NAND3_X1_102_ (
  .A1({ S6483 }),
  .A2({ S6494 }),
  .A3({ S6418 }),
  .ZN({ S6495 })
);
OAI211_X1 #() 
OAI211_X1_17_ (
  .A({ S6482 }),
  .B({ S3748 }),
  .C1({ S6451 }),
  .C2({ S25957[671] }),
  .ZN({ S6496 })
);
NAND3_X1 #() 
NAND3_X1_103_ (
  .A1({ S6486 }),
  .A2({ S6493 }),
  .A3({ S25957[741] }),
  .ZN({ S6497 })
);
NAND3_X1 #() 
NAND3_X1_104_ (
  .A1({ S6496 }),
  .A2({ S6497 }),
  .A3({ S25957[709] }),
  .ZN({ S6498 })
);
NAND3_X1 #() 
NAND3_X1_105_ (
  .A1({ S6495 }),
  .A2({ S6498 }),
  .A3({ S25957[677] }),
  .ZN({ S6499 })
);
INV_X1 #() 
INV_X1_71_ (
  .A({ S25957[677] }),
  .ZN({ S6500 })
);
NAND3_X1 #() 
NAND3_X1_106_ (
  .A1({ S6483 }),
  .A2({ S6494 }),
  .A3({ S25957[709] }),
  .ZN({ S6501 })
);
NAND3_X1 #() 
NAND3_X1_107_ (
  .A1({ S6496 }),
  .A2({ S6497 }),
  .A3({ S6418 }),
  .ZN({ S6503 })
);
NAND3_X1 #() 
NAND3_X1_108_ (
  .A1({ S6501 }),
  .A2({ S6503 }),
  .A3({ S6500 }),
  .ZN({ S6504 })
);
NAND3_X1 #() 
NAND3_X1_109_ (
  .A1({ S6499 }),
  .A2({ S6504 }),
  .A3({ S25957[645] }),
  .ZN({ S6505 })
);
NAND3_X1 #() 
NAND3_X1_110_ (
  .A1({ S6501 }),
  .A2({ S6503 }),
  .A3({ S25957[677] }),
  .ZN({ S6506 })
);
NAND3_X1 #() 
NAND3_X1_111_ (
  .A1({ S6495 }),
  .A2({ S6498 }),
  .A3({ S6500 }),
  .ZN({ S6507 })
);
NAND3_X1 #() 
NAND3_X1_112_ (
  .A1({ S6506 }),
  .A2({ S6507 }),
  .A3({ S5494 }),
  .ZN({ S6508 })
);
NAND2_X1 #() 
NAND2_X1_129_ (
  .A1({ S6505 }),
  .A2({ S6508 }),
  .ZN({ S25957[517] })
);
NAND2_X1 #() 
NAND2_X1_130_ (
  .A1({ S3842 }),
  .A2({ S3845 }),
  .ZN({ S6509 })
);
INV_X1 #() 
INV_X1_72_ (
  .A({ S6509 }),
  .ZN({ S25957[676] })
);
NAND3_X1 #() 
NAND3_X1_113_ (
  .A1({ S6232 }),
  .A2({ S25957[667] }),
  .A3({ S6208 }),
  .ZN({ S6510 })
);
NAND3_X1 #() 
NAND3_X1_114_ (
  .A1({ S6470 }),
  .A2({ S25957[668] }),
  .A3({ S6510 }),
  .ZN({ S6512 })
);
NAND2_X1 #() 
NAND2_X1_131_ (
  .A1({ S6223 }),
  .A2({ S6272 }),
  .ZN({ S6513 })
);
NAND3_X1 #() 
NAND3_X1_115_ (
  .A1({ S6315 }),
  .A2({ S6201 }),
  .A3({ S6513 }),
  .ZN({ S6514 })
);
NAND2_X1 #() 
NAND2_X1_132_ (
  .A1({ S6512 }),
  .A2({ S6514 }),
  .ZN({ S6515 })
);
NAND2_X1 #() 
NAND2_X1_133_ (
  .A1({ S6356 }),
  .A2({ S3 }),
  .ZN({ S6516 })
);
NAND3_X1 #() 
NAND3_X1_116_ (
  .A1({ S6286 }),
  .A2({ S3 }),
  .A3({ S6192 }),
  .ZN({ S6517 })
);
NOR2_X1 #() 
NOR2_X1_21_ (
  .A1({ S6320 }),
  .A2({ S25957[668] }),
  .ZN({ S6518 })
);
AOI22_X1 #() 
AOI22_X1_7_ (
  .A1({ S6518 }),
  .A2({ S6517 }),
  .B1({ S6516 }),
  .B2({ S6423 }),
  .ZN({ S6519 })
);
NAND2_X1 #() 
NAND2_X1_134_ (
  .A1({ S6519 }),
  .A2({ S25957[669] }),
  .ZN({ S6520 })
);
OAI211_X1 #() 
OAI211_X1_18_ (
  .A({ S6520 }),
  .B({ S25957[670] }),
  .C1({ S25957[669] }),
  .C2({ S6515 }),
  .ZN({ S6521 })
);
INV_X1 #() 
INV_X1_73_ (
  .A({ S6220 }),
  .ZN({ S6523 })
);
NAND2_X1 #() 
NAND2_X1_135_ (
  .A1({ S6256 }),
  .A2({ S6456 }),
  .ZN({ S6524 })
);
NAND2_X1 #() 
NAND2_X1_136_ (
  .A1({ S6524 }),
  .A2({ S3 }),
  .ZN({ S6525 })
);
OAI211_X1 #() 
OAI211_X1_19_ (
  .A({ S6525 }),
  .B({ S25957[668] }),
  .C1({ S6523 }),
  .C2({ S6379 }),
  .ZN({ S6526 })
);
NAND2_X1 #() 
NAND2_X1_137_ (
  .A1({ S6241 }),
  .A2({ S6253 }),
  .ZN({ S6527 })
);
OAI21_X1 #() 
OAI21_X1_90_ (
  .A({ S3 }),
  .B1({ S6386 }),
  .B2({ S6527 }),
  .ZN({ S6528 })
);
AOI21_X1 #() 
AOI21_X1_53_ (
  .A({ S25957[668] }),
  .B1({ S6287 }),
  .B2({ S6211 }),
  .ZN({ S6529 })
);
NAND2_X1 #() 
NAND2_X1_138_ (
  .A1({ S6528 }),
  .A2({ S6529 }),
  .ZN({ S6530 })
);
NAND3_X1 #() 
NAND3_X1_117_ (
  .A1({ S6530 }),
  .A2({ S6526 }),
  .A3({ S25957[669] }),
  .ZN({ S6531 })
);
NAND2_X1 #() 
NAND2_X1_139_ (
  .A1({ S6245 }),
  .A2({ S6207 }),
  .ZN({ S6532 })
);
AOI21_X1 #() 
AOI21_X1_54_ (
  .A({ S25957[667] }),
  .B1({ S6532 }),
  .B2({ S6258 }),
  .ZN({ S6534 })
);
OAI21_X1 #() 
OAI21_X1_91_ (
  .A({ S6201 }),
  .B1({ S6319 }),
  .B2({ S25957[665] }),
  .ZN({ S6535 })
);
NAND3_X1 #() 
NAND3_X1_118_ (
  .A1({ S6301 }),
  .A2({ S3 }),
  .A3({ S6258 }),
  .ZN({ S6536 })
);
NAND3_X1 #() 
NAND3_X1_119_ (
  .A1({ S6287 }),
  .A2({ S6241 }),
  .A3({ S6286 }),
  .ZN({ S6537 })
);
NAND3_X1 #() 
NAND3_X1_120_ (
  .A1({ S6536 }),
  .A2({ S25957[668] }),
  .A3({ S6537 }),
  .ZN({ S6538 })
);
OAI211_X1 #() 
OAI211_X1_20_ (
  .A({ S6538 }),
  .B({ S6306 }),
  .C1({ S6534 }),
  .C2({ S6535 }),
  .ZN({ S6539 })
);
NAND3_X1 #() 
NAND3_X1_121_ (
  .A1({ S6539 }),
  .A2({ S6531 }),
  .A3({ S4354 }),
  .ZN({ S6540 })
);
NAND3_X1 #() 
NAND3_X1_122_ (
  .A1({ S6521 }),
  .A2({ S25957[671] }),
  .A3({ S6540 }),
  .ZN({ S6541 })
);
AND2_X1 #() 
AND2_X1_5_ (
  .A1({ S6207 }),
  .A2({ S138 }),
  .ZN({ S6542 })
);
OAI21_X1 #() 
OAI21_X1_92_ (
  .A({ S6463 }),
  .B1({ S6219 }),
  .B2({ S25957[667] }),
  .ZN({ S6543 })
);
AOI21_X1 #() 
AOI21_X1_55_ (
  .A({ S3 }),
  .B1({ S6348 }),
  .B2({ S6210 }),
  .ZN({ S6545 })
);
NOR2_X1 #() 
NOR2_X1_22_ (
  .A1({ S6545 }),
  .A2({ S25957[668] }),
  .ZN({ S6546 })
);
INV_X1 #() 
INV_X1_74_ (
  .A({ S6546 }),
  .ZN({ S6547 })
);
OAI22_X1 #() 
OAI22_X1_4_ (
  .A1({ S6547 }),
  .A2({ S6543 }),
  .B1({ S6542 }),
  .B2({ S6201 }),
  .ZN({ S6548 })
);
NOR2_X1 #() 
NOR2_X1_23_ (
  .A1({ S6403 }),
  .A2({ S6224 }),
  .ZN({ S6549 })
);
INV_X1 #() 
INV_X1_75_ (
  .A({ S6301 }),
  .ZN({ S6550 })
);
NOR2_X1 #() 
NOR2_X1_24_ (
  .A1({ S6550 }),
  .A2({ S6273 }),
  .ZN({ S6551 })
);
NAND2_X1 #() 
NAND2_X1_140_ (
  .A1({ S6307 }),
  .A2({ S6201 }),
  .ZN({ S6552 })
);
OAI221_X1 #() 
OAI221_X1_4_ (
  .A({ S6306 }),
  .B1({ S6549 }),
  .B2({ S6234 }),
  .C1({ S6551 }),
  .C2({ S6552 }),
  .ZN({ S6553 })
);
OAI211_X1 #() 
OAI211_X1_21_ (
  .A({ S25957[670] }),
  .B({ S6553 }),
  .C1({ S6548 }),
  .C2({ S6306 }),
  .ZN({ S6554 })
);
NAND2_X1 #() 
NAND2_X1_141_ (
  .A1({ S6287 }),
  .A2({ S11 }),
  .ZN({ S6556 })
);
NAND3_X1 #() 
NAND3_X1_123_ (
  .A1({ S6401 }),
  .A2({ S6356 }),
  .A3({ S3 }),
  .ZN({ S6557 })
);
NAND2_X1 #() 
NAND2_X1_142_ (
  .A1({ S6557 }),
  .A2({ S6556 }),
  .ZN({ S6558 })
);
NAND2_X1 #() 
NAND2_X1_143_ (
  .A1({ S6470 }),
  .A2({ S25957[668] }),
  .ZN({ S6559 })
);
AOI21_X1 #() 
AOI21_X1_56_ (
  .A({ S3 }),
  .B1({ S6254 }),
  .B2({ S6253 }),
  .ZN({ S6560 })
);
OAI21_X1 #() 
OAI21_X1_93_ (
  .A({ S6306 }),
  .B1({ S6559 }),
  .B2({ S6560 }),
  .ZN({ S6561 })
);
AOI21_X1 #() 
AOI21_X1_57_ (
  .A({ S6561 }),
  .B1({ S6558 }),
  .B2({ S6201 }),
  .ZN({ S6562 })
);
NOR2_X1 #() 
NOR2_X1_25_ (
  .A1({ S6219 }),
  .A2({ S3 }),
  .ZN({ S6563 })
);
NOR2_X1 #() 
NOR2_X1_26_ (
  .A1({ S6183 }),
  .A2({ S25957[667] }),
  .ZN({ S6564 })
);
OAI21_X1 #() 
OAI21_X1_94_ (
  .A({ S6201 }),
  .B1({ S6563 }),
  .B2({ S6564 }),
  .ZN({ S6565 })
);
NAND3_X1 #() 
NAND3_X1_124_ (
  .A1({ S6276 }),
  .A2({ S25957[668] }),
  .A3({ S6463 }),
  .ZN({ S6567 })
);
AND2_X1 #() 
AND2_X1_6_ (
  .A1({ S6567 }),
  .A2({ S25957[669] }),
  .ZN({ S6568 })
);
AOI21_X1 #() 
AOI21_X1_58_ (
  .A({ S6562 }),
  .B1({ S6565 }),
  .B2({ S6568 }),
  .ZN({ S6569 })
);
OAI21_X1 #() 
OAI21_X1_95_ (
  .A({ S6554 }),
  .B1({ S6569 }),
  .B2({ S25957[670] }),
  .ZN({ S6570 })
);
OR2_X1 #() 
OR2_X1_3_ (
  .A1({ S6570 }),
  .A2({ S25957[671] }),
  .ZN({ S6571 })
);
NAND3_X1 #() 
NAND3_X1_125_ (
  .A1({ S6571 }),
  .A2({ S25957[1028] }),
  .A3({ S6541 }),
  .ZN({ S6572 })
);
NAND2_X1 #() 
NAND2_X1_144_ (
  .A1({ S6571 }),
  .A2({ S6541 }),
  .ZN({ S6573 })
);
NAND2_X1 #() 
NAND2_X1_145_ (
  .A1({ S6573 }),
  .A2({ S23396 }),
  .ZN({ S6574 })
);
NAND2_X1 #() 
NAND2_X1_146_ (
  .A1({ S6574 }),
  .A2({ S6572 }),
  .ZN({ S6575 })
);
INV_X1 #() 
INV_X1_76_ (
  .A({ S6575 }),
  .ZN({ S25957[516] })
);
NOR2_X1 #() 
NOR2_X1_27_ (
  .A1({ S3923 }),
  .A2({ S3924 }),
  .ZN({ S25957[707] })
);
NAND2_X1 #() 
NAND2_X1_147_ (
  .A1({ S24442 }),
  .A2({ S24441 }),
  .ZN({ S25957[995] })
);
NAND2_X1 #() 
NAND2_X1_148_ (
  .A1({ S1405 }),
  .A2({ S1416 }),
  .ZN({ S6577 })
);
XNOR2_X1 #() 
XNOR2_X1_4_ (
  .A({ S6577 }),
  .B({ S25957[995] }),
  .ZN({ S25957[867] })
);
NAND2_X1 #() 
NAND2_X1_149_ (
  .A1({ S3905 }),
  .A2({ S3919 }),
  .ZN({ S6578 })
);
XNOR2_X1 #() 
XNOR2_X1_5_ (
  .A({ S6578 }),
  .B({ S25957[867] }),
  .ZN({ S25957[739] })
);
INV_X1 #() 
INV_X1_77_ (
  .A({ S25957[739] }),
  .ZN({ S6579 })
);
AOI21_X1 #() 
AOI21_X1_59_ (
  .A({ S25957[666] }),
  .B1({ S6220 }),
  .B2({ S6245 }),
  .ZN({ S6580 })
);
INV_X1 #() 
INV_X1_78_ (
  .A({ S6253 }),
  .ZN({ S6581 })
);
AOI21_X1 #() 
AOI21_X1_60_ (
  .A({ S3 }),
  .B1({ S6581 }),
  .B2({ S6232 }),
  .ZN({ S6582 })
);
INV_X1 #() 
INV_X1_79_ (
  .A({ S6582 }),
  .ZN({ S6584 })
);
NAND4_X1 #() 
NAND4_X1_10_ (
  .A1({ S25957[664] }),
  .A2({ S4734 }),
  .A3({ S4737 }),
  .A4({ S25957[666] }),
  .ZN({ S6585 })
);
AOI21_X1 #() 
AOI21_X1_61_ (
  .A({ S6201 }),
  .B1({ S6585 }),
  .B2({ S6280 }),
  .ZN({ S6586 })
);
OAI21_X1 #() 
OAI21_X1_96_ (
  .A({ S6586 }),
  .B1({ S6584 }),
  .B2({ S6580 }),
  .ZN({ S6587 })
);
NAND3_X1 #() 
NAND3_X1_126_ (
  .A1({ S6203 }),
  .A2({ S3 }),
  .A3({ S6223 }),
  .ZN({ S6588 })
);
NAND4_X1 #() 
NAND4_X1_11_ (
  .A1({ S25957[665] }),
  .A2({ S25957[667] }),
  .A3({ S6253 }),
  .A4({ S6208 }),
  .ZN({ S6589 })
);
NAND3_X1 #() 
NAND3_X1_127_ (
  .A1({ S6588 }),
  .A2({ S6201 }),
  .A3({ S6589 }),
  .ZN({ S6590 })
);
NAND3_X1 #() 
NAND3_X1_128_ (
  .A1({ S6590 }),
  .A2({ S6587 }),
  .A3({ S25957[669] }),
  .ZN({ S6591 })
);
AOI21_X1 #() 
AOI21_X1_62_ (
  .A({ S3 }),
  .B1({ S6211 }),
  .B2({ S6209 }),
  .ZN({ S6592 })
);
NAND2_X1 #() 
NAND2_X1_150_ (
  .A1({ S6513 }),
  .A2({ S25957[668] }),
  .ZN({ S6593 })
);
NAND3_X1 #() 
NAND3_X1_129_ (
  .A1({ S6348 }),
  .A2({ S25957[667] }),
  .A3({ S6456 }),
  .ZN({ S6595 })
);
OAI211_X1 #() 
OAI211_X1_22_ (
  .A({ S6595 }),
  .B({ S6201 }),
  .C1({ S6246 }),
  .C2({ S6229 }),
  .ZN({ S6596 })
);
OAI211_X1 #() 
OAI211_X1_23_ (
  .A({ S6596 }),
  .B({ S6306 }),
  .C1({ S6592 }),
  .C2({ S6593 }),
  .ZN({ S6597 })
);
NAND3_X1 #() 
NAND3_X1_130_ (
  .A1({ S6591 }),
  .A2({ S4354 }),
  .A3({ S6597 }),
  .ZN({ S6598 })
);
NAND3_X1 #() 
NAND3_X1_131_ (
  .A1({ S6294 }),
  .A2({ S3 }),
  .A3({ S6254 }),
  .ZN({ S6599 })
);
AOI21_X1 #() 
AOI21_X1_63_ (
  .A({ S6201 }),
  .B1({ S6599 }),
  .B2({ S6396 }),
  .ZN({ S6600 })
);
NOR2_X1 #() 
NOR2_X1_28_ (
  .A1({ S6552 }),
  .A2({ S6350 }),
  .ZN({ S6601 })
);
OAI21_X1 #() 
OAI21_X1_97_ (
  .A({ S6306 }),
  .B1({ S6600 }),
  .B2({ S6601 }),
  .ZN({ S6602 })
);
OAI21_X1 #() 
OAI21_X1_98_ (
  .A({ S6556 }),
  .B1({ S6260 }),
  .B2({ S25957[667] }),
  .ZN({ S6603 })
);
NAND2_X1 #() 
NAND2_X1_151_ (
  .A1({ S6603 }),
  .A2({ S25957[668] }),
  .ZN({ S6604 })
);
NAND3_X1 #() 
NAND3_X1_132_ (
  .A1({ S6211 }),
  .A2({ S3 }),
  .A3({ S6245 }),
  .ZN({ S6606 })
);
OAI211_X1 #() 
OAI211_X1_24_ (
  .A({ S6201 }),
  .B({ S6606 }),
  .C1({ S6524 }),
  .C2({ S3 }),
  .ZN({ S6607 })
);
NAND3_X1 #() 
NAND3_X1_133_ (
  .A1({ S6604 }),
  .A2({ S25957[669] }),
  .A3({ S6607 }),
  .ZN({ S6608 })
);
AND2_X1 #() 
AND2_X1_7_ (
  .A1({ S6602 }),
  .A2({ S6608 }),
  .ZN({ S6609 })
);
OAI211_X1 #() 
OAI211_X1_25_ (
  .A({ S25957[671] }),
  .B({ S6598 }),
  .C1({ S6609 }),
  .C2({ S4354 }),
  .ZN({ S6610 })
);
NAND2_X1 #() 
NAND2_X1_152_ (
  .A1({ S6433 }),
  .A2({ S6202 }),
  .ZN({ S6611 })
);
NAND3_X1 #() 
NAND3_X1_134_ (
  .A1({ S6220 }),
  .A2({ S6286 }),
  .A3({ S3 }),
  .ZN({ S6612 })
);
NAND3_X1 #() 
NAND3_X1_135_ (
  .A1({ S6612 }),
  .A2({ S6201 }),
  .A3({ S6611 }),
  .ZN({ S6613 })
);
OAI211_X1 #() 
OAI211_X1_26_ (
  .A({ S25957[669] }),
  .B({ S6613 }),
  .C1({ S6304 }),
  .C2({ S6338 }),
  .ZN({ S6614 })
);
AOI21_X1 #() 
AOI21_X1_64_ (
  .A({ S25957[667] }),
  .B1({ S6223 }),
  .B2({ S25957[664] }),
  .ZN({ S6615 })
);
AND2_X1 #() 
AND2_X1_8_ (
  .A1({ S6615 }),
  .A2({ S25957[668] }),
  .ZN({ S6617 })
);
AOI21_X1 #() 
AOI21_X1_65_ (
  .A({ S25957[668] }),
  .B1({ S6394 }),
  .B2({ S6255 }),
  .ZN({ S6618 })
);
OAI21_X1 #() 
OAI21_X1_99_ (
  .A({ S6306 }),
  .B1({ S6618 }),
  .B2({ S6617 }),
  .ZN({ S6619 })
);
AOI21_X1 #() 
AOI21_X1_66_ (
  .A({ S4354 }),
  .B1({ S6614 }),
  .B2({ S6619 }),
  .ZN({ S6620 })
);
INV_X1 #() 
INV_X1_80_ (
  .A({ S6620 }),
  .ZN({ S6621 })
);
OAI211_X1 #() 
OAI211_X1_27_ (
  .A({ S25957[667] }),
  .B({ S11 }),
  .C1({ S6183 }),
  .C2({ S25957[666] }),
  .ZN({ S6622 })
);
NAND3_X1 #() 
NAND3_X1_136_ (
  .A1({ S6622 }),
  .A2({ S6431 }),
  .A3({ S25957[668] }),
  .ZN({ S6623 })
);
NAND2_X1 #() 
NAND2_X1_153_ (
  .A1({ S6253 }),
  .A2({ S25957[667] }),
  .ZN({ S6624 })
);
OAI21_X1 #() 
OAI21_X1_100_ (
  .A({ S6201 }),
  .B1({ S6550 }),
  .B2({ S6624 }),
  .ZN({ S6625 })
);
OAI211_X1 #() 
OAI211_X1_28_ (
  .A({ S6306 }),
  .B({ S6623 }),
  .C1({ S6625 }),
  .C2({ S6295 }),
  .ZN({ S6626 })
);
INV_X1 #() 
INV_X1_81_ (
  .A({ S11 }),
  .ZN({ S6628 })
);
OAI211_X1 #() 
OAI211_X1_29_ (
  .A({ S25957[668] }),
  .B({ S25957[666] }),
  .C1({ S6564 }),
  .C2({ S6628 }),
  .ZN({ S6629 })
);
NAND4_X1 #() 
NAND4_X1_12_ (
  .A1({ S6242 }),
  .A2({ S6286 }),
  .A3({ S6201 }),
  .A4({ S25957[664] }),
  .ZN({ S6630 })
);
NAND3_X1 #() 
NAND3_X1_137_ (
  .A1({ S6629 }),
  .A2({ S25957[669] }),
  .A3({ S6630 }),
  .ZN({ S6631 })
);
AOI21_X1 #() 
AOI21_X1_67_ (
  .A({ S25957[670] }),
  .B1({ S6626 }),
  .B2({ S6631 }),
  .ZN({ S6632 })
);
INV_X1 #() 
INV_X1_82_ (
  .A({ S6632 }),
  .ZN({ S6633 })
);
NAND3_X1 #() 
NAND3_X1_138_ (
  .A1({ S6621 }),
  .A2({ S4284 }),
  .A3({ S6633 }),
  .ZN({ S6634 })
);
NAND3_X1 #() 
NAND3_X1_139_ (
  .A1({ S6610 }),
  .A2({ S6579 }),
  .A3({ S6634 }),
  .ZN({ S6635 })
);
OAI21_X1 #() 
OAI21_X1_101_ (
  .A({ S4284 }),
  .B1({ S6620 }),
  .B2({ S6632 }),
  .ZN({ S6636 })
);
AND3_X1 #() 
AND3_X1_4_ (
  .A1({ S6591 }),
  .A2({ S4354 }),
  .A3({ S6597 }),
  .ZN({ S6637 })
);
AOI21_X1 #() 
AOI21_X1_68_ (
  .A({ S4354 }),
  .B1({ S6602 }),
  .B2({ S6608 }),
  .ZN({ S6639 })
);
OAI21_X1 #() 
OAI21_X1_102_ (
  .A({ S25957[671] }),
  .B1({ S6639 }),
  .B2({ S6637 }),
  .ZN({ S6640 })
);
NAND3_X1 #() 
NAND3_X1_140_ (
  .A1({ S6640 }),
  .A2({ S6636 }),
  .A3({ S25957[739] }),
  .ZN({ S6641 })
);
AOI21_X1 #() 
AOI21_X1_69_ (
  .A({ S25957[707] }),
  .B1({ S6635 }),
  .B2({ S6641 }),
  .ZN({ S6642 })
);
INV_X1 #() 
INV_X1_83_ (
  .A({ S25957[707] }),
  .ZN({ S6643 })
);
NAND3_X1 #() 
NAND3_X1_141_ (
  .A1({ S6610 }),
  .A2({ S25957[739] }),
  .A3({ S6634 }),
  .ZN({ S6644 })
);
NAND3_X1 #() 
NAND3_X1_142_ (
  .A1({ S6640 }),
  .A2({ S6636 }),
  .A3({ S6579 }),
  .ZN({ S6645 })
);
AOI21_X1 #() 
AOI21_X1_70_ (
  .A({ S6643 }),
  .B1({ S6644 }),
  .B2({ S6645 }),
  .ZN({ S6646 })
);
OAI21_X1 #() 
OAI21_X1_103_ (
  .A({ S104 }),
  .B1({ S6642 }),
  .B2({ S6646 }),
  .ZN({ S6647 })
);
NAND3_X1 #() 
NAND3_X1_143_ (
  .A1({ S6644 }),
  .A2({ S6645 }),
  .A3({ S6643 }),
  .ZN({ S6648 })
);
NAND3_X1 #() 
NAND3_X1_144_ (
  .A1({ S6635 }),
  .A2({ S6641 }),
  .A3({ S25957[707] }),
  .ZN({ S6650 })
);
NAND3_X1 #() 
NAND3_X1_145_ (
  .A1({ S6648 }),
  .A2({ S6650 }),
  .A3({ S25957[771] }),
  .ZN({ S6651 })
);
NAND2_X1 #() 
NAND2_X1_154_ (
  .A1({ S6647 }),
  .A2({ S6651 }),
  .ZN({ S12 })
);
OAI21_X1 #() 
OAI21_X1_104_ (
  .A({ S25957[771] }),
  .B1({ S6642 }),
  .B2({ S6646 }),
  .ZN({ S6652 })
);
NAND3_X1 #() 
NAND3_X1_146_ (
  .A1({ S6648 }),
  .A2({ S6650 }),
  .A3({ S104 }),
  .ZN({ S6653 })
);
NAND2_X1 #() 
NAND2_X1_155_ (
  .A1({ S6652 }),
  .A2({ S6653 }),
  .ZN({ S25957[515] })
);
NAND2_X1 #() 
NAND2_X1_156_ (
  .A1({ S24544 }),
  .A2({ S24541 }),
  .ZN({ S25957[928] })
);
XOR2_X1 #() 
XOR2_X1_2_ (
  .A({ S25957[832] }),
  .B({ S25957[928] }),
  .Z({ S25957[800] })
);
INV_X1 #() 
INV_X1_84_ (
  .A({ S25957[800] }),
  .ZN({ S6654 })
);
NAND2_X1 #() 
NAND2_X1_157_ (
  .A1({ S4013 }),
  .A2({ S4017 }),
  .ZN({ S6655 })
);
INV_X1 #() 
INV_X1_85_ (
  .A({ S6655 }),
  .ZN({ S25957[704] })
);
NAND2_X1 #() 
NAND2_X1_158_ (
  .A1({ S25957[704] }),
  .A2({ S6654 }),
  .ZN({ S6657 })
);
NAND2_X1 #() 
NAND2_X1_159_ (
  .A1({ S6655 }),
  .A2({ S25957[800] }),
  .ZN({ S6658 })
);
NAND2_X1 #() 
NAND2_X1_160_ (
  .A1({ S6657 }),
  .A2({ S6658 }),
  .ZN({ S25957[672] })
);
NAND3_X1 #() 
NAND3_X1_147_ (
  .A1({ S6254 }),
  .A2({ S3 }),
  .A3({ S6209 }),
  .ZN({ S6659 })
);
AND3_X1 #() 
AND3_X1_5_ (
  .A1({ S6659 }),
  .A2({ S6255 }),
  .A3({ S6201 }),
  .ZN({ S6660 })
);
NAND2_X1 #() 
NAND2_X1_161_ (
  .A1({ S6245 }),
  .A2({ S6278 }),
  .ZN({ S6661 })
);
AOI21_X1 #() 
AOI21_X1_71_ (
  .A({ S6201 }),
  .B1({ S6557 }),
  .B2({ S6661 }),
  .ZN({ S6662 })
);
OAI21_X1 #() 
OAI21_X1_105_ (
  .A({ S25957[669] }),
  .B1({ S6662 }),
  .B2({ S6660 }),
  .ZN({ S6663 })
);
NAND3_X1 #() 
NAND3_X1_148_ (
  .A1({ S6220 }),
  .A2({ S6245 }),
  .A3({ S6278 }),
  .ZN({ S6664 })
);
NAND3_X1 #() 
NAND3_X1_149_ (
  .A1({ S6525 }),
  .A2({ S25957[668] }),
  .A3({ S6664 }),
  .ZN({ S6666 })
);
INV_X1 #() 
INV_X1_86_ (
  .A({ S6349 }),
  .ZN({ S6667 })
);
NOR2_X1 #() 
NOR2_X1_29_ (
  .A1({ S6280 }),
  .A2({ S25957[668] }),
  .ZN({ S6668 })
);
OAI21_X1 #() 
OAI21_X1_106_ (
  .A({ S6668 }),
  .B1({ S6667 }),
  .B2({ S6373 }),
  .ZN({ S6669 })
);
NAND3_X1 #() 
NAND3_X1_150_ (
  .A1({ S6666 }),
  .A2({ S6306 }),
  .A3({ S6669 }),
  .ZN({ S6670 })
);
NAND3_X1 #() 
NAND3_X1_151_ (
  .A1({ S6663 }),
  .A2({ S6670 }),
  .A3({ S25957[670] }),
  .ZN({ S6671 })
);
INV_X1 #() 
INV_X1_87_ (
  .A({ S6254 }),
  .ZN({ S6672 })
);
INV_X1 #() 
INV_X1_88_ (
  .A({ S6258 }),
  .ZN({ S6673 })
);
OAI21_X1 #() 
OAI21_X1_107_ (
  .A({ S3 }),
  .B1({ S6672 }),
  .B2({ S6673 }),
  .ZN({ S6674 })
);
NAND3_X1 #() 
NAND3_X1_152_ (
  .A1({ S6674 }),
  .A2({ S25957[668] }),
  .A3({ S6584 }),
  .ZN({ S6675 })
);
AOI21_X1 #() 
AOI21_X1_72_ (
  .A({ S6306 }),
  .B1({ S6516 }),
  .B2({ S6529 }),
  .ZN({ S6677 })
);
NAND2_X1 #() 
NAND2_X1_162_ (
  .A1({ S6675 }),
  .A2({ S6677 }),
  .ZN({ S6678 })
);
NAND4_X1 #() 
NAND4_X1_13_ (
  .A1({ S11 }),
  .A2({ S3 }),
  .A3({ S6210 }),
  .A4({ S6228 }),
  .ZN({ S6679 })
);
AOI21_X1 #() 
AOI21_X1_73_ (
  .A({ S25957[668] }),
  .B1({ S6679 }),
  .B2({ S6611 }),
  .ZN({ S6680 })
);
NAND2_X1 #() 
NAND2_X1_163_ (
  .A1({ S6371 }),
  .A2({ S25957[668] }),
  .ZN({ S6681 })
);
AOI21_X1 #() 
AOI21_X1_74_ (
  .A({ S6681 }),
  .B1({ S6580 }),
  .B2({ S3 }),
  .ZN({ S6682 })
);
OAI21_X1 #() 
OAI21_X1_108_ (
  .A({ S6306 }),
  .B1({ S6682 }),
  .B2({ S6680 }),
  .ZN({ S6683 })
);
NAND3_X1 #() 
NAND3_X1_153_ (
  .A1({ S6678 }),
  .A2({ S6683 }),
  .A3({ S4354 }),
  .ZN({ S6684 })
);
NAND3_X1 #() 
NAND3_X1_154_ (
  .A1({ S6671 }),
  .A2({ S25957[671] }),
  .A3({ S6684 }),
  .ZN({ S6685 })
);
NAND4_X1 #() 
NAND4_X1_14_ (
  .A1({ S6348 }),
  .A2({ S6456 }),
  .A3({ S25957[667] }),
  .A4({ S6210 }),
  .ZN({ S6686 })
);
AOI21_X1 #() 
AOI21_X1_75_ (
  .A({ S6201 }),
  .B1({ S6245 }),
  .B2({ S6272 }),
  .ZN({ S6688 })
);
AOI22_X1 #() 
AOI22_X1_8_ (
  .A1({ S6366 }),
  .A2({ S6668 }),
  .B1({ S6688 }),
  .B2({ S6686 }),
  .ZN({ S6689 })
);
NAND3_X1 #() 
NAND3_X1_155_ (
  .A1({ S6419 }),
  .A2({ S6201 }),
  .A3({ S6457 }),
  .ZN({ S6690 })
);
INV_X1 #() 
INV_X1_89_ (
  .A({ S6433 }),
  .ZN({ S6691 })
);
NAND4_X1 #() 
NAND4_X1_15_ (
  .A1({ S6691 }),
  .A2({ S6378 }),
  .A3({ S6241 }),
  .A4({ S25957[668] }),
  .ZN({ S6692 })
);
NAND3_X1 #() 
NAND3_X1_156_ (
  .A1({ S6690 }),
  .A2({ S6306 }),
  .A3({ S6692 }),
  .ZN({ S6693 })
);
OAI211_X1 #() 
OAI211_X1_30_ (
  .A({ S6693 }),
  .B({ S25957[670] }),
  .C1({ S6306 }),
  .C2({ S6689 }),
  .ZN({ S6694 })
);
NAND4_X1 #() 
NAND4_X1_16_ (
  .A1({ S6232 }),
  .A2({ S25957[667] }),
  .A3({ S6253 }),
  .A4({ S6208 }),
  .ZN({ S6695 })
);
NAND3_X1 #() 
NAND3_X1_157_ (
  .A1({ S6439 }),
  .A2({ S6201 }),
  .A3({ S6695 }),
  .ZN({ S6696 })
);
NAND3_X1 #() 
NAND3_X1_158_ (
  .A1({ S6556 }),
  .A2({ S6434 }),
  .A3({ S25957[668] }),
  .ZN({ S6697 })
);
NAND3_X1 #() 
NAND3_X1_159_ (
  .A1({ S6696 }),
  .A2({ S25957[669] }),
  .A3({ S6697 }),
  .ZN({ S6699 })
);
AOI21_X1 #() 
AOI21_X1_76_ (
  .A({ S25957[667] }),
  .B1({ S6348 }),
  .B2({ S6456 }),
  .ZN({ S6700 })
);
OAI21_X1 #() 
OAI21_X1_109_ (
  .A({ S25957[668] }),
  .B1({ S6700 }),
  .B2({ S6592 }),
  .ZN({ S6701 })
);
NAND3_X1 #() 
NAND3_X1_160_ (
  .A1({ S6348 }),
  .A2({ S25957[667] }),
  .A3({ S11 }),
  .ZN({ S6702 })
);
OAI211_X1 #() 
OAI211_X1_31_ (
  .A({ S6254 }),
  .B({ S3 }),
  .C1({ S25957[665] }),
  .C2({ S6253 }),
  .ZN({ S6703 })
);
NAND3_X1 #() 
NAND3_X1_161_ (
  .A1({ S6703 }),
  .A2({ S6201 }),
  .A3({ S6702 }),
  .ZN({ S6704 })
);
NAND2_X1 #() 
NAND2_X1_164_ (
  .A1({ S6701 }),
  .A2({ S6704 }),
  .ZN({ S6705 })
);
NAND2_X1 #() 
NAND2_X1_165_ (
  .A1({ S6705 }),
  .A2({ S6306 }),
  .ZN({ S6706 })
);
NAND3_X1 #() 
NAND3_X1_162_ (
  .A1({ S6706 }),
  .A2({ S4354 }),
  .A3({ S6699 }),
  .ZN({ S6707 })
);
NAND3_X1 #() 
NAND3_X1_163_ (
  .A1({ S6707 }),
  .A2({ S4284 }),
  .A3({ S6694 }),
  .ZN({ S6708 })
);
NAND3_X1 #() 
NAND3_X1_164_ (
  .A1({ S6708 }),
  .A2({ S6685 }),
  .A3({ S4014 }),
  .ZN({ S6710 })
);
NAND3_X1 #() 
NAND3_X1_165_ (
  .A1({ S6255 }),
  .A2({ S6659 }),
  .A3({ S6201 }),
  .ZN({ S6711 })
);
AOI22_X1 #() 
AOI22_X1_9_ (
  .A1({ S6249 }),
  .A2({ S3 }),
  .B1({ S6278 }),
  .B2({ S6245 }),
  .ZN({ S6712 })
);
OAI211_X1 #() 
OAI211_X1_32_ (
  .A({ S25957[669] }),
  .B({ S6711 }),
  .C1({ S6712 }),
  .C2({ S6201 }),
  .ZN({ S6713 })
);
AOI21_X1 #() 
AOI21_X1_77_ (
  .A({ S25957[667] }),
  .B1({ S6256 }),
  .B2({ S6456 }),
  .ZN({ S6714 })
);
AOI21_X1 #() 
AOI21_X1_78_ (
  .A({ S6307 }),
  .B1({ S6183 }),
  .B2({ S11 }),
  .ZN({ S6715 })
);
OAI21_X1 #() 
OAI21_X1_110_ (
  .A({ S25957[668] }),
  .B1({ S6714 }),
  .B2({ S6715 }),
  .ZN({ S6716 })
);
AOI21_X1 #() 
AOI21_X1_79_ (
  .A({ S25957[667] }),
  .B1({ S25957[665] }),
  .B2({ S6372 }),
  .ZN({ S6717 })
);
OAI21_X1 #() 
OAI21_X1_111_ (
  .A({ S6201 }),
  .B1({ S6545 }),
  .B2({ S6717 }),
  .ZN({ S6718 })
);
NAND3_X1 #() 
NAND3_X1_166_ (
  .A1({ S6716 }),
  .A2({ S6718 }),
  .A3({ S6306 }),
  .ZN({ S6719 })
);
NAND3_X1 #() 
NAND3_X1_167_ (
  .A1({ S6713 }),
  .A2({ S6719 }),
  .A3({ S25957[670] }),
  .ZN({ S6721 })
);
AND2_X1 #() 
AND2_X1_9_ (
  .A1({ S6679 }),
  .A2({ S6611 }),
  .ZN({ S6722 })
);
OAI21_X1 #() 
OAI21_X1_112_ (
  .A({ S6279 }),
  .B1({ S6219 }),
  .B2({ S25957[667] }),
  .ZN({ S6723 })
);
OAI211_X1 #() 
OAI211_X1_33_ (
  .A({ S6306 }),
  .B({ S6723 }),
  .C1({ S6722 }),
  .C2({ S25957[668] }),
  .ZN({ S6724 })
);
NAND3_X1 #() 
NAND3_X1_168_ (
  .A1({ S6202 }),
  .A2({ S3 }),
  .A3({ S6192 }),
  .ZN({ S6725 })
);
OAI211_X1 #() 
OAI211_X1_34_ (
  .A({ S25957[668] }),
  .B({ S6725 }),
  .C1({ S6582 }),
  .C2({ S6615 }),
  .ZN({ S6726 })
);
NAND2_X1 #() 
NAND2_X1_166_ (
  .A1({ S6273 }),
  .A2({ S6230 }),
  .ZN({ S6727 })
);
AOI21_X1 #() 
AOI21_X1_80_ (
  .A({ S6319 }),
  .B1({ S6210 }),
  .B2({ S6232 }),
  .ZN({ S6728 })
);
OAI21_X1 #() 
OAI21_X1_113_ (
  .A({ S6201 }),
  .B1({ S6727 }),
  .B2({ S6728 }),
  .ZN({ S6729 })
);
NAND3_X1 #() 
NAND3_X1_169_ (
  .A1({ S6726 }),
  .A2({ S6729 }),
  .A3({ S25957[669] }),
  .ZN({ S6730 })
);
NAND3_X1 #() 
NAND3_X1_170_ (
  .A1({ S6724 }),
  .A2({ S6730 }),
  .A3({ S4354 }),
  .ZN({ S6732 })
);
NAND3_X1 #() 
NAND3_X1_171_ (
  .A1({ S6721 }),
  .A2({ S6732 }),
  .A3({ S25957[671] }),
  .ZN({ S6733 })
);
NAND2_X1 #() 
NAND2_X1_167_ (
  .A1({ S6378 }),
  .A2({ S6241 }),
  .ZN({ S6734 })
);
OAI21_X1 #() 
OAI21_X1_114_ (
  .A({ S25957[668] }),
  .B1({ S6734 }),
  .B2({ S6433 }),
  .ZN({ S6735 })
);
OAI21_X1 #() 
OAI21_X1_115_ (
  .A({ S6201 }),
  .B1({ S6459 }),
  .B2({ S6545 }),
  .ZN({ S6736 })
);
NAND3_X1 #() 
NAND3_X1_172_ (
  .A1({ S6736 }),
  .A2({ S6735 }),
  .A3({ S6306 }),
  .ZN({ S6737 })
);
NAND2_X1 #() 
NAND2_X1_168_ (
  .A1({ S6686 }),
  .A2({ S6688 }),
  .ZN({ S6738 })
);
NAND2_X1 #() 
NAND2_X1_169_ (
  .A1({ S6366 }),
  .A2({ S6668 }),
  .ZN({ S6739 })
);
NAND3_X1 #() 
NAND3_X1_173_ (
  .A1({ S6739 }),
  .A2({ S25957[669] }),
  .A3({ S6738 }),
  .ZN({ S6740 })
);
NAND3_X1 #() 
NAND3_X1_174_ (
  .A1({ S6737 }),
  .A2({ S6740 }),
  .A3({ S25957[670] }),
  .ZN({ S6741 })
);
AND3_X1 #() 
AND3_X1_6_ (
  .A1({ S6696 }),
  .A2({ S25957[669] }),
  .A3({ S6697 }),
  .ZN({ S6743 })
);
AOI21_X1 #() 
AOI21_X1_81_ (
  .A({ S25957[669] }),
  .B1({ S6701 }),
  .B2({ S6704 }),
  .ZN({ S6744 })
);
OAI21_X1 #() 
OAI21_X1_116_ (
  .A({ S4354 }),
  .B1({ S6744 }),
  .B2({ S6743 }),
  .ZN({ S6745 })
);
NAND3_X1 #() 
NAND3_X1_175_ (
  .A1({ S6745 }),
  .A2({ S6741 }),
  .A3({ S4284 }),
  .ZN({ S6746 })
);
NAND3_X1 #() 
NAND3_X1_176_ (
  .A1({ S6746 }),
  .A2({ S6733 }),
  .A3({ S25957[832] }),
  .ZN({ S6747 })
);
NAND3_X1 #() 
NAND3_X1_177_ (
  .A1({ S6710 }),
  .A2({ S25957[672] }),
  .A3({ S6747 }),
  .ZN({ S6748 })
);
INV_X1 #() 
INV_X1_90_ (
  .A({ S25957[672] }),
  .ZN({ S6749 })
);
AOI21_X1 #() 
AOI21_X1_82_ (
  .A({ S25957[832] }),
  .B1({ S6746 }),
  .B2({ S6733 }),
  .ZN({ S6750 })
);
AOI21_X1 #() 
AOI21_X1_83_ (
  .A({ S4014 }),
  .B1({ S6708 }),
  .B2({ S6685 }),
  .ZN({ S6751 })
);
OAI21_X1 #() 
OAI21_X1_117_ (
  .A({ S6749 }),
  .B1({ S6751 }),
  .B2({ S6750 }),
  .ZN({ S6752 })
);
NAND3_X1 #() 
NAND3_X1_178_ (
  .A1({ S6752 }),
  .A2({ S25957[640] }),
  .A3({ S6748 }),
  .ZN({ S6754 })
);
NAND2_X1 #() 
NAND2_X1_170_ (
  .A1({ S4016 }),
  .A2({ S4015 }),
  .ZN({ S25957[736] })
);
NAND3_X1 #() 
NAND3_X1_179_ (
  .A1({ S6708 }),
  .A2({ S6685 }),
  .A3({ S25957[736] }),
  .ZN({ S6755 })
);
INV_X1 #() 
INV_X1_91_ (
  .A({ S25957[736] }),
  .ZN({ S6756 })
);
NAND3_X1 #() 
NAND3_X1_180_ (
  .A1({ S6746 }),
  .A2({ S6733 }),
  .A3({ S6756 }),
  .ZN({ S6757 })
);
NAND3_X1 #() 
NAND3_X1_181_ (
  .A1({ S6755 }),
  .A2({ S25957[800] }),
  .A3({ S6757 }),
  .ZN({ S6758 })
);
NAND3_X1 #() 
NAND3_X1_182_ (
  .A1({ S6708 }),
  .A2({ S6685 }),
  .A3({ S6756 }),
  .ZN({ S6759 })
);
NAND3_X1 #() 
NAND3_X1_183_ (
  .A1({ S6746 }),
  .A2({ S6733 }),
  .A3({ S25957[736] }),
  .ZN({ S6760 })
);
NAND3_X1 #() 
NAND3_X1_184_ (
  .A1({ S6759 }),
  .A2({ S6654 }),
  .A3({ S6760 }),
  .ZN({ S6761 })
);
NAND3_X1 #() 
NAND3_X1_185_ (
  .A1({ S6758 }),
  .A2({ S6761 }),
  .A3({ S5479 }),
  .ZN({ S6762 })
);
NAND2_X1 #() 
NAND2_X1_171_ (
  .A1({ S6754 }),
  .A2({ S6762 }),
  .ZN({ S25957[512] })
);
NAND2_X1 #() 
NAND2_X1_172_ (
  .A1({ S1551 }),
  .A2({ S1556 }),
  .ZN({ S25957[801] })
);
NOR2_X1 #() 
NOR2_X1_30_ (
  .A1({ S4060 }),
  .A2({ S4061 }),
  .ZN({ S25957[705] })
);
XOR2_X1 #() 
XOR2_X1_3_ (
  .A({ S25957[705] }),
  .B({ S25957[801] }),
  .Z({ S25957[673] })
);
INV_X1 #() 
INV_X1_92_ (
  .A({ S25957[673] }),
  .ZN({ S6764 })
);
NAND2_X1 #() 
NAND2_X1_173_ (
  .A1({ S24630 }),
  .A2({ S24603 }),
  .ZN({ S25957[993] })
);
XNOR2_X1 #() 
XNOR2_X1_6_ (
  .A({ S1554 }),
  .B({ S25957[993] }),
  .ZN({ S25957[865] })
);
NAND2_X1 #() 
NAND2_X1_174_ (
  .A1({ S4059 }),
  .A2({ S4040 }),
  .ZN({ S6765 })
);
XNOR2_X1 #() 
XNOR2_X1_7_ (
  .A({ S6765 }),
  .B({ S25957[865] }),
  .ZN({ S25957[737] })
);
NAND2_X1 #() 
NAND2_X1_175_ (
  .A1({ S6286 }),
  .A2({ S25957[667] }),
  .ZN({ S6766 })
);
NAND2_X1 #() 
NAND2_X1_176_ (
  .A1({ S6734 }),
  .A2({ S3 }),
  .ZN({ S6768 })
);
NAND3_X1 #() 
NAND3_X1_186_ (
  .A1({ S6768 }),
  .A2({ S25957[668] }),
  .A3({ S6766 }),
  .ZN({ S6769 })
);
OAI21_X1 #() 
OAI21_X1_118_ (
  .A({ S6201 }),
  .B1({ S6293 }),
  .B2({ S6534 }),
  .ZN({ S6770 })
);
AOI21_X1 #() 
AOI21_X1_84_ (
  .A({ S25957[669] }),
  .B1({ S6770 }),
  .B2({ S6769 }),
  .ZN({ S6771 })
);
NAND2_X1 #() 
NAND2_X1_177_ (
  .A1({ S6294 }),
  .A2({ S6210 }),
  .ZN({ S6772 })
);
NAND2_X1 #() 
NAND2_X1_178_ (
  .A1({ S6282 }),
  .A2({ S25957[668] }),
  .ZN({ S6773 })
);
AOI21_X1 #() 
AOI21_X1_85_ (
  .A({ S6773 }),
  .B1({ S6772 }),
  .B2({ S25957[667] }),
  .ZN({ S6774 })
);
NAND3_X1 #() 
NAND3_X1_187_ (
  .A1({ S6612 }),
  .A2({ S6462 }),
  .A3({ S6201 }),
  .ZN({ S6775 })
);
NAND2_X1 #() 
NAND2_X1_179_ (
  .A1({ S6775 }),
  .A2({ S25957[669] }),
  .ZN({ S6776 })
);
OAI21_X1 #() 
OAI21_X1_119_ (
  .A({ S4354 }),
  .B1({ S6774 }),
  .B2({ S6776 }),
  .ZN({ S6777 })
);
AOI21_X1 #() 
AOI21_X1_86_ (
  .A({ S25957[668] }),
  .B1({ S6258 }),
  .B2({ S3 }),
  .ZN({ S6779 })
);
NAND2_X1 #() 
NAND2_X1_180_ (
  .A1({ S6686 }),
  .A2({ S6779 }),
  .ZN({ S6780 })
);
AOI21_X1 #() 
AOI21_X1_87_ (
  .A({ S6201 }),
  .B1({ S6241 }),
  .B2({ S6272 }),
  .ZN({ S6781 })
);
NAND2_X1 #() 
NAND2_X1_181_ (
  .A1({ S6781 }),
  .A2({ S6396 }),
  .ZN({ S6782 })
);
NAND3_X1 #() 
NAND3_X1_188_ (
  .A1({ S6780 }),
  .A2({ S25957[669] }),
  .A3({ S6782 }),
  .ZN({ S6783 })
);
NAND2_X1 #() 
NAND2_X1_182_ (
  .A1({ S6725 }),
  .A2({ S25957[668] }),
  .ZN({ S6784 })
);
AOI21_X1 #() 
AOI21_X1_88_ (
  .A({ S6784 }),
  .B1({ S6380 }),
  .B2({ S6294 }),
  .ZN({ S6785 })
);
AOI22_X1 #() 
AOI22_X1_10_ (
  .A1({ S6230 }),
  .A2({ S6235 }),
  .B1({ S6223 }),
  .B2({ S25957[664] }),
  .ZN({ S6786 })
);
NAND2_X1 #() 
NAND2_X1_183_ (
  .A1({ S6283 }),
  .A2({ S6201 }),
  .ZN({ S6787 })
);
OAI21_X1 #() 
OAI21_X1_120_ (
  .A({ S6306 }),
  .B1({ S6787 }),
  .B2({ S6786 }),
  .ZN({ S6788 })
);
OAI211_X1 #() 
OAI211_X1_35_ (
  .A({ S6783 }),
  .B({ S25957[670] }),
  .C1({ S6785 }),
  .C2({ S6788 }),
  .ZN({ S6790 })
);
OAI211_X1 #() 
OAI211_X1_36_ (
  .A({ S25957[671] }),
  .B({ S6790 }),
  .C1({ S6771 }),
  .C2({ S6777 }),
  .ZN({ S6791 })
);
AOI21_X1 #() 
AOI21_X1_89_ (
  .A({ S6201 }),
  .B1({ S6517 }),
  .B2({ S6589 }),
  .ZN({ S6792 })
);
OAI21_X1 #() 
OAI21_X1_121_ (
  .A({ S25957[669] }),
  .B1({ S6290 }),
  .B2({ S6792 }),
  .ZN({ S6793 })
);
NAND3_X1 #() 
NAND3_X1_189_ (
  .A1({ S6233 }),
  .A2({ S25957[668] }),
  .A3({ S6513 }),
  .ZN({ S6794 })
);
NAND2_X1 #() 
NAND2_X1_184_ (
  .A1({ S6225 }),
  .A2({ S6394 }),
  .ZN({ S6795 })
);
NAND3_X1 #() 
NAND3_X1_190_ (
  .A1({ S6795 }),
  .A2({ S6306 }),
  .A3({ S6794 }),
  .ZN({ S6796 })
);
NAND3_X1 #() 
NAND3_X1_191_ (
  .A1({ S6793 }),
  .A2({ S6796 }),
  .A3({ S4354 }),
  .ZN({ S6797 })
);
NAND2_X1 #() 
NAND2_X1_185_ (
  .A1({ S6236 }),
  .A2({ S6348 }),
  .ZN({ S6798 })
);
NAND3_X1 #() 
NAND3_X1_192_ (
  .A1({ S6798 }),
  .A2({ S6686 }),
  .A3({ S25957[668] }),
  .ZN({ S6799 })
);
OAI211_X1 #() 
OAI211_X1_37_ (
  .A({ S6664 }),
  .B({ S6201 }),
  .C1({ S6214 }),
  .C2({ S6527 }),
  .ZN({ S6801 })
);
NAND3_X1 #() 
NAND3_X1_193_ (
  .A1({ S6799 }),
  .A2({ S6801 }),
  .A3({ S6306 }),
  .ZN({ S6802 })
);
NAND3_X1 #() 
NAND3_X1_194_ (
  .A1({ S6287 }),
  .A2({ S6245 }),
  .A3({ S6220 }),
  .ZN({ S6803 })
);
NAND2_X1 #() 
NAND2_X1_186_ (
  .A1({ S6356 }),
  .A2({ S6216 }),
  .ZN({ S6804 })
);
NAND3_X1 #() 
NAND3_X1_195_ (
  .A1({ S6804 }),
  .A2({ S6803 }),
  .A3({ S25957[668] }),
  .ZN({ S6805 })
);
AOI21_X1 #() 
AOI21_X1_90_ (
  .A({ S6229 }),
  .B1({ S6232 }),
  .B2({ S6372 }),
  .ZN({ S6806 })
);
AOI21_X1 #() 
AOI21_X1_91_ (
  .A({ S6306 }),
  .B1({ S6471 }),
  .B2({ S6806 }),
  .ZN({ S6807 })
);
AOI21_X1 #() 
AOI21_X1_92_ (
  .A({ S4354 }),
  .B1({ S6805 }),
  .B2({ S6807 }),
  .ZN({ S6808 })
);
NAND2_X1 #() 
NAND2_X1_187_ (
  .A1({ S6808 }),
  .A2({ S6802 }),
  .ZN({ S6809 })
);
NAND3_X1 #() 
NAND3_X1_196_ (
  .A1({ S6797 }),
  .A2({ S6809 }),
  .A3({ S4284 }),
  .ZN({ S6810 })
);
NAND3_X1 #() 
NAND3_X1_197_ (
  .A1({ S6791 }),
  .A2({ S6810 }),
  .A3({ S25957[737] }),
  .ZN({ S6812 })
);
INV_X1 #() 
INV_X1_93_ (
  .A({ S25957[737] }),
  .ZN({ S6813 })
);
NAND2_X1 #() 
NAND2_X1_188_ (
  .A1({ S6791 }),
  .A2({ S6810 }),
  .ZN({ S6814 })
);
NAND2_X1 #() 
NAND2_X1_189_ (
  .A1({ S6814 }),
  .A2({ S6813 }),
  .ZN({ S6815 })
);
NAND3_X1 #() 
NAND3_X1_198_ (
  .A1({ S6815 }),
  .A2({ S25957[705] }),
  .A3({ S6812 }),
  .ZN({ S6816 })
);
INV_X1 #() 
INV_X1_94_ (
  .A({ S25957[705] }),
  .ZN({ S6817 })
);
NAND3_X1 #() 
NAND3_X1_199_ (
  .A1({ S6791 }),
  .A2({ S6810 }),
  .A3({ S6813 }),
  .ZN({ S6818 })
);
NAND2_X1 #() 
NAND2_X1_190_ (
  .A1({ S6814 }),
  .A2({ S25957[737] }),
  .ZN({ S6819 })
);
NAND3_X1 #() 
NAND3_X1_200_ (
  .A1({ S6819 }),
  .A2({ S6817 }),
  .A3({ S6818 }),
  .ZN({ S6820 })
);
NAND3_X1 #() 
NAND3_X1_201_ (
  .A1({ S6820 }),
  .A2({ S6816 }),
  .A3({ S6764 }),
  .ZN({ S6821 })
);
NAND3_X1 #() 
NAND3_X1_202_ (
  .A1({ S6815 }),
  .A2({ S6817 }),
  .A3({ S6812 }),
  .ZN({ S6823 })
);
NAND3_X1 #() 
NAND3_X1_203_ (
  .A1({ S6819 }),
  .A2({ S25957[705] }),
  .A3({ S6818 }),
  .ZN({ S6824 })
);
NAND3_X1 #() 
NAND3_X1_204_ (
  .A1({ S6823 }),
  .A2({ S6824 }),
  .A3({ S25957[673] }),
  .ZN({ S6825 })
);
NAND3_X1 #() 
NAND3_X1_205_ (
  .A1({ S6821 }),
  .A2({ S6825 }),
  .A3({ S25957[641] }),
  .ZN({ S6826 })
);
NAND3_X1 #() 
NAND3_X1_206_ (
  .A1({ S6820 }),
  .A2({ S6816 }),
  .A3({ S25957[673] }),
  .ZN({ S6827 })
);
NAND3_X1 #() 
NAND3_X1_207_ (
  .A1({ S6823 }),
  .A2({ S6824 }),
  .A3({ S6764 }),
  .ZN({ S6828 })
);
NAND3_X1 #() 
NAND3_X1_208_ (
  .A1({ S6827 }),
  .A2({ S6828 }),
  .A3({ S5464 }),
  .ZN({ S6829 })
);
NAND2_X1 #() 
NAND2_X1_191_ (
  .A1({ S6826 }),
  .A2({ S6829 }),
  .ZN({ S25957[513] })
);
NOR2_X1 #() 
NOR2_X1_31_ (
  .A1({ S1613 }),
  .A2({ S1617 }),
  .ZN({ S6830 })
);
NOR2_X1 #() 
NOR2_X1_32_ (
  .A1({ S4130 }),
  .A2({ S4159 }),
  .ZN({ S6831 })
);
NOR2_X1 #() 
NOR2_X1_33_ (
  .A1({ S6831 }),
  .A2({ S6830 }),
  .ZN({ S6833 })
);
INV_X1 #() 
INV_X1_95_ (
  .A({ S6830 }),
  .ZN({ S25957[802] })
);
INV_X1 #() 
INV_X1_96_ (
  .A({ S6831 }),
  .ZN({ S25957[706] })
);
NOR2_X1 #() 
NOR2_X1_34_ (
  .A1({ S25957[706] }),
  .A2({ S25957[802] }),
  .ZN({ S6834 })
);
NOR2_X1 #() 
NOR2_X1_35_ (
  .A1({ S6834 }),
  .A2({ S6833 }),
  .ZN({ S25957[674] })
);
NAND2_X1 #() 
NAND2_X1_192_ (
  .A1({ S1612 }),
  .A2({ S1606 }),
  .ZN({ S25957[866] })
);
XNOR2_X1 #() 
XNOR2_X1_8_ (
  .A({ S25957[866] }),
  .B({ S4131 }),
  .ZN({ S25957[834] })
);
OAI211_X1 #() 
OAI211_X1_38_ (
  .A({ S25957[667] }),
  .B({ S6245 }),
  .C1({ S6220 }),
  .C2({ S6207 }),
  .ZN({ S6835 })
);
AOI21_X1 #() 
AOI21_X1_93_ (
  .A({ S25957[668] }),
  .B1({ S6835 }),
  .B2({ S6403 }),
  .ZN({ S6836 })
);
NAND3_X1 #() 
NAND3_X1_209_ (
  .A1({ S6223 }),
  .A2({ S25957[667] }),
  .A3({ S25957[664] }),
  .ZN({ S6837 })
);
AOI21_X1 #() 
AOI21_X1_94_ (
  .A({ S6201 }),
  .B1({ S6394 }),
  .B2({ S6837 }),
  .ZN({ S6839 })
);
OAI21_X1 #() 
OAI21_X1_122_ (
  .A({ S25957[669] }),
  .B1({ S6836 }),
  .B2({ S6839 }),
  .ZN({ S6840 })
);
NAND3_X1 #() 
NAND3_X1_210_ (
  .A1({ S6374 }),
  .A2({ S6201 }),
  .A3({ S6371 }),
  .ZN({ S6841 })
);
NAND2_X1 #() 
NAND2_X1_193_ (
  .A1({ S6424 }),
  .A2({ S25957[667] }),
  .ZN({ S6842 })
);
OAI211_X1 #() 
OAI211_X1_39_ (
  .A({ S6842 }),
  .B({ S25957[668] }),
  .C1({ S25957[667] }),
  .C2({ S6359 }),
  .ZN({ S6843 })
);
NAND3_X1 #() 
NAND3_X1_211_ (
  .A1({ S6843 }),
  .A2({ S6306 }),
  .A3({ S6841 }),
  .ZN({ S6844 })
);
NAND3_X1 #() 
NAND3_X1_212_ (
  .A1({ S6840 }),
  .A2({ S6844 }),
  .A3({ S4354 }),
  .ZN({ S6845 })
);
NAND3_X1 #() 
NAND3_X1_213_ (
  .A1({ S6241 }),
  .A2({ S25957[667] }),
  .A3({ S6228 }),
  .ZN({ S6846 })
);
OAI211_X1 #() 
OAI211_X1_40_ (
  .A({ S6262 }),
  .B({ S6201 }),
  .C1({ S6580 }),
  .C2({ S6846 }),
  .ZN({ S6847 })
);
OAI21_X1 #() 
OAI21_X1_123_ (
  .A({ S3 }),
  .B1({ S6672 }),
  .B2({ S6424 }),
  .ZN({ S6848 })
);
NAND3_X1 #() 
NAND3_X1_214_ (
  .A1({ S6848 }),
  .A2({ S25957[668] }),
  .A3({ S6288 }),
  .ZN({ S6850 })
);
NAND3_X1 #() 
NAND3_X1_215_ (
  .A1({ S6850 }),
  .A2({ S25957[669] }),
  .A3({ S6847 }),
  .ZN({ S6851 })
);
NAND3_X1 #() 
NAND3_X1_216_ (
  .A1({ S6219 }),
  .A2({ S6221 }),
  .A3({ S25957[667] }),
  .ZN({ S6852 })
);
NAND3_X1 #() 
NAND3_X1_217_ (
  .A1({ S6852 }),
  .A2({ S25957[668] }),
  .A3({ S6476 }),
  .ZN({ S6853 })
);
NAND3_X1 #() 
NAND3_X1_218_ (
  .A1({ S6315 }),
  .A2({ S6201 }),
  .A3({ S6362 }),
  .ZN({ S6854 })
);
NAND3_X1 #() 
NAND3_X1_219_ (
  .A1({ S6853 }),
  .A2({ S6306 }),
  .A3({ S6854 }),
  .ZN({ S6855 })
);
NAND3_X1 #() 
NAND3_X1_220_ (
  .A1({ S6855 }),
  .A2({ S6851 }),
  .A3({ S25957[670] }),
  .ZN({ S6856 })
);
NAND3_X1 #() 
NAND3_X1_221_ (
  .A1({ S6856 }),
  .A2({ S25957[671] }),
  .A3({ S6845 }),
  .ZN({ S6857 })
);
NAND2_X1 #() 
NAND2_X1_194_ (
  .A1({ S6806 }),
  .A2({ S25957[667] }),
  .ZN({ S6858 })
);
NAND3_X1 #() 
NAND3_X1_222_ (
  .A1({ S6588 }),
  .A2({ S25957[668] }),
  .A3({ S6858 }),
  .ZN({ S6859 })
);
NAND2_X1 #() 
NAND2_X1_195_ (
  .A1({ S6348 }),
  .A2({ S25957[667] }),
  .ZN({ S6861 })
);
OAI211_X1 #() 
OAI211_X1_41_ (
  .A({ S6374 }),
  .B({ S6201 }),
  .C1({ S6316 }),
  .C2({ S6861 }),
  .ZN({ S6862 })
);
NAND3_X1 #() 
NAND3_X1_223_ (
  .A1({ S6859 }),
  .A2({ S25957[669] }),
  .A3({ S6862 }),
  .ZN({ S6863 })
);
NAND3_X1 #() 
NAND3_X1_224_ (
  .A1({ S6366 }),
  .A2({ S6201 }),
  .A3({ S6659 }),
  .ZN({ S6864 })
);
NAND3_X1 #() 
NAND3_X1_225_ (
  .A1({ S6536 }),
  .A2({ S6842 }),
  .A3({ S25957[668] }),
  .ZN({ S6865 })
);
NAND3_X1 #() 
NAND3_X1_226_ (
  .A1({ S6864 }),
  .A2({ S6306 }),
  .A3({ S6865 }),
  .ZN({ S6866 })
);
AOI21_X1 #() 
AOI21_X1_95_ (
  .A({ S25957[670] }),
  .B1({ S6863 }),
  .B2({ S6866 }),
  .ZN({ S6867 })
);
NAND3_X1 #() 
NAND3_X1_227_ (
  .A1({ S6301 }),
  .A2({ S3 }),
  .A3({ S6585 }),
  .ZN({ S6868 })
);
OAI211_X1 #() 
OAI211_X1_42_ (
  .A({ S25957[667] }),
  .B({ S6228 }),
  .C1({ S6232 }),
  .C2({ S6210 }),
  .ZN({ S6869 })
);
AOI21_X1 #() 
AOI21_X1_96_ (
  .A({ S6201 }),
  .B1({ S6868 }),
  .B2({ S6869 }),
  .ZN({ S6870 })
);
NAND3_X1 #() 
NAND3_X1_228_ (
  .A1({ S6256 }),
  .A2({ S3 }),
  .A3({ S6456 }),
  .ZN({ S6872 })
);
AND3_X1 #() 
AND3_X1_7_ (
  .A1({ S6872 }),
  .A2({ S6842 }),
  .A3({ S6201 }),
  .ZN({ S6873 })
);
NOR3_X1 #() 
NOR3_X1_6_ (
  .A1({ S6873 }),
  .A2({ S6870 }),
  .A3({ S25957[669] }),
  .ZN({ S6874 })
);
NAND3_X1 #() 
NAND3_X1_229_ (
  .A1({ S6286 }),
  .A2({ S3 }),
  .A3({ S25957[664] }),
  .ZN({ S6875 })
);
NAND2_X1 #() 
NAND2_X1_196_ (
  .A1({ S6875 }),
  .A2({ S6201 }),
  .ZN({ S6876 })
);
OAI211_X1 #() 
OAI211_X1_43_ (
  .A({ S6181 }),
  .B({ S6182 }),
  .C1({ S6192 }),
  .C2({ S25957[667] }),
  .ZN({ S6877 })
);
NAND3_X1 #() 
NAND3_X1_230_ (
  .A1({ S6362 }),
  .A2({ S6877 }),
  .A3({ S6253 }),
  .ZN({ S6878 })
);
AOI21_X1 #() 
AOI21_X1_97_ (
  .A({ S6306 }),
  .B1({ S6878 }),
  .B2({ S25957[668] }),
  .ZN({ S6879 })
);
OAI21_X1 #() 
OAI21_X1_124_ (
  .A({ S6879 }),
  .B1({ S6213 }),
  .B2({ S6876 }),
  .ZN({ S6880 })
);
NAND2_X1 #() 
NAND2_X1_197_ (
  .A1({ S6880 }),
  .A2({ S25957[670] }),
  .ZN({ S6881 })
);
NOR2_X1 #() 
NOR2_X1_36_ (
  .A1({ S6881 }),
  .A2({ S6874 }),
  .ZN({ S6883 })
);
OAI21_X1 #() 
OAI21_X1_125_ (
  .A({ S4284 }),
  .B1({ S6883 }),
  .B2({ S6867 }),
  .ZN({ S6884 })
);
AOI21_X1 #() 
AOI21_X1_98_ (
  .A({ S25957[834] }),
  .B1({ S6884 }),
  .B2({ S6857 }),
  .ZN({ S6885 })
);
AND3_X1 #() 
AND3_X1_8_ (
  .A1({ S6884 }),
  .A2({ S6857 }),
  .A3({ S25957[834] }),
  .ZN({ S6886 })
);
OAI21_X1 #() 
OAI21_X1_126_ (
  .A({ S25957[674] }),
  .B1({ S6886 }),
  .B2({ S6885 }),
  .ZN({ S6887 })
);
INV_X1 #() 
INV_X1_97_ (
  .A({ S25957[674] }),
  .ZN({ S6888 })
);
INV_X1 #() 
INV_X1_98_ (
  .A({ S25957[834] }),
  .ZN({ S6889 })
);
AND3_X1 #() 
AND3_X1_9_ (
  .A1({ S6856 }),
  .A2({ S6845 }),
  .A3({ S25957[671] }),
  .ZN({ S6890 })
);
NAND2_X1 #() 
NAND2_X1_198_ (
  .A1({ S6863 }),
  .A2({ S6866 }),
  .ZN({ S6891 })
);
NAND2_X1 #() 
NAND2_X1_199_ (
  .A1({ S6891 }),
  .A2({ S4354 }),
  .ZN({ S6892 })
);
AND2_X1 #() 
AND2_X1_10_ (
  .A1({ S6868 }),
  .A2({ S6869 }),
  .ZN({ S6894 })
);
NAND3_X1 #() 
NAND3_X1_231_ (
  .A1({ S6872 }),
  .A2({ S6842 }),
  .A3({ S6201 }),
  .ZN({ S6895 })
);
OAI211_X1 #() 
OAI211_X1_44_ (
  .A({ S6895 }),
  .B({ S6306 }),
  .C1({ S6894 }),
  .C2({ S6201 }),
  .ZN({ S6896 })
);
NAND3_X1 #() 
NAND3_X1_232_ (
  .A1({ S6896 }),
  .A2({ S25957[670] }),
  .A3({ S6880 }),
  .ZN({ S6897 })
);
AOI21_X1 #() 
AOI21_X1_99_ (
  .A({ S25957[671] }),
  .B1({ S6892 }),
  .B2({ S6897 }),
  .ZN({ S6898 })
);
OAI21_X1 #() 
OAI21_X1_127_ (
  .A({ S6889 }),
  .B1({ S6898 }),
  .B2({ S6890 }),
  .ZN({ S6899 })
);
NAND3_X1 #() 
NAND3_X1_233_ (
  .A1({ S6884 }),
  .A2({ S25957[834] }),
  .A3({ S6857 }),
  .ZN({ S6900 })
);
NAND3_X1 #() 
NAND3_X1_234_ (
  .A1({ S6899 }),
  .A2({ S6888 }),
  .A3({ S6900 }),
  .ZN({ S6901 })
);
NAND3_X1 #() 
NAND3_X1_235_ (
  .A1({ S6887 }),
  .A2({ S25957[642] }),
  .A3({ S6901 }),
  .ZN({ S6902 })
);
OAI21_X1 #() 
OAI21_X1_128_ (
  .A({ S6888 }),
  .B1({ S6886 }),
  .B2({ S6885 }),
  .ZN({ S6903 })
);
NAND3_X1 #() 
NAND3_X1_236_ (
  .A1({ S6899 }),
  .A2({ S25957[674] }),
  .A3({ S6900 }),
  .ZN({ S6905 })
);
NAND3_X1 #() 
NAND3_X1_237_ (
  .A1({ S6903 }),
  .A2({ S5471 }),
  .A3({ S6905 }),
  .ZN({ S6906 })
);
NAND2_X1 #() 
NAND2_X1_200_ (
  .A1({ S6902 }),
  .A2({ S6906 }),
  .ZN({ S25957[514] })
);
NAND3_X1 #() 
NAND3_X1_238_ (
  .A1({ S25957[656] }),
  .A2({ S5357 }),
  .A3({ S5358 }),
  .ZN({ S6907 })
);
INV_X1 #() 
INV_X1_99_ (
  .A({ S6907 }),
  .ZN({ S13 })
);
OAI211_X1 #() 
OAI211_X1_45_ (
  .A({ S2746 }),
  .B({ S2752 }),
  .C1({ S2819 }),
  .C2({ S2818 }),
  .ZN({ S14 })
);
AOI21_X1 #() 
AOI21_X1_100_ (
  .A({ S25957[658] }),
  .B1({ S5357 }),
  .B2({ S5358 }),
  .ZN({ S6908 })
);
NAND2_X1 #() 
NAND2_X1_201_ (
  .A1({ S25957[659] }),
  .A2({ S6908 }),
  .ZN({ S6909 })
);
AND3_X1 #() 
AND3_X1_10_ (
  .A1({ S25957[658] }),
  .A2({ S2752 }),
  .A3({ S2746 }),
  .ZN({ S6910 })
);
NOR2_X1 #() 
NOR2_X1_37_ (
  .A1({ S25957[659] }),
  .A2({ S6910 }),
  .ZN({ S6911 })
);
NAND4_X1 #() 
NAND4_X1_17_ (
  .A1({ S25957[656] }),
  .A2({ S5357 }),
  .A3({ S5358 }),
  .A4({ S5458 }),
  .ZN({ S6913 })
);
AOI21_X1 #() 
AOI21_X1_101_ (
  .A({ S2749 }),
  .B1({ S2750 }),
  .B2({ S2751 }),
  .ZN({ S6914 })
);
AOI21_X1 #() 
AOI21_X1_102_ (
  .A({ S25957[784] }),
  .B1({ S2742 }),
  .B2({ S2745 }),
  .ZN({ S6915 })
);
OAI21_X1 #() 
OAI21_X1_129_ (
  .A({ S5458 }),
  .B1({ S6914 }),
  .B2({ S6915 }),
  .ZN({ S6916 })
);
NAND2_X1 #() 
NAND2_X1_202_ (
  .A1({ S6916 }),
  .A2({ S5359 }),
  .ZN({ S6917 })
);
NAND2_X1 #() 
NAND2_X1_203_ (
  .A1({ S6917 }),
  .A2({ S6913 }),
  .ZN({ S6918 })
);
NAND2_X1 #() 
NAND2_X1_204_ (
  .A1({ S6918 }),
  .A2({ S6911 }),
  .ZN({ S6919 })
);
AOI21_X1 #() 
AOI21_X1_103_ (
  .A({ S25957[660] }),
  .B1({ S6919 }),
  .B2({ S6909 }),
  .ZN({ S6920 })
);
NAND2_X1 #() 
NAND2_X1_205_ (
  .A1({ S25957[656] }),
  .A2({ S25957[658] }),
  .ZN({ S6921 })
);
NAND2_X1 #() 
NAND2_X1_206_ (
  .A1({ S110 }),
  .A2({ S25957[657] }),
  .ZN({ S6922 })
);
INV_X1 #() 
INV_X1_100_ (
  .A({ S6922 }),
  .ZN({ S6924 })
);
NAND3_X1 #() 
NAND3_X1_239_ (
  .A1({ S5359 }),
  .A2({ S2662 }),
  .A3({ S2665 }),
  .ZN({ S6925 })
);
OAI211_X1 #() 
OAI211_X1_46_ (
  .A({ S25957[660] }),
  .B({ S6925 }),
  .C1({ S110 }),
  .C2({ S6921 }),
  .ZN({ S6926 })
);
AOI21_X1 #() 
AOI21_X1_104_ (
  .A({ S6926 }),
  .B1({ S6924 }),
  .B2({ S6921 }),
  .ZN({ S6927 })
);
NAND3_X1 #() 
NAND3_X1_240_ (
  .A1({ S2596 }),
  .A2({ S2597 }),
  .A3({ S2524 }),
  .ZN({ S6928 })
);
NAND2_X1 #() 
NAND2_X1_207_ (
  .A1({ S25957[692] }),
  .A2({ S25957[788] }),
  .ZN({ S6929 })
);
NAND2_X1 #() 
NAND2_X1_208_ (
  .A1({ S6929 }),
  .A2({ S6928 }),
  .ZN({ S6930 })
);
NAND3_X1 #() 
NAND3_X1_241_ (
  .A1({ S5458 }),
  .A2({ S2746 }),
  .A3({ S2752 }),
  .ZN({ S6931 })
);
OAI21_X1 #() 
OAI21_X1_130_ (
  .A({ S110 }),
  .B1({ S6931 }),
  .B2({ S25957[657] }),
  .ZN({ S6932 })
);
NAND4_X1 #() 
NAND4_X1_18_ (
  .A1({ S25957[657] }),
  .A2({ S25957[656] }),
  .A3({ S2665 }),
  .A4({ S2662 }),
  .ZN({ S6933 })
);
NAND3_X1 #() 
NAND3_X1_242_ (
  .A1({ S6932 }),
  .A2({ S6930 }),
  .A3({ S6933 }),
  .ZN({ S6935 })
);
NAND2_X1 #() 
NAND2_X1_209_ (
  .A1({ S25957[661] }),
  .A2({ S6935 }),
  .ZN({ S6936 })
);
NAND3_X1 #() 
NAND3_X1_243_ (
  .A1({ S6907 }),
  .A2({ S25957[658] }),
  .A3({ S14 }),
  .ZN({ S6937 })
);
NAND2_X1 #() 
NAND2_X1_210_ (
  .A1({ S5359 }),
  .A2({ S25957[656] }),
  .ZN({ S6938 })
);
OAI21_X1 #() 
OAI21_X1_131_ (
  .A({ S5458 }),
  .B1({ S2819 }),
  .B2({ S2818 }),
  .ZN({ S6939 })
);
NAND2_X1 #() 
NAND2_X1_211_ (
  .A1({ S6916 }),
  .A2({ S6939 }),
  .ZN({ S6940 })
);
NAND2_X1 #() 
NAND2_X1_212_ (
  .A1({ S6940 }),
  .A2({ S6938 }),
  .ZN({ S6941 })
);
AOI21_X1 #() 
AOI21_X1_105_ (
  .A({ S110 }),
  .B1({ S6941 }),
  .B2({ S6937 }),
  .ZN({ S6942 })
);
NAND3_X1 #() 
NAND3_X1_244_ (
  .A1({ S5357 }),
  .A2({ S5358 }),
  .A3({ S25957[658] }),
  .ZN({ S6943 })
);
INV_X1 #() 
INV_X1_101_ (
  .A({ S6943 }),
  .ZN({ S6944 })
);
NAND2_X1 #() 
NAND2_X1_213_ (
  .A1({ S6916 }),
  .A2({ S110 }),
  .ZN({ S6946 })
);
OAI21_X1 #() 
OAI21_X1_132_ (
  .A({ S25957[660] }),
  .B1({ S6946 }),
  .B2({ S6944 }),
  .ZN({ S6947 })
);
OAI21_X1 #() 
OAI21_X1_133_ (
  .A({ S4995 }),
  .B1({ S6942 }),
  .B2({ S6947 }),
  .ZN({ S6948 })
);
OAI22_X1 #() 
OAI22_X1_5_ (
  .A1({ S6948 }),
  .A2({ S6920 }),
  .B1({ S6927 }),
  .B2({ S6936 }),
  .ZN({ S6949 })
);
NOR2_X1 #() 
NOR2_X1_38_ (
  .A1({ S6949 }),
  .A2({ S25957[662] }),
  .ZN({ S6950 })
);
NAND2_X1 #() 
NAND2_X1_214_ (
  .A1({ S6910 }),
  .A2({ S5359 }),
  .ZN({ S6951 })
);
NAND2_X1 #() 
NAND2_X1_215_ (
  .A1({ S14 }),
  .A2({ S5458 }),
  .ZN({ S6952 })
);
NAND2_X1 #() 
NAND2_X1_216_ (
  .A1({ S6952 }),
  .A2({ S6951 }),
  .ZN({ S6953 })
);
AOI22_X1 #() 
AOI22_X1_11_ (
  .A1({ S5357 }),
  .A2({ S5358 }),
  .B1({ S2752 }),
  .B2({ S2746 }),
  .ZN({ S6954 })
);
NAND2_X1 #() 
NAND2_X1_217_ (
  .A1({ S25957[659] }),
  .A2({ S6954 }),
  .ZN({ S6955 })
);
AOI21_X1 #() 
AOI21_X1_106_ (
  .A({ S25957[660] }),
  .B1({ S6953 }),
  .B2({ S6955 }),
  .ZN({ S6957 })
);
NAND3_X1 #() 
NAND3_X1_245_ (
  .A1({ S6951 }),
  .A2({ S110 }),
  .A3({ S6913 }),
  .ZN({ S6958 })
);
NAND2_X1 #() 
NAND2_X1_218_ (
  .A1({ S6910 }),
  .A2({ S25957[657] }),
  .ZN({ S6959 })
);
NAND3_X1 #() 
NAND3_X1_246_ (
  .A1({ S6959 }),
  .A2({ S25957[659] }),
  .A3({ S6938 }),
  .ZN({ S6960 })
);
AOI21_X1 #() 
AOI21_X1_107_ (
  .A({ S25957[660] }),
  .B1({ S6958 }),
  .B2({ S6960 }),
  .ZN({ S6961 })
);
NAND2_X1 #() 
NAND2_X1_219_ (
  .A1({ S110 }),
  .A2({ S6931 }),
  .ZN({ S6962 })
);
NOR2_X1 #() 
NOR2_X1_39_ (
  .A1({ S6939 }),
  .A2({ S5282 }),
  .ZN({ S6963 })
);
NOR2_X1 #() 
NOR2_X1_40_ (
  .A1({ S6910 }),
  .A2({ S110 }),
  .ZN({ S6964 })
);
INV_X1 #() 
INV_X1_102_ (
  .A({ S6964 }),
  .ZN({ S6965 })
);
OAI22_X1 #() 
OAI22_X1_6_ (
  .A1({ S6963 }),
  .A2({ S6965 }),
  .B1({ S6962 }),
  .B2({ S5359 }),
  .ZN({ S6966 })
);
OAI21_X1 #() 
OAI21_X1_134_ (
  .A({ S25957[661] }),
  .B1({ S6966 }),
  .B2({ S6930 }),
  .ZN({ S6968 })
);
OAI21_X1 #() 
OAI21_X1_135_ (
  .A({ S25957[658] }),
  .B1({ S2819 }),
  .B2({ S2818 }),
  .ZN({ S6969 })
);
NAND2_X1 #() 
NAND2_X1_220_ (
  .A1({ S25957[659] }),
  .A2({ S6969 }),
  .ZN({ S6970 })
);
NOR2_X1 #() 
NOR2_X1_41_ (
  .A1({ S6970 }),
  .A2({ S13 }),
  .ZN({ S6971 })
);
NAND4_X1 #() 
NAND4_X1_19_ (
  .A1({ S5357 }),
  .A2({ S5358 }),
  .A3({ S2746 }),
  .A4({ S2752 }),
  .ZN({ S6972 })
);
INV_X1 #() 
INV_X1_103_ (
  .A({ S6972 }),
  .ZN({ S6973 })
);
OAI21_X1 #() 
OAI21_X1_136_ (
  .A({ S25957[660] }),
  .B1({ S6973 }),
  .B2({ S25957[659] }),
  .ZN({ S6974 })
);
OAI21_X1 #() 
OAI21_X1_137_ (
  .A({ S4995 }),
  .B1({ S6971 }),
  .B2({ S6974 }),
  .ZN({ S6975 })
);
OAI22_X1 #() 
OAI22_X1_7_ (
  .A1({ S6968 }),
  .A2({ S6961 }),
  .B1({ S6957 }),
  .B2({ S6975 }),
  .ZN({ S6976 })
);
OAI21_X1 #() 
OAI21_X1_138_ (
  .A({ S25957[663] }),
  .B1({ S6976 }),
  .B2({ S2444 }),
  .ZN({ S6977 })
);
NAND3_X1 #() 
NAND3_X1_247_ (
  .A1({ S5357 }),
  .A2({ S5458 }),
  .A3({ S5358 }),
  .ZN({ S6979 })
);
NAND2_X1 #() 
NAND2_X1_221_ (
  .A1({ S6938 }),
  .A2({ S6979 }),
  .ZN({ S6980 })
);
NOR2_X1 #() 
NOR2_X1_42_ (
  .A1({ S6980 }),
  .A2({ S110 }),
  .ZN({ S6981 })
);
AOI21_X1 #() 
AOI21_X1_108_ (
  .A({ S25957[659] }),
  .B1({ S6913 }),
  .B2({ S6969 }),
  .ZN({ S6982 })
);
OAI21_X1 #() 
OAI21_X1_139_ (
  .A({ S6930 }),
  .B1({ S6981 }),
  .B2({ S6982 }),
  .ZN({ S6983 })
);
AOI21_X1 #() 
AOI21_X1_109_ (
  .A({ S5458 }),
  .B1({ S2752 }),
  .B2({ S2746 }),
  .ZN({ S6984 })
);
NOR2_X1 #() 
NOR2_X1_43_ (
  .A1({ S6984 }),
  .A2({ S110 }),
  .ZN({ S6985 })
);
NAND2_X1 #() 
NAND2_X1_222_ (
  .A1({ S6985 }),
  .A2({ S6939 }),
  .ZN({ S6986 })
);
NAND2_X1 #() 
NAND2_X1_223_ (
  .A1({ S110 }),
  .A2({ S25957[656] }),
  .ZN({ S6987 })
);
NAND3_X1 #() 
NAND3_X1_248_ (
  .A1({ S6986 }),
  .A2({ S25957[660] }),
  .A3({ S6987 }),
  .ZN({ S6988 })
);
NAND3_X1 #() 
NAND3_X1_249_ (
  .A1({ S6983 }),
  .A2({ S2444 }),
  .A3({ S6988 }),
  .ZN({ S6990 })
);
NOR2_X1 #() 
NOR2_X1_44_ (
  .A1({ S6979 }),
  .A2({ S5282 }),
  .ZN({ S6991 })
);
NAND2_X1 #() 
NAND2_X1_224_ (
  .A1({ S6951 }),
  .A2({ S25957[659] }),
  .ZN({ S6992 })
);
OAI21_X1 #() 
OAI21_X1_140_ (
  .A({ S5282 }),
  .B1({ S25957[657] }),
  .B2({ S5458 }),
  .ZN({ S6993 })
);
NAND2_X1 #() 
NAND2_X1_225_ (
  .A1({ S6993 }),
  .A2({ S110 }),
  .ZN({ S6994 })
);
OAI211_X1 #() 
OAI211_X1_47_ (
  .A({ S6994 }),
  .B({ S25957[660] }),
  .C1({ S6992 }),
  .C2({ S6991 }),
  .ZN({ S6995 })
);
NAND2_X1 #() 
NAND2_X1_226_ (
  .A1({ S6979 }),
  .A2({ S6931 }),
  .ZN({ S6996 })
);
NAND3_X1 #() 
NAND3_X1_250_ (
  .A1({ S25957[658] }),
  .A2({ S2746 }),
  .A3({ S2752 }),
  .ZN({ S6997 })
);
NAND3_X1 #() 
NAND3_X1_251_ (
  .A1({ S6969 }),
  .A2({ S110 }),
  .A3({ S6997 }),
  .ZN({ S6998 })
);
OAI211_X1 #() 
OAI211_X1_48_ (
  .A({ S6930 }),
  .B({ S6998 }),
  .C1({ S6970 }),
  .C2({ S6996 }),
  .ZN({ S6999 })
);
NAND3_X1 #() 
NAND3_X1_252_ (
  .A1({ S6995 }),
  .A2({ S25957[662] }),
  .A3({ S6999 }),
  .ZN({ S7000 })
);
NAND2_X1 #() 
NAND2_X1_227_ (
  .A1({ S6990 }),
  .A2({ S7000 }),
  .ZN({ S7001 })
);
NAND2_X1 #() 
NAND2_X1_228_ (
  .A1({ S7001 }),
  .A2({ S25957[661] }),
  .ZN({ S7002 })
);
AOI21_X1 #() 
AOI21_X1_110_ (
  .A({ S110 }),
  .B1({ S6910 }),
  .B2({ S25957[657] }),
  .ZN({ S7003 })
);
INV_X1 #() 
INV_X1_104_ (
  .A({ S6937 }),
  .ZN({ S7004 })
);
NAND2_X1 #() 
NAND2_X1_229_ (
  .A1({ S6913 }),
  .A2({ S110 }),
  .ZN({ S7005 })
);
OAI21_X1 #() 
OAI21_X1_141_ (
  .A({ S25957[660] }),
  .B1({ S7004 }),
  .B2({ S7005 }),
  .ZN({ S7006 })
);
OR2_X1 #() 
OR2_X1_4_ (
  .A1({ S7006 }),
  .A2({ S7003 }),
  .ZN({ S7007 })
);
NAND2_X1 #() 
NAND2_X1_230_ (
  .A1({ S6907 }),
  .A2({ S14 }),
  .ZN({ S7008 })
);
NAND3_X1 #() 
NAND3_X1_253_ (
  .A1({ S7008 }),
  .A2({ S110 }),
  .A3({ S25957[658] }),
  .ZN({ S7009 })
);
NAND2_X1 #() 
NAND2_X1_231_ (
  .A1({ S6969 }),
  .A2({ S6997 }),
  .ZN({ S7010 })
);
AOI21_X1 #() 
AOI21_X1_111_ (
  .A({ S25957[660] }),
  .B1({ S7010 }),
  .B2({ S25957[659] }),
  .ZN({ S7011 })
);
AOI21_X1 #() 
AOI21_X1_112_ (
  .A({ S25957[662] }),
  .B1({ S7009 }),
  .B2({ S7011 }),
  .ZN({ S7012 })
);
NAND2_X1 #() 
NAND2_X1_232_ (
  .A1({ S6921 }),
  .A2({ S6979 }),
  .ZN({ S7013 })
);
NAND4_X1 #() 
NAND4_X1_20_ (
  .A1({ S6969 }),
  .A2({ S6979 }),
  .A3({ S6931 }),
  .A4({ S6997 }),
  .ZN({ S7014 })
);
AOI21_X1 #() 
AOI21_X1_113_ (
  .A({ S25957[660] }),
  .B1({ S7014 }),
  .B2({ S110 }),
  .ZN({ S7015 })
);
OAI21_X1 #() 
OAI21_X1_142_ (
  .A({ S7015 }),
  .B1({ S110 }),
  .B2({ S7013 }),
  .ZN({ S7016 })
);
AOI22_X1 #() 
AOI22_X1_12_ (
  .A1({ S6916 }),
  .A2({ S6939 }),
  .B1({ S5359 }),
  .B2({ S25957[656] }),
  .ZN({ S7017 })
);
OAI21_X1 #() 
OAI21_X1_143_ (
  .A({ S25957[659] }),
  .B1({ S7017 }),
  .B2({ S7010 }),
  .ZN({ S7018 })
);
NAND3_X1 #() 
NAND3_X1_254_ (
  .A1({ S6937 }),
  .A2({ S110 }),
  .A3({ S6916 }),
  .ZN({ S7019 })
);
NAND3_X1 #() 
NAND3_X1_255_ (
  .A1({ S7018 }),
  .A2({ S25957[660] }),
  .A3({ S7019 }),
  .ZN({ S7021 })
);
AOI21_X1 #() 
AOI21_X1_114_ (
  .A({ S2444 }),
  .B1({ S7021 }),
  .B2({ S7016 }),
  .ZN({ S7022 })
);
AOI21_X1 #() 
AOI21_X1_115_ (
  .A({ S7022 }),
  .B1({ S7012 }),
  .B2({ S7007 }),
  .ZN({ S7023 })
);
OAI211_X1 #() 
OAI211_X1_49_ (
  .A({ S4797 }),
  .B({ S7002 }),
  .C1({ S7023 }),
  .C2({ S25957[661] }),
  .ZN({ S7024 })
);
OAI21_X1 #() 
OAI21_X1_144_ (
  .A({ S7024 }),
  .B1({ S6950 }),
  .B2({ S6977 }),
  .ZN({ S7025 })
);
XNOR2_X1 #() 
XNOR2_X1_9_ (
  .A({ S7025 }),
  .B({ S22150 }),
  .ZN({ S7026 })
);
INV_X1 #() 
INV_X1_105_ (
  .A({ S7026 }),
  .ZN({ S25957[543] })
);
NAND2_X1 #() 
NAND2_X1_233_ (
  .A1({ S6921 }),
  .A2({ S6943 }),
  .ZN({ S7027 })
);
INV_X1 #() 
INV_X1_106_ (
  .A({ S7027 }),
  .ZN({ S7028 })
);
AOI21_X1 #() 
AOI21_X1_116_ (
  .A({ S25957[658] }),
  .B1({ S2752 }),
  .B2({ S2746 }),
  .ZN({ S7029 })
);
NOR2_X1 #() 
NOR2_X1_45_ (
  .A1({ S7029 }),
  .A2({ S25957[657] }),
  .ZN({ S7031 })
);
NAND2_X1 #() 
NAND2_X1_234_ (
  .A1({ S6964 }),
  .A2({ S7031 }),
  .ZN({ S7032 })
);
OAI21_X1 #() 
OAI21_X1_145_ (
  .A({ S7032 }),
  .B1({ S7028 }),
  .B2({ S25957[659] }),
  .ZN({ S7033 })
);
OAI21_X1 #() 
OAI21_X1_146_ (
  .A({ S6930 }),
  .B1({ S6971 }),
  .B2({ S6924 }),
  .ZN({ S7034 })
);
OAI211_X1 #() 
OAI211_X1_50_ (
  .A({ S7034 }),
  .B({ S25957[661] }),
  .C1({ S6930 }),
  .C2({ S7033 }),
  .ZN({ S7035 })
);
NAND3_X1 #() 
NAND3_X1_256_ (
  .A1({ S6916 }),
  .A2({ S6943 }),
  .A3({ S6997 }),
  .ZN({ S7036 })
);
NAND2_X1 #() 
NAND2_X1_235_ (
  .A1({ S7036 }),
  .A2({ S25957[659] }),
  .ZN({ S7037 })
);
NAND2_X1 #() 
NAND2_X1_236_ (
  .A1({ S6941 }),
  .A2({ S6911 }),
  .ZN({ S7038 })
);
AND2_X1 #() 
AND2_X1_11_ (
  .A1({ S7038 }),
  .A2({ S7037 }),
  .ZN({ S7039 })
);
NAND2_X1 #() 
NAND2_X1_237_ (
  .A1({ S6931 }),
  .A2({ S25957[657] }),
  .ZN({ S7040 })
);
NAND2_X1 #() 
NAND2_X1_238_ (
  .A1({ S7040 }),
  .A2({ S25957[659] }),
  .ZN({ S7042 })
);
NAND4_X1 #() 
NAND4_X1_21_ (
  .A1({ S6979 }),
  .A2({ S6969 }),
  .A3({ S110 }),
  .A4({ S25957[656] }),
  .ZN({ S7043 })
);
OAI211_X1 #() 
OAI211_X1_51_ (
  .A({ S6930 }),
  .B({ S7043 }),
  .C1({ S7042 }),
  .C2({ S6984 }),
  .ZN({ S7044 })
);
OAI21_X1 #() 
OAI21_X1_147_ (
  .A({ S7044 }),
  .B1({ S7039 }),
  .B2({ S6930 }),
  .ZN({ S7045 })
);
OAI21_X1 #() 
OAI21_X1_148_ (
  .A({ S7035 }),
  .B1({ S7045 }),
  .B2({ S25957[661] }),
  .ZN({ S7046 })
);
NAND2_X1 #() 
NAND2_X1_239_ (
  .A1({ S6959 }),
  .A2({ S6916 }),
  .ZN({ S7047 })
);
NAND2_X1 #() 
NAND2_X1_240_ (
  .A1({ S7047 }),
  .A2({ S25957[659] }),
  .ZN({ S7048 })
);
AOI21_X1 #() 
AOI21_X1_117_ (
  .A({ S25957[660] }),
  .B1({ S7038 }),
  .B2({ S7048 }),
  .ZN({ S7049 })
);
AOI21_X1 #() 
AOI21_X1_118_ (
  .A({ S6926 }),
  .B1({ S6996 }),
  .B2({ S110 }),
  .ZN({ S7050 })
);
NOR3_X1 #() 
NOR3_X1_7_ (
  .A1({ S7049 }),
  .A2({ S7050 }),
  .A3({ S25957[661] }),
  .ZN({ S7051 })
);
NAND2_X1 #() 
NAND2_X1_241_ (
  .A1({ S6944 }),
  .A2({ S25957[659] }),
  .ZN({ S7053 })
);
NAND3_X1 #() 
NAND3_X1_257_ (
  .A1({ S5282 }),
  .A2({ S25957[657] }),
  .A3({ S5458 }),
  .ZN({ S7054 })
);
OAI21_X1 #() 
OAI21_X1_149_ (
  .A({ S7053 }),
  .B1({ S25957[659] }),
  .B2({ S7054 }),
  .ZN({ S7055 })
);
INV_X1 #() 
INV_X1_107_ (
  .A({ S7055 }),
  .ZN({ S7056 })
);
AOI21_X1 #() 
AOI21_X1_119_ (
  .A({ S6930 }),
  .B1({ S7056 }),
  .B2({ S7009 }),
  .ZN({ S7057 })
);
NAND2_X1 #() 
NAND2_X1_242_ (
  .A1({ S6940 }),
  .A2({ S25957[659] }),
  .ZN({ S7058 })
);
NAND2_X1 #() 
NAND2_X1_243_ (
  .A1({ S7058 }),
  .A2({ S6930 }),
  .ZN({ S7059 })
);
NAND2_X1 #() 
NAND2_X1_244_ (
  .A1({ S6937 }),
  .A2({ S6952 }),
  .ZN({ S7060 })
);
OAI21_X1 #() 
OAI21_X1_150_ (
  .A({ S7053 }),
  .B1({ S7060 }),
  .B2({ S25957[659] }),
  .ZN({ S7061 })
);
OAI21_X1 #() 
OAI21_X1_151_ (
  .A({ S25957[661] }),
  .B1({ S7061 }),
  .B2({ S7059 }),
  .ZN({ S7062 })
);
OAI21_X1 #() 
OAI21_X1_152_ (
  .A({ S2444 }),
  .B1({ S7062 }),
  .B2({ S7057 }),
  .ZN({ S7064 })
);
OAI22_X1 #() 
OAI22_X1_8_ (
  .A1({ S7046 }),
  .A2({ S2444 }),
  .B1({ S7064 }),
  .B2({ S7051 }),
  .ZN({ S7065 })
);
NAND2_X1 #() 
NAND2_X1_245_ (
  .A1({ S6939 }),
  .A2({ S5282 }),
  .ZN({ S7066 })
);
INV_X1 #() 
INV_X1_108_ (
  .A({ S6979 }),
  .ZN({ S7067 })
);
AOI21_X1 #() 
AOI21_X1_120_ (
  .A({ S6930 }),
  .B1({ S7067 }),
  .B2({ S25957[659] }),
  .ZN({ S7068 })
);
OAI21_X1 #() 
OAI21_X1_153_ (
  .A({ S7068 }),
  .B1({ S25957[659] }),
  .B2({ S7066 }),
  .ZN({ S7069 })
);
NAND2_X1 #() 
NAND2_X1_246_ (
  .A1({ S6921 }),
  .A2({ S6972 }),
  .ZN({ S7070 })
);
INV_X1 #() 
INV_X1_109_ (
  .A({ S7070 }),
  .ZN({ S7071 })
);
NOR2_X1 #() 
NOR2_X1_46_ (
  .A1({ S7071 }),
  .A2({ S110 }),
  .ZN({ S7072 })
);
NAND2_X1 #() 
NAND2_X1_247_ (
  .A1({ S6907 }),
  .A2({ S25957[658] }),
  .ZN({ S7073 })
);
NAND3_X1 #() 
NAND3_X1_258_ (
  .A1({ S7073 }),
  .A2({ S110 }),
  .A3({ S6916 }),
  .ZN({ S7075 })
);
INV_X1 #() 
INV_X1_110_ (
  .A({ S7075 }),
  .ZN({ S7076 })
);
OAI21_X1 #() 
OAI21_X1_154_ (
  .A({ S25957[660] }),
  .B1({ S7076 }),
  .B2({ S7072 }),
  .ZN({ S7077 })
);
NOR2_X1 #() 
NOR2_X1_47_ (
  .A1({ S6922 }),
  .A2({ S7029 }),
  .ZN({ S7078 })
);
NOR2_X1 #() 
NOR2_X1_48_ (
  .A1({ S7072 }),
  .A2({ S7078 }),
  .ZN({ S7079 })
);
AOI21_X1 #() 
AOI21_X1_121_ (
  .A({ S4995 }),
  .B1({ S7079 }),
  .B2({ S6930 }),
  .ZN({ S7080 })
);
INV_X1 #() 
INV_X1_111_ (
  .A({ S7037 }),
  .ZN({ S7081 })
);
AOI21_X1 #() 
AOI21_X1_122_ (
  .A({ S7081 }),
  .B1({ S6937 }),
  .B2({ S110 }),
  .ZN({ S7082 })
);
AOI21_X1 #() 
AOI21_X1_123_ (
  .A({ S25957[661] }),
  .B1({ S7082 }),
  .B2({ S6930 }),
  .ZN({ S7083 })
);
AOI22_X1 #() 
AOI22_X1_13_ (
  .A1({ S7083 }),
  .A2({ S7069 }),
  .B1({ S7080 }),
  .B2({ S7077 }),
  .ZN({ S7084 })
);
NAND2_X1 #() 
NAND2_X1_248_ (
  .A1({ S6938 }),
  .A2({ S6931 }),
  .ZN({ S7086 })
);
OAI21_X1 #() 
OAI21_X1_155_ (
  .A({ S25957[659] }),
  .B1({ S7086 }),
  .B2({ S6973 }),
  .ZN({ S7087 })
);
NAND3_X1 #() 
NAND3_X1_259_ (
  .A1({ S7087 }),
  .A2({ S25957[660] }),
  .A3({ S6946 }),
  .ZN({ S7088 })
);
NAND3_X1 #() 
NAND3_X1_260_ (
  .A1({ S6969 }),
  .A2({ S6979 }),
  .A3({ S6931 }),
  .ZN({ S7089 })
);
NAND2_X1 #() 
NAND2_X1_249_ (
  .A1({ S7089 }),
  .A2({ S110 }),
  .ZN({ S7090 })
);
OAI21_X1 #() 
OAI21_X1_156_ (
  .A({ S7090 }),
  .B1({ S7067 }),
  .B2({ S6970 }),
  .ZN({ S7091 })
);
OAI21_X1 #() 
OAI21_X1_157_ (
  .A({ S7088 }),
  .B1({ S7091 }),
  .B2({ S25957[660] }),
  .ZN({ S7092 })
);
NAND2_X1 #() 
NAND2_X1_250_ (
  .A1({ S7092 }),
  .A2({ S25957[661] }),
  .ZN({ S7093 })
);
NAND2_X1 #() 
NAND2_X1_251_ (
  .A1({ S7089 }),
  .A2({ S25957[659] }),
  .ZN({ S7094 })
);
OAI211_X1 #() 
OAI211_X1_52_ (
  .A({ S6916 }),
  .B({ S6939 }),
  .C1({ S5359 }),
  .C2({ S6997 }),
  .ZN({ S7095 })
);
NAND2_X1 #() 
NAND2_X1_252_ (
  .A1({ S7095 }),
  .A2({ S25957[659] }),
  .ZN({ S7097 })
);
AOI21_X1 #() 
AOI21_X1_124_ (
  .A({ S6930 }),
  .B1({ S6963 }),
  .B2({ S110 }),
  .ZN({ S7098 })
);
AOI22_X1 #() 
AOI22_X1_14_ (
  .A1({ S7097 }),
  .A2({ S6930 }),
  .B1({ S7098 }),
  .B2({ S7094 }),
  .ZN({ S7099 })
);
OAI211_X1 #() 
OAI211_X1_53_ (
  .A({ S7093 }),
  .B({ S2444 }),
  .C1({ S25957[661] }),
  .C2({ S7099 }),
  .ZN({ S7100 })
);
OAI211_X1 #() 
OAI211_X1_54_ (
  .A({ S7100 }),
  .B({ S4797 }),
  .C1({ S7084 }),
  .C2({ S2444 }),
  .ZN({ S7101 })
);
OAI21_X1 #() 
OAI21_X1_158_ (
  .A({ S7101 }),
  .B1({ S4797 }),
  .B2({ S7065 }),
  .ZN({ S7102 })
);
NAND2_X1 #() 
NAND2_X1_253_ (
  .A1({ S7102 }),
  .A2({ S22219 }),
  .ZN({ S7103 })
);
INV_X1 #() 
INV_X1_112_ (
  .A({ S7103 }),
  .ZN({ S7104 })
);
NOR2_X1 #() 
NOR2_X1_49_ (
  .A1({ S7102 }),
  .A2({ S22219 }),
  .ZN({ S7105 })
);
NOR2_X1 #() 
NOR2_X1_50_ (
  .A1({ S7104 }),
  .A2({ S7105 }),
  .ZN({ S7106 })
);
INV_X1 #() 
INV_X1_113_ (
  .A({ S7106 }),
  .ZN({ S25957[542] })
);
NAND2_X1 #() 
NAND2_X1_254_ (
  .A1({ S24971 }),
  .A2({ S24969 }),
  .ZN({ S25957[957] })
);
XNOR2_X1 #() 
XNOR2_X1_10_ (
  .A({ S4355 }),
  .B({ S25957[957] }),
  .ZN({ S25957[829] })
);
NAND2_X1 #() 
NAND2_X1_255_ (
  .A1({ S4429 }),
  .A2({ S4432 }),
  .ZN({ S25957[733] })
);
XOR2_X1 #() 
XOR2_X1_4_ (
  .A({ S25957[733] }),
  .B({ S25957[829] }),
  .Z({ S25957[701] })
);
INV_X1 #() 
INV_X1_114_ (
  .A({ S25957[701] }),
  .ZN({ S7108 })
);
NOR2_X1 #() 
NOR2_X1_51_ (
  .A1({ S6931 }),
  .A2({ S5359 }),
  .ZN({ S7109 })
);
OAI211_X1 #() 
OAI211_X1_55_ (
  .A({ S6933 }),
  .B({ S25957[660] }),
  .C1({ S110 }),
  .C2({ S5458 }),
  .ZN({ S7110 })
);
AOI21_X1 #() 
AOI21_X1_125_ (
  .A({ S7110 }),
  .B1({ S7109 }),
  .B2({ S110 }),
  .ZN({ S7111 })
);
NOR2_X1 #() 
NOR2_X1_52_ (
  .A1({ S110 }),
  .A2({ S5458 }),
  .ZN({ S7112 })
);
OAI21_X1 #() 
OAI21_X1_159_ (
  .A({ S6997 }),
  .B1({ S7078 }),
  .B2({ S7112 }),
  .ZN({ S7114 })
);
NOR2_X1 #() 
NOR2_X1_53_ (
  .A1({ S7114 }),
  .A2({ S25957[660] }),
  .ZN({ S7115 })
);
NOR3_X1 #() 
NOR3_X1_8_ (
  .A1({ S7115 }),
  .A2({ S7111 }),
  .A3({ S4995 }),
  .ZN({ S7116 })
);
INV_X1 #() 
INV_X1_115_ (
  .A({ S7116 }),
  .ZN({ S7117 })
);
INV_X1 #() 
INV_X1_116_ (
  .A({ S6996 }),
  .ZN({ S7118 })
);
AOI21_X1 #() 
AOI21_X1_126_ (
  .A({ S110 }),
  .B1({ S6937 }),
  .B2({ S7118 }),
  .ZN({ S7119 })
);
NOR2_X1 #() 
NOR2_X1_54_ (
  .A1({ S6973 }),
  .A2({ S25957[659] }),
  .ZN({ S7120 })
);
NAND2_X1 #() 
NAND2_X1_256_ (
  .A1({ S6907 }),
  .A2({ S6997 }),
  .ZN({ S7121 })
);
NAND2_X1 #() 
NAND2_X1_257_ (
  .A1({ S7120 }),
  .A2({ S7121 }),
  .ZN({ S7122 })
);
INV_X1 #() 
INV_X1_117_ (
  .A({ S7122 }),
  .ZN({ S7123 })
);
NOR3_X1 #() 
NOR3_X1_9_ (
  .A1({ S7123 }),
  .A2({ S7119 }),
  .A3({ S6930 }),
  .ZN({ S7125 })
);
NAND3_X1 #() 
NAND3_X1_261_ (
  .A1({ S25957[657] }),
  .A2({ S25957[656] }),
  .A3({ S25957[658] }),
  .ZN({ S7126 })
);
OAI21_X1 #() 
OAI21_X1_160_ (
  .A({ S6955 }),
  .B1({ S25957[659] }),
  .B2({ S7126 }),
  .ZN({ S7127 })
);
NAND2_X1 #() 
NAND2_X1_258_ (
  .A1({ S7127 }),
  .A2({ S6930 }),
  .ZN({ S7128 })
);
NAND2_X1 #() 
NAND2_X1_259_ (
  .A1({ S7128 }),
  .A2({ S4995 }),
  .ZN({ S7129 })
);
NOR2_X1 #() 
NOR2_X1_55_ (
  .A1({ S7125 }),
  .A2({ S7129 }),
  .ZN({ S7130 })
);
INV_X1 #() 
INV_X1_118_ (
  .A({ S7130 }),
  .ZN({ S7131 })
);
NAND3_X1 #() 
NAND3_X1_262_ (
  .A1({ S7131 }),
  .A2({ S7117 }),
  .A3({ S2444 }),
  .ZN({ S7132 })
);
NAND3_X1 #() 
NAND3_X1_263_ (
  .A1({ S7073 }),
  .A2({ S25957[659] }),
  .A3({ S6916 }),
  .ZN({ S7133 })
);
INV_X1 #() 
INV_X1_119_ (
  .A({ S7133 }),
  .ZN({ S7134 })
);
NAND2_X1 #() 
NAND2_X1_260_ (
  .A1({ S6972 }),
  .A2({ S5458 }),
  .ZN({ S7136 })
);
AOI21_X1 #() 
AOI21_X1_127_ (
  .A({ S25957[659] }),
  .B1({ S7136 }),
  .B2({ S6997 }),
  .ZN({ S7137 })
);
OAI21_X1 #() 
OAI21_X1_161_ (
  .A({ S6930 }),
  .B1({ S7134 }),
  .B2({ S7137 }),
  .ZN({ S7138 })
);
NAND2_X1 #() 
NAND2_X1_261_ (
  .A1({ S6939 }),
  .A2({ S6931 }),
  .ZN({ S7139 })
);
AOI211_X1 #() 
AOI211_X1_2_ (
  .A({ S25957[659] }),
  .B({ S7139 }),
  .C1({ S25957[657] }),
  .C2({ S6984 }),
  .ZN({ S7140 })
);
NAND2_X1 #() 
NAND2_X1_262_ (
  .A1({ S6996 }),
  .A2({ S25957[659] }),
  .ZN({ S7141 })
);
NAND2_X1 #() 
NAND2_X1_263_ (
  .A1({ S7141 }),
  .A2({ S25957[660] }),
  .ZN({ S7142 })
);
OAI211_X1 #() 
OAI211_X1_56_ (
  .A({ S7138 }),
  .B({ S4995 }),
  .C1({ S7140 }),
  .C2({ S7142 }),
  .ZN({ S7143 })
);
NAND3_X1 #() 
NAND3_X1_264_ (
  .A1({ S6938 }),
  .A2({ S25957[658] }),
  .A3({ S6972 }),
  .ZN({ S7144 })
);
NAND3_X1 #() 
NAND3_X1_265_ (
  .A1({ S7144 }),
  .A2({ S25957[659] }),
  .A3({ S7054 }),
  .ZN({ S7145 })
);
OAI211_X1 #() 
OAI211_X1_57_ (
  .A({ S7145 }),
  .B({ S25957[660] }),
  .C1({ S25957[659] }),
  .C2({ S7089 }),
  .ZN({ S7147 })
);
NOR2_X1 #() 
NOR2_X1_56_ (
  .A1({ S6946 }),
  .A2({ S6973 }),
  .ZN({ S7148 })
);
AOI21_X1 #() 
AOI21_X1_128_ (
  .A({ S7148 }),
  .B1({ S5282 }),
  .B2({ S25957[659] }),
  .ZN({ S7149 })
);
OAI211_X1 #() 
OAI211_X1_58_ (
  .A({ S7147 }),
  .B({ S25957[661] }),
  .C1({ S25957[660] }),
  .C2({ S7149 }),
  .ZN({ S7150 })
);
NAND3_X1 #() 
NAND3_X1_266_ (
  .A1({ S7143 }),
  .A2({ S25957[662] }),
  .A3({ S7150 }),
  .ZN({ S7151 })
);
NAND3_X1 #() 
NAND3_X1_267_ (
  .A1({ S7132 }),
  .A2({ S4797 }),
  .A3({ S7151 }),
  .ZN({ S7152 })
);
OAI21_X1 #() 
OAI21_X1_162_ (
  .A({ S110 }),
  .B1({ S6997 }),
  .B2({ S5359 }),
  .ZN({ S7153 })
);
OAI22_X1 #() 
OAI22_X1_9_ (
  .A1({ S7153 }),
  .A2({ S6996 }),
  .B1({ S7066 }),
  .B2({ S110 }),
  .ZN({ S7154 })
);
NAND2_X1 #() 
NAND2_X1_264_ (
  .A1({ S7154 }),
  .A2({ S25957[660] }),
  .ZN({ S7155 })
);
NOR2_X1 #() 
NOR2_X1_57_ (
  .A1({ S25957[660] }),
  .A2({ S6984 }),
  .ZN({ S7156 })
);
NAND3_X1 #() 
NAND3_X1_268_ (
  .A1({ S7156 }),
  .A2({ S6922 }),
  .A3({ S7042 }),
  .ZN({ S7158 })
);
NAND3_X1 #() 
NAND3_X1_269_ (
  .A1({ S7155 }),
  .A2({ S25957[661] }),
  .A3({ S7158 }),
  .ZN({ S7159 })
);
AOI21_X1 #() 
AOI21_X1_129_ (
  .A({ S25957[660] }),
  .B1({ S7009 }),
  .B2({ S7037 }),
  .ZN({ S7160 })
);
NAND2_X1 #() 
NAND2_X1_265_ (
  .A1({ S6972 }),
  .A2({ S25957[658] }),
  .ZN({ S7161 })
);
AOI21_X1 #() 
AOI21_X1_130_ (
  .A({ S6930 }),
  .B1({ S7161 }),
  .B2({ S110 }),
  .ZN({ S7162 })
);
AND2_X1 #() 
AND2_X1_12_ (
  .A1({ S7162 }),
  .A2({ S7058 }),
  .ZN({ S7163 })
);
OAI21_X1 #() 
OAI21_X1_163_ (
  .A({ S4995 }),
  .B1({ S7163 }),
  .B2({ S7160 }),
  .ZN({ S7164 })
);
AND2_X1 #() 
AND2_X1_13_ (
  .A1({ S7164 }),
  .A2({ S7159 }),
  .ZN({ S7165 })
);
NAND2_X1 #() 
NAND2_X1_266_ (
  .A1({ S6938 }),
  .A2({ S6997 }),
  .ZN({ S7166 })
);
NAND2_X1 #() 
NAND2_X1_267_ (
  .A1({ S7166 }),
  .A2({ S110 }),
  .ZN({ S7167 })
);
OAI21_X1 #() 
OAI21_X1_164_ (
  .A({ S7167 }),
  .B1({ S110 }),
  .B2({ S7014 }),
  .ZN({ S7169 })
);
NAND2_X1 #() 
NAND2_X1_268_ (
  .A1({ S7169 }),
  .A2({ S25957[660] }),
  .ZN({ S7170 })
);
NAND3_X1 #() 
NAND3_X1_270_ (
  .A1({ S6972 }),
  .A2({ S6939 }),
  .A3({ S110 }),
  .ZN({ S7171 })
);
AND2_X1 #() 
AND2_X1_14_ (
  .A1({ S7171 }),
  .A2({ S6925 }),
  .ZN({ S7172 })
);
OAI211_X1 #() 
OAI211_X1_59_ (
  .A({ S7170 }),
  .B({ S25957[661] }),
  .C1({ S25957[660] }),
  .C2({ S7172 }),
  .ZN({ S7173 })
);
NAND3_X1 #() 
NAND3_X1_271_ (
  .A1({ S7144 }),
  .A2({ S25957[659] }),
  .A3({ S6952 }),
  .ZN({ S7174 })
);
AOI21_X1 #() 
AOI21_X1_131_ (
  .A({ S25957[660] }),
  .B1({ S7174 }),
  .B2({ S7005 }),
  .ZN({ S7175 })
);
NAND2_X1 #() 
NAND2_X1_269_ (
  .A1({ S7139 }),
  .A2({ S14 }),
  .ZN({ S7176 })
);
NOR2_X1 #() 
NOR2_X1_58_ (
  .A1({ S7176 }),
  .A2({ S110 }),
  .ZN({ S7177 })
);
AOI21_X1 #() 
AOI21_X1_132_ (
  .A({ S6930 }),
  .B1({ S7031 }),
  .B2({ S110 }),
  .ZN({ S7178 })
);
INV_X1 #() 
INV_X1_120_ (
  .A({ S7178 }),
  .ZN({ S7180 })
);
OAI21_X1 #() 
OAI21_X1_165_ (
  .A({ S4995 }),
  .B1({ S7180 }),
  .B2({ S7177 }),
  .ZN({ S7181 })
);
OAI211_X1 #() 
OAI211_X1_60_ (
  .A({ S7173 }),
  .B({ S2444 }),
  .C1({ S7175 }),
  .C2({ S7181 }),
  .ZN({ S7182 })
);
OAI211_X1 #() 
OAI211_X1_61_ (
  .A({ S7182 }),
  .B({ S25957[663] }),
  .C1({ S2444 }),
  .C2({ S7165 }),
  .ZN({ S7183 })
);
AOI21_X1 #() 
AOI21_X1_133_ (
  .A({ S4355 }),
  .B1({ S7152 }),
  .B2({ S7183 }),
  .ZN({ S7184 })
);
NAND3_X1 #() 
NAND3_X1_272_ (
  .A1({ S7171 }),
  .A2({ S6930 }),
  .A3({ S6925 }),
  .ZN({ S7185 })
);
OAI211_X1 #() 
OAI211_X1_62_ (
  .A({ S25957[661] }),
  .B({ S7185 }),
  .C1({ S7169 }),
  .C2({ S6930 }),
  .ZN({ S7186 })
);
NOR2_X1 #() 
NOR2_X1_59_ (
  .A1({ S7180 }),
  .A2({ S7177 }),
  .ZN({ S7187 })
);
NOR2_X1 #() 
NOR2_X1_60_ (
  .A1({ S7175 }),
  .A2({ S7187 }),
  .ZN({ S7188 })
);
OAI211_X1 #() 
OAI211_X1_63_ (
  .A({ S7186 }),
  .B({ S2444 }),
  .C1({ S25957[661] }),
  .C2({ S7188 }),
  .ZN({ S7189 })
);
NAND3_X1 #() 
NAND3_X1_273_ (
  .A1({ S7164 }),
  .A2({ S25957[662] }),
  .A3({ S7159 }),
  .ZN({ S7191 })
);
NAND3_X1 #() 
NAND3_X1_274_ (
  .A1({ S7189 }),
  .A2({ S25957[663] }),
  .A3({ S7191 }),
  .ZN({ S7192 })
);
OAI21_X1 #() 
OAI21_X1_166_ (
  .A({ S2444 }),
  .B1({ S7130 }),
  .B2({ S7116 }),
  .ZN({ S7193 })
);
AND2_X1 #() 
AND2_X1_15_ (
  .A1({ S7143 }),
  .A2({ S7150 }),
  .ZN({ S7194 })
);
OAI211_X1 #() 
OAI211_X1_64_ (
  .A({ S7193 }),
  .B({ S4797 }),
  .C1({ S7194 }),
  .C2({ S2444 }),
  .ZN({ S7195 })
);
AOI21_X1 #() 
AOI21_X1_134_ (
  .A({ S25957[861] }),
  .B1({ S7195 }),
  .B2({ S7192 }),
  .ZN({ S7196 })
);
OAI21_X1 #() 
OAI21_X1_167_ (
  .A({ S7108 }),
  .B1({ S7184 }),
  .B2({ S7196 }),
  .ZN({ S7197 })
);
NAND3_X1 #() 
NAND3_X1_275_ (
  .A1({ S7195 }),
  .A2({ S7192 }),
  .A3({ S25957[861] }),
  .ZN({ S7198 })
);
NAND3_X1 #() 
NAND3_X1_276_ (
  .A1({ S7152 }),
  .A2({ S4355 }),
  .A3({ S7183 }),
  .ZN({ S7199 })
);
NAND3_X1 #() 
NAND3_X1_277_ (
  .A1({ S7199 }),
  .A2({ S7198 }),
  .A3({ S25957[701] }),
  .ZN({ S7200 })
);
NAND3_X1 #() 
NAND3_X1_278_ (
  .A1({ S7197 }),
  .A2({ S25957[669] }),
  .A3({ S7200 }),
  .ZN({ S7202 })
);
OAI21_X1 #() 
OAI21_X1_168_ (
  .A({ S25957[701] }),
  .B1({ S7184 }),
  .B2({ S7196 }),
  .ZN({ S7203 })
);
NAND3_X1 #() 
NAND3_X1_279_ (
  .A1({ S7199 }),
  .A2({ S7198 }),
  .A3({ S7108 }),
  .ZN({ S7204 })
);
NAND3_X1 #() 
NAND3_X1_280_ (
  .A1({ S7203 }),
  .A2({ S6306 }),
  .A3({ S7204 }),
  .ZN({ S7205 })
);
NAND2_X1 #() 
NAND2_X1_270_ (
  .A1({ S7202 }),
  .A2({ S7205 }),
  .ZN({ S25957[541] })
);
NOR2_X1 #() 
NOR2_X1_61_ (
  .A1({ S6198 }),
  .A2({ S6199 }),
  .ZN({ S7206 })
);
INV_X1 #() 
INV_X1_121_ (
  .A({ S7206 }),
  .ZN({ S25957[700] })
);
NAND3_X1 #() 
NAND3_X1_281_ (
  .A1({ S7054 }),
  .A2({ S25957[659] }),
  .A3({ S6938 }),
  .ZN({ S7207 })
);
NAND2_X1 #() 
NAND2_X1_271_ (
  .A1({ S6943 }),
  .A2({ S6997 }),
  .ZN({ S7208 })
);
OAI21_X1 #() 
OAI21_X1_169_ (
  .A({ S110 }),
  .B1({ S6940 }),
  .B2({ S7208 }),
  .ZN({ S7209 })
);
AND3_X1 #() 
AND3_X1_11_ (
  .A1({ S7209 }),
  .A2({ S7207 }),
  .A3({ S25957[660] }),
  .ZN({ S7211 })
);
AOI21_X1 #() 
AOI21_X1_135_ (
  .A({ S25957[659] }),
  .B1({ S6941 }),
  .B2({ S7073 }),
  .ZN({ S7212 })
);
NOR2_X1 #() 
NOR2_X1_62_ (
  .A1({ S6997 }),
  .A2({ S5359 }),
  .ZN({ S7213 })
);
NAND2_X1 #() 
NAND2_X1_272_ (
  .A1({ S7213 }),
  .A2({ S25957[659] }),
  .ZN({ S7214 })
);
NAND3_X1 #() 
NAND3_X1_282_ (
  .A1({ S7214 }),
  .A2({ S7141 }),
  .A3({ S6930 }),
  .ZN({ S7215 })
);
OAI21_X1 #() 
OAI21_X1_170_ (
  .A({ S25957[661] }),
  .B1({ S7212 }),
  .B2({ S7215 }),
  .ZN({ S7216 })
);
NAND3_X1 #() 
NAND3_X1_283_ (
  .A1({ S25957[659] }),
  .A2({ S6921 }),
  .A3({ S5359 }),
  .ZN({ S7217 })
);
AOI21_X1 #() 
AOI21_X1_136_ (
  .A({ S25957[660] }),
  .B1({ S7095 }),
  .B2({ S110 }),
  .ZN({ S7218 })
);
NAND2_X1 #() 
NAND2_X1_273_ (
  .A1({ S7218 }),
  .A2({ S7217 }),
  .ZN({ S7219 })
);
NAND2_X1 #() 
NAND2_X1_274_ (
  .A1({ S6939 }),
  .A2({ S6997 }),
  .ZN({ S7220 })
);
NAND3_X1 #() 
NAND3_X1_284_ (
  .A1({ S7220 }),
  .A2({ S25957[659] }),
  .A3({ S6969 }),
  .ZN({ S7222 })
);
OAI211_X1 #() 
OAI211_X1_65_ (
  .A({ S7222 }),
  .B({ S25957[660] }),
  .C1({ S6991 }),
  .C2({ S7153 }),
  .ZN({ S7223 })
);
NAND3_X1 #() 
NAND3_X1_285_ (
  .A1({ S7219 }),
  .A2({ S7223 }),
  .A3({ S4995 }),
  .ZN({ S7224 })
);
OAI211_X1 #() 
OAI211_X1_66_ (
  .A({ S7224 }),
  .B({ S2444 }),
  .C1({ S7216 }),
  .C2({ S7211 }),
  .ZN({ S7225 })
);
NAND2_X1 #() 
NAND2_X1_275_ (
  .A1({ S6951 }),
  .A2({ S110 }),
  .ZN({ S7226 })
);
NAND3_X1 #() 
NAND3_X1_286_ (
  .A1({ S7226 }),
  .A2({ S7141 }),
  .A3({ S25957[660] }),
  .ZN({ S7227 })
);
NAND3_X1 #() 
NAND3_X1_287_ (
  .A1({ S6979 }),
  .A2({ S110 }),
  .A3({ S5282 }),
  .ZN({ S7228 })
);
NAND3_X1 #() 
NAND3_X1_288_ (
  .A1({ S6986 }),
  .A2({ S6930 }),
  .A3({ S7228 }),
  .ZN({ S7229 })
);
NAND3_X1 #() 
NAND3_X1_289_ (
  .A1({ S7229 }),
  .A2({ S25957[661] }),
  .A3({ S7227 }),
  .ZN({ S7230 })
);
OAI211_X1 #() 
OAI211_X1_67_ (
  .A({ S7171 }),
  .B({ S25957[660] }),
  .C1({ S6917 }),
  .C2({ S110 }),
  .ZN({ S7231 })
);
NAND2_X1 #() 
NAND2_X1_276_ (
  .A1({ S7013 }),
  .A2({ S110 }),
  .ZN({ S7233 })
);
OAI211_X1 #() 
OAI211_X1_68_ (
  .A({ S7233 }),
  .B({ S6930 }),
  .C1({ S110 }),
  .C2({ S6980 }),
  .ZN({ S7234 })
);
NAND3_X1 #() 
NAND3_X1_290_ (
  .A1({ S7234 }),
  .A2({ S4995 }),
  .A3({ S7231 }),
  .ZN({ S7235 })
);
NAND3_X1 #() 
NAND3_X1_291_ (
  .A1({ S7235 }),
  .A2({ S7230 }),
  .A3({ S25957[662] }),
  .ZN({ S7236 })
);
NAND3_X1 #() 
NAND3_X1_292_ (
  .A1({ S7225 }),
  .A2({ S25957[663] }),
  .A3({ S7236 }),
  .ZN({ S7237 })
);
NAND2_X1 #() 
NAND2_X1_277_ (
  .A1({ S7162 }),
  .A2({ S7094 }),
  .ZN({ S7238 })
);
OAI21_X1 #() 
OAI21_X1_171_ (
  .A({ S6930 }),
  .B1({ S25957[659] }),
  .B2({ S6907 }),
  .ZN({ S7239 })
);
OAI211_X1 #() 
OAI211_X1_69_ (
  .A({ S7238 }),
  .B({ S25957[661] }),
  .C1({ S7177 }),
  .C2({ S7239 }),
  .ZN({ S7240 })
);
NAND2_X1 #() 
NAND2_X1_278_ (
  .A1({ S6985 }),
  .A2({ S14 }),
  .ZN({ S7241 })
);
NAND3_X1 #() 
NAND3_X1_293_ (
  .A1({ S6952 }),
  .A2({ S6951 }),
  .A3({ S110 }),
  .ZN({ S7242 })
);
AOI21_X1 #() 
AOI21_X1_137_ (
  .A({ S25957[660] }),
  .B1({ S7241 }),
  .B2({ S7242 }),
  .ZN({ S7244 })
);
NAND4_X1 #() 
NAND4_X1_22_ (
  .A1({ S25957[659] }),
  .A2({ S6921 }),
  .A3({ S6979 }),
  .A4({ S6931 }),
  .ZN({ S7245 })
);
AND3_X1 #() 
AND3_X1_12_ (
  .A1({ S7245 }),
  .A2({ S7171 }),
  .A3({ S25957[660] }),
  .ZN({ S7246 })
);
OAI21_X1 #() 
OAI21_X1_172_ (
  .A({ S4995 }),
  .B1({ S7244 }),
  .B2({ S7246 }),
  .ZN({ S7247 })
);
NAND3_X1 #() 
NAND3_X1_294_ (
  .A1({ S7247 }),
  .A2({ S7240 }),
  .A3({ S2444 }),
  .ZN({ S7248 })
);
INV_X1 #() 
INV_X1_122_ (
  .A({ S139 }),
  .ZN({ S7249 })
);
OAI21_X1 #() 
OAI21_X1_173_ (
  .A({ S25957[660] }),
  .B1({ S7249 }),
  .B2({ S25957[658] }),
  .ZN({ S7250 })
);
AOI21_X1 #() 
AOI21_X1_138_ (
  .A({ S25957[659] }),
  .B1({ S7176 }),
  .B2({ S7161 }),
  .ZN({ S7251 })
);
NAND2_X1 #() 
NAND2_X1_279_ (
  .A1({ S7133 }),
  .A2({ S6930 }),
  .ZN({ S7252 })
);
OAI211_X1 #() 
OAI211_X1_70_ (
  .A({ S25957[661] }),
  .B({ S7250 }),
  .C1({ S7252 }),
  .C2({ S7251 }),
  .ZN({ S7253 })
);
NOR2_X1 #() 
NOR2_X1_63_ (
  .A1({ S7112 }),
  .A2({ S25957[660] }),
  .ZN({ S7255 })
);
OAI21_X1 #() 
OAI21_X1_174_ (
  .A({ S7255 }),
  .B1({ S6910 }),
  .B2({ S7005 }),
  .ZN({ S7256 })
);
NAND3_X1 #() 
NAND3_X1_295_ (
  .A1({ S6921 }),
  .A2({ S110 }),
  .A3({ S6943 }),
  .ZN({ S7257 })
);
NOR2_X1 #() 
NOR2_X1_64_ (
  .A1({ S7257 }),
  .A2({ S6908 }),
  .ZN({ S7258 })
);
OAI211_X1 #() 
OAI211_X1_71_ (
  .A({ S7256 }),
  .B({ S4995 }),
  .C1({ S6926 }),
  .C2({ S7258 }),
  .ZN({ S7259 })
);
NAND3_X1 #() 
NAND3_X1_296_ (
  .A1({ S7253 }),
  .A2({ S7259 }),
  .A3({ S25957[662] }),
  .ZN({ S7260 })
);
NAND3_X1 #() 
NAND3_X1_297_ (
  .A1({ S7248 }),
  .A2({ S7260 }),
  .A3({ S4797 }),
  .ZN({ S7261 })
);
NAND3_X1 #() 
NAND3_X1_298_ (
  .A1({ S7237 }),
  .A2({ S7261 }),
  .A3({ S4495 }),
  .ZN({ S7262 })
);
NAND2_X1 #() 
NAND2_X1_280_ (
  .A1({ S7237 }),
  .A2({ S7261 }),
  .ZN({ S7263 })
);
NAND2_X1 #() 
NAND2_X1_281_ (
  .A1({ S7263 }),
  .A2({ S25957[860] }),
  .ZN({ S7264 })
);
NAND3_X1 #() 
NAND3_X1_299_ (
  .A1({ S7264 }),
  .A2({ S7206 }),
  .A3({ S7262 }),
  .ZN({ S7266 })
);
AND3_X1 #() 
AND3_X1_13_ (
  .A1({ S7237 }),
  .A2({ S7261 }),
  .A3({ S4495 }),
  .ZN({ S7267 })
);
AOI21_X1 #() 
AOI21_X1_139_ (
  .A({ S4495 }),
  .B1({ S7237 }),
  .B2({ S7261 }),
  .ZN({ S7268 })
);
OAI21_X1 #() 
OAI21_X1_175_ (
  .A({ S25957[700] }),
  .B1({ S7267 }),
  .B2({ S7268 }),
  .ZN({ S7269 })
);
NAND3_X1 #() 
NAND3_X1_300_ (
  .A1({ S7269 }),
  .A2({ S7266 }),
  .A3({ S6201 }),
  .ZN({ S7270 })
);
OAI21_X1 #() 
OAI21_X1_176_ (
  .A({ S7206 }),
  .B1({ S7267 }),
  .B2({ S7268 }),
  .ZN({ S7271 })
);
NAND3_X1 #() 
NAND3_X1_301_ (
  .A1({ S7264 }),
  .A2({ S25957[700] }),
  .A3({ S7262 }),
  .ZN({ S7272 })
);
NAND3_X1 #() 
NAND3_X1_302_ (
  .A1({ S7271 }),
  .A2({ S7272 }),
  .A3({ S25957[668] }),
  .ZN({ S7273 })
);
NAND2_X1 #() 
NAND2_X1_282_ (
  .A1({ S7270 }),
  .A2({ S7273 }),
  .ZN({ S25957[540] })
);
NAND3_X1 #() 
NAND3_X1_303_ (
  .A1({ S6937 }),
  .A2({ S110 }),
  .A3({ S6939 }),
  .ZN({ S7274 })
);
NAND4_X1 #() 
NAND4_X1_23_ (
  .A1({ S25957[659] }),
  .A2({ S25957[657] }),
  .A3({ S6916 }),
  .A4({ S6997 }),
  .ZN({ S7276 })
);
NAND3_X1 #() 
NAND3_X1_304_ (
  .A1({ S7274 }),
  .A2({ S6930 }),
  .A3({ S7276 }),
  .ZN({ S7277 })
);
INV_X1 #() 
INV_X1_123_ (
  .A({ S7176 }),
  .ZN({ S7278 })
);
AOI21_X1 #() 
AOI21_X1_140_ (
  .A({ S6930 }),
  .B1({ S7036 }),
  .B2({ S110 }),
  .ZN({ S7279 })
);
OAI21_X1 #() 
OAI21_X1_177_ (
  .A({ S7279 }),
  .B1({ S6992 }),
  .B2({ S7278 }),
  .ZN({ S7280 })
);
NAND3_X1 #() 
NAND3_X1_305_ (
  .A1({ S7280 }),
  .A2({ S2444 }),
  .A3({ S7277 }),
  .ZN({ S7281 })
);
INV_X1 #() 
INV_X1_124_ (
  .A({ S7166 }),
  .ZN({ S7282 })
);
NOR3_X1 #() 
NOR3_X1_10_ (
  .A1({ S6940 }),
  .A2({ S7208 }),
  .A3({ S110 }),
  .ZN({ S7283 })
);
AOI21_X1 #() 
AOI21_X1_141_ (
  .A({ S7283 }),
  .B1({ S7282 }),
  .B2({ S7120 }),
  .ZN({ S7284 })
);
NAND3_X1 #() 
NAND3_X1_306_ (
  .A1({ S6959 }),
  .A2({ S110 }),
  .A3({ S6938 }),
  .ZN({ S7285 })
);
NAND3_X1 #() 
NAND3_X1_307_ (
  .A1({ S7241 }),
  .A2({ S7285 }),
  .A3({ S25957[660] }),
  .ZN({ S7287 })
);
OAI211_X1 #() 
OAI211_X1_72_ (
  .A({ S25957[662] }),
  .B({ S7287 }),
  .C1({ S7284 }),
  .C2({ S25957[660] }),
  .ZN({ S7288 })
);
AND2_X1 #() 
AND2_X1_16_ (
  .A1({ S7288 }),
  .A2({ S7281 }),
  .ZN({ S7289 })
);
NAND2_X1 #() 
NAND2_X1_283_ (
  .A1({ S6921 }),
  .A2({ S5359 }),
  .ZN({ S7290 })
);
NAND3_X1 #() 
NAND3_X1_308_ (
  .A1({ S7290 }),
  .A2({ S25957[659] }),
  .A3({ S7126 }),
  .ZN({ S7291 })
);
OAI211_X1 #() 
OAI211_X1_73_ (
  .A({ S7291 }),
  .B({ S6930 }),
  .C1({ S25957[659] }),
  .C2({ S7070 }),
  .ZN({ S7292 })
);
NAND2_X1 #() 
NAND2_X1_284_ (
  .A1({ S6941 }),
  .A2({ S25957[659] }),
  .ZN({ S7293 })
);
NAND3_X1 #() 
NAND3_X1_309_ (
  .A1({ S7293 }),
  .A2({ S25957[660] }),
  .A3({ S7233 }),
  .ZN({ S7294 })
);
NAND3_X1 #() 
NAND3_X1_310_ (
  .A1({ S7294 }),
  .A2({ S2444 }),
  .A3({ S7292 }),
  .ZN({ S7295 })
);
INV_X1 #() 
INV_X1_125_ (
  .A({ S7295 }),
  .ZN({ S7296 })
);
NAND2_X1 #() 
NAND2_X1_285_ (
  .A1({ S7029 }),
  .A2({ S5359 }),
  .ZN({ S7298 })
);
NAND3_X1 #() 
NAND3_X1_311_ (
  .A1({ S7144 }),
  .A2({ S110 }),
  .A3({ S7298 }),
  .ZN({ S7299 })
);
AOI21_X1 #() 
AOI21_X1_142_ (
  .A({ S6930 }),
  .B1({ S7299 }),
  .B2({ S7042 }),
  .ZN({ S7300 })
);
INV_X1 #() 
INV_X1_126_ (
  .A({ S7255 }),
  .ZN({ S7301 })
);
OAI21_X1 #() 
OAI21_X1_178_ (
  .A({ S25957[662] }),
  .B1({ S7301 }),
  .B2({ S7071 }),
  .ZN({ S7302 })
);
NOR2_X1 #() 
NOR2_X1_65_ (
  .A1({ S7302 }),
  .A2({ S7300 }),
  .ZN({ S7303 })
);
OAI21_X1 #() 
OAI21_X1_179_ (
  .A({ S4995 }),
  .B1({ S7296 }),
  .B2({ S7303 }),
  .ZN({ S7304 })
);
OAI211_X1 #() 
OAI211_X1_74_ (
  .A({ S25957[663] }),
  .B({ S7304 }),
  .C1({ S7289 }),
  .C2({ S4995 }),
  .ZN({ S7305 })
);
NAND4_X1 #() 
NAND4_X1_24_ (
  .A1({ S6970 }),
  .A2({ S6979 }),
  .A3({ S25957[656] }),
  .A4({ S6930 }),
  .ZN({ S7306 })
);
OAI21_X1 #() 
OAI21_X1_180_ (
  .A({ S25957[660] }),
  .B1({ S110 }),
  .B2({ S5282 }),
  .ZN({ S7307 })
);
OAI21_X1 #() 
OAI21_X1_181_ (
  .A({ S7306 }),
  .B1({ S7144 }),
  .B2({ S7307 }),
  .ZN({ S7309 })
);
OAI211_X1 #() 
OAI211_X1_75_ (
  .A({ S7019 }),
  .B({ S6930 }),
  .C1({ S6991 }),
  .C2({ S6965 }),
  .ZN({ S7310 })
);
NAND4_X1 #() 
NAND4_X1_25_ (
  .A1({ S6938 }),
  .A2({ S25957[659] }),
  .A3({ S6921 }),
  .A4({ S6972 }),
  .ZN({ S7311 })
);
NAND2_X1 #() 
NAND2_X1_286_ (
  .A1({ S7090 }),
  .A2({ S7311 }),
  .ZN({ S7312 })
);
AOI21_X1 #() 
AOI21_X1_143_ (
  .A({ S25957[661] }),
  .B1({ S7312 }),
  .B2({ S25957[660] }),
  .ZN({ S7313 })
);
NAND2_X1 #() 
NAND2_X1_287_ (
  .A1({ S7313 }),
  .A2({ S7310 }),
  .ZN({ S7314 })
);
OAI21_X1 #() 
OAI21_X1_182_ (
  .A({ S7314 }),
  .B1({ S4995 }),
  .B2({ S7309 }),
  .ZN({ S7315 })
);
AOI22_X1 #() 
AOI22_X1_15_ (
  .A1({ S6939 }),
  .A2({ S25957[656] }),
  .B1({ S2665 }),
  .B2({ S2662 }),
  .ZN({ S7316 })
);
OAI211_X1 #() 
OAI211_X1_76_ (
  .A({ S6930 }),
  .B({ S7043 }),
  .C1({ S6965 }),
  .C2({ S6963 }),
  .ZN({ S7317 })
);
OAI211_X1 #() 
OAI211_X1_77_ (
  .A({ S7317 }),
  .B({ S4995 }),
  .C1({ S6930 }),
  .C2({ S7316 }),
  .ZN({ S7318 })
);
NAND3_X1 #() 
NAND3_X1_312_ (
  .A1({ S6938 }),
  .A2({ S110 }),
  .A3({ S6979 }),
  .ZN({ S7320 })
);
NAND3_X1 #() 
NAND3_X1_313_ (
  .A1({ S25957[659] }),
  .A2({ S5282 }),
  .A3({ S6943 }),
  .ZN({ S7321 })
);
NAND3_X1 #() 
NAND3_X1_314_ (
  .A1({ S7320 }),
  .A2({ S7321 }),
  .A3({ S6930 }),
  .ZN({ S7322 })
);
OAI211_X1 #() 
OAI211_X1_78_ (
  .A({ S25957[661] }),
  .B({ S7322 }),
  .C1({ S7006 }),
  .C2({ S7081 }),
  .ZN({ S7323 })
);
NAND3_X1 #() 
NAND3_X1_315_ (
  .A1({ S7323 }),
  .A2({ S25957[662] }),
  .A3({ S7318 }),
  .ZN({ S7324 })
);
OAI211_X1 #() 
OAI211_X1_79_ (
  .A({ S7324 }),
  .B({ S4797 }),
  .C1({ S7315 }),
  .C2({ S25957[662] }),
  .ZN({ S7325 })
);
NAND3_X1 #() 
NAND3_X1_316_ (
  .A1({ S7305 }),
  .A2({ S83 }),
  .A3({ S7325 }),
  .ZN({ S7326 })
);
NAND2_X1 #() 
NAND2_X1_288_ (
  .A1({ S7323 }),
  .A2({ S7318 }),
  .ZN({ S7327 })
);
NAND2_X1 #() 
NAND2_X1_289_ (
  .A1({ S7327 }),
  .A2({ S25957[662] }),
  .ZN({ S7328 })
);
NAND2_X1 #() 
NAND2_X1_290_ (
  .A1({ S7315 }),
  .A2({ S2444 }),
  .ZN({ S7329 })
);
NAND3_X1 #() 
NAND3_X1_317_ (
  .A1({ S7329 }),
  .A2({ S7328 }),
  .A3({ S4797 }),
  .ZN({ S7331 })
);
AOI21_X1 #() 
AOI21_X1_144_ (
  .A({ S4995 }),
  .B1({ S7288 }),
  .B2({ S7281 }),
  .ZN({ S7332 })
);
OR2_X1 #() 
OR2_X1_5_ (
  .A1({ S7302 }),
  .A2({ S7300 }),
  .ZN({ S7333 })
);
AOI21_X1 #() 
AOI21_X1_145_ (
  .A({ S25957[661] }),
  .B1({ S7333 }),
  .B2({ S7295 }),
  .ZN({ S7334 })
);
OAI21_X1 #() 
OAI21_X1_183_ (
  .A({ S25957[663] }),
  .B1({ S7334 }),
  .B2({ S7332 }),
  .ZN({ S7335 })
);
NAND3_X1 #() 
NAND3_X1_318_ (
  .A1({ S7335 }),
  .A2({ S7331 }),
  .A3({ S25957[1051] }),
  .ZN({ S7336 })
);
AND2_X1 #() 
AND2_X1_17_ (
  .A1({ S7326 }),
  .A2({ S7336 }),
  .ZN({ S15 })
);
NAND2_X1 #() 
NAND2_X1_291_ (
  .A1({ S7326 }),
  .A2({ S7336 }),
  .ZN({ S25957[539] })
);
OAI21_X1 #() 
OAI21_X1_184_ (
  .A({ S110 }),
  .B1({ S6963 }),
  .B2({ S7213 }),
  .ZN({ S7337 })
);
NAND3_X1 #() 
NAND3_X1_319_ (
  .A1({ S7337 }),
  .A2({ S25957[660] }),
  .A3({ S6992 }),
  .ZN({ S7338 })
);
NAND4_X1 #() 
NAND4_X1_26_ (
  .A1({ S7226 }),
  .A2({ S7214 }),
  .A3({ S7141 }),
  .A4({ S6930 }),
  .ZN({ S7340 })
);
NAND3_X1 #() 
NAND3_X1_320_ (
  .A1({ S7338 }),
  .A2({ S25957[661] }),
  .A3({ S7340 }),
  .ZN({ S7341 })
);
OAI21_X1 #() 
OAI21_X1_185_ (
  .A({ S7053 }),
  .B1({ S7176 }),
  .B2({ S25957[659] }),
  .ZN({ S7342 })
);
NAND2_X1 #() 
NAND2_X1_292_ (
  .A1({ S7342 }),
  .A2({ S25957[660] }),
  .ZN({ S7343 })
);
NAND2_X1 #() 
NAND2_X1_293_ (
  .A1({ S7047 }),
  .A2({ S110 }),
  .ZN({ S7344 })
);
NAND3_X1 #() 
NAND3_X1_321_ (
  .A1({ S7344 }),
  .A2({ S6930 }),
  .A3({ S7321 }),
  .ZN({ S7345 })
);
NAND3_X1 #() 
NAND3_X1_322_ (
  .A1({ S7343 }),
  .A2({ S7345 }),
  .A3({ S4995 }),
  .ZN({ S7346 })
);
NAND3_X1 #() 
NAND3_X1_323_ (
  .A1({ S7346 }),
  .A2({ S7341 }),
  .A3({ S2444 }),
  .ZN({ S7347 })
);
AOI22_X1 #() 
AOI22_X1_16_ (
  .A1({ S7029 }),
  .A2({ S25957[657] }),
  .B1({ S2665 }),
  .B2({ S2662 }),
  .ZN({ S7348 })
);
AOI21_X1 #() 
AOI21_X1_146_ (
  .A({ S25957[660] }),
  .B1({ S7348 }),
  .B2({ S6917 }),
  .ZN({ S7349 })
);
NAND2_X1 #() 
NAND2_X1_294_ (
  .A1({ S7349 }),
  .A2({ S7245 }),
  .ZN({ S7351 })
);
NAND2_X1 #() 
NAND2_X1_295_ (
  .A1({ S7112 }),
  .A2({ S6972 }),
  .ZN({ S7352 })
);
NAND3_X1 #() 
NAND3_X1_324_ (
  .A1({ S7242 }),
  .A2({ S25957[660] }),
  .A3({ S7352 }),
  .ZN({ S7353 })
);
NAND3_X1 #() 
NAND3_X1_325_ (
  .A1({ S7351 }),
  .A2({ S25957[661] }),
  .A3({ S7353 }),
  .ZN({ S7354 })
);
OAI211_X1 #() 
OAI211_X1_80_ (
  .A({ S7209 }),
  .B({ S25957[660] }),
  .C1({ S6954 }),
  .C2({ S7352 }),
  .ZN({ S7355 })
);
AND2_X1 #() 
AND2_X1_18_ (
  .A1({ S6930 }),
  .A2({ S6962 }),
  .ZN({ S7356 })
);
NAND3_X1 #() 
NAND3_X1_326_ (
  .A1({ S7073 }),
  .A2({ S6916 }),
  .A3({ S6922 }),
  .ZN({ S7357 })
);
NAND2_X1 #() 
NAND2_X1_296_ (
  .A1({ S7357 }),
  .A2({ S7356 }),
  .ZN({ S7358 })
);
NAND3_X1 #() 
NAND3_X1_327_ (
  .A1({ S7355 }),
  .A2({ S4995 }),
  .A3({ S7358 }),
  .ZN({ S7359 })
);
NAND3_X1 #() 
NAND3_X1_328_ (
  .A1({ S7359 }),
  .A2({ S7354 }),
  .A3({ S25957[662] }),
  .ZN({ S7360 })
);
NAND3_X1 #() 
NAND3_X1_329_ (
  .A1({ S7347 }),
  .A2({ S7360 }),
  .A3({ S25957[663] }),
  .ZN({ S7362 })
);
NAND3_X1 #() 
NAND3_X1_330_ (
  .A1({ S7122 }),
  .A2({ S6930 }),
  .A3({ S7032 }),
  .ZN({ S7363 })
);
OAI211_X1 #() 
OAI211_X1_81_ (
  .A({ S7241 }),
  .B({ S25957[660] }),
  .C1({ S6973 }),
  .C2({ S6946 }),
  .ZN({ S7364 })
);
NAND3_X1 #() 
NAND3_X1_331_ (
  .A1({ S7363 }),
  .A2({ S7364 }),
  .A3({ S25957[661] }),
  .ZN({ S7365 })
);
OAI211_X1 #() 
OAI211_X1_82_ (
  .A({ S110 }),
  .B({ S5359 }),
  .C1({ S6910 }),
  .C2({ S7029 }),
  .ZN({ S7366 })
);
OAI211_X1 #() 
OAI211_X1_83_ (
  .A({ S6930 }),
  .B({ S7366 }),
  .C1({ S7060 }),
  .C2({ S110 }),
  .ZN({ S7367 })
);
NAND2_X1 #() 
NAND2_X1_297_ (
  .A1({ S6908 }),
  .A2({ S110 }),
  .ZN({ S7368 })
);
NAND4_X1 #() 
NAND4_X1_27_ (
  .A1({ S7293 }),
  .A2({ S7368 }),
  .A3({ S7009 }),
  .A4({ S25957[660] }),
  .ZN({ S7369 })
);
NAND3_X1 #() 
NAND3_X1_332_ (
  .A1({ S7369 }),
  .A2({ S7367 }),
  .A3({ S4995 }),
  .ZN({ S7370 })
);
NAND3_X1 #() 
NAND3_X1_333_ (
  .A1({ S7370 }),
  .A2({ S7365 }),
  .A3({ S2444 }),
  .ZN({ S7371 })
);
NAND4_X1 #() 
NAND4_X1_28_ (
  .A1({ S7290 }),
  .A2({ S7126 }),
  .A3({ S6931 }),
  .A4({ S25957[659] }),
  .ZN({ S7373 })
);
AOI21_X1 #() 
AOI21_X1_147_ (
  .A({ S6930 }),
  .B1({ S7066 }),
  .B2({ S110 }),
  .ZN({ S7374 })
);
AOI22_X1 #() 
AOI22_X1_17_ (
  .A1({ S7374 }),
  .A2({ S7373 }),
  .B1({ S7097 }),
  .B2({ S7356 }),
  .ZN({ S7375 })
);
AOI21_X1 #() 
AOI21_X1_148_ (
  .A({ S6930 }),
  .B1({ S25957[659] }),
  .B2({ S5282 }),
  .ZN({ S7376 })
);
NAND3_X1 #() 
NAND3_X1_334_ (
  .A1({ S7376 }),
  .A2({ S6969 }),
  .A3({ S7054 }),
  .ZN({ S7377 })
);
NAND2_X1 #() 
NAND2_X1_298_ (
  .A1({ S7290 }),
  .A2({ S110 }),
  .ZN({ S7378 })
);
NAND3_X1 #() 
NAND3_X1_335_ (
  .A1({ S7133 }),
  .A2({ S6930 }),
  .A3({ S7378 }),
  .ZN({ S7379 })
);
NAND3_X1 #() 
NAND3_X1_336_ (
  .A1({ S7377 }),
  .A2({ S7379 }),
  .A3({ S4995 }),
  .ZN({ S7380 })
);
OAI211_X1 #() 
OAI211_X1_84_ (
  .A({ S7380 }),
  .B({ S25957[662] }),
  .C1({ S7375 }),
  .C2({ S4995 }),
  .ZN({ S7381 })
);
NAND3_X1 #() 
NAND3_X1_337_ (
  .A1({ S7371 }),
  .A2({ S7381 }),
  .A3({ S4797 }),
  .ZN({ S7382 })
);
AND3_X1 #() 
AND3_X1_14_ (
  .A1({ S7382 }),
  .A2({ S7362 }),
  .A3({ S24021 }),
  .ZN({ S7384 })
);
AOI21_X1 #() 
AOI21_X1_149_ (
  .A({ S24021 }),
  .B1({ S7382 }),
  .B2({ S7362 }),
  .ZN({ S7385 })
);
NOR2_X1 #() 
NOR2_X1_66_ (
  .A1({ S7384 }),
  .A2({ S7385 }),
  .ZN({ S7386 })
);
INV_X1 #() 
INV_X1_127_ (
  .A({ S7386 }),
  .ZN({ S25957[536] })
);
NAND2_X1 #() 
NAND2_X1_299_ (
  .A1({ S4725 }),
  .A2({ S4728 }),
  .ZN({ S25957[729] })
);
NAND2_X1 #() 
NAND2_X1_300_ (
  .A1({ S4724 }),
  .A2({ S4722 }),
  .ZN({ S25957[761] })
);
NAND2_X1 #() 
NAND2_X1_301_ (
  .A1({ S6943 }),
  .A2({ S25957[656] }),
  .ZN({ S7387 })
);
NAND3_X1 #() 
NAND3_X1_338_ (
  .A1({ S6959 }),
  .A2({ S25957[659] }),
  .A3({ S7387 }),
  .ZN({ S7388 })
);
AOI21_X1 #() 
AOI21_X1_150_ (
  .A({ S6930 }),
  .B1({ S7388 }),
  .B2({ S6994 }),
  .ZN({ S7389 })
);
NAND2_X1 #() 
NAND2_X1_302_ (
  .A1({ S7136 }),
  .A2({ S25957[659] }),
  .ZN({ S7390 })
);
AOI21_X1 #() 
AOI21_X1_151_ (
  .A({ S25957[660] }),
  .B1({ S7390 }),
  .B2({ S7320 }),
  .ZN({ S7392 })
);
OAI21_X1 #() 
OAI21_X1_186_ (
  .A({ S25957[661] }),
  .B1({ S7389 }),
  .B2({ S7392 }),
  .ZN({ S7393 })
);
NAND2_X1 #() 
NAND2_X1_303_ (
  .A1({ S7018 }),
  .A2({ S7218 }),
  .ZN({ S7394 })
);
NAND3_X1 #() 
NAND3_X1_339_ (
  .A1({ S7054 }),
  .A2({ S110 }),
  .A3({ S6969 }),
  .ZN({ S7395 })
);
NAND2_X1 #() 
NAND2_X1_304_ (
  .A1({ S7068 }),
  .A2({ S7395 }),
  .ZN({ S7396 })
);
NAND3_X1 #() 
NAND3_X1_340_ (
  .A1({ S7394 }),
  .A2({ S4995 }),
  .A3({ S7396 }),
  .ZN({ S7397 })
);
NAND3_X1 #() 
NAND3_X1_341_ (
  .A1({ S7397 }),
  .A2({ S7393 }),
  .A3({ S2444 }),
  .ZN({ S7398 })
);
NOR2_X1 #() 
NOR2_X1_67_ (
  .A1({ S6944 }),
  .A2({ S25957[659] }),
  .ZN({ S7399 })
);
NAND2_X1 #() 
NAND2_X1_305_ (
  .A1({ S7399 }),
  .A2({ S5282 }),
  .ZN({ S7400 })
);
NAND3_X1 #() 
NAND3_X1_342_ (
  .A1({ S7145 }),
  .A2({ S7400 }),
  .A3({ S25957[660] }),
  .ZN({ S7401 })
);
NAND2_X1 #() 
NAND2_X1_306_ (
  .A1({ S6908 }),
  .A2({ S5282 }),
  .ZN({ S7403 })
);
NAND2_X1 #() 
NAND2_X1_307_ (
  .A1({ S7316 }),
  .A2({ S7403 }),
  .ZN({ S7404 })
);
AOI21_X1 #() 
AOI21_X1_152_ (
  .A({ S25957[660] }),
  .B1({ S7086 }),
  .B2({ S25957[659] }),
  .ZN({ S7405 })
);
AOI21_X1 #() 
AOI21_X1_153_ (
  .A({ S25957[661] }),
  .B1({ S7405 }),
  .B2({ S7404 }),
  .ZN({ S7406 })
);
NAND2_X1 #() 
NAND2_X1_308_ (
  .A1({ S7406 }),
  .A2({ S7401 }),
  .ZN({ S7407 })
);
NAND3_X1 #() 
NAND3_X1_343_ (
  .A1({ S7042 }),
  .A2({ S25957[660] }),
  .A3({ S6998 }),
  .ZN({ S7408 })
);
AOI21_X1 #() 
AOI21_X1_154_ (
  .A({ S25957[660] }),
  .B1({ S6959 }),
  .B2({ S110 }),
  .ZN({ S7409 })
);
NAND2_X1 #() 
NAND2_X1_309_ (
  .A1({ S7373 }),
  .A2({ S7409 }),
  .ZN({ S7410 })
);
NAND3_X1 #() 
NAND3_X1_344_ (
  .A1({ S7410 }),
  .A2({ S25957[661] }),
  .A3({ S7408 }),
  .ZN({ S7411 })
);
NAND3_X1 #() 
NAND3_X1_345_ (
  .A1({ S7407 }),
  .A2({ S25957[662] }),
  .A3({ S7411 }),
  .ZN({ S7412 })
);
NAND3_X1 #() 
NAND3_X1_346_ (
  .A1({ S7398 }),
  .A2({ S7412 }),
  .A3({ S25957[663] }),
  .ZN({ S7414 })
);
AOI21_X1 #() 
AOI21_X1_155_ (
  .A({ S6930 }),
  .B1({ S7276 }),
  .B2({ S7228 }),
  .ZN({ S7415 })
);
OAI21_X1 #() 
OAI21_X1_187_ (
  .A({ S25957[661] }),
  .B1({ S7415 }),
  .B2({ S7015 }),
  .ZN({ S7416 })
);
NAND3_X1 #() 
NAND3_X1_347_ (
  .A1({ S7043 }),
  .A2({ S6909 }),
  .A3({ S6930 }),
  .ZN({ S7417 })
);
OAI211_X1 #() 
OAI211_X1_85_ (
  .A({ S6925 }),
  .B({ S6921 }),
  .C1({ S25957[659] }),
  .C2({ S6979 }),
  .ZN({ S7418 })
);
OAI211_X1 #() 
OAI211_X1_86_ (
  .A({ S7417 }),
  .B({ S4995 }),
  .C1({ S6930 }),
  .C2({ S7418 }),
  .ZN({ S7419 })
);
NAND3_X1 #() 
NAND3_X1_348_ (
  .A1({ S7416 }),
  .A2({ S2444 }),
  .A3({ S7419 }),
  .ZN({ S7420 })
);
INV_X1 #() 
INV_X1_128_ (
  .A({ S7126 }),
  .ZN({ S7421 })
);
OAI211_X1 #() 
OAI211_X1_87_ (
  .A({ S7373 }),
  .B({ S25957[660] }),
  .C1({ S7421 }),
  .C2({ S6932 }),
  .ZN({ S7422 })
);
AOI21_X1 #() 
AOI21_X1_156_ (
  .A({ S25957[660] }),
  .B1({ S7008 }),
  .B2({ S7112 }),
  .ZN({ S7423 })
);
AOI21_X1 #() 
AOI21_X1_157_ (
  .A({ S25957[661] }),
  .B1({ S7423 }),
  .B2({ S7075 }),
  .ZN({ S7425 })
);
NAND2_X1 #() 
NAND2_X1_310_ (
  .A1({ S7425 }),
  .A2({ S7422 }),
  .ZN({ S7426 })
);
OAI211_X1 #() 
OAI211_X1_88_ (
  .A({ S25957[660] }),
  .B({ S7311 }),
  .C1({ S7226 }),
  .C2({ S7029 }),
  .ZN({ S7427 })
);
NAND2_X1 #() 
NAND2_X1_311_ (
  .A1({ S6962 }),
  .A2({ S5359 }),
  .ZN({ S7428 })
);
AOI21_X1 #() 
AOI21_X1_158_ (
  .A({ S4995 }),
  .B1({ S7156 }),
  .B2({ S7428 }),
  .ZN({ S7429 })
);
AOI21_X1 #() 
AOI21_X1_159_ (
  .A({ S2444 }),
  .B1({ S7429 }),
  .B2({ S7427 }),
  .ZN({ S7430 })
);
NAND2_X1 #() 
NAND2_X1_312_ (
  .A1({ S7426 }),
  .A2({ S7430 }),
  .ZN({ S7431 })
);
NAND3_X1 #() 
NAND3_X1_349_ (
  .A1({ S7431 }),
  .A2({ S4797 }),
  .A3({ S7420 }),
  .ZN({ S7432 })
);
NAND3_X1 #() 
NAND3_X1_350_ (
  .A1({ S7414 }),
  .A2({ S25957[761] }),
  .A3({ S7432 }),
  .ZN({ S7433 })
);
INV_X1 #() 
INV_X1_129_ (
  .A({ S25957[761] }),
  .ZN({ S7434 })
);
AOI22_X1 #() 
AOI22_X1_18_ (
  .A1({ S7425 }),
  .A2({ S7422 }),
  .B1({ S7429 }),
  .B2({ S7427 }),
  .ZN({ S7436 })
);
INV_X1 #() 
INV_X1_130_ (
  .A({ S7015 }),
  .ZN({ S7437 })
);
NAND2_X1 #() 
NAND2_X1_313_ (
  .A1({ S7276 }),
  .A2({ S7228 }),
  .ZN({ S7438 })
);
NAND2_X1 #() 
NAND2_X1_314_ (
  .A1({ S7438 }),
  .A2({ S25957[660] }),
  .ZN({ S7439 })
);
NAND3_X1 #() 
NAND3_X1_351_ (
  .A1({ S7439 }),
  .A2({ S7437 }),
  .A3({ S25957[661] }),
  .ZN({ S7440 })
);
NAND2_X1 #() 
NAND2_X1_315_ (
  .A1({ S7418 }),
  .A2({ S25957[660] }),
  .ZN({ S7441 })
);
NAND2_X1 #() 
NAND2_X1_316_ (
  .A1({ S7043 }),
  .A2({ S6909 }),
  .ZN({ S7442 })
);
NAND2_X1 #() 
NAND2_X1_317_ (
  .A1({ S7442 }),
  .A2({ S6930 }),
  .ZN({ S7443 })
);
NAND3_X1 #() 
NAND3_X1_352_ (
  .A1({ S7443 }),
  .A2({ S4995 }),
  .A3({ S7441 }),
  .ZN({ S7444 })
);
NAND3_X1 #() 
NAND3_X1_353_ (
  .A1({ S7440 }),
  .A2({ S2444 }),
  .A3({ S7444 }),
  .ZN({ S7445 })
);
OAI211_X1 #() 
OAI211_X1_89_ (
  .A({ S7445 }),
  .B({ S4797 }),
  .C1({ S7436 }),
  .C2({ S2444 }),
  .ZN({ S7447 })
);
AOI21_X1 #() 
AOI21_X1_160_ (
  .A({ S4995 }),
  .B1({ S7373 }),
  .B2({ S7409 }),
  .ZN({ S7448 })
);
AOI22_X1 #() 
AOI22_X1_19_ (
  .A1({ S7406 }),
  .A2({ S7401 }),
  .B1({ S7448 }),
  .B2({ S7408 }),
  .ZN({ S7449 })
);
AOI22_X1 #() 
AOI22_X1_20_ (
  .A1({ S7003 }),
  .A2({ S7387 }),
  .B1({ S6993 }),
  .B2({ S110 }),
  .ZN({ S7450 })
);
NAND3_X1 #() 
NAND3_X1_354_ (
  .A1({ S14 }),
  .A2({ S110 }),
  .A3({ S6943 }),
  .ZN({ S7451 })
);
NAND3_X1 #() 
NAND3_X1_355_ (
  .A1({ S7058 }),
  .A2({ S6930 }),
  .A3({ S7451 }),
  .ZN({ S7452 })
);
OAI211_X1 #() 
OAI211_X1_90_ (
  .A({ S7452 }),
  .B({ S25957[661] }),
  .C1({ S7450 }),
  .C2({ S6930 }),
  .ZN({ S7453 })
);
AOI22_X1 #() 
AOI22_X1_21_ (
  .A1({ S7018 }),
  .A2({ S7218 }),
  .B1({ S7068 }),
  .B2({ S7395 }),
  .ZN({ S7454 })
);
OAI211_X1 #() 
OAI211_X1_91_ (
  .A({ S7453 }),
  .B({ S2444 }),
  .C1({ S7454 }),
  .C2({ S25957[661] }),
  .ZN({ S7455 })
);
OAI211_X1 #() 
OAI211_X1_92_ (
  .A({ S7455 }),
  .B({ S25957[663] }),
  .C1({ S2444 }),
  .C2({ S7449 }),
  .ZN({ S7456 })
);
NAND3_X1 #() 
NAND3_X1_356_ (
  .A1({ S7456 }),
  .A2({ S7434 }),
  .A3({ S7447 }),
  .ZN({ S7458 })
);
NAND3_X1 #() 
NAND3_X1_357_ (
  .A1({ S7458 }),
  .A2({ S25957[729] }),
  .A3({ S7433 }),
  .ZN({ S7459 })
);
INV_X1 #() 
INV_X1_131_ (
  .A({ S25957[729] }),
  .ZN({ S7460 })
);
NAND3_X1 #() 
NAND3_X1_358_ (
  .A1({ S7414 }),
  .A2({ S7434 }),
  .A3({ S7432 }),
  .ZN({ S7461 })
);
NAND3_X1 #() 
NAND3_X1_359_ (
  .A1({ S7456 }),
  .A2({ S25957[761] }),
  .A3({ S7447 }),
  .ZN({ S7462 })
);
NAND3_X1 #() 
NAND3_X1_360_ (
  .A1({ S7462 }),
  .A2({ S7460 }),
  .A3({ S7461 }),
  .ZN({ S7463 })
);
NAND3_X1 #() 
NAND3_X1_361_ (
  .A1({ S7459 }),
  .A2({ S7463 }),
  .A3({ S3527 }),
  .ZN({ S7464 })
);
NAND3_X1 #() 
NAND3_X1_362_ (
  .A1({ S7458 }),
  .A2({ S7460 }),
  .A3({ S7433 }),
  .ZN({ S7465 })
);
NAND3_X1 #() 
NAND3_X1_363_ (
  .A1({ S7462 }),
  .A2({ S25957[729] }),
  .A3({ S7461 }),
  .ZN({ S7466 })
);
NAND3_X1 #() 
NAND3_X1_364_ (
  .A1({ S7465 }),
  .A2({ S7466 }),
  .A3({ S25957[793] }),
  .ZN({ S7467 })
);
NAND2_X1 #() 
NAND2_X1_318_ (
  .A1({ S7464 }),
  .A2({ S7467 }),
  .ZN({ S25957[537] })
);
NOR2_X1 #() 
NOR2_X1_68_ (
  .A1({ S4784 }),
  .A2({ S4787 }),
  .ZN({ S7469 })
);
INV_X1 #() 
INV_X1_132_ (
  .A({ S7469 }),
  .ZN({ S25957[730] })
);
NAND2_X1 #() 
NAND2_X1_319_ (
  .A1({ S2221 }),
  .A2({ S2220 }),
  .ZN({ S25957[890] })
);
NOR2_X1 #() 
NOR2_X1_69_ (
  .A1({ S4786 }),
  .A2({ S4785 }),
  .ZN({ S7470 })
);
XOR2_X1 #() 
XOR2_X1_5_ (
  .A({ S7470 }),
  .B({ S25957[890] }),
  .Z({ S25957[762] })
);
INV_X1 #() 
INV_X1_133_ (
  .A({ S25957[762] }),
  .ZN({ S7471 })
);
NAND3_X1 #() 
NAND3_X1_365_ (
  .A1({ S25957[659] }),
  .A2({ S25957[656] }),
  .A3({ S6939 }),
  .ZN({ S7472 })
);
NAND3_X1 #() 
NAND3_X1_366_ (
  .A1({ S7043 }),
  .A2({ S7472 }),
  .A3({ S25957[660] }),
  .ZN({ S7473 })
);
NAND4_X1 #() 
NAND4_X1_29_ (
  .A1({ S7217 }),
  .A2({ S7257 }),
  .A3({ S6933 }),
  .A4({ S6930 }),
  .ZN({ S7474 })
);
NAND3_X1 #() 
NAND3_X1_367_ (
  .A1({ S7474 }),
  .A2({ S7473 }),
  .A3({ S25957[661] }),
  .ZN({ S7476 })
);
NAND2_X1 #() 
NAND2_X1_320_ (
  .A1({ S6979 }),
  .A2({ S110 }),
  .ZN({ S7477 })
);
NAND4_X1 #() 
NAND4_X1_30_ (
  .A1({ S6916 }),
  .A2({ S25957[657] }),
  .A3({ S2665 }),
  .A4({ S2662 }),
  .ZN({ S7478 })
);
NAND3_X1 #() 
NAND3_X1_368_ (
  .A1({ S7478 }),
  .A2({ S25957[660] }),
  .A3({ S7477 }),
  .ZN({ S7479 })
);
OAI211_X1 #() 
OAI211_X1_93_ (
  .A({ S7053 }),
  .B({ S6930 }),
  .C1({ S6922 }),
  .C2({ S6931 }),
  .ZN({ S7480 })
);
NAND3_X1 #() 
NAND3_X1_369_ (
  .A1({ S7480 }),
  .A2({ S7479 }),
  .A3({ S4995 }),
  .ZN({ S7481 })
);
NAND3_X1 #() 
NAND3_X1_370_ (
  .A1({ S7476 }),
  .A2({ S7481 }),
  .A3({ S2444 }),
  .ZN({ S7482 })
);
NAND3_X1 #() 
NAND3_X1_371_ (
  .A1({ S7176 }),
  .A2({ S7161 }),
  .A3({ S25957[659] }),
  .ZN({ S7483 })
);
NOR2_X1 #() 
NOR2_X1_70_ (
  .A1({ S7399 }),
  .A2({ S25957[660] }),
  .ZN({ S7484 })
);
NAND2_X1 #() 
NAND2_X1_321_ (
  .A1({ S7483 }),
  .A2({ S7484 }),
  .ZN({ S7485 })
);
NAND4_X1 #() 
NAND4_X1_31_ (
  .A1({ S6913 }),
  .A2({ S6969 }),
  .A3({ S110 }),
  .A4({ S14 }),
  .ZN({ S7487 })
);
AOI21_X1 #() 
AOI21_X1_161_ (
  .A({ S6930 }),
  .B1({ S7220 }),
  .B2({ S25957[659] }),
  .ZN({ S7488 })
);
AOI21_X1 #() 
AOI21_X1_162_ (
  .A({ S4995 }),
  .B1({ S7488 }),
  .B2({ S7487 }),
  .ZN({ S7489 })
);
NAND2_X1 #() 
NAND2_X1_322_ (
  .A1({ S7489 }),
  .A2({ S7485 }),
  .ZN({ S7490 })
);
OAI211_X1 #() 
OAI211_X1_94_ (
  .A({ S6930 }),
  .B({ S7368 }),
  .C1({ S6980 }),
  .C2({ S110 }),
  .ZN({ S7491 })
);
NAND2_X1 #() 
NAND2_X1_323_ (
  .A1({ S6918 }),
  .A2({ S6964 }),
  .ZN({ S7492 })
);
NAND2_X1 #() 
NAND2_X1_324_ (
  .A1({ S7492 }),
  .A2({ S7178 }),
  .ZN({ S7493 })
);
NAND3_X1 #() 
NAND3_X1_372_ (
  .A1({ S7493 }),
  .A2({ S4995 }),
  .A3({ S7491 }),
  .ZN({ S7494 })
);
NAND3_X1 #() 
NAND3_X1_373_ (
  .A1({ S7490 }),
  .A2({ S7494 }),
  .A3({ S25957[662] }),
  .ZN({ S7495 })
);
NAND3_X1 #() 
NAND3_X1_374_ (
  .A1({ S7495 }),
  .A2({ S25957[663] }),
  .A3({ S7482 }),
  .ZN({ S7496 })
);
NAND3_X1 #() 
NAND3_X1_375_ (
  .A1({ S7176 }),
  .A2({ S7144 }),
  .A3({ S25957[659] }),
  .ZN({ S7498 })
);
OAI21_X1 #() 
OAI21_X1_188_ (
  .A({ S110 }),
  .B1({ S6908 }),
  .B2({ S5282 }),
  .ZN({ S7499 })
);
NAND3_X1 #() 
NAND3_X1_376_ (
  .A1({ S6938 }),
  .A2({ S25957[659] }),
  .A3({ S6939 }),
  .ZN({ S7500 })
);
AOI21_X1 #() 
AOI21_X1_163_ (
  .A({ S6930 }),
  .B1({ S7500 }),
  .B2({ S7499 }),
  .ZN({ S7501 })
);
OAI21_X1 #() 
OAI21_X1_189_ (
  .A({ S6930 }),
  .B1({ S6987 }),
  .B2({ S7067 }),
  .ZN({ S7502 })
);
INV_X1 #() 
INV_X1_134_ (
  .A({ S7502 }),
  .ZN({ S7503 })
);
AOI21_X1 #() 
AOI21_X1_164_ (
  .A({ S7501 }),
  .B1({ S7498 }),
  .B2({ S7503 }),
  .ZN({ S7504 })
);
NAND3_X1 #() 
NAND3_X1_377_ (
  .A1({ S25957[659] }),
  .A2({ S6943 }),
  .A3({ S6972 }),
  .ZN({ S7505 })
);
NAND3_X1 #() 
NAND3_X1_378_ (
  .A1({ S7209 }),
  .A2({ S6930 }),
  .A3({ S7505 }),
  .ZN({ S7506 })
);
NAND2_X1 #() 
NAND2_X1_325_ (
  .A1({ S6944 }),
  .A2({ S110 }),
  .ZN({ S7507 })
);
OAI211_X1 #() 
OAI211_X1_95_ (
  .A({ S25957[659] }),
  .B({ S6921 }),
  .C1({ S25957[656] }),
  .C2({ S6979 }),
  .ZN({ S7509 })
);
NAND4_X1 #() 
NAND4_X1_32_ (
  .A1({ S7509 }),
  .A2({ S7499 }),
  .A3({ S7507 }),
  .A4({ S25957[660] }),
  .ZN({ S7510 })
);
NAND3_X1 #() 
NAND3_X1_379_ (
  .A1({ S7506 }),
  .A2({ S4995 }),
  .A3({ S7510 }),
  .ZN({ S7511 })
);
OAI211_X1 #() 
OAI211_X1_96_ (
  .A({ S7511 }),
  .B({ S25957[662] }),
  .C1({ S7504 }),
  .C2({ S4995 }),
  .ZN({ S7512 })
);
NAND3_X1 #() 
NAND3_X1_380_ (
  .A1({ S6959 }),
  .A2({ S7136 }),
  .A3({ S25957[659] }),
  .ZN({ S7513 })
);
OAI21_X1 #() 
OAI21_X1_190_ (
  .A({ S7478 }),
  .B1({ S7153 }),
  .B2({ S6991 }),
  .ZN({ S7514 })
);
AOI22_X1 #() 
AOI22_X1_22_ (
  .A1({ S7349 }),
  .A2({ S7513 }),
  .B1({ S7514 }),
  .B2({ S25957[660] }),
  .ZN({ S7515 })
);
AOI211_X1 #() 
AOI211_X1_3_ (
  .A({ S6908 }),
  .B({ S25957[659] }),
  .C1({ S7010 }),
  .C2({ S14 }),
  .ZN({ S7516 })
);
AOI21_X1 #() 
AOI21_X1_165_ (
  .A({ S25957[660] }),
  .B1({ S7109 }),
  .B2({ S110 }),
  .ZN({ S7517 })
);
NAND4_X1 #() 
NAND4_X1_33_ (
  .A1({ S7126 }),
  .A2({ S6939 }),
  .A3({ S6931 }),
  .A4({ S25957[659] }),
  .ZN({ S7518 })
);
NAND2_X1 #() 
NAND2_X1_326_ (
  .A1({ S7517 }),
  .A2({ S7518 }),
  .ZN({ S7520 })
);
NAND2_X1 #() 
NAND2_X1_327_ (
  .A1({ S25957[659] }),
  .A2({ S6921 }),
  .ZN({ S7521 })
);
NOR2_X1 #() 
NOR2_X1_71_ (
  .A1({ S6931 }),
  .A2({ S25957[657] }),
  .ZN({ S7522 })
);
OAI21_X1 #() 
OAI21_X1_191_ (
  .A({ S25957[660] }),
  .B1({ S7521 }),
  .B2({ S7522 }),
  .ZN({ S7523 })
);
OAI211_X1 #() 
OAI211_X1_97_ (
  .A({ S7520 }),
  .B({ S25957[661] }),
  .C1({ S7516 }),
  .C2({ S7523 }),
  .ZN({ S7524 })
);
OAI211_X1 #() 
OAI211_X1_98_ (
  .A({ S7524 }),
  .B({ S2444 }),
  .C1({ S25957[661] }),
  .C2({ S7515 }),
  .ZN({ S7525 })
);
NAND3_X1 #() 
NAND3_X1_381_ (
  .A1({ S7525 }),
  .A2({ S7512 }),
  .A3({ S4797 }),
  .ZN({ S7526 })
);
NAND3_X1 #() 
NAND3_X1_382_ (
  .A1({ S7526 }),
  .A2({ S7471 }),
  .A3({ S7496 }),
  .ZN({ S7527 })
);
NOR3_X1 #() 
NOR3_X1_11_ (
  .A1({ S6954 }),
  .A2({ S6908 }),
  .A3({ S110 }),
  .ZN({ S7528 })
);
OAI21_X1 #() 
OAI21_X1_192_ (
  .A({ S25957[660] }),
  .B1({ S7528 }),
  .B2({ S7316 }),
  .ZN({ S7529 })
);
OAI21_X1 #() 
OAI21_X1_193_ (
  .A({ S7529 }),
  .B1({ S6942 }),
  .B2({ S7502 }),
  .ZN({ S7531 })
);
NOR2_X1 #() 
NOR2_X1_72_ (
  .A1({ S7316 }),
  .A2({ S6930 }),
  .ZN({ S7532 })
);
AOI22_X1 #() 
AOI22_X1_23_ (
  .A1({ S6985 }),
  .A2({ S7054 }),
  .B1({ S6944 }),
  .B2({ S110 }),
  .ZN({ S7533 })
);
AOI21_X1 #() 
AOI21_X1_166_ (
  .A({ S25957[661] }),
  .B1({ S7533 }),
  .B2({ S7532 }),
  .ZN({ S7534 })
);
AOI22_X1 #() 
AOI22_X1_24_ (
  .A1({ S7531 }),
  .A2({ S25957[661] }),
  .B1({ S7534 }),
  .B2({ S7506 }),
  .ZN({ S7535 })
);
AOI21_X1 #() 
AOI21_X1_167_ (
  .A({ S6930 }),
  .B1({ S6985 }),
  .B2({ S7403 }),
  .ZN({ S7536 })
);
AOI22_X1 #() 
AOI22_X1_25_ (
  .A1({ S7536 }),
  .A2({ S7274 }),
  .B1({ S7517 }),
  .B2({ S7518 }),
  .ZN({ S7537 })
);
NAND2_X1 #() 
NAND2_X1_328_ (
  .A1({ S7514 }),
  .A2({ S25957[660] }),
  .ZN({ S7538 })
);
NAND3_X1 #() 
NAND3_X1_383_ (
  .A1({ S7513 }),
  .A2({ S6930 }),
  .A3({ S7487 }),
  .ZN({ S7539 })
);
NAND3_X1 #() 
NAND3_X1_384_ (
  .A1({ S7538 }),
  .A2({ S7539 }),
  .A3({ S4995 }),
  .ZN({ S7540 })
);
OAI211_X1 #() 
OAI211_X1_99_ (
  .A({ S7540 }),
  .B({ S2444 }),
  .C1({ S4995 }),
  .C2({ S7537 }),
  .ZN({ S7542 })
);
OAI211_X1 #() 
OAI211_X1_100_ (
  .A({ S7542 }),
  .B({ S4797 }),
  .C1({ S7535 }),
  .C2({ S2444 }),
  .ZN({ S7543 })
);
AOI21_X1 #() 
AOI21_X1_168_ (
  .A({ S25957[661] }),
  .B1({ S7492 }),
  .B2({ S7178 }),
  .ZN({ S7544 })
);
AOI22_X1 #() 
AOI22_X1_26_ (
  .A1({ S7544 }),
  .A2({ S7491 }),
  .B1({ S7489 }),
  .B2({ S7485 }),
  .ZN({ S7545 })
);
NAND2_X1 #() 
NAND2_X1_329_ (
  .A1({ S7476 }),
  .A2({ S7481 }),
  .ZN({ S7546 })
);
NAND2_X1 #() 
NAND2_X1_330_ (
  .A1({ S7546 }),
  .A2({ S2444 }),
  .ZN({ S7547 })
);
OAI211_X1 #() 
OAI211_X1_101_ (
  .A({ S7547 }),
  .B({ S25957[663] }),
  .C1({ S7545 }),
  .C2({ S2444 }),
  .ZN({ S7548 })
);
NAND3_X1 #() 
NAND3_X1_385_ (
  .A1({ S7543 }),
  .A2({ S7548 }),
  .A3({ S25957[762] }),
  .ZN({ S7549 })
);
NAND3_X1 #() 
NAND3_X1_386_ (
  .A1({ S7549 }),
  .A2({ S25957[730] }),
  .A3({ S7527 }),
  .ZN({ S7550 })
);
NAND3_X1 #() 
NAND3_X1_387_ (
  .A1({ S7526 }),
  .A2({ S25957[762] }),
  .A3({ S7496 }),
  .ZN({ S7551 })
);
NAND3_X1 #() 
NAND3_X1_388_ (
  .A1({ S7543 }),
  .A2({ S7548 }),
  .A3({ S7471 }),
  .ZN({ S7553 })
);
NAND3_X1 #() 
NAND3_X1_389_ (
  .A1({ S7553 }),
  .A2({ S7469 }),
  .A3({ S7551 }),
  .ZN({ S7554 })
);
NAND3_X1 #() 
NAND3_X1_390_ (
  .A1({ S7550 }),
  .A2({ S7554 }),
  .A3({ S3488 }),
  .ZN({ S7555 })
);
NAND3_X1 #() 
NAND3_X1_391_ (
  .A1({ S7553 }),
  .A2({ S25957[730] }),
  .A3({ S7551 }),
  .ZN({ S7556 })
);
NAND3_X1 #() 
NAND3_X1_392_ (
  .A1({ S7549 }),
  .A2({ S7469 }),
  .A3({ S7527 }),
  .ZN({ S7557 })
);
NAND3_X1 #() 
NAND3_X1_393_ (
  .A1({ S7556 }),
  .A2({ S7557 }),
  .A3({ S25957[794] }),
  .ZN({ S7558 })
);
AND2_X1 #() 
AND2_X1_19_ (
  .A1({ S7558 }),
  .A2({ S7555 }),
  .ZN({ S25957[538] })
);
AOI22_X1 #() 
AOI22_X1_27_ (
  .A1({ S6012 }),
  .A2({ S6009 }),
  .B1({ S6096 }),
  .B2({ S6099 }),
  .ZN({ S16 })
);
NAND4_X1 #() 
NAND4_X1_34_ (
  .A1({ S6012 }),
  .A2({ S6009 }),
  .A3({ S6096 }),
  .A4({ S6099 }),
  .ZN({ S17 })
);
INV_X1 #() 
INV_X1_135_ (
  .A({ S25957[567] }),
  .ZN({ S7559 })
);
XOR2_X1 #() 
XOR2_X1_6_ (
  .A({ S25957[631] }),
  .B({ S25957[727] }),
  .Z({ S25957[599] })
);
INV_X1 #() 
INV_X1_136_ (
  .A({ S25957[599] }),
  .ZN({ S7561 })
);
INV_X1 #() 
INV_X1_137_ (
  .A({ S25957[527] }),
  .ZN({ S7562 })
);
OAI21_X1 #() 
OAI21_X1_194_ (
  .A({ S25957[648] }),
  .B1({ S6010 }),
  .B2({ S6011 }),
  .ZN({ S7563 })
);
NAND3_X1 #() 
NAND3_X1_394_ (
  .A1({ S6003 }),
  .A2({ S6008 }),
  .A3({ S4794 }),
  .ZN({ S7564 })
);
AOI21_X1 #() 
AOI21_X1_169_ (
  .A({ S25957[649] }),
  .B1({ S6097 }),
  .B2({ S6098 }),
  .ZN({ S7565 })
);
AOI21_X1 #() 
AOI21_X1_170_ (
  .A({ S4806 }),
  .B1({ S6091 }),
  .B2({ S6095 }),
  .ZN({ S7566 })
);
OAI211_X1 #() 
OAI211_X1_102_ (
  .A({ S7563 }),
  .B({ S7564 }),
  .C1({ S7566 }),
  .C2({ S7565 }),
  .ZN({ S7567 })
);
NAND3_X1 #() 
NAND3_X1_395_ (
  .A1({ S7567 }),
  .A2({ S25957[522] }),
  .A3({ S17 }),
  .ZN({ S7568 })
);
NAND3_X1 #() 
NAND3_X1_396_ (
  .A1({ S6179 }),
  .A2({ S25957[650] }),
  .A3({ S6178 }),
  .ZN({ S7569 })
);
NAND3_X1 #() 
NAND3_X1_397_ (
  .A1({ S6172 }),
  .A2({ S4816 }),
  .A3({ S6175 }),
  .ZN({ S7571 })
);
NAND2_X1 #() 
NAND2_X1_331_ (
  .A1({ S7569 }),
  .A2({ S7571 }),
  .ZN({ S7572 })
);
AOI21_X1 #() 
AOI21_X1_171_ (
  .A({ S25957[523] }),
  .B1({ S16 }),
  .B2({ S7572 }),
  .ZN({ S7573 })
);
NAND2_X1 #() 
NAND2_X1_332_ (
  .A1({ S7573 }),
  .A2({ S7568 }),
  .ZN({ S7574 })
);
OR2_X1 #() 
OR2_X1_6_ (
  .A1({ S5841 }),
  .A2({ S5840 }),
  .ZN({ S7575 })
);
NAND2_X1 #() 
NAND2_X1_333_ (
  .A1({ S7563 }),
  .A2({ S7564 }),
  .ZN({ S7576 })
);
NAND4_X1 #() 
NAND4_X1_35_ (
  .A1({ S7576 }),
  .A2({ S25957[521] }),
  .A3({ S7569 }),
  .A4({ S7571 }),
  .ZN({ S7577 })
);
AOI21_X1 #() 
AOI21_X1_172_ (
  .A({ S7575 }),
  .B1({ S7577 }),
  .B2({ S25957[523] }),
  .ZN({ S7578 })
);
OAI211_X1 #() 
OAI211_X1_103_ (
  .A({ S6009 }),
  .B({ S6012 }),
  .C1({ S7566 }),
  .C2({ S7565 }),
  .ZN({ S7579 })
);
NAND4_X1 #() 
NAND4_X1_36_ (
  .A1({ S7563 }),
  .A2({ S7564 }),
  .A3({ S6096 }),
  .A4({ S6099 }),
  .ZN({ S7580 })
);
NAND4_X1 #() 
NAND4_X1_37_ (
  .A1({ S7579 }),
  .A2({ S7580 }),
  .A3({ S9 }),
  .A4({ S25957[522] }),
  .ZN({ S7582 })
);
NAND2_X1 #() 
NAND2_X1_334_ (
  .A1({ S7567 }),
  .A2({ S25957[522] }),
  .ZN({ S7583 })
);
INV_X1 #() 
INV_X1_138_ (
  .A({ S7583 }),
  .ZN({ S7584 })
);
AOI21_X1 #() 
AOI21_X1_173_ (
  .A({ S25957[524] }),
  .B1({ S7584 }),
  .B2({ S25957[523] }),
  .ZN({ S7585 })
);
AOI22_X1 #() 
AOI22_X1_28_ (
  .A1({ S7585 }),
  .A2({ S7582 }),
  .B1({ S7574 }),
  .B2({ S7578 }),
  .ZN({ S7586 })
);
NAND3_X1 #() 
NAND3_X1_398_ (
  .A1({ S25957[521] }),
  .A2({ S6177 }),
  .A3({ S6180 }),
  .ZN({ S7587 })
);
NOR2_X1 #() 
NOR2_X1_73_ (
  .A1({ S7565 }),
  .A2({ S7566 }),
  .ZN({ S7588 })
);
AOI21_X1 #() 
AOI21_X1_174_ (
  .A({ S9 }),
  .B1({ S7588 }),
  .B2({ S25957[520] }),
  .ZN({ S7589 })
);
NAND2_X1 #() 
NAND2_X1_335_ (
  .A1({ S7589 }),
  .A2({ S7587 }),
  .ZN({ S7590 })
);
NAND2_X1 #() 
NAND2_X1_336_ (
  .A1({ S7567 }),
  .A2({ S7572 }),
  .ZN({ S7591 })
);
AOI21_X1 #() 
AOI21_X1_175_ (
  .A({ S25957[523] }),
  .B1({ S25957[522] }),
  .B2({ S25957[521] }),
  .ZN({ S7593 })
);
NAND2_X1 #() 
NAND2_X1_337_ (
  .A1({ S7593 }),
  .A2({ S7591 }),
  .ZN({ S7594 })
);
AOI21_X1 #() 
AOI21_X1_176_ (
  .A({ S25957[524] }),
  .B1({ S7594 }),
  .B2({ S7590 }),
  .ZN({ S7595 })
);
NAND4_X1 #() 
NAND4_X1_38_ (
  .A1({ S6177 }),
  .A2({ S6180 }),
  .A3({ S6096 }),
  .A4({ S6099 }),
  .ZN({ S7596 })
);
AOI21_X1 #() 
AOI21_X1_177_ (
  .A({ S9 }),
  .B1({ S25957[522] }),
  .B2({ S25957[520] }),
  .ZN({ S7597 })
);
NAND2_X1 #() 
NAND2_X1_338_ (
  .A1({ S7597 }),
  .A2({ S7596 }),
  .ZN({ S7598 })
);
NAND2_X1 #() 
NAND2_X1_339_ (
  .A1({ S25957[520] }),
  .A2({ S9 }),
  .ZN({ S7599 })
);
NAND3_X1 #() 
NAND3_X1_399_ (
  .A1({ S7598 }),
  .A2({ S25957[524] }),
  .A3({ S7599 }),
  .ZN({ S7600 })
);
INV_X1 #() 
INV_X1_139_ (
  .A({ S7600 }),
  .ZN({ S7601 })
);
OAI21_X1 #() 
OAI21_X1_195_ (
  .A({ S25957[525] }),
  .B1({ S7601 }),
  .B2({ S7595 }),
  .ZN({ S7602 })
);
OAI21_X1 #() 
OAI21_X1_196_ (
  .A({ S7602 }),
  .B1({ S7586 }),
  .B2({ S25957[525] }),
  .ZN({ S7604 })
);
INV_X1 #() 
INV_X1_140_ (
  .A({ S25957[525] }),
  .ZN({ S7605 })
);
NAND4_X1 #() 
NAND4_X1_39_ (
  .A1({ S7569 }),
  .A2({ S7571 }),
  .A3({ S7563 }),
  .A4({ S7564 }),
  .ZN({ S7606 })
);
AOI22_X1 #() 
AOI22_X1_29_ (
  .A1({ S7606 }),
  .A2({ S7580 }),
  .B1({ S25957[522] }),
  .B2({ S7588 }),
  .ZN({ S7607 })
);
OAI21_X1 #() 
OAI21_X1_197_ (
  .A({ S7575 }),
  .B1({ S7607 }),
  .B2({ S25957[523] }),
  .ZN({ S7608 })
);
AOI21_X1 #() 
AOI21_X1_178_ (
  .A({ S7608 }),
  .B1({ S7597 }),
  .B2({ S7587 }),
  .ZN({ S7609 })
);
NAND4_X1 #() 
NAND4_X1_40_ (
  .A1({ S6177 }),
  .A2({ S6180 }),
  .A3({ S6009 }),
  .A4({ S6012 }),
  .ZN({ S7610 })
);
NAND3_X1 #() 
NAND3_X1_400_ (
  .A1({ S7579 }),
  .A2({ S25957[522] }),
  .A3({ S7580 }),
  .ZN({ S7611 })
);
AOI21_X1 #() 
AOI21_X1_179_ (
  .A({ S25957[523] }),
  .B1({ S7611 }),
  .B2({ S7610 }),
  .ZN({ S7612 })
);
NAND3_X1 #() 
NAND3_X1_401_ (
  .A1({ S7579 }),
  .A2({ S7572 }),
  .A3({ S7580 }),
  .ZN({ S7613 })
);
AOI21_X1 #() 
AOI21_X1_180_ (
  .A({ S9 }),
  .B1({ S7613 }),
  .B2({ S7583 }),
  .ZN({ S7615 })
);
NOR3_X1 #() 
NOR3_X1_12_ (
  .A1({ S7615 }),
  .A2({ S7612 }),
  .A3({ S7575 }),
  .ZN({ S7616 })
);
OAI21_X1 #() 
OAI21_X1_198_ (
  .A({ S7605 }),
  .B1({ S7609 }),
  .B2({ S7616 }),
  .ZN({ S7617 })
);
NAND3_X1 #() 
NAND3_X1_402_ (
  .A1({ S25957[522] }),
  .A2({ S25957[523] }),
  .A3({ S25957[521] }),
  .ZN({ S7618 })
);
NAND2_X1 #() 
NAND2_X1_340_ (
  .A1({ S7618 }),
  .A2({ S25957[524] }),
  .ZN({ S7619 })
);
NAND4_X1 #() 
NAND4_X1_41_ (
  .A1({ S7569 }),
  .A2({ S7571 }),
  .A3({ S6009 }),
  .A4({ S6012 }),
  .ZN({ S7620 })
);
NAND3_X1 #() 
NAND3_X1_403_ (
  .A1({ S7620 }),
  .A2({ S7567 }),
  .A3({ S25957[523] }),
  .ZN({ S7621 })
);
AOI21_X1 #() 
AOI21_X1_181_ (
  .A({ S25957[520] }),
  .B1({ S25957[522] }),
  .B2({ S7588 }),
  .ZN({ S7622 })
);
OAI21_X1 #() 
OAI21_X1_199_ (
  .A({ S7621 }),
  .B1({ S7622 }),
  .B2({ S25957[523] }),
  .ZN({ S7623 })
);
NAND4_X1 #() 
NAND4_X1_42_ (
  .A1({ S7569 }),
  .A2({ S7571 }),
  .A3({ S6096 }),
  .A4({ S6099 }),
  .ZN({ S7624 })
);
NAND2_X1 #() 
NAND2_X1_341_ (
  .A1({ S7580 }),
  .A2({ S7572 }),
  .ZN({ S7626 })
);
NAND3_X1 #() 
NAND3_X1_404_ (
  .A1({ S7626 }),
  .A2({ S25957[523] }),
  .A3({ S7624 }),
  .ZN({ S7627 })
);
OAI21_X1 #() 
OAI21_X1_200_ (
  .A({ S9 }),
  .B1({ S16 }),
  .B2({ S7572 }),
  .ZN({ S7628 })
);
NAND3_X1 #() 
NAND3_X1_405_ (
  .A1({ S7627 }),
  .A2({ S7575 }),
  .A3({ S7628 }),
  .ZN({ S7629 })
);
OAI211_X1 #() 
OAI211_X1_104_ (
  .A({ S25957[525] }),
  .B({ S7629 }),
  .C1({ S7623 }),
  .C2({ S7619 }),
  .ZN({ S7630 })
);
NAND2_X1 #() 
NAND2_X1_342_ (
  .A1({ S7617 }),
  .A2({ S7630 }),
  .ZN({ S7631 })
);
NAND2_X1 #() 
NAND2_X1_343_ (
  .A1({ S7631 }),
  .A2({ S25957[526] }),
  .ZN({ S7632 })
);
OAI211_X1 #() 
OAI211_X1_105_ (
  .A({ S7632 }),
  .B({ S7562 }),
  .C1({ S25957[526] }),
  .C2({ S7604 }),
  .ZN({ S7633 })
);
AOI21_X1 #() 
AOI21_X1_182_ (
  .A({ S25957[523] }),
  .B1({ S7572 }),
  .B2({ S7576 }),
  .ZN({ S7634 })
);
INV_X1 #() 
INV_X1_141_ (
  .A({ S7634 }),
  .ZN({ S7635 })
);
NAND3_X1 #() 
NAND3_X1_406_ (
  .A1({ S7572 }),
  .A2({ S7588 }),
  .A3({ S25957[520] }),
  .ZN({ S7637 })
);
AOI21_X1 #() 
AOI21_X1_183_ (
  .A({ S9 }),
  .B1({ S25957[522] }),
  .B2({ S7576 }),
  .ZN({ S7638 })
);
NAND2_X1 #() 
NAND2_X1_344_ (
  .A1({ S7638 }),
  .A2({ S7637 }),
  .ZN({ S7639 })
);
OAI21_X1 #() 
OAI21_X1_201_ (
  .A({ S7639 }),
  .B1({ S7635 }),
  .B2({ S7588 }),
  .ZN({ S7640 })
);
AOI21_X1 #() 
AOI21_X1_184_ (
  .A({ S9 }),
  .B1({ S7577 }),
  .B2({ S7580 }),
  .ZN({ S7641 })
);
NAND2_X1 #() 
NAND2_X1_345_ (
  .A1({ S7620 }),
  .A2({ S7567 }),
  .ZN({ S7642 })
);
AOI21_X1 #() 
AOI21_X1_185_ (
  .A({ S7641 }),
  .B1({ S7642 }),
  .B2({ S7593 }),
  .ZN({ S7643 })
);
AOI21_X1 #() 
AOI21_X1_186_ (
  .A({ S7605 }),
  .B1({ S7643 }),
  .B2({ S7575 }),
  .ZN({ S7644 })
);
OAI21_X1 #() 
OAI21_X1_202_ (
  .A({ S7644 }),
  .B1({ S7575 }),
  .B2({ S7640 }),
  .ZN({ S7645 })
);
AOI21_X1 #() 
AOI21_X1_187_ (
  .A({ S25957[523] }),
  .B1({ S7576 }),
  .B2({ S25957[521] }),
  .ZN({ S7646 })
);
NAND2_X1 #() 
NAND2_X1_346_ (
  .A1({ S7624 }),
  .A2({ S25957[523] }),
  .ZN({ S7648 })
);
NOR2_X1 #() 
NOR2_X1_74_ (
  .A1({ S7648 }),
  .A2({ S16 }),
  .ZN({ S7649 })
);
OAI21_X1 #() 
OAI21_X1_203_ (
  .A({ S25957[524] }),
  .B1({ S7649 }),
  .B2({ S7646 }),
  .ZN({ S7650 })
);
NAND3_X1 #() 
NAND3_X1_407_ (
  .A1({ S7572 }),
  .A2({ S7588 }),
  .A3({ S7576 }),
  .ZN({ S7651 })
);
NAND2_X1 #() 
NAND2_X1_347_ (
  .A1({ S17 }),
  .A2({ S25957[522] }),
  .ZN({ S7652 })
);
NOR2_X1 #() 
NOR2_X1_75_ (
  .A1({ S25957[521] }),
  .A2({ S9 }),
  .ZN({ S7653 })
);
AOI21_X1 #() 
AOI21_X1_188_ (
  .A({ S25957[524] }),
  .B1({ S7653 }),
  .B2({ S25957[520] }),
  .ZN({ S7654 })
);
NAND3_X1 #() 
NAND3_X1_408_ (
  .A1({ S7654 }),
  .A2({ S7651 }),
  .A3({ S7652 }),
  .ZN({ S7655 })
);
AND2_X1 #() 
AND2_X1_20_ (
  .A1({ S7650 }),
  .A2({ S7655 }),
  .ZN({ S7656 })
);
OAI21_X1 #() 
OAI21_X1_204_ (
  .A({ S7645 }),
  .B1({ S7656 }),
  .B2({ S25957[525] }),
  .ZN({ S7657 })
);
NAND2_X1 #() 
NAND2_X1_348_ (
  .A1({ S7657 }),
  .A2({ S25957[526] }),
  .ZN({ S7659 })
);
INV_X1 #() 
INV_X1_142_ (
  .A({ S25957[526] }),
  .ZN({ S7660 })
);
NAND2_X1 #() 
NAND2_X1_349_ (
  .A1({ S25957[521] }),
  .A2({ S9 }),
  .ZN({ S7661 })
);
INV_X1 #() 
INV_X1_143_ (
  .A({ S7661 }),
  .ZN({ S7662 })
);
AOI21_X1 #() 
AOI21_X1_189_ (
  .A({ S9 }),
  .B1({ S6177 }),
  .B2({ S6180 }),
  .ZN({ S7663 })
);
AOI21_X1 #() 
AOI21_X1_190_ (
  .A({ S7653 }),
  .B1({ S7663 }),
  .B2({ S25957[520] }),
  .ZN({ S7664 })
);
NAND2_X1 #() 
NAND2_X1_350_ (
  .A1({ S7664 }),
  .A2({ S25957[524] }),
  .ZN({ S7665 })
);
AOI21_X1 #() 
AOI21_X1_191_ (
  .A({ S7665 }),
  .B1({ S7662 }),
  .B2({ S7606 }),
  .ZN({ S7666 })
);
OAI21_X1 #() 
OAI21_X1_205_ (
  .A({ S9 }),
  .B1({ S17 }),
  .B2({ S25957[522] }),
  .ZN({ S7667 })
);
NAND3_X1 #() 
NAND3_X1_409_ (
  .A1({ S7667 }),
  .A2({ S7575 }),
  .A3({ S7567 }),
  .ZN({ S7668 })
);
INV_X1 #() 
INV_X1_144_ (
  .A({ S7668 }),
  .ZN({ S7670 })
);
OAI21_X1 #() 
OAI21_X1_206_ (
  .A({ S25957[525] }),
  .B1({ S7666 }),
  .B2({ S7670 }),
  .ZN({ S7671 })
);
AOI21_X1 #() 
AOI21_X1_192_ (
  .A({ S9 }),
  .B1({ S7613 }),
  .B2({ S7568 }),
  .ZN({ S7672 })
);
INV_X1 #() 
INV_X1_145_ (
  .A({ S7672 }),
  .ZN({ S7673 })
);
NAND4_X1 #() 
NAND4_X1_43_ (
  .A1({ S6177 }),
  .A2({ S6180 }),
  .A3({ S7563 }),
  .A4({ S7564 }),
  .ZN({ S7674 })
);
NAND3_X1 #() 
NAND3_X1_410_ (
  .A1({ S25957[521] }),
  .A2({ S7569 }),
  .A3({ S7571 }),
  .ZN({ S7675 })
);
NAND3_X1 #() 
NAND3_X1_411_ (
  .A1({ S7674 }),
  .A2({ S7675 }),
  .A3({ S9 }),
  .ZN({ S7676 })
);
AOI21_X1 #() 
AOI21_X1_193_ (
  .A({ S7575 }),
  .B1({ S7673 }),
  .B2({ S7676 }),
  .ZN({ S7677 })
);
AOI21_X1 #() 
AOI21_X1_194_ (
  .A({ S25957[523] }),
  .B1({ S25957[522] }),
  .B2({ S7576 }),
  .ZN({ S7678 })
);
NAND2_X1 #() 
NAND2_X1_351_ (
  .A1({ S7674 }),
  .A2({ S25957[521] }),
  .ZN({ S7679 })
);
NAND3_X1 #() 
NAND3_X1_412_ (
  .A1({ S7679 }),
  .A2({ S7678 }),
  .A3({ S7637 }),
  .ZN({ S7681 })
);
AOI21_X1 #() 
AOI21_X1_195_ (
  .A({ S25957[524] }),
  .B1({ S7653 }),
  .B2({ S7572 }),
  .ZN({ S7682 })
);
NAND2_X1 #() 
NAND2_X1_352_ (
  .A1({ S7681 }),
  .A2({ S7682 }),
  .ZN({ S7683 })
);
NAND2_X1 #() 
NAND2_X1_353_ (
  .A1({ S7683 }),
  .A2({ S7605 }),
  .ZN({ S7684 })
);
OAI211_X1 #() 
OAI211_X1_106_ (
  .A({ S7671 }),
  .B({ S7660 }),
  .C1({ S7677 }),
  .C2({ S7684 }),
  .ZN({ S7685 })
);
NAND2_X1 #() 
NAND2_X1_354_ (
  .A1({ S7659 }),
  .A2({ S7685 }),
  .ZN({ S7686 })
);
NAND2_X1 #() 
NAND2_X1_355_ (
  .A1({ S7686 }),
  .A2({ S25957[527] }),
  .ZN({ S7687 })
);
NAND3_X1 #() 
NAND3_X1_413_ (
  .A1({ S7687 }),
  .A2({ S4920 }),
  .A3({ S7633 }),
  .ZN({ S7688 })
);
NAND3_X1 #() 
NAND3_X1_414_ (
  .A1({ S7659 }),
  .A2({ S25957[527] }),
  .A3({ S7685 }),
  .ZN({ S7689 })
);
OAI21_X1 #() 
OAI21_X1_207_ (
  .A({ S7632 }),
  .B1({ S25957[526] }),
  .B2({ S7604 }),
  .ZN({ S7690 })
);
NAND2_X1 #() 
NAND2_X1_356_ (
  .A1({ S7690 }),
  .A2({ S7562 }),
  .ZN({ S7692 })
);
NAND3_X1 #() 
NAND3_X1_415_ (
  .A1({ S7692 }),
  .A2({ S7689 }),
  .A3({ S25957[631] }),
  .ZN({ S7693 })
);
NAND3_X1 #() 
NAND3_X1_416_ (
  .A1({ S7688 }),
  .A2({ S7693 }),
  .A3({ S7561 }),
  .ZN({ S7694 })
);
NAND3_X1 #() 
NAND3_X1_417_ (
  .A1({ S7687 }),
  .A2({ S25957[631] }),
  .A3({ S7633 }),
  .ZN({ S7695 })
);
NAND3_X1 #() 
NAND3_X1_418_ (
  .A1({ S7692 }),
  .A2({ S7689 }),
  .A3({ S4920 }),
  .ZN({ S7696 })
);
NAND3_X1 #() 
NAND3_X1_419_ (
  .A1({ S7695 }),
  .A2({ S7696 }),
  .A3({ S25957[599] }),
  .ZN({ S7697 })
);
NAND3_X1 #() 
NAND3_X1_420_ (
  .A1({ S7694 }),
  .A2({ S7697 }),
  .A3({ S7559 }),
  .ZN({ S7698 })
);
AOI21_X1 #() 
AOI21_X1_196_ (
  .A({ S25957[599] }),
  .B1({ S7695 }),
  .B2({ S7696 }),
  .ZN({ S7699 })
);
AOI21_X1 #() 
AOI21_X1_197_ (
  .A({ S7561 }),
  .B1({ S7688 }),
  .B2({ S7693 }),
  .ZN({ S7700 })
);
OAI21_X1 #() 
OAI21_X1_208_ (
  .A({ S25957[567] }),
  .B1({ S7699 }),
  .B2({ S7700 }),
  .ZN({ S7701 })
);
NAND3_X1 #() 
NAND3_X1_421_ (
  .A1({ S7701 }),
  .A2({ S4924 }),
  .A3({ S7698 }),
  .ZN({ S7703 })
);
OAI21_X1 #() 
OAI21_X1_209_ (
  .A({ S7559 }),
  .B1({ S7699 }),
  .B2({ S7700 }),
  .ZN({ S7704 })
);
NAND3_X1 #() 
NAND3_X1_422_ (
  .A1({ S7694 }),
  .A2({ S7697 }),
  .A3({ S25957[567] }),
  .ZN({ S7705 })
);
NAND3_X1 #() 
NAND3_X1_423_ (
  .A1({ S7704 }),
  .A2({ S25957[535] }),
  .A3({ S7705 }),
  .ZN({ S7706 })
);
NAND2_X1 #() 
NAND2_X1_357_ (
  .A1({ S7703 }),
  .A2({ S7706 }),
  .ZN({ S7707 })
);
INV_X1 #() 
INV_X1_146_ (
  .A({ S7707 }),
  .ZN({ S25957[407] })
);
INV_X1 #() 
INV_X1_147_ (
  .A({ S25957[534] }),
  .ZN({ S7708 })
);
XNOR2_X1 #() 
XNOR2_X1_11_ (
  .A({ S2439 }),
  .B({ S25957[854] }),
  .ZN({ S25957[726] })
);
INV_X1 #() 
INV_X1_148_ (
  .A({ S25957[726] }),
  .ZN({ S7709 })
);
INV_X1 #() 
INV_X1_149_ (
  .A({ S7652 }),
  .ZN({ S7710 })
);
INV_X1 #() 
INV_X1_150_ (
  .A({ S7653 }),
  .ZN({ S7711 })
);
NAND2_X1 #() 
NAND2_X1_358_ (
  .A1({ S7674 }),
  .A2({ S7620 }),
  .ZN({ S7712 })
);
NOR2_X1 #() 
NOR2_X1_76_ (
  .A1({ S7712 }),
  .A2({ S7711 }),
  .ZN({ S7713 })
);
AOI21_X1 #() 
AOI21_X1_198_ (
  .A({ S7713 }),
  .B1({ S7710 }),
  .B2({ S9 }),
  .ZN({ S7714 })
);
NAND2_X1 #() 
NAND2_X1_359_ (
  .A1({ S7575 }),
  .A2({ S7661 }),
  .ZN({ S7715 })
);
OAI22_X1 #() 
OAI22_X1_10_ (
  .A1({ S7714 }),
  .A2({ S7575 }),
  .B1({ S7649 }),
  .B2({ S7715 }),
  .ZN({ S7716 })
);
NAND2_X1 #() 
NAND2_X1_360_ (
  .A1({ S7716 }),
  .A2({ S25957[526] }),
  .ZN({ S7717 })
);
NAND2_X1 #() 
NAND2_X1_361_ (
  .A1({ S7579 }),
  .A2({ S7572 }),
  .ZN({ S7718 })
);
NAND2_X1 #() 
NAND2_X1_362_ (
  .A1({ S7718 }),
  .A2({ S7675 }),
  .ZN({ S7719 })
);
INV_X1 #() 
INV_X1_151_ (
  .A({ S7719 }),
  .ZN({ S7720 })
);
NAND2_X1 #() 
NAND2_X1_363_ (
  .A1({ S7567 }),
  .A2({ S17 }),
  .ZN({ S7721 })
);
NAND3_X1 #() 
NAND3_X1_424_ (
  .A1({ S7721 }),
  .A2({ S9 }),
  .A3({ S7674 }),
  .ZN({ S7722 })
);
OAI21_X1 #() 
OAI21_X1_210_ (
  .A({ S7722 }),
  .B1({ S7720 }),
  .B2({ S9 }),
  .ZN({ S7723 })
);
NOR2_X1 #() 
NOR2_X1_77_ (
  .A1({ S25957[522] }),
  .A2({ S25957[520] }),
  .ZN({ S7724 })
);
NAND2_X1 #() 
NAND2_X1_364_ (
  .A1({ S7724 }),
  .A2({ S7662 }),
  .ZN({ S7725 })
);
AND4_X1 #() 
AND4_X1_1_ (
  .A1({ S25957[524] }),
  .A2({ S7725 }),
  .A3({ S7582 }),
  .A4({ S7618 }),
  .ZN({ S7726 })
);
AOI21_X1 #() 
AOI21_X1_199_ (
  .A({ S7726 }),
  .B1({ S7723 }),
  .B2({ S7575 }),
  .ZN({ S7727 })
);
OAI21_X1 #() 
OAI21_X1_211_ (
  .A({ S7717 }),
  .B1({ S7727 }),
  .B2({ S25957[526] }),
  .ZN({ S7728 })
);
NAND2_X1 #() 
NAND2_X1_365_ (
  .A1({ S7728 }),
  .A2({ S25957[525] }),
  .ZN({ S7729 })
);
NAND3_X1 #() 
NAND3_X1_425_ (
  .A1({ S7674 }),
  .A2({ S7620 }),
  .A3({ S7567 }),
  .ZN({ S7730 })
);
NAND2_X1 #() 
NAND2_X1_366_ (
  .A1({ S7730 }),
  .A2({ S25957[523] }),
  .ZN({ S7731 })
);
NAND2_X1 #() 
NAND2_X1_367_ (
  .A1({ S7613 }),
  .A2({ S7678 }),
  .ZN({ S7732 })
);
NAND3_X1 #() 
NAND3_X1_426_ (
  .A1({ S7731 }),
  .A2({ S25957[524] }),
  .A3({ S7732 }),
  .ZN({ S7733 })
);
AOI21_X1 #() 
AOI21_X1_200_ (
  .A({ S9 }),
  .B1({ S7652 }),
  .B2({ S7567 }),
  .ZN({ S7734 })
);
OAI21_X1 #() 
OAI21_X1_212_ (
  .A({ S7733 }),
  .B1({ S7608 }),
  .B2({ S7734 }),
  .ZN({ S7735 })
);
NAND2_X1 #() 
NAND2_X1_368_ (
  .A1({ S7579 }),
  .A2({ S25957[522] }),
  .ZN({ S7736 })
);
NAND3_X1 #() 
NAND3_X1_427_ (
  .A1({ S7736 }),
  .A2({ S25957[523] }),
  .A3({ S7610 }),
  .ZN({ S7737 })
);
AOI21_X1 #() 
AOI21_X1_201_ (
  .A({ S25957[524] }),
  .B1({ S7732 }),
  .B2({ S7737 }),
  .ZN({ S7738 })
);
INV_X1 #() 
INV_X1_152_ (
  .A({ S7626 }),
  .ZN({ S7739 })
);
AOI21_X1 #() 
AOI21_X1_202_ (
  .A({ S7665 }),
  .B1({ S9 }),
  .B2({ S7739 }),
  .ZN({ S7740 })
);
NOR3_X1 #() 
NOR3_X1_13_ (
  .A1({ S7740 }),
  .A2({ S7738 }),
  .A3({ S25957[526] }),
  .ZN({ S7742 })
);
AOI21_X1 #() 
AOI21_X1_203_ (
  .A({ S7742 }),
  .B1({ S7735 }),
  .B2({ S25957[526] }),
  .ZN({ S7743 })
);
OAI211_X1 #() 
OAI211_X1_107_ (
  .A({ S7729 }),
  .B({ S25957[527] }),
  .C1({ S25957[525] }),
  .C2({ S7743 }),
  .ZN({ S7744 })
);
AOI22_X1 #() 
AOI22_X1_30_ (
  .A1({ S7569 }),
  .A2({ S7571 }),
  .B1({ S6099 }),
  .B2({ S6096 }),
  .ZN({ S7745 })
);
AOI21_X1 #() 
AOI21_X1_204_ (
  .A({ S7575 }),
  .B1({ S7745 }),
  .B2({ S25957[523] }),
  .ZN({ S7746 })
);
INV_X1 #() 
INV_X1_153_ (
  .A({ S7746 }),
  .ZN({ S7747 })
);
AOI21_X1 #() 
AOI21_X1_205_ (
  .A({ S9 }),
  .B1({ S7718 }),
  .B2({ S7577 }),
  .ZN({ S7748 })
);
INV_X1 #() 
INV_X1_154_ (
  .A({ S7674 }),
  .ZN({ S7749 })
);
OAI22_X1 #() 
OAI22_X1_11_ (
  .A1({ S7711 }),
  .A2({ S7749 }),
  .B1({ S7637 }),
  .B2({ S25957[523] }),
  .ZN({ S7750 })
);
OAI22_X1 #() 
OAI22_X1_12_ (
  .A1({ S7747 }),
  .A2({ S7750 }),
  .B1({ S7748 }),
  .B2({ S25957[524] }),
  .ZN({ S7751 })
);
NAND2_X1 #() 
NAND2_X1_369_ (
  .A1({ S7593 }),
  .A2({ S7637 }),
  .ZN({ S7752 })
);
OAI211_X1 #() 
OAI211_X1_108_ (
  .A({ S7752 }),
  .B({ S7575 }),
  .C1({ S7745 }),
  .C2({ S7648 }),
  .ZN({ S7753 })
);
NAND3_X1 #() 
NAND3_X1_428_ (
  .A1({ S25957[522] }),
  .A2({ S7588 }),
  .A3({ S7576 }),
  .ZN({ S7754 })
);
NAND3_X1 #() 
NAND3_X1_429_ (
  .A1({ S7754 }),
  .A2({ S25957[523] }),
  .A3({ S7567 }),
  .ZN({ S7755 })
);
AOI21_X1 #() 
AOI21_X1_206_ (
  .A({ S7575 }),
  .B1({ S9 }),
  .B2({ S7674 }),
  .ZN({ S7756 })
);
AOI21_X1 #() 
AOI21_X1_207_ (
  .A({ S7605 }),
  .B1({ S7755 }),
  .B2({ S7756 }),
  .ZN({ S7757 })
);
NAND2_X1 #() 
NAND2_X1_370_ (
  .A1({ S7753 }),
  .A2({ S7757 }),
  .ZN({ S7758 })
);
OAI21_X1 #() 
OAI21_X1_213_ (
  .A({ S7758 }),
  .B1({ S7751 }),
  .B2({ S25957[525] }),
  .ZN({ S7759 })
);
NAND2_X1 #() 
NAND2_X1_371_ (
  .A1({ S7606 }),
  .A2({ S7579 }),
  .ZN({ S7760 })
);
OAI211_X1 #() 
OAI211_X1_109_ (
  .A({ S7674 }),
  .B({ S9 }),
  .C1({ S16 }),
  .C2({ S7572 }),
  .ZN({ S7761 })
);
NAND2_X1 #() 
NAND2_X1_372_ (
  .A1({ S7761 }),
  .A2({ S25957[524] }),
  .ZN({ S7763 })
);
AOI21_X1 #() 
AOI21_X1_208_ (
  .A({ S7763 }),
  .B1({ S7760 }),
  .B2({ S25957[523] }),
  .ZN({ S7764 })
);
INV_X1 #() 
INV_X1_155_ (
  .A({ S7760 }),
  .ZN({ S7765 })
);
AOI211_X1 #() 
AOI211_X1_4_ (
  .A({ S25957[524] }),
  .B({ S7765 }),
  .C1({ S9 }),
  .C2({ S7588 }),
  .ZN({ S7766 })
);
OAI21_X1 #() 
OAI21_X1_214_ (
  .A({ S25957[525] }),
  .B1({ S7766 }),
  .B2({ S7764 }),
  .ZN({ S7767 })
);
INV_X1 #() 
INV_X1_156_ (
  .A({ S7568 }),
  .ZN({ S7768 })
);
OAI211_X1 #() 
OAI211_X1_110_ (
  .A({ S7731 }),
  .B({ S7575 }),
  .C1({ S25957[523] }),
  .C2({ S7768 }),
  .ZN({ S7769 })
);
NAND2_X1 #() 
NAND2_X1_373_ (
  .A1({ S7596 }),
  .A2({ S7576 }),
  .ZN({ S7770 })
);
OAI21_X1 #() 
OAI21_X1_215_ (
  .A({ S7746 }),
  .B1({ S25957[523] }),
  .B2({ S7770 }),
  .ZN({ S7771 })
);
NAND3_X1 #() 
NAND3_X1_430_ (
  .A1({ S7769 }),
  .A2({ S7605 }),
  .A3({ S7771 }),
  .ZN({ S7772 })
);
NAND3_X1 #() 
NAND3_X1_431_ (
  .A1({ S7767 }),
  .A2({ S25957[526] }),
  .A3({ S7772 }),
  .ZN({ S7774 })
);
OAI211_X1 #() 
OAI211_X1_111_ (
  .A({ S7774 }),
  .B({ S7562 }),
  .C1({ S25957[526] }),
  .C2({ S7759 }),
  .ZN({ S7775 })
);
NAND3_X1 #() 
NAND3_X1_432_ (
  .A1({ S7744 }),
  .A2({ S7775 }),
  .A3({ S7709 }),
  .ZN({ S7776 })
);
NAND2_X1 #() 
NAND2_X1_374_ (
  .A1({ S7744 }),
  .A2({ S7775 }),
  .ZN({ S7777 })
);
NAND2_X1 #() 
NAND2_X1_375_ (
  .A1({ S7777 }),
  .A2({ S25957[726] }),
  .ZN({ S7778 })
);
NAND2_X1 #() 
NAND2_X1_376_ (
  .A1({ S7778 }),
  .A2({ S7776 }),
  .ZN({ S25957[470] })
);
OAI21_X1 #() 
OAI21_X1_216_ (
  .A({ S25957[470] }),
  .B1({ S4991 }),
  .B2({ S4992 }),
  .ZN({ S7779 })
);
NAND3_X1 #() 
NAND3_X1_433_ (
  .A1({ S7778 }),
  .A2({ S25957[566] }),
  .A3({ S7776 }),
  .ZN({ S7780 })
);
NAND3_X1 #() 
NAND3_X1_434_ (
  .A1({ S7779 }),
  .A2({ S7708 }),
  .A3({ S7780 }),
  .ZN({ S7781 })
);
NAND2_X1 #() 
NAND2_X1_377_ (
  .A1({ S7779 }),
  .A2({ S7780 }),
  .ZN({ S25957[438] })
);
NAND2_X1 #() 
NAND2_X1_378_ (
  .A1({ S25957[438] }),
  .A2({ S25957[534] }),
  .ZN({ S7783 })
);
NAND2_X1 #() 
NAND2_X1_379_ (
  .A1({ S7783 }),
  .A2({ S7781 }),
  .ZN({ S7784 })
);
INV_X1 #() 
INV_X1_157_ (
  .A({ S7784 }),
  .ZN({ S25957[406] })
);
NOR2_X1 #() 
NOR2_X1_78_ (
  .A1({ S5056 }),
  .A2({ S5057 }),
  .ZN({ S25957[597] })
);
NAND2_X1 #() 
NAND2_X1_380_ (
  .A1({ S2516 }),
  .A2({ S2517 }),
  .ZN({ S25957[757] })
);
XOR2_X1 #() 
XOR2_X1_7_ (
  .A({ S5060 }),
  .B({ S25957[757] }),
  .Z({ S25957[629] })
);
OAI221_X1 #() 
OAI221_X1_5_ (
  .A({ S7575 }),
  .B1({ S7606 }),
  .B2({ S9 }),
  .C1({ S7712 }),
  .C2({ S7661 }),
  .ZN({ S7785 })
);
NOR2_X1 #() 
NOR2_X1_79_ (
  .A1({ S16 }),
  .A2({ S25957[522] }),
  .ZN({ S7786 })
);
OAI21_X1 #() 
OAI21_X1_217_ (
  .A({ S7725 }),
  .B1({ S7786 }),
  .B2({ S9 }),
  .ZN({ S7787 })
);
AOI21_X1 #() 
AOI21_X1_209_ (
  .A({ S7605 }),
  .B1({ S7787 }),
  .B2({ S25957[524] }),
  .ZN({ S7788 })
);
AND2_X1 #() 
AND2_X1_21_ (
  .A1({ S7788 }),
  .A2({ S7785 }),
  .ZN({ S7790 })
);
NAND3_X1 #() 
NAND3_X1_435_ (
  .A1({ S7611 }),
  .A2({ S25957[523] }),
  .A3({ S7637 }),
  .ZN({ S7791 })
);
AOI21_X1 #() 
AOI21_X1_210_ (
  .A({ S25957[523] }),
  .B1({ S7754 }),
  .B2({ S7567 }),
  .ZN({ S7792 })
);
INV_X1 #() 
INV_X1_158_ (
  .A({ S7792 }),
  .ZN({ S7793 })
);
NAND3_X1 #() 
NAND3_X1_436_ (
  .A1({ S7793 }),
  .A2({ S25957[524] }),
  .A3({ S7791 }),
  .ZN({ S7794 })
);
INV_X1 #() 
INV_X1_159_ (
  .A({ S7589 }),
  .ZN({ S7795 })
);
NOR2_X1 #() 
NOR2_X1_80_ (
  .A1({ S7567 }),
  .A2({ S7572 }),
  .ZN({ S7796 })
);
OAI211_X1 #() 
OAI211_X1_112_ (
  .A({ S7575 }),
  .B({ S7795 }),
  .C1({ S7796 }),
  .C2({ S25957[523] }),
  .ZN({ S7797 })
);
AOI21_X1 #() 
AOI21_X1_211_ (
  .A({ S25957[525] }),
  .B1({ S7794 }),
  .B2({ S7797 }),
  .ZN({ S7798 })
);
OAI21_X1 #() 
OAI21_X1_218_ (
  .A({ S7660 }),
  .B1({ S7790 }),
  .B2({ S7798 }),
  .ZN({ S7799 })
);
AOI22_X1 #() 
AOI22_X1_31_ (
  .A1({ S7563 }),
  .A2({ S7564 }),
  .B1({ S6099 }),
  .B2({ S6096 }),
  .ZN({ S7801 })
);
NAND2_X1 #() 
NAND2_X1_381_ (
  .A1({ S7801 }),
  .A2({ S7572 }),
  .ZN({ S7802 })
);
AND3_X1 #() 
AND3_X1_15_ (
  .A1({ S7611 }),
  .A2({ S7802 }),
  .A3({ S25957[523] }),
  .ZN({ S7803 })
);
NOR2_X1 #() 
NOR2_X1_81_ (
  .A1({ S25957[520] }),
  .A2({ S9 }),
  .ZN({ S7804 })
);
NAND2_X1 #() 
NAND2_X1_382_ (
  .A1({ S7579 }),
  .A2({ S9 }),
  .ZN({ S7805 })
);
NOR2_X1 #() 
NOR2_X1_82_ (
  .A1({ S7805 }),
  .A2({ S7749 }),
  .ZN({ S7806 })
);
OAI21_X1 #() 
OAI21_X1_219_ (
  .A({ S7575 }),
  .B1({ S7806 }),
  .B2({ S7804 }),
  .ZN({ S7807 })
);
NAND2_X1 #() 
NAND2_X1_383_ (
  .A1({ S7624 }),
  .A2({ S17 }),
  .ZN({ S7808 })
);
NAND2_X1 #() 
NAND2_X1_384_ (
  .A1({ S7587 }),
  .A2({ S9 }),
  .ZN({ S7809 })
);
OAI21_X1 #() 
OAI21_X1_220_ (
  .A({ S25957[524] }),
  .B1({ S7808 }),
  .B2({ S7809 }),
  .ZN({ S7810 })
);
OAI211_X1 #() 
OAI211_X1_113_ (
  .A({ S7807 }),
  .B({ S25957[525] }),
  .C1({ S7803 }),
  .C2({ S7810 }),
  .ZN({ S7812 })
);
NAND2_X1 #() 
NAND2_X1_385_ (
  .A1({ S7739 }),
  .A2({ S25957[523] }),
  .ZN({ S7813 })
);
NAND2_X1 #() 
NAND2_X1_386_ (
  .A1({ S16 }),
  .A2({ S25957[522] }),
  .ZN({ S7814 })
);
NAND3_X1 #() 
NAND3_X1_437_ (
  .A1({ S7591 }),
  .A2({ S7814 }),
  .A3({ S9 }),
  .ZN({ S7815 })
);
NAND3_X1 #() 
NAND3_X1_438_ (
  .A1({ S7813 }),
  .A2({ S7815 }),
  .A3({ S25957[524] }),
  .ZN({ S7816 })
);
NAND3_X1 #() 
NAND3_X1_439_ (
  .A1({ S7583 }),
  .A2({ S25957[523] }),
  .A3({ S7674 }),
  .ZN({ S7817 })
);
NAND3_X1 #() 
NAND3_X1_440_ (
  .A1({ S7802 }),
  .A2({ S9 }),
  .A3({ S7606 }),
  .ZN({ S7818 })
);
AND2_X1 #() 
AND2_X1_22_ (
  .A1({ S7817 }),
  .A2({ S7818 }),
  .ZN({ S7819 })
);
OAI211_X1 #() 
OAI211_X1_114_ (
  .A({ S7605 }),
  .B({ S7816 }),
  .C1({ S7819 }),
  .C2({ S25957[524] }),
  .ZN({ S7820 })
);
NAND3_X1 #() 
NAND3_X1_441_ (
  .A1({ S7820 }),
  .A2({ S7812 }),
  .A3({ S25957[526] }),
  .ZN({ S7821 })
);
NAND3_X1 #() 
NAND3_X1_442_ (
  .A1({ S7799 }),
  .A2({ S7562 }),
  .A3({ S7821 }),
  .ZN({ S7823 })
);
NAND3_X1 #() 
NAND3_X1_443_ (
  .A1({ S7626 }),
  .A2({ S7577 }),
  .A3({ S9 }),
  .ZN({ S7824 })
);
OAI211_X1 #() 
OAI211_X1_115_ (
  .A({ S7824 }),
  .B({ S25957[524] }),
  .C1({ S9 }),
  .C2({ S7770 }),
  .ZN({ S7825 })
);
AOI21_X1 #() 
AOI21_X1_212_ (
  .A({ S7588 }),
  .B1({ S7674 }),
  .B2({ S7620 }),
  .ZN({ S7826 })
);
NAND2_X1 #() 
NAND2_X1_387_ (
  .A1({ S7606 }),
  .A2({ S7588 }),
  .ZN({ S7827 })
);
NAND2_X1 #() 
NAND2_X1_388_ (
  .A1({ S7827 }),
  .A2({ S9 }),
  .ZN({ S7828 })
);
OAI21_X1 #() 
OAI21_X1_221_ (
  .A({ S7828 }),
  .B1({ S7826 }),
  .B2({ S9 }),
  .ZN({ S7829 })
);
NAND2_X1 #() 
NAND2_X1_389_ (
  .A1({ S7829 }),
  .A2({ S7575 }),
  .ZN({ S7830 })
);
NAND2_X1 #() 
NAND2_X1_390_ (
  .A1({ S7830 }),
  .A2({ S7825 }),
  .ZN({ S7831 })
);
NAND2_X1 #() 
NAND2_X1_391_ (
  .A1({ S7831 }),
  .A2({ S25957[525] }),
  .ZN({ S7832 })
);
NAND3_X1 #() 
NAND3_X1_444_ (
  .A1({ S7731 }),
  .A2({ S7575 }),
  .A3({ S7582 }),
  .ZN({ S7834 })
);
OAI21_X1 #() 
OAI21_X1_222_ (
  .A({ S25957[523] }),
  .B1({ S7801 }),
  .B2({ S25957[522] }),
  .ZN({ S7835 })
);
NAND2_X1 #() 
NAND2_X1_392_ (
  .A1({ S7646 }),
  .A2({ S25957[522] }),
  .ZN({ S7836 })
);
NAND2_X1 #() 
NAND2_X1_393_ (
  .A1({ S7836 }),
  .A2({ S7835 }),
  .ZN({ S7837 })
);
OAI211_X1 #() 
OAI211_X1_116_ (
  .A({ S7834 }),
  .B({ S7605 }),
  .C1({ S7575 }),
  .C2({ S7837 }),
  .ZN({ S7838 })
);
AOI21_X1 #() 
AOI21_X1_213_ (
  .A({ S7660 }),
  .B1({ S7832 }),
  .B2({ S7838 }),
  .ZN({ S7839 })
);
INV_X1 #() 
INV_X1_160_ (
  .A({ S7839 }),
  .ZN({ S7840 })
);
AOI21_X1 #() 
AOI21_X1_214_ (
  .A({ S7653 }),
  .B1({ S7646 }),
  .B2({ S7596 }),
  .ZN({ S7841 })
);
NOR2_X1 #() 
NOR2_X1_83_ (
  .A1({ S7661 }),
  .A2({ S7576 }),
  .ZN({ S7842 })
);
NAND2_X1 #() 
NAND2_X1_394_ (
  .A1({ S7583 }),
  .A2({ S7626 }),
  .ZN({ S7843 })
);
OAI21_X1 #() 
OAI21_X1_223_ (
  .A({ S7635 }),
  .B1({ S7843 }),
  .B2({ S9 }),
  .ZN({ S7845 })
);
NAND2_X1 #() 
NAND2_X1_395_ (
  .A1({ S7845 }),
  .A2({ S25957[524] }),
  .ZN({ S7846 })
);
OAI221_X1 #() 
OAI221_X1_6_ (
  .A({ S25957[525] }),
  .B1({ S7841 }),
  .B2({ S25957[524] }),
  .C1({ S7846 }),
  .C2({ S7842 }),
  .ZN({ S7847 })
);
NAND2_X1 #() 
NAND2_X1_396_ (
  .A1({ S7568 }),
  .A2({ S7651 }),
  .ZN({ S7848 })
);
AOI21_X1 #() 
AOI21_X1_215_ (
  .A({ S7573 }),
  .B1({ S7848 }),
  .B2({ S25957[523] }),
  .ZN({ S7849 })
);
INV_X1 #() 
INV_X1_161_ (
  .A({ S17 }),
  .ZN({ S7850 })
);
NOR2_X1 #() 
NOR2_X1_84_ (
  .A1({ S7591 }),
  .A2({ S7850 }),
  .ZN({ S7851 })
);
NAND2_X1 #() 
NAND2_X1_397_ (
  .A1({ S7851 }),
  .A2({ S25957[523] }),
  .ZN({ S7852 })
);
AOI21_X1 #() 
AOI21_X1_216_ (
  .A({ S7575 }),
  .B1({ S7808 }),
  .B2({ S9 }),
  .ZN({ S7853 })
);
NAND2_X1 #() 
NAND2_X1_398_ (
  .A1({ S7852 }),
  .A2({ S7853 }),
  .ZN({ S7854 })
);
OAI211_X1 #() 
OAI211_X1_117_ (
  .A({ S7854 }),
  .B({ S7605 }),
  .C1({ S25957[524] }),
  .C2({ S7849 }),
  .ZN({ S7856 })
);
NAND3_X1 #() 
NAND3_X1_445_ (
  .A1({ S7847 }),
  .A2({ S7856 }),
  .A3({ S7660 }),
  .ZN({ S7857 })
);
NAND3_X1 #() 
NAND3_X1_446_ (
  .A1({ S7840 }),
  .A2({ S25957[527] }),
  .A3({ S7857 }),
  .ZN({ S7858 })
);
NAND3_X1 #() 
NAND3_X1_447_ (
  .A1({ S7858 }),
  .A2({ S25957[629] }),
  .A3({ S7823 }),
  .ZN({ S7859 })
);
INV_X1 #() 
INV_X1_162_ (
  .A({ S25957[629] }),
  .ZN({ S7860 })
);
INV_X1 #() 
INV_X1_163_ (
  .A({ S7857 }),
  .ZN({ S7861 })
);
OAI21_X1 #() 
OAI21_X1_224_ (
  .A({ S25957[527] }),
  .B1({ S7861 }),
  .B2({ S7839 }),
  .ZN({ S7862 })
);
NAND2_X1 #() 
NAND2_X1_399_ (
  .A1({ S7799 }),
  .A2({ S7821 }),
  .ZN({ S7863 })
);
NAND2_X1 #() 
NAND2_X1_400_ (
  .A1({ S7863 }),
  .A2({ S7562 }),
  .ZN({ S7864 })
);
NAND3_X1 #() 
NAND3_X1_448_ (
  .A1({ S7862 }),
  .A2({ S7860 }),
  .A3({ S7864 }),
  .ZN({ S7865 })
);
NAND2_X1 #() 
NAND2_X1_401_ (
  .A1({ S7865 }),
  .A2({ S7859 }),
  .ZN({ S25957[501] })
);
NAND2_X1 #() 
NAND2_X1_402_ (
  .A1({ S25957[501] }),
  .A2({ S25957[597] }),
  .ZN({ S7867 })
);
INV_X1 #() 
INV_X1_164_ (
  .A({ S25957[597] }),
  .ZN({ S7868 })
);
NAND3_X1 #() 
NAND3_X1_449_ (
  .A1({ S7865 }),
  .A2({ S7859 }),
  .A3({ S7868 }),
  .ZN({ S7869 })
);
NAND3_X1 #() 
NAND3_X1_450_ (
  .A1({ S7867 }),
  .A2({ S7869 }),
  .A3({ S4995 }),
  .ZN({ S7870 })
);
NAND3_X1 #() 
NAND3_X1_451_ (
  .A1({ S7858 }),
  .A2({ S7860 }),
  .A3({ S7823 }),
  .ZN({ S7871 })
);
NAND3_X1 #() 
NAND3_X1_452_ (
  .A1({ S7862 }),
  .A2({ S25957[629] }),
  .A3({ S7864 }),
  .ZN({ S7872 })
);
NAND3_X1 #() 
NAND3_X1_453_ (
  .A1({ S7872 }),
  .A2({ S7871 }),
  .A3({ S7868 }),
  .ZN({ S7873 })
);
NAND3_X1 #() 
NAND3_X1_454_ (
  .A1({ S7865 }),
  .A2({ S7859 }),
  .A3({ S25957[597] }),
  .ZN({ S7874 })
);
NAND3_X1 #() 
NAND3_X1_455_ (
  .A1({ S7873 }),
  .A2({ S7874 }),
  .A3({ S25957[661] }),
  .ZN({ S7875 })
);
NAND2_X1 #() 
NAND2_X1_403_ (
  .A1({ S7870 }),
  .A2({ S7875 }),
  .ZN({ S25957[405] })
);
NAND2_X1 #() 
NAND2_X1_404_ (
  .A1({ S5123 }),
  .A2({ S5121 }),
  .ZN({ S25957[596] })
);
XOR2_X1 #() 
XOR2_X1_8_ (
  .A({ S25957[596] }),
  .B({ S25957[692] }),
  .Z({ S25957[564] })
);
INV_X1 #() 
INV_X1_165_ (
  .A({ S25957[564] }),
  .ZN({ S7877 })
);
NAND2_X1 #() 
NAND2_X1_405_ (
  .A1({ S2590 }),
  .A2({ S2579 }),
  .ZN({ S25957[756] })
);
XNOR2_X1 #() 
XNOR2_X1_12_ (
  .A({ S25957[756] }),
  .B({ S5067 }),
  .ZN({ S25957[724] })
);
INV_X1 #() 
INV_X1_166_ (
  .A({ S25957[724] }),
  .ZN({ S7878 })
);
NAND2_X1 #() 
NAND2_X1_406_ (
  .A1({ S7754 }),
  .A2({ S9 }),
  .ZN({ S7879 })
);
NAND3_X1 #() 
NAND3_X1_456_ (
  .A1({ S7813 }),
  .A2({ S25957[524] }),
  .A3({ S7879 }),
  .ZN({ S7880 })
);
NAND3_X1 #() 
NAND3_X1_457_ (
  .A1({ S7587 }),
  .A2({ S9 }),
  .A3({ S7576 }),
  .ZN({ S7881 })
);
NAND3_X1 #() 
NAND3_X1_458_ (
  .A1({ S7598 }),
  .A2({ S7881 }),
  .A3({ S7575 }),
  .ZN({ S7883 })
);
NAND3_X1 #() 
NAND3_X1_459_ (
  .A1({ S7880 }),
  .A2({ S25957[525] }),
  .A3({ S7883 }),
  .ZN({ S7884 })
);
NAND2_X1 #() 
NAND2_X1_407_ (
  .A1({ S7674 }),
  .A2({ S7588 }),
  .ZN({ S7885 })
);
AOI21_X1 #() 
AOI21_X1_217_ (
  .A({ S7575 }),
  .B1({ S7646 }),
  .B2({ S7596 }),
  .ZN({ S7886 })
);
OAI21_X1 #() 
OAI21_X1_225_ (
  .A({ S7886 }),
  .B1({ S9 }),
  .B2({ S7885 }),
  .ZN({ S7887 })
);
NAND3_X1 #() 
NAND3_X1_460_ (
  .A1({ S7596 }),
  .A2({ S7620 }),
  .A3({ S9 }),
  .ZN({ S7888 })
);
AOI21_X1 #() 
AOI21_X1_218_ (
  .A({ S25957[524] }),
  .B1({ S7589 }),
  .B2({ S7587 }),
  .ZN({ S7889 })
);
NAND2_X1 #() 
NAND2_X1_408_ (
  .A1({ S7889 }),
  .A2({ S7888 }),
  .ZN({ S7890 })
);
NAND3_X1 #() 
NAND3_X1_461_ (
  .A1({ S7887 }),
  .A2({ S7890 }),
  .A3({ S7605 }),
  .ZN({ S7891 })
);
NAND2_X1 #() 
NAND2_X1_409_ (
  .A1({ S7884 }),
  .A2({ S7891 }),
  .ZN({ S7892 })
);
NAND2_X1 #() 
NAND2_X1_410_ (
  .A1({ S7892 }),
  .A2({ S25957[526] }),
  .ZN({ S7894 })
);
NAND3_X1 #() 
NAND3_X1_462_ (
  .A1({ S7802 }),
  .A2({ S25957[523] }),
  .A3({ S7580 }),
  .ZN({ S7895 })
);
INV_X1 #() 
INV_X1_167_ (
  .A({ S7596 }),
  .ZN({ S7896 })
);
OAI21_X1 #() 
OAI21_X1_226_ (
  .A({ S9 }),
  .B1({ S7642 }),
  .B2({ S7896 }),
  .ZN({ S7897 })
);
NAND3_X1 #() 
NAND3_X1_463_ (
  .A1({ S7897 }),
  .A2({ S25957[524] }),
  .A3({ S7895 }),
  .ZN({ S7898 })
);
NAND2_X1 #() 
NAND2_X1_411_ (
  .A1({ S7606 }),
  .A2({ S7653 }),
  .ZN({ S7899 })
);
AOI21_X1 #() 
AOI21_X1_219_ (
  .A({ S25957[523] }),
  .B1({ S7718 }),
  .B2({ S7577 }),
  .ZN({ S7900 })
);
NOR2_X1 #() 
NOR2_X1_85_ (
  .A1({ S7900 }),
  .A2({ S25957[524] }),
  .ZN({ S7901 })
);
NAND2_X1 #() 
NAND2_X1_412_ (
  .A1({ S7736 }),
  .A2({ S25957[523] }),
  .ZN({ S7902 })
);
NOR2_X1 #() 
NOR2_X1_86_ (
  .A1({ S7902 }),
  .A2({ S7745 }),
  .ZN({ S7903 })
);
AOI21_X1 #() 
AOI21_X1_220_ (
  .A({ S25957[523] }),
  .B1({ S7736 }),
  .B2({ S7591 }),
  .ZN({ S7905 })
);
NOR2_X1 #() 
NOR2_X1_87_ (
  .A1({ S7903 }),
  .A2({ S7905 }),
  .ZN({ S7906 })
);
AOI22_X1 #() 
AOI22_X1_32_ (
  .A1({ S7906 }),
  .A2({ S25957[524] }),
  .B1({ S7899 }),
  .B2({ S7901 }),
  .ZN({ S7907 })
);
OAI21_X1 #() 
OAI21_X1_227_ (
  .A({ S9 }),
  .B1({ S7826 }),
  .B2({ S7808 }),
  .ZN({ S7908 })
);
AOI21_X1 #() 
AOI21_X1_221_ (
  .A({ S25957[524] }),
  .B1({ S7736 }),
  .B2({ S7589 }),
  .ZN({ S7909 })
);
AOI21_X1 #() 
AOI21_X1_222_ (
  .A({ S7605 }),
  .B1({ S7908 }),
  .B2({ S7909 }),
  .ZN({ S7910 })
);
AOI22_X1 #() 
AOI22_X1_33_ (
  .A1({ S7907 }),
  .A2({ S7605 }),
  .B1({ S7910 }),
  .B2({ S7898 }),
  .ZN({ S7911 })
);
OAI21_X1 #() 
OAI21_X1_228_ (
  .A({ S7894 }),
  .B1({ S7911 }),
  .B2({ S25957[526] }),
  .ZN({ S7912 })
);
NAND2_X1 #() 
NAND2_X1_413_ (
  .A1({ S7912 }),
  .A2({ S25957[527] }),
  .ZN({ S7913 })
);
INV_X1 #() 
INV_X1_168_ (
  .A({ S140 }),
  .ZN({ S7914 })
);
OAI21_X1 #() 
OAI21_X1_229_ (
  .A({ S25957[524] }),
  .B1({ S25957[522] }),
  .B2({ S7914 }),
  .ZN({ S7916 })
);
NAND3_X1 #() 
NAND3_X1_464_ (
  .A1({ S7786 }),
  .A2({ S9 }),
  .A3({ S17 }),
  .ZN({ S7917 })
);
NAND4_X1 #() 
NAND4_X1_44_ (
  .A1({ S7917 }),
  .A2({ S7817 }),
  .A3({ S7836 }),
  .A4({ S7575 }),
  .ZN({ S7918 })
);
AOI21_X1 #() 
AOI21_X1_223_ (
  .A({ S7660 }),
  .B1({ S7918 }),
  .B2({ S7916 }),
  .ZN({ S7919 })
);
NAND2_X1 #() 
NAND2_X1_414_ (
  .A1({ S7627 }),
  .A2({ S7836 }),
  .ZN({ S7920 })
);
NAND2_X1 #() 
NAND2_X1_415_ (
  .A1({ S7920 }),
  .A2({ S25957[524] }),
  .ZN({ S7921 })
);
OAI211_X1 #() 
OAI211_X1_118_ (
  .A({ S7852 }),
  .B({ S7575 }),
  .C1({ S25957[523] }),
  .C2({ S7567 }),
  .ZN({ S7922 })
);
AOI21_X1 #() 
AOI21_X1_224_ (
  .A({ S25957[526] }),
  .B1({ S7922 }),
  .B2({ S7921 }),
  .ZN({ S7923 })
);
OAI21_X1 #() 
OAI21_X1_230_ (
  .A({ S25957[525] }),
  .B1({ S7919 }),
  .B2({ S7923 }),
  .ZN({ S7924 })
);
NAND2_X1 #() 
NAND2_X1_416_ (
  .A1({ S16 }),
  .A2({ S7572 }),
  .ZN({ S7925 })
);
NAND2_X1 #() 
NAND2_X1_417_ (
  .A1({ S7678 }),
  .A2({ S7925 }),
  .ZN({ S7927 })
);
NOR2_X1 #() 
NOR2_X1_88_ (
  .A1({ S7663 }),
  .A2({ S25957[524] }),
  .ZN({ S7928 })
);
NAND2_X1 #() 
NAND2_X1_418_ (
  .A1({ S7927 }),
  .A2({ S7928 }),
  .ZN({ S7929 })
);
NAND2_X1 #() 
NAND2_X1_419_ (
  .A1({ S7652 }),
  .A2({ S9 }),
  .ZN({ S7930 })
);
NOR2_X1 #() 
NOR2_X1_89_ (
  .A1({ S7930 }),
  .A2({ S7896 }),
  .ZN({ S7931 })
);
OAI21_X1 #() 
OAI21_X1_231_ (
  .A({ S7929 }),
  .B1({ S7931 }),
  .B2({ S7665 }),
  .ZN({ S7932 })
);
NAND3_X1 #() 
NAND3_X1_465_ (
  .A1({ S7606 }),
  .A2({ S25957[523] }),
  .A3({ S17 }),
  .ZN({ S7933 })
);
NAND2_X1 #() 
NAND2_X1_420_ (
  .A1({ S17 }),
  .A2({ S7572 }),
  .ZN({ S7934 })
);
NAND3_X1 #() 
NAND3_X1_466_ (
  .A1({ S7754 }),
  .A2({ S7934 }),
  .A3({ S9 }),
  .ZN({ S7935 })
);
NAND2_X1 #() 
NAND2_X1_421_ (
  .A1({ S7935 }),
  .A2({ S7933 }),
  .ZN({ S7936 })
);
NAND2_X1 #() 
NAND2_X1_422_ (
  .A1({ S7936 }),
  .A2({ S7575 }),
  .ZN({ S7938 })
);
NAND2_X1 #() 
NAND2_X1_423_ (
  .A1({ S7597 }),
  .A2({ S7626 }),
  .ZN({ S7939 })
);
AOI21_X1 #() 
AOI21_X1_225_ (
  .A({ S25957[526] }),
  .B1({ S7886 }),
  .B2({ S7939 }),
  .ZN({ S7940 })
);
AOI22_X1 #() 
AOI22_X1_34_ (
  .A1({ S7940 }),
  .A2({ S7938 }),
  .B1({ S7932 }),
  .B2({ S25957[526] }),
  .ZN({ S7941 })
);
OAI211_X1 #() 
OAI211_X1_119_ (
  .A({ S7924 }),
  .B({ S7562 }),
  .C1({ S7941 }),
  .C2({ S25957[525] }),
  .ZN({ S7942 })
);
NAND3_X1 #() 
NAND3_X1_467_ (
  .A1({ S7913 }),
  .A2({ S7942 }),
  .A3({ S7878 }),
  .ZN({ S7943 })
);
OAI211_X1 #() 
OAI211_X1_120_ (
  .A({ S7894 }),
  .B({ S25957[527] }),
  .C1({ S7911 }),
  .C2({ S25957[526] }),
  .ZN({ S7944 })
);
NAND3_X1 #() 
NAND3_X1_468_ (
  .A1({ S7918 }),
  .A2({ S25957[525] }),
  .A3({ S7916 }),
  .ZN({ S7945 })
);
OAI21_X1 #() 
OAI21_X1_232_ (
  .A({ S7945 }),
  .B1({ S7932 }),
  .B2({ S25957[525] }),
  .ZN({ S7946 })
);
NAND2_X1 #() 
NAND2_X1_424_ (
  .A1({ S7946 }),
  .A2({ S25957[526] }),
  .ZN({ S7947 })
);
AND2_X1 #() 
AND2_X1_23_ (
  .A1({ S7922 }),
  .A2({ S7921 }),
  .ZN({ S7949 })
);
NAND2_X1 #() 
NAND2_X1_425_ (
  .A1({ S7886 }),
  .A2({ S7939 }),
  .ZN({ S7950 })
);
NAND3_X1 #() 
NAND3_X1_469_ (
  .A1({ S7938 }),
  .A2({ S7605 }),
  .A3({ S7950 }),
  .ZN({ S7951 })
);
OAI211_X1 #() 
OAI211_X1_121_ (
  .A({ S7951 }),
  .B({ S7660 }),
  .C1({ S7949 }),
  .C2({ S7605 }),
  .ZN({ S7952 })
);
NAND3_X1 #() 
NAND3_X1_470_ (
  .A1({ S7952 }),
  .A2({ S7562 }),
  .A3({ S7947 }),
  .ZN({ S7953 })
);
NAND3_X1 #() 
NAND3_X1_471_ (
  .A1({ S7953 }),
  .A2({ S7944 }),
  .A3({ S25957[724] }),
  .ZN({ S7954 })
);
NAND3_X1 #() 
NAND3_X1_472_ (
  .A1({ S7943 }),
  .A2({ S7954 }),
  .A3({ S7877 }),
  .ZN({ S7955 })
);
AOI21_X1 #() 
AOI21_X1_226_ (
  .A({ S25957[724] }),
  .B1({ S7953 }),
  .B2({ S7944 }),
  .ZN({ S7956 })
);
INV_X1 #() 
INV_X1_169_ (
  .A({ S7954 }),
  .ZN({ S7957 })
);
OAI21_X1 #() 
OAI21_X1_233_ (
  .A({ S25957[564] }),
  .B1({ S7957 }),
  .B2({ S7956 }),
  .ZN({ S7958 })
);
NAND3_X1 #() 
NAND3_X1_473_ (
  .A1({ S7958 }),
  .A2({ S5128 }),
  .A3({ S7955 }),
  .ZN({ S7960 })
);
OAI21_X1 #() 
OAI21_X1_234_ (
  .A({ S7877 }),
  .B1({ S7957 }),
  .B2({ S7956 }),
  .ZN({ S7961 })
);
NAND3_X1 #() 
NAND3_X1_474_ (
  .A1({ S7943 }),
  .A2({ S7954 }),
  .A3({ S25957[564] }),
  .ZN({ S7962 })
);
NAND3_X1 #() 
NAND3_X1_475_ (
  .A1({ S7961 }),
  .A2({ S25957[532] }),
  .A3({ S7962 }),
  .ZN({ S7963 })
);
NAND2_X1 #() 
NAND2_X1_426_ (
  .A1({ S7960 }),
  .A2({ S7963 }),
  .ZN({ S25957[404] })
);
NAND2_X1 #() 
NAND2_X1_427_ (
  .A1({ S5219 }),
  .A2({ S5216 }),
  .ZN({ S25957[563] })
);
INV_X1 #() 
INV_X1_170_ (
  .A({ S25957[563] }),
  .ZN({ S7964 })
);
NOR2_X1 #() 
NOR2_X1_90_ (
  .A1({ S5218 }),
  .A2({ S5217 }),
  .ZN({ S7965 })
);
INV_X1 #() 
INV_X1_171_ (
  .A({ S7965 }),
  .ZN({ S25957[595] })
);
NAND2_X1 #() 
NAND2_X1_428_ (
  .A1({ S23083 }),
  .A2({ S23084 }),
  .ZN({ S25957[1011] })
);
NAND2_X1 #() 
NAND2_X1_429_ (
  .A1({ S25810 }),
  .A2({ S25824 }),
  .ZN({ S7967 })
);
XNOR2_X1 #() 
XNOR2_X1_13_ (
  .A({ S7967 }),
  .B({ S25957[1011] }),
  .ZN({ S25957[883] })
);
NAND2_X1 #() 
NAND2_X1_430_ (
  .A1({ S2650 }),
  .A2({ S2655 }),
  .ZN({ S7968 })
);
XNOR2_X1 #() 
XNOR2_X1_14_ (
  .A({ S7968 }),
  .B({ S25957[883] }),
  .ZN({ S25957[755] })
);
NAND2_X1 #() 
NAND2_X1_431_ (
  .A1({ S5214 }),
  .A2({ S5203 }),
  .ZN({ S7969 })
);
XOR2_X1 #() 
XOR2_X1_9_ (
  .A({ S7969 }),
  .B({ S25957[755] }),
  .Z({ S25957[627] })
);
INV_X1 #() 
INV_X1_172_ (
  .A({ S25957[627] }),
  .ZN({ S7970 })
);
NAND2_X1 #() 
NAND2_X1_432_ (
  .A1({ S7754 }),
  .A2({ S25957[523] }),
  .ZN({ S7971 })
);
AOI21_X1 #() 
AOI21_X1_227_ (
  .A({ S7575 }),
  .B1({ S7730 }),
  .B2({ S9 }),
  .ZN({ S7972 })
);
OAI21_X1 #() 
OAI21_X1_235_ (
  .A({ S7972 }),
  .B1({ S7851 }),
  .B2({ S7971 }),
  .ZN({ S7973 })
);
NAND3_X1 #() 
NAND3_X1_476_ (
  .A1({ S7568 }),
  .A2({ S9 }),
  .A3({ S7596 }),
  .ZN({ S7975 })
);
AOI21_X1 #() 
AOI21_X1_228_ (
  .A({ S9 }),
  .B1({ S6096 }),
  .B2({ S6099 }),
  .ZN({ S7976 })
);
NAND3_X1 #() 
NAND3_X1_477_ (
  .A1({ S7976 }),
  .A2({ S7674 }),
  .A3({ S7620 }),
  .ZN({ S7977 })
);
NAND3_X1 #() 
NAND3_X1_478_ (
  .A1({ S7975 }),
  .A2({ S7575 }),
  .A3({ S7977 }),
  .ZN({ S7978 })
);
NAND3_X1 #() 
NAND3_X1_479_ (
  .A1({ S7973 }),
  .A2({ S7978 }),
  .A3({ S25957[525] }),
  .ZN({ S7979 })
);
NAND2_X1 #() 
NAND2_X1_433_ (
  .A1({ S7613 }),
  .A2({ S25957[523] }),
  .ZN({ S7980 })
);
AOI21_X1 #() 
AOI21_X1_229_ (
  .A({ S7575 }),
  .B1({ S7678 }),
  .B2({ S7596 }),
  .ZN({ S7981 })
);
AOI21_X1 #() 
AOI21_X1_230_ (
  .A({ S9 }),
  .B1({ S7588 }),
  .B2({ S7576 }),
  .ZN({ S7982 })
);
NAND3_X1 #() 
NAND3_X1_480_ (
  .A1({ S7814 }),
  .A2({ S7982 }),
  .A3({ S7596 }),
  .ZN({ S7983 })
);
AOI21_X1 #() 
AOI21_X1_231_ (
  .A({ S25957[524] }),
  .B1({ S7646 }),
  .B2({ S7606 }),
  .ZN({ S7984 })
);
AOI22_X1 #() 
AOI22_X1_35_ (
  .A1({ S7981 }),
  .A2({ S7980 }),
  .B1({ S7983 }),
  .B2({ S7984 }),
  .ZN({ S7986 })
);
AOI21_X1 #() 
AOI21_X1_232_ (
  .A({ S25957[526] }),
  .B1({ S7986 }),
  .B2({ S7605 }),
  .ZN({ S7987 })
);
NAND3_X1 #() 
NAND3_X1_481_ (
  .A1({ S7675 }),
  .A2({ S7567 }),
  .A3({ S25957[523] }),
  .ZN({ S7988 })
);
NAND3_X1 #() 
NAND3_X1_482_ (
  .A1({ S7611 }),
  .A2({ S9 }),
  .A3({ S7637 }),
  .ZN({ S7989 })
);
AOI21_X1 #() 
AOI21_X1_233_ (
  .A({ S7575 }),
  .B1({ S7989 }),
  .B2({ S7988 }),
  .ZN({ S7990 })
);
NAND2_X1 #() 
NAND2_X1_434_ (
  .A1({ S7928 }),
  .A2({ S7760 }),
  .ZN({ S7991 })
);
INV_X1 #() 
INV_X1_173_ (
  .A({ S7991 }),
  .ZN({ S7992 })
);
OAI21_X1 #() 
OAI21_X1_236_ (
  .A({ S7605 }),
  .B1({ S7990 }),
  .B2({ S7992 }),
  .ZN({ S7993 })
);
OAI211_X1 #() 
OAI211_X1_122_ (
  .A({ S9 }),
  .B({ S7580 }),
  .C1({ S7579 }),
  .C2({ S7572 }),
  .ZN({ S7994 })
);
AND3_X1 #() 
AND3_X1_16_ (
  .A1({ S7994 }),
  .A2({ S7933 }),
  .A3({ S25957[524] }),
  .ZN({ S7995 })
);
NAND4_X1 #() 
NAND4_X1_45_ (
  .A1({ S7620 }),
  .A2({ S7596 }),
  .A3({ S7567 }),
  .A4({ S25957[523] }),
  .ZN({ S7997 })
);
NAND4_X1 #() 
NAND4_X1_46_ (
  .A1({ S7620 }),
  .A2({ S7579 }),
  .A3({ S7580 }),
  .A4({ S9 }),
  .ZN({ S7998 })
);
AOI21_X1 #() 
AOI21_X1_234_ (
  .A({ S25957[524] }),
  .B1({ S7997 }),
  .B2({ S7998 }),
  .ZN({ S7999 })
);
OAI21_X1 #() 
OAI21_X1_237_ (
  .A({ S25957[525] }),
  .B1({ S7995 }),
  .B2({ S7999 }),
  .ZN({ S8000 })
);
NAND2_X1 #() 
NAND2_X1_435_ (
  .A1({ S7993 }),
  .A2({ S8000 }),
  .ZN({ S8001 })
);
AOI22_X1 #() 
AOI22_X1_36_ (
  .A1({ S8001 }),
  .A2({ S25957[526] }),
  .B1({ S7987 }),
  .B2({ S7979 }),
  .ZN({ S8002 })
);
NAND2_X1 #() 
NAND2_X1_436_ (
  .A1({ S7638 }),
  .A2({ S7925 }),
  .ZN({ S8003 })
);
NAND2_X1 #() 
NAND2_X1_437_ (
  .A1({ S8003 }),
  .A2({ S7575 }),
  .ZN({ S8004 })
);
OAI211_X1 #() 
OAI211_X1_123_ (
  .A({ S25957[523] }),
  .B({ S17 }),
  .C1({ S7567 }),
  .C2({ S25957[522] }),
  .ZN({ S8005 })
);
OAI211_X1 #() 
OAI211_X1_124_ (
  .A({ S8005 }),
  .B({ S25957[524] }),
  .C1({ S7808 }),
  .C2({ S7809 }),
  .ZN({ S8006 })
);
OAI211_X1 #() 
OAI211_X1_125_ (
  .A({ S8006 }),
  .B({ S7605 }),
  .C1({ S8004 }),
  .C2({ S7612 }),
  .ZN({ S8008 })
);
NAND2_X1 #() 
NAND2_X1_438_ (
  .A1({ S7606 }),
  .A2({ S7580 }),
  .ZN({ S8009 })
);
AOI21_X1 #() 
AOI21_X1_235_ (
  .A({ S25957[524] }),
  .B1({ S7648 }),
  .B2({ S8009 }),
  .ZN({ S8010 })
);
NAND4_X1 #() 
NAND4_X1_47_ (
  .A1({ S25957[522] }),
  .A2({ S7588 }),
  .A3({ S7576 }),
  .A4({ S25957[523] }),
  .ZN({ S8011 })
);
NAND3_X1 #() 
NAND3_X1_483_ (
  .A1({ S7582 }),
  .A2({ S25957[524] }),
  .A3({ S8011 }),
  .ZN({ S8012 })
);
INV_X1 #() 
INV_X1_174_ (
  .A({ S8012 }),
  .ZN({ S8013 })
);
OAI21_X1 #() 
OAI21_X1_238_ (
  .A({ S25957[525] }),
  .B1({ S8013 }),
  .B2({ S8010 }),
  .ZN({ S8014 })
);
AOI21_X1 #() 
AOI21_X1_236_ (
  .A({ S25957[526] }),
  .B1({ S8008 }),
  .B2({ S8014 }),
  .ZN({ S8015 })
);
NAND4_X1 #() 
NAND4_X1_48_ (
  .A1({ S7624 }),
  .A2({ S7587 }),
  .A3({ S9 }),
  .A4({ S25957[520] }),
  .ZN({ S8016 })
);
NAND3_X1 #() 
NAND3_X1_484_ (
  .A1({ S7639 }),
  .A2({ S7575 }),
  .A3({ S8016 }),
  .ZN({ S8017 })
);
NAND3_X1 #() 
NAND3_X1_485_ (
  .A1({ S7606 }),
  .A2({ S7567 }),
  .A3({ S9 }),
  .ZN({ S8019 })
);
NAND2_X1 #() 
NAND2_X1_439_ (
  .A1({ S8019 }),
  .A2({ S25957[524] }),
  .ZN({ S8020 })
);
NAND3_X1 #() 
NAND3_X1_486_ (
  .A1({ S8017 }),
  .A2({ S7605 }),
  .A3({ S8020 }),
  .ZN({ S8021 })
);
NAND3_X1 #() 
NAND3_X1_487_ (
  .A1({ S7731 }),
  .A2({ S7574 }),
  .A3({ S25957[524] }),
  .ZN({ S8022 })
);
NAND3_X1 #() 
NAND3_X1_488_ (
  .A1({ S7587 }),
  .A2({ S9 }),
  .A3({ S7580 }),
  .ZN({ S8023 })
);
AOI21_X1 #() 
AOI21_X1_237_ (
  .A({ S25957[524] }),
  .B1({ S7804 }),
  .B2({ S7675 }),
  .ZN({ S8024 })
);
AOI21_X1 #() 
AOI21_X1_238_ (
  .A({ S7605 }),
  .B1({ S8024 }),
  .B2({ S8023 }),
  .ZN({ S8025 })
);
NAND2_X1 #() 
NAND2_X1_440_ (
  .A1({ S8022 }),
  .A2({ S8025 }),
  .ZN({ S8026 })
);
AOI21_X1 #() 
AOI21_X1_239_ (
  .A({ S7660 }),
  .B1({ S8026 }),
  .B2({ S8021 }),
  .ZN({ S8027 })
);
OAI21_X1 #() 
OAI21_X1_239_ (
  .A({ S7562 }),
  .B1({ S8015 }),
  .B2({ S8027 }),
  .ZN({ S8028 })
);
OAI211_X1 #() 
OAI211_X1_126_ (
  .A({ S8028 }),
  .B({ S7970 }),
  .C1({ S8002 }),
  .C2({ S7562 }),
  .ZN({ S8030 })
);
NAND2_X1 #() 
NAND2_X1_441_ (
  .A1({ S7987 }),
  .A2({ S7979 }),
  .ZN({ S8031 })
);
INV_X1 #() 
INV_X1_175_ (
  .A({ S7988 }),
  .ZN({ S8032 })
);
AOI21_X1 #() 
AOI21_X1_240_ (
  .A({ S25957[523] }),
  .B1({ S7568 }),
  .B2({ S7626 }),
  .ZN({ S8033 })
);
OAI21_X1 #() 
OAI21_X1_240_ (
  .A({ S25957[524] }),
  .B1({ S8033 }),
  .B2({ S8032 }),
  .ZN({ S8034 })
);
AOI21_X1 #() 
AOI21_X1_241_ (
  .A({ S25957[525] }),
  .B1({ S8034 }),
  .B2({ S7991 }),
  .ZN({ S8035 })
);
AOI21_X1 #() 
AOI21_X1_242_ (
  .A({ S7575 }),
  .B1({ S7994 }),
  .B2({ S7933 }),
  .ZN({ S8036 })
);
AND3_X1 #() 
AND3_X1_17_ (
  .A1({ S7997 }),
  .A2({ S7998 }),
  .A3({ S7575 }),
  .ZN({ S8037 })
);
NOR3_X1 #() 
NOR3_X1_14_ (
  .A1({ S8037 }),
  .A2({ S8036 }),
  .A3({ S7605 }),
  .ZN({ S8038 })
);
OAI21_X1 #() 
OAI21_X1_241_ (
  .A({ S25957[526] }),
  .B1({ S8035 }),
  .B2({ S8038 }),
  .ZN({ S8039 })
);
AOI21_X1 #() 
AOI21_X1_243_ (
  .A({ S7562 }),
  .B1({ S8039 }),
  .B2({ S8031 }),
  .ZN({ S8041 })
);
INV_X1 #() 
INV_X1_176_ (
  .A({ S7612 }),
  .ZN({ S8042 })
);
AOI21_X1 #() 
AOI21_X1_244_ (
  .A({ S25957[524] }),
  .B1({ S8042 }),
  .B2({ S8003 }),
  .ZN({ S8043 })
);
NAND4_X1 #() 
NAND4_X1_49_ (
  .A1({ S7606 }),
  .A2({ S7579 }),
  .A3({ S25957[523] }),
  .A4({ S7580 }),
  .ZN({ S8044 })
);
NAND3_X1 #() 
NAND3_X1_489_ (
  .A1({ S7752 }),
  .A2({ S25957[524] }),
  .A3({ S8044 }),
  .ZN({ S8045 })
);
NAND2_X1 #() 
NAND2_X1_442_ (
  .A1({ S8045 }),
  .A2({ S7605 }),
  .ZN({ S8046 })
);
INV_X1 #() 
INV_X1_177_ (
  .A({ S8010 }),
  .ZN({ S8047 })
);
NAND3_X1 #() 
NAND3_X1_490_ (
  .A1({ S8047 }),
  .A2({ S25957[525] }),
  .A3({ S8012 }),
  .ZN({ S8048 })
);
OAI211_X1 #() 
OAI211_X1_127_ (
  .A({ S8048 }),
  .B({ S7660 }),
  .C1({ S8043 }),
  .C2({ S8046 }),
  .ZN({ S8049 })
);
NAND2_X1 #() 
NAND2_X1_443_ (
  .A1({ S8026 }),
  .A2({ S8021 }),
  .ZN({ S8050 })
);
NAND2_X1 #() 
NAND2_X1_444_ (
  .A1({ S8050 }),
  .A2({ S25957[526] }),
  .ZN({ S8052 })
);
AOI21_X1 #() 
AOI21_X1_245_ (
  .A({ S25957[527] }),
  .B1({ S8052 }),
  .B2({ S8049 }),
  .ZN({ S8053 })
);
OAI21_X1 #() 
OAI21_X1_242_ (
  .A({ S25957[627] }),
  .B1({ S8041 }),
  .B2({ S8053 }),
  .ZN({ S8054 })
);
NAND3_X1 #() 
NAND3_X1_491_ (
  .A1({ S8054 }),
  .A2({ S25957[595] }),
  .A3({ S8030 }),
  .ZN({ S8055 })
);
OAI21_X1 #() 
OAI21_X1_243_ (
  .A({ S7970 }),
  .B1({ S8041 }),
  .B2({ S8053 }),
  .ZN({ S8056 })
);
OAI211_X1 #() 
OAI211_X1_128_ (
  .A({ S8028 }),
  .B({ S25957[627] }),
  .C1({ S8002 }),
  .C2({ S7562 }),
  .ZN({ S8057 })
);
NAND3_X1 #() 
NAND3_X1_492_ (
  .A1({ S8056 }),
  .A2({ S7965 }),
  .A3({ S8057 }),
  .ZN({ S8058 })
);
AOI21_X1 #() 
AOI21_X1_246_ (
  .A({ S7964 }),
  .B1({ S8055 }),
  .B2({ S8058 }),
  .ZN({ S8059 })
);
NAND3_X1 #() 
NAND3_X1_493_ (
  .A1({ S8056 }),
  .A2({ S25957[595] }),
  .A3({ S8057 }),
  .ZN({ S8060 })
);
NAND3_X1 #() 
NAND3_X1_494_ (
  .A1({ S8054 }),
  .A2({ S7965 }),
  .A3({ S8030 }),
  .ZN({ S8061 })
);
AOI21_X1 #() 
AOI21_X1_247_ (
  .A({ S25957[563] }),
  .B1({ S8060 }),
  .B2({ S8061 }),
  .ZN({ S8063 })
);
OAI21_X1 #() 
OAI21_X1_244_ (
  .A({ S6 }),
  .B1({ S8059 }),
  .B2({ S8063 }),
  .ZN({ S8064 })
);
NAND3_X1 #() 
NAND3_X1_495_ (
  .A1({ S8060 }),
  .A2({ S8061 }),
  .A3({ S25957[563] }),
  .ZN({ S8065 })
);
NAND3_X1 #() 
NAND3_X1_496_ (
  .A1({ S8055 }),
  .A2({ S8058 }),
  .A3({ S7964 }),
  .ZN({ S8066 })
);
NAND3_X1 #() 
NAND3_X1_497_ (
  .A1({ S8065 }),
  .A2({ S8066 }),
  .A3({ S25957[531] }),
  .ZN({ S8067 })
);
NAND2_X1 #() 
NAND2_X1_445_ (
  .A1({ S8064 }),
  .A2({ S8067 }),
  .ZN({ S18 })
);
OAI21_X1 #() 
OAI21_X1_245_ (
  .A({ S25957[531] }),
  .B1({ S8059 }),
  .B2({ S8063 }),
  .ZN({ S8068 })
);
NAND3_X1 #() 
NAND3_X1_498_ (
  .A1({ S8065 }),
  .A2({ S8066 }),
  .A3({ S6 }),
  .ZN({ S8069 })
);
NAND2_X1 #() 
NAND2_X1_446_ (
  .A1({ S8068 }),
  .A2({ S8069 }),
  .ZN({ S25957[403] })
);
NAND2_X1 #() 
NAND2_X1_447_ (
  .A1({ S25913 }),
  .A2({ S25882 }),
  .ZN({ S25957[848] })
);
XOR2_X1 #() 
XOR2_X1_10_ (
  .A({ S25957[752] }),
  .B({ S25957[848] }),
  .Z({ S25957[720] })
);
AND2_X1 #() 
AND2_X1_24_ (
  .A1({ S7804 }),
  .A2({ S7675 }),
  .ZN({ S8071 })
);
AOI21_X1 #() 
AOI21_X1_248_ (
  .A({ S25957[523] }),
  .B1({ S7577 }),
  .B2({ S7674 }),
  .ZN({ S8072 })
);
OAI21_X1 #() 
OAI21_X1_246_ (
  .A({ S7575 }),
  .B1({ S8072 }),
  .B2({ S8071 }),
  .ZN({ S8073 })
);
INV_X1 #() 
INV_X1_178_ (
  .A({ S7619 }),
  .ZN({ S8074 })
);
AOI21_X1 #() 
AOI21_X1_249_ (
  .A({ S25957[525] }),
  .B1({ S8074 }),
  .B2({ S7917 }),
  .ZN({ S8075 })
);
NAND2_X1 #() 
NAND2_X1_448_ (
  .A1({ S7971 }),
  .A2({ S8019 }),
  .ZN({ S8076 })
);
NAND3_X1 #() 
NAND3_X1_499_ (
  .A1({ S7675 }),
  .A2({ S9 }),
  .A3({ S7576 }),
  .ZN({ S8077 })
);
NAND3_X1 #() 
NAND3_X1_500_ (
  .A1({ S8076 }),
  .A2({ S25957[524] }),
  .A3({ S8077 }),
  .ZN({ S8078 })
);
NAND2_X1 #() 
NAND2_X1_449_ (
  .A1({ S7736 }),
  .A2({ S7589 }),
  .ZN({ S8079 })
);
NAND2_X1 #() 
NAND2_X1_450_ (
  .A1({ S8079 }),
  .A2({ S7879 }),
  .ZN({ S8081 })
);
AOI21_X1 #() 
AOI21_X1_250_ (
  .A({ S7605 }),
  .B1({ S8081 }),
  .B2({ S7575 }),
  .ZN({ S8082 })
);
AOI22_X1 #() 
AOI22_X1_37_ (
  .A1({ S8082 }),
  .A2({ S8078 }),
  .B1({ S8075 }),
  .B2({ S8073 }),
  .ZN({ S8083 })
);
NAND2_X1 #() 
NAND2_X1_451_ (
  .A1({ S7573 }),
  .A2({ S7885 }),
  .ZN({ S8084 })
);
NAND3_X1 #() 
NAND3_X1_501_ (
  .A1({ S8084 }),
  .A2({ S7575 }),
  .A3({ S7939 }),
  .ZN({ S8085 })
);
OAI211_X1 #() 
OAI211_X1_129_ (
  .A({ S7935 }),
  .B({ S25957[524] }),
  .C1({ S9 }),
  .C2({ S7736 }),
  .ZN({ S8086 })
);
NAND3_X1 #() 
NAND3_X1_502_ (
  .A1({ S8086 }),
  .A2({ S8085 }),
  .A3({ S25957[525] }),
  .ZN({ S8087 })
);
NAND3_X1 #() 
NAND3_X1_503_ (
  .A1({ S7663 }),
  .A2({ S7579 }),
  .A3({ S7580 }),
  .ZN({ S8088 })
);
NAND3_X1 #() 
NAND3_X1_504_ (
  .A1({ S7897 }),
  .A2({ S25957[524] }),
  .A3({ S8088 }),
  .ZN({ S8089 })
);
NAND3_X1 #() 
NAND3_X1_505_ (
  .A1({ S7583 }),
  .A2({ S7661 }),
  .A3({ S7674 }),
  .ZN({ S8090 })
);
NOR2_X1 #() 
NOR2_X1_91_ (
  .A1({ S7634 }),
  .A2({ S25957[524] }),
  .ZN({ S8092 })
);
AOI21_X1 #() 
AOI21_X1_251_ (
  .A({ S25957[525] }),
  .B1({ S8092 }),
  .B2({ S8090 }),
  .ZN({ S8093 })
);
NAND2_X1 #() 
NAND2_X1_452_ (
  .A1({ S8089 }),
  .A2({ S8093 }),
  .ZN({ S8094 })
);
NAND3_X1 #() 
NAND3_X1_506_ (
  .A1({ S8087 }),
  .A2({ S8094 }),
  .A3({ S25957[526] }),
  .ZN({ S8095 })
);
OAI211_X1 #() 
OAI211_X1_130_ (
  .A({ S8095 }),
  .B({ S25957[527] }),
  .C1({ S8083 }),
  .C2({ S25957[526] }),
  .ZN({ S8096 })
);
NAND3_X1 #() 
NAND3_X1_507_ (
  .A1({ S7721 }),
  .A2({ S25957[523] }),
  .A3({ S7572 }),
  .ZN({ S8097 })
);
AOI21_X1 #() 
AOI21_X1_252_ (
  .A({ S25957[523] }),
  .B1({ S16 }),
  .B2({ S25957[522] }),
  .ZN({ S8098 })
);
AOI21_X1 #() 
AOI21_X1_253_ (
  .A({ S7575 }),
  .B1({ S8098 }),
  .B2({ S7827 }),
  .ZN({ S8099 })
);
NAND3_X1 #() 
NAND3_X1_508_ (
  .A1({ S7637 }),
  .A2({ S7754 }),
  .A3({ S9 }),
  .ZN({ S8100 })
);
AOI21_X1 #() 
AOI21_X1_254_ (
  .A({ S25957[524] }),
  .B1({ S7814 }),
  .B2({ S7982 }),
  .ZN({ S8101 })
);
AOI22_X1 #() 
AOI22_X1_38_ (
  .A1({ S8099 }),
  .A2({ S8097 }),
  .B1({ S8101 }),
  .B2({ S8100 }),
  .ZN({ S8103 })
);
OAI211_X1 #() 
OAI211_X1_131_ (
  .A({ S7933 }),
  .B({ S25957[524] }),
  .C1({ S7749 }),
  .C2({ S7805 }),
  .ZN({ S8104 })
);
OAI21_X1 #() 
OAI21_X1_247_ (
  .A({ S7575 }),
  .B1({ S7712 }),
  .B2({ S7711 }),
  .ZN({ S8105 })
);
OAI211_X1 #() 
OAI211_X1_132_ (
  .A({ S8104 }),
  .B({ S25957[525] }),
  .C1({ S8105 }),
  .C2({ S7792 }),
  .ZN({ S8106 })
);
OAI211_X1 #() 
OAI211_X1_133_ (
  .A({ S8106 }),
  .B({ S7660 }),
  .C1({ S8103 }),
  .C2({ S25957[525] }),
  .ZN({ S8107 })
);
NOR2_X1 #() 
NOR2_X1_92_ (
  .A1({ S7801 }),
  .A2({ S25957[522] }),
  .ZN({ S8108 })
);
NOR2_X1 #() 
NOR2_X1_93_ (
  .A1({ S7579 }),
  .A2({ S7572 }),
  .ZN({ S8109 })
);
OAI21_X1 #() 
OAI21_X1_248_ (
  .A({ S25957[523] }),
  .B1({ S8109 }),
  .B2({ S8108 }),
  .ZN({ S8110 })
);
NAND4_X1 #() 
NAND4_X1_50_ (
  .A1({ S7814 }),
  .A2({ S7982 }),
  .A3({ S7596 }),
  .A4({ S7610 }),
  .ZN({ S8111 })
);
AOI21_X1 #() 
AOI21_X1_255_ (
  .A({ S7575 }),
  .B1({ S7678 }),
  .B2({ S7579 }),
  .ZN({ S8112 })
);
AOI22_X1 #() 
AOI22_X1_39_ (
  .A1({ S8110 }),
  .A2({ S8092 }),
  .B1({ S8112 }),
  .B2({ S8111 }),
  .ZN({ S8114 })
);
NAND3_X1 #() 
NAND3_X1_509_ (
  .A1({ S7817 }),
  .A2({ S7828 }),
  .A3({ S7575 }),
  .ZN({ S8115 })
);
OAI211_X1 #() 
OAI211_X1_134_ (
  .A({ S7719 }),
  .B({ S25957[524] }),
  .C1({ S9 }),
  .C2({ S25957[520] }),
  .ZN({ S8116 })
);
NAND3_X1 #() 
NAND3_X1_510_ (
  .A1({ S8116 }),
  .A2({ S8115 }),
  .A3({ S7605 }),
  .ZN({ S8117 })
);
OAI211_X1 #() 
OAI211_X1_135_ (
  .A({ S8117 }),
  .B({ S25957[526] }),
  .C1({ S8114 }),
  .C2({ S7605 }),
  .ZN({ S8118 })
);
NAND3_X1 #() 
NAND3_X1_511_ (
  .A1({ S8118 }),
  .A2({ S8107 }),
  .A3({ S7562 }),
  .ZN({ S8119 })
);
NAND3_X1 #() 
NAND3_X1_512_ (
  .A1({ S8096 }),
  .A2({ S8119 }),
  .A3({ S25957[720] }),
  .ZN({ S8120 })
);
INV_X1 #() 
INV_X1_179_ (
  .A({ S8120 }),
  .ZN({ S8121 })
);
AOI21_X1 #() 
AOI21_X1_256_ (
  .A({ S25957[720] }),
  .B1({ S8096 }),
  .B2({ S8119 }),
  .ZN({ S8122 })
);
OAI21_X1 #() 
OAI21_X1_249_ (
  .A({ S25957[656] }),
  .B1({ S8121 }),
  .B2({ S8122 }),
  .ZN({ S8123 })
);
INV_X1 #() 
INV_X1_180_ (
  .A({ S25957[720] }),
  .ZN({ S8125 })
);
NAND2_X1 #() 
NAND2_X1_453_ (
  .A1({ S8096 }),
  .A2({ S8119 }),
  .ZN({ S8126 })
);
NAND2_X1 #() 
NAND2_X1_454_ (
  .A1({ S8126 }),
  .A2({ S8125 }),
  .ZN({ S8127 })
);
NAND3_X1 #() 
NAND3_X1_513_ (
  .A1({ S8127 }),
  .A2({ S5282 }),
  .A3({ S8120 }),
  .ZN({ S8128 })
);
NAND2_X1 #() 
NAND2_X1_455_ (
  .A1({ S8123 }),
  .A2({ S8128 }),
  .ZN({ S25957[400] })
);
NOR2_X1 #() 
NOR2_X1_94_ (
  .A1({ S5355 }),
  .A2({ S5356 }),
  .ZN({ S25957[721] })
);
NAND3_X1 #() 
NAND3_X1_514_ (
  .A1({ S5333 }),
  .A2({ S5349 }),
  .A3({ S25957[721] }),
  .ZN({ S8129 })
);
INV_X1 #() 
INV_X1_181_ (
  .A({ S25957[721] }),
  .ZN({ S8130 })
);
NAND3_X1 #() 
NAND3_X1_515_ (
  .A1({ S5352 }),
  .A2({ S5351 }),
  .A3({ S8130 }),
  .ZN({ S8131 })
);
NAND3_X1 #() 
NAND3_X1_516_ (
  .A1({ S8129 }),
  .A2({ S8131 }),
  .A3({ S25957[785] }),
  .ZN({ S8132 })
);
NAND3_X1 #() 
NAND3_X1_517_ (
  .A1({ S5333 }),
  .A2({ S5349 }),
  .A3({ S8130 }),
  .ZN({ S8134 })
);
NAND3_X1 #() 
NAND3_X1_518_ (
  .A1({ S5352 }),
  .A2({ S5351 }),
  .A3({ S25957[721] }),
  .ZN({ S8135 })
);
NAND3_X1 #() 
NAND3_X1_519_ (
  .A1({ S8134 }),
  .A2({ S8135 }),
  .A3({ S4249 }),
  .ZN({ S8136 })
);
NAND2_X1 #() 
NAND2_X1_456_ (
  .A1({ S8132 }),
  .A2({ S8136 }),
  .ZN({ S8137 })
);
XNOR2_X1 #() 
XNOR2_X1_15_ (
  .A({ S25957[721] }),
  .B({ S5286 }),
  .ZN({ S25957[689] })
);
NAND2_X1 #() 
NAND2_X1_457_ (
  .A1({ S5352 }),
  .A2({ S5351 }),
  .ZN({ S25957[625] })
);
INV_X1 #() 
INV_X1_182_ (
  .A({ S25957[625] }),
  .ZN({ S8138 })
);
NOR3_X1 #() 
NOR3_X1_15_ (
  .A1({ S7615 }),
  .A2({ S7900 }),
  .A3({ S25957[524] }),
  .ZN({ S8139 })
);
NAND3_X1 #() 
NAND3_X1_520_ (
  .A1({ S7802 }),
  .A2({ S9 }),
  .A3({ S7624 }),
  .ZN({ S8140 })
);
NAND2_X1 #() 
NAND2_X1_458_ (
  .A1({ S8140 }),
  .A2({ S7746 }),
  .ZN({ S8141 })
);
NAND2_X1 #() 
NAND2_X1_459_ (
  .A1({ S8141 }),
  .A2({ S7605 }),
  .ZN({ S8143 })
);
AOI21_X1 #() 
AOI21_X1_257_ (
  .A({ S9 }),
  .B1({ S7611 }),
  .B2({ S7610 }),
  .ZN({ S8144 })
);
NAND3_X1 #() 
NAND3_X1_521_ (
  .A1({ S7835 }),
  .A2({ S8023 }),
  .A3({ S7575 }),
  .ZN({ S8145 })
);
OAI21_X1 #() 
OAI21_X1_250_ (
  .A({ S25957[524] }),
  .B1({ S7622 }),
  .B2({ S25957[523] }),
  .ZN({ S8146 })
);
OAI211_X1 #() 
OAI211_X1_136_ (
  .A({ S25957[525] }),
  .B({ S8145 }),
  .C1({ S8144 }),
  .C2({ S8146 }),
  .ZN({ S8147 })
);
OAI21_X1 #() 
OAI21_X1_251_ (
  .A({ S8147 }),
  .B1({ S8139 }),
  .B2({ S8143 }),
  .ZN({ S8148 })
);
NAND2_X1 #() 
NAND2_X1_460_ (
  .A1({ S8077 }),
  .A2({ S25957[524] }),
  .ZN({ S8149 })
);
NAND2_X1 #() 
NAND2_X1_461_ (
  .A1({ S7606 }),
  .A2({ S7567 }),
  .ZN({ S8150 })
);
OAI211_X1 #() 
OAI211_X1_137_ (
  .A({ S7621 }),
  .B({ S7575 }),
  .C1({ S7667 }),
  .C2({ S8150 }),
  .ZN({ S8151 })
);
OAI211_X1 #() 
OAI211_X1_138_ (
  .A({ S8151 }),
  .B({ S7605 }),
  .C1({ S7803 }),
  .C2({ S8149 }),
  .ZN({ S8152 })
);
AOI21_X1 #() 
AOI21_X1_258_ (
  .A({ S9 }),
  .B1({ S7568 }),
  .B2({ S7925 }),
  .ZN({ S8154 })
);
NAND3_X1 #() 
NAND3_X1_522_ (
  .A1({ S7628 }),
  .A2({ S7988 }),
  .A3({ S25957[524] }),
  .ZN({ S8155 })
);
OAI21_X1 #() 
OAI21_X1_252_ (
  .A({ S7575 }),
  .B1({ S8109 }),
  .B2({ S25957[523] }),
  .ZN({ S8156 })
);
OAI211_X1 #() 
OAI211_X1_139_ (
  .A({ S25957[525] }),
  .B({ S8155 }),
  .C1({ S8154 }),
  .C2({ S8156 }),
  .ZN({ S8157 })
);
NAND3_X1 #() 
NAND3_X1_523_ (
  .A1({ S8152 }),
  .A2({ S8157 }),
  .A3({ S25957[526] }),
  .ZN({ S8158 })
);
OAI211_X1 #() 
OAI211_X1_140_ (
  .A({ S8158 }),
  .B({ S25957[527] }),
  .C1({ S8148 }),
  .C2({ S25957[526] }),
  .ZN({ S8159 })
);
AOI21_X1 #() 
AOI21_X1_259_ (
  .A({ S25957[524] }),
  .B1({ S7843 }),
  .B2({ S9 }),
  .ZN({ S8160 })
);
AOI21_X1 #() 
AOI21_X1_260_ (
  .A({ S7575 }),
  .B1({ S7977 }),
  .B2({ S7881 }),
  .ZN({ S8161 })
);
OAI21_X1 #() 
OAI21_X1_253_ (
  .A({ S25957[525] }),
  .B1({ S8160 }),
  .B2({ S8161 }),
  .ZN({ S8162 })
);
NAND3_X1 #() 
NAND3_X1_524_ (
  .A1({ S7664 }),
  .A2({ S25957[524] }),
  .A3({ S7888 }),
  .ZN({ S8163 })
);
NAND2_X1 #() 
NAND2_X1_462_ (
  .A1({ S8016 }),
  .A2({ S7682 }),
  .ZN({ S8165 })
);
NAND3_X1 #() 
NAND3_X1_525_ (
  .A1({ S8163 }),
  .A2({ S7605 }),
  .A3({ S8165 }),
  .ZN({ S8166 })
);
NAND3_X1 #() 
NAND3_X1_526_ (
  .A1({ S8162 }),
  .A2({ S7660 }),
  .A3({ S8166 }),
  .ZN({ S8167 })
);
NAND3_X1 #() 
NAND3_X1_527_ (
  .A1({ S7754 }),
  .A2({ S9 }),
  .A3({ S7674 }),
  .ZN({ S8168 })
);
NAND3_X1 #() 
NAND3_X1_528_ (
  .A1({ S8168 }),
  .A2({ S25957[524] }),
  .A3({ S8044 }),
  .ZN({ S8169 })
);
OAI211_X1 #() 
OAI211_X1_141_ (
  .A({ S7575 }),
  .B({ S7606 }),
  .C1({ S7634 }),
  .C2({ S25957[521] }),
  .ZN({ S8170 })
);
NAND3_X1 #() 
NAND3_X1_529_ (
  .A1({ S8169 }),
  .A2({ S25957[525] }),
  .A3({ S8170 }),
  .ZN({ S8171 })
);
OAI21_X1 #() 
OAI21_X1_254_ (
  .A({ S25957[524] }),
  .B1({ S7667 }),
  .B2({ S7796 }),
  .ZN({ S8172 })
);
NAND3_X1 #() 
NAND3_X1_530_ (
  .A1({ S7761 }),
  .A2({ S7575 }),
  .A3({ S8088 }),
  .ZN({ S8173 })
);
OAI211_X1 #() 
OAI211_X1_142_ (
  .A({ S8173 }),
  .B({ S7605 }),
  .C1({ S8172 }),
  .C2({ S8154 }),
  .ZN({ S8174 })
);
NAND3_X1 #() 
NAND3_X1_531_ (
  .A1({ S8174 }),
  .A2({ S8171 }),
  .A3({ S25957[526] }),
  .ZN({ S8176 })
);
NAND3_X1 #() 
NAND3_X1_532_ (
  .A1({ S8167 }),
  .A2({ S8176 }),
  .A3({ S7562 }),
  .ZN({ S8177 })
);
NAND3_X1 #() 
NAND3_X1_533_ (
  .A1({ S8159 }),
  .A2({ S8177 }),
  .A3({ S8138 }),
  .ZN({ S8178 })
);
NAND2_X1 #() 
NAND2_X1_463_ (
  .A1({ S8152 }),
  .A2({ S8157 }),
  .ZN({ S8179 })
);
NAND2_X1 #() 
NAND2_X1_464_ (
  .A1({ S8179 }),
  .A2({ S25957[526] }),
  .ZN({ S8180 })
);
NAND2_X1 #() 
NAND2_X1_465_ (
  .A1({ S8148 }),
  .A2({ S7660 }),
  .ZN({ S8181 })
);
NAND3_X1 #() 
NAND3_X1_534_ (
  .A1({ S8181 }),
  .A2({ S8180 }),
  .A3({ S25957[527] }),
  .ZN({ S8182 })
);
NAND2_X1 #() 
NAND2_X1_466_ (
  .A1({ S8174 }),
  .A2({ S8171 }),
  .ZN({ S8183 })
);
NAND2_X1 #() 
NAND2_X1_467_ (
  .A1({ S8183 }),
  .A2({ S25957[526] }),
  .ZN({ S8184 })
);
NAND2_X1 #() 
NAND2_X1_468_ (
  .A1({ S7977 }),
  .A2({ S7881 }),
  .ZN({ S8185 })
);
NAND2_X1 #() 
NAND2_X1_469_ (
  .A1({ S8185 }),
  .A2({ S25957[524] }),
  .ZN({ S8187 })
);
AOI21_X1 #() 
AOI21_X1_261_ (
  .A({ S7605 }),
  .B1({ S8187 }),
  .B2({ S7608 }),
  .ZN({ S8188 })
);
AND3_X1 #() 
AND3_X1_18_ (
  .A1({ S8163 }),
  .A2({ S7605 }),
  .A3({ S8165 }),
  .ZN({ S8189 })
);
OAI21_X1 #() 
OAI21_X1_255_ (
  .A({ S7660 }),
  .B1({ S8188 }),
  .B2({ S8189 }),
  .ZN({ S8190 })
);
NAND3_X1 #() 
NAND3_X1_535_ (
  .A1({ S8184 }),
  .A2({ S8190 }),
  .A3({ S7562 }),
  .ZN({ S8191 })
);
NAND3_X1 #() 
NAND3_X1_536_ (
  .A1({ S8182 }),
  .A2({ S8191 }),
  .A3({ S25957[625] }),
  .ZN({ S8192 })
);
AOI21_X1 #() 
AOI21_X1_262_ (
  .A({ S25957[689] }),
  .B1({ S8192 }),
  .B2({ S8178 }),
  .ZN({ S8193 })
);
INV_X1 #() 
INV_X1_183_ (
  .A({ S25957[689] }),
  .ZN({ S8194 })
);
NAND3_X1 #() 
NAND3_X1_537_ (
  .A1({ S8182 }),
  .A2({ S8191 }),
  .A3({ S8138 }),
  .ZN({ S8195 })
);
NAND3_X1 #() 
NAND3_X1_538_ (
  .A1({ S8159 }),
  .A2({ S8177 }),
  .A3({ S25957[625] }),
  .ZN({ S8196 })
);
AOI21_X1 #() 
AOI21_X1_263_ (
  .A({ S8194 }),
  .B1({ S8195 }),
  .B2({ S8196 }),
  .ZN({ S8198 })
);
OAI21_X1 #() 
OAI21_X1_256_ (
  .A({ S8137 }),
  .B1({ S8193 }),
  .B2({ S8198 }),
  .ZN({ S8199 })
);
NAND3_X1 #() 
NAND3_X1_539_ (
  .A1({ S8195 }),
  .A2({ S8194 }),
  .A3({ S8196 }),
  .ZN({ S8200 })
);
NAND3_X1 #() 
NAND3_X1_540_ (
  .A1({ S8192 }),
  .A2({ S25957[689] }),
  .A3({ S8178 }),
  .ZN({ S8201 })
);
NAND3_X1 #() 
NAND3_X1_541_ (
  .A1({ S8200 }),
  .A2({ S8201 }),
  .A3({ S25957[529] }),
  .ZN({ S8202 })
);
NAND2_X1 #() 
NAND2_X1_470_ (
  .A1({ S8199 }),
  .A2({ S8202 }),
  .ZN({ S25957[401] })
);
NAND2_X1 #() 
NAND2_X1_471_ (
  .A1({ S5451 }),
  .A2({ S5454 }),
  .ZN({ S25957[562] })
);
NOR2_X1 #() 
NOR2_X1_95_ (
  .A1({ S2886 }),
  .A2({ S2865 }),
  .ZN({ S8203 })
);
INV_X1 #() 
INV_X1_184_ (
  .A({ S8203 }),
  .ZN({ S25957[722] })
);
NOR2_X1 #() 
NOR2_X1_96_ (
  .A1({ S7593 }),
  .A2({ S25957[524] }),
  .ZN({ S8204 })
);
OAI21_X1 #() 
OAI21_X1_257_ (
  .A({ S8204 }),
  .B1({ S7851 }),
  .B2({ S7902 }),
  .ZN({ S8206 })
);
AOI21_X1 #() 
AOI21_X1_264_ (
  .A({ S7575 }),
  .B1({ S7597 }),
  .B2({ S7587 }),
  .ZN({ S8207 })
);
AOI21_X1 #() 
AOI21_X1_265_ (
  .A({ S7605 }),
  .B1({ S8207 }),
  .B2({ S8084 }),
  .ZN({ S8208 })
);
NAND2_X1 #() 
NAND2_X1_472_ (
  .A1({ S8208 }),
  .A2({ S8206 }),
  .ZN({ S8209 })
);
NAND2_X1 #() 
NAND2_X1_473_ (
  .A1({ S7896 }),
  .A2({ S9 }),
  .ZN({ S8210 })
);
NAND3_X1 #() 
NAND3_X1_542_ (
  .A1({ S7679 }),
  .A2({ S7638 }),
  .A3({ S7637 }),
  .ZN({ S8211 })
);
AOI22_X1 #() 
AOI22_X1_40_ (
  .A1({ S7853 }),
  .A2({ S8211 }),
  .B1({ S7889 }),
  .B2({ S8210 }),
  .ZN({ S8212 })
);
NAND2_X1 #() 
NAND2_X1_474_ (
  .A1({ S8212 }),
  .A2({ S7605 }),
  .ZN({ S8213 })
);
NAND3_X1 #() 
NAND3_X1_543_ (
  .A1({ S8213 }),
  .A2({ S25957[526] }),
  .A3({ S8209 }),
  .ZN({ S8214 })
);
NAND3_X1 #() 
NAND3_X1_544_ (
  .A1({ S7596 }),
  .A2({ S25957[523] }),
  .A3({ S25957[520] }),
  .ZN({ S8215 })
);
NAND3_X1 #() 
NAND3_X1_545_ (
  .A1({ S8016 }),
  .A2({ S25957[524] }),
  .A3({ S8215 }),
  .ZN({ S8217 })
);
AOI21_X1 #() 
AOI21_X1_266_ (
  .A({ S25957[524] }),
  .B1({ S16 }),
  .B2({ S25957[523] }),
  .ZN({ S8218 })
);
NAND3_X1 #() 
NAND3_X1_546_ (
  .A1({ S7930 }),
  .A2({ S8218 }),
  .A3({ S7899 }),
  .ZN({ S8219 })
);
NAND3_X1 #() 
NAND3_X1_547_ (
  .A1({ S8217 }),
  .A2({ S8219 }),
  .A3({ S25957[525] }),
  .ZN({ S8220 })
);
NAND2_X1 #() 
NAND2_X1_475_ (
  .A1({ S7976 }),
  .A2({ S7674 }),
  .ZN({ S8221 })
);
NAND3_X1 #() 
NAND3_X1_548_ (
  .A1({ S8221 }),
  .A2({ S7809 }),
  .A3({ S25957[524] }),
  .ZN({ S8222 })
);
OAI211_X1 #() 
OAI211_X1_143_ (
  .A({ S7618 }),
  .B({ S7575 }),
  .C1({ S7661 }),
  .C2({ S7610 }),
  .ZN({ S8223 })
);
NAND3_X1 #() 
NAND3_X1_549_ (
  .A1({ S8223 }),
  .A2({ S8222 }),
  .A3({ S7605 }),
  .ZN({ S8224 })
);
NAND3_X1 #() 
NAND3_X1_550_ (
  .A1({ S7660 }),
  .A2({ S8220 }),
  .A3({ S8224 }),
  .ZN({ S8225 })
);
NAND3_X1 #() 
NAND3_X1_551_ (
  .A1({ S8214 }),
  .A2({ S25957[527] }),
  .A3({ S8225 }),
  .ZN({ S8226 })
);
AOI21_X1 #() 
AOI21_X1_267_ (
  .A({ S25957[524] }),
  .B1({ S7724 }),
  .B2({ S7662 }),
  .ZN({ S8228 })
);
NAND3_X1 #() 
NAND3_X1_552_ (
  .A1({ S7591 }),
  .A2({ S7814 }),
  .A3({ S25957[523] }),
  .ZN({ S8229 })
);
NAND2_X1 #() 
NAND2_X1_476_ (
  .A1({ S8229 }),
  .A2({ S8228 }),
  .ZN({ S8230 })
);
AOI21_X1 #() 
AOI21_X1_268_ (
  .A({ S7575 }),
  .B1({ S7597 }),
  .B2({ S7651 }),
  .ZN({ S8231 })
);
NAND2_X1 #() 
NAND2_X1_477_ (
  .A1({ S8231 }),
  .A2({ S7975 }),
  .ZN({ S8232 })
);
NAND3_X1 #() 
NAND3_X1_553_ (
  .A1({ S8232 }),
  .A2({ S8230 }),
  .A3({ S25957[525] }),
  .ZN({ S8233 })
);
NAND3_X1 #() 
NAND3_X1_554_ (
  .A1({ S7679 }),
  .A2({ S9 }),
  .A3({ S7637 }),
  .ZN({ S8234 })
);
NAND3_X1 #() 
NAND3_X1_555_ (
  .A1({ S8110 }),
  .A2({ S7575 }),
  .A3({ S8234 }),
  .ZN({ S8235 })
);
OAI211_X1 #() 
OAI211_X1_144_ (
  .A({ S25957[524] }),
  .B({ S8221 }),
  .C1({ S7826 }),
  .C2({ S25957[523] }),
  .ZN({ S8236 })
);
NAND3_X1 #() 
NAND3_X1_556_ (
  .A1({ S8235 }),
  .A2({ S7605 }),
  .A3({ S8236 }),
  .ZN({ S8237 })
);
NAND3_X1 #() 
NAND3_X1_557_ (
  .A1({ S8237 }),
  .A2({ S7660 }),
  .A3({ S8233 }),
  .ZN({ S8239 })
);
OAI21_X1 #() 
OAI21_X1_258_ (
  .A({ S25957[525] }),
  .B1({ S7745 }),
  .B2({ S7599 }),
  .ZN({ S8240 })
);
NOR2_X1 #() 
NOR2_X1_97_ (
  .A1({ S7672 }),
  .A2({ S8240 }),
  .ZN({ S8241 })
);
NAND4_X1 #() 
NAND4_X1_51_ (
  .A1({ S7620 }),
  .A2({ S7596 }),
  .A3({ S7567 }),
  .A4({ S9 }),
  .ZN({ S8242 })
);
AOI21_X1 #() 
AOI21_X1_269_ (
  .A({ S25957[525] }),
  .B1({ S7976 }),
  .B2({ S7674 }),
  .ZN({ S8243 })
);
NAND2_X1 #() 
NAND2_X1_478_ (
  .A1({ S8243 }),
  .A2({ S8242 }),
  .ZN({ S8244 })
);
NAND2_X1 #() 
NAND2_X1_479_ (
  .A1({ S8244 }),
  .A2({ S7575 }),
  .ZN({ S8245 })
);
NAND2_X1 #() 
NAND2_X1_480_ (
  .A1({ S7597 }),
  .A2({ S7802 }),
  .ZN({ S8246 })
);
AOI21_X1 #() 
AOI21_X1_270_ (
  .A({ S25957[525] }),
  .B1({ S7662 }),
  .B2({ S25957[522] }),
  .ZN({ S8247 })
);
NAND2_X1 #() 
NAND2_X1_481_ (
  .A1({ S7589 }),
  .A2({ S7596 }),
  .ZN({ S8248 })
);
AOI22_X1 #() 
AOI22_X1_41_ (
  .A1({ S8247 }),
  .A2({ S8246 }),
  .B1({ S8248 }),
  .B2({ S25957[525] }),
  .ZN({ S8250 })
);
OAI22_X1 #() 
OAI22_X1_13_ (
  .A1({ S8241 }),
  .A2({ S8245 }),
  .B1({ S8250 }),
  .B2({ S8020 }),
  .ZN({ S8251 })
);
NAND2_X1 #() 
NAND2_X1_482_ (
  .A1({ S8251 }),
  .A2({ S25957[526] }),
  .ZN({ S8252 })
);
NAND3_X1 #() 
NAND3_X1_558_ (
  .A1({ S8252 }),
  .A2({ S8239 }),
  .A3({ S7562 }),
  .ZN({ S8253 })
);
NAND3_X1 #() 
NAND3_X1_559_ (
  .A1({ S8253 }),
  .A2({ S8226 }),
  .A3({ S25957[722] }),
  .ZN({ S8254 })
);
AOI22_X1 #() 
AOI22_X1_42_ (
  .A1({ S8212 }),
  .A2({ S7605 }),
  .B1({ S8208 }),
  .B2({ S8206 }),
  .ZN({ S8255 })
);
NAND2_X1 #() 
NAND2_X1_483_ (
  .A1({ S8220 }),
  .A2({ S8224 }),
  .ZN({ S8256 })
);
NAND2_X1 #() 
NAND2_X1_484_ (
  .A1({ S8256 }),
  .A2({ S7660 }),
  .ZN({ S8257 })
);
OAI211_X1 #() 
OAI211_X1_145_ (
  .A({ S8257 }),
  .B({ S25957[527] }),
  .C1({ S8255 }),
  .C2({ S7660 }),
  .ZN({ S8258 })
);
OAI221_X1 #() 
OAI221_X1_7_ (
  .A({ S25957[526] }),
  .B1({ S8250 }),
  .B2({ S8020 }),
  .C1({ S8245 }),
  .C2({ S8241 }),
  .ZN({ S8259 })
);
INV_X1 #() 
INV_X1_185_ (
  .A({ S8221 }),
  .ZN({ S8261 })
);
OAI21_X1 #() 
OAI21_X1_259_ (
  .A({ S25957[524] }),
  .B1({ S7905 }),
  .B2({ S8261 }),
  .ZN({ S8262 })
);
AND3_X1 #() 
AND3_X1_19_ (
  .A1({ S7679 }),
  .A2({ S7637 }),
  .A3({ S9 }),
  .ZN({ S8263 })
);
OAI21_X1 #() 
OAI21_X1_260_ (
  .A({ S7575 }),
  .B1({ S8263 }),
  .B2({ S7748 }),
  .ZN({ S8264 })
);
NAND3_X1 #() 
NAND3_X1_560_ (
  .A1({ S8264 }),
  .A2({ S7605 }),
  .A3({ S8262 }),
  .ZN({ S8265 })
);
NAND2_X1 #() 
NAND2_X1_485_ (
  .A1({ S8232 }),
  .A2({ S8230 }),
  .ZN({ S8266 })
);
NAND2_X1 #() 
NAND2_X1_486_ (
  .A1({ S8266 }),
  .A2({ S25957[525] }),
  .ZN({ S8267 })
);
NAND3_X1 #() 
NAND3_X1_561_ (
  .A1({ S8265 }),
  .A2({ S8267 }),
  .A3({ S7660 }),
  .ZN({ S8268 })
);
NAND3_X1 #() 
NAND3_X1_562_ (
  .A1({ S8268 }),
  .A2({ S7562 }),
  .A3({ S8259 }),
  .ZN({ S8269 })
);
NAND3_X1 #() 
NAND3_X1_563_ (
  .A1({ S8269 }),
  .A2({ S8203 }),
  .A3({ S8258 }),
  .ZN({ S8270 })
);
AOI21_X1 #() 
AOI21_X1_271_ (
  .A({ S25957[562] }),
  .B1({ S8270 }),
  .B2({ S8254 }),
  .ZN({ S8272 })
);
AND3_X1 #() 
AND3_X1_20_ (
  .A1({ S8270 }),
  .A2({ S8254 }),
  .A3({ S25957[562] }),
  .ZN({ S8273 })
);
OAI21_X1 #() 
OAI21_X1_261_ (
  .A({ S25957[530] }),
  .B1({ S8273 }),
  .B2({ S8272 }),
  .ZN({ S8274 })
);
NAND3_X1 #() 
NAND3_X1_564_ (
  .A1({ S5452 }),
  .A2({ S5453 }),
  .A3({ S25957[722] }),
  .ZN({ S8275 })
);
NAND3_X1 #() 
NAND3_X1_565_ (
  .A1({ S5418 }),
  .A2({ S5450 }),
  .A3({ S8203 }),
  .ZN({ S8276 })
);
NAND3_X1 #() 
NAND3_X1_566_ (
  .A1({ S8275 }),
  .A2({ S8276 }),
  .A3({ S4170 }),
  .ZN({ S8277 })
);
NAND3_X1 #() 
NAND3_X1_567_ (
  .A1({ S5418 }),
  .A2({ S5450 }),
  .A3({ S25957[722] }),
  .ZN({ S8278 })
);
NAND3_X1 #() 
NAND3_X1_568_ (
  .A1({ S5452 }),
  .A2({ S5453 }),
  .A3({ S8203 }),
  .ZN({ S8279 })
);
NAND3_X1 #() 
NAND3_X1_569_ (
  .A1({ S8278 }),
  .A2({ S8279 }),
  .A3({ S25957[786] }),
  .ZN({ S8280 })
);
NAND2_X1 #() 
NAND2_X1_487_ (
  .A1({ S8277 }),
  .A2({ S8280 }),
  .ZN({ S8281 })
);
INV_X1 #() 
INV_X1_186_ (
  .A({ S25957[562] }),
  .ZN({ S8283 })
);
AOI21_X1 #() 
AOI21_X1_272_ (
  .A({ S8203 }),
  .B1({ S8269 }),
  .B2({ S8258 }),
  .ZN({ S8284 })
);
AOI21_X1 #() 
AOI21_X1_273_ (
  .A({ S25957[722] }),
  .B1({ S8253 }),
  .B2({ S8226 }),
  .ZN({ S8285 })
);
OAI21_X1 #() 
OAI21_X1_262_ (
  .A({ S8283 }),
  .B1({ S8284 }),
  .B2({ S8285 }),
  .ZN({ S8286 })
);
NAND3_X1 #() 
NAND3_X1_570_ (
  .A1({ S8270 }),
  .A2({ S8254 }),
  .A3({ S25957[562] }),
  .ZN({ S8287 })
);
NAND3_X1 #() 
NAND3_X1_571_ (
  .A1({ S8286 }),
  .A2({ S8281 }),
  .A3({ S8287 }),
  .ZN({ S8288 })
);
NAND2_X1 #() 
NAND2_X1_488_ (
  .A1({ S8274 }),
  .A2({ S8288 }),
  .ZN({ S25957[402] })
);
NAND3_X1 #() 
NAND3_X1_572_ (
  .A1({ S6752 }),
  .A2({ S5479 }),
  .A3({ S6748 }),
  .ZN({ S8289 })
);
NAND3_X1 #() 
NAND3_X1_573_ (
  .A1({ S6758 }),
  .A2({ S6761 }),
  .A3({ S25957[640] }),
  .ZN({ S8290 })
);
NAND2_X1 #() 
NAND2_X1_489_ (
  .A1({ S8289 }),
  .A2({ S8290 }),
  .ZN({ S8291 })
);
AOI21_X1 #() 
AOI21_X1_274_ (
  .A({ S8291 }),
  .B1({ S6826 }),
  .B2({ S6829 }),
  .ZN({ S19 })
);
NAND3_X1 #() 
NAND3_X1_574_ (
  .A1({ S6826 }),
  .A2({ S6829 }),
  .A3({ S8291 }),
  .ZN({ S20 })
);
XNOR2_X1 #() 
XNOR2_X1_16_ (
  .A({ S25957[719] }),
  .B({ S25957[815] }),
  .ZN({ S8293 })
);
NAND2_X1 #() 
NAND2_X1_490_ (
  .A1({ S6335 }),
  .A2({ S6333 }),
  .ZN({ S8294 })
);
INV_X1 #() 
INV_X1_187_ (
  .A({ S25957[517] }),
  .ZN({ S8295 })
);
AOI21_X1 #() 
AOI21_X1_275_ (
  .A({ S5464 }),
  .B1({ S6827 }),
  .B2({ S6828 }),
  .ZN({ S8296 })
);
AOI21_X1 #() 
AOI21_X1_276_ (
  .A({ S25957[641] }),
  .B1({ S6821 }),
  .B2({ S6825 }),
  .ZN({ S8297 })
);
OAI21_X1 #() 
OAI21_X1_263_ (
  .A({ S25957[514] }),
  .B1({ S8296 }),
  .B2({ S8297 }),
  .ZN({ S8298 })
);
AOI21_X1 #() 
AOI21_X1_277_ (
  .A({ S12 }),
  .B1({ S8298 }),
  .B2({ S20 }),
  .ZN({ S8299 })
);
NAND4_X1 #() 
NAND4_X1_52_ (
  .A1({ S6826 }),
  .A2({ S6829 }),
  .A3({ S6902 }),
  .A4({ S6906 }),
  .ZN({ S8300 })
);
NAND3_X1 #() 
NAND3_X1_575_ (
  .A1({ S8291 }),
  .A2({ S6902 }),
  .A3({ S6906 }),
  .ZN({ S8302 })
);
NAND2_X1 #() 
NAND2_X1_491_ (
  .A1({ S8300 }),
  .A2({ S8302 }),
  .ZN({ S8303 })
);
NAND2_X1 #() 
NAND2_X1_492_ (
  .A1({ S8298 }),
  .A2({ S12 }),
  .ZN({ S8304 })
);
NOR2_X1 #() 
NOR2_X1_98_ (
  .A1({ S8304 }),
  .A2({ S8303 }),
  .ZN({ S8305 })
);
OAI21_X1 #() 
OAI21_X1_264_ (
  .A({ S6575 }),
  .B1({ S8305 }),
  .B2({ S8299 }),
  .ZN({ S8306 })
);
AOI22_X1 #() 
AOI22_X1_43_ (
  .A1({ S6902 }),
  .A2({ S6906 }),
  .B1({ S6762 }),
  .B2({ S6754 }),
  .ZN({ S8307 })
);
NOR2_X1 #() 
NOR2_X1_99_ (
  .A1({ S8307 }),
  .A2({ S12 }),
  .ZN({ S8308 })
);
NAND2_X1 #() 
NAND2_X1_493_ (
  .A1({ S8308 }),
  .A2({ S8300 }),
  .ZN({ S8309 })
);
NAND2_X1 #() 
NAND2_X1_494_ (
  .A1({ S12 }),
  .A2({ S25957[512] }),
  .ZN({ S8310 })
);
NAND3_X1 #() 
NAND3_X1_576_ (
  .A1({ S8309 }),
  .A2({ S25957[516] }),
  .A3({ S8310 }),
  .ZN({ S8311 })
);
AOI21_X1 #() 
AOI21_X1_278_ (
  .A({ S8295 }),
  .B1({ S8306 }),
  .B2({ S8311 }),
  .ZN({ S8313 })
);
AND2_X1 #() 
AND2_X1_25_ (
  .A1({ S6906 }),
  .A2({ S6902 }),
  .ZN({ S8314 })
);
OAI21_X1 #() 
OAI21_X1_265_ (
  .A({ S25957[512] }),
  .B1({ S8296 }),
  .B2({ S8297 }),
  .ZN({ S8315 })
);
AOI21_X1 #() 
AOI21_X1_279_ (
  .A({ S8314 }),
  .B1({ S8315 }),
  .B2({ S20 }),
  .ZN({ S8316 })
);
NOR2_X1 #() 
NOR2_X1_100_ (
  .A1({ S8316 }),
  .A2({ S25957[515] }),
  .ZN({ S8317 })
);
AOI21_X1 #() 
AOI21_X1_280_ (
  .A({ S5471 }),
  .B1({ S6903 }),
  .B2({ S6905 }),
  .ZN({ S8318 })
);
AOI21_X1 #() 
AOI21_X1_281_ (
  .A({ S25957[642] }),
  .B1({ S6887 }),
  .B2({ S6901 }),
  .ZN({ S8319 })
);
OAI21_X1 #() 
OAI21_X1_266_ (
  .A({ S8291 }),
  .B1({ S8318 }),
  .B2({ S8319 }),
  .ZN({ S8320 })
);
OAI211_X1 #() 
OAI211_X1_146_ (
  .A({ S6826 }),
  .B({ S6829 }),
  .C1({ S8319 }),
  .C2({ S8318 }),
  .ZN({ S8321 })
);
NAND2_X1 #() 
NAND2_X1_495_ (
  .A1({ S8321 }),
  .A2({ S25957[515] }),
  .ZN({ S8322 })
);
INV_X1 #() 
INV_X1_188_ (
  .A({ S8322 }),
  .ZN({ S8324 })
);
AOI21_X1 #() 
AOI21_X1_282_ (
  .A({ S8317 }),
  .B1({ S8320 }),
  .B2({ S8324 }),
  .ZN({ S8325 })
);
NAND2_X1 #() 
NAND2_X1_496_ (
  .A1({ S20 }),
  .A2({ S25957[514] }),
  .ZN({ S8326 })
);
NOR2_X1 #() 
NOR2_X1_101_ (
  .A1({ S8326 }),
  .A2({ S19 }),
  .ZN({ S8327 })
);
AND3_X1 #() 
AND3_X1_21_ (
  .A1({ S25957[512] }),
  .A2({ S6902 }),
  .A3({ S6906 }),
  .ZN({ S8328 })
);
NAND2_X1 #() 
NAND2_X1_497_ (
  .A1({ S8328 }),
  .A2({ S25957[513] }),
  .ZN({ S8329 })
);
NAND2_X1 #() 
NAND2_X1_498_ (
  .A1({ S8329 }),
  .A2({ S12 }),
  .ZN({ S8330 })
);
NOR2_X1 #() 
NOR2_X1_102_ (
  .A1({ S8327 }),
  .A2({ S8330 }),
  .ZN({ S8331 })
);
AOI22_X1 #() 
AOI22_X1_44_ (
  .A1({ S6902 }),
  .A2({ S6906 }),
  .B1({ S8290 }),
  .B2({ S8289 }),
  .ZN({ S8332 })
);
NOR2_X1 #() 
NOR2_X1_103_ (
  .A1({ S8332 }),
  .A2({ S12 }),
  .ZN({ S8333 })
);
INV_X1 #() 
INV_X1_189_ (
  .A({ S8333 }),
  .ZN({ S8335 })
);
NAND3_X1 #() 
NAND3_X1_577_ (
  .A1({ S25957[515] }),
  .A2({ S6826 }),
  .A3({ S6829 }),
  .ZN({ S8336 })
);
NAND3_X1 #() 
NAND3_X1_578_ (
  .A1({ S8335 }),
  .A2({ S25957[516] }),
  .A3({ S8336 }),
  .ZN({ S8337 })
);
OAI22_X1 #() 
OAI22_X1_14_ (
  .A1({ S8325 }),
  .A2({ S25957[516] }),
  .B1({ S8331 }),
  .B2({ S8337 }),
  .ZN({ S8338 })
);
AOI21_X1 #() 
AOI21_X1_283_ (
  .A({ S8313 }),
  .B1({ S8338 }),
  .B2({ S8295 }),
  .ZN({ S8339 })
);
AOI21_X1 #() 
AOI21_X1_284_ (
  .A({ S12 }),
  .B1({ S8300 }),
  .B2({ S8320 }),
  .ZN({ S8340 })
);
AND2_X1 #() 
AND2_X1_26_ (
  .A1({ S6829 }),
  .A2({ S6826 }),
  .ZN({ S8341 })
);
NAND3_X1 #() 
NAND3_X1_579_ (
  .A1({ S6826 }),
  .A2({ S6829 }),
  .A3({ S25957[512] }),
  .ZN({ S8342 })
);
OAI21_X1 #() 
OAI21_X1_267_ (
  .A({ S25957[512] }),
  .B1({ S8318 }),
  .B2({ S8319 }),
  .ZN({ S8343 })
);
AOI22_X1 #() 
AOI22_X1_45_ (
  .A1({ S25957[514] }),
  .A2({ S8341 }),
  .B1({ S8342 }),
  .B2({ S8343 }),
  .ZN({ S8344 })
);
OAI21_X1 #() 
OAI21_X1_268_ (
  .A({ S6575 }),
  .B1({ S8344 }),
  .B2({ S25957[515] }),
  .ZN({ S8345 })
);
NAND2_X1 #() 
NAND2_X1_499_ (
  .A1({ S8321 }),
  .A2({ S8320 }),
  .ZN({ S8346 })
);
AOI21_X1 #() 
AOI21_X1_285_ (
  .A({ S25957[514] }),
  .B1({ S8315 }),
  .B2({ S20 }),
  .ZN({ S8347 })
);
OAI21_X1 #() 
OAI21_X1_269_ (
  .A({ S25957[515] }),
  .B1({ S8347 }),
  .B2({ S8346 }),
  .ZN({ S8348 })
);
NAND3_X1 #() 
NAND3_X1_580_ (
  .A1({ S8315 }),
  .A2({ S25957[514] }),
  .A3({ S20 }),
  .ZN({ S8349 })
);
NAND3_X1 #() 
NAND3_X1_581_ (
  .A1({ S25957[512] }),
  .A2({ S6902 }),
  .A3({ S6906 }),
  .ZN({ S8350 })
);
AND2_X1 #() 
AND2_X1_27_ (
  .A1({ S8350 }),
  .A2({ S12 }),
  .ZN({ S8351 })
);
NAND2_X1 #() 
NAND2_X1_500_ (
  .A1({ S8349 }),
  .A2({ S8351 }),
  .ZN({ S8352 })
);
NAND3_X1 #() 
NAND3_X1_582_ (
  .A1({ S8348 }),
  .A2({ S25957[516] }),
  .A3({ S8352 }),
  .ZN({ S8353 })
);
OAI211_X1 #() 
OAI211_X1_147_ (
  .A({ S8353 }),
  .B({ S8295 }),
  .C1({ S8340 }),
  .C2({ S8345 }),
  .ZN({ S8354 })
);
NAND2_X1 #() 
NAND2_X1_501_ (
  .A1({ S8315 }),
  .A2({ S8314 }),
  .ZN({ S8355 })
);
NAND2_X1 #() 
NAND2_X1_502_ (
  .A1({ S8355 }),
  .A2({ S8326 }),
  .ZN({ S8356 })
);
NAND2_X1 #() 
NAND2_X1_503_ (
  .A1({ S8332 }),
  .A2({ S25957[513] }),
  .ZN({ S8357 })
);
AND2_X1 #() 
AND2_X1_28_ (
  .A1({ S8302 }),
  .A2({ S12 }),
  .ZN({ S8358 })
);
NAND2_X1 #() 
NAND2_X1_504_ (
  .A1({ S8358 }),
  .A2({ S8357 }),
  .ZN({ S8359 })
);
NAND2_X1 #() 
NAND2_X1_505_ (
  .A1({ S8359 }),
  .A2({ S25957[516] }),
  .ZN({ S8360 })
);
AOI21_X1 #() 
AOI21_X1_286_ (
  .A({ S8360 }),
  .B1({ S8356 }),
  .B2({ S25957[515] }),
  .ZN({ S8361 })
);
NAND2_X1 #() 
NAND2_X1_506_ (
  .A1({ S8342 }),
  .A2({ S8314 }),
  .ZN({ S8362 })
);
AOI21_X1 #() 
AOI21_X1_287_ (
  .A({ S12 }),
  .B1({ S8362 }),
  .B2({ S8321 }),
  .ZN({ S8363 })
);
INV_X1 #() 
INV_X1_190_ (
  .A({ S8363 }),
  .ZN({ S8364 })
);
NAND2_X1 #() 
NAND2_X1_507_ (
  .A1({ S8346 }),
  .A2({ S12 }),
  .ZN({ S8365 })
);
AOI21_X1 #() 
AOI21_X1_288_ (
  .A({ S25957[516] }),
  .B1({ S8364 }),
  .B2({ S8365 }),
  .ZN({ S8366 })
);
OAI21_X1 #() 
OAI21_X1_270_ (
  .A({ S25957[517] }),
  .B1({ S8361 }),
  .B2({ S8366 }),
  .ZN({ S8367 })
);
NAND2_X1 #() 
NAND2_X1_508_ (
  .A1({ S8354 }),
  .A2({ S8367 }),
  .ZN({ S8368 })
);
NAND2_X1 #() 
NAND2_X1_509_ (
  .A1({ S8368 }),
  .A2({ S25957[518] }),
  .ZN({ S8369 })
);
OAI211_X1 #() 
OAI211_X1_148_ (
  .A({ S8369 }),
  .B({ S8294 }),
  .C1({ S25957[518] }),
  .C2({ S8339 }),
  .ZN({ S8370 })
);
NAND2_X1 #() 
NAND2_X1_510_ (
  .A1({ S25957[513] }),
  .A2({ S8350 }),
  .ZN({ S8371 })
);
NAND2_X1 #() 
NAND2_X1_511_ (
  .A1({ S8341 }),
  .A2({ S8328 }),
  .ZN({ S8372 })
);
NAND3_X1 #() 
NAND3_X1_583_ (
  .A1({ S8372 }),
  .A2({ S12 }),
  .A3({ S8371 }),
  .ZN({ S8373 })
);
OAI21_X1 #() 
OAI21_X1_271_ (
  .A({ S6575 }),
  .B1({ S8300 }),
  .B2({ S12 }),
  .ZN({ S8374 })
);
INV_X1 #() 
INV_X1_191_ (
  .A({ S8374 }),
  .ZN({ S8375 })
);
OAI21_X1 #() 
OAI21_X1_272_ (
  .A({ S8375 }),
  .B1({ S8373 }),
  .B2({ S8332 }),
  .ZN({ S8376 })
);
OAI21_X1 #() 
OAI21_X1_273_ (
  .A({ S8291 }),
  .B1({ S8296 }),
  .B2({ S8297 }),
  .ZN({ S8377 })
);
NAND3_X1 #() 
NAND3_X1_584_ (
  .A1({ S8377 }),
  .A2({ S8314 }),
  .A3({ S8342 }),
  .ZN({ S8378 })
);
AOI21_X1 #() 
AOI21_X1_289_ (
  .A({ S12 }),
  .B1({ S8349 }),
  .B2({ S8378 }),
  .ZN({ S8379 })
);
AOI22_X1 #() 
AOI22_X1_46_ (
  .A1({ S6829 }),
  .A2({ S6826 }),
  .B1({ S6902 }),
  .B2({ S6906 }),
  .ZN({ S8380 })
);
NAND2_X1 #() 
NAND2_X1_512_ (
  .A1({ S8350 }),
  .A2({ S12 }),
  .ZN({ S8381 })
);
NOR2_X1 #() 
NOR2_X1_104_ (
  .A1({ S8381 }),
  .A2({ S8380 }),
  .ZN({ S8382 })
);
OAI21_X1 #() 
OAI21_X1_274_ (
  .A({ S25957[516] }),
  .B1({ S8379 }),
  .B2({ S8382 }),
  .ZN({ S8383 })
);
AOI21_X1 #() 
AOI21_X1_290_ (
  .A({ S25957[517] }),
  .B1({ S8383 }),
  .B2({ S8376 }),
  .ZN({ S8384 })
);
NAND3_X1 #() 
NAND3_X1_585_ (
  .A1({ S8343 }),
  .A2({ S12 }),
  .A3({ S25957[513] }),
  .ZN({ S8386 })
);
OAI21_X1 #() 
OAI21_X1_275_ (
  .A({ S25957[515] }),
  .B1({ S8341 }),
  .B2({ S8307 }),
  .ZN({ S8387 })
);
NAND2_X1 #() 
NAND2_X1_513_ (
  .A1({ S8387 }),
  .A2({ S25957[516] }),
  .ZN({ S8388 })
);
INV_X1 #() 
INV_X1_192_ (
  .A({ S8388 }),
  .ZN({ S8389 })
);
NAND2_X1 #() 
NAND2_X1_514_ (
  .A1({ S8302 }),
  .A2({ S12 }),
  .ZN({ S8390 })
);
NAND2_X1 #() 
NAND2_X1_515_ (
  .A1({ S25957[513] }),
  .A2({ S12 }),
  .ZN({ S8391 })
);
NAND2_X1 #() 
NAND2_X1_516_ (
  .A1({ S8391 }),
  .A2({ S8390 }),
  .ZN({ S8392 })
);
NOR3_X1 #() 
NOR3_X1_16_ (
  .A1({ S8392 }),
  .A2({ S19 }),
  .A3({ S25957[516] }),
  .ZN({ S8393 })
);
AOI211_X1 #() 
AOI211_X1_5_ (
  .A({ S8295 }),
  .B({ S8393 }),
  .C1({ S8386 }),
  .C2({ S8389 }),
  .ZN({ S8394 })
);
NOR2_X1 #() 
NOR2_X1_105_ (
  .A1({ S8384 }),
  .A2({ S8394 }),
  .ZN({ S8395 })
);
NAND3_X1 #() 
NAND3_X1_586_ (
  .A1({ S8357 }),
  .A2({ S25957[515] }),
  .A3({ S8342 }),
  .ZN({ S8397 })
);
NAND2_X1 #() 
NAND2_X1_517_ (
  .A1({ S8356 }),
  .A2({ S12 }),
  .ZN({ S8398 })
);
AOI21_X1 #() 
AOI21_X1_291_ (
  .A({ S25957[516] }),
  .B1({ S8398 }),
  .B2({ S8397 }),
  .ZN({ S8399 })
);
OAI211_X1 #() 
OAI211_X1_149_ (
  .A({ S8320 }),
  .B({ S25957[515] }),
  .C1({ S25957[513] }),
  .C2({ S8350 }),
  .ZN({ S8400 })
);
NAND2_X1 #() 
NAND2_X1_518_ (
  .A1({ S25957[513] }),
  .A2({ S8302 }),
  .ZN({ S8401 })
);
OAI21_X1 #() 
OAI21_X1_276_ (
  .A({ S8400 }),
  .B1({ S25957[515] }),
  .B2({ S8401 }),
  .ZN({ S8402 })
);
OAI21_X1 #() 
OAI21_X1_277_ (
  .A({ S25957[517] }),
  .B1({ S8402 }),
  .B2({ S6575 }),
  .ZN({ S8403 })
);
NOR2_X1 #() 
NOR2_X1_106_ (
  .A1({ S8322 }),
  .A2({ S19 }),
  .ZN({ S8404 })
);
AOI21_X1 #() 
AOI21_X1_292_ (
  .A({ S25957[512] }),
  .B1({ S6826 }),
  .B2({ S6829 }),
  .ZN({ S8405 })
);
NOR2_X1 #() 
NOR2_X1_107_ (
  .A1({ S8405 }),
  .A2({ S25957[515] }),
  .ZN({ S8406 })
);
OAI21_X1 #() 
OAI21_X1_278_ (
  .A({ S25957[516] }),
  .B1({ S8404 }),
  .B2({ S8406 }),
  .ZN({ S8408 })
);
NAND4_X1 #() 
NAND4_X1_53_ (
  .A1({ S8314 }),
  .A2({ S6829 }),
  .A3({ S6826 }),
  .A4({ S8291 }),
  .ZN({ S8409 })
);
NOR2_X1 #() 
NOR2_X1_108_ (
  .A1({ S25957[513] }),
  .A2({ S12 }),
  .ZN({ S8410 })
);
AOI21_X1 #() 
AOI21_X1_293_ (
  .A({ S25957[516] }),
  .B1({ S8410 }),
  .B2({ S25957[512] }),
  .ZN({ S8411 })
);
NAND3_X1 #() 
NAND3_X1_587_ (
  .A1({ S8411 }),
  .A2({ S8326 }),
  .A3({ S8409 }),
  .ZN({ S8412 })
);
AND2_X1 #() 
AND2_X1_29_ (
  .A1({ S8408 }),
  .A2({ S8412 }),
  .ZN({ S8413 })
);
OAI22_X1 #() 
OAI22_X1_15_ (
  .A1({ S8413 }),
  .A2({ S25957[517] }),
  .B1({ S8399 }),
  .B2({ S8403 }),
  .ZN({ S8414 })
);
NAND2_X1 #() 
NAND2_X1_519_ (
  .A1({ S8414 }),
  .A2({ S25957[518] }),
  .ZN({ S8415 })
);
OAI211_X1 #() 
OAI211_X1_150_ (
  .A({ S25957[519] }),
  .B({ S8415 }),
  .C1({ S8395 }),
  .C2({ S25957[518] }),
  .ZN({ S8416 })
);
NAND2_X1 #() 
NAND2_X1_520_ (
  .A1({ S8370 }),
  .A2({ S8416 }),
  .ZN({ S8417 })
);
NAND2_X1 #() 
NAND2_X1_521_ (
  .A1({ S8417 }),
  .A2({ S25957[623] }),
  .ZN({ S8419 })
);
OR2_X1 #() 
OR2_X1_7_ (
  .A1({ S8417 }),
  .A2({ S25957[623] }),
  .ZN({ S8420 })
);
NAND2_X1 #() 
NAND2_X1_522_ (
  .A1({ S8420 }),
  .A2({ S8419 }),
  .ZN({ S8421 })
);
NOR2_X1 #() 
NOR2_X1_109_ (
  .A1({ S8421 }),
  .A2({ S8293 }),
  .ZN({ S8422 })
);
INV_X1 #() 
INV_X1_193_ (
  .A({ S8293 }),
  .ZN({ S25957[687] })
);
INV_X1 #() 
INV_X1_194_ (
  .A({ S8421 }),
  .ZN({ S25957[495] })
);
NOR2_X1 #() 
NOR2_X1_110_ (
  .A1({ S25957[495] }),
  .A2({ S25957[687] }),
  .ZN({ S8423 })
);
OAI21_X1 #() 
OAI21_X1_279_ (
  .A({ S7562 }),
  .B1({ S8423 }),
  .B2({ S8422 }),
  .ZN({ S8424 })
);
INV_X1 #() 
INV_X1_195_ (
  .A({ S8424 }),
  .ZN({ S8425 })
);
NOR3_X1 #() 
NOR3_X1_17_ (
  .A1({ S8423 }),
  .A2({ S8422 }),
  .A3({ S7562 }),
  .ZN({ S8426 })
);
NOR2_X1 #() 
NOR2_X1_111_ (
  .A1({ S8425 }),
  .A2({ S8426 }),
  .ZN({ S25957[399] })
);
NAND4_X1 #() 
NAND4_X1_54_ (
  .A1({ S8315 }),
  .A2({ S20 }),
  .A3({ S12 }),
  .A4({ S8314 }),
  .ZN({ S8428 })
);
NAND2_X1 #() 
NAND2_X1_523_ (
  .A1({ S8307 }),
  .A2({ S12 }),
  .ZN({ S8429 })
);
NAND2_X1 #() 
NAND2_X1_524_ (
  .A1({ S8428 }),
  .A2({ S8429 }),
  .ZN({ S8430 })
);
AOI21_X1 #() 
AOI21_X1_294_ (
  .A({ S12 }),
  .B1({ S8357 }),
  .B2({ S8350 }),
  .ZN({ S8431 })
);
OAI21_X1 #() 
OAI21_X1_280_ (
  .A({ S6575 }),
  .B1({ S8430 }),
  .B2({ S8431 }),
  .ZN({ S8432 })
);
OAI21_X1 #() 
OAI21_X1_281_ (
  .A({ S8389 }),
  .B1({ S25957[515] }),
  .B2({ S8362 }),
  .ZN({ S8433 })
);
AND3_X1 #() 
AND3_X1_22_ (
  .A1({ S8433 }),
  .A2({ S8432 }),
  .A3({ S8295 }),
  .ZN({ S8434 })
);
NAND3_X1 #() 
NAND3_X1_588_ (
  .A1({ S8307 }),
  .A2({ S6826 }),
  .A3({ S6829 }),
  .ZN({ S8435 })
);
NAND3_X1 #() 
NAND3_X1_589_ (
  .A1({ S8435 }),
  .A2({ S25957[515] }),
  .A3({ S8302 }),
  .ZN({ S8436 })
);
INV_X1 #() 
INV_X1_196_ (
  .A({ S8436 }),
  .ZN({ S8438 })
);
OAI21_X1 #() 
OAI21_X1_282_ (
  .A({ S25957[516] }),
  .B1({ S8438 }),
  .B2({ S8430 }),
  .ZN({ S8439 })
);
NAND4_X1 #() 
NAND4_X1_55_ (
  .A1({ S25957[514] }),
  .A2({ S6829 }),
  .A3({ S6826 }),
  .A4({ S8291 }),
  .ZN({ S8440 })
);
NAND2_X1 #() 
NAND2_X1_525_ (
  .A1({ S8440 }),
  .A2({ S25957[515] }),
  .ZN({ S8441 })
);
OAI21_X1 #() 
OAI21_X1_283_ (
  .A({ S8441 }),
  .B1({ S8344 }),
  .B2({ S25957[515] }),
  .ZN({ S8442 })
);
NAND2_X1 #() 
NAND2_X1_526_ (
  .A1({ S8303 }),
  .A2({ S25957[515] }),
  .ZN({ S8443 })
);
NAND3_X1 #() 
NAND3_X1_590_ (
  .A1({ S8442 }),
  .A2({ S6575 }),
  .A3({ S8443 }),
  .ZN({ S8444 })
);
NAND3_X1 #() 
NAND3_X1_591_ (
  .A1({ S8444 }),
  .A2({ S8439 }),
  .A3({ S8295 }),
  .ZN({ S8445 })
);
NAND4_X1 #() 
NAND4_X1_56_ (
  .A1({ S8341 }),
  .A2({ S8320 }),
  .A3({ S25957[515] }),
  .A4({ S8350 }),
  .ZN({ S8446 })
);
INV_X1 #() 
INV_X1_197_ (
  .A({ S8446 }),
  .ZN({ S8447 })
);
OAI21_X1 #() 
OAI21_X1_284_ (
  .A({ S25957[516] }),
  .B1({ S8326 }),
  .B2({ S25957[515] }),
  .ZN({ S8449 })
);
AOI21_X1 #() 
AOI21_X1_295_ (
  .A({ S8404 }),
  .B1({ S25957[513] }),
  .B2({ S12 }),
  .ZN({ S8450 })
);
OAI22_X1 #() 
OAI22_X1_16_ (
  .A1({ S8450 }),
  .A2({ S25957[516] }),
  .B1({ S8447 }),
  .B2({ S8449 }),
  .ZN({ S8451 })
);
OAI21_X1 #() 
OAI21_X1_285_ (
  .A({ S8445 }),
  .B1({ S8451 }),
  .B2({ S8295 }),
  .ZN({ S8452 })
);
NAND4_X1 #() 
NAND4_X1_57_ (
  .A1({ S8377 }),
  .A2({ S8342 }),
  .A3({ S25957[514] }),
  .A4({ S12 }),
  .ZN({ S8453 })
);
INV_X1 #() 
INV_X1_198_ (
  .A({ S8453 }),
  .ZN({ S8454 })
);
AOI22_X1 #() 
AOI22_X1_47_ (
  .A1({ S6652 }),
  .A2({ S6653 }),
  .B1({ S6906 }),
  .B2({ S6902 }),
  .ZN({ S8455 })
);
NAND2_X1 #() 
NAND2_X1_527_ (
  .A1({ S8455 }),
  .A2({ S25957[513] }),
  .ZN({ S8456 })
);
NAND3_X1 #() 
NAND3_X1_592_ (
  .A1({ S8405 }),
  .A2({ S12 }),
  .A3({ S8314 }),
  .ZN({ S8457 })
);
NAND2_X1 #() 
NAND2_X1_528_ (
  .A1({ S8457 }),
  .A2({ S8456 }),
  .ZN({ S8458 })
);
OAI21_X1 #() 
OAI21_X1_286_ (
  .A({ S25957[516] }),
  .B1({ S8454 }),
  .B2({ S8458 }),
  .ZN({ S8460 })
);
NAND2_X1 #() 
NAND2_X1_529_ (
  .A1({ S8307 }),
  .A2({ S25957[513] }),
  .ZN({ S8461 })
);
AOI21_X1 #() 
AOI21_X1_296_ (
  .A({ S25957[515] }),
  .B1({ S8461 }),
  .B2({ S20 }),
  .ZN({ S8462 })
);
NOR2_X1 #() 
NOR2_X1_112_ (
  .A1({ S8341 }),
  .A2({ S8302 }),
  .ZN({ S8463 })
);
OAI21_X1 #() 
OAI21_X1_287_ (
  .A({ S6575 }),
  .B1({ S8463 }),
  .B2({ S8322 }),
  .ZN({ S8464 })
);
OAI21_X1 #() 
OAI21_X1_288_ (
  .A({ S8460 }),
  .B1({ S8462 }),
  .B2({ S8464 }),
  .ZN({ S8465 })
);
OAI21_X1 #() 
OAI21_X1_289_ (
  .A({ S6416 }),
  .B1({ S8465 }),
  .B2({ S8295 }),
  .ZN({ S8466 })
);
OAI221_X1 #() 
OAI221_X1_8_ (
  .A({ S25957[519] }),
  .B1({ S8434 }),
  .B2({ S8466 }),
  .C1({ S6416 }),
  .C2({ S8452 }),
  .ZN({ S8467 })
);
NOR2_X1 #() 
NOR2_X1_113_ (
  .A1({ S25957[513] }),
  .A2({ S8350 }),
  .ZN({ S8468 })
);
NOR2_X1 #() 
NOR2_X1_114_ (
  .A1({ S8304 }),
  .A2({ S8468 }),
  .ZN({ S8469 })
);
AOI21_X1 #() 
AOI21_X1_297_ (
  .A({ S25957[514] }),
  .B1({ S6829 }),
  .B2({ S6826 }),
  .ZN({ S8471 })
);
OAI21_X1 #() 
OAI21_X1_290_ (
  .A({ S6575 }),
  .B1({ S8322 }),
  .B2({ S8471 }),
  .ZN({ S8472 })
);
OAI21_X1 #() 
OAI21_X1_291_ (
  .A({ S8381 }),
  .B1({ S8441 }),
  .B2({ S19 }),
  .ZN({ S8473 })
);
OAI221_X1 #() 
OAI221_X1_9_ (
  .A({ S25957[517] }),
  .B1({ S8469 }),
  .B2({ S8472 }),
  .C1({ S6575 }),
  .C2({ S8473 }),
  .ZN({ S8474 })
);
AND3_X1 #() 
AND3_X1_23_ (
  .A1({ S8332 }),
  .A2({ S25957[513] }),
  .A3({ S25957[515] }),
  .ZN({ S8475 })
);
OAI21_X1 #() 
OAI21_X1_292_ (
  .A({ S25957[516] }),
  .B1({ S8310 }),
  .B2({ S8300 }),
  .ZN({ S8476 })
);
NAND4_X1 #() 
NAND4_X1_58_ (
  .A1({ S6647 }),
  .A2({ S6651 }),
  .A3({ S6902 }),
  .A4({ S6906 }),
  .ZN({ S8477 })
);
OAI21_X1 #() 
OAI21_X1_293_ (
  .A({ S6575 }),
  .B1({ S8405 }),
  .B2({ S8477 }),
  .ZN({ S8478 })
);
OAI221_X1 #() 
OAI221_X1_10_ (
  .A({ S8295 }),
  .B1({ S8478 }),
  .B2({ S8475 }),
  .C1({ S8363 }),
  .C2({ S8476 }),
  .ZN({ S8479 })
);
AND2_X1 #() 
AND2_X1_30_ (
  .A1({ S8474 }),
  .A2({ S8479 }),
  .ZN({ S8480 })
);
NAND2_X1 #() 
NAND2_X1_530_ (
  .A1({ S8300 }),
  .A2({ S8291 }),
  .ZN({ S8482 })
);
AOI21_X1 #() 
AOI21_X1_298_ (
  .A({ S6575 }),
  .B1({ S8471 }),
  .B2({ S25957[515] }),
  .ZN({ S8483 })
);
OAI21_X1 #() 
OAI21_X1_294_ (
  .A({ S8483 }),
  .B1({ S25957[515] }),
  .B2({ S8482 }),
  .ZN({ S8484 })
);
OAI21_X1 #() 
OAI21_X1_295_ (
  .A({ S8436 }),
  .B1({ S8327 }),
  .B2({ S25957[515] }),
  .ZN({ S8485 })
);
OAI21_X1 #() 
OAI21_X1_296_ (
  .A({ S8484 }),
  .B1({ S8485 }),
  .B2({ S25957[516] }),
  .ZN({ S8486 })
);
NAND2_X1 #() 
NAND2_X1_531_ (
  .A1({ S8486 }),
  .A2({ S8295 }),
  .ZN({ S8487 })
);
NAND2_X1 #() 
NAND2_X1_532_ (
  .A1({ S20 }),
  .A2({ S8350 }),
  .ZN({ S8488 })
);
NOR2_X1 #() 
NOR2_X1_115_ (
  .A1({ S8488 }),
  .A2({ S12 }),
  .ZN({ S8489 })
);
NAND4_X1 #() 
NAND4_X1_59_ (
  .A1({ S8321 }),
  .A2({ S12 }),
  .A3({ S8320 }),
  .A4({ S8350 }),
  .ZN({ S8490 })
);
NAND2_X1 #() 
NAND2_X1_533_ (
  .A1({ S8490 }),
  .A2({ S25957[516] }),
  .ZN({ S8491 })
);
AOI22_X1 #() 
AOI22_X1_48_ (
  .A1({ S8314 }),
  .A2({ S25957[512] }),
  .B1({ S6826 }),
  .B2({ S6829 }),
  .ZN({ S8493 })
);
AOI21_X1 #() 
AOI21_X1_299_ (
  .A({ S8489 }),
  .B1({ S8493 }),
  .B2({ S12 }),
  .ZN({ S8494 })
);
OAI221_X1 #() 
OAI221_X1_11_ (
  .A({ S25957[517] }),
  .B1({ S8489 }),
  .B2({ S8491 }),
  .C1({ S8494 }),
  .C2({ S25957[516] }),
  .ZN({ S8495 })
);
NAND3_X1 #() 
NAND3_X1_593_ (
  .A1({ S8495 }),
  .A2({ S8487 }),
  .A3({ S25957[518] }),
  .ZN({ S8496 })
);
OAI211_X1 #() 
OAI211_X1_151_ (
  .A({ S8294 }),
  .B({ S8496 }),
  .C1({ S8480 }),
  .C2({ S25957[518] }),
  .ZN({ S8497 })
);
NAND2_X1 #() 
NAND2_X1_534_ (
  .A1({ S8467 }),
  .A2({ S8497 }),
  .ZN({ S8498 })
);
NAND2_X1 #() 
NAND2_X1_535_ (
  .A1({ S8498 }),
  .A2({ S5652 }),
  .ZN({ S8499 })
);
INV_X1 #() 
INV_X1_199_ (
  .A({ S8499 }),
  .ZN({ S8500 })
);
NAND3_X1 #() 
NAND3_X1_594_ (
  .A1({ S8467 }),
  .A2({ S8497 }),
  .A3({ S25957[718] }),
  .ZN({ S8501 })
);
INV_X1 #() 
INV_X1_200_ (
  .A({ S8501 }),
  .ZN({ S8502 })
);
NOR2_X1 #() 
NOR2_X1_116_ (
  .A1({ S8500 }),
  .A2({ S8502 }),
  .ZN({ S8504 })
);
NOR2_X1 #() 
NOR2_X1_117_ (
  .A1({ S8504 }),
  .A2({ S25957[654] }),
  .ZN({ S8505 })
);
INV_X1 #() 
INV_X1_201_ (
  .A({ S8504 }),
  .ZN({ S25957[462] })
);
NOR2_X1 #() 
NOR2_X1_118_ (
  .A1({ S25957[462] }),
  .A2({ S4862 }),
  .ZN({ S8506 })
);
NOR2_X1 #() 
NOR2_X1_119_ (
  .A1({ S8506 }),
  .A2({ S8505 }),
  .ZN({ S8507 })
);
INV_X1 #() 
INV_X1_202_ (
  .A({ S8507 }),
  .ZN({ S25957[398] })
);
NAND2_X1 #() 
NAND2_X1_536_ (
  .A1({ S3148 }),
  .A2({ S3151 }),
  .ZN({ S25957[717] })
);
XNOR2_X1 #() 
XNOR2_X1_17_ (
  .A({ S25957[717] }),
  .B({ S5736 }),
  .ZN({ S25957[685] })
);
NAND2_X1 #() 
NAND2_X1_537_ (
  .A1({ S5734 }),
  .A2({ S5729 }),
  .ZN({ S8508 })
);
NAND2_X1 #() 
NAND2_X1_538_ (
  .A1({ S8443 }),
  .A2({ S6575 }),
  .ZN({ S8509 })
);
NAND2_X1 #() 
NAND2_X1_539_ (
  .A1({ S8357 }),
  .A2({ S12 }),
  .ZN({ S8511 })
);
INV_X1 #() 
INV_X1_203_ (
  .A({ S8511 }),
  .ZN({ S8512 })
);
NOR2_X1 #() 
NOR2_X1_120_ (
  .A1({ S8482 }),
  .A2({ S12 }),
  .ZN({ S8513 })
);
AOI21_X1 #() 
AOI21_X1_300_ (
  .A({ S8513 }),
  .B1({ S8362 }),
  .B2({ S8512 }),
  .ZN({ S8514 })
);
OAI21_X1 #() 
OAI21_X1_297_ (
  .A({ S12 }),
  .B1({ S8307 }),
  .B2({ S25957[513] }),
  .ZN({ S8515 })
);
NAND2_X1 #() 
NAND2_X1_540_ (
  .A1({ S8377 }),
  .A2({ S8455 }),
  .ZN({ S8516 })
);
NAND2_X1 #() 
NAND2_X1_541_ (
  .A1({ S8516 }),
  .A2({ S8515 }),
  .ZN({ S8517 })
);
OAI22_X1 #() 
OAI22_X1_17_ (
  .A1({ S8514 }),
  .A2({ S6575 }),
  .B1({ S8509 }),
  .B2({ S8517 }),
  .ZN({ S8518 })
);
AOI21_X1 #() 
AOI21_X1_301_ (
  .A({ S25957[516] }),
  .B1({ S8436 }),
  .B2({ S8453 }),
  .ZN({ S8519 })
);
NAND2_X1 #() 
NAND2_X1_542_ (
  .A1({ S8300 }),
  .A2({ S8350 }),
  .ZN({ S8520 })
);
NAND2_X1 #() 
NAND2_X1_543_ (
  .A1({ S8321 }),
  .A2({ S8343 }),
  .ZN({ S8522 })
);
OAI21_X1 #() 
OAI21_X1_298_ (
  .A({ S25957[516] }),
  .B1({ S8522 }),
  .B2({ S25957[515] }),
  .ZN({ S8523 })
);
AOI21_X1 #() 
AOI21_X1_302_ (
  .A({ S8523 }),
  .B1({ S8520 }),
  .B2({ S25957[515] }),
  .ZN({ S8524 })
);
OAI21_X1 #() 
OAI21_X1_299_ (
  .A({ S8295 }),
  .B1({ S8524 }),
  .B2({ S8519 }),
  .ZN({ S8525 })
);
OAI21_X1 #() 
OAI21_X1_300_ (
  .A({ S8525 }),
  .B1({ S8518 }),
  .B2({ S8295 }),
  .ZN({ S8526 })
);
NAND2_X1 #() 
NAND2_X1_544_ (
  .A1({ S8526 }),
  .A2({ S25957[518] }),
  .ZN({ S8527 })
);
NAND2_X1 #() 
NAND2_X1_545_ (
  .A1({ S8406 }),
  .A2({ S8300 }),
  .ZN({ S8528 })
);
NOR2_X1 #() 
NOR2_X1_121_ (
  .A1({ S8410 }),
  .A2({ S25957[516] }),
  .ZN({ S8529 })
);
AOI22_X1 #() 
AOI22_X1_49_ (
  .A1({ S8344 }),
  .A2({ S25957[515] }),
  .B1({ S8315 }),
  .B2({ S8358 }),
  .ZN({ S8530 })
);
AOI22_X1 #() 
AOI22_X1_50_ (
  .A1({ S8530 }),
  .A2({ S25957[516] }),
  .B1({ S8528 }),
  .B2({ S8529 }),
  .ZN({ S8531 })
);
INV_X1 #() 
INV_X1_204_ (
  .A({ S8330 }),
  .ZN({ S8533 })
);
AOI21_X1 #() 
AOI21_X1_303_ (
  .A({ S12 }),
  .B1({ S8349 }),
  .B2({ S8409 }),
  .ZN({ S8534 })
);
OAI21_X1 #() 
OAI21_X1_301_ (
  .A({ S6575 }),
  .B1({ S8534 }),
  .B2({ S8533 }),
  .ZN({ S8535 })
);
NAND3_X1 #() 
NAND3_X1_595_ (
  .A1({ S8315 }),
  .A2({ S8314 }),
  .A3({ S20 }),
  .ZN({ S8536 })
);
NOR2_X1 #() 
NOR2_X1_122_ (
  .A1({ S8536 }),
  .A2({ S12 }),
  .ZN({ S8537 })
);
OAI21_X1 #() 
OAI21_X1_302_ (
  .A({ S25957[516] }),
  .B1({ S8381 }),
  .B2({ S25957[513] }),
  .ZN({ S8538 })
);
OAI211_X1 #() 
OAI211_X1_152_ (
  .A({ S8535 }),
  .B({ S8295 }),
  .C1({ S8537 }),
  .C2({ S8538 }),
  .ZN({ S8539 })
);
OAI211_X1 #() 
OAI211_X1_153_ (
  .A({ S8539 }),
  .B({ S6416 }),
  .C1({ S8295 }),
  .C2({ S8531 }),
  .ZN({ S8540 })
);
AOI21_X1 #() 
AOI21_X1_304_ (
  .A({ S8294 }),
  .B1({ S8527 }),
  .B2({ S8540 }),
  .ZN({ S8541 })
);
OAI21_X1 #() 
OAI21_X1_303_ (
  .A({ S25957[515] }),
  .B1({ S8341 }),
  .B2({ S8302 }),
  .ZN({ S8542 })
);
NOR2_X1 #() 
NOR2_X1_123_ (
  .A1({ S8316 }),
  .A2({ S8542 }),
  .ZN({ S8544 })
);
NOR2_X1 #() 
NOR2_X1_124_ (
  .A1({ S12 }),
  .A2({ S25957[512] }),
  .ZN({ S8545 })
);
NOR2_X1 #() 
NOR2_X1_125_ (
  .A1({ S8381 }),
  .A2({ S8405 }),
  .ZN({ S8546 })
);
OAI21_X1 #() 
OAI21_X1_304_ (
  .A({ S6575 }),
  .B1({ S8546 }),
  .B2({ S8545 }),
  .ZN({ S8547 })
);
NAND3_X1 #() 
NAND3_X1_596_ (
  .A1({ S8362 }),
  .A2({ S12 }),
  .A3({ S8321 }),
  .ZN({ S8548 })
);
NAND2_X1 #() 
NAND2_X1_546_ (
  .A1({ S8548 }),
  .A2({ S25957[516] }),
  .ZN({ S8549 })
);
OAI211_X1 #() 
OAI211_X1_154_ (
  .A({ S25957[517] }),
  .B({ S8547 }),
  .C1({ S8544 }),
  .C2({ S8549 }),
  .ZN({ S8550 })
);
OAI21_X1 #() 
OAI21_X1_305_ (
  .A({ S12 }),
  .B1({ S8341 }),
  .B2({ S8302 }),
  .ZN({ S8551 })
);
NAND4_X1 #() 
NAND4_X1_60_ (
  .A1({ S8321 }),
  .A2({ S25957[515] }),
  .A3({ S8320 }),
  .A4({ S8350 }),
  .ZN({ S8552 })
);
NAND2_X1 #() 
NAND2_X1_547_ (
  .A1({ S8552 }),
  .A2({ S8551 }),
  .ZN({ S8553 })
);
NAND3_X1 #() 
NAND3_X1_597_ (
  .A1({ S8553 }),
  .A2({ S6575 }),
  .A3({ S8429 }),
  .ZN({ S8555 })
);
NAND3_X1 #() 
NAND3_X1_598_ (
  .A1({ S8355 }),
  .A2({ S12 }),
  .A3({ S8461 }),
  .ZN({ S8556 })
);
NAND3_X1 #() 
NAND3_X1_599_ (
  .A1({ S8342 }),
  .A2({ S25957[515] }),
  .A3({ S8314 }),
  .ZN({ S8557 })
);
NAND3_X1 #() 
NAND3_X1_600_ (
  .A1({ S8556 }),
  .A2({ S25957[516] }),
  .A3({ S8557 }),
  .ZN({ S8558 })
);
NAND3_X1 #() 
NAND3_X1_601_ (
  .A1({ S8555 }),
  .A2({ S8558 }),
  .A3({ S8295 }),
  .ZN({ S8559 })
);
NAND3_X1 #() 
NAND3_X1_602_ (
  .A1({ S8559 }),
  .A2({ S25957[518] }),
  .A3({ S8550 }),
  .ZN({ S8560 })
);
NOR3_X1 #() 
NOR3_X1_18_ (
  .A1({ S8316 }),
  .A2({ S8468 }),
  .A3({ S12 }),
  .ZN({ S8561 })
);
NAND4_X1 #() 
NAND4_X1_61_ (
  .A1({ S8377 }),
  .A2({ S8302 }),
  .A3({ S8342 }),
  .A4({ S12 }),
  .ZN({ S8562 })
);
NAND2_X1 #() 
NAND2_X1_548_ (
  .A1({ S8562 }),
  .A2({ S25957[516] }),
  .ZN({ S8563 })
);
AOI21_X1 #() 
AOI21_X1_305_ (
  .A({ S8291 }),
  .B1({ S6647 }),
  .B2({ S6651 }),
  .ZN({ S8564 })
);
AOI22_X1 #() 
AOI22_X1_51_ (
  .A1({ S8410 }),
  .A2({ S25957[512] }),
  .B1({ S8380 }),
  .B2({ S8564 }),
  .ZN({ S8566 })
);
OAI221_X1 #() 
OAI221_X1_12_ (
  .A({ S8295 }),
  .B1({ S25957[516] }),
  .B2({ S8566 }),
  .C1({ S8561 }),
  .C2({ S8563 }),
  .ZN({ S8567 })
);
NAND2_X1 #() 
NAND2_X1_549_ (
  .A1({ S8307 }),
  .A2({ S25957[515] }),
  .ZN({ S8568 })
);
NAND3_X1 #() 
NAND3_X1_603_ (
  .A1({ S8351 }),
  .A2({ S25957[513] }),
  .A3({ S8320 }),
  .ZN({ S8569 })
);
AOI21_X1 #() 
AOI21_X1_306_ (
  .A({ S25957[516] }),
  .B1({ S8569 }),
  .B2({ S8568 }),
  .ZN({ S8570 })
);
AOI21_X1 #() 
AOI21_X1_307_ (
  .A({ S6575 }),
  .B1({ S8443 }),
  .B2({ S8551 }),
  .ZN({ S8571 })
);
OR3_X1 #() 
OR3_X1_1_ (
  .A1({ S8570 }),
  .A2({ S8571 }),
  .A3({ S8295 }),
  .ZN({ S8572 })
);
NAND3_X1 #() 
NAND3_X1_604_ (
  .A1({ S8572 }),
  .A2({ S6416 }),
  .A3({ S8567 }),
  .ZN({ S8573 })
);
AOI21_X1 #() 
AOI21_X1_308_ (
  .A({ S25957[519] }),
  .B1({ S8573 }),
  .B2({ S8560 }),
  .ZN({ S8574 })
);
NOR2_X1 #() 
NOR2_X1_126_ (
  .A1({ S8541 }),
  .A2({ S8574 }),
  .ZN({ S8575 })
);
NAND2_X1 #() 
NAND2_X1_550_ (
  .A1({ S8575 }),
  .A2({ S8508 }),
  .ZN({ S8577 })
);
INV_X1 #() 
INV_X1_205_ (
  .A({ S8508 }),
  .ZN({ S25957[621] })
);
OAI21_X1 #() 
OAI21_X1_306_ (
  .A({ S25957[621] }),
  .B1({ S8541 }),
  .B2({ S8574 }),
  .ZN({ S8578 })
);
AOI21_X1 #() 
AOI21_X1_309_ (
  .A({ S25957[685] }),
  .B1({ S8577 }),
  .B2({ S8578 }),
  .ZN({ S8579 })
);
INV_X1 #() 
INV_X1_206_ (
  .A({ S25957[685] }),
  .ZN({ S8580 })
);
NAND2_X1 #() 
NAND2_X1_551_ (
  .A1({ S8575 }),
  .A2({ S25957[621] }),
  .ZN({ S8581 })
);
OAI21_X1 #() 
OAI21_X1_307_ (
  .A({ S8508 }),
  .B1({ S8541 }),
  .B2({ S8574 }),
  .ZN({ S8582 })
);
AOI21_X1 #() 
AOI21_X1_310_ (
  .A({ S8580 }),
  .B1({ S8581 }),
  .B2({ S8582 }),
  .ZN({ S8583 })
);
OAI21_X1 #() 
OAI21_X1_308_ (
  .A({ S7605 }),
  .B1({ S8579 }),
  .B2({ S8583 }),
  .ZN({ S8584 })
);
NAND3_X1 #() 
NAND3_X1_605_ (
  .A1({ S8581 }),
  .A2({ S8582 }),
  .A3({ S8580 }),
  .ZN({ S8585 })
);
NAND3_X1 #() 
NAND3_X1_606_ (
  .A1({ S8577 }),
  .A2({ S8578 }),
  .A3({ S25957[685] }),
  .ZN({ S8587 })
);
NAND3_X1 #() 
NAND3_X1_607_ (
  .A1({ S8585 }),
  .A2({ S8587 }),
  .A3({ S25957[525] }),
  .ZN({ S8588 })
);
NAND2_X1 #() 
NAND2_X1_552_ (
  .A1({ S8584 }),
  .A2({ S8588 }),
  .ZN({ S25957[397] })
);
NAND2_X1 #() 
NAND2_X1_553_ (
  .A1({ S5835 }),
  .A2({ S5839 }),
  .ZN({ S25957[556] })
);
INV_X1 #() 
INV_X1_207_ (
  .A({ S5745 }),
  .ZN({ S25957[716] })
);
OAI211_X1 #() 
OAI211_X1_155_ (
  .A({ S25957[515] }),
  .B({ S8342 }),
  .C1({ S8377 }),
  .C2({ S25957[514] }),
  .ZN({ S8589 })
);
OAI21_X1 #() 
OAI21_X1_309_ (
  .A({ S12 }),
  .B1({ S8488 }),
  .B2({ S8380 }),
  .ZN({ S8590 })
);
NAND3_X1 #() 
NAND3_X1_608_ (
  .A1({ S8590 }),
  .A2({ S8589 }),
  .A3({ S25957[516] }),
  .ZN({ S8591 })
);
NAND2_X1 #() 
NAND2_X1_554_ (
  .A1({ S8315 }),
  .A2({ S25957[514] }),
  .ZN({ S8592 })
);
AOI21_X1 #() 
AOI21_X1_311_ (
  .A({ S25957[515] }),
  .B1({ S8378 }),
  .B2({ S8592 }),
  .ZN({ S8593 })
);
NAND2_X1 #() 
NAND2_X1_555_ (
  .A1({ S8405 }),
  .A2({ S8455 }),
  .ZN({ S8595 })
);
NAND3_X1 #() 
NAND3_X1_609_ (
  .A1({ S8595 }),
  .A2({ S8557 }),
  .A3({ S6575 }),
  .ZN({ S8596 })
);
OAI211_X1 #() 
OAI211_X1_156_ (
  .A({ S8591 }),
  .B({ S25957[517] }),
  .C1({ S8593 }),
  .C2({ S8596 }),
  .ZN({ S8597 })
);
NAND2_X1 #() 
NAND2_X1_556_ (
  .A1({ S25957[513] }),
  .A2({ S8314 }),
  .ZN({ S8598 })
);
AND2_X1 #() 
AND2_X1_31_ (
  .A1({ S8598 }),
  .A2({ S8321 }),
  .ZN({ S8599 })
);
NAND2_X1 #() 
NAND2_X1_557_ (
  .A1({ S8599 }),
  .A2({ S8308 }),
  .ZN({ S8600 })
);
NAND4_X1 #() 
NAND4_X1_62_ (
  .A1({ S8321 }),
  .A2({ S8300 }),
  .A3({ S8302 }),
  .A4({ S8343 }),
  .ZN({ S8601 })
);
NAND2_X1 #() 
NAND2_X1_558_ (
  .A1({ S8601 }),
  .A2({ S12 }),
  .ZN({ S8602 })
);
NAND3_X1 #() 
NAND3_X1_610_ (
  .A1({ S8600 }),
  .A2({ S25957[516] }),
  .A3({ S8602 }),
  .ZN({ S8603 })
);
NAND2_X1 #() 
NAND2_X1_559_ (
  .A1({ S8410 }),
  .A2({ S8343 }),
  .ZN({ S8604 })
);
NAND2_X1 #() 
NAND2_X1_560_ (
  .A1({ S8377 }),
  .A2({ S25957[514] }),
  .ZN({ S8606 })
);
AOI21_X1 #() 
AOI21_X1_312_ (
  .A({ S25957[515] }),
  .B1({ S8405 }),
  .B2({ S8314 }),
  .ZN({ S8607 })
);
AOI21_X1 #() 
AOI21_X1_313_ (
  .A({ S25957[516] }),
  .B1({ S8607 }),
  .B2({ S8606 }),
  .ZN({ S8608 })
);
NAND2_X1 #() 
NAND2_X1_561_ (
  .A1({ S8608 }),
  .A2({ S8604 }),
  .ZN({ S8609 })
);
NAND3_X1 #() 
NAND3_X1_611_ (
  .A1({ S8603 }),
  .A2({ S8295 }),
  .A3({ S8609 }),
  .ZN({ S8610 })
);
NAND3_X1 #() 
NAND3_X1_612_ (
  .A1({ S8610 }),
  .A2({ S6416 }),
  .A3({ S8597 }),
  .ZN({ S8611 })
);
NAND2_X1 #() 
NAND2_X1_562_ (
  .A1({ S8440 }),
  .A2({ S12 }),
  .ZN({ S8612 })
);
NAND3_X1 #() 
NAND3_X1_613_ (
  .A1({ S8612 }),
  .A2({ S25957[516] }),
  .A3({ S8557 }),
  .ZN({ S8613 })
);
NAND3_X1 #() 
NAND3_X1_614_ (
  .A1({ S8598 }),
  .A2({ S12 }),
  .A3({ S8291 }),
  .ZN({ S8614 })
);
NAND3_X1 #() 
NAND3_X1_615_ (
  .A1({ S8614 }),
  .A2({ S8309 }),
  .A3({ S6575 }),
  .ZN({ S8615 })
);
NAND3_X1 #() 
NAND3_X1_616_ (
  .A1({ S8615 }),
  .A2({ S25957[517] }),
  .A3({ S8613 }),
  .ZN({ S8617 })
);
OAI21_X1 #() 
OAI21_X1_310_ (
  .A({ S8528 }),
  .B1({ S8328 }),
  .B2({ S8336 }),
  .ZN({ S8618 })
);
NAND3_X1 #() 
NAND3_X1_617_ (
  .A1({ S8598 }),
  .A2({ S25957[515] }),
  .A3({ S8342 }),
  .ZN({ S8619 })
);
NAND3_X1 #() 
NAND3_X1_618_ (
  .A1({ S8300 }),
  .A2({ S12 }),
  .A3({ S8320 }),
  .ZN({ S8620 })
);
NAND3_X1 #() 
NAND3_X1_619_ (
  .A1({ S8619 }),
  .A2({ S6575 }),
  .A3({ S8620 }),
  .ZN({ S8621 })
);
OAI211_X1 #() 
OAI211_X1_157_ (
  .A({ S8295 }),
  .B({ S8621 }),
  .C1({ S8618 }),
  .C2({ S6575 }),
  .ZN({ S8622 })
);
NAND3_X1 #() 
NAND3_X1_620_ (
  .A1({ S8622 }),
  .A2({ S25957[518] }),
  .A3({ S8617 }),
  .ZN({ S8623 })
);
NAND3_X1 #() 
NAND3_X1_621_ (
  .A1({ S8611 }),
  .A2({ S8623 }),
  .A3({ S25957[519] }),
  .ZN({ S8624 })
);
AOI21_X1 #() 
AOI21_X1_314_ (
  .A({ S25957[516] }),
  .B1({ S19 }),
  .B2({ S12 }),
  .ZN({ S8625 })
);
OAI21_X1 #() 
OAI21_X1_311_ (
  .A({ S8625 }),
  .B1({ S8536 }),
  .B2({ S12 }),
  .ZN({ S8626 })
);
OAI211_X1 #() 
OAI211_X1_158_ (
  .A({ S8626 }),
  .B({ S25957[517] }),
  .C1({ S8363 }),
  .C2({ S8523 }),
  .ZN({ S8628 })
);
AND4_X1 #() 
AND4_X1_2_ (
  .A1({ S6829 }),
  .A2({ S6826 }),
  .A3({ S6902 }),
  .A4({ S6906 }),
  .ZN({ S8629 })
);
OAI21_X1 #() 
OAI21_X1_312_ (
  .A({ S12 }),
  .B1({ S8629 }),
  .B2({ S8405 }),
  .ZN({ S8630 })
);
NAND3_X1 #() 
NAND3_X1_622_ (
  .A1({ S8630 }),
  .A2({ S25957[516] }),
  .A3({ S8400 }),
  .ZN({ S8631 })
);
NAND3_X1 #() 
NAND3_X1_623_ (
  .A1({ S20 }),
  .A2({ S8343 }),
  .A3({ S25957[515] }),
  .ZN({ S8632 })
);
NAND2_X1 #() 
NAND2_X1_563_ (
  .A1({ S20 }),
  .A2({ S8314 }),
  .ZN({ S8633 })
);
NAND3_X1 #() 
NAND3_X1_624_ (
  .A1({ S8633 }),
  .A2({ S12 }),
  .A3({ S8440 }),
  .ZN({ S8634 })
);
NAND3_X1 #() 
NAND3_X1_625_ (
  .A1({ S8634 }),
  .A2({ S6575 }),
  .A3({ S8632 }),
  .ZN({ S8635 })
);
NAND3_X1 #() 
NAND3_X1_626_ (
  .A1({ S8631 }),
  .A2({ S8635 }),
  .A3({ S8295 }),
  .ZN({ S8636 })
);
NAND3_X1 #() 
NAND3_X1_627_ (
  .A1({ S8628 }),
  .A2({ S8636 }),
  .A3({ S6416 }),
  .ZN({ S8637 })
);
AOI21_X1 #() 
AOI21_X1_315_ (
  .A({ S25957[515] }),
  .B1({ S8598 }),
  .B2({ S8440 }),
  .ZN({ S8639 })
);
NAND3_X1 #() 
NAND3_X1_628_ (
  .A1({ S8329 }),
  .A2({ S12 }),
  .A3({ S8320 }),
  .ZN({ S8640 })
);
NOR2_X1 #() 
NOR2_X1_127_ (
  .A1({ S8455 }),
  .A2({ S25957[516] }),
  .ZN({ S8641 })
);
AOI21_X1 #() 
AOI21_X1_316_ (
  .A({ S25957[517] }),
  .B1({ S8640 }),
  .B2({ S8641 }),
  .ZN({ S8642 })
);
OAI21_X1 #() 
OAI21_X1_313_ (
  .A({ S8642 }),
  .B1({ S8388 }),
  .B2({ S8639 }),
  .ZN({ S8643 })
);
AOI21_X1 #() 
AOI21_X1_317_ (
  .A({ S6575 }),
  .B1({ S8314 }),
  .B2({ S141 }),
  .ZN({ S8644 })
);
AOI21_X1 #() 
AOI21_X1_318_ (
  .A({ S25957[514] }),
  .B1({ S8377 }),
  .B2({ S8342 }),
  .ZN({ S8645 })
);
OAI21_X1 #() 
OAI21_X1_314_ (
  .A({ S12 }),
  .B1({ S8645 }),
  .B2({ S8522 }),
  .ZN({ S8646 })
);
AND2_X1 #() 
AND2_X1_32_ (
  .A1({ S8350 }),
  .A2({ S25957[515] }),
  .ZN({ S8647 })
);
AOI21_X1 #() 
AOI21_X1_319_ (
  .A({ S25957[516] }),
  .B1({ S8592 }),
  .B2({ S8647 }),
  .ZN({ S8648 })
);
AOI21_X1 #() 
AOI21_X1_320_ (
  .A({ S8644 }),
  .B1({ S8646 }),
  .B2({ S8648 }),
  .ZN({ S8650 })
);
NAND2_X1 #() 
NAND2_X1_564_ (
  .A1({ S8650 }),
  .A2({ S25957[517] }),
  .ZN({ S8651 })
);
NAND3_X1 #() 
NAND3_X1_629_ (
  .A1({ S8651 }),
  .A2({ S25957[518] }),
  .A3({ S8643 }),
  .ZN({ S8652 })
);
NAND3_X1 #() 
NAND3_X1_630_ (
  .A1({ S8652 }),
  .A2({ S8294 }),
  .A3({ S8637 }),
  .ZN({ S8653 })
);
NAND3_X1 #() 
NAND3_X1_631_ (
  .A1({ S8653 }),
  .A2({ S8624 }),
  .A3({ S25957[716] }),
  .ZN({ S8654 })
);
NAND2_X1 #() 
NAND2_X1_565_ (
  .A1({ S8653 }),
  .A2({ S8624 }),
  .ZN({ S8655 })
);
NAND2_X1 #() 
NAND2_X1_566_ (
  .A1({ S8655 }),
  .A2({ S5745 }),
  .ZN({ S8656 })
);
AOI21_X1 #() 
AOI21_X1_321_ (
  .A({ S25957[556] }),
  .B1({ S8656 }),
  .B2({ S8654 }),
  .ZN({ S8657 })
);
INV_X1 #() 
INV_X1_208_ (
  .A({ S25957[556] }),
  .ZN({ S8658 })
);
AND2_X1 #() 
AND2_X1_33_ (
  .A1({ S8628 }),
  .A2({ S8636 }),
  .ZN({ S8659 })
);
AND2_X1 #() 
AND2_X1_34_ (
  .A1({ S8640 }),
  .A2({ S8641 }),
  .ZN({ S8661 })
);
NOR2_X1 #() 
NOR2_X1_128_ (
  .A1({ S8388 }),
  .A2({ S8639 }),
  .ZN({ S8662 })
);
OAI21_X1 #() 
OAI21_X1_315_ (
  .A({ S8295 }),
  .B1({ S8662 }),
  .B2({ S8661 }),
  .ZN({ S8663 })
);
OAI211_X1 #() 
OAI211_X1_159_ (
  .A({ S8663 }),
  .B({ S25957[518] }),
  .C1({ S8295 }),
  .C2({ S8650 }),
  .ZN({ S8664 })
);
OAI211_X1 #() 
OAI211_X1_160_ (
  .A({ S8664 }),
  .B({ S8294 }),
  .C1({ S25957[518] }),
  .C2({ S8659 }),
  .ZN({ S8665 })
);
NAND2_X1 #() 
NAND2_X1_567_ (
  .A1({ S8622 }),
  .A2({ S8617 }),
  .ZN({ S8666 })
);
NAND2_X1 #() 
NAND2_X1_568_ (
  .A1({ S8666 }),
  .A2({ S25957[518] }),
  .ZN({ S8667 })
);
AOI22_X1 #() 
AOI22_X1_52_ (
  .A1({ S8599 }),
  .A2({ S8308 }),
  .B1({ S8601 }),
  .B2({ S12 }),
  .ZN({ S8668 })
);
OAI21_X1 #() 
OAI21_X1_316_ (
  .A({ S8604 }),
  .B1({ S8551 }),
  .B2({ S8522 }),
  .ZN({ S8669 })
);
NAND2_X1 #() 
NAND2_X1_569_ (
  .A1({ S8669 }),
  .A2({ S6575 }),
  .ZN({ S8670 })
);
OAI211_X1 #() 
OAI211_X1_161_ (
  .A({ S8670 }),
  .B({ S8295 }),
  .C1({ S8668 }),
  .C2({ S6575 }),
  .ZN({ S8672 })
);
OAI21_X1 #() 
OAI21_X1_317_ (
  .A({ S8591 }),
  .B1({ S8593 }),
  .B2({ S8596 }),
  .ZN({ S8673 })
);
NAND2_X1 #() 
NAND2_X1_570_ (
  .A1({ S8673 }),
  .A2({ S25957[517] }),
  .ZN({ S8674 })
);
NAND3_X1 #() 
NAND3_X1_632_ (
  .A1({ S8674 }),
  .A2({ S8672 }),
  .A3({ S6416 }),
  .ZN({ S8675 })
);
NAND3_X1 #() 
NAND3_X1_633_ (
  .A1({ S8667 }),
  .A2({ S8675 }),
  .A3({ S25957[519] }),
  .ZN({ S8676 })
);
AOI21_X1 #() 
AOI21_X1_322_ (
  .A({ S5745 }),
  .B1({ S8665 }),
  .B2({ S8676 }),
  .ZN({ S8677 })
);
AOI21_X1 #() 
AOI21_X1_323_ (
  .A({ S25957[716] }),
  .B1({ S8653 }),
  .B2({ S8624 }),
  .ZN({ S8678 })
);
NOR3_X1 #() 
NOR3_X1_19_ (
  .A1({ S8677 }),
  .A2({ S8678 }),
  .A3({ S8658 }),
  .ZN({ S8679 })
);
OAI21_X1 #() 
OAI21_X1_318_ (
  .A({ S25957[524] }),
  .B1({ S8679 }),
  .B2({ S8657 }),
  .ZN({ S8680 })
);
OAI21_X1 #() 
OAI21_X1_319_ (
  .A({ S8658 }),
  .B1({ S8677 }),
  .B2({ S8678 }),
  .ZN({ S8681 })
);
NAND3_X1 #() 
NAND3_X1_634_ (
  .A1({ S8656 }),
  .A2({ S8654 }),
  .A3({ S25957[556] }),
  .ZN({ S8683 })
);
NAND3_X1 #() 
NAND3_X1_635_ (
  .A1({ S8681 }),
  .A2({ S8683 }),
  .A3({ S7575 }),
  .ZN({ S8684 })
);
NAND2_X1 #() 
NAND2_X1_571_ (
  .A1({ S8680 }),
  .A2({ S8684 }),
  .ZN({ S25957[396] })
);
NAND2_X1 #() 
NAND2_X1_572_ (
  .A1({ S789 }),
  .A2({ S790 }),
  .ZN({ S25957[811] })
);
NOR2_X1 #() 
NOR2_X1_129_ (
  .A1({ S3271 }),
  .A2({ S3259 }),
  .ZN({ S25957[715] })
);
XOR2_X1 #() 
XOR2_X1_11_ (
  .A({ S25957[715] }),
  .B({ S25957[811] }),
  .Z({ S25957[683] })
);
INV_X1 #() 
INV_X1_209_ (
  .A({ S25957[683] }),
  .ZN({ S8685 })
);
NAND2_X1 #() 
NAND2_X1_573_ (
  .A1({ S3270 }),
  .A2({ S3265 }),
  .ZN({ S8686 })
);
XNOR2_X1 #() 
XNOR2_X1_18_ (
  .A({ S8686 }),
  .B({ S25957[875] }),
  .ZN({ S25957[747] })
);
XOR2_X1 #() 
XOR2_X1_12_ (
  .A({ S5899 }),
  .B({ S25957[747] }),
  .Z({ S25957[619] })
);
INV_X1 #() 
INV_X1_210_ (
  .A({ S25957[619] }),
  .ZN({ S8688 })
);
NAND2_X1 #() 
NAND2_X1_574_ (
  .A1({ S8342 }),
  .A2({ S8343 }),
  .ZN({ S8689 })
);
NAND2_X1 #() 
NAND2_X1_575_ (
  .A1({ S8435 }),
  .A2({ S25957[515] }),
  .ZN({ S8690 })
);
OAI211_X1 #() 
OAI211_X1_162_ (
  .A({ S8690 }),
  .B({ S6575 }),
  .C1({ S8689 }),
  .C2({ S25957[515] }),
  .ZN({ S8691 })
);
NAND2_X1 #() 
NAND2_X1_576_ (
  .A1({ S8441 }),
  .A2({ S25957[516] }),
  .ZN({ S8692 })
);
OAI211_X1 #() 
OAI211_X1_163_ (
  .A({ S8691 }),
  .B({ S25957[517] }),
  .C1({ S8317 }),
  .C2({ S8692 }),
  .ZN({ S8693 })
);
OAI211_X1 #() 
OAI211_X1_164_ (
  .A({ S25957[515] }),
  .B({ S20 }),
  .C1({ S8315 }),
  .C2({ S25957[514] }),
  .ZN({ S8694 })
);
NAND3_X1 #() 
NAND3_X1_636_ (
  .A1({ S8694 }),
  .A2({ S8548 }),
  .A3({ S25957[516] }),
  .ZN({ S8695 })
);
NAND2_X1 #() 
NAND2_X1_577_ (
  .A1({ S8352 }),
  .A2({ S8568 }),
  .ZN({ S8696 })
);
OAI211_X1 #() 
OAI211_X1_165_ (
  .A({ S8295 }),
  .B({ S8695 }),
  .C1({ S8696 }),
  .C2({ S8509 }),
  .ZN({ S8697 })
);
NAND3_X1 #() 
NAND3_X1_637_ (
  .A1({ S8697 }),
  .A2({ S8693 }),
  .A3({ S6416 }),
  .ZN({ S8699 })
);
NAND4_X1 #() 
NAND4_X1_63_ (
  .A1({ S8315 }),
  .A2({ S8343 }),
  .A3({ S25957[516] }),
  .A4({ S12 }),
  .ZN({ S8700 })
);
INV_X1 #() 
INV_X1_211_ (
  .A({ S8700 }),
  .ZN({ S8701 })
);
NAND3_X1 #() 
NAND3_X1_638_ (
  .A1({ S8598 }),
  .A2({ S8321 }),
  .A3({ S8564 }),
  .ZN({ S8702 })
);
AOI21_X1 #() 
AOI21_X1_324_ (
  .A({ S25957[516] }),
  .B1({ S8702 }),
  .B2({ S8400 }),
  .ZN({ S8703 })
);
OAI21_X1 #() 
OAI21_X1_320_ (
  .A({ S8295 }),
  .B1({ S8703 }),
  .B2({ S8701 }),
  .ZN({ S8704 })
);
NAND2_X1 #() 
NAND2_X1_578_ (
  .A1({ S8436 }),
  .A2({ S25957[516] }),
  .ZN({ S8705 })
);
AOI21_X1 #() 
AOI21_X1_325_ (
  .A({ S25957[515] }),
  .B1({ S25957[513] }),
  .B2({ S8314 }),
  .ZN({ S8706 })
);
NAND2_X1 #() 
NAND2_X1_579_ (
  .A1({ S8706 }),
  .A2({ S8342 }),
  .ZN({ S8707 })
);
AOI21_X1 #() 
AOI21_X1_326_ (
  .A({ S25957[516] }),
  .B1({ S8545 }),
  .B2({ S8298 }),
  .ZN({ S8708 })
);
AOI21_X1 #() 
AOI21_X1_327_ (
  .A({ S8295 }),
  .B1({ S8707 }),
  .B2({ S8708 }),
  .ZN({ S8710 })
);
OAI21_X1 #() 
OAI21_X1_321_ (
  .A({ S8710 }),
  .B1({ S8331 }),
  .B2({ S8705 }),
  .ZN({ S8711 })
);
NAND3_X1 #() 
NAND3_X1_639_ (
  .A1({ S8711 }),
  .A2({ S8704 }),
  .A3({ S25957[518] }),
  .ZN({ S8712 })
);
NAND3_X1 #() 
NAND3_X1_640_ (
  .A1({ S8699 }),
  .A2({ S8712 }),
  .A3({ S8294 }),
  .ZN({ S8713 })
);
AOI21_X1 #() 
AOI21_X1_328_ (
  .A({ S12 }),
  .B1({ S8520 }),
  .B2({ S8342 }),
  .ZN({ S8714 })
);
NAND3_X1 #() 
NAND3_X1_641_ (
  .A1({ S25957[513] }),
  .A2({ S8314 }),
  .A3({ S12 }),
  .ZN({ S8715 })
);
AOI21_X1 #() 
AOI21_X1_329_ (
  .A({ S6575 }),
  .B1({ S8307 }),
  .B2({ S12 }),
  .ZN({ S8716 })
);
NAND2_X1 #() 
NAND2_X1_580_ (
  .A1({ S8716 }),
  .A2({ S8715 }),
  .ZN({ S8717 })
);
NAND2_X1 #() 
NAND2_X1_581_ (
  .A1({ S8300 }),
  .A2({ S25957[515] }),
  .ZN({ S8718 })
);
AOI21_X1 #() 
AOI21_X1_330_ (
  .A({ S25957[516] }),
  .B1({ S8488 }),
  .B2({ S12 }),
  .ZN({ S8719 })
);
OAI21_X1 #() 
OAI21_X1_322_ (
  .A({ S8719 }),
  .B1({ S8718 }),
  .B2({ S8316 }),
  .ZN({ S8721 })
);
OAI211_X1 #() 
OAI211_X1_166_ (
  .A({ S8721 }),
  .B({ S8295 }),
  .C1({ S8714 }),
  .C2({ S8717 }),
  .ZN({ S8722 })
);
OAI211_X1 #() 
OAI211_X1_167_ (
  .A({ S12 }),
  .B({ S8300 }),
  .C1({ S8326 }),
  .C2({ S19 }),
  .ZN({ S8723 })
);
AOI21_X1 #() 
AOI21_X1_331_ (
  .A({ S12 }),
  .B1({ S8341 }),
  .B2({ S8332 }),
  .ZN({ S8724 })
);
NAND2_X1 #() 
NAND2_X1_582_ (
  .A1({ S8536 }),
  .A2({ S8724 }),
  .ZN({ S8725 })
);
AOI21_X1 #() 
AOI21_X1_332_ (
  .A({ S6575 }),
  .B1({ S8358 }),
  .B2({ S8435 }),
  .ZN({ S8726 })
);
AOI21_X1 #() 
AOI21_X1_333_ (
  .A({ S25957[516] }),
  .B1({ S8493 }),
  .B2({ S8333 }),
  .ZN({ S8727 })
);
AOI22_X1 #() 
AOI22_X1_53_ (
  .A1({ S8727 }),
  .A2({ S8723 }),
  .B1({ S8725 }),
  .B2({ S8726 }),
  .ZN({ S8728 })
);
AOI21_X1 #() 
AOI21_X1_334_ (
  .A({ S25957[518] }),
  .B1({ S8728 }),
  .B2({ S25957[517] }),
  .ZN({ S8729 })
);
NAND2_X1 #() 
NAND2_X1_583_ (
  .A1({ S8315 }),
  .A2({ S20 }),
  .ZN({ S8730 })
);
AOI21_X1 #() 
AOI21_X1_335_ (
  .A({ S8468 }),
  .B1({ S8730 }),
  .B2({ S25957[514] }),
  .ZN({ S8732 })
);
NAND2_X1 #() 
NAND2_X1_584_ (
  .A1({ S8401 }),
  .A2({ S25957[515] }),
  .ZN({ S8733 })
);
INV_X1 #() 
INV_X1_212_ (
  .A({ S8733 }),
  .ZN({ S8734 })
);
AOI21_X1 #() 
AOI21_X1_336_ (
  .A({ S8734 }),
  .B1({ S8732 }),
  .B2({ S12 }),
  .ZN({ S8735 })
);
NAND3_X1 #() 
NAND3_X1_642_ (
  .A1({ S8641 }),
  .A2({ S20 }),
  .A3({ S8350 }),
  .ZN({ S8736 })
);
OAI211_X1 #() 
OAI211_X1_168_ (
  .A({ S8295 }),
  .B({ S8736 }),
  .C1({ S8735 }),
  .C2({ S6575 }),
  .ZN({ S8737 })
);
NAND3_X1 #() 
NAND3_X1_643_ (
  .A1({ S8357 }),
  .A2({ S12 }),
  .A3({ S8342 }),
  .ZN({ S8738 })
);
AOI21_X1 #() 
AOI21_X1_337_ (
  .A({ S6575 }),
  .B1({ S8308 }),
  .B2({ S20 }),
  .ZN({ S8739 })
);
NAND2_X1 #() 
NAND2_X1_585_ (
  .A1({ S8392 }),
  .A2({ S8315 }),
  .ZN({ S8740 })
);
NAND3_X1 #() 
NAND3_X1_644_ (
  .A1({ S8298 }),
  .A2({ S20 }),
  .A3({ S8350 }),
  .ZN({ S8741 })
);
AOI21_X1 #() 
AOI21_X1_338_ (
  .A({ S25957[516] }),
  .B1({ S8741 }),
  .B2({ S25957[515] }),
  .ZN({ S8743 })
);
AOI22_X1 #() 
AOI22_X1_54_ (
  .A1({ S8743 }),
  .A2({ S8740 }),
  .B1({ S8739 }),
  .B2({ S8738 }),
  .ZN({ S8744 })
);
AOI21_X1 #() 
AOI21_X1_339_ (
  .A({ S6416 }),
  .B1({ S8744 }),
  .B2({ S25957[517] }),
  .ZN({ S8745 })
);
AOI22_X1 #() 
AOI22_X1_55_ (
  .A1({ S8737 }),
  .A2({ S8745 }),
  .B1({ S8729 }),
  .B2({ S8722 }),
  .ZN({ S8746 })
);
OAI211_X1 #() 
OAI211_X1_169_ (
  .A({ S8688 }),
  .B({ S8713 }),
  .C1({ S8746 }),
  .C2({ S8294 }),
  .ZN({ S8747 })
);
AND3_X1 #() 
AND3_X1_24_ (
  .A1({ S8699 }),
  .A2({ S8294 }),
  .A3({ S8712 }),
  .ZN({ S8748 })
);
NAND2_X1 #() 
NAND2_X1_586_ (
  .A1({ S8728 }),
  .A2({ S25957[517] }),
  .ZN({ S8749 })
);
NAND3_X1 #() 
NAND3_X1_645_ (
  .A1({ S8749 }),
  .A2({ S6416 }),
  .A3({ S8722 }),
  .ZN({ S8750 })
);
NAND2_X1 #() 
NAND2_X1_587_ (
  .A1({ S8745 }),
  .A2({ S8737 }),
  .ZN({ S8751 })
);
AOI21_X1 #() 
AOI21_X1_340_ (
  .A({ S8294 }),
  .B1({ S8751 }),
  .B2({ S8750 }),
  .ZN({ S8752 })
);
OAI21_X1 #() 
OAI21_X1_323_ (
  .A({ S25957[619] }),
  .B1({ S8752 }),
  .B2({ S8748 }),
  .ZN({ S8754 })
);
AOI21_X1 #() 
AOI21_X1_341_ (
  .A({ S8685 }),
  .B1({ S8754 }),
  .B2({ S8747 }),
  .ZN({ S8755 })
);
OAI21_X1 #() 
OAI21_X1_324_ (
  .A({ S8688 }),
  .B1({ S8752 }),
  .B2({ S8748 }),
  .ZN({ S8756 })
);
OAI211_X1 #() 
OAI211_X1_170_ (
  .A({ S25957[619] }),
  .B({ S8713 }),
  .C1({ S8746 }),
  .C2({ S8294 }),
  .ZN({ S8757 })
);
AOI21_X1 #() 
AOI21_X1_342_ (
  .A({ S25957[683] }),
  .B1({ S8756 }),
  .B2({ S8757 }),
  .ZN({ S8758 })
);
OAI21_X1 #() 
OAI21_X1_325_ (
  .A({ S9 }),
  .B1({ S8755 }),
  .B2({ S8758 }),
  .ZN({ S8759 })
);
NAND3_X1 #() 
NAND3_X1_646_ (
  .A1({ S8756 }),
  .A2({ S25957[683] }),
  .A3({ S8757 }),
  .ZN({ S8760 })
);
NAND3_X1 #() 
NAND3_X1_647_ (
  .A1({ S8754 }),
  .A2({ S8685 }),
  .A3({ S8747 }),
  .ZN({ S8761 })
);
NAND3_X1 #() 
NAND3_X1_648_ (
  .A1({ S8760 }),
  .A2({ S8761 }),
  .A3({ S25957[523] }),
  .ZN({ S8762 })
);
NAND2_X1 #() 
NAND2_X1_588_ (
  .A1({ S8759 }),
  .A2({ S8762 }),
  .ZN({ S21 })
);
AOI21_X1 #() 
AOI21_X1_343_ (
  .A({ S25957[523] }),
  .B1({ S8760 }),
  .B2({ S8761 }),
  .ZN({ S8764 })
);
AND3_X1 #() 
AND3_X1_25_ (
  .A1({ S8761 }),
  .A2({ S8760 }),
  .A3({ S25957[523] }),
  .ZN({ S8765 })
);
NOR2_X1 #() 
NOR2_X1_130_ (
  .A1({ S8765 }),
  .A2({ S8764 }),
  .ZN({ S25957[395] })
);
NOR2_X1 #() 
NOR2_X1_131_ (
  .A1({ S6010 }),
  .A2({ S6011 }),
  .ZN({ S8766 })
);
INV_X1 #() 
INV_X1_213_ (
  .A({ S8766 }),
  .ZN({ S25957[552] })
);
NAND2_X1 #() 
NAND2_X1_589_ (
  .A1({ S867 }),
  .A2({ S868 }),
  .ZN({ S25957[840] })
);
XOR2_X1 #() 
XOR2_X1_13_ (
  .A({ S25957[744] }),
  .B({ S25957[840] }),
  .Z({ S25957[712] })
);
AND2_X1 #() 
AND2_X1_35_ (
  .A1({ S8428 }),
  .A2({ S8456 }),
  .ZN({ S8767 })
);
NAND4_X1 #() 
NAND4_X1_64_ (
  .A1({ S20 }),
  .A2({ S8343 }),
  .A3({ S12 }),
  .A4({ S8302 }),
  .ZN({ S8768 })
);
AOI21_X1 #() 
AOI21_X1_344_ (
  .A({ S25957[517] }),
  .B1({ S8708 }),
  .B2({ S8768 }),
  .ZN({ S8769 })
);
OAI21_X1 #() 
OAI21_X1_326_ (
  .A({ S8769 }),
  .B1({ S8767 }),
  .B2({ S6575 }),
  .ZN({ S8771 })
);
NAND2_X1 #() 
NAND2_X1_590_ (
  .A1({ S20 }),
  .A2({ S8343 }),
  .ZN({ S8772 })
);
NAND2_X1 #() 
NAND2_X1_591_ (
  .A1({ S8598 }),
  .A2({ S12 }),
  .ZN({ S8773 })
);
OAI211_X1 #() 
OAI211_X1_171_ (
  .A({ S25957[516] }),
  .B({ S8441 }),
  .C1({ S8773 }),
  .C2({ S8772 }),
  .ZN({ S8774 })
);
NAND4_X1 #() 
NAND4_X1_65_ (
  .A1({ S8612 }),
  .A2({ S8595 }),
  .A3({ S8557 }),
  .A4({ S6575 }),
  .ZN({ S8775 })
);
NAND3_X1 #() 
NAND3_X1_649_ (
  .A1({ S8774 }),
  .A2({ S25957[517] }),
  .A3({ S8775 }),
  .ZN({ S8776 })
);
NAND3_X1 #() 
NAND3_X1_650_ (
  .A1({ S8771 }),
  .A2({ S8776 }),
  .A3({ S6416 }),
  .ZN({ S8777 })
);
NAND4_X1 #() 
NAND4_X1_66_ (
  .A1({ S8298 }),
  .A2({ S8350 }),
  .A3({ S12 }),
  .A4({ S20 }),
  .ZN({ S8778 })
);
OAI211_X1 #() 
OAI211_X1_172_ (
  .A({ S25957[516] }),
  .B({ S8778 }),
  .C1({ S8316 }),
  .C2({ S12 }),
  .ZN({ S8779 })
);
AOI21_X1 #() 
AOI21_X1_345_ (
  .A({ S25957[517] }),
  .B1({ S8553 }),
  .B2({ S6575 }),
  .ZN({ S8780 })
);
NAND3_X1 #() 
NAND3_X1_651_ (
  .A1({ S8373 }),
  .A2({ S6575 }),
  .A3({ S8400 }),
  .ZN({ S8782 })
);
NAND2_X1 #() 
NAND2_X1_592_ (
  .A1({ S8634 }),
  .A2({ S8516 }),
  .ZN({ S8783 })
);
AOI21_X1 #() 
AOI21_X1_346_ (
  .A({ S8295 }),
  .B1({ S8783 }),
  .B2({ S25957[516] }),
  .ZN({ S8784 })
);
AOI22_X1 #() 
AOI22_X1_56_ (
  .A1({ S8784 }),
  .A2({ S8782 }),
  .B1({ S8780 }),
  .B2({ S8779 }),
  .ZN({ S8785 })
);
OAI211_X1 #() 
OAI211_X1_173_ (
  .A({ S25957[519] }),
  .B({ S8777 }),
  .C1({ S8785 }),
  .C2({ S6416 }),
  .ZN({ S8786 })
);
NAND3_X1 #() 
NAND3_X1_652_ (
  .A1({ S8377 }),
  .A2({ S25957[514] }),
  .A3({ S8342 }),
  .ZN({ S8787 })
);
NAND3_X1 #() 
NAND3_X1_653_ (
  .A1({ S8787 }),
  .A2({ S25957[515] }),
  .A3({ S8355 }),
  .ZN({ S8788 })
);
AOI21_X1 #() 
AOI21_X1_347_ (
  .A({ S6575 }),
  .B1({ S8482 }),
  .B2({ S12 }),
  .ZN({ S8789 })
);
NAND2_X1 #() 
NAND2_X1_593_ (
  .A1({ S8788 }),
  .A2({ S8789 }),
  .ZN({ S8790 })
);
NOR2_X1 #() 
NOR2_X1_132_ (
  .A1({ S8478 }),
  .A2({ S8475 }),
  .ZN({ S8791 })
);
AOI21_X1 #() 
AOI21_X1_348_ (
  .A({ S8295 }),
  .B1({ S8791 }),
  .B2({ S8390 }),
  .ZN({ S8793 })
);
NAND3_X1 #() 
NAND3_X1_654_ (
  .A1({ S8552 }),
  .A2({ S6575 }),
  .A3({ S8515 }),
  .ZN({ S8794 })
);
OAI211_X1 #() 
OAI211_X1_174_ (
  .A({ S25957[516] }),
  .B({ S8321 }),
  .C1({ S8706 }),
  .C2({ S25957[512] }),
  .ZN({ S8795 })
);
NAND2_X1 #() 
NAND2_X1_594_ (
  .A1({ S8795 }),
  .A2({ S8794 }),
  .ZN({ S8796 })
);
AOI22_X1 #() 
AOI22_X1_57_ (
  .A1({ S8793 }),
  .A2({ S8790 }),
  .B1({ S8796 }),
  .B2({ S8295 }),
  .ZN({ S8797 })
);
NAND2_X1 #() 
NAND2_X1_595_ (
  .A1({ S8629 }),
  .A2({ S12 }),
  .ZN({ S8798 })
);
NAND3_X1 #() 
NAND3_X1_655_ (
  .A1({ S8453 }),
  .A2({ S25957[516] }),
  .A3({ S8798 }),
  .ZN({ S8799 })
);
NAND4_X1 #() 
NAND4_X1_67_ (
  .A1({ S8377 }),
  .A2({ S8350 }),
  .A3({ S8342 }),
  .A4({ S25957[515] }),
  .ZN({ S8800 })
);
OAI211_X1 #() 
OAI211_X1_175_ (
  .A({ S8341 }),
  .B({ S12 }),
  .C1({ S8328 }),
  .C2({ S8332 }),
  .ZN({ S8801 })
);
NAND3_X1 #() 
NAND3_X1_656_ (
  .A1({ S8800 }),
  .A2({ S8801 }),
  .A3({ S6575 }),
  .ZN({ S8802 })
);
OAI211_X1 #() 
OAI211_X1_176_ (
  .A({ S8295 }),
  .B({ S8802 }),
  .C1({ S8799 }),
  .C2({ S8714 }),
  .ZN({ S8804 })
);
OAI211_X1 #() 
OAI211_X1_177_ (
  .A({ S8632 }),
  .B({ S25957[516] }),
  .C1({ S8405 }),
  .C2({ S8381 }),
  .ZN({ S8805 })
);
NAND3_X1 #() 
NAND3_X1_657_ (
  .A1({ S8562 }),
  .A2({ S6575 }),
  .A3({ S8446 }),
  .ZN({ S8806 })
);
NAND3_X1 #() 
NAND3_X1_658_ (
  .A1({ S8806 }),
  .A2({ S25957[517] }),
  .A3({ S8805 }),
  .ZN({ S8807 })
);
NAND3_X1 #() 
NAND3_X1_659_ (
  .A1({ S8804 }),
  .A2({ S6416 }),
  .A3({ S8807 }),
  .ZN({ S8808 })
);
OAI211_X1 #() 
OAI211_X1_178_ (
  .A({ S8808 }),
  .B({ S8294 }),
  .C1({ S8797 }),
  .C2({ S6416 }),
  .ZN({ S8809 })
);
AOI21_X1 #() 
AOI21_X1_349_ (
  .A({ S25957[712] }),
  .B1({ S8786 }),
  .B2({ S8809 }),
  .ZN({ S8810 })
);
INV_X1 #() 
INV_X1_214_ (
  .A({ S25957[712] }),
  .ZN({ S8811 })
);
NAND2_X1 #() 
NAND2_X1_596_ (
  .A1({ S8793 }),
  .A2({ S8790 }),
  .ZN({ S8812 })
);
NAND2_X1 #() 
NAND2_X1_597_ (
  .A1({ S8796 }),
  .A2({ S8295 }),
  .ZN({ S8813 })
);
NAND3_X1 #() 
NAND3_X1_660_ (
  .A1({ S8812 }),
  .A2({ S25957[518] }),
  .A3({ S8813 }),
  .ZN({ S8815 })
);
NAND2_X1 #() 
NAND2_X1_598_ (
  .A1({ S8804 }),
  .A2({ S8807 }),
  .ZN({ S8816 })
);
NAND2_X1 #() 
NAND2_X1_599_ (
  .A1({ S8816 }),
  .A2({ S6416 }),
  .ZN({ S8817 })
);
NAND3_X1 #() 
NAND3_X1_661_ (
  .A1({ S8817 }),
  .A2({ S8815 }),
  .A3({ S8294 }),
  .ZN({ S8818 })
);
NAND2_X1 #() 
NAND2_X1_600_ (
  .A1({ S8780 }),
  .A2({ S8779 }),
  .ZN({ S8819 })
);
NAND2_X1 #() 
NAND2_X1_601_ (
  .A1({ S8783 }),
  .A2({ S25957[516] }),
  .ZN({ S8820 })
);
NAND3_X1 #() 
NAND3_X1_662_ (
  .A1({ S8820 }),
  .A2({ S25957[517] }),
  .A3({ S8782 }),
  .ZN({ S8821 })
);
NAND3_X1 #() 
NAND3_X1_663_ (
  .A1({ S8821 }),
  .A2({ S8819 }),
  .A3({ S25957[518] }),
  .ZN({ S8822 })
);
NAND3_X1 #() 
NAND3_X1_664_ (
  .A1({ S8428 }),
  .A2({ S25957[516] }),
  .A3({ S8456 }),
  .ZN({ S8823 })
);
NAND2_X1 #() 
NAND2_X1_602_ (
  .A1({ S8545 }),
  .A2({ S8298 }),
  .ZN({ S8824 })
);
NAND2_X1 #() 
NAND2_X1_603_ (
  .A1({ S8824 }),
  .A2({ S8768 }),
  .ZN({ S8826 })
);
NAND2_X1 #() 
NAND2_X1_604_ (
  .A1({ S8826 }),
  .A2({ S6575 }),
  .ZN({ S8827 })
);
NAND3_X1 #() 
NAND3_X1_665_ (
  .A1({ S8827 }),
  .A2({ S8823 }),
  .A3({ S8295 }),
  .ZN({ S8828 })
);
NAND2_X1 #() 
NAND2_X1_605_ (
  .A1({ S8774 }),
  .A2({ S8775 }),
  .ZN({ S8829 })
);
NAND2_X1 #() 
NAND2_X1_606_ (
  .A1({ S8829 }),
  .A2({ S25957[517] }),
  .ZN({ S8830 })
);
NAND3_X1 #() 
NAND3_X1_666_ (
  .A1({ S8830 }),
  .A2({ S6416 }),
  .A3({ S8828 }),
  .ZN({ S8831 })
);
NAND3_X1 #() 
NAND3_X1_667_ (
  .A1({ S8822 }),
  .A2({ S8831 }),
  .A3({ S25957[519] }),
  .ZN({ S8832 })
);
AOI21_X1 #() 
AOI21_X1_350_ (
  .A({ S8811 }),
  .B1({ S8818 }),
  .B2({ S8832 }),
  .ZN({ S8833 })
);
OAI21_X1 #() 
OAI21_X1_327_ (
  .A({ S25957[552] }),
  .B1({ S8833 }),
  .B2({ S8810 }),
  .ZN({ S8834 })
);
NAND3_X1 #() 
NAND3_X1_668_ (
  .A1({ S8818 }),
  .A2({ S8832 }),
  .A3({ S8811 }),
  .ZN({ S8835 })
);
NAND3_X1 #() 
NAND3_X1_669_ (
  .A1({ S8786 }),
  .A2({ S8809 }),
  .A3({ S25957[712] }),
  .ZN({ S8837 })
);
NAND3_X1 #() 
NAND3_X1_670_ (
  .A1({ S8835 }),
  .A2({ S8837 }),
  .A3({ S8766 }),
  .ZN({ S8838 })
);
NAND3_X1 #() 
NAND3_X1_671_ (
  .A1({ S8834 }),
  .A2({ S25957[520] }),
  .A3({ S8838 }),
  .ZN({ S8839 })
);
OAI21_X1 #() 
OAI21_X1_328_ (
  .A({ S8766 }),
  .B1({ S8833 }),
  .B2({ S8810 }),
  .ZN({ S8840 })
);
NAND3_X1 #() 
NAND3_X1_672_ (
  .A1({ S8835 }),
  .A2({ S8837 }),
  .A3({ S25957[552] }),
  .ZN({ S8841 })
);
NAND3_X1 #() 
NAND3_X1_673_ (
  .A1({ S8840 }),
  .A2({ S7576 }),
  .A3({ S8841 }),
  .ZN({ S8842 })
);
NAND2_X1 #() 
NAND2_X1_607_ (
  .A1({ S8839 }),
  .A2({ S8842 }),
  .ZN({ S25957[392] })
);
NOR2_X1 #() 
NOR2_X1_133_ (
  .A1({ S3404 }),
  .A2({ S3405 }),
  .ZN({ S25957[713] })
);
NAND2_X1 #() 
NAND2_X1_608_ (
  .A1({ S6090 }),
  .A2({ S6054 }),
  .ZN({ S25957[617] })
);
AND2_X1 #() 
AND2_X1_36_ (
  .A1({ S25957[617] }),
  .A2({ S25957[713] }),
  .ZN({ S8843 })
);
NOR2_X1 #() 
NOR2_X1_134_ (
  .A1({ S25957[617] }),
  .A2({ S25957[713] }),
  .ZN({ S8845 })
);
NOR2_X1 #() 
NOR2_X1_135_ (
  .A1({ S8843 }),
  .A2({ S8845 }),
  .ZN({ S25957[585] })
);
NAND2_X1 #() 
NAND2_X1_609_ (
  .A1({ S8689 }),
  .A2({ S8321 }),
  .ZN({ S8846 })
);
AOI21_X1 #() 
AOI21_X1_351_ (
  .A({ S25957[516] }),
  .B1({ S8846 }),
  .B2({ S12 }),
  .ZN({ S8847 })
);
NAND4_X1 #() 
NAND4_X1_68_ (
  .A1({ S8320 }),
  .A2({ S25957[513] }),
  .A3({ S8350 }),
  .A4({ S25957[515] }),
  .ZN({ S8848 })
);
AOI21_X1 #() 
AOI21_X1_352_ (
  .A({ S6575 }),
  .B1({ S8614 }),
  .B2({ S8848 }),
  .ZN({ S8849 })
);
OAI21_X1 #() 
OAI21_X1_329_ (
  .A({ S25957[517] }),
  .B1({ S8847 }),
  .B2({ S8849 }),
  .ZN({ S8850 })
);
AND3_X1 #() 
AND3_X1_26_ (
  .A1({ S8598 }),
  .A2({ S8321 }),
  .A3({ S8564 }),
  .ZN({ S8851 })
);
NAND4_X1 #() 
NAND4_X1_69_ (
  .A1({ S8716 }),
  .A2({ S8715 }),
  .A3({ S8568 }),
  .A4({ S8336 }),
  .ZN({ S8852 })
);
OAI211_X1 #() 
OAI211_X1_179_ (
  .A({ S8852 }),
  .B({ S8295 }),
  .C1({ S8851 }),
  .C2({ S8374 }),
  .ZN({ S8853 })
);
NAND3_X1 #() 
NAND3_X1_674_ (
  .A1({ S8850 }),
  .A2({ S6416 }),
  .A3({ S8853 }),
  .ZN({ S8855 })
);
NAND3_X1 #() 
NAND3_X1_675_ (
  .A1({ S8377 }),
  .A2({ S8350 }),
  .A3({ S8320 }),
  .ZN({ S8856 })
);
NAND2_X1 #() 
NAND2_X1_610_ (
  .A1({ S8529 }),
  .A2({ S8856 }),
  .ZN({ S8857 })
);
NAND3_X1 #() 
NAND3_X1_676_ (
  .A1({ S8372 }),
  .A2({ S8308 }),
  .A3({ S8371 }),
  .ZN({ S8858 })
);
AOI21_X1 #() 
AOI21_X1_353_ (
  .A({ S6575 }),
  .B1({ S8351 }),
  .B2({ S8440 }),
  .ZN({ S8859 })
);
NAND2_X1 #() 
NAND2_X1_611_ (
  .A1({ S8859 }),
  .A2({ S8858 }),
  .ZN({ S8860 })
);
NAND3_X1 #() 
NAND3_X1_677_ (
  .A1({ S8860 }),
  .A2({ S25957[517] }),
  .A3({ S8857 }),
  .ZN({ S8861 })
);
NAND2_X1 #() 
NAND2_X1_612_ (
  .A1({ S8392 }),
  .A2({ S8461 }),
  .ZN({ S8862 })
);
AND3_X1 #() 
AND3_X1_27_ (
  .A1({ S8788 }),
  .A2({ S25957[516] }),
  .A3({ S8862 }),
  .ZN({ S8863 })
);
NAND3_X1 #() 
NAND3_X1_678_ (
  .A1({ S8377 }),
  .A2({ S8342 }),
  .A3({ S8455 }),
  .ZN({ S8864 })
);
NAND3_X1 #() 
NAND3_X1_679_ (
  .A1({ S8864 }),
  .A2({ S8490 }),
  .A3({ S6575 }),
  .ZN({ S8866 })
);
NAND2_X1 #() 
NAND2_X1_613_ (
  .A1({ S8866 }),
  .A2({ S8295 }),
  .ZN({ S8867 })
);
OAI211_X1 #() 
OAI211_X1_180_ (
  .A({ S8861 }),
  .B({ S25957[518] }),
  .C1({ S8863 }),
  .C2({ S8867 }),
  .ZN({ S8868 })
);
NAND3_X1 #() 
NAND3_X1_680_ (
  .A1({ S8868 }),
  .A2({ S8855 }),
  .A3({ S8294 }),
  .ZN({ S8869 })
);
NAND2_X1 #() 
NAND2_X1_614_ (
  .A1({ S8332 }),
  .A2({ S12 }),
  .ZN({ S8870 })
);
NAND2_X1 #() 
NAND2_X1_615_ (
  .A1({ S8333 }),
  .A2({ S8315 }),
  .ZN({ S8871 })
);
NAND4_X1 #() 
NAND4_X1_70_ (
  .A1({ S8428 }),
  .A2({ S8871 }),
  .A3({ S6575 }),
  .A4({ S8870 }),
  .ZN({ S8872 })
);
NAND3_X1 #() 
NAND3_X1_681_ (
  .A1({ S8298 }),
  .A2({ S12 }),
  .A3({ S8291 }),
  .ZN({ S8873 })
);
OAI211_X1 #() 
OAI211_X1_181_ (
  .A({ S25957[516] }),
  .B({ S8873 }),
  .C1({ S8316 }),
  .C2({ S8542 }),
  .ZN({ S8874 })
);
NAND3_X1 #() 
NAND3_X1_682_ (
  .A1({ S8874 }),
  .A2({ S8872 }),
  .A3({ S8295 }),
  .ZN({ S8875 })
);
OAI211_X1 #() 
OAI211_X1_182_ (
  .A({ S8733 }),
  .B({ S25957[516] }),
  .C1({ S8346 }),
  .C2({ S25957[515] }),
  .ZN({ S8877 })
);
NAND3_X1 #() 
NAND3_X1_683_ (
  .A1({ S8788 }),
  .A2({ S6575 }),
  .A3({ S8511 }),
  .ZN({ S8878 })
);
NAND3_X1 #() 
NAND3_X1_684_ (
  .A1({ S8878 }),
  .A2({ S25957[517] }),
  .A3({ S8877 }),
  .ZN({ S8879 })
);
NAND3_X1 #() 
NAND3_X1_685_ (
  .A1({ S8879 }),
  .A2({ S25957[518] }),
  .A3({ S8875 }),
  .ZN({ S8880 })
);
OAI21_X1 #() 
OAI21_X1_330_ (
  .A({ S8647 }),
  .B1({ S8326 }),
  .B2({ S19 }),
  .ZN({ S8881 })
);
AOI21_X1 #() 
AOI21_X1_354_ (
  .A({ S6575 }),
  .B1({ S8881 }),
  .B2({ S8359 }),
  .ZN({ S8882 })
);
INV_X1 #() 
INV_X1_215_ (
  .A({ S8477 }),
  .ZN({ S8883 })
);
AOI21_X1 #() 
AOI21_X1_355_ (
  .A({ S25957[516] }),
  .B1({ S8883 }),
  .B2({ S8377 }),
  .ZN({ S8884 })
);
NAND3_X1 #() 
NAND3_X1_686_ (
  .A1({ S8298 }),
  .A2({ S12 }),
  .A3({ S20 }),
  .ZN({ S8885 })
);
AND2_X1 #() 
AND2_X1_37_ (
  .A1({ S8884 }),
  .A2({ S8885 }),
  .ZN({ S8886 })
);
OAI21_X1 #() 
OAI21_X1_331_ (
  .A({ S25957[517] }),
  .B1({ S8882 }),
  .B2({ S8886 }),
  .ZN({ S8888 })
);
AOI21_X1 #() 
AOI21_X1_356_ (
  .A({ S12 }),
  .B1({ S8378 }),
  .B2({ S8592 }),
  .ZN({ S8889 })
);
OAI21_X1 #() 
OAI21_X1_332_ (
  .A({ S6575 }),
  .B1({ S8551 }),
  .B2({ S8522 }),
  .ZN({ S8890 })
);
OAI211_X1 #() 
OAI211_X1_183_ (
  .A({ S8321 }),
  .B({ S12 }),
  .C1({ S8341 }),
  .C2({ S8302 }),
  .ZN({ S8891 })
);
AOI21_X1 #() 
AOI21_X1_357_ (
  .A({ S25957[517] }),
  .B1({ S8483 }),
  .B2({ S8891 }),
  .ZN({ S8892 })
);
OAI21_X1 #() 
OAI21_X1_333_ (
  .A({ S8892 }),
  .B1({ S8889 }),
  .B2({ S8890 }),
  .ZN({ S8893 })
);
NAND3_X1 #() 
NAND3_X1_687_ (
  .A1({ S8888 }),
  .A2({ S6416 }),
  .A3({ S8893 }),
  .ZN({ S8894 })
);
NAND3_X1 #() 
NAND3_X1_688_ (
  .A1({ S8880 }),
  .A2({ S8894 }),
  .A3({ S25957[519] }),
  .ZN({ S8895 })
);
NAND3_X1 #() 
NAND3_X1_689_ (
  .A1({ S8895 }),
  .A2({ S8869 }),
  .A3({ S25957[617] }),
  .ZN({ S8896 })
);
INV_X1 #() 
INV_X1_216_ (
  .A({ S25957[617] }),
  .ZN({ S8897 })
);
AOI21_X1 #() 
AOI21_X1_358_ (
  .A({ S8295 }),
  .B1({ S8859 }),
  .B2({ S8858 }),
  .ZN({ S8899 })
);
NAND3_X1 #() 
NAND3_X1_690_ (
  .A1({ S8788 }),
  .A2({ S25957[516] }),
  .A3({ S8862 }),
  .ZN({ S8900 })
);
AND2_X1 #() 
AND2_X1_38_ (
  .A1({ S8866 }),
  .A2({ S8295 }),
  .ZN({ S8901 })
);
AOI22_X1 #() 
AOI22_X1_58_ (
  .A1({ S8901 }),
  .A2({ S8900 }),
  .B1({ S8899 }),
  .B2({ S8857 }),
  .ZN({ S8902 })
);
OAI21_X1 #() 
OAI21_X1_334_ (
  .A({ S8852 }),
  .B1({ S8851 }),
  .B2({ S8374 }),
  .ZN({ S8903 })
);
NAND2_X1 #() 
NAND2_X1_616_ (
  .A1({ S8903 }),
  .A2({ S8295 }),
  .ZN({ S8904 })
);
NAND2_X1 #() 
NAND2_X1_617_ (
  .A1({ S8614 }),
  .A2({ S8848 }),
  .ZN({ S8905 })
);
NAND2_X1 #() 
NAND2_X1_618_ (
  .A1({ S8905 }),
  .A2({ S25957[516] }),
  .ZN({ S8906 })
);
NAND3_X1 #() 
NAND3_X1_691_ (
  .A1({ S8906 }),
  .A2({ S25957[517] }),
  .A3({ S8345 }),
  .ZN({ S8907 })
);
NAND3_X1 #() 
NAND3_X1_692_ (
  .A1({ S8907 }),
  .A2({ S8904 }),
  .A3({ S6416 }),
  .ZN({ S8908 })
);
OAI211_X1 #() 
OAI211_X1_184_ (
  .A({ S8908 }),
  .B({ S8294 }),
  .C1({ S8902 }),
  .C2({ S6416 }),
  .ZN({ S8910 })
);
OAI211_X1 #() 
OAI211_X1_185_ (
  .A({ S8733 }),
  .B({ S25957[517] }),
  .C1({ S8346 }),
  .C2({ S25957[515] }),
  .ZN({ S8911 })
);
NAND2_X1 #() 
NAND2_X1_619_ (
  .A1({ S8873 }),
  .A2({ S8295 }),
  .ZN({ S8912 })
);
OAI21_X1 #() 
OAI21_X1_335_ (
  .A({ S8911 }),
  .B1({ S8544 }),
  .B2({ S8912 }),
  .ZN({ S8913 })
);
NAND2_X1 #() 
NAND2_X1_620_ (
  .A1({ S8913 }),
  .A2({ S25957[516] }),
  .ZN({ S8914 })
);
NAND3_X1 #() 
NAND3_X1_693_ (
  .A1({ S6499 }),
  .A2({ S6504 }),
  .A3({ S5494 }),
  .ZN({ S8915 })
);
NAND2_X1 #() 
NAND2_X1_621_ (
  .A1({ S6499 }),
  .A2({ S6504 }),
  .ZN({ S25957[549] })
);
NAND2_X1 #() 
NAND2_X1_622_ (
  .A1({ S25957[549] }),
  .A2({ S25957[645] }),
  .ZN({ S8916 })
);
AOI22_X1 #() 
AOI22_X1_59_ (
  .A1({ S8916 }),
  .A2({ S8915 }),
  .B1({ S8332 }),
  .B2({ S12 }),
  .ZN({ S8917 })
);
AND3_X1 #() 
AND3_X1_28_ (
  .A1({ S8428 }),
  .A2({ S8871 }),
  .A3({ S8917 }),
  .ZN({ S8918 })
);
OAI21_X1 #() 
OAI21_X1_336_ (
  .A({ S8329 }),
  .B1({ S8326 }),
  .B2({ S19 }),
  .ZN({ S8920 })
);
OAI211_X1 #() 
OAI211_X1_186_ (
  .A({ S25957[517] }),
  .B({ S8310 }),
  .C1({ S8380 }),
  .C2({ S25957[515] }),
  .ZN({ S8921 })
);
AOI21_X1 #() 
AOI21_X1_359_ (
  .A({ S8921 }),
  .B1({ S8920 }),
  .B2({ S25957[515] }),
  .ZN({ S8922 })
);
OAI21_X1 #() 
OAI21_X1_337_ (
  .A({ S6575 }),
  .B1({ S8922 }),
  .B2({ S8918 }),
  .ZN({ S8923 })
);
NAND3_X1 #() 
NAND3_X1_694_ (
  .A1({ S8914 }),
  .A2({ S8923 }),
  .A3({ S25957[518] }),
  .ZN({ S8924 })
);
AOI22_X1 #() 
AOI22_X1_60_ (
  .A1({ S8349 }),
  .A2({ S8647 }),
  .B1({ S8357 }),
  .B2({ S8358 }),
  .ZN({ S8925 })
);
AOI21_X1 #() 
AOI21_X1_360_ (
  .A({ S8295 }),
  .B1({ S8884 }),
  .B2({ S8885 }),
  .ZN({ S8926 })
);
OAI21_X1 #() 
OAI21_X1_338_ (
  .A({ S8926 }),
  .B1({ S8925 }),
  .B2({ S6575 }),
  .ZN({ S8927 })
);
AOI22_X1 #() 
AOI22_X1_61_ (
  .A1({ S8348 }),
  .A2({ S8608 }),
  .B1({ S8483 }),
  .B2({ S8891 }),
  .ZN({ S8928 })
);
OAI211_X1 #() 
OAI211_X1_187_ (
  .A({ S6416 }),
  .B({ S8927 }),
  .C1({ S8928 }),
  .C2({ S25957[517] }),
  .ZN({ S8929 })
);
NAND3_X1 #() 
NAND3_X1_695_ (
  .A1({ S8924 }),
  .A2({ S8929 }),
  .A3({ S25957[519] }),
  .ZN({ S8931 })
);
NAND3_X1 #() 
NAND3_X1_696_ (
  .A1({ S8931 }),
  .A2({ S8910 }),
  .A3({ S8897 }),
  .ZN({ S8932 })
);
NAND3_X1 #() 
NAND3_X1_697_ (
  .A1({ S8932 }),
  .A2({ S8896 }),
  .A3({ S25957[585] }),
  .ZN({ S8933 })
);
INV_X1 #() 
INV_X1_217_ (
  .A({ S25957[585] }),
  .ZN({ S8934 })
);
NAND3_X1 #() 
NAND3_X1_698_ (
  .A1({ S8895 }),
  .A2({ S8869 }),
  .A3({ S8897 }),
  .ZN({ S8935 })
);
NAND3_X1 #() 
NAND3_X1_699_ (
  .A1({ S8931 }),
  .A2({ S8910 }),
  .A3({ S25957[617] }),
  .ZN({ S8936 })
);
NAND3_X1 #() 
NAND3_X1_700_ (
  .A1({ S8936 }),
  .A2({ S8935 }),
  .A3({ S8934 }),
  .ZN({ S8937 })
);
NAND3_X1 #() 
NAND3_X1_701_ (
  .A1({ S8933 }),
  .A2({ S8937 }),
  .A3({ S25957[649] }),
  .ZN({ S8938 })
);
NAND3_X1 #() 
NAND3_X1_702_ (
  .A1({ S8932 }),
  .A2({ S8896 }),
  .A3({ S8934 }),
  .ZN({ S8939 })
);
NAND3_X1 #() 
NAND3_X1_703_ (
  .A1({ S8936 }),
  .A2({ S8935 }),
  .A3({ S25957[585] }),
  .ZN({ S8940 })
);
NAND3_X1 #() 
NAND3_X1_704_ (
  .A1({ S8939 }),
  .A2({ S8940 }),
  .A3({ S4806 }),
  .ZN({ S8942 })
);
AND2_X1 #() 
AND2_X1_39_ (
  .A1({ S8942 }),
  .A2({ S8938 }),
  .ZN({ S25957[393] })
);
NOR2_X1 #() 
NOR2_X1_136_ (
  .A1({ S6157 }),
  .A2({ S6171 }),
  .ZN({ S25957[586] })
);
NAND2_X1 #() 
NAND2_X1_623_ (
  .A1({ S3459 }),
  .A2({ S3435 }),
  .ZN({ S8943 })
);
XNOR2_X1 #() 
XNOR2_X1_19_ (
  .A({ S8943 }),
  .B({ S25957[874] }),
  .ZN({ S25957[746] })
);
NAND2_X1 #() 
NAND2_X1_624_ (
  .A1({ S6156 }),
  .A2({ S6127 }),
  .ZN({ S8944 })
);
XOR2_X1 #() 
XOR2_X1_14_ (
  .A({ S8944 }),
  .B({ S25957[746] }),
  .Z({ S25957[618] })
);
INV_X1 #() 
INV_X1_218_ (
  .A({ S25957[618] }),
  .ZN({ S8945 })
);
NOR2_X1 #() 
NOR2_X1_137_ (
  .A1({ S8493 }),
  .A2({ S8468 }),
  .ZN({ S8946 })
);
AOI21_X1 #() 
AOI21_X1_361_ (
  .A({ S8538 }),
  .B1({ S8946 }),
  .B2({ S8333 }),
  .ZN({ S8947 })
);
NOR2_X1 #() 
NOR2_X1_138_ (
  .A1({ S8300 }),
  .A2({ S25957[515] }),
  .ZN({ S8949 })
);
NOR3_X1 #() 
NOR3_X1_20_ (
  .A1({ S8299 }),
  .A2({ S8949 }),
  .A3({ S25957[516] }),
  .ZN({ S8950 })
);
OAI21_X1 #() 
OAI21_X1_339_ (
  .A({ S8295 }),
  .B1({ S8947 }),
  .B2({ S8950 }),
  .ZN({ S8951 })
);
NAND3_X1 #() 
NAND3_X1_705_ (
  .A1({ S8536 }),
  .A2({ S25957[515] }),
  .A3({ S8606 }),
  .ZN({ S8952 })
);
AOI21_X1 #() 
AOI21_X1_362_ (
  .A({ S25957[516] }),
  .B1({ S8952 }),
  .B2({ S8304 }),
  .ZN({ S8953 })
);
OAI21_X1 #() 
OAI21_X1_340_ (
  .A({ S8371 }),
  .B1({ S25957[514] }),
  .B2({ S8342 }),
  .ZN({ S8954 })
);
AOI21_X1 #() 
AOI21_X1_363_ (
  .A({ S8340 }),
  .B1({ S8954 }),
  .B2({ S12 }),
  .ZN({ S8955 })
);
OAI21_X1 #() 
OAI21_X1_341_ (
  .A({ S25957[517] }),
  .B1({ S8955 }),
  .B2({ S6575 }),
  .ZN({ S8956 })
);
OAI211_X1 #() 
OAI211_X1_188_ (
  .A({ S8951 }),
  .B({ S25957[518] }),
  .C1({ S8953 }),
  .C2({ S8956 }),
  .ZN({ S8957 })
);
NAND2_X1 #() 
NAND2_X1_625_ (
  .A1({ S8371 }),
  .A2({ S25957[515] }),
  .ZN({ S8958 })
);
NAND3_X1 #() 
NAND3_X1_706_ (
  .A1({ S8958 }),
  .A2({ S25957[516] }),
  .A3({ S8715 }),
  .ZN({ S8960 })
);
NAND2_X1 #() 
NAND2_X1_626_ (
  .A1({ S8458 }),
  .A2({ S6575 }),
  .ZN({ S8961 })
);
NAND3_X1 #() 
NAND3_X1_707_ (
  .A1({ S8961 }),
  .A2({ S8295 }),
  .A3({ S8960 }),
  .ZN({ S8962 })
);
NAND2_X1 #() 
NAND2_X1_627_ (
  .A1({ S8326 }),
  .A2({ S12 }),
  .ZN({ S8963 })
);
NAND3_X1 #() 
NAND3_X1_708_ (
  .A1({ S8435 }),
  .A2({ S25957[515] }),
  .A3({ S8377 }),
  .ZN({ S8964 })
);
AOI21_X1 #() 
AOI21_X1_364_ (
  .A({ S25957[516] }),
  .B1({ S8964 }),
  .B2({ S8963 }),
  .ZN({ S8965 })
);
NAND3_X1 #() 
NAND3_X1_709_ (
  .A1({ S8300 }),
  .A2({ S25957[515] }),
  .A3({ S25957[512] }),
  .ZN({ S8966 })
);
AND2_X1 #() 
AND2_X1_40_ (
  .A1({ S8702 }),
  .A2({ S8966 }),
  .ZN({ S8967 })
);
OAI21_X1 #() 
OAI21_X1_342_ (
  .A({ S25957[517] }),
  .B1({ S8967 }),
  .B2({ S6575 }),
  .ZN({ S8968 })
);
OAI211_X1 #() 
OAI211_X1_189_ (
  .A({ S6416 }),
  .B({ S8962 }),
  .C1({ S8968 }),
  .C2({ S8965 }),
  .ZN({ S8969 })
);
NAND3_X1 #() 
NAND3_X1_710_ (
  .A1({ S8957 }),
  .A2({ S25957[519] }),
  .A3({ S8969 }),
  .ZN({ S8971 })
);
AOI21_X1 #() 
AOI21_X1_365_ (
  .A({ S25957[516] }),
  .B1({ S8689 }),
  .B2({ S12 }),
  .ZN({ S8972 })
);
INV_X1 #() 
INV_X1_219_ (
  .A({ S8972 }),
  .ZN({ S8973 })
);
OAI211_X1 #() 
OAI211_X1_190_ (
  .A({ S25957[516] }),
  .B({ S25957[515] }),
  .C1({ S8332 }),
  .C2({ S25957[513] }),
  .ZN({ S8974 })
);
NAND3_X1 #() 
NAND3_X1_711_ (
  .A1({ S8700 }),
  .A2({ S25957[517] }),
  .A3({ S8974 }),
  .ZN({ S8975 })
);
INV_X1 #() 
INV_X1_220_ (
  .A({ S8975 }),
  .ZN({ S8976 })
);
OAI21_X1 #() 
OAI21_X1_343_ (
  .A({ S8976 }),
  .B1({ S8379 }),
  .B2({ S8973 }),
  .ZN({ S8977 })
);
AOI21_X1 #() 
AOI21_X1_366_ (
  .A({ S12 }),
  .B1({ S8405 }),
  .B2({ S8314 }),
  .ZN({ S8978 })
);
NAND4_X1 #() 
NAND4_X1_71_ (
  .A1({ S8298 }),
  .A2({ S8300 }),
  .A3({ S8302 }),
  .A4({ S8320 }),
  .ZN({ S8979 })
);
AOI22_X1 #() 
AOI22_X1_62_ (
  .A1({ S8979 }),
  .A2({ S12 }),
  .B1({ S8978 }),
  .B2({ S8343 }),
  .ZN({ S8980 })
);
AND3_X1 #() 
AND3_X1_29_ (
  .A1({ S25957[513] }),
  .A2({ S8350 }),
  .A3({ S25957[515] }),
  .ZN({ S8981 })
);
INV_X1 #() 
INV_X1_221_ (
  .A({ S8981 }),
  .ZN({ S8982 })
);
NAND3_X1 #() 
NAND3_X1_712_ (
  .A1({ S8982 }),
  .A2({ S8778 }),
  .A3({ S6575 }),
  .ZN({ S8983 })
);
OAI211_X1 #() 
OAI211_X1_191_ (
  .A({ S8295 }),
  .B({ S8983 }),
  .C1({ S8980 }),
  .C2({ S6575 }),
  .ZN({ S8984 })
);
NAND3_X1 #() 
NAND3_X1_713_ (
  .A1({ S8984 }),
  .A2({ S8977 }),
  .A3({ S25957[518] }),
  .ZN({ S8985 })
);
AOI21_X1 #() 
AOI21_X1_367_ (
  .A({ S6575 }),
  .B1({ S8409 }),
  .B2({ S8308 }),
  .ZN({ S8986 })
);
NAND2_X1 #() 
NAND2_X1_628_ (
  .A1({ S8723 }),
  .A2({ S8986 }),
  .ZN({ S8987 })
);
NAND4_X1 #() 
NAND4_X1_72_ (
  .A1({ S8461 }),
  .A2({ S8302 }),
  .A3({ S8300 }),
  .A4({ S25957[515] }),
  .ZN({ S8988 })
);
NAND3_X1 #() 
NAND3_X1_714_ (
  .A1({ S8988 }),
  .A2({ S6575 }),
  .A3({ S8457 }),
  .ZN({ S8989 })
);
NAND2_X1 #() 
NAND2_X1_629_ (
  .A1({ S8987 }),
  .A2({ S8989 }),
  .ZN({ S8990 })
);
NAND2_X1 #() 
NAND2_X1_630_ (
  .A1({ S8990 }),
  .A2({ S25957[517] }),
  .ZN({ S8992 })
);
AOI211_X1 #() 
AOI211_X1_6_ (
  .A({ S6575 }),
  .B({ S8981 }),
  .C1({ S8601 }),
  .C2({ S12 }),
  .ZN({ S8993 })
);
AND3_X1 #() 
AND3_X1_30_ (
  .A1({ S8373 }),
  .A2({ S8884 }),
  .A3({ S8595 }),
  .ZN({ S8994 })
);
OAI21_X1 #() 
OAI21_X1_344_ (
  .A({ S8295 }),
  .B1({ S8993 }),
  .B2({ S8994 }),
  .ZN({ S8995 })
);
NAND3_X1 #() 
NAND3_X1_715_ (
  .A1({ S8995 }),
  .A2({ S8992 }),
  .A3({ S6416 }),
  .ZN({ S8996 })
);
NAND3_X1 #() 
NAND3_X1_716_ (
  .A1({ S8996 }),
  .A2({ S8294 }),
  .A3({ S8985 }),
  .ZN({ S8997 })
);
NAND3_X1 #() 
NAND3_X1_717_ (
  .A1({ S8997 }),
  .A2({ S8971 }),
  .A3({ S8945 }),
  .ZN({ S8998 })
);
AOI21_X1 #() 
AOI21_X1_368_ (
  .A({ S6575 }),
  .B1({ S8702 }),
  .B2({ S8966 }),
  .ZN({ S8999 })
);
OAI21_X1 #() 
OAI21_X1_345_ (
  .A({ S25957[517] }),
  .B1({ S8965 }),
  .B2({ S8999 }),
  .ZN({ S9000 })
);
NAND3_X1 #() 
NAND3_X1_718_ (
  .A1({ S8982 }),
  .A2({ S25957[516] }),
  .A3({ S8773 }),
  .ZN({ S9001 })
);
OAI211_X1 #() 
OAI211_X1_192_ (
  .A({ S9001 }),
  .B({ S8295 }),
  .C1({ S25957[516] }),
  .C2({ S8458 }),
  .ZN({ S9003 })
);
NAND3_X1 #() 
NAND3_X1_719_ (
  .A1({ S9000 }),
  .A2({ S9003 }),
  .A3({ S6416 }),
  .ZN({ S9004 })
);
NAND3_X1 #() 
NAND3_X1_720_ (
  .A1({ S8952 }),
  .A2({ S6575 }),
  .A3({ S8304 }),
  .ZN({ S9005 })
);
INV_X1 #() 
INV_X1_222_ (
  .A({ S8340 }),
  .ZN({ S9006 })
);
OAI21_X1 #() 
OAI21_X1_346_ (
  .A({ S12 }),
  .B1({ S8493 }),
  .B2({ S8468 }),
  .ZN({ S9007 })
);
NAND3_X1 #() 
NAND3_X1_721_ (
  .A1({ S9007 }),
  .A2({ S25957[516] }),
  .A3({ S9006 }),
  .ZN({ S9008 })
);
NAND3_X1 #() 
NAND3_X1_722_ (
  .A1({ S9005 }),
  .A2({ S25957[517] }),
  .A3({ S9008 }),
  .ZN({ S9009 })
);
NOR2_X1 #() 
NOR2_X1_139_ (
  .A1({ S8954 }),
  .A2({ S8335 }),
  .ZN({ S9010 })
);
NAND3_X1 #() 
NAND3_X1_723_ (
  .A1({ S8619 }),
  .A2({ S8798 }),
  .A3({ S6575 }),
  .ZN({ S9011 })
);
OAI211_X1 #() 
OAI211_X1_193_ (
  .A({ S8295 }),
  .B({ S9011 }),
  .C1({ S9010 }),
  .C2({ S8538 }),
  .ZN({ S9012 })
);
NAND3_X1 #() 
NAND3_X1_724_ (
  .A1({ S9009 }),
  .A2({ S25957[518] }),
  .A3({ S9012 }),
  .ZN({ S9014 })
);
NAND3_X1 #() 
NAND3_X1_725_ (
  .A1({ S9014 }),
  .A2({ S9004 }),
  .A3({ S25957[519] }),
  .ZN({ S9015 })
);
OAI21_X1 #() 
OAI21_X1_347_ (
  .A({ S25957[515] }),
  .B1({ S8327 }),
  .B2({ S8347 }),
  .ZN({ S9016 })
);
AOI21_X1 #() 
AOI21_X1_369_ (
  .A({ S8975 }),
  .B1({ S9016 }),
  .B2({ S8972 }),
  .ZN({ S9017 })
);
NAND3_X1 #() 
NAND3_X1_726_ (
  .A1({ S8590 }),
  .A2({ S6575 }),
  .A3({ S8958 }),
  .ZN({ S9018 })
);
OAI211_X1 #() 
OAI211_X1_194_ (
  .A({ S25957[515] }),
  .B({ S8343 }),
  .C1({ S8341 }),
  .C2({ S8302 }),
  .ZN({ S9019 })
);
AOI21_X1 #() 
AOI21_X1_370_ (
  .A({ S8291 }),
  .B1({ S8598 }),
  .B2({ S8321 }),
  .ZN({ S9020 })
);
OAI211_X1 #() 
OAI211_X1_195_ (
  .A({ S25957[516] }),
  .B({ S9019 }),
  .C1({ S9020 }),
  .C2({ S25957[515] }),
  .ZN({ S9021 })
);
AOI21_X1 #() 
AOI21_X1_371_ (
  .A({ S25957[517] }),
  .B1({ S9021 }),
  .B2({ S9018 }),
  .ZN({ S9022 })
);
OAI21_X1 #() 
OAI21_X1_348_ (
  .A({ S25957[518] }),
  .B1({ S9022 }),
  .B2({ S9017 }),
  .ZN({ S9023 })
);
NAND3_X1 #() 
NAND3_X1_727_ (
  .A1({ S8987 }),
  .A2({ S8989 }),
  .A3({ S25957[517] }),
  .ZN({ S9024 })
);
NAND3_X1 #() 
NAND3_X1_728_ (
  .A1({ S8602 }),
  .A2({ S25957[516] }),
  .A3({ S8982 }),
  .ZN({ S9025 })
);
NAND2_X1 #() 
NAND2_X1_631_ (
  .A1({ S8791 }),
  .A2({ S8373 }),
  .ZN({ S9026 })
);
NAND3_X1 #() 
NAND3_X1_729_ (
  .A1({ S9025 }),
  .A2({ S9026 }),
  .A3({ S8295 }),
  .ZN({ S9027 })
);
NAND3_X1 #() 
NAND3_X1_730_ (
  .A1({ S9027 }),
  .A2({ S6416 }),
  .A3({ S9024 }),
  .ZN({ S9028 })
);
NAND3_X1 #() 
NAND3_X1_731_ (
  .A1({ S9023 }),
  .A2({ S8294 }),
  .A3({ S9028 }),
  .ZN({ S9029 })
);
NAND3_X1 #() 
NAND3_X1_732_ (
  .A1({ S9029 }),
  .A2({ S9015 }),
  .A3({ S25957[618] }),
  .ZN({ S9030 })
);
NAND3_X1 #() 
NAND3_X1_733_ (
  .A1({ S8998 }),
  .A2({ S25957[586] }),
  .A3({ S9030 }),
  .ZN({ S9031 })
);
INV_X1 #() 
INV_X1_223_ (
  .A({ S25957[586] }),
  .ZN({ S9032 })
);
NAND3_X1 #() 
NAND3_X1_734_ (
  .A1({ S9029 }),
  .A2({ S9015 }),
  .A3({ S8945 }),
  .ZN({ S9033 })
);
NAND3_X1 #() 
NAND3_X1_735_ (
  .A1({ S8997 }),
  .A2({ S8971 }),
  .A3({ S25957[618] }),
  .ZN({ S9035 })
);
NAND3_X1 #() 
NAND3_X1_736_ (
  .A1({ S9035 }),
  .A2({ S9032 }),
  .A3({ S9033 }),
  .ZN({ S9036 })
);
NAND3_X1 #() 
NAND3_X1_737_ (
  .A1({ S9031 }),
  .A2({ S9036 }),
  .A3({ S25957[650] }),
  .ZN({ S9037 })
);
NAND3_X1 #() 
NAND3_X1_738_ (
  .A1({ S8998 }),
  .A2({ S9032 }),
  .A3({ S9030 }),
  .ZN({ S9038 })
);
NAND3_X1 #() 
NAND3_X1_739_ (
  .A1({ S9035 }),
  .A2({ S25957[586] }),
  .A3({ S9033 }),
  .ZN({ S9039 })
);
NAND3_X1 #() 
NAND3_X1_740_ (
  .A1({ S9038 }),
  .A2({ S9039 }),
  .A3({ S4816 }),
  .ZN({ S9040 })
);
AND2_X1 #() 
AND2_X1_41_ (
  .A1({ S9040 }),
  .A2({ S9037 }),
  .ZN({ S25957[394] })
);
AOI21_X1 #() 
AOI21_X1_372_ (
  .A({ S7386 }),
  .B1({ S7464 }),
  .B2({ S7467 }),
  .ZN({ S22 })
);
NAND3_X1 #() 
NAND3_X1_741_ (
  .A1({ S7464 }),
  .A2({ S7467 }),
  .A3({ S7386 }),
  .ZN({ S23 })
);
NAND2_X1 #() 
NAND2_X1_632_ (
  .A1({ S3594 }),
  .A2({ S3596 }),
  .ZN({ S9041 })
);
AOI21_X1 #() 
AOI21_X1_373_ (
  .A({ S25957[825] }),
  .B1({ S7458 }),
  .B2({ S7433 }),
  .ZN({ S9043 })
);
AOI21_X1 #() 
AOI21_X1_374_ (
  .A({ S4730 }),
  .B1({ S7462 }),
  .B2({ S7461 }),
  .ZN({ S9044 })
);
OAI21_X1 #() 
OAI21_X1_349_ (
  .A({ S6232 }),
  .B1({ S9043 }),
  .B2({ S9044 }),
  .ZN({ S9045 })
);
NAND3_X1 #() 
NAND3_X1_742_ (
  .A1({ S7462 }),
  .A2({ S4730 }),
  .A3({ S7461 }),
  .ZN({ S9046 })
);
NAND3_X1 #() 
NAND3_X1_743_ (
  .A1({ S7458 }),
  .A2({ S25957[825] }),
  .A3({ S7433 }),
  .ZN({ S9047 })
);
NAND3_X1 #() 
NAND3_X1_744_ (
  .A1({ S9046 }),
  .A2({ S9047 }),
  .A3({ S25957[665] }),
  .ZN({ S9048 })
);
NAND3_X1 #() 
NAND3_X1_745_ (
  .A1({ S9045 }),
  .A2({ S25957[536] }),
  .A3({ S9048 }),
  .ZN({ S9049 })
);
NOR2_X1 #() 
NOR2_X1_140_ (
  .A1({ S9049 }),
  .A2({ S25957[538] }),
  .ZN({ S9050 })
);
NAND2_X1 #() 
NAND2_X1_633_ (
  .A1({ S7555 }),
  .A2({ S7558 }),
  .ZN({ S9051 })
);
NOR2_X1 #() 
NOR2_X1_141_ (
  .A1({ S23 }),
  .A2({ S9051 }),
  .ZN({ S9052 })
);
NOR3_X1 #() 
NOR3_X1_21_ (
  .A1({ S9050 }),
  .A2({ S9052 }),
  .A3({ S15 }),
  .ZN({ S9054 })
);
AOI21_X1 #() 
AOI21_X1_375_ (
  .A({ S25957[794] }),
  .B1({ S7556 }),
  .B2({ S7557 }),
  .ZN({ S9055 })
);
AOI21_X1 #() 
AOI21_X1_376_ (
  .A({ S3488 }),
  .B1({ S7550 }),
  .B2({ S7554 }),
  .ZN({ S9056 })
);
OAI21_X1 #() 
OAI21_X1_350_ (
  .A({ S7386 }),
  .B1({ S9055 }),
  .B2({ S9056 }),
  .ZN({ S9057 })
);
NAND3_X1 #() 
NAND3_X1_746_ (
  .A1({ S9045 }),
  .A2({ S7386 }),
  .A3({ S9048 }),
  .ZN({ S9058 })
);
OAI211_X1 #() 
OAI211_X1_196_ (
  .A({ S9057 }),
  .B({ S15 }),
  .C1({ S9058 }),
  .C2({ S9051 }),
  .ZN({ S9059 })
);
NAND2_X1 #() 
NAND2_X1_634_ (
  .A1({ S9059 }),
  .A2({ S25957[540] }),
  .ZN({ S9060 })
);
NAND3_X1 #() 
NAND3_X1_747_ (
  .A1({ S7271 }),
  .A2({ S7272 }),
  .A3({ S6201 }),
  .ZN({ S9061 })
);
NAND3_X1 #() 
NAND3_X1_748_ (
  .A1({ S7269 }),
  .A2({ S7266 }),
  .A3({ S25957[668] }),
  .ZN({ S9062 })
);
NAND2_X1 #() 
NAND2_X1_635_ (
  .A1({ S9061 }),
  .A2({ S9062 }),
  .ZN({ S9063 })
);
NAND4_X1 #() 
NAND4_X1_73_ (
  .A1({ S9045 }),
  .A2({ S9048 }),
  .A3({ S7555 }),
  .A4({ S7558 }),
  .ZN({ S9065 })
);
AND3_X1 #() 
AND3_X1_31_ (
  .A1({ S7467 }),
  .A2({ S7464 }),
  .A3({ S25957[536] }),
  .ZN({ S9066 })
);
NAND2_X1 #() 
NAND2_X1_636_ (
  .A1({ S9066 }),
  .A2({ S9051 }),
  .ZN({ S9067 })
);
NAND2_X1 #() 
NAND2_X1_637_ (
  .A1({ S9067 }),
  .A2({ S9065 }),
  .ZN({ S9068 })
);
NAND2_X1 #() 
NAND2_X1_638_ (
  .A1({ S9068 }),
  .A2({ S25957[539] }),
  .ZN({ S9069 })
);
NAND4_X1 #() 
NAND4_X1_74_ (
  .A1({ S7555 }),
  .A2({ S7558 }),
  .A3({ S7464 }),
  .A4({ S7467 }),
  .ZN({ S9070 })
);
NAND3_X1 #() 
NAND3_X1_749_ (
  .A1({ S7555 }),
  .A2({ S7558 }),
  .A3({ S7386 }),
  .ZN({ S9071 })
);
NAND3_X1 #() 
NAND3_X1_750_ (
  .A1({ S9070 }),
  .A2({ S15 }),
  .A3({ S9071 }),
  .ZN({ S9072 })
);
NAND3_X1 #() 
NAND3_X1_751_ (
  .A1({ S9069 }),
  .A2({ S9063 }),
  .A3({ S9072 }),
  .ZN({ S9073 })
);
OAI21_X1 #() 
OAI21_X1_351_ (
  .A({ S9073 }),
  .B1({ S9054 }),
  .B2({ S9060 }),
  .ZN({ S9074 })
);
NAND2_X1 #() 
NAND2_X1_639_ (
  .A1({ S9051 }),
  .A2({ S25957[537] }),
  .ZN({ S9076 })
);
INV_X1 #() 
INV_X1_224_ (
  .A({ S9076 }),
  .ZN({ S9077 })
);
NAND3_X1 #() 
NAND3_X1_752_ (
  .A1({ S7555 }),
  .A2({ S7558 }),
  .A3({ S25957[536] }),
  .ZN({ S9078 })
);
NAND2_X1 #() 
NAND2_X1_640_ (
  .A1({ S9078 }),
  .A2({ S25957[539] }),
  .ZN({ S9079 })
);
NAND3_X1 #() 
NAND3_X1_753_ (
  .A1({ S7464 }),
  .A2({ S7467 }),
  .A3({ S25957[536] }),
  .ZN({ S9080 })
);
NAND2_X1 #() 
NAND2_X1_641_ (
  .A1({ S9080 }),
  .A2({ S9051 }),
  .ZN({ S9081 })
);
NAND3_X1 #() 
NAND3_X1_754_ (
  .A1({ S9081 }),
  .A2({ S9070 }),
  .A3({ S9071 }),
  .ZN({ S9082 })
);
AOI21_X1 #() 
AOI21_X1_377_ (
  .A({ S25957[540] }),
  .B1({ S9082 }),
  .B2({ S15 }),
  .ZN({ S9083 })
);
OAI21_X1 #() 
OAI21_X1_352_ (
  .A({ S9083 }),
  .B1({ S9077 }),
  .B2({ S9079 }),
  .ZN({ S9084 })
);
NAND2_X1 #() 
NAND2_X1_642_ (
  .A1({ S9049 }),
  .A2({ S25957[538] }),
  .ZN({ S9085 })
);
NAND3_X1 #() 
NAND3_X1_755_ (
  .A1({ S9058 }),
  .A2({ S9051 }),
  .A3({ S9080 }),
  .ZN({ S9087 })
);
AOI21_X1 #() 
AOI21_X1_378_ (
  .A({ S15 }),
  .B1({ S9087 }),
  .B2({ S9085 }),
  .ZN({ S9088 })
);
NAND3_X1 #() 
NAND3_X1_756_ (
  .A1({ S9049 }),
  .A2({ S25957[538] }),
  .A3({ S23 }),
  .ZN({ S9089 })
);
AOI21_X1 #() 
AOI21_X1_379_ (
  .A({ S25957[539] }),
  .B1({ S9051 }),
  .B2({ S25957[536] }),
  .ZN({ S9090 })
);
NAND2_X1 #() 
NAND2_X1_643_ (
  .A1({ S9089 }),
  .A2({ S9090 }),
  .ZN({ S9091 })
);
NAND2_X1 #() 
NAND2_X1_644_ (
  .A1({ S9091 }),
  .A2({ S25957[540] }),
  .ZN({ S9092 })
);
OAI21_X1 #() 
OAI21_X1_353_ (
  .A({ S9084 }),
  .B1({ S9088 }),
  .B2({ S9092 }),
  .ZN({ S9093 })
);
NOR2_X1 #() 
NOR2_X1_142_ (
  .A1({ S9093 }),
  .A2({ S25957[541] }),
  .ZN({ S9094 })
);
AOI21_X1 #() 
AOI21_X1_380_ (
  .A({ S9094 }),
  .B1({ S9074 }),
  .B2({ S25957[541] }),
  .ZN({ S9095 })
);
NAND3_X1 #() 
NAND3_X1_757_ (
  .A1({ S7197 }),
  .A2({ S6306 }),
  .A3({ S7200 }),
  .ZN({ S9096 })
);
NAND3_X1 #() 
NAND3_X1_758_ (
  .A1({ S7203 }),
  .A2({ S25957[669] }),
  .A3({ S7204 }),
  .ZN({ S9098 })
);
NAND2_X1 #() 
NAND2_X1_645_ (
  .A1({ S9096 }),
  .A2({ S9098 }),
  .ZN({ S9099 })
);
NOR2_X1 #() 
NOR2_X1_143_ (
  .A1({ S9058 }),
  .A2({ S9051 }),
  .ZN({ S9100 })
);
NAND2_X1 #() 
NAND2_X1_646_ (
  .A1({ S22 }),
  .A2({ S9051 }),
  .ZN({ S9101 })
);
NAND3_X1 #() 
NAND3_X1_759_ (
  .A1({ S9089 }),
  .A2({ S15 }),
  .A3({ S9101 }),
  .ZN({ S9102 })
);
OAI211_X1 #() 
OAI211_X1_197_ (
  .A({ S9102 }),
  .B({ S25957[540] }),
  .C1({ S15 }),
  .C2({ S9100 }),
  .ZN({ S9103 })
);
NAND2_X1 #() 
NAND2_X1_647_ (
  .A1({ S9070 }),
  .A2({ S9071 }),
  .ZN({ S9104 })
);
NOR2_X1 #() 
NOR2_X1_144_ (
  .A1({ S9104 }),
  .A2({ S15 }),
  .ZN({ S9105 })
);
NAND3_X1 #() 
NAND3_X1_760_ (
  .A1({ S9058 }),
  .A2({ S25957[538] }),
  .A3({ S9080 }),
  .ZN({ S9106 })
);
INV_X1 #() 
INV_X1_225_ (
  .A({ S9106 }),
  .ZN({ S9107 })
);
NOR2_X1 #() 
NOR2_X1_145_ (
  .A1({ S9107 }),
  .A2({ S25957[539] }),
  .ZN({ S9109 })
);
OAI21_X1 #() 
OAI21_X1_354_ (
  .A({ S9063 }),
  .B1({ S9109 }),
  .B2({ S9105 }),
  .ZN({ S9110 })
);
NAND3_X1 #() 
NAND3_X1_761_ (
  .A1({ S9110 }),
  .A2({ S9099 }),
  .A3({ S9103 }),
  .ZN({ S9111 })
);
NAND3_X1 #() 
NAND3_X1_762_ (
  .A1({ S7555 }),
  .A2({ S7558 }),
  .A3({ S25957[539] }),
  .ZN({ S9112 })
);
NAND3_X1 #() 
NAND3_X1_763_ (
  .A1({ S7464 }),
  .A2({ S7467 }),
  .A3({ S25957[539] }),
  .ZN({ S9113 })
);
NAND2_X1 #() 
NAND2_X1_648_ (
  .A1({ S9112 }),
  .A2({ S9113 }),
  .ZN({ S9114 })
);
NAND2_X1 #() 
NAND2_X1_649_ (
  .A1({ S9114 }),
  .A2({ S9080 }),
  .ZN({ S9115 })
);
NAND2_X1 #() 
NAND2_X1_650_ (
  .A1({ S9049 }),
  .A2({ S9051 }),
  .ZN({ S9116 })
);
AOI21_X1 #() 
AOI21_X1_381_ (
  .A({ S25957[539] }),
  .B1({ S25957[538] }),
  .B2({ S25957[537] }),
  .ZN({ S9117 })
);
NAND2_X1 #() 
NAND2_X1_651_ (
  .A1({ S9117 }),
  .A2({ S9116 }),
  .ZN({ S9118 })
);
AOI21_X1 #() 
AOI21_X1_382_ (
  .A({ S25957[540] }),
  .B1({ S9118 }),
  .B2({ S9115 }),
  .ZN({ S9120 })
);
NAND2_X1 #() 
NAND2_X1_652_ (
  .A1({ S25957[537] }),
  .A2({ S25957[539] }),
  .ZN({ S9121 })
);
NAND2_X1 #() 
NAND2_X1_653_ (
  .A1({ S9121 }),
  .A2({ S9112 }),
  .ZN({ S9122 })
);
NOR2_X1 #() 
NOR2_X1_146_ (
  .A1({ S25957[539] }),
  .A2({ S7386 }),
  .ZN({ S9123 })
);
AOI211_X1 #() 
AOI211_X1_7_ (
  .A({ S9123 }),
  .B({ S9063 }),
  .C1({ S9122 }),
  .C2({ S9078 }),
  .ZN({ S9124 })
);
OR3_X1 #() 
OR3_X1_2_ (
  .A1({ S9120 }),
  .A2({ S9124 }),
  .A3({ S9099 }),
  .ZN({ S9125 })
);
NAND3_X1 #() 
NAND3_X1_764_ (
  .A1({ S9125 }),
  .A2({ S9111 }),
  .A3({ S7106 }),
  .ZN({ S9126 })
);
OAI211_X1 #() 
OAI211_X1_198_ (
  .A({ S7026 }),
  .B({ S9126 }),
  .C1({ S9095 }),
  .C2({ S7106 }),
  .ZN({ S9127 })
);
AND3_X1 #() 
AND3_X1_32_ (
  .A1({ S7467 }),
  .A2({ S7464 }),
  .A3({ S7386 }),
  .ZN({ S9128 })
);
NAND2_X1 #() 
NAND2_X1_654_ (
  .A1({ S9128 }),
  .A2({ S25957[538] }),
  .ZN({ S9129 })
);
OAI211_X1 #() 
OAI211_X1_199_ (
  .A({ S9129 }),
  .B({ S9076 }),
  .C1({ S9090 }),
  .C2({ S25957[539] }),
  .ZN({ S9130 })
);
NAND2_X1 #() 
NAND2_X1_655_ (
  .A1({ S25957[539] }),
  .A2({ S7386 }),
  .ZN({ S9131 })
);
NAND2_X1 #() 
NAND2_X1_656_ (
  .A1({ S9113 }),
  .A2({ S9131 }),
  .ZN({ S9132 })
);
NAND2_X1 #() 
NAND2_X1_657_ (
  .A1({ S9132 }),
  .A2({ S9070 }),
  .ZN({ S9133 })
);
NAND2_X1 #() 
NAND2_X1_658_ (
  .A1({ S9058 }),
  .A2({ S15 }),
  .ZN({ S9134 })
);
NAND3_X1 #() 
NAND3_X1_765_ (
  .A1({ S9133 }),
  .A2({ S25957[540] }),
  .A3({ S9134 }),
  .ZN({ S9135 })
);
OAI21_X1 #() 
OAI21_X1_355_ (
  .A({ S9135 }),
  .B1({ S9130 }),
  .B2({ S25957[540] }),
  .ZN({ S9136 })
);
OAI211_X1 #() 
OAI211_X1_200_ (
  .A({ S25957[539] }),
  .B({ S9071 }),
  .C1({ S25957[538] }),
  .C2({ S9080 }),
  .ZN({ S9137 })
);
AOI21_X1 #() 
AOI21_X1_383_ (
  .A({ S25957[536] }),
  .B1({ S7555 }),
  .B2({ S7558 }),
  .ZN({ S9138 })
);
NOR2_X1 #() 
NOR2_X1_147_ (
  .A1({ S9138 }),
  .A2({ S25957[539] }),
  .ZN({ S9139 })
);
NAND2_X1 #() 
NAND2_X1_659_ (
  .A1({ S9139 }),
  .A2({ S25957[537] }),
  .ZN({ S9141 })
);
NAND3_X1 #() 
NAND3_X1_766_ (
  .A1({ S9141 }),
  .A2({ S25957[540] }),
  .A3({ S9137 }),
  .ZN({ S9142 })
);
NAND2_X1 #() 
NAND2_X1_660_ (
  .A1({ S9058 }),
  .A2({ S9078 }),
  .ZN({ S9143 })
);
AOI21_X1 #() 
AOI21_X1_384_ (
  .A({ S25957[536] }),
  .B1({ S7464 }),
  .B2({ S7467 }),
  .ZN({ S9144 })
);
AOI21_X1 #() 
AOI21_X1_385_ (
  .A({ S9066 }),
  .B1({ S25957[538] }),
  .B2({ S9144 }),
  .ZN({ S9145 })
);
OAI21_X1 #() 
OAI21_X1_356_ (
  .A({ S15 }),
  .B1({ S25957[538] }),
  .B2({ S25957[537] }),
  .ZN({ S9146 })
);
OAI221_X1 #() 
OAI221_X1_13_ (
  .A({ S9063 }),
  .B1({ S9146 }),
  .B2({ S9143 }),
  .C1({ S9145 }),
  .C2({ S15 }),
  .ZN({ S9147 })
);
NAND3_X1 #() 
NAND3_X1_767_ (
  .A1({ S9147 }),
  .A2({ S25957[541] }),
  .A3({ S9142 }),
  .ZN({ S9148 })
);
OAI21_X1 #() 
OAI21_X1_357_ (
  .A({ S9148 }),
  .B1({ S25957[541] }),
  .B2({ S9136 }),
  .ZN({ S9149 })
);
NAND2_X1 #() 
NAND2_X1_661_ (
  .A1({ S9149 }),
  .A2({ S25957[542] }),
  .ZN({ S9150 })
);
NAND3_X1 #() 
NAND3_X1_768_ (
  .A1({ S9049 }),
  .A2({ S9051 }),
  .A3({ S23 }),
  .ZN({ S9152 })
);
NAND3_X1 #() 
NAND3_X1_769_ (
  .A1({ S9106 }),
  .A2({ S9152 }),
  .A3({ S25957[539] }),
  .ZN({ S9153 })
);
NAND2_X1 #() 
NAND2_X1_662_ (
  .A1({ S9090 }),
  .A2({ S9065 }),
  .ZN({ S9154 })
);
AOI21_X1 #() 
AOI21_X1_386_ (
  .A({ S9063 }),
  .B1({ S9153 }),
  .B2({ S9154 }),
  .ZN({ S9155 })
);
INV_X1 #() 
INV_X1_226_ (
  .A({ S9122 }),
  .ZN({ S9156 })
);
NAND2_X1 #() 
NAND2_X1_663_ (
  .A1({ S9065 }),
  .A2({ S9071 }),
  .ZN({ S9157 })
);
AOI22_X1 #() 
AOI22_X1_63_ (
  .A1({ S9058 }),
  .A2({ S9080 }),
  .B1({ S7558 }),
  .B2({ S7555 }),
  .ZN({ S9158 })
);
OAI21_X1 #() 
OAI21_X1_358_ (
  .A({ S15 }),
  .B1({ S9158 }),
  .B2({ S9157 }),
  .ZN({ S9159 })
);
AOI21_X1 #() 
AOI21_X1_387_ (
  .A({ S25957[540] }),
  .B1({ S9159 }),
  .B2({ S9156 }),
  .ZN({ S9160 })
);
OR2_X1 #() 
OR2_X1_8_ (
  .A1({ S9160 }),
  .A2({ S9155 }),
  .ZN({ S9161 })
);
AOI21_X1 #() 
AOI21_X1_388_ (
  .A({ S25957[539] }),
  .B1({ S7464 }),
  .B2({ S7467 }),
  .ZN({ S9163 })
);
NAND2_X1 #() 
NAND2_X1_664_ (
  .A1({ S9163 }),
  .A2({ S9078 }),
  .ZN({ S9164 })
);
NAND4_X1 #() 
NAND4_X1_75_ (
  .A1({ S7558 }),
  .A2({ S7555 }),
  .A3({ S25957[536] }),
  .A4({ S25957[539] }),
  .ZN({ S9165 })
);
NAND3_X1 #() 
NAND3_X1_770_ (
  .A1({ S25957[540] }),
  .A2({ S9165 }),
  .A3({ S9113 }),
  .ZN({ S9166 })
);
INV_X1 #() 
INV_X1_227_ (
  .A({ S9166 }),
  .ZN({ S9167 })
);
INV_X1 #() 
INV_X1_228_ (
  .A({ S9132 }),
  .ZN({ S9168 })
);
NAND2_X1 #() 
NAND2_X1_665_ (
  .A1({ S9045 }),
  .A2({ S9048 }),
  .ZN({ S9169 })
);
NAND3_X1 #() 
NAND3_X1_771_ (
  .A1({ S9169 }),
  .A2({ S7386 }),
  .A3({ S9051 }),
  .ZN({ S9170 })
);
AOI21_X1 #() 
AOI21_X1_389_ (
  .A({ S25957[540] }),
  .B1({ S9168 }),
  .B2({ S9170 }),
  .ZN({ S9171 })
);
AOI211_X1 #() 
AOI211_X1_8_ (
  .A({ S9099 }),
  .B({ S9171 }),
  .C1({ S9164 }),
  .C2({ S9167 }),
  .ZN({ S9172 })
);
AOI21_X1 #() 
AOI21_X1_390_ (
  .A({ S9172 }),
  .B1({ S9161 }),
  .B2({ S9099 }),
  .ZN({ S9174 })
);
OAI211_X1 #() 
OAI211_X1_201_ (
  .A({ S25957[543] }),
  .B({ S9150 }),
  .C1({ S9174 }),
  .C2({ S25957[542] }),
  .ZN({ S9175 })
);
AOI21_X1 #() 
AOI21_X1_391_ (
  .A({ S9041 }),
  .B1({ S9127 }),
  .B2({ S9175 }),
  .ZN({ S9176 })
);
NAND3_X1 #() 
NAND3_X1_772_ (
  .A1({ S9127 }),
  .A2({ S9175 }),
  .A3({ S9041 }),
  .ZN({ S9177 })
);
INV_X1 #() 
INV_X1_229_ (
  .A({ S9177 }),
  .ZN({ S9178 })
);
OAI21_X1 #() 
OAI21_X1_359_ (
  .A({ S25957[551] }),
  .B1({ S9178 }),
  .B2({ S9176 }),
  .ZN({ S9179 })
);
INV_X1 #() 
INV_X1_230_ (
  .A({ S9176 }),
  .ZN({ S9180 })
);
NAND3_X1 #() 
NAND3_X1_773_ (
  .A1({ S9180 }),
  .A2({ S9177 }),
  .A3({ S6332 }),
  .ZN({ S9181 })
);
NAND3_X1 #() 
NAND3_X1_774_ (
  .A1({ S9179 }),
  .A2({ S9181 }),
  .A3({ S8294 }),
  .ZN({ S9182 })
);
NAND2_X1 #() 
NAND2_X1_666_ (
  .A1({ S9179 }),
  .A2({ S9181 }),
  .ZN({ S25957[423] })
);
NAND2_X1 #() 
NAND2_X1_667_ (
  .A1({ S25957[423] }),
  .A2({ S25957[519] }),
  .ZN({ S9184 })
);
AND2_X1 #() 
AND2_X1_42_ (
  .A1({ S9184 }),
  .A2({ S9182 }),
  .ZN({ S25957[391] })
);
INV_X1 #() 
INV_X1_231_ (
  .A({ S25957[678] }),
  .ZN({ S9185 })
);
INV_X1 #() 
INV_X1_232_ (
  .A({ S6336 }),
  .ZN({ S25957[870] })
);
XNOR2_X1 #() 
XNOR2_X1_20_ (
  .A({ S3675 }),
  .B({ S25957[870] }),
  .ZN({ S25957[742] })
);
XNOR2_X1 #() 
XNOR2_X1_21_ (
  .A({ S6411 }),
  .B({ S25957[742] }),
  .ZN({ S25957[614] })
);
INV_X1 #() 
INV_X1_233_ (
  .A({ S25957[614] }),
  .ZN({ S9186 })
);
NAND2_X1 #() 
NAND2_X1_668_ (
  .A1({ S9058 }),
  .A2({ S9080 }),
  .ZN({ S9187 })
);
INV_X1 #() 
INV_X1_234_ (
  .A({ S9090 }),
  .ZN({ S9188 })
);
AOI21_X1 #() 
AOI21_X1_392_ (
  .A({ S15 }),
  .B1({ S9144 }),
  .B2({ S9051 }),
  .ZN({ S9189 })
);
AOI21_X1 #() 
AOI21_X1_393_ (
  .A({ S25957[540] }),
  .B1({ S9189 }),
  .B2({ S9070 }),
  .ZN({ S9191 })
);
OAI21_X1 #() 
OAI21_X1_360_ (
  .A({ S9191 }),
  .B1({ S9187 }),
  .B2({ S9188 }),
  .ZN({ S9192 })
);
NAND4_X1 #() 
NAND4_X1_76_ (
  .A1({ S9058 }),
  .A2({ S25957[538] }),
  .A3({ S9080 }),
  .A4({ S15 }),
  .ZN({ S9193 })
);
INV_X1 #() 
INV_X1_235_ (
  .A({ S9193 }),
  .ZN({ S9194 })
);
NAND2_X1 #() 
NAND2_X1_669_ (
  .A1({ S9138 }),
  .A2({ S9163 }),
  .ZN({ S9195 })
);
OAI21_X1 #() 
OAI21_X1_361_ (
  .A({ S9195 }),
  .B1({ S15 }),
  .B2({ S9065 }),
  .ZN({ S9196 })
);
OAI21_X1 #() 
OAI21_X1_362_ (
  .A({ S25957[540] }),
  .B1({ S9194 }),
  .B2({ S9196 }),
  .ZN({ S9197 })
);
NAND3_X1 #() 
NAND3_X1_775_ (
  .A1({ S9192 }),
  .A2({ S25957[541] }),
  .A3({ S9197 }),
  .ZN({ S9198 })
);
NAND2_X1 #() 
NAND2_X1_670_ (
  .A1({ S9071 }),
  .A2({ S15 }),
  .ZN({ S9199 })
);
INV_X1 #() 
INV_X1_236_ (
  .A({ S9087 }),
  .ZN({ S9200 })
);
NOR2_X1 #() 
NOR2_X1_148_ (
  .A1({ S9200 }),
  .A2({ S9199 }),
  .ZN({ S9202 })
);
OAI21_X1 #() 
OAI21_X1_363_ (
  .A({ S25957[539] }),
  .B1({ S25957[538] }),
  .B2({ S22 }),
  .ZN({ S9203 })
);
OAI21_X1 #() 
OAI21_X1_364_ (
  .A({ S9083 }),
  .B1({ S9128 }),
  .B2({ S9203 }),
  .ZN({ S9204 })
);
OAI21_X1 #() 
OAI21_X1_365_ (
  .A({ S25957[539] }),
  .B1({ S9080 }),
  .B2({ S9051 }),
  .ZN({ S9205 })
);
OAI21_X1 #() 
OAI21_X1_366_ (
  .A({ S25957[540] }),
  .B1({ S9205 }),
  .B2({ S9138 }),
  .ZN({ S9206 })
);
OAI21_X1 #() 
OAI21_X1_367_ (
  .A({ S9204 }),
  .B1({ S9202 }),
  .B2({ S9206 }),
  .ZN({ S9207 })
);
NAND2_X1 #() 
NAND2_X1_671_ (
  .A1({ S9065 }),
  .A2({ S9078 }),
  .ZN({ S9208 })
);
AOI21_X1 #() 
AOI21_X1_394_ (
  .A({ S7386 }),
  .B1({ S7555 }),
  .B2({ S7558 }),
  .ZN({ S9209 })
);
NOR2_X1 #() 
NOR2_X1_149_ (
  .A1({ S9209 }),
  .A2({ S9113 }),
  .ZN({ S9210 })
);
NAND2_X1 #() 
NAND2_X1_672_ (
  .A1({ S9210 }),
  .A2({ S9071 }),
  .ZN({ S9211 })
);
INV_X1 #() 
INV_X1_237_ (
  .A({ S9211 }),
  .ZN({ S9213 })
);
AOI211_X1 #() 
AOI211_X1_9_ (
  .A({ S9063 }),
  .B({ S9213 }),
  .C1({ S15 }),
  .C2({ S9208 }),
  .ZN({ S9214 })
);
INV_X1 #() 
INV_X1_238_ (
  .A({ S9163 }),
  .ZN({ S9215 })
);
AOI21_X1 #() 
AOI21_X1_395_ (
  .A({ S25957[540] }),
  .B1({ S9133 }),
  .B2({ S9215 }),
  .ZN({ S9216 })
);
OAI21_X1 #() 
OAI21_X1_368_ (
  .A({ S25957[541] }),
  .B1({ S9214 }),
  .B2({ S9216 }),
  .ZN({ S9217 })
);
OAI21_X1 #() 
OAI21_X1_369_ (
  .A({ S9217 }),
  .B1({ S9207 }),
  .B2({ S25957[541] }),
  .ZN({ S9218 })
);
AOI21_X1 #() 
AOI21_X1_396_ (
  .A({ S9209 }),
  .B1({ S25957[538] }),
  .B2({ S9144 }),
  .ZN({ S9219 })
);
NOR2_X1 #() 
NOR2_X1_150_ (
  .A1({ S9219 }),
  .A2({ S15 }),
  .ZN({ S9220 })
);
OAI21_X1 #() 
OAI21_X1_370_ (
  .A({ S9063 }),
  .B1({ S9202 }),
  .B2({ S9220 }),
  .ZN({ S9221 })
);
NOR2_X1 #() 
NOR2_X1_151_ (
  .A1({ S9081 }),
  .A2({ S25957[539] }),
  .ZN({ S9222 })
);
OAI211_X1 #() 
OAI211_X1_202_ (
  .A({ S9221 }),
  .B({ S9099 }),
  .C1({ S9166 }),
  .C2({ S9222 }),
  .ZN({ S9224 })
);
AND2_X1 #() 
AND2_X1_43_ (
  .A1({ S9224 }),
  .A2({ S7106 }),
  .ZN({ S9225 })
);
AOI22_X1 #() 
AOI22_X1_64_ (
  .A1({ S9225 }),
  .A2({ S9198 }),
  .B1({ S25957[542] }),
  .B2({ S9218 }),
  .ZN({ S9226 })
);
NOR2_X1 #() 
NOR2_X1_152_ (
  .A1({ S9090 }),
  .A2({ S9063 }),
  .ZN({ S9227 })
);
AOI21_X1 #() 
AOI21_X1_397_ (
  .A({ S15 }),
  .B1({ S9128 }),
  .B2({ S25957[538] }),
  .ZN({ S9228 })
);
NAND2_X1 #() 
NAND2_X1_673_ (
  .A1({ S9228 }),
  .A2({ S9049 }),
  .ZN({ S9229 })
);
AOI22_X1 #() 
AOI22_X1_65_ (
  .A1({ S9117 }),
  .A2({ S9067 }),
  .B1({ S9114 }),
  .B2({ S9070 }),
  .ZN({ S9230 })
);
AOI22_X1 #() 
AOI22_X1_66_ (
  .A1({ S9230 }),
  .A2({ S9063 }),
  .B1({ S9227 }),
  .B2({ S9229 }),
  .ZN({ S9231 })
);
NAND3_X1 #() 
NAND3_X1_776_ (
  .A1({ S9069 }),
  .A2({ S9215 }),
  .A3({ S9227 }),
  .ZN({ S9232 })
);
AOI22_X1 #() 
AOI22_X1_67_ (
  .A1({ S25957[537] }),
  .A2({ S7386 }),
  .B1({ S7555 }),
  .B2({ S7558 }),
  .ZN({ S9233 })
);
OAI21_X1 #() 
OAI21_X1_371_ (
  .A({ S25957[539] }),
  .B1({ S9100 }),
  .B2({ S9233 }),
  .ZN({ S9235 })
);
OAI211_X1 #() 
OAI211_X1_203_ (
  .A({ S9232 }),
  .B({ S9099 }),
  .C1({ S25957[540] }),
  .C2({ S9235 }),
  .ZN({ S9236 })
);
OAI21_X1 #() 
OAI21_X1_372_ (
  .A({ S9236 }),
  .B1({ S9231 }),
  .B2({ S9099 }),
  .ZN({ S9237 })
);
OAI21_X1 #() 
OAI21_X1_373_ (
  .A({ S25957[536] }),
  .B1({ S9055 }),
  .B2({ S9056 }),
  .ZN({ S9238 })
);
NAND3_X1 #() 
NAND3_X1_777_ (
  .A1({ S9238 }),
  .A2({ S25957[539] }),
  .A3({ S23 }),
  .ZN({ S9239 })
);
INV_X1 #() 
INV_X1_239_ (
  .A({ S9239 }),
  .ZN({ S9240 })
);
NAND2_X1 #() 
NAND2_X1_674_ (
  .A1({ S9238 }),
  .A2({ S25957[537] }),
  .ZN({ S9241 })
);
NOR2_X1 #() 
NOR2_X1_153_ (
  .A1({ S9241 }),
  .A2({ S25957[539] }),
  .ZN({ S9242 })
);
OAI21_X1 #() 
OAI21_X1_374_ (
  .A({ S9063 }),
  .B1({ S9242 }),
  .B2({ S9240 }),
  .ZN({ S9243 })
);
NAND4_X1 #() 
NAND4_X1_77_ (
  .A1({ S9238 }),
  .A2({ S9070 }),
  .A3({ S15 }),
  .A4({ S9071 }),
  .ZN({ S9244 })
);
NAND3_X1 #() 
NAND3_X1_778_ (
  .A1({ S9244 }),
  .A2({ S25957[540] }),
  .A3({ S9239 }),
  .ZN({ S9246 })
);
NAND3_X1 #() 
NAND3_X1_779_ (
  .A1({ S9243 }),
  .A2({ S25957[541] }),
  .A3({ S9246 }),
  .ZN({ S9247 })
);
AOI21_X1 #() 
AOI21_X1_398_ (
  .A({ S9051 }),
  .B1({ S9058 }),
  .B2({ S9080 }),
  .ZN({ S9248 })
);
NOR2_X1 #() 
NOR2_X1_154_ (
  .A1({ S9248 }),
  .A2({ S25957[539] }),
  .ZN({ S9249 })
);
OAI21_X1 #() 
OAI21_X1_375_ (
  .A({ S9063 }),
  .B1({ S9205 }),
  .B2({ S9138 }),
  .ZN({ S9250 })
);
NAND3_X1 #() 
NAND3_X1_780_ (
  .A1({ S9051 }),
  .A2({ S25957[537] }),
  .A3({ S25957[539] }),
  .ZN({ S9251 })
);
OAI211_X1 #() 
OAI211_X1_204_ (
  .A({ S25957[540] }),
  .B({ S9251 }),
  .C1({ S9146 }),
  .C2({ S25957[536] }),
  .ZN({ S9252 })
);
OAI21_X1 #() 
OAI21_X1_376_ (
  .A({ S9252 }),
  .B1({ S9249 }),
  .B2({ S9250 }),
  .ZN({ S9253 })
);
NAND2_X1 #() 
NAND2_X1_675_ (
  .A1({ S9253 }),
  .A2({ S9099 }),
  .ZN({ S9254 })
);
NAND3_X1 #() 
NAND3_X1_781_ (
  .A1({ S9254 }),
  .A2({ S25957[542] }),
  .A3({ S9247 }),
  .ZN({ S9255 })
);
OAI21_X1 #() 
OAI21_X1_377_ (
  .A({ S9255 }),
  .B1({ S9237 }),
  .B2({ S25957[542] }),
  .ZN({ S9257 })
);
NAND2_X1 #() 
NAND2_X1_676_ (
  .A1({ S9257 }),
  .A2({ S7026 }),
  .ZN({ S9258 })
);
OAI211_X1 #() 
OAI211_X1_205_ (
  .A({ S9186 }),
  .B({ S9258 }),
  .C1({ S9226 }),
  .C2({ S7026 }),
  .ZN({ S9259 })
);
OR2_X1 #() 
OR2_X1_9_ (
  .A1({ S9257 }),
  .A2({ S25957[543] }),
  .ZN({ S9260 })
);
NAND2_X1 #() 
NAND2_X1_677_ (
  .A1({ S9226 }),
  .A2({ S25957[543] }),
  .ZN({ S9261 })
);
NAND3_X1 #() 
NAND3_X1_782_ (
  .A1({ S9261 }),
  .A2({ S9260 }),
  .A3({ S25957[614] }),
  .ZN({ S9262 })
);
NAND3_X1 #() 
NAND3_X1_783_ (
  .A1({ S9262 }),
  .A2({ S9185 }),
  .A3({ S9259 }),
  .ZN({ S9263 })
);
NAND2_X1 #() 
NAND2_X1_678_ (
  .A1({ S9262 }),
  .A2({ S9259 }),
  .ZN({ S25957[486] })
);
NAND2_X1 #() 
NAND2_X1_679_ (
  .A1({ S25957[486] }),
  .A2({ S25957[678] }),
  .ZN({ S9264 })
);
NAND3_X1 #() 
NAND3_X1_784_ (
  .A1({ S9264 }),
  .A2({ S6416 }),
  .A3({ S9263 }),
  .ZN({ S9265 })
);
NAND2_X1 #() 
NAND2_X1_680_ (
  .A1({ S25957[486] }),
  .A2({ S9185 }),
  .ZN({ S9267 })
);
NAND3_X1 #() 
NAND3_X1_785_ (
  .A1({ S9262 }),
  .A2({ S25957[678] }),
  .A3({ S9259 }),
  .ZN({ S9268 })
);
NAND3_X1 #() 
NAND3_X1_786_ (
  .A1({ S9267 }),
  .A2({ S9268 }),
  .A3({ S25957[518] }),
  .ZN({ S9269 })
);
NAND2_X1 #() 
NAND2_X1_681_ (
  .A1({ S9265 }),
  .A2({ S9269 }),
  .ZN({ S25957[390] })
);
AOI21_X1 #() 
AOI21_X1_399_ (
  .A({ S9233 }),
  .B1({ S9144 }),
  .B2({ S15 }),
  .ZN({ S9270 })
);
OAI221_X1 #() 
OAI221_X1_14_ (
  .A({ S9099 }),
  .B1({ S9250 }),
  .B2({ S9194 }),
  .C1({ S9270 }),
  .C2({ S9063 }),
  .ZN({ S9271 })
);
AOI21_X1 #() 
AOI21_X1_400_ (
  .A({ S25957[539] }),
  .B1({ S25957[537] }),
  .B2({ S7386 }),
  .ZN({ S9272 })
);
AOI22_X1 #() 
AOI22_X1_68_ (
  .A1({ S9122 }),
  .A2({ S7386 }),
  .B1({ S9272 }),
  .B2({ S9081 }),
  .ZN({ S9273 })
);
NAND2_X1 #() 
NAND2_X1_682_ (
  .A1({ S9132 }),
  .A2({ S9065 }),
  .ZN({ S9274 })
);
NAND4_X1 #() 
NAND4_X1_78_ (
  .A1({ S9274 }),
  .A2({ S9215 }),
  .A3({ S9078 }),
  .A4({ S9063 }),
  .ZN({ S9275 })
);
OAI211_X1 #() 
OAI211_X1_206_ (
  .A({ S9275 }),
  .B({ S25957[541] }),
  .C1({ S9273 }),
  .C2({ S9063 }),
  .ZN({ S9277 })
);
AOI21_X1 #() 
AOI21_X1_401_ (
  .A({ S7106 }),
  .B1({ S9271 }),
  .B2({ S9277 }),
  .ZN({ S9278 })
);
AOI22_X1 #() 
AOI22_X1_69_ (
  .A1({ S9105 }),
  .A2({ S9081 }),
  .B1({ S9049 }),
  .B2({ S9139 }),
  .ZN({ S9279 })
);
INV_X1 #() 
INV_X1_240_ (
  .A({ S9113 }),
  .ZN({ S9280 })
);
OAI211_X1 #() 
OAI211_X1_207_ (
  .A({ S7464 }),
  .B({ S7467 }),
  .C1({ S9056 }),
  .C2({ S9055 }),
  .ZN({ S9281 })
);
INV_X1 #() 
INV_X1_241_ (
  .A({ S9281 }),
  .ZN({ S9282 })
);
NOR2_X1 #() 
NOR2_X1_155_ (
  .A1({ S9282 }),
  .A2({ S9134 }),
  .ZN({ S9283 })
);
OAI21_X1 #() 
OAI21_X1_378_ (
  .A({ S9063 }),
  .B1({ S9283 }),
  .B2({ S9280 }),
  .ZN({ S9284 })
);
OAI21_X1 #() 
OAI21_X1_379_ (
  .A({ S9284 }),
  .B1({ S9279 }),
  .B2({ S9063 }),
  .ZN({ S9285 })
);
NAND2_X1 #() 
NAND2_X1_683_ (
  .A1({ S9285 }),
  .A2({ S25957[541] }),
  .ZN({ S9286 })
);
NAND2_X1 #() 
NAND2_X1_684_ (
  .A1({ S25957[537] }),
  .A2({ S9123 }),
  .ZN({ S9288 })
);
NAND3_X1 #() 
NAND3_X1_787_ (
  .A1({ S9089 }),
  .A2({ S25957[539] }),
  .A3({ S9170 }),
  .ZN({ S9289 })
);
OAI211_X1 #() 
OAI211_X1_208_ (
  .A({ S9289 }),
  .B({ S9063 }),
  .C1({ S25957[538] }),
  .C2({ S9288 }),
  .ZN({ S9290 })
);
NAND2_X1 #() 
NAND2_X1_685_ (
  .A1({ S9158 }),
  .A2({ S25957[539] }),
  .ZN({ S9291 })
);
AOI21_X1 #() 
AOI21_X1_402_ (
  .A({ S9063 }),
  .B1({ S9090 }),
  .B2({ S9169 }),
  .ZN({ S9292 })
);
NAND2_X1 #() 
NAND2_X1_686_ (
  .A1({ S9291 }),
  .A2({ S9292 }),
  .ZN({ S9293 })
);
NAND2_X1 #() 
NAND2_X1_687_ (
  .A1({ S9290 }),
  .A2({ S9293 }),
  .ZN({ S9294 })
);
NAND2_X1 #() 
NAND2_X1_688_ (
  .A1({ S9294 }),
  .A2({ S9099 }),
  .ZN({ S9295 })
);
AOI21_X1 #() 
AOI21_X1_403_ (
  .A({ S25957[542] }),
  .B1({ S9286 }),
  .B2({ S9295 }),
  .ZN({ S9296 })
);
OAI21_X1 #() 
OAI21_X1_380_ (
  .A({ S25957[543] }),
  .B1({ S9296 }),
  .B2({ S9278 }),
  .ZN({ S9297 })
);
AOI22_X1 #() 
AOI22_X1_70_ (
  .A1({ S9068 }),
  .A2({ S15 }),
  .B1({ S9106 }),
  .B2({ S9189 }),
  .ZN({ S9299 })
);
NAND2_X1 #() 
NAND2_X1_689_ (
  .A1({ S9078 }),
  .A2({ S23 }),
  .ZN({ S9300 })
);
NAND2_X1 #() 
NAND2_X1_690_ (
  .A1({ S9300 }),
  .A2({ S15 }),
  .ZN({ S9301 })
);
NAND3_X1 #() 
NAND3_X1_788_ (
  .A1({ S9301 }),
  .A2({ S9063 }),
  .A3({ S9131 }),
  .ZN({ S9302 })
);
OAI211_X1 #() 
OAI211_X1_209_ (
  .A({ S9302 }),
  .B({ S25957[541] }),
  .C1({ S9063 }),
  .C2({ S9299 }),
  .ZN({ S9303 })
);
NOR2_X1 #() 
NOR2_X1_156_ (
  .A1({ S9049 }),
  .A2({ S9051 }),
  .ZN({ S9304 })
);
NOR2_X1 #() 
NOR2_X1_157_ (
  .A1({ S9304 }),
  .A2({ S25957[539] }),
  .ZN({ S9305 })
);
OAI21_X1 #() 
OAI21_X1_381_ (
  .A({ S25957[540] }),
  .B1({ S9081 }),
  .B2({ S15 }),
  .ZN({ S9306 })
);
AOI21_X1 #() 
AOI21_X1_404_ (
  .A({ S9306 }),
  .B1({ S9305 }),
  .B2({ S9116 }),
  .ZN({ S9307 })
);
NAND4_X1 #() 
NAND4_X1_79_ (
  .A1({ S9238 }),
  .A2({ S9070 }),
  .A3({ S25957[539] }),
  .A4({ S9071 }),
  .ZN({ S9308 })
);
AOI21_X1 #() 
AOI21_X1_405_ (
  .A({ S25957[539] }),
  .B1({ S9051 }),
  .B2({ S25957[537] }),
  .ZN({ S9310 })
);
OAI21_X1 #() 
OAI21_X1_382_ (
  .A({ S9078 }),
  .B1({ S9310 }),
  .B2({ S9123 }),
  .ZN({ S9311 })
);
AOI21_X1 #() 
AOI21_X1_406_ (
  .A({ S25957[540] }),
  .B1({ S9311 }),
  .B2({ S9308 }),
  .ZN({ S9312 })
);
OAI21_X1 #() 
OAI21_X1_383_ (
  .A({ S9099 }),
  .B1({ S9312 }),
  .B2({ S9307 }),
  .ZN({ S9313 })
);
AOI21_X1 #() 
AOI21_X1_407_ (
  .A({ S7106 }),
  .B1({ S9303 }),
  .B2({ S9313 }),
  .ZN({ S9314 })
);
NAND3_X1 #() 
NAND3_X1_789_ (
  .A1({ S9238 }),
  .A2({ S25957[537] }),
  .A3({ S9071 }),
  .ZN({ S9315 })
);
OAI211_X1 #() 
OAI211_X1_210_ (
  .A({ S9063 }),
  .B({ S9165 }),
  .C1({ S9315 }),
  .C2({ S25957[539] }),
  .ZN({ S9316 })
);
OAI21_X1 #() 
OAI21_X1_384_ (
  .A({ S15 }),
  .B1({ S9058 }),
  .B2({ S25957[538] }),
  .ZN({ S9317 })
);
OAI211_X1 #() 
OAI211_X1_211_ (
  .A({ S9317 }),
  .B({ S25957[540] }),
  .C1({ S9168 }),
  .C2({ S25957[538] }),
  .ZN({ S9318 })
);
NAND3_X1 #() 
NAND3_X1_790_ (
  .A1({ S9318 }),
  .A2({ S9316 }),
  .A3({ S25957[541] }),
  .ZN({ S9319 })
);
AOI21_X1 #() 
AOI21_X1_408_ (
  .A({ S7386 }),
  .B1({ S25957[537] }),
  .B2({ S25957[539] }),
  .ZN({ S9321 })
);
AOI21_X1 #() 
AOI21_X1_409_ (
  .A({ S25957[540] }),
  .B1({ S9065 }),
  .B2({ S15 }),
  .ZN({ S9322 })
);
NAND2_X1 #() 
NAND2_X1_691_ (
  .A1({ S9322 }),
  .A2({ S9321 }),
  .ZN({ S9323 })
);
NOR2_X1 #() 
NOR2_X1_158_ (
  .A1({ S25957[538] }),
  .A2({ S9080 }),
  .ZN({ S9324 })
);
NOR3_X1 #() 
NOR3_X1_22_ (
  .A1({ S9107 }),
  .A2({ S9324 }),
  .A3({ S15 }),
  .ZN({ S9325 })
);
NOR2_X1 #() 
NOR2_X1_159_ (
  .A1({ S9066 }),
  .A2({ S9144 }),
  .ZN({ S9326 })
);
NAND2_X1 #() 
NAND2_X1_692_ (
  .A1({ S9326 }),
  .A2({ S9139 }),
  .ZN({ S9327 })
);
NAND2_X1 #() 
NAND2_X1_693_ (
  .A1({ S9327 }),
  .A2({ S25957[540] }),
  .ZN({ S9328 })
);
OAI21_X1 #() 
OAI21_X1_385_ (
  .A({ S9323 }),
  .B1({ S9325 }),
  .B2({ S9328 }),
  .ZN({ S9329 })
);
NAND2_X1 #() 
NAND2_X1_694_ (
  .A1({ S9329 }),
  .A2({ S9099 }),
  .ZN({ S9330 })
);
AOI21_X1 #() 
AOI21_X1_410_ (
  .A({ S25957[542] }),
  .B1({ S9330 }),
  .B2({ S9319 }),
  .ZN({ S9332 })
);
OAI21_X1 #() 
OAI21_X1_386_ (
  .A({ S7026 }),
  .B1({ S9332 }),
  .B2({ S9314 }),
  .ZN({ S9333 })
);
AOI21_X1 #() 
AOI21_X1_411_ (
  .A({ S6418 }),
  .B1({ S9297 }),
  .B2({ S9333 }),
  .ZN({ S9334 })
);
NAND3_X1 #() 
NAND3_X1_791_ (
  .A1({ S9297 }),
  .A2({ S9333 }),
  .A3({ S6418 }),
  .ZN({ S9335 })
);
INV_X1 #() 
INV_X1_242_ (
  .A({ S9335 }),
  .ZN({ S9336 })
);
OAI21_X1 #() 
OAI21_X1_387_ (
  .A({ S5494 }),
  .B1({ S9336 }),
  .B2({ S9334 }),
  .ZN({ S9337 })
);
INV_X1 #() 
INV_X1_243_ (
  .A({ S9334 }),
  .ZN({ S9338 })
);
NAND3_X1 #() 
NAND3_X1_792_ (
  .A1({ S9338 }),
  .A2({ S9335 }),
  .A3({ S25957[645] }),
  .ZN({ S9339 })
);
NAND2_X1 #() 
NAND2_X1_695_ (
  .A1({ S9337 }),
  .A2({ S9339 }),
  .ZN({ S25957[389] })
);
XNOR2_X1 #() 
XNOR2_X1_22_ (
  .A({ S6573 }),
  .B({ S25957[836] }),
  .ZN({ S25957[580] })
);
XNOR2_X1 #() 
XNOR2_X1_23_ (
  .A({ S25957[580] }),
  .B({ S6509 }),
  .ZN({ S25957[548] })
);
NAND2_X1 #() 
NAND2_X1_696_ (
  .A1({ S3843 }),
  .A2({ S3844 }),
  .ZN({ S9341 })
);
INV_X1 #() 
INV_X1_244_ (
  .A({ S9341 }),
  .ZN({ S25957[708] })
);
OAI21_X1 #() 
OAI21_X1_388_ (
  .A({ S15 }),
  .B1({ S9058 }),
  .B2({ S9051 }),
  .ZN({ S9342 })
);
OAI21_X1 #() 
OAI21_X1_389_ (
  .A({ S25957[539] }),
  .B1({ S9282 }),
  .B2({ S9100 }),
  .ZN({ S9343 })
);
OAI211_X1 #() 
OAI211_X1_212_ (
  .A({ S9343 }),
  .B({ S25957[540] }),
  .C1({ S9050 }),
  .C2({ S9342 }),
  .ZN({ S9344 })
);
OAI21_X1 #() 
OAI21_X1_390_ (
  .A({ S15 }),
  .B1({ S9200 }),
  .B2({ S9104 }),
  .ZN({ S9345 })
);
AND2_X1 #() 
AND2_X1_44_ (
  .A1({ S9080 }),
  .A2({ S9051 }),
  .ZN({ S9346 })
);
OAI21_X1 #() 
OAI21_X1_391_ (
  .A({ S25957[539] }),
  .B1({ S9100 }),
  .B2({ S9346 }),
  .ZN({ S9347 })
);
NAND3_X1 #() 
NAND3_X1_793_ (
  .A1({ S9345 }),
  .A2({ S9063 }),
  .A3({ S9347 }),
  .ZN({ S9348 })
);
AOI21_X1 #() 
AOI21_X1_412_ (
  .A({ S25957[539] }),
  .B1({ S7555 }),
  .B2({ S7558 }),
  .ZN({ S9350 })
);
OAI22_X1 #() 
OAI22_X1_18_ (
  .A1({ S9058 }),
  .A2({ S25957[538] }),
  .B1({ S9350 }),
  .B2({ S9080 }),
  .ZN({ S9351 })
);
AOI21_X1 #() 
AOI21_X1_413_ (
  .A({ S9099 }),
  .B1({ S9351 }),
  .B2({ S25957[540] }),
  .ZN({ S9352 })
);
NAND4_X1 #() 
NAND4_X1_80_ (
  .A1({ S25957[537] }),
  .A2({ S7386 }),
  .A3({ S7555 }),
  .A4({ S7558 }),
  .ZN({ S9353 })
);
NAND2_X1 #() 
NAND2_X1_697_ (
  .A1({ S9058 }),
  .A2({ S9051 }),
  .ZN({ S9354 })
);
AOI21_X1 #() 
AOI21_X1_414_ (
  .A({ S25957[539] }),
  .B1({ S9354 }),
  .B2({ S9353 }),
  .ZN({ S9355 })
);
INV_X1 #() 
INV_X1_245_ (
  .A({ S9355 }),
  .ZN({ S9356 })
);
AOI21_X1 #() 
AOI21_X1_415_ (
  .A({ S25957[540] }),
  .B1({ S9280 }),
  .B2({ S9078 }),
  .ZN({ S9357 })
);
AOI21_X1 #() 
AOI21_X1_416_ (
  .A({ S25957[541] }),
  .B1({ S9356 }),
  .B2({ S9357 }),
  .ZN({ S9358 })
);
AOI22_X1 #() 
AOI22_X1_71_ (
  .A1({ S9358 }),
  .A2({ S9344 }),
  .B1({ S9348 }),
  .B2({ S9352 }),
  .ZN({ S9359 })
);
NAND2_X1 #() 
NAND2_X1_698_ (
  .A1({ S9359 }),
  .A2({ S7106 }),
  .ZN({ S9361 })
);
INV_X1 #() 
INV_X1_246_ (
  .A({ S9210 }),
  .ZN({ S9362 })
);
NOR2_X1 #() 
NOR2_X1_160_ (
  .A1({ S9283 }),
  .A2({ S9063 }),
  .ZN({ S9363 })
);
NAND3_X1 #() 
NAND3_X1_794_ (
  .A1({ S9281 }),
  .A2({ S15 }),
  .A3({ S9071 }),
  .ZN({ S9364 })
);
AOI21_X1 #() 
AOI21_X1_417_ (
  .A({ S25957[540] }),
  .B1({ S9114 }),
  .B2({ S9080 }),
  .ZN({ S9365 })
);
AOI22_X1 #() 
AOI22_X1_72_ (
  .A1({ S9363 }),
  .A2({ S9362 }),
  .B1({ S9364 }),
  .B2({ S9365 }),
  .ZN({ S9366 })
);
OAI21_X1 #() 
OAI21_X1_392_ (
  .A({ S15 }),
  .B1({ S23 }),
  .B2({ S9051 }),
  .ZN({ S9367 })
);
OAI211_X1 #() 
OAI211_X1_213_ (
  .A({ S9367 }),
  .B({ S25957[540] }),
  .C1({ S15 }),
  .C2({ S9081 }),
  .ZN({ S9368 })
);
NAND3_X1 #() 
NAND3_X1_795_ (
  .A1({ S9076 }),
  .A2({ S15 }),
  .A3({ S7386 }),
  .ZN({ S9369 })
);
OAI21_X1 #() 
OAI21_X1_393_ (
  .A({ S9369 }),
  .B1({ S9282 }),
  .B2({ S9079 }),
  .ZN({ S9370 })
);
OAI21_X1 #() 
OAI21_X1_394_ (
  .A({ S9368 }),
  .B1({ S9370 }),
  .B2({ S25957[540] }),
  .ZN({ S9372 })
);
NAND2_X1 #() 
NAND2_X1_699_ (
  .A1({ S9372 }),
  .A2({ S25957[541] }),
  .ZN({ S9373 })
);
OAI21_X1 #() 
OAI21_X1_395_ (
  .A({ S9373 }),
  .B1({ S9366 }),
  .B2({ S25957[541] }),
  .ZN({ S9374 })
);
NAND2_X1 #() 
NAND2_X1_700_ (
  .A1({ S9374 }),
  .A2({ S25957[542] }),
  .ZN({ S9375 })
);
NAND3_X1 #() 
NAND3_X1_796_ (
  .A1({ S9375 }),
  .A2({ S9361 }),
  .A3({ S25957[543] }),
  .ZN({ S9376 })
);
OAI21_X1 #() 
OAI21_X1_396_ (
  .A({ S9167 }),
  .B1({ S9146 }),
  .B2({ S9208 }),
  .ZN({ S9377 })
);
OAI21_X1 #() 
OAI21_X1_397_ (
  .A({ S9078 }),
  .B1({ S25957[538] }),
  .B2({ S22 }),
  .ZN({ S9378 })
);
INV_X1 #() 
INV_X1_247_ (
  .A({ S9378 }),
  .ZN({ S9379 })
);
AND2_X1 #() 
AND2_X1_45_ (
  .A1({ S9063 }),
  .A2({ S9112 }),
  .ZN({ S9380 })
);
OAI21_X1 #() 
OAI21_X1_398_ (
  .A({ S9380 }),
  .B1({ S9379 }),
  .B2({ S25957[539] }),
  .ZN({ S9381 })
);
NAND2_X1 #() 
NAND2_X1_701_ (
  .A1({ S9381 }),
  .A2({ S9377 }),
  .ZN({ S9383 })
);
INV_X1 #() 
INV_X1_248_ (
  .A({ S142 }),
  .ZN({ S9384 })
);
OAI21_X1 #() 
OAI21_X1_399_ (
  .A({ S25957[540] }),
  .B1({ S25957[538] }),
  .B2({ S9384 }),
  .ZN({ S9385 })
);
OAI211_X1 #() 
OAI211_X1_214_ (
  .A({ S9063 }),
  .B({ S9308 }),
  .C1({ S9200 }),
  .C2({ S9342 }),
  .ZN({ S9386 })
);
NAND3_X1 #() 
NAND3_X1_797_ (
  .A1({ S9386 }),
  .A2({ S25957[541] }),
  .A3({ S9385 }),
  .ZN({ S9387 })
);
OAI21_X1 #() 
OAI21_X1_400_ (
  .A({ S9387 }),
  .B1({ S9383 }),
  .B2({ S25957[541] }),
  .ZN({ S9388 })
);
NAND2_X1 #() 
NAND2_X1_702_ (
  .A1({ S9388 }),
  .A2({ S25957[542] }),
  .ZN({ S9389 })
);
AND2_X1 #() 
AND2_X1_46_ (
  .A1({ S9291 }),
  .A2({ S9288 }),
  .ZN({ S9390 })
);
AOI21_X1 #() 
AOI21_X1_418_ (
  .A({ S9063 }),
  .B1({ S9272 }),
  .B2({ S25957[538] }),
  .ZN({ S9391 })
);
AOI21_X1 #() 
AOI21_X1_419_ (
  .A({ S9099 }),
  .B1({ S9069 }),
  .B2({ S9391 }),
  .ZN({ S9392 })
);
OAI21_X1 #() 
OAI21_X1_401_ (
  .A({ S9392 }),
  .B1({ S25957[540] }),
  .B2({ S9390 }),
  .ZN({ S9394 })
);
NAND3_X1 #() 
NAND3_X1_798_ (
  .A1({ S9129 }),
  .A2({ S9076 }),
  .A3({ S9090 }),
  .ZN({ S9395 })
);
NAND3_X1 #() 
NAND3_X1_799_ (
  .A1({ S9078 }),
  .A2({ S23 }),
  .A3({ S25957[539] }),
  .ZN({ S9396 })
);
AND2_X1 #() 
AND2_X1_47_ (
  .A1({ S9395 }),
  .A2({ S9396 }),
  .ZN({ S9397 })
);
OAI21_X1 #() 
OAI21_X1_402_ (
  .A({ S25957[540] }),
  .B1({ S9282 }),
  .B2({ S9134 }),
  .ZN({ S9398 })
);
AOI21_X1 #() 
AOI21_X1_420_ (
  .A({ S15 }),
  .B1({ S9067 }),
  .B2({ S9071 }),
  .ZN({ S9399 })
);
OAI221_X1 #() 
OAI221_X1_15_ (
  .A({ S9099 }),
  .B1({ S9398 }),
  .B2({ S9399 }),
  .C1({ S9397 }),
  .C2({ S25957[540] }),
  .ZN({ S9400 })
);
NAND3_X1 #() 
NAND3_X1_800_ (
  .A1({ S9400 }),
  .A2({ S7106 }),
  .A3({ S9394 }),
  .ZN({ S9401 })
);
NAND2_X1 #() 
NAND2_X1_703_ (
  .A1({ S9401 }),
  .A2({ S9389 }),
  .ZN({ S9402 })
);
NAND2_X1 #() 
NAND2_X1_704_ (
  .A1({ S9402 }),
  .A2({ S7026 }),
  .ZN({ S9403 })
);
NAND3_X1 #() 
NAND3_X1_801_ (
  .A1({ S9403 }),
  .A2({ S25957[708] }),
  .A3({ S9376 }),
  .ZN({ S9405 })
);
NAND3_X1 #() 
NAND3_X1_802_ (
  .A1({ S9401 }),
  .A2({ S9389 }),
  .A3({ S7026 }),
  .ZN({ S9406 })
);
OAI211_X1 #() 
OAI211_X1_215_ (
  .A({ S9373 }),
  .B({ S25957[542] }),
  .C1({ S9366 }),
  .C2({ S25957[541] }),
  .ZN({ S9407 })
);
OAI211_X1 #() 
OAI211_X1_216_ (
  .A({ S9407 }),
  .B({ S25957[543] }),
  .C1({ S25957[542] }),
  .C2({ S9359 }),
  .ZN({ S9408 })
);
NAND3_X1 #() 
NAND3_X1_803_ (
  .A1({ S9408 }),
  .A2({ S9406 }),
  .A3({ S9341 }),
  .ZN({ S9409 })
);
AOI21_X1 #() 
AOI21_X1_421_ (
  .A({ S25957[644] }),
  .B1({ S9405 }),
  .B2({ S9409 }),
  .ZN({ S9410 })
);
AOI21_X1 #() 
AOI21_X1_422_ (
  .A({ S9341 }),
  .B1({ S9408 }),
  .B2({ S9406 }),
  .ZN({ S9411 })
);
INV_X1 #() 
INV_X1_249_ (
  .A({ S9409 }),
  .ZN({ S9412 })
);
NOR3_X1 #() 
NOR3_X1_23_ (
  .A1({ S9412 }),
  .A2({ S9411 }),
  .A3({ S5495 }),
  .ZN({ S9413 })
);
NOR2_X1 #() 
NOR2_X1_161_ (
  .A1({ S9413 }),
  .A2({ S9410 }),
  .ZN({ S25957[388] })
);
NOR2_X1 #() 
NOR2_X1_162_ (
  .A1({ S3925 }),
  .A2({ S3921 }),
  .ZN({ S25957[675] })
);
INV_X1 #() 
INV_X1_250_ (
  .A({ S25957[675] }),
  .ZN({ S9415 })
);
NOR2_X1 #() 
NOR2_X1_163_ (
  .A1({ S6642 }),
  .A2({ S6646 }),
  .ZN({ S25957[579] })
);
XNOR2_X1 #() 
XNOR2_X1_24_ (
  .A({ S25957[579] }),
  .B({ S9415 }),
  .ZN({ S25957[547] })
);
AOI21_X1 #() 
AOI21_X1_423_ (
  .A({ S15 }),
  .B1({ S9081 }),
  .B2({ S9078 }),
  .ZN({ S9416 })
);
NAND2_X1 #() 
NAND2_X1_705_ (
  .A1({ S9051 }),
  .A2({ S15 }),
  .ZN({ S9417 })
);
AOI22_X1 #() 
AOI22_X1_73_ (
  .A1({ S9417 }),
  .A2({ S9288 }),
  .B1({ S9080 }),
  .B2({ S9051 }),
  .ZN({ S9418 })
);
OAI21_X1 #() 
OAI21_X1_403_ (
  .A({ S9063 }),
  .B1({ S9418 }),
  .B2({ S9416 }),
  .ZN({ S9419 })
);
NAND3_X1 #() 
NAND3_X1_804_ (
  .A1({ S9049 }),
  .A2({ S15 }),
  .A3({ S9078 }),
  .ZN({ S9420 })
);
NOR2_X1 #() 
NOR2_X1_164_ (
  .A1({ S9420 }),
  .A2({ S9063 }),
  .ZN({ S9421 })
);
NOR2_X1 #() 
NOR2_X1_165_ (
  .A1({ S9421 }),
  .A2({ S25957[541] }),
  .ZN({ S9423 })
);
NAND2_X1 #() 
NAND2_X1_706_ (
  .A1({ S9419 }),
  .A2({ S9423 }),
  .ZN({ S9424 })
);
NAND2_X1 #() 
NAND2_X1_707_ (
  .A1({ S9079 }),
  .A2({ S9121 }),
  .ZN({ S9425 })
);
AOI21_X1 #() 
AOI21_X1_424_ (
  .A({ S9063 }),
  .B1({ S9425 }),
  .B2({ S9057 }),
  .ZN({ S9426 })
);
NAND3_X1 #() 
NAND3_X1_805_ (
  .A1({ S9076 }),
  .A2({ S15 }),
  .A3({ S9080 }),
  .ZN({ S9427 })
);
INV_X1 #() 
INV_X1_251_ (
  .A({ S9131 }),
  .ZN({ S9428 })
);
AOI21_X1 #() 
AOI21_X1_425_ (
  .A({ S25957[540] }),
  .B1({ S9065 }),
  .B2({ S9428 }),
  .ZN({ S9429 })
);
AOI22_X1 #() 
AOI22_X1_74_ (
  .A1({ S9426 }),
  .A2({ S9102 }),
  .B1({ S9427 }),
  .B2({ S9429 }),
  .ZN({ S9430 })
);
OAI211_X1 #() 
OAI211_X1_217_ (
  .A({ S9424 }),
  .B({ S25957[542] }),
  .C1({ S9430 }),
  .C2({ S9099 }),
  .ZN({ S9431 })
);
NAND2_X1 #() 
NAND2_X1_708_ (
  .A1({ S9065 }),
  .A2({ S15 }),
  .ZN({ S9432 })
);
NAND4_X1 #() 
NAND4_X1_81_ (
  .A1({ S9058 }),
  .A2({ S9078 }),
  .A3({ S9080 }),
  .A4({ S25957[539] }),
  .ZN({ S9434 })
);
OAI211_X1 #() 
OAI211_X1_218_ (
  .A({ S9434 }),
  .B({ S25957[540] }),
  .C1({ S9432 }),
  .C2({ S9324 }),
  .ZN({ S9435 })
);
AOI22_X1 #() 
AOI22_X1_75_ (
  .A1({ S9378 }),
  .A2({ S25957[539] }),
  .B1({ S9089 }),
  .B2({ S9090 }),
  .ZN({ S9436 })
);
OAI211_X1 #() 
OAI211_X1_219_ (
  .A({ S9099 }),
  .B({ S9435 }),
  .C1({ S9436 }),
  .C2({ S25957[540] }),
  .ZN({ S9437 })
);
AOI21_X1 #() 
AOI21_X1_426_ (
  .A({ S9228 }),
  .B1({ S9106 }),
  .B2({ S15 }),
  .ZN({ S9438 })
);
NAND3_X1 #() 
NAND3_X1_806_ (
  .A1({ S9078 }),
  .A2({ S9080 }),
  .A3({ S15 }),
  .ZN({ S9439 })
);
NAND2_X1 #() 
NAND2_X1_709_ (
  .A1({ S9205 }),
  .A2({ S9439 }),
  .ZN({ S9440 })
);
AOI21_X1 #() 
AOI21_X1_427_ (
  .A({ S9099 }),
  .B1({ S9440 }),
  .B2({ S9063 }),
  .ZN({ S9441 })
);
OAI21_X1 #() 
OAI21_X1_404_ (
  .A({ S9441 }),
  .B1({ S9438 }),
  .B2({ S9063 }),
  .ZN({ S9442 })
);
NAND3_X1 #() 
NAND3_X1_807_ (
  .A1({ S9437 }),
  .A2({ S9442 }),
  .A3({ S7106 }),
  .ZN({ S9443 })
);
NAND3_X1 #() 
NAND3_X1_808_ (
  .A1({ S9431 }),
  .A2({ S9443 }),
  .A3({ S7026 }),
  .ZN({ S9445 })
);
OAI211_X1 #() 
OAI211_X1_220_ (
  .A({ S25957[540] }),
  .B({ S9396 }),
  .C1({ S9342 }),
  .C2({ S9066 }),
  .ZN({ S9446 })
);
INV_X1 #() 
INV_X1_252_ (
  .A({ S9199 }),
  .ZN({ S9447 })
);
AOI21_X1 #() 
AOI21_X1_428_ (
  .A({ S15 }),
  .B1({ S9057 }),
  .B2({ S25957[537] }),
  .ZN({ S9448 })
);
NAND2_X1 #() 
NAND2_X1_710_ (
  .A1({ S9169 }),
  .A2({ S9078 }),
  .ZN({ S9449 })
);
AOI22_X1 #() 
AOI22_X1_76_ (
  .A1({ S9449 }),
  .A2({ S9448 }),
  .B1({ S9447 }),
  .B2({ S9326 }),
  .ZN({ S9450 })
);
OAI211_X1 #() 
OAI211_X1_221_ (
  .A({ S25957[541] }),
  .B({ S9446 }),
  .C1({ S9450 }),
  .C2({ S25957[540] }),
  .ZN({ S9451 })
);
NAND3_X1 #() 
NAND3_X1_809_ (
  .A1({ S9106 }),
  .A2({ S9067 }),
  .A3({ S15 }),
  .ZN({ S9452 })
);
NAND2_X1 #() 
NAND2_X1_711_ (
  .A1({ S9452 }),
  .A2({ S9274 }),
  .ZN({ S9453 })
);
NAND2_X1 #() 
NAND2_X1_712_ (
  .A1({ S9453 }),
  .A2({ S25957[540] }),
  .ZN({ S9454 })
);
AND2_X1 #() 
AND2_X1_48_ (
  .A1({ S9380 }),
  .A2({ S9143 }),
  .ZN({ S9456 })
);
NOR2_X1 #() 
NOR2_X1_166_ (
  .A1({ S9456 }),
  .A2({ S25957[541] }),
  .ZN({ S9457 })
);
NAND2_X1 #() 
NAND2_X1_713_ (
  .A1({ S9454 }),
  .A2({ S9457 }),
  .ZN({ S9458 })
);
NAND3_X1 #() 
NAND3_X1_810_ (
  .A1({ S9458 }),
  .A2({ S25957[542] }),
  .A3({ S9451 }),
  .ZN({ S9459 })
);
NAND3_X1 #() 
NAND3_X1_811_ (
  .A1({ S9106 }),
  .A2({ S25957[539] }),
  .A3({ S9281 }),
  .ZN({ S9460 })
);
AOI21_X1 #() 
AOI21_X1_429_ (
  .A({ S25957[540] }),
  .B1({ S9272 }),
  .B2({ S9078 }),
  .ZN({ S9461 })
);
NAND2_X1 #() 
NAND2_X1_714_ (
  .A1({ S9460 }),
  .A2({ S9461 }),
  .ZN({ S9462 })
);
NAND2_X1 #() 
NAND2_X1_715_ (
  .A1({ S9087 }),
  .A2({ S25957[539] }),
  .ZN({ S9463 })
);
NAND3_X1 #() 
NAND3_X1_812_ (
  .A1({ S9463 }),
  .A2({ S25957[540] }),
  .A3({ S9364 }),
  .ZN({ S9464 })
);
NAND3_X1 #() 
NAND3_X1_813_ (
  .A1({ S9462 }),
  .A2({ S9464 }),
  .A3({ S9099 }),
  .ZN({ S9465 })
);
AOI21_X1 #() 
AOI21_X1_430_ (
  .A({ S15 }),
  .B1({ S7464 }),
  .B2({ S7467 }),
  .ZN({ S9467 })
);
NAND3_X1 #() 
NAND3_X1_814_ (
  .A1({ S9238 }),
  .A2({ S9467 }),
  .A3({ S9071 }),
  .ZN({ S9468 })
);
OAI211_X1 #() 
OAI211_X1_222_ (
  .A({ S9063 }),
  .B({ S9468 }),
  .C1({ S9248 }),
  .C2({ S9146 }),
  .ZN({ S9469 })
);
OAI21_X1 #() 
OAI21_X1_405_ (
  .A({ S25957[539] }),
  .B1({ S23 }),
  .B2({ S9051 }),
  .ZN({ S9470 })
);
OAI211_X1 #() 
OAI211_X1_223_ (
  .A({ S9057 }),
  .B({ S15 }),
  .C1({ S9051 }),
  .C2({ S9080 }),
  .ZN({ S9471 })
);
OAI211_X1 #() 
OAI211_X1_224_ (
  .A({ S9471 }),
  .B({ S25957[540] }),
  .C1({ S9158 }),
  .C2({ S9470 }),
  .ZN({ S9472 })
);
NAND3_X1 #() 
NAND3_X1_815_ (
  .A1({ S9472 }),
  .A2({ S9469 }),
  .A3({ S25957[541] }),
  .ZN({ S9473 })
);
NAND3_X1 #() 
NAND3_X1_816_ (
  .A1({ S9465 }),
  .A2({ S9473 }),
  .A3({ S7106 }),
  .ZN({ S9474 })
);
NAND3_X1 #() 
NAND3_X1_817_ (
  .A1({ S9459 }),
  .A2({ S25957[543] }),
  .A3({ S9474 }),
  .ZN({ S9475 })
);
AOI21_X1 #() 
AOI21_X1_431_ (
  .A({ S25957[707] }),
  .B1({ S9475 }),
  .B2({ S9445 }),
  .ZN({ S9476 })
);
NAND2_X1 #() 
NAND2_X1_716_ (
  .A1({ S9465 }),
  .A2({ S9473 }),
  .ZN({ S9478 })
);
NAND2_X1 #() 
NAND2_X1_717_ (
  .A1({ S9478 }),
  .A2({ S7106 }),
  .ZN({ S9479 })
);
NAND2_X1 #() 
NAND2_X1_718_ (
  .A1({ S9300 }),
  .A2({ S25957[539] }),
  .ZN({ S9480 })
);
OAI211_X1 #() 
OAI211_X1_225_ (
  .A({ S25957[540] }),
  .B({ S9480 }),
  .C1({ S9145 }),
  .C2({ S25957[539] }),
  .ZN({ S9481 })
);
NAND3_X1 #() 
NAND3_X1_818_ (
  .A1({ S9449 }),
  .A2({ S9132 }),
  .A3({ S9065 }),
  .ZN({ S9482 })
);
OAI211_X1 #() 
OAI211_X1_226_ (
  .A({ S9482 }),
  .B({ S9063 }),
  .C1({ S9199 }),
  .C2({ S9187 }),
  .ZN({ S9483 })
);
NAND3_X1 #() 
NAND3_X1_819_ (
  .A1({ S9483 }),
  .A2({ S9481 }),
  .A3({ S25957[541] }),
  .ZN({ S9484 })
);
AOI21_X1 #() 
AOI21_X1_432_ (
  .A({ S9456 }),
  .B1({ S9453 }),
  .B2({ S25957[540] }),
  .ZN({ S9485 })
);
OAI211_X1 #() 
OAI211_X1_227_ (
  .A({ S25957[542] }),
  .B({ S9484 }),
  .C1({ S9485 }),
  .C2({ S25957[541] }),
  .ZN({ S9486 })
);
NAND3_X1 #() 
NAND3_X1_820_ (
  .A1({ S9479 }),
  .A2({ S9486 }),
  .A3({ S25957[543] }),
  .ZN({ S9487 })
);
OAI21_X1 #() 
OAI21_X1_406_ (
  .A({ S9434 }),
  .B1({ S9432 }),
  .B2({ S9324 }),
  .ZN({ S9489 })
);
NAND2_X1 #() 
NAND2_X1_719_ (
  .A1({ S9489 }),
  .A2({ S25957[540] }),
  .ZN({ S9490 })
);
NAND2_X1 #() 
NAND2_X1_720_ (
  .A1({ S9378 }),
  .A2({ S25957[539] }),
  .ZN({ S9491 })
);
NAND3_X1 #() 
NAND3_X1_821_ (
  .A1({ S9491 }),
  .A2({ S9063 }),
  .A3({ S9091 }),
  .ZN({ S9492 })
);
NAND3_X1 #() 
NAND3_X1_822_ (
  .A1({ S9490 }),
  .A2({ S9492 }),
  .A3({ S9099 }),
  .ZN({ S9493 })
);
NAND3_X1 #() 
NAND3_X1_823_ (
  .A1({ S9205 }),
  .A2({ S9439 }),
  .A3({ S9063 }),
  .ZN({ S9494 })
);
NAND2_X1 #() 
NAND2_X1_721_ (
  .A1({ S9470 }),
  .A2({ S25957[540] }),
  .ZN({ S9495 })
);
OAI211_X1 #() 
OAI211_X1_228_ (
  .A({ S25957[541] }),
  .B({ S9494 }),
  .C1({ S9109 }),
  .C2({ S9495 }),
  .ZN({ S9496 })
);
NAND3_X1 #() 
NAND3_X1_824_ (
  .A1({ S9493 }),
  .A2({ S9496 }),
  .A3({ S7106 }),
  .ZN({ S9497 })
);
INV_X1 #() 
INV_X1_253_ (
  .A({ S9102 }),
  .ZN({ S9498 })
);
NAND2_X1 #() 
NAND2_X1_722_ (
  .A1({ S9429 }),
  .A2({ S9427 }),
  .ZN({ S9500 })
);
OAI211_X1 #() 
OAI211_X1_229_ (
  .A({ S9500 }),
  .B({ S25957[541] }),
  .C1({ S9498 }),
  .C2({ S9206 }),
  .ZN({ S9501 })
);
NAND2_X1 #() 
NAND2_X1_723_ (
  .A1({ S9417 }),
  .A2({ S9288 }),
  .ZN({ S9502 })
);
NAND2_X1 #() 
NAND2_X1_724_ (
  .A1({ S9502 }),
  .A2({ S9081 }),
  .ZN({ S9503 })
);
AOI21_X1 #() 
AOI21_X1_433_ (
  .A({ S25957[540] }),
  .B1({ S9503 }),
  .B2({ S9137 }),
  .ZN({ S9504 })
);
OAI21_X1 #() 
OAI21_X1_407_ (
  .A({ S9099 }),
  .B1({ S9504 }),
  .B2({ S9421 }),
  .ZN({ S9505 })
);
NAND3_X1 #() 
NAND3_X1_825_ (
  .A1({ S9505 }),
  .A2({ S25957[542] }),
  .A3({ S9501 }),
  .ZN({ S9506 })
);
NAND3_X1 #() 
NAND3_X1_826_ (
  .A1({ S9506 }),
  .A2({ S9497 }),
  .A3({ S7026 }),
  .ZN({ S9507 })
);
AOI21_X1 #() 
AOI21_X1_434_ (
  .A({ S6643 }),
  .B1({ S9487 }),
  .B2({ S9507 }),
  .ZN({ S9508 })
);
OAI21_X1 #() 
OAI21_X1_408_ (
  .A({ S25957[547] }),
  .B1({ S9508 }),
  .B2({ S9476 }),
  .ZN({ S9509 })
);
INV_X1 #() 
INV_X1_254_ (
  .A({ S25957[547] }),
  .ZN({ S9511 })
);
NAND3_X1 #() 
NAND3_X1_827_ (
  .A1({ S9487 }),
  .A2({ S6643 }),
  .A3({ S9507 }),
  .ZN({ S9512 })
);
NAND3_X1 #() 
NAND3_X1_828_ (
  .A1({ S9475 }),
  .A2({ S25957[707] }),
  .A3({ S9445 }),
  .ZN({ S9513 })
);
NAND3_X1 #() 
NAND3_X1_829_ (
  .A1({ S9512 }),
  .A2({ S9513 }),
  .A3({ S9511 }),
  .ZN({ S9514 })
);
NAND3_X1 #() 
NAND3_X1_830_ (
  .A1({ S9509 }),
  .A2({ S25957[515] }),
  .A3({ S9514 }),
  .ZN({ S9515 })
);
NAND2_X1 #() 
NAND2_X1_725_ (
  .A1({ S6644 }),
  .A2({ S6645 }),
  .ZN({ S25957[611] })
);
NAND3_X1 #() 
NAND3_X1_831_ (
  .A1({ S9487 }),
  .A2({ S25957[611] }),
  .A3({ S9507 }),
  .ZN({ S9516 })
);
INV_X1 #() 
INV_X1_255_ (
  .A({ S25957[611] }),
  .ZN({ S9517 })
);
NAND3_X1 #() 
NAND3_X1_832_ (
  .A1({ S9475 }),
  .A2({ S9517 }),
  .A3({ S9445 }),
  .ZN({ S9518 })
);
NAND3_X1 #() 
NAND3_X1_833_ (
  .A1({ S9516 }),
  .A2({ S9518 }),
  .A3({ S9415 }),
  .ZN({ S9519 })
);
NAND3_X1 #() 
NAND3_X1_834_ (
  .A1({ S9487 }),
  .A2({ S9517 }),
  .A3({ S9507 }),
  .ZN({ S9521 })
);
NAND3_X1 #() 
NAND3_X1_835_ (
  .A1({ S9475 }),
  .A2({ S25957[611] }),
  .A3({ S9445 }),
  .ZN({ S9522 })
);
NAND3_X1 #() 
NAND3_X1_836_ (
  .A1({ S9521 }),
  .A2({ S9522 }),
  .A3({ S25957[675] }),
  .ZN({ S9523 })
);
NAND3_X1 #() 
NAND3_X1_837_ (
  .A1({ S9519 }),
  .A2({ S9523 }),
  .A3({ S12 }),
  .ZN({ S9524 })
);
NAND2_X1 #() 
NAND2_X1_726_ (
  .A1({ S9515 }),
  .A2({ S9524 }),
  .ZN({ S24 })
);
AOI21_X1 #() 
AOI21_X1_435_ (
  .A({ S12 }),
  .B1({ S9519 }),
  .B2({ S9523 }),
  .ZN({ S9525 })
);
AND3_X1 #() 
AND3_X1_33_ (
  .A1({ S9523 }),
  .A2({ S9519 }),
  .A3({ S12 }),
  .ZN({ S9526 })
);
NOR2_X1 #() 
NOR2_X1_167_ (
  .A1({ S9526 }),
  .A2({ S9525 }),
  .ZN({ S25957[387] })
);
NAND3_X1 #() 
NAND3_X1_838_ (
  .A1({ S9301 }),
  .A2({ S25957[540] }),
  .A3({ S9396 }),
  .ZN({ S9527 })
);
NAND3_X1 #() 
NAND3_X1_839_ (
  .A1({ S9327 }),
  .A2({ S9211 }),
  .A3({ S9063 }),
  .ZN({ S9528 })
);
NAND3_X1 #() 
NAND3_X1_840_ (
  .A1({ S9528 }),
  .A2({ S25957[541] }),
  .A3({ S9527 }),
  .ZN({ S9530 })
);
NAND4_X1 #() 
NAND4_X1_82_ (
  .A1({ S9076 }),
  .A2({ S9058 }),
  .A3({ S25957[539] }),
  .A4({ S9080 }),
  .ZN({ S9531 })
);
OAI21_X1 #() 
OAI21_X1_409_ (
  .A({ S15 }),
  .B1({ S9324 }),
  .B2({ S9052 }),
  .ZN({ S9532 })
);
NAND3_X1 #() 
NAND3_X1_841_ (
  .A1({ S9532 }),
  .A2({ S9063 }),
  .A3({ S9531 }),
  .ZN({ S9533 })
);
AOI21_X1 #() 
AOI21_X1_436_ (
  .A({ S9063 }),
  .B1({ S9169 }),
  .B2({ S9350 }),
  .ZN({ S9534 })
);
NAND3_X1 #() 
NAND3_X1_842_ (
  .A1({ S9463 }),
  .A2({ S9193 }),
  .A3({ S9534 }),
  .ZN({ S9535 })
);
NAND3_X1 #() 
NAND3_X1_843_ (
  .A1({ S9533 }),
  .A2({ S9099 }),
  .A3({ S9535 }),
  .ZN({ S9536 })
);
NAND3_X1 #() 
NAND3_X1_844_ (
  .A1({ S9536 }),
  .A2({ S9530 }),
  .A3({ S7106 }),
  .ZN({ S9537 })
);
NOR2_X1 #() 
NOR2_X1_168_ (
  .A1({ S9139 }),
  .A2({ S25957[540] }),
  .ZN({ S9538 })
);
AOI21_X1 #() 
AOI21_X1_437_ (
  .A({ S15 }),
  .B1({ S9049 }),
  .B2({ S9051 }),
  .ZN({ S9539 })
);
NAND2_X1 #() 
NAND2_X1_727_ (
  .A1({ S9539 }),
  .A2({ S9106 }),
  .ZN({ S9541 })
);
AOI21_X1 #() 
AOI21_X1_438_ (
  .A({ S9063 }),
  .B1({ S9272 }),
  .B2({ S9071 }),
  .ZN({ S9542 })
);
AOI22_X1 #() 
AOI22_X1_77_ (
  .A1({ S9538 }),
  .A2({ S9235 }),
  .B1({ S9541 }),
  .B2({ S9542 }),
  .ZN({ S9543 })
);
OAI211_X1 #() 
OAI211_X1_230_ (
  .A({ S9308 }),
  .B({ S9063 }),
  .C1({ S9146 }),
  .C2({ S9128 }),
  .ZN({ S9544 })
);
INV_X1 #() 
INV_X1_256_ (
  .A({ S9065 }),
  .ZN({ S9545 })
);
OAI211_X1 #() 
OAI211_X1_231_ (
  .A({ S25957[540] }),
  .B({ S9131 }),
  .C1({ S9545 }),
  .C2({ S9233 }),
  .ZN({ S9546 })
);
NAND3_X1 #() 
NAND3_X1_845_ (
  .A1({ S9544 }),
  .A2({ S9546 }),
  .A3({ S9099 }),
  .ZN({ S9547 })
);
OAI211_X1 #() 
OAI211_X1_232_ (
  .A({ S9547 }),
  .B({ S25957[542] }),
  .C1({ S9543 }),
  .C2({ S9099 }),
  .ZN({ S9548 })
);
NAND3_X1 #() 
NAND3_X1_846_ (
  .A1({ S9537 }),
  .A2({ S9548 }),
  .A3({ S7026 }),
  .ZN({ S9549 })
);
NAND3_X1 #() 
NAND3_X1_847_ (
  .A1({ S9065 }),
  .A2({ S15 }),
  .A3({ S7386 }),
  .ZN({ S9550 })
);
NAND2_X1 #() 
NAND2_X1_728_ (
  .A1({ S9420 }),
  .A2({ S9470 }),
  .ZN({ S9552 })
);
AOI21_X1 #() 
AOI21_X1_439_ (
  .A({ S9063 }),
  .B1({ S9552 }),
  .B2({ S9550 }),
  .ZN({ S9553 })
);
INV_X1 #() 
INV_X1_257_ (
  .A({ S9367 }),
  .ZN({ S9554 })
);
NAND2_X1 #() 
NAND2_X1_729_ (
  .A1({ S9144 }),
  .A2({ S25957[539] }),
  .ZN({ S9555 })
);
OAI211_X1 #() 
OAI211_X1_233_ (
  .A({ S9555 }),
  .B({ S9063 }),
  .C1({ S9081 }),
  .C2({ S15 }),
  .ZN({ S9556 })
);
OAI21_X1 #() 
OAI21_X1_410_ (
  .A({ S25957[541] }),
  .B1({ S9556 }),
  .B2({ S9554 }),
  .ZN({ S9557 })
);
OAI21_X1 #() 
OAI21_X1_411_ (
  .A({ S9429 }),
  .B1({ S9219 }),
  .B2({ S25957[539] }),
  .ZN({ S9558 })
);
NAND2_X1 #() 
NAND2_X1_730_ (
  .A1({ S9065 }),
  .A2({ S25957[539] }),
  .ZN({ S9559 })
);
OAI211_X1 #() 
OAI211_X1_234_ (
  .A({ S25957[540] }),
  .B({ S9559 }),
  .C1({ S9158 }),
  .C2({ S25957[539] }),
  .ZN({ S9560 })
);
NAND3_X1 #() 
NAND3_X1_848_ (
  .A1({ S9560 }),
  .A2({ S9558 }),
  .A3({ S9099 }),
  .ZN({ S9561 })
);
OAI211_X1 #() 
OAI211_X1_235_ (
  .A({ S9561 }),
  .B({ S7106 }),
  .C1({ S9553 }),
  .C2({ S9557 }),
  .ZN({ S9563 })
);
NOR2_X1 #() 
NOR2_X1_169_ (
  .A1({ S9144 }),
  .A2({ S9112 }),
  .ZN({ S9564 })
);
INV_X1 #() 
INV_X1_258_ (
  .A({ S9564 }),
  .ZN({ S9565 })
);
NAND3_X1 #() 
NAND3_X1_849_ (
  .A1({ S9395 }),
  .A2({ S9565 }),
  .A3({ S25957[540] }),
  .ZN({ S9566 })
);
NAND2_X1 #() 
NAND2_X1_731_ (
  .A1({ S9566 }),
  .A2({ S25957[541] }),
  .ZN({ S9567 })
);
NAND2_X1 #() 
NAND2_X1_732_ (
  .A1({ S9117 }),
  .A2({ S9152 }),
  .ZN({ S9568 })
);
AOI21_X1 #() 
AOI21_X1_440_ (
  .A({ S25957[540] }),
  .B1({ S9568 }),
  .B2({ S9137 }),
  .ZN({ S9569 })
);
NAND3_X1 #() 
NAND3_X1_850_ (
  .A1({ S9080 }),
  .A2({ S7555 }),
  .A3({ S7558 }),
  .ZN({ S9570 })
);
AOI21_X1 #() 
AOI21_X1_441_ (
  .A({ S25957[539] }),
  .B1({ S9354 }),
  .B2({ S9570 }),
  .ZN({ S9571 })
);
NAND3_X1 #() 
NAND3_X1_851_ (
  .A1({ S9308 }),
  .A2({ S9317 }),
  .A3({ S9063 }),
  .ZN({ S9572 })
);
NAND4_X1 #() 
NAND4_X1_83_ (
  .A1({ S9058 }),
  .A2({ S25957[538] }),
  .A3({ S9080 }),
  .A4({ S25957[539] }),
  .ZN({ S9574 })
);
NAND2_X1 #() 
NAND2_X1_733_ (
  .A1({ S9574 }),
  .A2({ S25957[540] }),
  .ZN({ S9575 })
);
OAI211_X1 #() 
OAI211_X1_236_ (
  .A({ S9572 }),
  .B({ S9099 }),
  .C1({ S9575 }),
  .C2({ S9571 }),
  .ZN({ S9576 })
);
OAI211_X1 #() 
OAI211_X1_237_ (
  .A({ S9576 }),
  .B({ S25957[542] }),
  .C1({ S9567 }),
  .C2({ S9569 }),
  .ZN({ S9577 })
);
NAND3_X1 #() 
NAND3_X1_852_ (
  .A1({ S9577 }),
  .A2({ S9563 }),
  .A3({ S25957[543] }),
  .ZN({ S9578 })
);
AND3_X1 #() 
AND3_X1_34_ (
  .A1({ S9578 }),
  .A2({ S9549 }),
  .A3({ S6655 }),
  .ZN({ S9579 })
);
AOI21_X1 #() 
AOI21_X1_442_ (
  .A({ S6655 }),
  .B1({ S9578 }),
  .B2({ S9549 }),
  .ZN({ S9580 })
);
OAI21_X1 #() 
OAI21_X1_412_ (
  .A({ S5479 }),
  .B1({ S9579 }),
  .B2({ S9580 }),
  .ZN({ S9581 })
);
NAND3_X1 #() 
NAND3_X1_853_ (
  .A1({ S9578 }),
  .A2({ S9549 }),
  .A3({ S6655 }),
  .ZN({ S9582 })
);
NAND3_X1 #() 
NAND3_X1_854_ (
  .A1({ S9536 }),
  .A2({ S9530 }),
  .A3({ S7026 }),
  .ZN({ S9583 })
);
OAI211_X1 #() 
OAI211_X1_238_ (
  .A({ S9561 }),
  .B({ S25957[543] }),
  .C1({ S9553 }),
  .C2({ S9557 }),
  .ZN({ S9585 })
);
NAND2_X1 #() 
NAND2_X1_734_ (
  .A1({ S9583 }),
  .A2({ S9585 }),
  .ZN({ S9586 })
);
NAND2_X1 #() 
NAND2_X1_735_ (
  .A1({ S9586 }),
  .A2({ S7106 }),
  .ZN({ S9587 })
);
OAI21_X1 #() 
OAI21_X1_413_ (
  .A({ S9057 }),
  .B1({ S9049 }),
  .B2({ S9051 }),
  .ZN({ S9588 })
);
AOI21_X1 #() 
AOI21_X1_443_ (
  .A({ S25957[539] }),
  .B1({ S9169 }),
  .B2({ S9078 }),
  .ZN({ S9589 })
);
AOI21_X1 #() 
AOI21_X1_444_ (
  .A({ S9589 }),
  .B1({ S9588 }),
  .B2({ S25957[539] }),
  .ZN({ S9590 })
);
NAND2_X1 #() 
NAND2_X1_736_ (
  .A1({ S25957[538] }),
  .A2({ S9163 }),
  .ZN({ S9591 })
);
NAND3_X1 #() 
NAND3_X1_855_ (
  .A1({ S9058 }),
  .A2({ S15 }),
  .A3({ S9051 }),
  .ZN({ S9592 })
);
OAI211_X1 #() 
OAI211_X1_239_ (
  .A({ S25957[539] }),
  .B({ S25957[536] }),
  .C1({ S9051 }),
  .C2({ S25957[537] }),
  .ZN({ S9593 })
);
NAND4_X1 #() 
NAND4_X1_84_ (
  .A1({ S9593 }),
  .A2({ S9592 }),
  .A3({ S9591 }),
  .A4({ S25957[540] }),
  .ZN({ S9594 })
);
OAI211_X1 #() 
OAI211_X1_240_ (
  .A({ S9099 }),
  .B({ S9594 }),
  .C1({ S9590 }),
  .C2({ S25957[540] }),
  .ZN({ S9596 })
);
NAND2_X1 #() 
NAND2_X1_737_ (
  .A1({ S9235 }),
  .A2({ S9538 }),
  .ZN({ S9597 })
);
AOI21_X1 #() 
AOI21_X1_445_ (
  .A({ S9099 }),
  .B1({ S9541 }),
  .B2({ S9542 }),
  .ZN({ S9598 })
);
NAND2_X1 #() 
NAND2_X1_738_ (
  .A1({ S9598 }),
  .A2({ S9597 }),
  .ZN({ S9599 })
);
AOI21_X1 #() 
AOI21_X1_446_ (
  .A({ S25957[543] }),
  .B1({ S9599 }),
  .B2({ S9596 }),
  .ZN({ S9600 })
);
NOR2_X1 #() 
NOR2_X1_170_ (
  .A1({ S9187 }),
  .A2({ S9112 }),
  .ZN({ S9601 })
);
OAI21_X1 #() 
OAI21_X1_414_ (
  .A({ S25957[540] }),
  .B1({ S9571 }),
  .B2({ S9601 }),
  .ZN({ S9602 })
);
NAND2_X1 #() 
NAND2_X1_739_ (
  .A1({ S9308 }),
  .A2({ S9317 }),
  .ZN({ S9603 })
);
NAND2_X1 #() 
NAND2_X1_740_ (
  .A1({ S9603 }),
  .A2({ S9063 }),
  .ZN({ S9604 })
);
NAND3_X1 #() 
NAND3_X1_856_ (
  .A1({ S9602 }),
  .A2({ S9099 }),
  .A3({ S9604 }),
  .ZN({ S9605 })
);
NAND3_X1 #() 
NAND3_X1_857_ (
  .A1({ S9281 }),
  .A2({ S9065 }),
  .A3({ S9078 }),
  .ZN({ S9607 })
);
AOI21_X1 #() 
AOI21_X1_447_ (
  .A({ S9564 }),
  .B1({ S9607 }),
  .B2({ S9090 }),
  .ZN({ S9608 })
);
OAI211_X1 #() 
OAI211_X1_241_ (
  .A({ S9063 }),
  .B({ S9137 }),
  .C1({ S9158 }),
  .C2({ S9432 }),
  .ZN({ S9609 })
);
OAI211_X1 #() 
OAI211_X1_242_ (
  .A({ S9609 }),
  .B({ S25957[541] }),
  .C1({ S9608 }),
  .C2({ S9063 }),
  .ZN({ S9610 })
);
AOI21_X1 #() 
AOI21_X1_448_ (
  .A({ S7026 }),
  .B1({ S9605 }),
  .B2({ S9610 }),
  .ZN({ S9611 })
);
OAI21_X1 #() 
OAI21_X1_415_ (
  .A({ S25957[542] }),
  .B1({ S9611 }),
  .B2({ S9600 }),
  .ZN({ S9612 })
);
NAND3_X1 #() 
NAND3_X1_858_ (
  .A1({ S9587 }),
  .A2({ S9612 }),
  .A3({ S25957[704] }),
  .ZN({ S9613 })
);
NAND3_X1 #() 
NAND3_X1_859_ (
  .A1({ S9613 }),
  .A2({ S25957[640] }),
  .A3({ S9582 }),
  .ZN({ S9614 })
);
NAND2_X1 #() 
NAND2_X1_741_ (
  .A1({ S9581 }),
  .A2({ S9614 }),
  .ZN({ S25957[384] })
);
NAND2_X1 #() 
NAND2_X1_742_ (
  .A1({ S9189 }),
  .A2({ S9106 }),
  .ZN({ S9615 })
);
INV_X1 #() 
INV_X1_259_ (
  .A({ S9615 }),
  .ZN({ S9617 })
);
NOR2_X1 #() 
NOR2_X1_171_ (
  .A1({ S25957[538] }),
  .A2({ S23 }),
  .ZN({ S9618 })
);
NAND3_X1 #() 
NAND3_X1_860_ (
  .A1({ S9049 }),
  .A2({ S25957[539] }),
  .A3({ S9071 }),
  .ZN({ S9619 })
);
OAI211_X1 #() 
OAI211_X1_243_ (
  .A({ S9063 }),
  .B({ S9619 }),
  .C1({ S9420 }),
  .C2({ S9618 }),
  .ZN({ S9620 })
);
NAND2_X1 #() 
NAND2_X1_743_ (
  .A1({ S9550 }),
  .A2({ S25957[540] }),
  .ZN({ S9621 })
);
OAI211_X1 #() 
OAI211_X1_244_ (
  .A({ S9620 }),
  .B({ S9099 }),
  .C1({ S9617 }),
  .C2({ S9621 }),
  .ZN({ S9622 })
);
AOI21_X1 #() 
AOI21_X1_449_ (
  .A({ S15 }),
  .B1({ S9089 }),
  .B2({ S9101 }),
  .ZN({ S9623 })
);
NAND2_X1 #() 
NAND2_X1_744_ (
  .A1({ S9342 }),
  .A2({ S9063 }),
  .ZN({ S9624 })
);
NAND3_X1 #() 
NAND3_X1_861_ (
  .A1({ S9274 }),
  .A2({ S25957[540] }),
  .A3({ S9072 }),
  .ZN({ S9625 })
);
OAI211_X1 #() 
OAI211_X1_245_ (
  .A({ S9625 }),
  .B({ S25957[541] }),
  .C1({ S9623 }),
  .C2({ S9624 }),
  .ZN({ S9626 })
);
NAND3_X1 #() 
NAND3_X1_862_ (
  .A1({ S9622 }),
  .A2({ S25957[542] }),
  .A3({ S9626 }),
  .ZN({ S9628 })
);
NOR3_X1 #() 
NOR3_X1_24_ (
  .A1({ S9088 }),
  .A2({ S9355 }),
  .A3({ S25957[540] }),
  .ZN({ S9629 })
);
NAND3_X1 #() 
NAND3_X1_863_ (
  .A1({ S9592 }),
  .A2({ S9251 }),
  .A3({ S9591 }),
  .ZN({ S9630 })
);
OAI21_X1 #() 
OAI21_X1_416_ (
  .A({ S9099 }),
  .B1({ S9630 }),
  .B2({ S9063 }),
  .ZN({ S9631 })
);
NAND2_X1 #() 
NAND2_X1_745_ (
  .A1({ S9238 }),
  .A2({ S25957[539] }),
  .ZN({ S9632 })
);
NOR2_X1 #() 
NOR2_X1_172_ (
  .A1({ S9248 }),
  .A2({ S9632 }),
  .ZN({ S9633 })
);
NAND3_X1 #() 
NAND3_X1_864_ (
  .A1({ S9427 }),
  .A2({ S9380 }),
  .A3({ S9555 }),
  .ZN({ S9634 })
);
OAI211_X1 #() 
OAI211_X1_246_ (
  .A({ S25957[541] }),
  .B({ S9634 }),
  .C1({ S9060 }),
  .C2({ S9633 }),
  .ZN({ S9635 })
);
OAI211_X1 #() 
OAI211_X1_247_ (
  .A({ S9635 }),
  .B({ S7106 }),
  .C1({ S9629 }),
  .C2({ S9631 }),
  .ZN({ S9636 })
);
NAND3_X1 #() 
NAND3_X1_865_ (
  .A1({ S9636 }),
  .A2({ S9628 }),
  .A3({ S25957[543] }),
  .ZN({ S9637 })
);
AOI21_X1 #() 
AOI21_X1_450_ (
  .A({ S9063 }),
  .B1({ S9369 }),
  .B2({ S9468 }),
  .ZN({ S9639 })
);
OAI21_X1 #() 
OAI21_X1_417_ (
  .A({ S25957[541] }),
  .B1({ S9083 }),
  .B2({ S9639 }),
  .ZN({ S9640 })
);
NAND2_X1 #() 
NAND2_X1_746_ (
  .A1({ S9167 }),
  .A2({ S9364 }),
  .ZN({ S9641 })
);
OAI21_X1 #() 
OAI21_X1_418_ (
  .A({ S9063 }),
  .B1({ S25957[538] }),
  .B2({ S9113 }),
  .ZN({ S9642 })
);
OAI211_X1 #() 
OAI211_X1_248_ (
  .A({ S9641 }),
  .B({ S9099 }),
  .C1({ S9418 }),
  .C2({ S9642 }),
  .ZN({ S9643 })
);
NAND3_X1 #() 
NAND3_X1_866_ (
  .A1({ S9640 }),
  .A2({ S9643 }),
  .A3({ S7106 }),
  .ZN({ S9644 })
);
NOR2_X1 #() 
NOR2_X1_173_ (
  .A1({ S9367 }),
  .A2({ S9209 }),
  .ZN({ S9645 })
);
NAND2_X1 #() 
NAND2_X1_747_ (
  .A1({ S9434 }),
  .A2({ S25957[540] }),
  .ZN({ S9646 })
);
NAND4_X1 #() 
NAND4_X1_85_ (
  .A1({ S9170 }),
  .A2({ S9078 }),
  .A3({ S9113 }),
  .A4({ S9063 }),
  .ZN({ S9647 })
);
OAI211_X1 #() 
OAI211_X1_249_ (
  .A({ S25957[541] }),
  .B({ S9647 }),
  .C1({ S9646 }),
  .C2({ S9645 }),
  .ZN({ S9648 })
);
NAND4_X1 #() 
NAND4_X1_86_ (
  .A1({ S25957[537] }),
  .A2({ S25957[536] }),
  .A3({ S7555 }),
  .A4({ S7558 }),
  .ZN({ S9650 })
);
NAND3_X1 #() 
NAND3_X1_867_ (
  .A1({ S9170 }),
  .A2({ S9650 }),
  .A3({ S15 }),
  .ZN({ S9651 })
);
AND3_X1 #() 
AND3_X1_35_ (
  .A1({ S9541 }),
  .A2({ S25957[540] }),
  .A3({ S9651 }),
  .ZN({ S9652 })
);
NAND3_X1 #() 
NAND3_X1_868_ (
  .A1({ S9244 }),
  .A2({ S9574 }),
  .A3({ S9063 }),
  .ZN({ S9653 })
);
NAND2_X1 #() 
NAND2_X1_748_ (
  .A1({ S9653 }),
  .A2({ S9099 }),
  .ZN({ S9654 })
);
OAI211_X1 #() 
OAI211_X1_250_ (
  .A({ S9648 }),
  .B({ S25957[542] }),
  .C1({ S9652 }),
  .C2({ S9654 }),
  .ZN({ S9655 })
);
NAND3_X1 #() 
NAND3_X1_869_ (
  .A1({ S9644 }),
  .A2({ S9655 }),
  .A3({ S7026 }),
  .ZN({ S9656 })
);
NAND3_X1 #() 
NAND3_X1_870_ (
  .A1({ S9637 }),
  .A2({ S9656 }),
  .A3({ S6817 }),
  .ZN({ S9657 })
);
AOI21_X1 #() 
AOI21_X1_451_ (
  .A({ S9063 }),
  .B1({ S9541 }),
  .B2({ S9651 }),
  .ZN({ S9658 })
);
AND2_X1 #() 
AND2_X1_49_ (
  .A1({ S9244 }),
  .A2({ S9574 }),
  .ZN({ S9659 })
);
OAI21_X1 #() 
OAI21_X1_419_ (
  .A({ S9099 }),
  .B1({ S9659 }),
  .B2({ S25957[540] }),
  .ZN({ S9661 })
);
INV_X1 #() 
INV_X1_260_ (
  .A({ S9079 }),
  .ZN({ S9662 })
);
AOI22_X1 #() 
AOI22_X1_78_ (
  .A1({ S9662 }),
  .A2({ S9326 }),
  .B1({ S9129 }),
  .B2({ S9090 }),
  .ZN({ S9663 })
);
NAND3_X1 #() 
NAND3_X1_871_ (
  .A1({ S9170 }),
  .A2({ S9113 }),
  .A3({ S9078 }),
  .ZN({ S9664 })
);
NAND2_X1 #() 
NAND2_X1_749_ (
  .A1({ S9664 }),
  .A2({ S9063 }),
  .ZN({ S9665 })
);
OAI211_X1 #() 
OAI211_X1_251_ (
  .A({ S9665 }),
  .B({ S25957[541] }),
  .C1({ S9663 }),
  .C2({ S9063 }),
  .ZN({ S9666 })
);
OAI211_X1 #() 
OAI211_X1_252_ (
  .A({ S9666 }),
  .B({ S25957[542] }),
  .C1({ S9661 }),
  .C2({ S9658 }),
  .ZN({ S9667 })
);
OAI21_X1 #() 
OAI21_X1_420_ (
  .A({ S15 }),
  .B1({ S9346 }),
  .B2({ S9104 }),
  .ZN({ S9668 })
);
NAND2_X1 #() 
NAND2_X1_750_ (
  .A1({ S9668 }),
  .A2({ S9063 }),
  .ZN({ S9669 })
);
NAND2_X1 #() 
NAND2_X1_751_ (
  .A1({ S9369 }),
  .A2({ S9468 }),
  .ZN({ S9670 })
);
NAND2_X1 #() 
NAND2_X1_752_ (
  .A1({ S9670 }),
  .A2({ S25957[540] }),
  .ZN({ S9671 })
);
NAND3_X1 #() 
NAND3_X1_872_ (
  .A1({ S9669 }),
  .A2({ S9671 }),
  .A3({ S25957[541] }),
  .ZN({ S9672 })
);
AOI21_X1 #() 
AOI21_X1_452_ (
  .A({ S25957[539] }),
  .B1({ S9076 }),
  .B2({ S9078 }),
  .ZN({ S9673 })
);
OAI22_X1 #() 
OAI22_X1_19_ (
  .A1({ S9418 }),
  .A2({ S9642 }),
  .B1({ S9673 }),
  .B2({ S9166 }),
  .ZN({ S9674 })
);
AOI21_X1 #() 
AOI21_X1_453_ (
  .A({ S25957[542] }),
  .B1({ S9674 }),
  .B2({ S9099 }),
  .ZN({ S9675 })
);
NAND2_X1 #() 
NAND2_X1_753_ (
  .A1({ S9675 }),
  .A2({ S9672 }),
  .ZN({ S9676 })
);
NAND3_X1 #() 
NAND3_X1_873_ (
  .A1({ S9667 }),
  .A2({ S7026 }),
  .A3({ S9676 }),
  .ZN({ S9677 })
);
OAI21_X1 #() 
OAI21_X1_421_ (
  .A({ S25957[540] }),
  .B1({ S9448 }),
  .B2({ S9502 }),
  .ZN({ S9678 })
);
AOI22_X1 #() 
AOI22_X1_79_ (
  .A1({ S9539 }),
  .A2({ S9106 }),
  .B1({ S9353 }),
  .B2({ S15 }),
  .ZN({ S9679 })
);
OAI211_X1 #() 
OAI211_X1_253_ (
  .A({ S9678 }),
  .B({ S25957[541] }),
  .C1({ S9679 }),
  .C2({ S25957[540] }),
  .ZN({ S9680 })
);
NAND4_X1 #() 
NAND4_X1_87_ (
  .A1({ S9170 }),
  .A2({ S9078 }),
  .A3({ S9049 }),
  .A4({ S15 }),
  .ZN({ S9682 })
);
AOI21_X1 #() 
AOI21_X1_454_ (
  .A({ S25957[540] }),
  .B1({ S9132 }),
  .B2({ S9071 }),
  .ZN({ S9683 })
);
AOI21_X1 #() 
AOI21_X1_455_ (
  .A({ S9063 }),
  .B1({ S9117 }),
  .B2({ S7386 }),
  .ZN({ S9684 })
);
AOI22_X1 #() 
AOI22_X1_80_ (
  .A1({ S9684 }),
  .A2({ S9615 }),
  .B1({ S9682 }),
  .B2({ S9683 }),
  .ZN({ S9685 })
);
OAI211_X1 #() 
OAI211_X1_254_ (
  .A({ S9680 }),
  .B({ S25957[542] }),
  .C1({ S25957[541] }),
  .C2({ S9685 }),
  .ZN({ S9686 })
);
OAI21_X1 #() 
OAI21_X1_422_ (
  .A({ S7386 }),
  .B1({ S9051 }),
  .B2({ S25957[537] }),
  .ZN({ S9687 })
);
NOR2_X1 #() 
NOR2_X1_174_ (
  .A1({ S9209 }),
  .A2({ S15 }),
  .ZN({ S9688 })
);
AOI22_X1 #() 
AOI22_X1_81_ (
  .A1({ S9089 }),
  .A2({ S9688 }),
  .B1({ S9687 }),
  .B2({ S15 }),
  .ZN({ S9689 })
);
AOI21_X1 #() 
AOI21_X1_456_ (
  .A({ S15 }),
  .B1({ S9058 }),
  .B2({ S9051 }),
  .ZN({ S9690 })
);
AOI21_X1 #() 
AOI21_X1_457_ (
  .A({ S25957[539] }),
  .B1({ S9065 }),
  .B2({ S23 }),
  .ZN({ S9691 })
);
OAI21_X1 #() 
OAI21_X1_423_ (
  .A({ S9063 }),
  .B1({ S9691 }),
  .B2({ S9690 }),
  .ZN({ S9693 })
);
OAI211_X1 #() 
OAI211_X1_255_ (
  .A({ S9693 }),
  .B({ S25957[541] }),
  .C1({ S9689 }),
  .C2({ S9063 }),
  .ZN({ S9694 })
);
NAND2_X1 #() 
NAND2_X1_754_ (
  .A1({ S9630 }),
  .A2({ S25957[540] }),
  .ZN({ S9695 })
);
OAI21_X1 #() 
OAI21_X1_424_ (
  .A({ S9063 }),
  .B1({ S9088 }),
  .B2({ S9355 }),
  .ZN({ S9696 })
);
NAND3_X1 #() 
NAND3_X1_874_ (
  .A1({ S9696 }),
  .A2({ S9099 }),
  .A3({ S9695 }),
  .ZN({ S9697 })
);
NAND3_X1 #() 
NAND3_X1_875_ (
  .A1({ S9697 }),
  .A2({ S7106 }),
  .A3({ S9694 }),
  .ZN({ S9698 })
);
NAND3_X1 #() 
NAND3_X1_876_ (
  .A1({ S9698 }),
  .A2({ S25957[543] }),
  .A3({ S9686 }),
  .ZN({ S9699 })
);
NAND3_X1 #() 
NAND3_X1_877_ (
  .A1({ S9699 }),
  .A2({ S9677 }),
  .A3({ S25957[705] }),
  .ZN({ S9700 })
);
AOI21_X1 #() 
AOI21_X1_458_ (
  .A({ S5464 }),
  .B1({ S9700 }),
  .B2({ S9657 }),
  .ZN({ S9701 })
);
AND3_X1 #() 
AND3_X1_36_ (
  .A1({ S9700 }),
  .A2({ S9657 }),
  .A3({ S5464 }),
  .ZN({ S9702 })
);
NOR2_X1 #() 
NOR2_X1_175_ (
  .A1({ S9702 }),
  .A2({ S9701 }),
  .ZN({ S25957[385] })
);
NAND2_X1 #() 
NAND2_X1_755_ (
  .A1({ S9122 }),
  .A2({ S9071 }),
  .ZN({ S9704 })
);
NAND2_X1 #() 
NAND2_X1_756_ (
  .A1({ S9568 }),
  .A2({ S9704 }),
  .ZN({ S9705 })
);
NAND2_X1 #() 
NAND2_X1_757_ (
  .A1({ S9705 }),
  .A2({ S25957[540] }),
  .ZN({ S9706 })
);
NAND3_X1 #() 
NAND3_X1_878_ (
  .A1({ S9152 }),
  .A2({ S25957[539] }),
  .A3({ S9570 }),
  .ZN({ S9707 })
);
NAND2_X1 #() 
NAND2_X1_758_ (
  .A1({ S9707 }),
  .A2({ S9292 }),
  .ZN({ S9708 })
);
NAND2_X1 #() 
NAND2_X1_759_ (
  .A1({ S9058 }),
  .A2({ S25957[538] }),
  .ZN({ S9709 })
);
NAND3_X1 #() 
NAND3_X1_879_ (
  .A1({ S9152 }),
  .A2({ S25957[539] }),
  .A3({ S9709 }),
  .ZN({ S9710 })
);
AOI21_X1 #() 
AOI21_X1_459_ (
  .A({ S9099 }),
  .B1({ S9710 }),
  .B2({ S9322 }),
  .ZN({ S9711 })
);
NAND2_X1 #() 
NAND2_X1_760_ (
  .A1({ S9350 }),
  .A2({ S9169 }),
  .ZN({ S9712 })
);
AOI21_X1 #() 
AOI21_X1_460_ (
  .A({ S25957[541] }),
  .B1({ S9365 }),
  .B2({ S9712 }),
  .ZN({ S9714 })
);
AOI22_X1 #() 
AOI22_X1_82_ (
  .A1({ S9706 }),
  .A2({ S9711 }),
  .B1({ S9714 }),
  .B2({ S9708 }),
  .ZN({ S9715 })
);
NOR2_X1 #() 
NOR2_X1_176_ (
  .A1({ S9121 }),
  .A2({ S9209 }),
  .ZN({ S9716 })
);
OAI21_X1 #() 
OAI21_X1_425_ (
  .A({ S25957[540] }),
  .B1({ S9716 }),
  .B2({ S9310 }),
  .ZN({ S9717 })
);
NAND2_X1 #() 
NAND2_X1_761_ (
  .A1({ S9196 }),
  .A2({ S9063 }),
  .ZN({ S9718 })
);
NAND3_X1 #() 
NAND3_X1_880_ (
  .A1({ S9718 }),
  .A2({ S9717 }),
  .A3({ S9099 }),
  .ZN({ S9719 })
);
AOI21_X1 #() 
AOI21_X1_461_ (
  .A({ S9063 }),
  .B1({ S9132 }),
  .B2({ S9078 }),
  .ZN({ S9720 })
);
NAND2_X1 #() 
NAND2_X1_762_ (
  .A1({ S9668 }),
  .A2({ S9720 }),
  .ZN({ S9721 })
);
OAI22_X1 #() 
OAI22_X1_20_ (
  .A1({ S9321 }),
  .A2({ S9144 }),
  .B1({ S9467 }),
  .B2({ S25957[538] }),
  .ZN({ S9722 })
);
AOI21_X1 #() 
AOI21_X1_462_ (
  .A({ S9099 }),
  .B1({ S9722 }),
  .B2({ S9063 }),
  .ZN({ S9723 })
);
NAND2_X1 #() 
NAND2_X1_763_ (
  .A1({ S9723 }),
  .A2({ S9721 }),
  .ZN({ S9725 })
);
NAND3_X1 #() 
NAND3_X1_881_ (
  .A1({ S9725 }),
  .A2({ S7106 }),
  .A3({ S9719 }),
  .ZN({ S9726 })
);
OAI211_X1 #() 
OAI211_X1_256_ (
  .A({ S9726 }),
  .B({ S25957[543] }),
  .C1({ S9715 }),
  .C2({ S7106 }),
  .ZN({ S9727 })
);
OAI211_X1 #() 
OAI211_X1_257_ (
  .A({ S25957[539] }),
  .B({ S9078 }),
  .C1({ S9058 }),
  .C2({ S25957[538] }),
  .ZN({ S9728 })
);
NAND3_X1 #() 
NAND3_X1_882_ (
  .A1({ S9728 }),
  .A2({ S9420 }),
  .A3({ S9591 }),
  .ZN({ S9729 })
);
NAND2_X1 #() 
NAND2_X1_764_ (
  .A1({ S9729 }),
  .A2({ S25957[540] }),
  .ZN({ S9730 })
);
AOI21_X1 #() 
AOI21_X1_463_ (
  .A({ S15 }),
  .B1({ S9238 }),
  .B2({ S25957[537] }),
  .ZN({ S9731 })
);
OAI21_X1 #() 
OAI21_X1_426_ (
  .A({ S9063 }),
  .B1({ S9571 }),
  .B2({ S9731 }),
  .ZN({ S9732 })
);
NAND3_X1 #() 
NAND3_X1_883_ (
  .A1({ S9730 }),
  .A2({ S9732 }),
  .A3({ S9099 }),
  .ZN({ S9733 })
);
NAND3_X1 #() 
NAND3_X1_884_ (
  .A1({ S9076 }),
  .A2({ S15 }),
  .A3({ S25957[536] }),
  .ZN({ S9734 })
);
NAND3_X1 #() 
NAND3_X1_885_ (
  .A1({ S9153 }),
  .A2({ S9063 }),
  .A3({ S9734 }),
  .ZN({ S9736 })
);
AOI21_X1 #() 
AOI21_X1_464_ (
  .A({ S25957[539] }),
  .B1({ S9169 }),
  .B2({ S9051 }),
  .ZN({ S9737 })
);
NAND2_X1 #() 
NAND2_X1_765_ (
  .A1({ S9281 }),
  .A2({ S7386 }),
  .ZN({ S9738 })
);
OAI21_X1 #() 
OAI21_X1_427_ (
  .A({ S9738 }),
  .B1({ S9737 }),
  .B2({ S9280 }),
  .ZN({ S9739 })
);
AOI21_X1 #() 
AOI21_X1_465_ (
  .A({ S9099 }),
  .B1({ S9739 }),
  .B2({ S25957[540] }),
  .ZN({ S9740 })
);
NAND2_X1 #() 
NAND2_X1_766_ (
  .A1({ S9740 }),
  .A2({ S9736 }),
  .ZN({ S9741 })
);
NAND3_X1 #() 
NAND3_X1_886_ (
  .A1({ S9733 }),
  .A2({ S9741 }),
  .A3({ S25957[542] }),
  .ZN({ S9742 })
);
OAI211_X1 #() 
OAI211_X1_258_ (
  .A({ S9063 }),
  .B({ S9195 }),
  .C1({ S9203 }),
  .C2({ S9304 }),
  .ZN({ S9743 })
);
OAI211_X1 #() 
OAI211_X1_259_ (
  .A({ S25957[539] }),
  .B({ S9078 }),
  .C1({ S25957[538] }),
  .C2({ S23 }),
  .ZN({ S9744 })
);
OAI211_X1 #() 
OAI211_X1_260_ (
  .A({ S25957[540] }),
  .B({ S9744 }),
  .C1({ S9248 }),
  .C2({ S9146 }),
  .ZN({ S9745 })
);
NAND3_X1 #() 
NAND3_X1_887_ (
  .A1({ S9745 }),
  .A2({ S9743 }),
  .A3({ S25957[541] }),
  .ZN({ S9747 })
);
AOI21_X1 #() 
AOI21_X1_466_ (
  .A({ S15 }),
  .B1({ S9354 }),
  .B2({ S9353 }),
  .ZN({ S9748 })
);
OAI21_X1 #() 
OAI21_X1_428_ (
  .A({ S9063 }),
  .B1({ S9158 }),
  .B2({ S9432 }),
  .ZN({ S9749 })
);
AOI21_X1 #() 
AOI21_X1_467_ (
  .A({ S9063 }),
  .B1({ S9238 }),
  .B2({ S9467 }),
  .ZN({ S9750 })
);
OAI21_X1 #() 
OAI21_X1_429_ (
  .A({ S9750 }),
  .B1({ S9342 }),
  .B2({ S9050 }),
  .ZN({ S9751 })
);
OAI211_X1 #() 
OAI211_X1_261_ (
  .A({ S9099 }),
  .B({ S9751 }),
  .C1({ S9749 }),
  .C2({ S9748 }),
  .ZN({ S9752 })
);
NAND2_X1 #() 
NAND2_X1_767_ (
  .A1({ S9752 }),
  .A2({ S9747 }),
  .ZN({ S9753 })
);
NAND2_X1 #() 
NAND2_X1_768_ (
  .A1({ S9753 }),
  .A2({ S7106 }),
  .ZN({ S9754 })
);
NAND3_X1 #() 
NAND3_X1_888_ (
  .A1({ S9754 }),
  .A2({ S9742 }),
  .A3({ S7026 }),
  .ZN({ S9755 })
);
AOI21_X1 #() 
AOI21_X1_468_ (
  .A({ S6831 }),
  .B1({ S9755 }),
  .B2({ S9727 }),
  .ZN({ S9756 })
);
OAI211_X1 #() 
OAI211_X1_262_ (
  .A({ S25957[541] }),
  .B({ S9738 }),
  .C1({ S9737 }),
  .C2({ S9280 }),
  .ZN({ S9758 })
);
NAND4_X1 #() 
NAND4_X1_88_ (
  .A1({ S9728 }),
  .A2({ S9591 }),
  .A3({ S9420 }),
  .A4({ S9099 }),
  .ZN({ S9759 })
);
AOI21_X1 #() 
AOI21_X1_469_ (
  .A({ S9063 }),
  .B1({ S9759 }),
  .B2({ S9758 }),
  .ZN({ S9760 })
);
NAND3_X1 #() 
NAND3_X1_889_ (
  .A1({ S9089 }),
  .A2({ S9087 }),
  .A3({ S25957[539] }),
  .ZN({ S9761 })
);
NAND3_X1 #() 
NAND3_X1_890_ (
  .A1({ S9761 }),
  .A2({ S25957[541] }),
  .A3({ S9439 }),
  .ZN({ S9762 })
);
OAI21_X1 #() 
OAI21_X1_430_ (
  .A({ S15 }),
  .B1({ S9157 }),
  .B2({ S9233 }),
  .ZN({ S9763 })
);
INV_X1 #() 
INV_X1_261_ (
  .A({ S9731 }),
  .ZN({ S9764 })
);
NAND3_X1 #() 
NAND3_X1_891_ (
  .A1({ S9763 }),
  .A2({ S9099 }),
  .A3({ S9764 }),
  .ZN({ S9765 })
);
NAND2_X1 #() 
NAND2_X1_769_ (
  .A1({ S9765 }),
  .A2({ S9762 }),
  .ZN({ S9766 })
);
AOI21_X1 #() 
AOI21_X1_470_ (
  .A({ S9760 }),
  .B1({ S9766 }),
  .B2({ S9063 }),
  .ZN({ S9767 })
);
NAND3_X1 #() 
NAND3_X1_892_ (
  .A1({ S9752 }),
  .A2({ S9747 }),
  .A3({ S7106 }),
  .ZN({ S9769 })
);
OAI211_X1 #() 
OAI211_X1_263_ (
  .A({ S7026 }),
  .B({ S9769 }),
  .C1({ S9767 }),
  .C2({ S7106 }),
  .ZN({ S9770 })
);
AOI22_X1 #() 
AOI22_X1_83_ (
  .A1({ S9668 }),
  .A2({ S9720 }),
  .B1({ S9722 }),
  .B2({ S9063 }),
  .ZN({ S9771 })
);
OAI21_X1 #() 
OAI21_X1_431_ (
  .A({ S9750 }),
  .B1({ S25957[539] }),
  .B2({ S9077 }),
  .ZN({ S9772 })
);
OAI211_X1 #() 
OAI211_X1_264_ (
  .A({ S9772 }),
  .B({ S9099 }),
  .C1({ S25957[540] }),
  .C2({ S9196 }),
  .ZN({ S9773 })
);
OAI211_X1 #() 
OAI211_X1_265_ (
  .A({ S9773 }),
  .B({ S7106 }),
  .C1({ S9771 }),
  .C2({ S9099 }),
  .ZN({ S9774 })
);
AOI22_X1 #() 
AOI22_X1_84_ (
  .A1({ S9152 }),
  .A2({ S9117 }),
  .B1({ S9122 }),
  .B2({ S9071 }),
  .ZN({ S9775 })
);
OAI21_X1 #() 
OAI21_X1_432_ (
  .A({ S9711 }),
  .B1({ S9063 }),
  .B2({ S9775 }),
  .ZN({ S9776 })
);
NAND2_X1 #() 
NAND2_X1_770_ (
  .A1({ S9714 }),
  .A2({ S9708 }),
  .ZN({ S9777 })
);
NAND3_X1 #() 
NAND3_X1_893_ (
  .A1({ S9776 }),
  .A2({ S9777 }),
  .A3({ S25957[542] }),
  .ZN({ S9778 })
);
NAND3_X1 #() 
NAND3_X1_894_ (
  .A1({ S9778 }),
  .A2({ S9774 }),
  .A3({ S25957[543] }),
  .ZN({ S9779 })
);
AOI21_X1 #() 
AOI21_X1_471_ (
  .A({ S25957[706] }),
  .B1({ S9770 }),
  .B2({ S9779 }),
  .ZN({ S9780 })
);
OAI21_X1 #() 
OAI21_X1_433_ (
  .A({ S25957[642] }),
  .B1({ S9780 }),
  .B2({ S9756 }),
  .ZN({ S9781 })
);
AOI21_X1 #() 
AOI21_X1_472_ (
  .A({ S7106 }),
  .B1({ S9740 }),
  .B2({ S9736 }),
  .ZN({ S9782 })
);
AOI22_X1 #() 
AOI22_X1_85_ (
  .A1({ S7106 }),
  .A2({ S9753 }),
  .B1({ S9782 }),
  .B2({ S9733 }),
  .ZN({ S9783 })
);
OAI211_X1 #() 
OAI211_X1_266_ (
  .A({ S25957[706] }),
  .B({ S9779 }),
  .C1({ S9783 }),
  .C2({ S25957[543] }),
  .ZN({ S9784 })
);
NAND3_X1 #() 
NAND3_X1_895_ (
  .A1({ S9755 }),
  .A2({ S9727 }),
  .A3({ S6831 }),
  .ZN({ S9785 })
);
NAND3_X1 #() 
NAND3_X1_896_ (
  .A1({ S9784 }),
  .A2({ S9785 }),
  .A3({ S5471 }),
  .ZN({ S9786 })
);
NAND2_X1 #() 
NAND2_X1_771_ (
  .A1({ S9781 }),
  .A2({ S9786 }),
  .ZN({ S25957[386] })
);
OAI21_X1 #() 
OAI21_X1_434_ (
  .A({ S25957[656] }),
  .B1({ S5283 }),
  .B2({ S5284 }),
  .ZN({ S9787 })
);
NAND3_X1 #() 
NAND3_X1_897_ (
  .A1({ S5277 }),
  .A2({ S5280 }),
  .A3({ S5282 }),
  .ZN({ S9788 })
);
NAND4_X1 #() 
NAND4_X1_89_ (
  .A1({ S8136 }),
  .A2({ S9787 }),
  .A3({ S8132 }),
  .A4({ S9788 }),
  .ZN({ S9789 })
);
INV_X1 #() 
INV_X1_262_ (
  .A({ S9789 }),
  .ZN({ S25 })
);
NAND4_X1 #() 
NAND4_X1_90_ (
  .A1({ S5362 }),
  .A2({ S5354 }),
  .A3({ S5285 }),
  .A4({ S5281 }),
  .ZN({ S26 })
);
XOR2_X1 #() 
XOR2_X1_15_ (
  .A({ S25957[863] }),
  .B({ S25957[959] }),
  .Z({ S25957[831] })
);
XNOR2_X1 #() 
XNOR2_X1_25_ (
  .A({ S4281 }),
  .B({ S25957[831] }),
  .ZN({ S25957[703] })
);
XNOR2_X1 #() 
XNOR2_X1_26_ (
  .A({ S7025 }),
  .B({ S25957[863] }),
  .ZN({ S25957[607] })
);
XOR2_X1 #() 
XOR2_X1_16_ (
  .A({ S25957[607] }),
  .B({ S25957[703] }),
  .Z({ S25957[575] })
);
NAND2_X1 #() 
NAND2_X1_772_ (
  .A1({ S5063 }),
  .A2({ S5066 }),
  .ZN({ S9790 })
);
NAND3_X1 #() 
NAND3_X1_898_ (
  .A1({ S26 }),
  .A2({ S25957[530] }),
  .A3({ S9789 }),
  .ZN({ S9791 })
);
AOI22_X1 #() 
AOI22_X1_86_ (
  .A1({ S5285 }),
  .A2({ S5281 }),
  .B1({ S8277 }),
  .B2({ S8280 }),
  .ZN({ S9793 })
);
AOI21_X1 #() 
AOI21_X1_473_ (
  .A({ S25957[531] }),
  .B1({ S9793 }),
  .B2({ S25957[529] }),
  .ZN({ S9794 })
);
NAND2_X1 #() 
NAND2_X1_773_ (
  .A1({ S9794 }),
  .A2({ S9791 }),
  .ZN({ S9795 })
);
INV_X1 #() 
INV_X1_263_ (
  .A({ S9795 }),
  .ZN({ S9796 })
);
NAND4_X1 #() 
NAND4_X1_91_ (
  .A1({ S5285 }),
  .A2({ S8277 }),
  .A3({ S8280 }),
  .A4({ S5281 }),
  .ZN({ S9797 })
);
NOR2_X1 #() 
NOR2_X1_177_ (
  .A1({ S9797 }),
  .A2({ S8137 }),
  .ZN({ S9798 })
);
OAI21_X1 #() 
OAI21_X1_435_ (
  .A({ S25957[532] }),
  .B1({ S9798 }),
  .B2({ S6 }),
  .ZN({ S9799 })
);
NAND4_X1 #() 
NAND4_X1_92_ (
  .A1({ S8136 }),
  .A2({ S5285 }),
  .A3({ S8132 }),
  .A4({ S5281 }),
  .ZN({ S9800 })
);
NAND4_X1 #() 
NAND4_X1_93_ (
  .A1({ S5362 }),
  .A2({ S5354 }),
  .A3({ S9788 }),
  .A4({ S9787 }),
  .ZN({ S9801 })
);
NAND4_X1 #() 
NAND4_X1_94_ (
  .A1({ S9801 }),
  .A2({ S9800 }),
  .A3({ S25957[530] }),
  .A4({ S6 }),
  .ZN({ S9802 })
);
NAND2_X1 #() 
NAND2_X1_774_ (
  .A1({ S9789 }),
  .A2({ S25957[530] }),
  .ZN({ S9804 })
);
OAI211_X1 #() 
OAI211_X1_267_ (
  .A({ S9802 }),
  .B({ S5128 }),
  .C1({ S6 }),
  .C2({ S9804 }),
  .ZN({ S9805 })
);
OAI211_X1 #() 
OAI211_X1_268_ (
  .A({ S9790 }),
  .B({ S9805 }),
  .C1({ S9796 }),
  .C2({ S9799 }),
  .ZN({ S9806 })
);
NAND4_X1 #() 
NAND4_X1_95_ (
  .A1({ S5461 }),
  .A2({ S8136 }),
  .A3({ S8132 }),
  .A4({ S5455 }),
  .ZN({ S9807 })
);
NAND3_X1 #() 
NAND3_X1_899_ (
  .A1({ S9801 }),
  .A2({ S25957[531] }),
  .A3({ S9807 }),
  .ZN({ S9808 })
);
INV_X1 #() 
INV_X1_264_ (
  .A({ S9808 }),
  .ZN({ S9809 })
);
NAND2_X1 #() 
NAND2_X1_775_ (
  .A1({ S9789 }),
  .A2({ S8281 }),
  .ZN({ S9810 })
);
AOI21_X1 #() 
AOI21_X1_474_ (
  .A({ S25957[531] }),
  .B1({ S25957[529] }),
  .B2({ S25957[530] }),
  .ZN({ S9811 })
);
AOI21_X1 #() 
AOI21_X1_475_ (
  .A({ S9809 }),
  .B1({ S9810 }),
  .B2({ S9811 }),
  .ZN({ S9812 })
);
NAND4_X1 #() 
NAND4_X1_96_ (
  .A1({ S5362 }),
  .A2({ S5461 }),
  .A3({ S5354 }),
  .A4({ S5455 }),
  .ZN({ S9813 })
);
AOI21_X1 #() 
AOI21_X1_476_ (
  .A({ S6 }),
  .B1({ S25957[530] }),
  .B2({ S25957[528] }),
  .ZN({ S9815 })
);
NAND2_X1 #() 
NAND2_X1_776_ (
  .A1({ S9815 }),
  .A2({ S9813 }),
  .ZN({ S9816 })
);
NAND2_X1 #() 
NAND2_X1_777_ (
  .A1({ S6 }),
  .A2({ S25957[528] }),
  .ZN({ S9817 })
);
NAND3_X1 #() 
NAND3_X1_900_ (
  .A1({ S9816 }),
  .A2({ S25957[532] }),
  .A3({ S9817 }),
  .ZN({ S9818 })
);
OAI21_X1 #() 
OAI21_X1_436_ (
  .A({ S9818 }),
  .B1({ S9812 }),
  .B2({ S25957[532] }),
  .ZN({ S9819 })
);
OAI21_X1 #() 
OAI21_X1_437_ (
  .A({ S9806 }),
  .B1({ S9819 }),
  .B2({ S9790 }),
  .ZN({ S9820 })
);
NAND2_X1 #() 
NAND2_X1_778_ (
  .A1({ S9815 }),
  .A2({ S9807 }),
  .ZN({ S9821 })
);
NAND4_X1 #() 
NAND4_X1_97_ (
  .A1({ S5362 }),
  .A2({ S5354 }),
  .A3({ S8277 }),
  .A4({ S8280 }),
  .ZN({ S9822 })
);
NAND4_X1 #() 
NAND4_X1_98_ (
  .A1({ S5461 }),
  .A2({ S5285 }),
  .A3({ S5455 }),
  .A4({ S5281 }),
  .ZN({ S9823 })
);
NAND4_X1 #() 
NAND4_X1_99_ (
  .A1({ S9822 }),
  .A2({ S9807 }),
  .A3({ S9823 }),
  .A4({ S9797 }),
  .ZN({ S9824 })
);
AOI21_X1 #() 
AOI21_X1_477_ (
  .A({ S25957[532] }),
  .B1({ S9824 }),
  .B2({ S6 }),
  .ZN({ S9826 })
);
NAND3_X1 #() 
NAND3_X1_901_ (
  .A1({ S9801 }),
  .A2({ S8281 }),
  .A3({ S9800 }),
  .ZN({ S9827 })
);
AOI21_X1 #() 
AOI21_X1_478_ (
  .A({ S6 }),
  .B1({ S9827 }),
  .B2({ S9804 }),
  .ZN({ S9828 })
);
NAND3_X1 #() 
NAND3_X1_902_ (
  .A1({ S9801 }),
  .A2({ S25957[530] }),
  .A3({ S9800 }),
  .ZN({ S9829 })
);
AOI21_X1 #() 
AOI21_X1_479_ (
  .A({ S25957[531] }),
  .B1({ S9829 }),
  .B2({ S9823 }),
  .ZN({ S9830 })
);
NOR3_X1 #() 
NOR3_X1_25_ (
  .A1({ S9830 }),
  .A2({ S9828 }),
  .A3({ S5128 }),
  .ZN({ S9831 })
);
AOI21_X1 #() 
AOI21_X1_480_ (
  .A({ S9831 }),
  .B1({ S9826 }),
  .B2({ S9821 }),
  .ZN({ S9832 })
);
AOI21_X1 #() 
AOI21_X1_481_ (
  .A({ S25957[528] }),
  .B1({ S25957[530] }),
  .B2({ S8137 }),
  .ZN({ S9833 })
);
OAI21_X1 #() 
OAI21_X1_438_ (
  .A({ S25957[532] }),
  .B1({ S9833 }),
  .B2({ S25957[531] }),
  .ZN({ S9834 })
);
NAND4_X1 #() 
NAND4_X1_100_ (
  .A1({ S25957[528] }),
  .A2({ S8281 }),
  .A3({ S8132 }),
  .A4({ S8136 }),
  .ZN({ S9835 })
);
NAND2_X1 #() 
NAND2_X1_779_ (
  .A1({ S9787 }),
  .A2({ S9788 }),
  .ZN({ S9837 })
);
NAND3_X1 #() 
NAND3_X1_903_ (
  .A1({ S25957[530] }),
  .A2({ S8137 }),
  .A3({ S9837 }),
  .ZN({ S9838 })
);
NAND2_X1 #() 
NAND2_X1_780_ (
  .A1({ S9838 }),
  .A2({ S9835 }),
  .ZN({ S9839 })
);
NOR2_X1 #() 
NOR2_X1_178_ (
  .A1({ S9839 }),
  .A2({ S6 }),
  .ZN({ S9840 })
);
NAND4_X1 #() 
NAND4_X1_101_ (
  .A1({ S8132 }),
  .A2({ S8136 }),
  .A3({ S8277 }),
  .A4({ S8280 }),
  .ZN({ S9841 })
);
NAND3_X1 #() 
NAND3_X1_904_ (
  .A1({ S8137 }),
  .A2({ S25957[528] }),
  .A3({ S8281 }),
  .ZN({ S9842 })
);
NAND2_X1 #() 
NAND2_X1_781_ (
  .A1({ S9842 }),
  .A2({ S9841 }),
  .ZN({ S9843 })
);
NAND2_X1 #() 
NAND2_X1_782_ (
  .A1({ S9843 }),
  .A2({ S25957[531] }),
  .ZN({ S9844 })
);
NAND2_X1 #() 
NAND2_X1_783_ (
  .A1({ S9804 }),
  .A2({ S6 }),
  .ZN({ S9845 })
);
NAND3_X1 #() 
NAND3_X1_905_ (
  .A1({ S9844 }),
  .A2({ S5128 }),
  .A3({ S9845 }),
  .ZN({ S9846 })
);
OAI211_X1 #() 
OAI211_X1_269_ (
  .A({ S9846 }),
  .B({ S25957[533] }),
  .C1({ S9834 }),
  .C2({ S9840 }),
  .ZN({ S9848 })
);
OAI21_X1 #() 
OAI21_X1_439_ (
  .A({ S9848 }),
  .B1({ S9832 }),
  .B2({ S25957[533] }),
  .ZN({ S9849 })
);
MUX2_X1 #() 
MUX2_X1_2_ (
  .A({ S9820 }),
  .B({ S9849 }),
  .S({ S25957[534] }),
  .Z({ S9850 })
);
NOR2_X1 #() 
NOR2_X1_179_ (
  .A1({ S9850 }),
  .A2({ S25957[535] }),
  .ZN({ S9851 })
);
AOI22_X1 #() 
AOI22_X1_87_ (
  .A1({ S8136 }),
  .A2({ S8132 }),
  .B1({ S8277 }),
  .B2({ S8280 }),
  .ZN({ S9852 })
);
NAND2_X1 #() 
NAND2_X1_784_ (
  .A1({ S9797 }),
  .A2({ S6 }),
  .ZN({ S9853 })
);
NAND4_X1 #() 
NAND4_X1_102_ (
  .A1({ S5461 }),
  .A2({ S9787 }),
  .A3({ S5455 }),
  .A4({ S9788 }),
  .ZN({ S9854 })
);
NAND2_X1 #() 
NAND2_X1_785_ (
  .A1({ S9854 }),
  .A2({ S8137 }),
  .ZN({ S9855 })
);
AOI21_X1 #() 
AOI21_X1_482_ (
  .A({ S9853 }),
  .B1({ S9855 }),
  .B2({ S9835 }),
  .ZN({ S9856 })
);
AOI21_X1 #() 
AOI21_X1_483_ (
  .A({ S9856 }),
  .B1({ S9852 }),
  .B2({ S25957[531] }),
  .ZN({ S9857 })
);
AOI21_X1 #() 
AOI21_X1_484_ (
  .A({ S6 }),
  .B1({ S9791 }),
  .B2({ S9827 }),
  .ZN({ S9859 })
);
INV_X1 #() 
INV_X1_265_ (
  .A({ S9841 }),
  .ZN({ S9860 })
);
AOI22_X1 #() 
AOI22_X1_88_ (
  .A1({ S25957[528] }),
  .A2({ S8281 }),
  .B1({ S5223 }),
  .B2({ S5220 }),
  .ZN({ S9861 })
);
INV_X1 #() 
INV_X1_266_ (
  .A({ S9861 }),
  .ZN({ S9862 })
);
OAI21_X1 #() 
OAI21_X1_440_ (
  .A({ S25957[532] }),
  .B1({ S9862 }),
  .B2({ S9860 }),
  .ZN({ S9863 })
);
OAI22_X1 #() 
OAI22_X1_21_ (
  .A1({ S9857 }),
  .A2({ S25957[532] }),
  .B1({ S9859 }),
  .B2({ S9863 }),
  .ZN({ S9864 })
);
NAND4_X1 #() 
NAND4_X1_103_ (
  .A1({ S9787 }),
  .A2({ S8277 }),
  .A3({ S8280 }),
  .A4({ S9788 }),
  .ZN({ S9865 })
);
INV_X1 #() 
INV_X1_267_ (
  .A({ S9865 }),
  .ZN({ S9866 })
);
NAND4_X1 #() 
NAND4_X1_104_ (
  .A1({ S8132 }),
  .A2({ S8136 }),
  .A3({ S5224 }),
  .A4({ S5225 }),
  .ZN({ S9867 })
);
OAI21_X1 #() 
OAI21_X1_441_ (
  .A({ S25957[531] }),
  .B1({ S9866 }),
  .B2({ S8137 }),
  .ZN({ S9868 })
);
OAI211_X1 #() 
OAI211_X1_270_ (
  .A({ S9868 }),
  .B({ S25957[532] }),
  .C1({ S9866 }),
  .C2({ S9867 }),
  .ZN({ S9870 })
);
AOI21_X1 #() 
AOI21_X1_485_ (
  .A({ S25957[531] }),
  .B1({ S9837 }),
  .B2({ S8281 }),
  .ZN({ S9871 })
);
NAND3_X1 #() 
NAND3_X1_906_ (
  .A1({ S9789 }),
  .A2({ S9867 }),
  .A3({ S5128 }),
  .ZN({ S9872 })
);
OAI211_X1 #() 
OAI211_X1_271_ (
  .A({ S9870 }),
  .B({ S25957[533] }),
  .C1({ S9871 }),
  .C2({ S9872 }),
  .ZN({ S9873 })
);
OAI211_X1 #() 
OAI211_X1_272_ (
  .A({ S7708 }),
  .B({ S9873 }),
  .C1({ S9864 }),
  .C2({ S25957[533] }),
  .ZN({ S9874 })
);
AND2_X1 #() 
AND2_X1_50_ (
  .A1({ S8137 }),
  .A2({ S25957[528] }),
  .ZN({ S9875 })
);
OAI21_X1 #() 
OAI21_X1_442_ (
  .A({ S25957[531] }),
  .B1({ S9798 }),
  .B2({ S9875 }),
  .ZN({ S9876 })
);
AOI21_X1 #() 
AOI21_X1_486_ (
  .A({ S25957[532] }),
  .B1({ S9839 }),
  .B2({ S6 }),
  .ZN({ S9877 })
);
AOI22_X1 #() 
AOI22_X1_89_ (
  .A1({ S8137 }),
  .A2({ S25957[528] }),
  .B1({ S8277 }),
  .B2({ S8280 }),
  .ZN({ S9878 })
);
OAI21_X1 #() 
OAI21_X1_443_ (
  .A({ S25957[531] }),
  .B1({ S9878 }),
  .B2({ S9866 }),
  .ZN({ S9879 })
);
NOR2_X1 #() 
NOR2_X1_180_ (
  .A1({ S8137 }),
  .A2({ S25957[531] }),
  .ZN({ S9881 })
);
AOI21_X1 #() 
AOI21_X1_487_ (
  .A({ S5128 }),
  .B1({ S9881 }),
  .B2({ S9823 }),
  .ZN({ S9882 })
);
AOI22_X1 #() 
AOI22_X1_90_ (
  .A1({ S9877 }),
  .A2({ S9876 }),
  .B1({ S9879 }),
  .B2({ S9882 }),
  .ZN({ S9883 })
);
INV_X1 #() 
INV_X1_268_ (
  .A({ S9822 }),
  .ZN({ S9884 })
);
NAND2_X1 #() 
NAND2_X1_786_ (
  .A1({ S9789 }),
  .A2({ S25957[531] }),
  .ZN({ S9885 })
);
NAND2_X1 #() 
NAND2_X1_787_ (
  .A1({ S9800 }),
  .A2({ S6 }),
  .ZN({ S9886 })
);
OAI211_X1 #() 
OAI211_X1_273_ (
  .A({ S25957[532] }),
  .B({ S9886 }),
  .C1({ S9884 }),
  .C2({ S9885 }),
  .ZN({ S9887 })
);
NAND2_X1 #() 
NAND2_X1_788_ (
  .A1({ S26 }),
  .A2({ S25957[530] }),
  .ZN({ S9888 })
);
AOI22_X1 #() 
AOI22_X1_91_ (
  .A1({ S9788 }),
  .A2({ S9787 }),
  .B1({ S8277 }),
  .B2({ S8280 }),
  .ZN({ S9889 })
);
NAND2_X1 #() 
NAND2_X1_789_ (
  .A1({ S9889 }),
  .A2({ S8137 }),
  .ZN({ S9890 })
);
OAI211_X1 #() 
OAI211_X1_274_ (
  .A({ S9888 }),
  .B({ S9890 }),
  .C1({ S9801 }),
  .C2({ S6 }),
  .ZN({ S9892 })
);
AOI21_X1 #() 
AOI21_X1_488_ (
  .A({ S25957[533] }),
  .B1({ S9892 }),
  .B2({ S5128 }),
  .ZN({ S9893 })
);
AOI22_X1 #() 
AOI22_X1_92_ (
  .A1({ S9883 }),
  .A2({ S25957[533] }),
  .B1({ S9887 }),
  .B2({ S9893 }),
  .ZN({ S9894 })
);
NAND2_X1 #() 
NAND2_X1_790_ (
  .A1({ S9894 }),
  .A2({ S25957[534] }),
  .ZN({ S9895 })
);
NAND3_X1 #() 
NAND3_X1_907_ (
  .A1({ S9895 }),
  .A2({ S9874 }),
  .A3({ S25957[535] }),
  .ZN({ S9896 })
);
INV_X1 #() 
INV_X1_269_ (
  .A({ S9896 }),
  .ZN({ S9897 })
);
NOR3_X1 #() 
NOR3_X1_26_ (
  .A1({ S9851 }),
  .A2({ S9897 }),
  .A3({ S4281 }),
  .ZN({ S9898 })
);
NOR2_X1 #() 
NOR2_X1_181_ (
  .A1({ S9851 }),
  .A2({ S9897 }),
  .ZN({ S9899 })
);
NOR2_X1 #() 
NOR2_X1_182_ (
  .A1({ S9899 }),
  .A2({ S25957[735] }),
  .ZN({ S9900 })
);
NOR2_X1 #() 
NOR2_X1_183_ (
  .A1({ S9900 }),
  .A2({ S9898 }),
  .ZN({ S25957[479] })
);
NAND2_X1 #() 
NAND2_X1_791_ (
  .A1({ S25957[479] }),
  .A2({ S25957[575] }),
  .ZN({ S9902 })
);
INV_X1 #() 
INV_X1_270_ (
  .A({ S25957[575] }),
  .ZN({ S9903 })
);
INV_X1 #() 
INV_X1_271_ (
  .A({ S25957[479] }),
  .ZN({ S9904 })
);
NAND2_X1 #() 
NAND2_X1_792_ (
  .A1({ S9904 }),
  .A2({ S9903 }),
  .ZN({ S9905 })
);
NAND3_X1 #() 
NAND3_X1_908_ (
  .A1({ S9905 }),
  .A2({ S25957[543] }),
  .A3({ S9902 }),
  .ZN({ S9906 })
);
NAND2_X1 #() 
NAND2_X1_793_ (
  .A1({ S9904 }),
  .A2({ S25957[575] }),
  .ZN({ S9907 })
);
NAND2_X1 #() 
NAND2_X1_794_ (
  .A1({ S25957[479] }),
  .A2({ S9903 }),
  .ZN({ S9908 })
);
NAND3_X1 #() 
NAND3_X1_909_ (
  .A1({ S9907 }),
  .A2({ S7026 }),
  .A3({ S9908 }),
  .ZN({ S9909 })
);
NAND2_X1 #() 
NAND2_X1_795_ (
  .A1({ S9906 }),
  .A2({ S9909 }),
  .ZN({ S9910 })
);
INV_X1 #() 
INV_X1_272_ (
  .A({ S9910 }),
  .ZN({ S25957[415] })
);
NAND2_X1 #() 
NAND2_X1_796_ (
  .A1({ S4352 }),
  .A2({ S4349 }),
  .ZN({ S25957[702] })
);
XNOR2_X1 #() 
XNOR2_X1_27_ (
  .A({ S7102 }),
  .B({ S1804 }),
  .ZN({ S25957[606] })
);
XOR2_X1 #() 
XOR2_X1_17_ (
  .A({ S25957[606] }),
  .B({ S25957[702] }),
  .Z({ S25957[574] })
);
NAND2_X1 #() 
NAND2_X1_797_ (
  .A1({ S4344 }),
  .A2({ S4347 }),
  .ZN({ S25957[766] })
);
XOR2_X1 #() 
XOR2_X1_18_ (
  .A({ S7102 }),
  .B({ S25957[766] }),
  .Z({ S25957[638] })
);
AOI22_X1 #() 
AOI22_X1_93_ (
  .A1({ S25957[528] }),
  .A2({ S8281 }),
  .B1({ S5362 }),
  .B2({ S5354 }),
  .ZN({ S9912 })
);
OAI21_X1 #() 
OAI21_X1_444_ (
  .A({ S5128 }),
  .B1({ S9865 }),
  .B2({ S6 }),
  .ZN({ S9913 })
);
AOI21_X1 #() 
AOI21_X1_489_ (
  .A({ S25957[531] }),
  .B1({ S9789 }),
  .B2({ S25957[530] }),
  .ZN({ S9914 })
);
NAND2_X1 #() 
NAND2_X1_798_ (
  .A1({ S26 }),
  .A2({ S9854 }),
  .ZN({ S9915 })
);
NOR2_X1 #() 
NOR2_X1_184_ (
  .A1({ S9915 }),
  .A2({ S6 }),
  .ZN({ S9916 })
);
AOI21_X1 #() 
AOI21_X1_490_ (
  .A({ S9916 }),
  .B1({ S9914 }),
  .B2({ S9854 }),
  .ZN({ S9918 })
);
OAI221_X1 #() 
OAI221_X1_16_ (
  .A({ S25957[533] }),
  .B1({ S9912 }),
  .B2({ S9913 }),
  .C1({ S9918 }),
  .C2({ S5128 }),
  .ZN({ S9919 })
);
NAND2_X1 #() 
NAND2_X1_799_ (
  .A1({ S9791 }),
  .A2({ S6 }),
  .ZN({ S9920 })
);
NAND3_X1 #() 
NAND3_X1_910_ (
  .A1({ S9854 }),
  .A2({ S9841 }),
  .A3({ S9797 }),
  .ZN({ S9921 })
);
AOI21_X1 #() 
AOI21_X1_491_ (
  .A({ S25957[532] }),
  .B1({ S9921 }),
  .B2({ S25957[531] }),
  .ZN({ S9922 })
);
NAND2_X1 #() 
NAND2_X1_800_ (
  .A1({ S9807 }),
  .A2({ S25957[531] }),
  .ZN({ S9923 })
);
NAND3_X1 #() 
NAND3_X1_911_ (
  .A1({ S9800 }),
  .A2({ S6 }),
  .A3({ S9797 }),
  .ZN({ S9924 })
);
AOI21_X1 #() 
AOI21_X1_492_ (
  .A({ S5128 }),
  .B1({ S9924 }),
  .B2({ S9923 }),
  .ZN({ S9925 })
);
AOI21_X1 #() 
AOI21_X1_493_ (
  .A({ S9925 }),
  .B1({ S9922 }),
  .B2({ S9920 }),
  .ZN({ S9926 })
);
NAND2_X1 #() 
NAND2_X1_801_ (
  .A1({ S9926 }),
  .A2({ S9790 }),
  .ZN({ S9927 })
);
AOI21_X1 #() 
AOI21_X1_494_ (
  .A({ S7708 }),
  .B1({ S9919 }),
  .B2({ S9927 }),
  .ZN({ S9929 })
);
AOI21_X1 #() 
AOI21_X1_495_ (
  .A({ S25957[531] }),
  .B1({ S9852 }),
  .B2({ S25957[528] }),
  .ZN({ S9930 })
);
NOR2_X1 #() 
NOR2_X1_185_ (
  .A1({ S9930 }),
  .A2({ S5128 }),
  .ZN({ S9931 })
);
NAND2_X1 #() 
NAND2_X1_802_ (
  .A1({ S9813 }),
  .A2({ S9854 }),
  .ZN({ S9932 })
);
OAI21_X1 #() 
OAI21_X1_445_ (
  .A({ S25957[531] }),
  .B1({ S9932 }),
  .B2({ S9798 }),
  .ZN({ S9933 })
);
NOR2_X1 #() 
NOR2_X1_186_ (
  .A1({ S9933 }),
  .A2({ S25957[532] }),
  .ZN({ S9934 })
);
AOI211_X1 #() 
AOI211_X1_10_ (
  .A({ S25957[533] }),
  .B({ S9934 }),
  .C1({ S9844 }),
  .C2({ S9931 }),
  .ZN({ S9935 })
);
NAND3_X1 #() 
NAND3_X1_912_ (
  .A1({ S9838 }),
  .A2({ S25957[531] }),
  .A3({ S9789 }),
  .ZN({ S9936 })
);
NAND3_X1 #() 
NAND3_X1_913_ (
  .A1({ S9936 }),
  .A2({ S25957[532] }),
  .A3({ S9862 }),
  .ZN({ S9937 })
);
NAND2_X1 #() 
NAND2_X1_803_ (
  .A1({ S9811 }),
  .A2({ S9842 }),
  .ZN({ S9938 })
);
OAI21_X1 #() 
OAI21_X1_446_ (
  .A({ S9938 }),
  .B1({ S9884 }),
  .B2({ S9923 }),
  .ZN({ S9940 })
);
OR2_X1 #() 
OR2_X1_10_ (
  .A1({ S9940 }),
  .A2({ S25957[532] }),
  .ZN({ S9941 })
);
AOI21_X1 #() 
AOI21_X1_496_ (
  .A({ S9790 }),
  .B1({ S9941 }),
  .B2({ S9937 }),
  .ZN({ S9942 })
);
NOR3_X1 #() 
NOR3_X1_27_ (
  .A1({ S9935 }),
  .A2({ S9942 }),
  .A3({ S25957[534] }),
  .ZN({ S9943 })
);
OAI21_X1 #() 
OAI21_X1_447_ (
  .A({ S4924 }),
  .B1({ S9943 }),
  .B2({ S9929 }),
  .ZN({ S9944 })
);
AOI21_X1 #() 
AOI21_X1_497_ (
  .A({ S6 }),
  .B1({ S25957[530] }),
  .B2({ S9837 }),
  .ZN({ S9945 })
);
AOI22_X1 #() 
AOI22_X1_94_ (
  .A1({ S25957[528] }),
  .A2({ S8281 }),
  .B1({ S8132 }),
  .B2({ S8136 }),
  .ZN({ S9946 })
);
NAND2_X1 #() 
NAND2_X1_804_ (
  .A1({ S9945 }),
  .A2({ S9946 }),
  .ZN({ S9947 })
);
NAND2_X1 #() 
NAND2_X1_805_ (
  .A1({ S9841 }),
  .A2({ S9865 }),
  .ZN({ S9948 })
);
NAND2_X1 #() 
NAND2_X1_806_ (
  .A1({ S9948 }),
  .A2({ S6 }),
  .ZN({ S9949 })
);
AOI21_X1 #() 
AOI21_X1_498_ (
  .A({ S5128 }),
  .B1({ S9947 }),
  .B2({ S9949 }),
  .ZN({ S9951 })
);
OAI21_X1 #() 
OAI21_X1_448_ (
  .A({ S9867 }),
  .B1({ S9884 }),
  .B2({ S9885 }),
  .ZN({ S9952 })
);
OAI21_X1 #() 
OAI21_X1_449_ (
  .A({ S25957[533] }),
  .B1({ S9952 }),
  .B2({ S25957[532] }),
  .ZN({ S9953 })
);
AOI21_X1 #() 
AOI21_X1_499_ (
  .A({ S25957[530] }),
  .B1({ S26 }),
  .B2({ S9789 }),
  .ZN({ S9954 })
);
AOI21_X1 #() 
AOI21_X1_500_ (
  .A({ S5128 }),
  .B1({ S9921 }),
  .B2({ S25957[531] }),
  .ZN({ S9955 })
);
OAI21_X1 #() 
OAI21_X1_450_ (
  .A({ S9955 }),
  .B1({ S9853 }),
  .B2({ S9954 }),
  .ZN({ S9956 })
);
AOI22_X1 #() 
AOI22_X1_95_ (
  .A1({ S8136 }),
  .A2({ S8132 }),
  .B1({ S9787 }),
  .B2({ S9788 }),
  .ZN({ S9957 })
);
NAND3_X1 #() 
NAND3_X1_914_ (
  .A1({ S9813 }),
  .A2({ S25957[531] }),
  .A3({ S9823 }),
  .ZN({ S9958 })
);
OAI21_X1 #() 
OAI21_X1_451_ (
  .A({ S9826 }),
  .B1({ S9957 }),
  .B2({ S9958 }),
  .ZN({ S9959 })
);
NAND3_X1 #() 
NAND3_X1_915_ (
  .A1({ S9959 }),
  .A2({ S9790 }),
  .A3({ S9956 }),
  .ZN({ S9960 })
);
OAI21_X1 #() 
OAI21_X1_452_ (
  .A({ S9960 }),
  .B1({ S9951 }),
  .B2({ S9953 }),
  .ZN({ S9962 })
);
NAND2_X1 #() 
NAND2_X1_807_ (
  .A1({ S9962 }),
  .A2({ S25957[534] }),
  .ZN({ S9963 })
);
NOR2_X1 #() 
NOR2_X1_187_ (
  .A1({ S9954 }),
  .A2({ S9853 }),
  .ZN({ S9964 })
);
NAND3_X1 #() 
NAND3_X1_916_ (
  .A1({ S25957[529] }),
  .A2({ S25957[530] }),
  .A3({ S9837 }),
  .ZN({ S9965 })
);
AOI21_X1 #() 
AOI21_X1_501_ (
  .A({ S6 }),
  .B1({ S9965 }),
  .B2({ S9854 }),
  .ZN({ S9966 })
);
OAI21_X1 #() 
OAI21_X1_453_ (
  .A({ S5128 }),
  .B1({ S9964 }),
  .B2({ S9966 }),
  .ZN({ S9967 })
);
NAND2_X1 #() 
NAND2_X1_808_ (
  .A1({ S9801 }),
  .A2({ S8281 }),
  .ZN({ S9968 })
);
OAI211_X1 #() 
OAI211_X1_275_ (
  .A({ S9868 }),
  .B({ S25957[532] }),
  .C1({ S25957[531] }),
  .C2({ S9968 }),
  .ZN({ S9969 })
);
NAND3_X1 #() 
NAND3_X1_917_ (
  .A1({ S9967 }),
  .A2({ S9790 }),
  .A3({ S9969 }),
  .ZN({ S9970 })
);
NAND4_X1 #() 
NAND4_X1_105_ (
  .A1({ S5220 }),
  .A2({ S5223 }),
  .A3({ S8277 }),
  .A4({ S8280 }),
  .ZN({ S9971 })
);
INV_X1 #() 
INV_X1_273_ (
  .A({ S9971 }),
  .ZN({ S9973 })
);
NAND2_X1 #() 
NAND2_X1_809_ (
  .A1({ S9973 }),
  .A2({ S25957[529] }),
  .ZN({ S9974 })
);
NAND2_X1 #() 
NAND2_X1_810_ (
  .A1({ S9881 }),
  .A2({ S9889 }),
  .ZN({ S9975 })
);
NAND2_X1 #() 
NAND2_X1_811_ (
  .A1({ S9975 }),
  .A2({ S9974 }),
  .ZN({ S9976 })
);
NAND2_X1 #() 
NAND2_X1_812_ (
  .A1({ S9802 }),
  .A2({ S25957[532] }),
  .ZN({ S9977 })
);
NAND3_X1 #() 
NAND3_X1_918_ (
  .A1({ S25957[529] }),
  .A2({ S25957[530] }),
  .A3({ S25957[528] }),
  .ZN({ S9978 })
);
NAND3_X1 #() 
NAND3_X1_919_ (
  .A1({ S9978 }),
  .A2({ S6 }),
  .A3({ S26 }),
  .ZN({ S9979 })
);
NAND2_X1 #() 
NAND2_X1_813_ (
  .A1({ S9800 }),
  .A2({ S8281 }),
  .ZN({ S9980 })
);
NAND3_X1 #() 
NAND3_X1_920_ (
  .A1({ S9980 }),
  .A2({ S25957[531] }),
  .A3({ S9841 }),
  .ZN({ S9981 })
);
NAND3_X1 #() 
NAND3_X1_921_ (
  .A1({ S9979 }),
  .A2({ S9981 }),
  .A3({ S5128 }),
  .ZN({ S9982 })
);
OAI21_X1 #() 
OAI21_X1_454_ (
  .A({ S9982 }),
  .B1({ S9976 }),
  .B2({ S9977 }),
  .ZN({ S9984 })
);
NAND2_X1 #() 
NAND2_X1_814_ (
  .A1({ S9984 }),
  .A2({ S25957[533] }),
  .ZN({ S9985 })
);
NAND3_X1 #() 
NAND3_X1_922_ (
  .A1({ S9970 }),
  .A2({ S9985 }),
  .A3({ S7708 }),
  .ZN({ S9986 })
);
AOI21_X1 #() 
AOI21_X1_502_ (
  .A({ S4924 }),
  .B1({ S9963 }),
  .B2({ S9986 }),
  .ZN({ S9987 })
);
INV_X1 #() 
INV_X1_274_ (
  .A({ S9987 }),
  .ZN({ S9988 })
);
NAND3_X1 #() 
NAND3_X1_923_ (
  .A1({ S9988 }),
  .A2({ S9944 }),
  .A3({ S25957[638] }),
  .ZN({ S9989 })
);
INV_X1 #() 
INV_X1_275_ (
  .A({ S25957[638] }),
  .ZN({ S9990 })
);
INV_X1 #() 
INV_X1_276_ (
  .A({ S9944 }),
  .ZN({ S9991 })
);
OAI21_X1 #() 
OAI21_X1_455_ (
  .A({ S9990 }),
  .B1({ S9991 }),
  .B2({ S9987 }),
  .ZN({ S9992 })
);
NAND2_X1 #() 
NAND2_X1_815_ (
  .A1({ S9992 }),
  .A2({ S9989 }),
  .ZN({ S25957[510] })
);
NAND2_X1 #() 
NAND2_X1_816_ (
  .A1({ S25957[510] }),
  .A2({ S25957[606] }),
  .ZN({ S9994 })
);
INV_X1 #() 
INV_X1_277_ (
  .A({ S25957[606] }),
  .ZN({ S9995 })
);
NAND3_X1 #() 
NAND3_X1_924_ (
  .A1({ S9992 }),
  .A2({ S9989 }),
  .A3({ S9995 }),
  .ZN({ S9996 })
);
NAND3_X1 #() 
NAND3_X1_925_ (
  .A1({ S9994 }),
  .A2({ S9996 }),
  .A3({ S25957[574] }),
  .ZN({ S9997 })
);
INV_X1 #() 
INV_X1_278_ (
  .A({ S25957[574] }),
  .ZN({ S9998 })
);
NAND3_X1 #() 
NAND3_X1_926_ (
  .A1({ S9988 }),
  .A2({ S9944 }),
  .A3({ S9990 }),
  .ZN({ S9999 })
);
OAI21_X1 #() 
OAI21_X1_456_ (
  .A({ S25957[638] }),
  .B1({ S9991 }),
  .B2({ S9987 }),
  .ZN({ S10000 })
);
NAND3_X1 #() 
NAND3_X1_927_ (
  .A1({ S10000 }),
  .A2({ S9999 }),
  .A3({ S9995 }),
  .ZN({ S10001 })
);
NAND3_X1 #() 
NAND3_X1_928_ (
  .A1({ S9992 }),
  .A2({ S9989 }),
  .A3({ S25957[606] }),
  .ZN({ S10002 })
);
NAND3_X1 #() 
NAND3_X1_929_ (
  .A1({ S10001 }),
  .A2({ S10002 }),
  .A3({ S9998 }),
  .ZN({ S10003 })
);
NAND3_X1 #() 
NAND3_X1_930_ (
  .A1({ S9997 }),
  .A2({ S10003 }),
  .A3({ S25957[542] }),
  .ZN({ S10005 })
);
NAND3_X1 #() 
NAND3_X1_931_ (
  .A1({ S9994 }),
  .A2({ S9996 }),
  .A3({ S9998 }),
  .ZN({ S10006 })
);
NAND3_X1 #() 
NAND3_X1_932_ (
  .A1({ S10001 }),
  .A2({ S10002 }),
  .A3({ S25957[574] }),
  .ZN({ S10007 })
);
NAND3_X1 #() 
NAND3_X1_933_ (
  .A1({ S10006 }),
  .A2({ S10007 }),
  .A3({ S7106 }),
  .ZN({ S10008 })
);
AND2_X1 #() 
AND2_X1_51_ (
  .A1({ S10008 }),
  .A2({ S10005 }),
  .ZN({ S25957[414] })
);
NOR2_X1 #() 
NOR2_X1_188_ (
  .A1({ S7184 }),
  .A2({ S7196 }),
  .ZN({ S10009 })
);
INV_X1 #() 
INV_X1_279_ (
  .A({ S10009 }),
  .ZN({ S25957[605] })
);
NAND2_X1 #() 
NAND2_X1_817_ (
  .A1({ S4426 }),
  .A2({ S4428 }),
  .ZN({ S25957[765] })
);
NAND3_X1 #() 
NAND3_X1_934_ (
  .A1({ S7195 }),
  .A2({ S7192 }),
  .A3({ S25957[765] }),
  .ZN({ S10010 })
);
NAND4_X1 #() 
NAND4_X1_106_ (
  .A1({ S7152 }),
  .A2({ S7183 }),
  .A3({ S4426 }),
  .A4({ S4428 }),
  .ZN({ S10011 })
);
NAND2_X1 #() 
NAND2_X1_818_ (
  .A1({ S10011 }),
  .A2({ S10010 }),
  .ZN({ S25957[637] })
);
INV_X1 #() 
INV_X1_280_ (
  .A({ S25957[637] }),
  .ZN({ S10013 })
);
AOI21_X1 #() 
AOI21_X1_503_ (
  .A({ S6 }),
  .B1({ S9823 }),
  .B2({ S25957[529] }),
  .ZN({ S10014 })
);
INV_X1 #() 
INV_X1_281_ (
  .A({ S10014 }),
  .ZN({ S10015 })
);
NAND4_X1 #() 
NAND4_X1_107_ (
  .A1({ S10015 }),
  .A2({ S9867 }),
  .A3({ S9865 }),
  .A4({ S5128 }),
  .ZN({ S10016 })
);
NAND3_X1 #() 
NAND3_X1_935_ (
  .A1({ S9800 }),
  .A2({ S6 }),
  .A3({ S25957[530] }),
  .ZN({ S10017 })
);
OAI21_X1 #() 
OAI21_X1_457_ (
  .A({ S10017 }),
  .B1({ S9932 }),
  .B2({ S6 }),
  .ZN({ S10018 })
);
NOR2_X1 #() 
NOR2_X1_189_ (
  .A1({ S10018 }),
  .A2({ S5128 }),
  .ZN({ S10019 })
);
AOI21_X1 #() 
AOI21_X1_504_ (
  .A({ S10019 }),
  .B1({ S9922 }),
  .B2({ S9802 }),
  .ZN({ S10020 })
);
AOI22_X1 #() 
AOI22_X1_96_ (
  .A1({ S5362 }),
  .A2({ S5354 }),
  .B1({ S9787 }),
  .B2({ S9788 }),
  .ZN({ S10021 })
);
OAI21_X1 #() 
OAI21_X1_458_ (
  .A({ S6 }),
  .B1({ S9878 }),
  .B2({ S10021 }),
  .ZN({ S10023 })
);
AOI21_X1 #() 
AOI21_X1_505_ (
  .A({ S5128 }),
  .B1({ S9945 }),
  .B2({ S9800 }),
  .ZN({ S10024 })
);
AOI21_X1 #() 
AOI21_X1_506_ (
  .A({ S9790 }),
  .B1({ S10024 }),
  .B2({ S10023 }),
  .ZN({ S10025 })
);
AOI22_X1 #() 
AOI22_X1_97_ (
  .A1({ S10020 }),
  .A2({ S9790 }),
  .B1({ S10025 }),
  .B2({ S10016 }),
  .ZN({ S10026 })
);
INV_X1 #() 
INV_X1_282_ (
  .A({ S9797 }),
  .ZN({ S10027 })
);
OAI21_X1 #() 
OAI21_X1_459_ (
  .A({ S6 }),
  .B1({ S9875 }),
  .B2({ S10027 }),
  .ZN({ S10028 })
);
OAI211_X1 #() 
OAI211_X1_276_ (
  .A({ S10028 }),
  .B({ S25957[532] }),
  .C1({ S9824 }),
  .C2({ S6 }),
  .ZN({ S10029 })
);
NAND3_X1 #() 
NAND3_X1_936_ (
  .A1({ S9813 }),
  .A2({ S6 }),
  .A3({ S9800 }),
  .ZN({ S10030 })
);
AOI21_X1 #() 
AOI21_X1_507_ (
  .A({ S25957[532] }),
  .B1({ S25957[531] }),
  .B2({ S8137 }),
  .ZN({ S10031 })
);
AOI21_X1 #() 
AOI21_X1_508_ (
  .A({ S9790 }),
  .B1({ S10030 }),
  .B2({ S10031 }),
  .ZN({ S10032 })
);
OAI21_X1 #() 
OAI21_X1_460_ (
  .A({ S6 }),
  .B1({ S9789 }),
  .B2({ S25957[530] }),
  .ZN({ S10034 })
);
AOI21_X1 #() 
AOI21_X1_509_ (
  .A({ S8281 }),
  .B1({ S9801 }),
  .B2({ S9800 }),
  .ZN({ S10035 })
);
NOR2_X1 #() 
NOR2_X1_190_ (
  .A1({ S9823 }),
  .A2({ S25957[529] }),
  .ZN({ S10036 })
);
OAI21_X1 #() 
OAI21_X1_461_ (
  .A({ S25957[531] }),
  .B1({ S10035 }),
  .B2({ S10036 }),
  .ZN({ S10037 })
);
NAND3_X1 #() 
NAND3_X1_937_ (
  .A1({ S10037 }),
  .A2({ S5128 }),
  .A3({ S10034 }),
  .ZN({ S10038 })
);
NAND4_X1 #() 
NAND4_X1_108_ (
  .A1({ S26 }),
  .A2({ S9789 }),
  .A3({ S8281 }),
  .A4({ S25957[531] }),
  .ZN({ S10039 })
);
OAI21_X1 #() 
OAI21_X1_462_ (
  .A({ S10039 }),
  .B1({ S25957[531] }),
  .B2({ S9855 }),
  .ZN({ S10040 })
);
AOI21_X1 #() 
AOI21_X1_510_ (
  .A({ S25957[533] }),
  .B1({ S10040 }),
  .B2({ S25957[532] }),
  .ZN({ S10041 })
);
AOI22_X1 #() 
AOI22_X1_98_ (
  .A1({ S10041 }),
  .A2({ S10038 }),
  .B1({ S10032 }),
  .B2({ S10029 }),
  .ZN({ S10042 })
);
OR2_X1 #() 
OR2_X1_11_ (
  .A1({ S10042 }),
  .A2({ S25957[534] }),
  .ZN({ S10043 })
);
OAI211_X1 #() 
OAI211_X1_277_ (
  .A({ S10043 }),
  .B({ S25957[535] }),
  .C1({ S10026 }),
  .C2({ S7708 }),
  .ZN({ S10045 })
);
NAND4_X1 #() 
NAND4_X1_109_ (
  .A1({ S9822 }),
  .A2({ S9854 }),
  .A3({ S9797 }),
  .A4({ S25957[531] }),
  .ZN({ S10046 })
);
AOI21_X1 #() 
AOI21_X1_511_ (
  .A({ S25957[531] }),
  .B1({ S9889 }),
  .B2({ S25957[529] }),
  .ZN({ S10047 })
);
NAND4_X1 #() 
NAND4_X1_110_ (
  .A1({ S5285 }),
  .A2({ S5223 }),
  .A3({ S5220 }),
  .A4({ S5281 }),
  .ZN({ S10048 })
);
AOI22_X1 #() 
AOI22_X1_99_ (
  .A1({ S9971 }),
  .A2({ S10048 }),
  .B1({ S9789 }),
  .B2({ S25957[530] }),
  .ZN({ S10049 })
);
OAI21_X1 #() 
OAI21_X1_463_ (
  .A({ S5128 }),
  .B1({ S10049 }),
  .B2({ S10047 }),
  .ZN({ S10050 })
);
AOI21_X1 #() 
AOI21_X1_512_ (
  .A({ S10050 }),
  .B1({ S10046 }),
  .B2({ S9866 }),
  .ZN({ S10051 })
);
NAND3_X1 #() 
NAND3_X1_938_ (
  .A1({ S9801 }),
  .A2({ S25957[531] }),
  .A3({ S8281 }),
  .ZN({ S10052 })
);
NAND2_X1 #() 
NAND2_X1_819_ (
  .A1({ S10052 }),
  .A2({ S25957[532] }),
  .ZN({ S10053 })
);
AOI21_X1 #() 
AOI21_X1_513_ (
  .A({ S25957[531] }),
  .B1({ S9804 }),
  .B2({ S9835 }),
  .ZN({ S10054 })
);
OAI21_X1 #() 
OAI21_X1_464_ (
  .A({ S9790 }),
  .B1({ S10053 }),
  .B2({ S10054 }),
  .ZN({ S10056 })
);
AOI21_X1 #() 
AOI21_X1_514_ (
  .A({ S8281 }),
  .B1({ S26 }),
  .B2({ S9789 }),
  .ZN({ S10057 })
);
NAND2_X1 #() 
NAND2_X1_820_ (
  .A1({ S9843 }),
  .A2({ S6 }),
  .ZN({ S10058 })
);
OAI21_X1 #() 
OAI21_X1_465_ (
  .A({ S25957[531] }),
  .B1({ S9800 }),
  .B2({ S25957[530] }),
  .ZN({ S10059 })
);
OAI21_X1 #() 
OAI21_X1_466_ (
  .A({ S10058 }),
  .B1({ S10057 }),
  .B2({ S10059 }),
  .ZN({ S10060 })
);
OAI21_X1 #() 
OAI21_X1_467_ (
  .A({ S10048 }),
  .B1({ S9886 }),
  .B2({ S9793 }),
  .ZN({ S10061 })
);
NAND2_X1 #() 
NAND2_X1_821_ (
  .A1({ S10061 }),
  .A2({ S5128 }),
  .ZN({ S10062 })
);
OAI211_X1 #() 
OAI211_X1_278_ (
  .A({ S25957[533] }),
  .B({ S10062 }),
  .C1({ S10060 }),
  .C2({ S5128 }),
  .ZN({ S10063 })
);
OAI211_X1 #() 
OAI211_X1_279_ (
  .A({ S10063 }),
  .B({ S25957[534] }),
  .C1({ S10051 }),
  .C2({ S10056 }),
  .ZN({ S10064 })
);
NAND3_X1 #() 
NAND3_X1_939_ (
  .A1({ S9829 }),
  .A2({ S25957[531] }),
  .A3({ S9842 }),
  .ZN({ S10065 })
);
NAND2_X1 #() 
NAND2_X1_822_ (
  .A1({ S26 }),
  .A2({ S9789 }),
  .ZN({ S10067 })
);
NAND2_X1 #() 
NAND2_X1_823_ (
  .A1({ S10067 }),
  .A2({ S9871 }),
  .ZN({ S10068 })
);
NAND3_X1 #() 
NAND3_X1_940_ (
  .A1({ S10065 }),
  .A2({ S25957[532] }),
  .A3({ S10068 }),
  .ZN({ S10069 })
);
NOR2_X1 #() 
NOR2_X1_191_ (
  .A1({ S9801 }),
  .A2({ S6 }),
  .ZN({ S10070 })
);
NOR2_X1 #() 
NOR2_X1_192_ (
  .A1({ S9841 }),
  .A2({ S9837 }),
  .ZN({ S10071 })
);
AOI21_X1 #() 
AOI21_X1_515_ (
  .A({ S10070 }),
  .B1({ S6 }),
  .B2({ S10071 }),
  .ZN({ S10072 })
);
OAI21_X1 #() 
OAI21_X1_468_ (
  .A({ S10069 }),
  .B1({ S25957[532] }),
  .B2({ S10072 }),
  .ZN({ S10073 })
);
NAND2_X1 #() 
NAND2_X1_824_ (
  .A1({ S9854 }),
  .A2({ S25957[529] }),
  .ZN({ S10074 })
);
NOR2_X1 #() 
NOR2_X1_193_ (
  .A1({ S10074 }),
  .A2({ S9853 }),
  .ZN({ S10075 })
);
OAI21_X1 #() 
OAI21_X1_469_ (
  .A({ S25957[532] }),
  .B1({ S9885 }),
  .B2({ S25957[530] }),
  .ZN({ S10076 })
);
OAI22_X1 #() 
OAI22_X1_22_ (
  .A1({ S10076 }),
  .A2({ S10047 }),
  .B1({ S10075 }),
  .B2({ S9913 }),
  .ZN({ S10078 })
);
AOI21_X1 #() 
AOI21_X1_516_ (
  .A({ S25957[534] }),
  .B1({ S10078 }),
  .B2({ S25957[533] }),
  .ZN({ S10079 })
);
OAI21_X1 #() 
OAI21_X1_470_ (
  .A({ S10079 }),
  .B1({ S25957[533] }),
  .B2({ S10073 }),
  .ZN({ S10080 })
);
NAND3_X1 #() 
NAND3_X1_941_ (
  .A1({ S10064 }),
  .A2({ S10080 }),
  .A3({ S4924 }),
  .ZN({ S10081 })
);
NAND2_X1 #() 
NAND2_X1_825_ (
  .A1({ S10045 }),
  .A2({ S10081 }),
  .ZN({ S10082 })
);
NAND2_X1 #() 
NAND2_X1_826_ (
  .A1({ S10082 }),
  .A2({ S10013 }),
  .ZN({ S10083 })
);
NAND3_X1 #() 
NAND3_X1_942_ (
  .A1({ S10045 }),
  .A2({ S10081 }),
  .A3({ S25957[637] }),
  .ZN({ S10084 })
);
NAND3_X1 #() 
NAND3_X1_943_ (
  .A1({ S10083 }),
  .A2({ S10084 }),
  .A3({ S25957[605] }),
  .ZN({ S10085 })
);
NAND2_X1 #() 
NAND2_X1_827_ (
  .A1({ S10083 }),
  .A2({ S10084 }),
  .ZN({ S25957[509] })
);
NAND2_X1 #() 
NAND2_X1_828_ (
  .A1({ S25957[509] }),
  .A2({ S10009 }),
  .ZN({ S10086 })
);
NAND3_X1 #() 
NAND3_X1_944_ (
  .A1({ S10086 }),
  .A2({ S25957[669] }),
  .A3({ S10085 }),
  .ZN({ S10088 })
);
NAND2_X1 #() 
NAND2_X1_829_ (
  .A1({ S25957[509] }),
  .A2({ S25957[605] }),
  .ZN({ S10089 })
);
NAND3_X1 #() 
NAND3_X1_945_ (
  .A1({ S10083 }),
  .A2({ S10084 }),
  .A3({ S10009 }),
  .ZN({ S10090 })
);
NAND3_X1 #() 
NAND3_X1_946_ (
  .A1({ S10089 }),
  .A2({ S10090 }),
  .A3({ S6306 }),
  .ZN({ S10091 })
);
NAND2_X1 #() 
NAND2_X1_830_ (
  .A1({ S10088 }),
  .A2({ S10091 }),
  .ZN({ S25957[413] })
);
NAND2_X1 #() 
NAND2_X1_831_ (
  .A1({ S7269 }),
  .A2({ S7266 }),
  .ZN({ S10092 })
);
INV_X1 #() 
INV_X1_283_ (
  .A({ S10092 }),
  .ZN({ S25957[572] })
);
NAND2_X1 #() 
NAND2_X1_832_ (
  .A1({ S4494 }),
  .A2({ S4496 }),
  .ZN({ S10093 })
);
NAND2_X1 #() 
NAND2_X1_833_ (
  .A1({ S10017 }),
  .A2({ S25957[532] }),
  .ZN({ S10094 })
);
AOI21_X1 #() 
AOI21_X1_517_ (
  .A({ S10094 }),
  .B1({ S9843 }),
  .B2({ S25957[531] }),
  .ZN({ S10095 })
);
NAND2_X1 #() 
NAND2_X1_834_ (
  .A1({ S25 }),
  .A2({ S6 }),
  .ZN({ S10097 })
);
AOI21_X1 #() 
AOI21_X1_518_ (
  .A({ S25957[532] }),
  .B1({ S10097 }),
  .B2({ S10039 }),
  .ZN({ S10098 })
);
OAI21_X1 #() 
OAI21_X1_471_ (
  .A({ S25957[533] }),
  .B1({ S10095 }),
  .B2({ S10098 }),
  .ZN({ S10099 })
);
OAI21_X1 #() 
OAI21_X1_472_ (
  .A({ S6 }),
  .B1({ S10036 }),
  .B2({ S9948 }),
  .ZN({ S10100 })
);
NAND2_X1 #() 
NAND2_X1_835_ (
  .A1({ S9815 }),
  .A2({ S26 }),
  .ZN({ S10101 })
);
AOI21_X1 #() 
AOI21_X1_519_ (
  .A({ S25957[532] }),
  .B1({ S10100 }),
  .B2({ S10101 }),
  .ZN({ S10102 })
);
NAND4_X1 #() 
NAND4_X1_111_ (
  .A1({ S9807 }),
  .A2({ S9823 }),
  .A3({ S25957[531] }),
  .A4({ S9865 }),
  .ZN({ S10103 })
);
AND3_X1 #() 
AND3_X1_37_ (
  .A1({ S10103 }),
  .A2({ S10030 }),
  .A3({ S25957[532] }),
  .ZN({ S10104 })
);
OAI21_X1 #() 
OAI21_X1_473_ (
  .A({ S9790 }),
  .B1({ S10102 }),
  .B2({ S10104 }),
  .ZN({ S10105 })
);
NAND3_X1 #() 
NAND3_X1_947_ (
  .A1({ S10105 }),
  .A2({ S10099 }),
  .A3({ S7708 }),
  .ZN({ S10106 })
);
AND2_X1 #() 
AND2_X1_52_ (
  .A1({ S8281 }),
  .A2({ S143 }),
  .ZN({ S10108 })
);
NAND4_X1 #() 
NAND4_X1_112_ (
  .A1({ S26 }),
  .A2({ S9789 }),
  .A3({ S8281 }),
  .A4({ S6 }),
  .ZN({ S10109 })
);
NAND4_X1 #() 
NAND4_X1_113_ (
  .A1({ S10046 }),
  .A2({ S10109 }),
  .A3({ S5128 }),
  .A4({ S10017 }),
  .ZN({ S10110 })
);
OAI211_X1 #() 
OAI211_X1_280_ (
  .A({ S10110 }),
  .B({ S25957[533] }),
  .C1({ S5128 }),
  .C2({ S10108 }),
  .ZN({ S10111 })
);
NAND2_X1 #() 
NAND2_X1_836_ (
  .A1({ S9971 }),
  .A2({ S5128 }),
  .ZN({ S10112 })
);
NAND3_X1 #() 
NAND3_X1_948_ (
  .A1({ S9835 }),
  .A2({ S6 }),
  .A3({ S9797 }),
  .ZN({ S10113 })
);
INV_X1 #() 
INV_X1_284_ (
  .A({ S10113 }),
  .ZN({ S10114 })
);
NAND3_X1 #() 
NAND3_X1_949_ (
  .A1({ S9888 }),
  .A2({ S6 }),
  .A3({ S9813 }),
  .ZN({ S10115 })
);
NAND3_X1 #() 
NAND3_X1_950_ (
  .A1({ S10115 }),
  .A2({ S25957[532] }),
  .A3({ S9868 }),
  .ZN({ S10116 })
);
OAI211_X1 #() 
OAI211_X1_281_ (
  .A({ S10116 }),
  .B({ S9790 }),
  .C1({ S10112 }),
  .C2({ S10114 }),
  .ZN({ S10117 })
);
NAND3_X1 #() 
NAND3_X1_951_ (
  .A1({ S10117 }),
  .A2({ S10111 }),
  .A3({ S25957[534] }),
  .ZN({ S10119 })
);
NAND3_X1 #() 
NAND3_X1_952_ (
  .A1({ S10106 }),
  .A2({ S4924 }),
  .A3({ S10119 }),
  .ZN({ S10120 })
);
NAND3_X1 #() 
NAND3_X1_953_ (
  .A1({ S9813 }),
  .A2({ S6 }),
  .A3({ S9797 }),
  .ZN({ S10121 })
);
NAND3_X1 #() 
NAND3_X1_954_ (
  .A1({ S9808 }),
  .A2({ S10121 }),
  .A3({ S5128 }),
  .ZN({ S10122 })
);
OAI211_X1 #() 
OAI211_X1_282_ (
  .A({ S10030 }),
  .B({ S25957[532] }),
  .C1({ S6 }),
  .C2({ S9855 }),
  .ZN({ S10123 })
);
NAND3_X1 #() 
NAND3_X1_955_ (
  .A1({ S10123 }),
  .A2({ S10122 }),
  .A3({ S9790 }),
  .ZN({ S10124 })
);
NAND2_X1 #() 
NAND2_X1_837_ (
  .A1({ S9838 }),
  .A2({ S6 }),
  .ZN({ S10125 })
);
NAND3_X1 #() 
NAND3_X1_956_ (
  .A1({ S10125 }),
  .A2({ S25957[532] }),
  .A3({ S10052 }),
  .ZN({ S10126 })
);
NAND3_X1 #() 
NAND3_X1_957_ (
  .A1({ S9807 }),
  .A2({ S6 }),
  .A3({ S9837 }),
  .ZN({ S10127 })
);
NAND3_X1 #() 
NAND3_X1_958_ (
  .A1({ S9816 }),
  .A2({ S5128 }),
  .A3({ S10127 }),
  .ZN({ S10128 })
);
NAND3_X1 #() 
NAND3_X1_959_ (
  .A1({ S10128 }),
  .A2({ S25957[533] }),
  .A3({ S10126 }),
  .ZN({ S10130 })
);
NAND3_X1 #() 
NAND3_X1_960_ (
  .A1({ S10130 }),
  .A2({ S10124 }),
  .A3({ S25957[534] }),
  .ZN({ S10131 })
);
AOI21_X1 #() 
AOI21_X1_520_ (
  .A({ S25957[531] }),
  .B1({ S9827 }),
  .B2({ S9804 }),
  .ZN({ S10132 })
);
NAND4_X1 #() 
NAND4_X1_114_ (
  .A1({ S9822 }),
  .A2({ S9801 }),
  .A3({ S9865 }),
  .A4({ S25957[531] }),
  .ZN({ S10133 })
);
NAND2_X1 #() 
NAND2_X1_838_ (
  .A1({ S10133 }),
  .A2({ S5128 }),
  .ZN({ S10134 })
);
NAND4_X1 #() 
NAND4_X1_115_ (
  .A1({ S9837 }),
  .A2({ S8281 }),
  .A3({ S8132 }),
  .A4({ S8136 }),
  .ZN({ S10135 })
);
NAND3_X1 #() 
NAND3_X1_961_ (
  .A1({ S10135 }),
  .A2({ S25957[531] }),
  .A3({ S9801 }),
  .ZN({ S10136 })
);
AOI22_X1 #() 
AOI22_X1_100_ (
  .A1({ S9865 }),
  .A2({ S9800 }),
  .B1({ S25957[529] }),
  .B2({ S25957[530] }),
  .ZN({ S10137 })
);
OAI211_X1 #() 
OAI211_X1_283_ (
  .A({ S10136 }),
  .B({ S25957[532] }),
  .C1({ S10137 }),
  .C2({ S25957[531] }),
  .ZN({ S10138 })
);
OAI211_X1 #() 
OAI211_X1_284_ (
  .A({ S10138 }),
  .B({ S25957[533] }),
  .C1({ S10132 }),
  .C2({ S10134 }),
  .ZN({ S10139 })
);
NAND2_X1 #() 
NAND2_X1_839_ (
  .A1({ S9865 }),
  .A2({ S25957[531] }),
  .ZN({ S10141 })
);
OAI21_X1 #() 
OAI21_X1_474_ (
  .A({ S6 }),
  .B1({ S9932 }),
  .B2({ S9798 }),
  .ZN({ S10142 })
);
OAI21_X1 #() 
OAI21_X1_475_ (
  .A({ S10142 }),
  .B1({ S25957[529] }),
  .B2({ S10141 }),
  .ZN({ S10143 })
);
OAI21_X1 #() 
OAI21_X1_476_ (
  .A({ S25957[531] }),
  .B1({ S9798 }),
  .B2({ S9852 }),
  .ZN({ S10144 })
);
OAI211_X1 #() 
OAI211_X1_285_ (
  .A({ S10144 }),
  .B({ S25957[532] }),
  .C1({ S10034 }),
  .C2({ S9798 }),
  .ZN({ S10145 })
);
OAI211_X1 #() 
OAI211_X1_286_ (
  .A({ S9790 }),
  .B({ S10145 }),
  .C1({ S10143 }),
  .C2({ S25957[532] }),
  .ZN({ S10146 })
);
NAND3_X1 #() 
NAND3_X1_962_ (
  .A1({ S10146 }),
  .A2({ S10139 }),
  .A3({ S7708 }),
  .ZN({ S10147 })
);
NAND3_X1 #() 
NAND3_X1_963_ (
  .A1({ S10147 }),
  .A2({ S25957[535] }),
  .A3({ S10131 }),
  .ZN({ S10148 })
);
NAND3_X1 #() 
NAND3_X1_964_ (
  .A1({ S10148 }),
  .A2({ S10120 }),
  .A3({ S10093 }),
  .ZN({ S10149 })
);
AOI21_X1 #() 
AOI21_X1_521_ (
  .A({ S10093 }),
  .B1({ S10148 }),
  .B2({ S10120 }),
  .ZN({ S10150 })
);
INV_X1 #() 
INV_X1_285_ (
  .A({ S10150 }),
  .ZN({ S10152 })
);
NAND3_X1 #() 
NAND3_X1_965_ (
  .A1({ S10152 }),
  .A2({ S25957[572] }),
  .A3({ S10149 }),
  .ZN({ S10153 })
);
INV_X1 #() 
INV_X1_286_ (
  .A({ S10149 }),
  .ZN({ S10154 })
);
OAI21_X1 #() 
OAI21_X1_477_ (
  .A({ S10092 }),
  .B1({ S10154 }),
  .B2({ S10150 }),
  .ZN({ S10155 })
);
NAND3_X1 #() 
NAND3_X1_966_ (
  .A1({ S10153 }),
  .A2({ S10155 }),
  .A3({ S25957[540] }),
  .ZN({ S10156 })
);
OAI21_X1 #() 
OAI21_X1_478_ (
  .A({ S25957[572] }),
  .B1({ S10154 }),
  .B2({ S10150 }),
  .ZN({ S10157 })
);
NAND3_X1 #() 
NAND3_X1_967_ (
  .A1({ S10152 }),
  .A2({ S10092 }),
  .A3({ S10149 }),
  .ZN({ S10158 })
);
NAND3_X1 #() 
NAND3_X1_968_ (
  .A1({ S10158 }),
  .A2({ S10157 }),
  .A3({ S9063 }),
  .ZN({ S10159 })
);
NAND2_X1 #() 
NAND2_X1_840_ (
  .A1({ S10156 }),
  .A2({ S10159 }),
  .ZN({ S25957[412] })
);
NAND2_X1 #() 
NAND2_X1_841_ (
  .A1({ S4589 }),
  .A2({ S4592 }),
  .ZN({ S25957[699] })
);
NAND2_X1 #() 
NAND2_X1_842_ (
  .A1({ S4591 }),
  .A2({ S4590 }),
  .ZN({ S25957[763] })
);
NAND2_X1 #() 
NAND2_X1_843_ (
  .A1({ S7335 }),
  .A2({ S7331 }),
  .ZN({ S10161 })
);
XOR2_X1 #() 
XOR2_X1_19_ (
  .A({ S10161 }),
  .B({ S25957[763] }),
  .Z({ S25957[635] })
);
NAND3_X1 #() 
NAND3_X1_969_ (
  .A1({ S9835 }),
  .A2({ S25957[531] }),
  .A3({ S9797 }),
  .ZN({ S10162 })
);
INV_X1 #() 
INV_X1_287_ (
  .A({ S10162 }),
  .ZN({ S10163 })
);
OAI21_X1 #() 
OAI21_X1_479_ (
  .A({ S5128 }),
  .B1({ S9830 }),
  .B2({ S10163 }),
  .ZN({ S10164 })
);
AOI21_X1 #() 
AOI21_X1_522_ (
  .A({ S5128 }),
  .B1({ S10067 }),
  .B2({ S9815 }),
  .ZN({ S10165 })
);
NAND2_X1 #() 
NAND2_X1_844_ (
  .A1({ S10165 }),
  .A2({ S9938 }),
  .ZN({ S10166 })
);
NAND3_X1 #() 
NAND3_X1_970_ (
  .A1({ S10164 }),
  .A2({ S9790 }),
  .A3({ S10166 }),
  .ZN({ S10167 })
);
NAND2_X1 #() 
NAND2_X1_845_ (
  .A1({ S9807 }),
  .A2({ S6 }),
  .ZN({ S10168 })
);
AOI21_X1 #() 
AOI21_X1_523_ (
  .A({ S9837 }),
  .B1({ S10168 }),
  .B2({ S9822 }),
  .ZN({ S10170 })
);
NAND3_X1 #() 
NAND3_X1_971_ (
  .A1({ S9957 }),
  .A2({ S25957[531] }),
  .A3({ S25957[530] }),
  .ZN({ S10171 })
);
NAND3_X1 #() 
NAND3_X1_972_ (
  .A1({ S9802 }),
  .A2({ S10171 }),
  .A3({ S25957[532] }),
  .ZN({ S10172 })
);
OAI211_X1 #() 
OAI211_X1_287_ (
  .A({ S10172 }),
  .B({ S25957[533] }),
  .C1({ S25957[532] }),
  .C2({ S10170 }),
  .ZN({ S10173 })
);
NAND3_X1 #() 
NAND3_X1_973_ (
  .A1({ S10167 }),
  .A2({ S7708 }),
  .A3({ S10173 }),
  .ZN({ S10174 })
);
NAND3_X1 #() 
NAND3_X1_974_ (
  .A1({ S9789 }),
  .A2({ S6 }),
  .A3({ S9865 }),
  .ZN({ S10175 })
);
NOR2_X1 #() 
NOR2_X1_194_ (
  .A1({ S10175 }),
  .A2({ S5128 }),
  .ZN({ S10176 })
);
INV_X1 #() 
INV_X1_288_ (
  .A({ S10176 }),
  .ZN({ S10177 })
);
NAND2_X1 #() 
NAND2_X1_846_ (
  .A1({ S9826 }),
  .A2({ S10103 }),
  .ZN({ S10178 })
);
AOI21_X1 #() 
AOI21_X1_524_ (
  .A({ S25957[533] }),
  .B1({ S10178 }),
  .B2({ S10177 }),
  .ZN({ S10179 })
);
AOI21_X1 #() 
AOI21_X1_525_ (
  .A({ S25957[531] }),
  .B1({ S26 }),
  .B2({ S9841 }),
  .ZN({ S10181 })
);
NAND3_X1 #() 
NAND3_X1_975_ (
  .A1({ S9841 }),
  .A2({ S25957[531] }),
  .A3({ S9837 }),
  .ZN({ S10182 })
);
NAND2_X1 #() 
NAND2_X1_847_ (
  .A1({ S10182 }),
  .A2({ S5128 }),
  .ZN({ S10183 })
);
OAI21_X1 #() 
OAI21_X1_480_ (
  .A({ S25957[533] }),
  .B1({ S10183 }),
  .B2({ S10181 }),
  .ZN({ S10184 })
);
AOI21_X1 #() 
AOI21_X1_526_ (
  .A({ S10184 }),
  .B1({ S9955 }),
  .B2({ S9795 }),
  .ZN({ S10185 })
);
OAI21_X1 #() 
OAI21_X1_481_ (
  .A({ S25957[534] }),
  .B1({ S10179 }),
  .B2({ S10185 }),
  .ZN({ S10186 })
);
NAND3_X1 #() 
NAND3_X1_976_ (
  .A1({ S10186 }),
  .A2({ S4924 }),
  .A3({ S10174 }),
  .ZN({ S10187 })
);
NAND3_X1 #() 
NAND3_X1_977_ (
  .A1({ S26 }),
  .A2({ S8281 }),
  .A3({ S9789 }),
  .ZN({ S10188 })
);
NAND3_X1 #() 
NAND3_X1_978_ (
  .A1({ S10188 }),
  .A2({ S25957[531] }),
  .A3({ S9838 }),
  .ZN({ S10189 })
);
AOI21_X1 #() 
AOI21_X1_527_ (
  .A({ S5128 }),
  .B1({ S9921 }),
  .B2({ S6 }),
  .ZN({ S10190 })
);
NAND2_X1 #() 
NAND2_X1_848_ (
  .A1({ S10190 }),
  .A2({ S10189 }),
  .ZN({ S10192 })
);
NAND3_X1 #() 
NAND3_X1_979_ (
  .A1({ S9791 }),
  .A2({ S6 }),
  .A3({ S9813 }),
  .ZN({ S10193 })
);
AOI21_X1 #() 
AOI21_X1_528_ (
  .A({ S25957[532] }),
  .B1({ S9945 }),
  .B2({ S9912 }),
  .ZN({ S10194 })
);
NAND2_X1 #() 
NAND2_X1_849_ (
  .A1({ S10193 }),
  .A2({ S10194 }),
  .ZN({ S10195 })
);
NAND3_X1 #() 
NAND3_X1_980_ (
  .A1({ S10192 }),
  .A2({ S10195 }),
  .A3({ S25957[533] }),
  .ZN({ S10196 })
);
NAND2_X1 #() 
NAND2_X1_850_ (
  .A1({ S9813 }),
  .A2({ S25957[531] }),
  .ZN({ S10197 })
);
NAND3_X1 #() 
NAND3_X1_981_ (
  .A1({ S9800 }),
  .A2({ S6 }),
  .A3({ S9865 }),
  .ZN({ S10198 })
);
OAI211_X1 #() 
OAI211_X1_288_ (
  .A({ S5128 }),
  .B({ S10198 }),
  .C1({ S10057 }),
  .C2({ S10197 }),
  .ZN({ S10199 })
);
OAI211_X1 #() 
OAI211_X1_289_ (
  .A({ S25957[532] }),
  .B({ S10121 }),
  .C1({ S9954 }),
  .C2({ S6 }),
  .ZN({ S10200 })
);
NAND3_X1 #() 
NAND3_X1_982_ (
  .A1({ S10199 }),
  .A2({ S10200 }),
  .A3({ S9790 }),
  .ZN({ S10201 })
);
NAND3_X1 #() 
NAND3_X1_983_ (
  .A1({ S10196 }),
  .A2({ S7708 }),
  .A3({ S10201 }),
  .ZN({ S10203 })
);
AOI21_X1 #() 
AOI21_X1_529_ (
  .A({ S10014 }),
  .B1({ S9930 }),
  .B2({ S9829 }),
  .ZN({ S10204 })
);
OAI22_X1 #() 
OAI22_X1_23_ (
  .A1({ S10204 }),
  .A2({ S5128 }),
  .B1({ S10112 }),
  .B2({ S9915 }),
  .ZN({ S10205 })
);
NAND3_X1 #() 
NAND3_X1_984_ (
  .A1({ S26 }),
  .A2({ S9854 }),
  .A3({ S9841 }),
  .ZN({ S10206 })
);
OAI221_X1 #() 
OAI221_X1_17_ (
  .A({ S5128 }),
  .B1({ S9924 }),
  .B2({ S9875 }),
  .C1({ S6 }),
  .C2({ S10206 }),
  .ZN({ S10207 })
);
NAND3_X1 #() 
NAND3_X1_985_ (
  .A1({ S9965 }),
  .A2({ S6 }),
  .A3({ S9801 }),
  .ZN({ S10208 })
);
NAND2_X1 #() 
NAND2_X1_851_ (
  .A1({ S10208 }),
  .A2({ S10101 }),
  .ZN({ S10209 })
);
AOI21_X1 #() 
AOI21_X1_530_ (
  .A({ S9790 }),
  .B1({ S10209 }),
  .B2({ S25957[532] }),
  .ZN({ S10210 })
);
AOI22_X1 #() 
AOI22_X1_101_ (
  .A1({ S9790 }),
  .A2({ S10205 }),
  .B1({ S10210 }),
  .B2({ S10207 }),
  .ZN({ S10211 })
);
OAI211_X1 #() 
OAI211_X1_290_ (
  .A({ S25957[535] }),
  .B({ S10203 }),
  .C1({ S10211 }),
  .C2({ S7708 }),
  .ZN({ S10212 })
);
NAND3_X1 #() 
NAND3_X1_986_ (
  .A1({ S10187 }),
  .A2({ S10212 }),
  .A3({ S25957[635] }),
  .ZN({ S10214 })
);
INV_X1 #() 
INV_X1_289_ (
  .A({ S25957[635] }),
  .ZN({ S10215 })
);
OAI21_X1 #() 
OAI21_X1_482_ (
  .A({ S6 }),
  .B1({ S10057 }),
  .B2({ S9889 }),
  .ZN({ S10216 })
);
NAND2_X1 #() 
NAND2_X1_852_ (
  .A1({ S10216 }),
  .A2({ S10162 }),
  .ZN({ S10217 })
);
AOI22_X1 #() 
AOI22_X1_102_ (
  .A1({ S10217 }),
  .A2({ S5128 }),
  .B1({ S10165 }),
  .B2({ S9938 }),
  .ZN({ S10218 })
);
NAND2_X1 #() 
NAND2_X1_853_ (
  .A1({ S10173 }),
  .A2({ S7708 }),
  .ZN({ S10219 })
);
AOI21_X1 #() 
AOI21_X1_531_ (
  .A({ S10219 }),
  .B1({ S10218 }),
  .B2({ S9790 }),
  .ZN({ S10220 })
);
NAND4_X1 #() 
NAND4_X1_116_ (
  .A1({ S9822 }),
  .A2({ S9807 }),
  .A3({ S6 }),
  .A4({ S25957[528] }),
  .ZN({ S10221 })
);
AOI21_X1 #() 
AOI21_X1_532_ (
  .A({ S25957[532] }),
  .B1({ S9879 }),
  .B2({ S10221 }),
  .ZN({ S10222 })
);
OAI21_X1 #() 
OAI21_X1_483_ (
  .A({ S9790 }),
  .B1({ S10222 }),
  .B2({ S10176 }),
  .ZN({ S10223 })
);
NAND2_X1 #() 
NAND2_X1_854_ (
  .A1({ S9955 }),
  .A2({ S9795 }),
  .ZN({ S10225 })
);
OAI211_X1 #() 
OAI211_X1_291_ (
  .A({ S10225 }),
  .B({ S25957[533] }),
  .C1({ S10181 }),
  .C2({ S10183 }),
  .ZN({ S10226 })
);
AOI21_X1 #() 
AOI21_X1_533_ (
  .A({ S7708 }),
  .B1({ S10223 }),
  .B2({ S10226 }),
  .ZN({ S10227 })
);
OAI21_X1 #() 
OAI21_X1_484_ (
  .A({ S4924 }),
  .B1({ S10220 }),
  .B2({ S10227 }),
  .ZN({ S10228 })
);
AND3_X1 #() 
AND3_X1_38_ (
  .A1({ S10196 }),
  .A2({ S7708 }),
  .A3({ S10201 }),
  .ZN({ S10229 })
);
NAND2_X1 #() 
NAND2_X1_855_ (
  .A1({ S9930 }),
  .A2({ S9829 }),
  .ZN({ S10230 })
);
AOI21_X1 #() 
AOI21_X1_534_ (
  .A({ S5128 }),
  .B1({ S10230 }),
  .B2({ S10015 }),
  .ZN({ S10231 })
);
NOR2_X1 #() 
NOR2_X1_195_ (
  .A1({ S9915 }),
  .A2({ S10112 }),
  .ZN({ S10232 })
);
OAI21_X1 #() 
OAI21_X1_485_ (
  .A({ S9790 }),
  .B1({ S10231 }),
  .B2({ S10232 }),
  .ZN({ S10233 })
);
NAND2_X1 #() 
NAND2_X1_856_ (
  .A1({ S10209 }),
  .A2({ S25957[532] }),
  .ZN({ S10234 })
);
NAND3_X1 #() 
NAND3_X1_987_ (
  .A1({ S10234 }),
  .A2({ S10207 }),
  .A3({ S25957[533] }),
  .ZN({ S10236 })
);
AOI21_X1 #() 
AOI21_X1_535_ (
  .A({ S7708 }),
  .B1({ S10233 }),
  .B2({ S10236 }),
  .ZN({ S10237 })
);
OAI21_X1 #() 
OAI21_X1_486_ (
  .A({ S25957[535] }),
  .B1({ S10237 }),
  .B2({ S10229 }),
  .ZN({ S10238 })
);
NAND3_X1 #() 
NAND3_X1_988_ (
  .A1({ S10228 }),
  .A2({ S10238 }),
  .A3({ S10215 }),
  .ZN({ S10239 })
);
AOI21_X1 #() 
AOI21_X1_536_ (
  .A({ S25957[699] }),
  .B1({ S10239 }),
  .B2({ S10214 }),
  .ZN({ S10240 })
);
INV_X1 #() 
INV_X1_290_ (
  .A({ S25957[699] }),
  .ZN({ S10241 })
);
NAND3_X1 #() 
NAND3_X1_989_ (
  .A1({ S10187 }),
  .A2({ S10212 }),
  .A3({ S10215 }),
  .ZN({ S10242 })
);
NAND3_X1 #() 
NAND3_X1_990_ (
  .A1({ S10228 }),
  .A2({ S10238 }),
  .A3({ S25957[635] }),
  .ZN({ S10243 })
);
AOI21_X1 #() 
AOI21_X1_537_ (
  .A({ S10241 }),
  .B1({ S10243 }),
  .B2({ S10242 }),
  .ZN({ S10244 })
);
OAI21_X1 #() 
OAI21_X1_487_ (
  .A({ S25957[539] }),
  .B1({ S10240 }),
  .B2({ S10244 }),
  .ZN({ S10245 })
);
NAND3_X1 #() 
NAND3_X1_991_ (
  .A1({ S10243 }),
  .A2({ S10242 }),
  .A3({ S10241 }),
  .ZN({ S10247 })
);
NAND3_X1 #() 
NAND3_X1_992_ (
  .A1({ S10239 }),
  .A2({ S10214 }),
  .A3({ S25957[699] }),
  .ZN({ S10248 })
);
NAND3_X1 #() 
NAND3_X1_993_ (
  .A1({ S10247 }),
  .A2({ S10248 }),
  .A3({ S15 }),
  .ZN({ S10249 })
);
NAND2_X1 #() 
NAND2_X1_857_ (
  .A1({ S10245 }),
  .A2({ S10249 }),
  .ZN({ S28 })
);
AOI21_X1 #() 
AOI21_X1_538_ (
  .A({ S15 }),
  .B1({ S10247 }),
  .B2({ S10248 }),
  .ZN({ S10250 })
);
AND3_X1 #() 
AND3_X1_39_ (
  .A1({ S10248 }),
  .A2({ S10247 }),
  .A3({ S15 }),
  .ZN({ S10251 })
);
NOR2_X1 #() 
NOR2_X1_196_ (
  .A1({ S10251 }),
  .A2({ S10250 }),
  .ZN({ S25957[411] })
);
XNOR2_X1 #() 
XNOR2_X1_28_ (
  .A({ S25957[856] }),
  .B({ S4597 }),
  .ZN({ S25957[824] })
);
NAND2_X1 #() 
NAND2_X1_858_ (
  .A1({ S4671 }),
  .A2({ S4645 }),
  .ZN({ S25957[760] })
);
NAND2_X1 #() 
NAND2_X1_859_ (
  .A1({ S7382 }),
  .A2({ S7362 }),
  .ZN({ S10252 })
);
XNOR2_X1 #() 
XNOR2_X1_29_ (
  .A({ S10252 }),
  .B({ S25957[760] }),
  .ZN({ S25957[632] })
);
OR2_X1 #() 
OR2_X1_12_ (
  .A1({ S25957[632] }),
  .A2({ S25957[824] }),
  .ZN({ S10254 })
);
NAND2_X1 #() 
NAND2_X1_860_ (
  .A1({ S25957[632] }),
  .A2({ S25957[824] }),
  .ZN({ S10255 })
);
NAND2_X1 #() 
NAND2_X1_861_ (
  .A1({ S10254 }),
  .A2({ S10255 }),
  .ZN({ S10256 })
);
NAND2_X1 #() 
NAND2_X1_862_ (
  .A1({ S6185 }),
  .A2({ S6187 }),
  .ZN({ S25957[728] })
);
INV_X1 #() 
INV_X1_291_ (
  .A({ S25957[728] }),
  .ZN({ S10257 })
);
NAND4_X1 #() 
NAND4_X1_117_ (
  .A1({ S9801 }),
  .A2({ S9854 }),
  .A3({ S9800 }),
  .A4({ S25957[531] }),
  .ZN({ S10258 })
);
AND2_X1 #() 
AND2_X1_53_ (
  .A1({ S9838 }),
  .A2({ S9842 }),
  .ZN({ S10259 })
);
OAI211_X1 #() 
OAI211_X1_292_ (
  .A({ S10258 }),
  .B({ S5128 }),
  .C1({ S10259 }),
  .C2({ S25957[531] }),
  .ZN({ S10260 })
);
NAND2_X1 #() 
NAND2_X1_863_ (
  .A1({ S9827 }),
  .A2({ S25957[531] }),
  .ZN({ S10261 })
);
NOR2_X1 #() 
NOR2_X1_197_ (
  .A1({ S9813 }),
  .A2({ S25957[531] }),
  .ZN({ S10263 })
);
INV_X1 #() 
INV_X1_292_ (
  .A({ S10263 }),
  .ZN({ S10264 })
);
NAND4_X1 #() 
NAND4_X1_118_ (
  .A1({ S10261 }),
  .A2({ S10264 }),
  .A3({ S25957[532] }),
  .A4({ S9802 }),
  .ZN({ S10265 })
);
NAND3_X1 #() 
NAND3_X1_994_ (
  .A1({ S10260 }),
  .A2({ S10265 }),
  .A3({ S9790 }),
  .ZN({ S10266 })
);
NAND3_X1 #() 
NAND3_X1_995_ (
  .A1({ S10068 }),
  .A2({ S9947 }),
  .A3({ S5128 }),
  .ZN({ S10267 })
);
AOI21_X1 #() 
AOI21_X1_539_ (
  .A({ S5128 }),
  .B1({ S9861 }),
  .B2({ S9800 }),
  .ZN({ S10268 })
);
AOI21_X1 #() 
AOI21_X1_540_ (
  .A({ S9790 }),
  .B1({ S10268 }),
  .B2({ S10101 }),
  .ZN({ S10269 })
);
AOI21_X1 #() 
AOI21_X1_541_ (
  .A({ S25957[534] }),
  .B1({ S10269 }),
  .B2({ S10267 }),
  .ZN({ S10270 })
);
NAND2_X1 #() 
NAND2_X1_864_ (
  .A1({ S10266 }),
  .A2({ S10270 }),
  .ZN({ S10271 })
);
NOR2_X1 #() 
NOR2_X1_198_ (
  .A1({ S9871 }),
  .A2({ S25957[532] }),
  .ZN({ S10272 })
);
NAND3_X1 #() 
NAND3_X1_996_ (
  .A1({ S9829 }),
  .A2({ S25957[531] }),
  .A3({ S9810 }),
  .ZN({ S10274 })
);
AND2_X1 #() 
AND2_X1_54_ (
  .A1({ S9924 }),
  .A2({ S25957[532] }),
  .ZN({ S10275 })
);
AOI22_X1 #() 
AOI22_X1_103_ (
  .A1({ S10274 }),
  .A2({ S10275 }),
  .B1({ S9933 }),
  .B2({ S10272 }),
  .ZN({ S10276 })
);
OAI211_X1 #() 
OAI211_X1_293_ (
  .A({ S9867 }),
  .B({ S5128 }),
  .C1({ S9865 }),
  .C2({ S25957[531] }),
  .ZN({ S10277 })
);
NAND4_X1 #() 
NAND4_X1_119_ (
  .A1({ S10135 }),
  .A2({ S10048 }),
  .A3({ S9822 }),
  .A4({ S25957[532] }),
  .ZN({ S10278 })
);
OAI211_X1 #() 
OAI211_X1_294_ (
  .A({ S10278 }),
  .B({ S9790 }),
  .C1({ S10049 }),
  .C2({ S10277 }),
  .ZN({ S10279 })
);
OAI211_X1 #() 
OAI211_X1_295_ (
  .A({ S25957[534] }),
  .B({ S10279 }),
  .C1({ S10276 }),
  .C2({ S9790 }),
  .ZN({ S10280 })
);
NAND3_X1 #() 
NAND3_X1_997_ (
  .A1({ S10280 }),
  .A2({ S10271 }),
  .A3({ S4924 }),
  .ZN({ S10281 })
);
OAI21_X1 #() 
OAI21_X1_488_ (
  .A({ S25957[532] }),
  .B1({ S10021 }),
  .B2({ S9971 }),
  .ZN({ S10282 })
);
INV_X1 #() 
INV_X1_293_ (
  .A({ S10282 }),
  .ZN({ S10283 })
);
NAND2_X1 #() 
NAND2_X1_865_ (
  .A1({ S10100 }),
  .A2({ S10283 }),
  .ZN({ S10285 })
);
OAI211_X1 #() 
OAI211_X1_296_ (
  .A({ S10103 }),
  .B({ S5128 }),
  .C1({ S10034 }),
  .C2({ S9946 }),
  .ZN({ S10286 })
);
NAND3_X1 #() 
NAND3_X1_998_ (
  .A1({ S10285 }),
  .A2({ S25957[533] }),
  .A3({ S10286 }),
  .ZN({ S10287 })
);
OAI21_X1 #() 
OAI21_X1_489_ (
  .A({ S6 }),
  .B1({ S9800 }),
  .B2({ S25957[530] }),
  .ZN({ S10288 })
);
AOI21_X1 #() 
AOI21_X1_542_ (
  .A({ S25957[532] }),
  .B1({ S10046 }),
  .B2({ S10288 }),
  .ZN({ S10289 })
);
NAND3_X1 #() 
NAND3_X1_999_ (
  .A1({ S9973 }),
  .A2({ S9800 }),
  .A3({ S9801 }),
  .ZN({ S10290 })
);
OAI21_X1 #() 
OAI21_X1_490_ (
  .A({ S10290 }),
  .B1({ S10137 }),
  .B2({ S25957[531] }),
  .ZN({ S10291 })
);
AOI21_X1 #() 
AOI21_X1_543_ (
  .A({ S10289 }),
  .B1({ S25957[532] }),
  .B2({ S10291 }),
  .ZN({ S10292 })
);
OAI211_X1 #() 
OAI211_X1_297_ (
  .A({ S25957[534] }),
  .B({ S10287 }),
  .C1({ S10292 }),
  .C2({ S25957[533] }),
  .ZN({ S10293 })
);
NAND4_X1 #() 
NAND4_X1_120_ (
  .A1({ S9822 }),
  .A2({ S9823 }),
  .A3({ S6 }),
  .A4({ S9865 }),
  .ZN({ S10294 })
);
AOI21_X1 #() 
AOI21_X1_544_ (
  .A({ S25957[532] }),
  .B1({ S10294 }),
  .B2({ S10182 }),
  .ZN({ S10296 })
);
AND3_X1 #() 
AND3_X1_40_ (
  .A1({ S10109 }),
  .A2({ S9974 }),
  .A3({ S25957[532] }),
  .ZN({ S10297 })
);
OAI21_X1 #() 
OAI21_X1_491_ (
  .A({ S9790 }),
  .B1({ S10297 }),
  .B2({ S10296 }),
  .ZN({ S10298 })
);
NAND3_X1 #() 
NAND3_X1_1000_ (
  .A1({ S10133 }),
  .A2({ S10125 }),
  .A3({ S5128 }),
  .ZN({ S10299 })
);
OAI21_X1 #() 
OAI21_X1_492_ (
  .A({ S25957[531] }),
  .B1({ S25957[529] }),
  .B2({ S9797 }),
  .ZN({ S10300 })
);
AOI22_X1 #() 
AOI22_X1_104_ (
  .A1({ S10300 }),
  .A2({ S10175 }),
  .B1({ S9811 }),
  .B2({ S9837 }),
  .ZN({ S10301 })
);
OAI211_X1 #() 
OAI211_X1_298_ (
  .A({ S25957[533] }),
  .B({ S10299 }),
  .C1({ S10301 }),
  .C2({ S5128 }),
  .ZN({ S10302 })
);
NAND3_X1 #() 
NAND3_X1_1001_ (
  .A1({ S10298 }),
  .A2({ S10302 }),
  .A3({ S7708 }),
  .ZN({ S10303 })
);
NAND3_X1 #() 
NAND3_X1_1002_ (
  .A1({ S10293 }),
  .A2({ S25957[535] }),
  .A3({ S10303 }),
  .ZN({ S10304 })
);
NAND3_X1 #() 
NAND3_X1_1003_ (
  .A1({ S10304 }),
  .A2({ S10281 }),
  .A3({ S10257 }),
  .ZN({ S10305 })
);
AND2_X1 #() 
AND2_X1_55_ (
  .A1({ S10266 }),
  .A2({ S10270 }),
  .ZN({ S10307 })
);
NAND2_X1 #() 
NAND2_X1_866_ (
  .A1({ S9933 }),
  .A2({ S10272 }),
  .ZN({ S10308 })
);
OAI211_X1 #() 
OAI211_X1_299_ (
  .A({ S25957[532] }),
  .B({ S9924 }),
  .C1({ S10057 }),
  .C2({ S9958 }),
  .ZN({ S10309 })
);
AOI21_X1 #() 
AOI21_X1_545_ (
  .A({ S9790 }),
  .B1({ S10308 }),
  .B2({ S10309 }),
  .ZN({ S10310 })
);
NAND2_X1 #() 
NAND2_X1_867_ (
  .A1({ S10279 }),
  .A2({ S25957[534] }),
  .ZN({ S10311 })
);
OAI21_X1 #() 
OAI21_X1_493_ (
  .A({ S4924 }),
  .B1({ S10310 }),
  .B2({ S10311 }),
  .ZN({ S10312 })
);
NOR2_X1 #() 
NOR2_X1_199_ (
  .A1({ S10307 }),
  .A2({ S10312 }),
  .ZN({ S10313 })
);
AOI22_X1 #() 
AOI22_X1_105_ (
  .A1({ S10206 }),
  .A2({ S6 }),
  .B1({ S10067 }),
  .B2({ S9973 }),
  .ZN({ S10314 })
);
OAI211_X1 #() 
OAI211_X1_300_ (
  .A({ S10050 }),
  .B({ S9790 }),
  .C1({ S10314 }),
  .C2({ S5128 }),
  .ZN({ S10315 })
);
NAND2_X1 #() 
NAND2_X1_868_ (
  .A1({ S9888 }),
  .A2({ S9890 }),
  .ZN({ S10316 })
);
AOI21_X1 #() 
AOI21_X1_546_ (
  .A({ S10282 }),
  .B1({ S10316 }),
  .B2({ S6 }),
  .ZN({ S10317 })
);
NOR2_X1 #() 
NOR2_X1_200_ (
  .A1({ S10034 }),
  .A2({ S9946 }),
  .ZN({ S10318 })
);
OAI21_X1 #() 
OAI21_X1_494_ (
  .A({ S5128 }),
  .B1({ S9878 }),
  .B2({ S10141 }),
  .ZN({ S10319 })
);
NOR2_X1 #() 
NOR2_X1_201_ (
  .A1({ S10318 }),
  .A2({ S10319 }),
  .ZN({ S10320 })
);
OAI21_X1 #() 
OAI21_X1_495_ (
  .A({ S25957[533] }),
  .B1({ S10320 }),
  .B2({ S10317 }),
  .ZN({ S10321 })
);
NAND3_X1 #() 
NAND3_X1_1004_ (
  .A1({ S10321 }),
  .A2({ S25957[534] }),
  .A3({ S10315 }),
  .ZN({ S10322 })
);
NAND2_X1 #() 
NAND2_X1_869_ (
  .A1({ S10294 }),
  .A2({ S10182 }),
  .ZN({ S10323 })
);
NAND2_X1 #() 
NAND2_X1_870_ (
  .A1({ S10323 }),
  .A2({ S5128 }),
  .ZN({ S10324 })
);
NAND3_X1 #() 
NAND3_X1_1005_ (
  .A1({ S10109 }),
  .A2({ S9974 }),
  .A3({ S25957[532] }),
  .ZN({ S10325 })
);
AOI21_X1 #() 
AOI21_X1_547_ (
  .A({ S25957[533] }),
  .B1({ S10324 }),
  .B2({ S10325 }),
  .ZN({ S10326 })
);
NAND3_X1 #() 
NAND3_X1_1006_ (
  .A1({ S9841 }),
  .A2({ S6 }),
  .A3({ S9837 }),
  .ZN({ S10328 })
);
NAND2_X1 #() 
NAND2_X1_871_ (
  .A1({ S10300 }),
  .A2({ S10175 }),
  .ZN({ S10329 })
);
NAND3_X1 #() 
NAND3_X1_1007_ (
  .A1({ S10329 }),
  .A2({ S25957[532] }),
  .A3({ S10328 }),
  .ZN({ S10330 })
);
NAND2_X1 #() 
NAND2_X1_872_ (
  .A1({ S10133 }),
  .A2({ S10125 }),
  .ZN({ S10331 })
);
NAND2_X1 #() 
NAND2_X1_873_ (
  .A1({ S10331 }),
  .A2({ S5128 }),
  .ZN({ S10332 })
);
AOI21_X1 #() 
AOI21_X1_548_ (
  .A({ S9790 }),
  .B1({ S10332 }),
  .B2({ S10330 }),
  .ZN({ S10333 })
);
OAI21_X1 #() 
OAI21_X1_496_ (
  .A({ S7708 }),
  .B1({ S10333 }),
  .B2({ S10326 }),
  .ZN({ S10334 })
);
AOI21_X1 #() 
AOI21_X1_549_ (
  .A({ S4924 }),
  .B1({ S10334 }),
  .B2({ S10322 }),
  .ZN({ S10335 })
);
OAI21_X1 #() 
OAI21_X1_497_ (
  .A({ S25957[728] }),
  .B1({ S10335 }),
  .B2({ S10313 }),
  .ZN({ S10336 })
);
AOI21_X1 #() 
AOI21_X1_550_ (
  .A({ S10256 }),
  .B1({ S10336 }),
  .B2({ S10305 }),
  .ZN({ S10337 })
);
INV_X1 #() 
INV_X1_294_ (
  .A({ S10256 }),
  .ZN({ S25957[568] })
);
AND3_X1 #() 
AND3_X1_41_ (
  .A1({ S10304 }),
  .A2({ S10281 }),
  .A3({ S10257 }),
  .ZN({ S10339 })
);
AOI21_X1 #() 
AOI21_X1_551_ (
  .A({ S10257 }),
  .B1({ S10304 }),
  .B2({ S10281 }),
  .ZN({ S10340 })
);
NOR3_X1 #() 
NOR3_X1_28_ (
  .A1({ S10339 }),
  .A2({ S10340 }),
  .A3({ S25957[568] }),
  .ZN({ S10341 })
);
OAI21_X1 #() 
OAI21_X1_498_ (
  .A({ S25957[536] }),
  .B1({ S10341 }),
  .B2({ S10337 }),
  .ZN({ S10342 })
);
OAI21_X1 #() 
OAI21_X1_499_ (
  .A({ S25957[568] }),
  .B1({ S10339 }),
  .B2({ S10340 }),
  .ZN({ S10343 })
);
NAND3_X1 #() 
NAND3_X1_1008_ (
  .A1({ S10336 }),
  .A2({ S10256 }),
  .A3({ S10305 }),
  .ZN({ S10344 })
);
NAND3_X1 #() 
NAND3_X1_1009_ (
  .A1({ S10343 }),
  .A2({ S10344 }),
  .A3({ S7386 }),
  .ZN({ S10345 })
);
NAND2_X1 #() 
NAND2_X1_874_ (
  .A1({ S10342 }),
  .A2({ S10345 }),
  .ZN({ S25957[408] })
);
NOR2_X1 #() 
NOR2_X1_202_ (
  .A1({ S9043 }),
  .A2({ S9044 }),
  .ZN({ S25957[569] })
);
AOI21_X1 #() 
AOI21_X1_552_ (
  .A({ S25957[531] }),
  .B1({ S9965 }),
  .B2({ S9980 }),
  .ZN({ S10347 })
);
NOR3_X1 #() 
NOR3_X1_29_ (
  .A1({ S9828 }),
  .A2({ S10347 }),
  .A3({ S25957[532] }),
  .ZN({ S10348 })
);
INV_X1 #() 
INV_X1_295_ (
  .A({ S9807 }),
  .ZN({ S10349 })
);
NAND2_X1 #() 
NAND2_X1_875_ (
  .A1({ S10349 }),
  .A2({ S25957[531] }),
  .ZN({ S10350 })
);
NAND3_X1 #() 
NAND3_X1_1010_ (
  .A1({ S10135 }),
  .A2({ S6 }),
  .A3({ S9822 }),
  .ZN({ S10351 })
);
NAND3_X1 #() 
NAND3_X1_1011_ (
  .A1({ S10351 }),
  .A2({ S10350 }),
  .A3({ S25957[532] }),
  .ZN({ S10352 })
);
NAND2_X1 #() 
NAND2_X1_876_ (
  .A1({ S10352 }),
  .A2({ S9790 }),
  .ZN({ S10353 })
);
AOI21_X1 #() 
AOI21_X1_553_ (
  .A({ S6 }),
  .B1({ S9829 }),
  .B2({ S9823 }),
  .ZN({ S10354 })
);
NAND3_X1 #() 
NAND3_X1_1012_ (
  .A1({ S9801 }),
  .A2({ S6 }),
  .A3({ S9807 }),
  .ZN({ S10355 })
);
OAI211_X1 #() 
OAI211_X1_301_ (
  .A({ S10355 }),
  .B({ S5128 }),
  .C1({ S9932 }),
  .C2({ S6 }),
  .ZN({ S10356 })
);
OAI211_X1 #() 
OAI211_X1_302_ (
  .A({ S10356 }),
  .B({ S25957[533] }),
  .C1({ S10354 }),
  .C2({ S9834 }),
  .ZN({ S10358 })
);
OAI211_X1 #() 
OAI211_X1_303_ (
  .A({ S10358 }),
  .B({ S7708 }),
  .C1({ S10348 }),
  .C2({ S10353 }),
  .ZN({ S10359 })
);
OAI211_X1 #() 
OAI211_X1_304_ (
  .A({ S25957[532] }),
  .B({ S10328 }),
  .C1({ S10057 }),
  .C2({ S10059 }),
  .ZN({ S10360 })
);
NAND3_X1 #() 
NAND3_X1_1013_ (
  .A1({ S9789 }),
  .A2({ S25957[531] }),
  .A3({ S9797 }),
  .ZN({ S10361 })
);
AOI21_X1 #() 
AOI21_X1_554_ (
  .A({ S25957[532] }),
  .B1({ S10027 }),
  .B2({ S6 }),
  .ZN({ S10362 })
);
NAND3_X1 #() 
NAND3_X1_1014_ (
  .A1({ S10362 }),
  .A2({ S10109 }),
  .A3({ S10361 }),
  .ZN({ S10363 })
);
NAND3_X1 #() 
NAND3_X1_1015_ (
  .A1({ S10360 }),
  .A2({ S9790 }),
  .A3({ S10363 }),
  .ZN({ S10364 })
);
NAND2_X1 #() 
NAND2_X1_877_ (
  .A1({ S9965 }),
  .A2({ S6 }),
  .ZN({ S10365 })
);
OAI211_X1 #() 
OAI211_X1_305_ (
  .A({ S10365 }),
  .B({ S5128 }),
  .C1({ S10057 }),
  .C2({ S9958 }),
  .ZN({ S10366 })
);
NAND3_X1 #() 
NAND3_X1_1016_ (
  .A1({ S10015 }),
  .A2({ S9845 }),
  .A3({ S25957[532] }),
  .ZN({ S10367 })
);
NAND3_X1 #() 
NAND3_X1_1017_ (
  .A1({ S10366 }),
  .A2({ S10367 }),
  .A3({ S25957[533] }),
  .ZN({ S10369 })
);
NAND3_X1 #() 
NAND3_X1_1018_ (
  .A1({ S10369 }),
  .A2({ S10364 }),
  .A3({ S25957[534] }),
  .ZN({ S10370 })
);
NAND3_X1 #() 
NAND3_X1_1019_ (
  .A1({ S10359 }),
  .A2({ S25957[535] }),
  .A3({ S10370 }),
  .ZN({ S10371 })
);
NAND2_X1 #() 
NAND2_X1_878_ (
  .A1({ S10067 }),
  .A2({ S9815 }),
  .ZN({ S10372 })
);
NAND3_X1 #() 
NAND3_X1_1020_ (
  .A1({ S9838 }),
  .A2({ S6 }),
  .A3({ S9854 }),
  .ZN({ S10373 })
);
NAND3_X1 #() 
NAND3_X1_1021_ (
  .A1({ S10372 }),
  .A2({ S10373 }),
  .A3({ S25957[532] }),
  .ZN({ S10374 })
);
OAI21_X1 #() 
OAI21_X1_500_ (
  .A({ S9854 }),
  .B1({ S9852 }),
  .B2({ S25957[528] }),
  .ZN({ S10375 })
);
AOI21_X1 #() 
AOI21_X1_555_ (
  .A({ S9790 }),
  .B1({ S10031 }),
  .B2({ S10375 }),
  .ZN({ S10376 })
);
NAND2_X1 #() 
NAND2_X1_879_ (
  .A1({ S10376 }),
  .A2({ S10374 }),
  .ZN({ S10377 })
);
NAND3_X1 #() 
NAND3_X1_1022_ (
  .A1({ S9890 }),
  .A2({ S9978 }),
  .A3({ S6 }),
  .ZN({ S10378 })
);
AND3_X1 #() 
AND3_X1_42_ (
  .A1({ S10274 }),
  .A2({ S25957[532] }),
  .A3({ S10378 }),
  .ZN({ S10380 })
);
NAND2_X1 #() 
NAND2_X1_880_ (
  .A1({ S9804 }),
  .A2({ S9861 }),
  .ZN({ S10381 })
);
NAND3_X1 #() 
NAND3_X1_1023_ (
  .A1({ S10381 }),
  .A2({ S10290 }),
  .A3({ S5128 }),
  .ZN({ S10382 })
);
NAND2_X1 #() 
NAND2_X1_881_ (
  .A1({ S10382 }),
  .A2({ S9790 }),
  .ZN({ S10383 })
);
OAI211_X1 #() 
OAI211_X1_306_ (
  .A({ S10377 }),
  .B({ S25957[534] }),
  .C1({ S10380 }),
  .C2({ S10383 }),
  .ZN({ S10384 })
);
NAND3_X1 #() 
NAND3_X1_1024_ (
  .A1({ S9868 }),
  .A2({ S25957[532] }),
  .A3({ S10121 }),
  .ZN({ S10385 })
);
AOI21_X1 #() 
AOI21_X1_556_ (
  .A({ S25957[532] }),
  .B1({ S9852 }),
  .B2({ S25957[531] }),
  .ZN({ S10386 })
);
NAND2_X1 #() 
NAND2_X1_882_ (
  .A1({ S10386 }),
  .A2({ S10221 }),
  .ZN({ S10387 })
);
NAND3_X1 #() 
NAND3_X1_1025_ (
  .A1({ S10385 }),
  .A2({ S10387 }),
  .A3({ S9790 }),
  .ZN({ S10388 })
);
NAND4_X1 #() 
NAND4_X1_121_ (
  .A1({ S9854 }),
  .A2({ S25957[529] }),
  .A3({ S9797 }),
  .A4({ S25957[531] }),
  .ZN({ S10389 })
);
AOI21_X1 #() 
AOI21_X1_557_ (
  .A({ S5128 }),
  .B1({ S10389 }),
  .B2({ S10127 }),
  .ZN({ S10391 })
);
OAI21_X1 #() 
OAI21_X1_501_ (
  .A({ S25957[533] }),
  .B1({ S9826 }),
  .B2({ S10391 }),
  .ZN({ S10392 })
);
NAND3_X1 #() 
NAND3_X1_1026_ (
  .A1({ S10392 }),
  .A2({ S7708 }),
  .A3({ S10388 }),
  .ZN({ S10393 })
);
NAND3_X1 #() 
NAND3_X1_1027_ (
  .A1({ S10384 }),
  .A2({ S10393 }),
  .A3({ S4924 }),
  .ZN({ S10394 })
);
AOI21_X1 #() 
AOI21_X1_558_ (
  .A({ S25957[729] }),
  .B1({ S10371 }),
  .B2({ S10394 }),
  .ZN({ S10395 })
);
AND3_X1 #() 
AND3_X1_43_ (
  .A1({ S10371 }),
  .A2({ S10394 }),
  .A3({ S25957[729] }),
  .ZN({ S10396 })
);
OAI21_X1 #() 
OAI21_X1_502_ (
  .A({ S25957[569] }),
  .B1({ S10396 }),
  .B2({ S10395 }),
  .ZN({ S10397 })
);
INV_X1 #() 
INV_X1_296_ (
  .A({ S25957[569] }),
  .ZN({ S10398 })
);
NAND2_X1 #() 
NAND2_X1_883_ (
  .A1({ S10371 }),
  .A2({ S10394 }),
  .ZN({ S10399 })
);
NAND2_X1 #() 
NAND2_X1_884_ (
  .A1({ S10399 }),
  .A2({ S7460 }),
  .ZN({ S10400 })
);
NAND3_X1 #() 
NAND3_X1_1028_ (
  .A1({ S10371 }),
  .A2({ S10394 }),
  .A3({ S25957[729] }),
  .ZN({ S10401 })
);
NAND3_X1 #() 
NAND3_X1_1029_ (
  .A1({ S10400 }),
  .A2({ S10398 }),
  .A3({ S10401 }),
  .ZN({ S10402 })
);
NAND3_X1 #() 
NAND3_X1_1030_ (
  .A1({ S10397 }),
  .A2({ S10402 }),
  .A3({ S25957[537] }),
  .ZN({ S10403 })
);
NAND3_X1 #() 
NAND3_X1_1031_ (
  .A1({ S10400 }),
  .A2({ S25957[569] }),
  .A3({ S10401 }),
  .ZN({ S10404 })
);
OAI21_X1 #() 
OAI21_X1_503_ (
  .A({ S10398 }),
  .B1({ S10396 }),
  .B2({ S10395 }),
  .ZN({ S10405 })
);
NAND3_X1 #() 
NAND3_X1_1032_ (
  .A1({ S10405 }),
  .A2({ S10404 }),
  .A3({ S9169 }),
  .ZN({ S10406 })
);
NAND2_X1 #() 
NAND2_X1_885_ (
  .A1({ S10403 }),
  .A2({ S10406 }),
  .ZN({ S25957[409] })
);
NAND2_X1 #() 
NAND2_X1_886_ (
  .A1({ S2223 }),
  .A2({ S2226 }),
  .ZN({ S25957[826] })
);
XNOR2_X1 #() 
XNOR2_X1_30_ (
  .A({ S7469 }),
  .B({ S25957[826] }),
  .ZN({ S25957[698] })
);
NAND2_X1 #() 
NAND2_X1_887_ (
  .A1({ S7550 }),
  .A2({ S7554 }),
  .ZN({ S25957[602] })
);
AND2_X1 #() 
AND2_X1_56_ (
  .A1({ S25957[602] }),
  .A2({ S25957[698] }),
  .ZN({ S10408 })
);
NOR2_X1 #() 
NOR2_X1_203_ (
  .A1({ S25957[602] }),
  .A2({ S25957[698] }),
  .ZN({ S10409 })
);
NOR2_X1 #() 
NOR2_X1_204_ (
  .A1({ S10408 }),
  .A2({ S10409 }),
  .ZN({ S25957[570] })
);
NAND2_X1 #() 
NAND2_X1_888_ (
  .A1({ S9912 }),
  .A2({ S25957[531] }),
  .ZN({ S10410 })
);
OAI211_X1 #() 
OAI211_X1_307_ (
  .A({ S10410 }),
  .B({ S5128 }),
  .C1({ S25957[531] }),
  .C2({ S10206 }),
  .ZN({ S10411 })
);
NAND2_X1 #() 
NAND2_X1_889_ (
  .A1({ S9875 }),
  .A2({ S25957[530] }),
  .ZN({ S10412 })
);
AOI22_X1 #() 
AOI22_X1_106_ (
  .A1({ S10412 }),
  .A2({ S9794 }),
  .B1({ S9815 }),
  .B2({ S10135 }),
  .ZN({ S10413 })
);
OAI211_X1 #() 
OAI211_X1_308_ (
  .A({ S10411 }),
  .B({ S9790 }),
  .C1({ S10413 }),
  .C2({ S5128 }),
  .ZN({ S10414 })
);
OAI21_X1 #() 
OAI21_X1_504_ (
  .A({ S5128 }),
  .B1({ S10349 }),
  .B2({ S9817 }),
  .ZN({ S10415 })
);
NAND3_X1 #() 
NAND3_X1_1033_ (
  .A1({ S9801 }),
  .A2({ S9813 }),
  .A3({ S25957[531] }),
  .ZN({ S10416 })
);
AOI21_X1 #() 
AOI21_X1_559_ (
  .A({ S5128 }),
  .B1({ S10416 }),
  .B2({ S10175 }),
  .ZN({ S10418 })
);
INV_X1 #() 
INV_X1_297_ (
  .A({ S10418 }),
  .ZN({ S10419 })
);
OAI211_X1 #() 
OAI211_X1_309_ (
  .A({ S10419 }),
  .B({ S25957[533] }),
  .C1({ S9859 }),
  .C2({ S10415 }),
  .ZN({ S10420 })
);
NAND3_X1 #() 
NAND3_X1_1034_ (
  .A1({ S10420 }),
  .A2({ S10414 }),
  .A3({ S25957[534] }),
  .ZN({ S10421 })
);
OAI21_X1 #() 
OAI21_X1_505_ (
  .A({ S10410 }),
  .B1({ S10034 }),
  .B2({ S9798 }),
  .ZN({ S10422 })
);
NAND2_X1 #() 
NAND2_X1_890_ (
  .A1({ S10422 }),
  .A2({ S25957[532] }),
  .ZN({ S10423 })
);
AOI21_X1 #() 
AOI21_X1_560_ (
  .A({ S6 }),
  .B1({ S9965 }),
  .B2({ S9980 }),
  .ZN({ S10424 })
);
AOI21_X1 #() 
AOI21_X1_561_ (
  .A({ S25957[531] }),
  .B1({ S9855 }),
  .B2({ S9835 }),
  .ZN({ S10425 })
);
OAI21_X1 #() 
OAI21_X1_506_ (
  .A({ S5128 }),
  .B1({ S10424 }),
  .B2({ S10425 }),
  .ZN({ S10426 })
);
NAND3_X1 #() 
NAND3_X1_1035_ (
  .A1({ S10426 }),
  .A2({ S10423 }),
  .A3({ S9790 }),
  .ZN({ S10427 })
);
NAND2_X1 #() 
NAND2_X1_891_ (
  .A1({ S9890 }),
  .A2({ S9815 }),
  .ZN({ S10428 })
);
NAND2_X1 #() 
NAND2_X1_892_ (
  .A1({ S10193 }),
  .A2({ S10428 }),
  .ZN({ S10429 })
);
NAND2_X1 #() 
NAND2_X1_893_ (
  .A1({ S10429 }),
  .A2({ S25957[532] }),
  .ZN({ S10430 })
);
OAI21_X1 #() 
OAI21_X1_507_ (
  .A({ S9975 }),
  .B1({ S9958 }),
  .B2({ S10071 }),
  .ZN({ S10431 })
);
AOI21_X1 #() 
AOI21_X1_562_ (
  .A({ S9790 }),
  .B1({ S10431 }),
  .B2({ S5128 }),
  .ZN({ S10432 })
);
NAND2_X1 #() 
NAND2_X1_894_ (
  .A1({ S10430 }),
  .A2({ S10432 }),
  .ZN({ S10433 })
);
NAND3_X1 #() 
NAND3_X1_1036_ (
  .A1({ S10433 }),
  .A2({ S10427 }),
  .A3({ S7708 }),
  .ZN({ S10434 })
);
NAND3_X1 #() 
NAND3_X1_1037_ (
  .A1({ S10434 }),
  .A2({ S10421 }),
  .A3({ S4924 }),
  .ZN({ S10435 })
);
NOR2_X1 #() 
NOR2_X1_205_ (
  .A1({ S10263 }),
  .A2({ S25957[532] }),
  .ZN({ S10436 })
);
NAND4_X1 #() 
NAND4_X1_122_ (
  .A1({ S9945 }),
  .A2({ S9842 }),
  .A3({ S9800 }),
  .A4({ S9841 }),
  .ZN({ S10437 })
);
AOI21_X1 #() 
AOI21_X1_563_ (
  .A({ S5128 }),
  .B1({ S9946 }),
  .B2({ S6 }),
  .ZN({ S10439 })
);
AOI22_X1 #() 
AOI22_X1_107_ (
  .A1({ S10436 }),
  .A2({ S9808 }),
  .B1({ S10437 }),
  .B2({ S10439 }),
  .ZN({ S10440 })
);
OAI211_X1 #() 
OAI211_X1_310_ (
  .A({ S9821 }),
  .B({ S25957[532] }),
  .C1({ S10034 }),
  .C2({ S9946 }),
  .ZN({ S10441 })
);
NOR2_X1 #() 
NOR2_X1_206_ (
  .A1({ S9811 }),
  .A2({ S25957[532] }),
  .ZN({ S10442 })
);
AOI21_X1 #() 
AOI21_X1_564_ (
  .A({ S6 }),
  .B1({ S9800 }),
  .B2({ S25957[530] }),
  .ZN({ S10443 })
);
NAND2_X1 #() 
NAND2_X1_895_ (
  .A1({ S10188 }),
  .A2({ S10443 }),
  .ZN({ S10444 })
);
AOI21_X1 #() 
AOI21_X1_565_ (
  .A({ S9790 }),
  .B1({ S10444 }),
  .B2({ S10442 }),
  .ZN({ S10445 })
);
AOI22_X1 #() 
AOI22_X1_108_ (
  .A1({ S10440 }),
  .A2({ S9790 }),
  .B1({ S10445 }),
  .B2({ S10441 }),
  .ZN({ S10446 })
);
INV_X1 #() 
INV_X1_298_ (
  .A({ S10168 }),
  .ZN({ S10447 })
);
AOI21_X1 #() 
AOI21_X1_566_ (
  .A({ S8137 }),
  .B1({ S10048 }),
  .B2({ S9971 }),
  .ZN({ S10448 })
);
OAI21_X1 #() 
OAI21_X1_508_ (
  .A({ S25957[532] }),
  .B1({ S10447 }),
  .B2({ S10448 }),
  .ZN({ S10450 })
);
NAND2_X1 #() 
NAND2_X1_896_ (
  .A1({ S9976 }),
  .A2({ S5128 }),
  .ZN({ S10451 })
);
NAND3_X1 #() 
NAND3_X1_1038_ (
  .A1({ S10451 }),
  .A2({ S10450 }),
  .A3({ S9790 }),
  .ZN({ S10452 })
);
AOI21_X1 #() 
AOI21_X1_567_ (
  .A({ S9837 }),
  .B1({ S8137 }),
  .B2({ S8281 }),
  .ZN({ S10453 })
);
AOI22_X1 #() 
AOI22_X1_109_ (
  .A1({ S9914 }),
  .A2({ S9968 }),
  .B1({ S10453 }),
  .B2({ S25957[531] }),
  .ZN({ S10454 })
);
OAI211_X1 #() 
OAI211_X1_311_ (
  .A({ S9949 }),
  .B({ S5128 }),
  .C1({ S10067 }),
  .C2({ S10197 }),
  .ZN({ S10455 })
);
OAI211_X1 #() 
OAI211_X1_312_ (
  .A({ S10455 }),
  .B({ S25957[533] }),
  .C1({ S5128 }),
  .C2({ S10454 }),
  .ZN({ S10456 })
);
NAND3_X1 #() 
NAND3_X1_1039_ (
  .A1({ S10456 }),
  .A2({ S10452 }),
  .A3({ S7708 }),
  .ZN({ S10457 })
);
OAI211_X1 #() 
OAI211_X1_313_ (
  .A({ S10457 }),
  .B({ S25957[535] }),
  .C1({ S10446 }),
  .C2({ S7708 }),
  .ZN({ S10458 })
);
AOI21_X1 #() 
AOI21_X1_568_ (
  .A({ S7469 }),
  .B1({ S10435 }),
  .B2({ S10458 }),
  .ZN({ S10459 })
);
NAND3_X1 #() 
NAND3_X1_1040_ (
  .A1({ S10188 }),
  .A2({ S6 }),
  .A3({ S9841 }),
  .ZN({ S10461 })
);
NAND3_X1 #() 
NAND3_X1_1041_ (
  .A1({ S10461 }),
  .A2({ S9933 }),
  .A3({ S5128 }),
  .ZN({ S10462 })
);
OAI211_X1 #() 
OAI211_X1_314_ (
  .A({ S10410 }),
  .B({ S25957[532] }),
  .C1({ S10034 }),
  .C2({ S9798 }),
  .ZN({ S10463 })
);
NAND3_X1 #() 
NAND3_X1_1042_ (
  .A1({ S10462 }),
  .A2({ S9790 }),
  .A3({ S10463 }),
  .ZN({ S10464 })
);
OAI211_X1 #() 
OAI211_X1_315_ (
  .A({ S9975 }),
  .B({ S5128 }),
  .C1({ S9958 }),
  .C2({ S10071 }),
  .ZN({ S10465 })
);
NAND3_X1 #() 
NAND3_X1_1043_ (
  .A1({ S10193 }),
  .A2({ S25957[532] }),
  .A3({ S10428 }),
  .ZN({ S10466 })
);
NAND3_X1 #() 
NAND3_X1_1044_ (
  .A1({ S10466 }),
  .A2({ S25957[533] }),
  .A3({ S10465 }),
  .ZN({ S10467 })
);
NAND3_X1 #() 
NAND3_X1_1045_ (
  .A1({ S10464 }),
  .A2({ S10467 }),
  .A3({ S7708 }),
  .ZN({ S10468 })
);
OAI21_X1 #() 
OAI21_X1_509_ (
  .A({ S25957[531] }),
  .B1({ S10035 }),
  .B2({ S9954 }),
  .ZN({ S10469 })
);
INV_X1 #() 
INV_X1_299_ (
  .A({ S10415 }),
  .ZN({ S10470 })
);
AOI21_X1 #() 
AOI21_X1_569_ (
  .A({ S10418 }),
  .B1({ S10469 }),
  .B2({ S10470 }),
  .ZN({ S10472 })
);
NAND2_X1 #() 
NAND2_X1_897_ (
  .A1({ S10074 }),
  .A2({ S25957[531] }),
  .ZN({ S10473 })
);
OAI211_X1 #() 
OAI211_X1_316_ (
  .A({ S10473 }),
  .B({ S5128 }),
  .C1({ S10137 }),
  .C2({ S25957[531] }),
  .ZN({ S10474 })
);
NOR2_X1 #() 
NOR2_X1_207_ (
  .A1({ S9801 }),
  .A2({ S8281 }),
  .ZN({ S10475 })
);
NAND2_X1 #() 
NAND2_X1_898_ (
  .A1({ S9815 }),
  .A2({ S10135 }),
  .ZN({ S10476 })
);
OAI211_X1 #() 
OAI211_X1_317_ (
  .A({ S10476 }),
  .B({ S25957[532] }),
  .C1({ S10034 }),
  .C2({ S10475 }),
  .ZN({ S10477 })
);
NAND3_X1 #() 
NAND3_X1_1046_ (
  .A1({ S10477 }),
  .A2({ S10474 }),
  .A3({ S9790 }),
  .ZN({ S10478 })
);
OAI211_X1 #() 
OAI211_X1_318_ (
  .A({ S10478 }),
  .B({ S25957[534] }),
  .C1({ S10472 }),
  .C2({ S9790 }),
  .ZN({ S10479 })
);
NAND3_X1 #() 
NAND3_X1_1047_ (
  .A1({ S10479 }),
  .A2({ S10468 }),
  .A3({ S4924 }),
  .ZN({ S10480 })
);
OAI211_X1 #() 
OAI211_X1_319_ (
  .A({ S25957[531] }),
  .B({ S9800 }),
  .C1({ S9801 }),
  .C2({ S8281 }),
  .ZN({ S10481 })
);
OAI211_X1 #() 
OAI211_X1_320_ (
  .A({ S10481 }),
  .B({ S5128 }),
  .C1({ S25957[531] }),
  .C2({ S9948 }),
  .ZN({ S10483 })
);
NAND2_X1 #() 
NAND2_X1_899_ (
  .A1({ S10453 }),
  .A2({ S25957[531] }),
  .ZN({ S10484 })
);
NAND3_X1 #() 
NAND3_X1_1048_ (
  .A1({ S10484 }),
  .A2({ S25957[532] }),
  .A3({ S10221 }),
  .ZN({ S10485 })
);
NAND3_X1 #() 
NAND3_X1_1049_ (
  .A1({ S10483 }),
  .A2({ S25957[533] }),
  .A3({ S10485 }),
  .ZN({ S10486 })
);
NAND3_X1 #() 
NAND3_X1_1050_ (
  .A1({ S10410 }),
  .A2({ S25957[532] }),
  .A3({ S10168 }),
  .ZN({ S10487 })
);
OAI211_X1 #() 
OAI211_X1_321_ (
  .A({ S10487 }),
  .B({ S9790 }),
  .C1({ S25957[532] }),
  .C2({ S9976 }),
  .ZN({ S10488 })
);
NAND3_X1 #() 
NAND3_X1_1051_ (
  .A1({ S10486 }),
  .A2({ S10488 }),
  .A3({ S7708 }),
  .ZN({ S10489 })
);
NAND2_X1 #() 
NAND2_X1_900_ (
  .A1({ S10436 }),
  .A2({ S9808 }),
  .ZN({ S10490 })
);
NAND2_X1 #() 
NAND2_X1_901_ (
  .A1({ S10437 }),
  .A2({ S10439 }),
  .ZN({ S10491 })
);
NAND3_X1 #() 
NAND3_X1_1052_ (
  .A1({ S10490 }),
  .A2({ S10491 }),
  .A3({ S9790 }),
  .ZN({ S10492 })
);
NAND2_X1 #() 
NAND2_X1_902_ (
  .A1({ S10445 }),
  .A2({ S10441 }),
  .ZN({ S10494 })
);
NAND3_X1 #() 
NAND3_X1_1053_ (
  .A1({ S10494 }),
  .A2({ S10492 }),
  .A3({ S25957[534] }),
  .ZN({ S10495 })
);
NAND3_X1 #() 
NAND3_X1_1054_ (
  .A1({ S10495 }),
  .A2({ S10489 }),
  .A3({ S25957[535] }),
  .ZN({ S10496 })
);
AOI21_X1 #() 
AOI21_X1_570_ (
  .A({ S25957[730] }),
  .B1({ S10480 }),
  .B2({ S10496 }),
  .ZN({ S10497 })
);
OAI21_X1 #() 
OAI21_X1_510_ (
  .A({ S25957[570] }),
  .B1({ S10459 }),
  .B2({ S10497 }),
  .ZN({ S10498 })
);
INV_X1 #() 
INV_X1_300_ (
  .A({ S25957[570] }),
  .ZN({ S10499 })
);
NAND3_X1 #() 
NAND3_X1_1055_ (
  .A1({ S10480 }),
  .A2({ S25957[730] }),
  .A3({ S10496 }),
  .ZN({ S10500 })
);
NAND3_X1 #() 
NAND3_X1_1056_ (
  .A1({ S10435 }),
  .A2({ S10458 }),
  .A3({ S7469 }),
  .ZN({ S10501 })
);
NAND3_X1 #() 
NAND3_X1_1057_ (
  .A1({ S10501 }),
  .A2({ S10500 }),
  .A3({ S10499 }),
  .ZN({ S10502 })
);
NAND3_X1 #() 
NAND3_X1_1058_ (
  .A1({ S10498 }),
  .A2({ S25957[538] }),
  .A3({ S10502 }),
  .ZN({ S10503 })
);
OAI21_X1 #() 
OAI21_X1_511_ (
  .A({ S10499 }),
  .B1({ S10459 }),
  .B2({ S10497 }),
  .ZN({ S10505 })
);
NAND3_X1 #() 
NAND3_X1_1059_ (
  .A1({ S10501 }),
  .A2({ S10500 }),
  .A3({ S25957[570] }),
  .ZN({ S10506 })
);
NAND3_X1 #() 
NAND3_X1_1060_ (
  .A1({ S10505 }),
  .A2({ S9051 }),
  .A3({ S10506 }),
  .ZN({ S10507 })
);
NAND2_X1 #() 
NAND2_X1_903_ (
  .A1({ S10503 }),
  .A2({ S10507 }),
  .ZN({ S25957[410] })
);
NAND3_X1 #() 
NAND3_X1_1061_ (
  .A1({ S8834 }),
  .A2({ S7576 }),
  .A3({ S8838 }),
  .ZN({ S10508 })
);
NAND3_X1 #() 
NAND3_X1_1062_ (
  .A1({ S8840 }),
  .A2({ S25957[520] }),
  .A3({ S8841 }),
  .ZN({ S10509 })
);
AND4_X1 #() 
AND4_X1_3_ (
  .A1({ S10509 }),
  .A2({ S10508 }),
  .A3({ S8938 }),
  .A4({ S8942 }),
  .ZN({ S30 })
);
AOI21_X1 #() 
AOI21_X1_571_ (
  .A({ S4806 }),
  .B1({ S8939 }),
  .B2({ S8940 }),
  .ZN({ S10510 })
);
AOI21_X1 #() 
AOI21_X1_572_ (
  .A({ S25957[649] }),
  .B1({ S8933 }),
  .B2({ S8937 }),
  .ZN({ S10511 })
);
OAI211_X1 #() 
OAI211_X1_322_ (
  .A({ S8839 }),
  .B({ S8842 }),
  .C1({ S10511 }),
  .C2({ S10510 }),
  .ZN({ S31 })
);
NAND2_X1 #() 
NAND2_X1_904_ (
  .A1({ S7701 }),
  .A2({ S7698 }),
  .ZN({ S25957[439] })
);
NAND4_X1 #() 
NAND4_X1_123_ (
  .A1({ S10508 }),
  .A2({ S10509 }),
  .A3({ S9037 }),
  .A4({ S9040 }),
  .ZN({ S10513 })
);
INV_X1 #() 
INV_X1_301_ (
  .A({ S10513 }),
  .ZN({ S10514 })
);
OAI21_X1 #() 
OAI21_X1_512_ (
  .A({ S25957[393] }),
  .B1({ S8765 }),
  .B2({ S8764 }),
  .ZN({ S10515 })
);
NAND2_X1 #() 
NAND2_X1_905_ (
  .A1({ S8938 }),
  .A2({ S8942 }),
  .ZN({ S10516 })
);
NAND3_X1 #() 
NAND3_X1_1063_ (
  .A1({ S8759 }),
  .A2({ S8762 }),
  .A3({ S10516 }),
  .ZN({ S10517 })
);
INV_X1 #() 
INV_X1_302_ (
  .A({ S10517 }),
  .ZN({ S10518 })
);
NOR2_X1 #() 
NOR2_X1_208_ (
  .A1({ S21 }),
  .A2({ S10513 }),
  .ZN({ S10519 })
);
NOR2_X1 #() 
NOR2_X1_209_ (
  .A1({ S10519 }),
  .A2({ S10518 }),
  .ZN({ S10520 })
);
OAI211_X1 #() 
OAI211_X1_323_ (
  .A({ S10520 }),
  .B({ S25957[396] }),
  .C1({ S10514 }),
  .C2({ S10515 }),
  .ZN({ S10521 })
);
NAND2_X1 #() 
NAND2_X1_906_ (
  .A1({ S8681 }),
  .A2({ S8683 }),
  .ZN({ S10523 })
);
NAND2_X1 #() 
NAND2_X1_907_ (
  .A1({ S10523 }),
  .A2({ S7575 }),
  .ZN({ S10524 })
);
NAND3_X1 #() 
NAND3_X1_1064_ (
  .A1({ S8681 }),
  .A2({ S8683 }),
  .A3({ S25957[524] }),
  .ZN({ S10525 })
);
NAND2_X1 #() 
NAND2_X1_908_ (
  .A1({ S10524 }),
  .A2({ S10525 }),
  .ZN({ S10526 })
);
NAND4_X1 #() 
NAND4_X1_124_ (
  .A1({ S10508 }),
  .A2({ S10509 }),
  .A3({ S8938 }),
  .A4({ S8942 }),
  .ZN({ S10527 })
);
NAND2_X1 #() 
NAND2_X1_909_ (
  .A1({ S10508 }),
  .A2({ S10509 }),
  .ZN({ S10528 })
);
NAND2_X1 #() 
NAND2_X1_910_ (
  .A1({ S9037 }),
  .A2({ S9040 }),
  .ZN({ S10529 })
);
NAND3_X1 #() 
NAND3_X1_1065_ (
  .A1({ S10528 }),
  .A2({ S10529 }),
  .A3({ S10516 }),
  .ZN({ S10530 })
);
NAND2_X1 #() 
NAND2_X1_911_ (
  .A1({ S10530 }),
  .A2({ S21 }),
  .ZN({ S10531 })
);
OAI211_X1 #() 
OAI211_X1_324_ (
  .A({ S10531 }),
  .B({ S10526 }),
  .C1({ S21 }),
  .C2({ S10527 }),
  .ZN({ S10532 })
);
NAND3_X1 #() 
NAND3_X1_1066_ (
  .A1({ S10521 }),
  .A2({ S25957[397] }),
  .A3({ S10532 }),
  .ZN({ S10534 })
);
NAND4_X1 #() 
NAND4_X1_125_ (
  .A1({ S9037 }),
  .A2({ S9040 }),
  .A3({ S8938 }),
  .A4({ S8942 }),
  .ZN({ S10535 })
);
NAND3_X1 #() 
NAND3_X1_1067_ (
  .A1({ S31 }),
  .A2({ S10529 }),
  .A3({ S10527 }),
  .ZN({ S10536 })
);
AOI21_X1 #() 
AOI21_X1_573_ (
  .A({ S25957[395] }),
  .B1({ S10536 }),
  .B2({ S10535 }),
  .ZN({ S10537 })
);
NAND4_X1 #() 
NAND4_X1_126_ (
  .A1({ S8839 }),
  .A2({ S8842 }),
  .A3({ S9037 }),
  .A4({ S9040 }),
  .ZN({ S10538 })
);
NAND2_X1 #() 
NAND2_X1_912_ (
  .A1({ S21 }),
  .A2({ S10538 }),
  .ZN({ S10539 })
);
INV_X1 #() 
INV_X1_303_ (
  .A({ S10539 }),
  .ZN({ S10540 })
);
NAND2_X1 #() 
NAND2_X1_913_ (
  .A1({ S10529 }),
  .A2({ S10516 }),
  .ZN({ S10541 })
);
NOR2_X1 #() 
NOR2_X1_210_ (
  .A1({ S21 }),
  .A2({ S10541 }),
  .ZN({ S10542 })
);
OAI21_X1 #() 
OAI21_X1_513_ (
  .A({ S10526 }),
  .B1({ S10540 }),
  .B2({ S10542 }),
  .ZN({ S10543 })
);
NAND3_X1 #() 
NAND3_X1_1068_ (
  .A1({ S31 }),
  .A2({ S25957[394] }),
  .A3({ S10527 }),
  .ZN({ S10545 })
);
NAND4_X1 #() 
NAND4_X1_127_ (
  .A1({ S8839 }),
  .A2({ S8842 }),
  .A3({ S8938 }),
  .A4({ S8942 }),
  .ZN({ S10546 })
);
OAI211_X1 #() 
OAI211_X1_325_ (
  .A({ S10508 }),
  .B({ S10509 }),
  .C1({ S10511 }),
  .C2({ S10510 }),
  .ZN({ S10547 })
);
NAND3_X1 #() 
NAND3_X1_1069_ (
  .A1({ S10547 }),
  .A2({ S10529 }),
  .A3({ S10546 }),
  .ZN({ S10548 })
);
AOI21_X1 #() 
AOI21_X1_574_ (
  .A({ S21 }),
  .B1({ S10545 }),
  .B2({ S10548 }),
  .ZN({ S10549 })
);
INV_X1 #() 
INV_X1_304_ (
  .A({ S10535 }),
  .ZN({ S10550 })
);
AOI22_X1 #() 
AOI22_X1_110_ (
  .A1({ S10529 }),
  .A2({ S25957[392] }),
  .B1({ S8759 }),
  .B2({ S8762 }),
  .ZN({ S10551 })
);
INV_X1 #() 
INV_X1_305_ (
  .A({ S10551 }),
  .ZN({ S10552 })
);
OAI21_X1 #() 
OAI21_X1_514_ (
  .A({ S25957[396] }),
  .B1({ S10552 }),
  .B2({ S10550 }),
  .ZN({ S10553 })
);
OAI22_X1 #() 
OAI22_X1_24_ (
  .A1({ S10553 }),
  .A2({ S10549 }),
  .B1({ S10543 }),
  .B2({ S10537 }),
  .ZN({ S10554 })
);
OAI211_X1 #() 
OAI211_X1_326_ (
  .A({ S10534 }),
  .B({ S8507 }),
  .C1({ S25957[397] }),
  .C2({ S10554 }),
  .ZN({ S10556 })
);
NAND3_X1 #() 
NAND3_X1_1070_ (
  .A1({ S8585 }),
  .A2({ S8587 }),
  .A3({ S7605 }),
  .ZN({ S10557 })
);
OAI21_X1 #() 
OAI21_X1_515_ (
  .A({ S25957[525] }),
  .B1({ S8579 }),
  .B2({ S8583 }),
  .ZN({ S10558 })
);
NAND2_X1 #() 
NAND2_X1_914_ (
  .A1({ S10558 }),
  .A2({ S10557 }),
  .ZN({ S10559 })
);
INV_X1 #() 
INV_X1_306_ (
  .A({ S10546 }),
  .ZN({ S10560 })
);
NOR2_X1 #() 
NOR2_X1_211_ (
  .A1({ S10560 }),
  .A2({ S25957[395] }),
  .ZN({ S10561 })
);
OAI211_X1 #() 
OAI211_X1_327_ (
  .A({ S9037 }),
  .B({ S9040 }),
  .C1({ S10511 }),
  .C2({ S10510 }),
  .ZN({ S10562 })
);
NAND2_X1 #() 
NAND2_X1_915_ (
  .A1({ S10562 }),
  .A2({ S10527 }),
  .ZN({ S10563 })
);
NOR2_X1 #() 
NOR2_X1_212_ (
  .A1({ S10563 }),
  .A2({ S21 }),
  .ZN({ S10564 })
);
OR2_X1 #() 
OR2_X1_13_ (
  .A1({ S10564 }),
  .A2({ S10561 }),
  .ZN({ S10565 })
);
OAI21_X1 #() 
OAI21_X1_516_ (
  .A({ S10559 }),
  .B1({ S10565 }),
  .B2({ S10526 }),
  .ZN({ S10567 })
);
NAND3_X1 #() 
NAND3_X1_1071_ (
  .A1({ S10529 }),
  .A2({ S8938 }),
  .A3({ S8942 }),
  .ZN({ S10568 })
);
NAND2_X1 #() 
NAND2_X1_916_ (
  .A1({ S25957[392] }),
  .A2({ S10529 }),
  .ZN({ S10569 })
);
AOI22_X1 #() 
AOI22_X1_111_ (
  .A1({ S10509 }),
  .A2({ S10508 }),
  .B1({ S8938 }),
  .B2({ S8942 }),
  .ZN({ S10570 })
);
NAND2_X1 #() 
NAND2_X1_917_ (
  .A1({ S10570 }),
  .A2({ S25957[394] }),
  .ZN({ S10571 })
);
NAND4_X1 #() 
NAND4_X1_128_ (
  .A1({ S10571 }),
  .A2({ S10569 }),
  .A3({ S10568 }),
  .A4({ S21 }),
  .ZN({ S10572 })
);
NAND3_X1 #() 
NAND3_X1_1072_ (
  .A1({ S10571 }),
  .A2({ S25957[395] }),
  .A3({ S10568 }),
  .ZN({ S10573 })
);
AOI21_X1 #() 
AOI21_X1_575_ (
  .A({ S25957[396] }),
  .B1({ S10572 }),
  .B2({ S10573 }),
  .ZN({ S10574 })
);
NAND2_X1 #() 
NAND2_X1_918_ (
  .A1({ S10528 }),
  .A2({ S10529 }),
  .ZN({ S10575 })
);
NAND2_X1 #() 
NAND2_X1_919_ (
  .A1({ S10575 }),
  .A2({ S25957[393] }),
  .ZN({ S10576 })
);
NAND2_X1 #() 
NAND2_X1_920_ (
  .A1({ S10514 }),
  .A2({ S25957[395] }),
  .ZN({ S10578 })
);
AOI22_X1 #() 
AOI22_X1_112_ (
  .A1({ S8842 }),
  .A2({ S8839 }),
  .B1({ S8938 }),
  .B2({ S8942 }),
  .ZN({ S10579 })
);
NOR2_X1 #() 
NOR2_X1_213_ (
  .A1({ S10579 }),
  .A2({ S25957[394] }),
  .ZN({ S10580 })
);
AOI21_X1 #() 
AOI21_X1_576_ (
  .A({ S10526 }),
  .B1({ S10580 }),
  .B2({ S25957[395] }),
  .ZN({ S10581 })
);
OAI211_X1 #() 
OAI211_X1_328_ (
  .A({ S10581 }),
  .B({ S10578 }),
  .C1({ S10576 }),
  .C2({ S25957[395] }),
  .ZN({ S10582 })
);
AOI21_X1 #() 
AOI21_X1_577_ (
  .A({ S10529 }),
  .B1({ S10547 }),
  .B2({ S10546 }),
  .ZN({ S10583 })
);
AOI22_X1 #() 
AOI22_X1_113_ (
  .A1({ S9037 }),
  .A2({ S9040 }),
  .B1({ S8942 }),
  .B2({ S8938 }),
  .ZN({ S10584 })
);
NAND2_X1 #() 
NAND2_X1_921_ (
  .A1({ S10584 }),
  .A2({ S25957[392] }),
  .ZN({ S10585 })
);
INV_X1 #() 
INV_X1_307_ (
  .A({ S10585 }),
  .ZN({ S10586 })
);
OAI21_X1 #() 
OAI21_X1_517_ (
  .A({ S25957[395] }),
  .B1({ S10586 }),
  .B2({ S10583 }),
  .ZN({ S10587 })
);
AOI22_X1 #() 
AOI22_X1_114_ (
  .A1({ S8842 }),
  .A2({ S8839 }),
  .B1({ S9037 }),
  .B2({ S9040 }),
  .ZN({ S10589 })
);
NAND2_X1 #() 
NAND2_X1_922_ (
  .A1({ S10589 }),
  .A2({ S25957[393] }),
  .ZN({ S10590 })
);
NAND2_X1 #() 
NAND2_X1_923_ (
  .A1({ S10590 }),
  .A2({ S10571 }),
  .ZN({ S10591 })
);
NAND2_X1 #() 
NAND2_X1_924_ (
  .A1({ S10591 }),
  .A2({ S21 }),
  .ZN({ S10592 })
);
NAND3_X1 #() 
NAND3_X1_1073_ (
  .A1({ S10587 }),
  .A2({ S10592 }),
  .A3({ S10526 }),
  .ZN({ S10593 })
);
NAND3_X1 #() 
NAND3_X1_1074_ (
  .A1({ S10593 }),
  .A2({ S25957[397] }),
  .A3({ S10582 }),
  .ZN({ S10594 })
);
OAI211_X1 #() 
OAI211_X1_329_ (
  .A({ S10594 }),
  .B({ S25957[398] }),
  .C1({ S10567 }),
  .C2({ S10574 }),
  .ZN({ S10595 })
);
NAND3_X1 #() 
NAND3_X1_1075_ (
  .A1({ S10595 }),
  .A2({ S10556 }),
  .A3({ S25957[399] }),
  .ZN({ S10596 })
);
INV_X1 #() 
INV_X1_308_ (
  .A({ S8426 }),
  .ZN({ S10597 })
);
NAND2_X1 #() 
NAND2_X1_925_ (
  .A1({ S10597 }),
  .A2({ S8424 }),
  .ZN({ S10598 })
);
AOI21_X1 #() 
AOI21_X1_578_ (
  .A({ S25957[392] }),
  .B1({ S25957[394] }),
  .B2({ S10516 }),
  .ZN({ S10600 })
);
OAI21_X1 #() 
OAI21_X1_518_ (
  .A({ S25957[396] }),
  .B1({ S10600 }),
  .B2({ S25957[395] }),
  .ZN({ S10601 })
);
NOR2_X1 #() 
NOR2_X1_214_ (
  .A1({ S10591 }),
  .A2({ S21 }),
  .ZN({ S10602 })
);
NAND2_X1 #() 
NAND2_X1_926_ (
  .A1({ S10585 }),
  .A2({ S10535 }),
  .ZN({ S10603 })
);
NAND2_X1 #() 
NAND2_X1_927_ (
  .A1({ S10603 }),
  .A2({ S25957[395] }),
  .ZN({ S10604 })
);
NAND3_X1 #() 
NAND3_X1_1076_ (
  .A1({ S21 }),
  .A2({ S10562 }),
  .A3({ S10538 }),
  .ZN({ S10605 })
);
NAND3_X1 #() 
NAND3_X1_1077_ (
  .A1({ S10604 }),
  .A2({ S10526 }),
  .A3({ S10605 }),
  .ZN({ S10606 })
);
OAI21_X1 #() 
OAI21_X1_519_ (
  .A({ S10606 }),
  .B1({ S10602 }),
  .B2({ S10601 }),
  .ZN({ S10607 })
);
NAND2_X1 #() 
NAND2_X1_928_ (
  .A1({ S10607 }),
  .A2({ S25957[397] }),
  .ZN({ S10608 })
);
NAND2_X1 #() 
NAND2_X1_929_ (
  .A1({ S10527 }),
  .A2({ S25957[394] }),
  .ZN({ S10609 })
);
AOI21_X1 #() 
AOI21_X1_579_ (
  .A({ S21 }),
  .B1({ S10548 }),
  .B2({ S10609 }),
  .ZN({ S10611 })
);
NAND3_X1 #() 
NAND3_X1_1078_ (
  .A1({ S10547 }),
  .A2({ S25957[394] }),
  .A3({ S10546 }),
  .ZN({ S10612 })
);
AOI21_X1 #() 
AOI21_X1_580_ (
  .A({ S25957[395] }),
  .B1({ S10612 }),
  .B2({ S10575 }),
  .ZN({ S10613 })
);
OR3_X1 #() 
OR3_X1_3_ (
  .A1({ S10613 }),
  .A2({ S10611 }),
  .A3({ S10526 }),
  .ZN({ S10614 })
);
NAND2_X1 #() 
NAND2_X1_930_ (
  .A1({ S10568 }),
  .A2({ S25957[395] }),
  .ZN({ S10615 })
);
OAI211_X1 #() 
OAI211_X1_330_ (
  .A({ S10562 }),
  .B({ S10538 }),
  .C1({ S10579 }),
  .C2({ S25957[394] }),
  .ZN({ S10616 })
);
AOI21_X1 #() 
AOI21_X1_581_ (
  .A({ S25957[396] }),
  .B1({ S10616 }),
  .B2({ S21 }),
  .ZN({ S10617 })
);
OAI21_X1 #() 
OAI21_X1_520_ (
  .A({ S10617 }),
  .B1({ S10514 }),
  .B2({ S10615 }),
  .ZN({ S10618 })
);
NAND3_X1 #() 
NAND3_X1_1079_ (
  .A1({ S10614 }),
  .A2({ S10559 }),
  .A3({ S10618 }),
  .ZN({ S10619 })
);
AOI21_X1 #() 
AOI21_X1_582_ (
  .A({ S8507 }),
  .B1({ S10608 }),
  .B2({ S10619 }),
  .ZN({ S10620 })
);
NAND2_X1 #() 
NAND2_X1_931_ (
  .A1({ S10527 }),
  .A2({ S10529 }),
  .ZN({ S10622 })
);
NAND3_X1 #() 
NAND3_X1_1080_ (
  .A1({ S10568 }),
  .A2({ S25957[395] }),
  .A3({ S10547 }),
  .ZN({ S10623 })
);
INV_X1 #() 
INV_X1_309_ (
  .A({ S10623 }),
  .ZN({ S10624 })
);
NOR2_X1 #() 
NOR2_X1_215_ (
  .A1({ S10550 }),
  .A2({ S25957[395] }),
  .ZN({ S10625 })
);
AOI21_X1 #() 
AOI21_X1_583_ (
  .A({ S10624 }),
  .B1({ S10622 }),
  .B2({ S10625 }),
  .ZN({ S10626 })
);
OAI21_X1 #() 
OAI21_X1_521_ (
  .A({ S25957[392] }),
  .B1({ S8765 }),
  .B2({ S8764 }),
  .ZN({ S10627 })
);
NOR2_X1 #() 
NOR2_X1_216_ (
  .A1({ S10514 }),
  .A2({ S21 }),
  .ZN({ S10628 })
);
NAND2_X1 #() 
NAND2_X1_932_ (
  .A1({ S10628 }),
  .A2({ S10541 }),
  .ZN({ S10629 })
);
NAND3_X1 #() 
NAND3_X1_1081_ (
  .A1({ S10629 }),
  .A2({ S25957[396] }),
  .A3({ S10627 }),
  .ZN({ S10630 })
);
OAI211_X1 #() 
OAI211_X1_331_ (
  .A({ S25957[397] }),
  .B({ S10630 }),
  .C1({ S10626 }),
  .C2({ S25957[396] }),
  .ZN({ S10631 })
);
AOI21_X1 #() 
AOI21_X1_584_ (
  .A({ S10529 }),
  .B1({ S31 }),
  .B2({ S10527 }),
  .ZN({ S10633 })
);
NOR2_X1 #() 
NOR2_X1_217_ (
  .A1({ S10633 }),
  .A2({ S25957[395] }),
  .ZN({ S10634 })
);
AOI21_X1 #() 
AOI21_X1_585_ (
  .A({ S10634 }),
  .B1({ S10609 }),
  .B2({ S25957[395] }),
  .ZN({ S10635 })
);
NOR2_X1 #() 
NOR2_X1_218_ (
  .A1({ S10535 }),
  .A2({ S25957[392] }),
  .ZN({ S10636 })
);
NOR2_X1 #() 
NOR2_X1_219_ (
  .A1({ S10636 }),
  .A2({ S21 }),
  .ZN({ S10637 })
);
NAND2_X1 #() 
NAND2_X1_933_ (
  .A1({ S10590 }),
  .A2({ S21 }),
  .ZN({ S10638 })
);
OAI21_X1 #() 
OAI21_X1_522_ (
  .A({ S25957[396] }),
  .B1({ S10638 }),
  .B2({ S10583 }),
  .ZN({ S10639 })
);
OAI221_X1 #() 
OAI221_X1_18_ (
  .A({ S10559 }),
  .B1({ S10637 }),
  .B2({ S10639 }),
  .C1({ S10635 }),
  .C2({ S25957[396] }),
  .ZN({ S10640 })
);
AND3_X1 #() 
AND3_X1_44_ (
  .A1({ S10640 }),
  .A2({ S10631 }),
  .A3({ S8507 }),
  .ZN({ S10641 })
);
OAI21_X1 #() 
OAI21_X1_523_ (
  .A({ S10598 }),
  .B1({ S10641 }),
  .B2({ S10620 }),
  .ZN({ S10642 })
);
NAND2_X1 #() 
NAND2_X1_934_ (
  .A1({ S10642 }),
  .A2({ S10596 }),
  .ZN({ S10644 })
);
NAND2_X1 #() 
NAND2_X1_935_ (
  .A1({ S10644 }),
  .A2({ S25957[599] }),
  .ZN({ S10645 })
);
INV_X1 #() 
INV_X1_310_ (
  .A({ S10645 }),
  .ZN({ S10646 })
);
NOR2_X1 #() 
NOR2_X1_220_ (
  .A1({ S10644 }),
  .A2({ S25957[599] }),
  .ZN({ S10647 })
);
NOR2_X1 #() 
NOR2_X1_221_ (
  .A1({ S10646 }),
  .A2({ S10647 }),
  .ZN({ S10648 })
);
INV_X1 #() 
INV_X1_311_ (
  .A({ S10648 }),
  .ZN({ S25957[343] })
);
NAND2_X1 #() 
NAND2_X1_936_ (
  .A1({ S25957[343] }),
  .A2({ S25957[439] }),
  .ZN({ S10649 })
);
NAND3_X1 #() 
NAND3_X1_1082_ (
  .A1({ S10648 }),
  .A2({ S7698 }),
  .A3({ S7701 }),
  .ZN({ S10650 })
);
NAND2_X1 #() 
NAND2_X1_937_ (
  .A1({ S10649 }),
  .A2({ S10650 }),
  .ZN({ S10651 })
);
NAND2_X1 #() 
NAND2_X1_938_ (
  .A1({ S10651 }),
  .A2({ S7707 }),
  .ZN({ S10652 })
);
NAND3_X1 #() 
NAND3_X1_1083_ (
  .A1({ S10649 }),
  .A2({ S25957[407] }),
  .A3({ S10650 }),
  .ZN({ S10654 })
);
AND2_X1 #() 
AND2_X1_57_ (
  .A1({ S10652 }),
  .A2({ S10654 }),
  .ZN({ S25957[279] })
);
XNOR2_X1 #() 
XNOR2_X1_31_ (
  .A({ S25957[630] }),
  .B({ S7709 }),
  .ZN({ S25957[598] })
);
OAI22_X1 #() 
OAI22_X1_25_ (
  .A1({ S10515 }),
  .A2({ S10575 }),
  .B1({ S10535 }),
  .B2({ S21 }),
  .ZN({ S10655 })
);
INV_X1 #() 
INV_X1_312_ (
  .A({ S10655 }),
  .ZN({ S10656 })
);
OAI21_X1 #() 
OAI21_X1_524_ (
  .A({ S10656 }),
  .B1({ S25957[395] }),
  .B2({ S10612 }),
  .ZN({ S10657 })
);
NAND2_X1 #() 
NAND2_X1_939_ (
  .A1({ S10657 }),
  .A2({ S25957[396] }),
  .ZN({ S10658 })
);
NAND3_X1 #() 
NAND3_X1_1084_ (
  .A1({ S25957[393] }),
  .A2({ S10528 }),
  .A3({ S10529 }),
  .ZN({ S10659 })
);
NAND2_X1 #() 
NAND2_X1_940_ (
  .A1({ S10659 }),
  .A2({ S10562 }),
  .ZN({ S10660 })
);
NAND2_X1 #() 
NAND2_X1_941_ (
  .A1({ S21 }),
  .A2({ S10547 }),
  .ZN({ S10661 })
);
NAND2_X1 #() 
NAND2_X1_942_ (
  .A1({ S10569 }),
  .A2({ S10546 }),
  .ZN({ S10663 })
);
OAI221_X1 #() 
OAI221_X1_19_ (
  .A({ S10526 }),
  .B1({ S10663 }),
  .B2({ S10661 }),
  .C1({ S10660 }),
  .C2({ S21 }),
  .ZN({ S10664 })
);
AND2_X1 #() 
AND2_X1_58_ (
  .A1({ S10664 }),
  .A2({ S10658 }),
  .ZN({ S10665 })
);
INV_X1 #() 
INV_X1_313_ (
  .A({ S10548 }),
  .ZN({ S10666 })
);
NAND4_X1 #() 
NAND4_X1_129_ (
  .A1({ S25957[395] }),
  .A2({ S10575 }),
  .A3({ S31 }),
  .A4({ S10513 }),
  .ZN({ S10667 })
);
OAI21_X1 #() 
OAI21_X1_525_ (
  .A({ S10667 }),
  .B1({ S10666 }),
  .B2({ S10539 }),
  .ZN({ S10668 })
);
NAND2_X1 #() 
NAND2_X1_943_ (
  .A1({ S10547 }),
  .A2({ S10529 }),
  .ZN({ S10669 })
);
OAI21_X1 #() 
OAI21_X1_526_ (
  .A({ S10520 }),
  .B1({ S25957[395] }),
  .B2({ S10669 }),
  .ZN({ S10670 })
);
AOI21_X1 #() 
AOI21_X1_586_ (
  .A({ S25957[397] }),
  .B1({ S10670 }),
  .B2({ S25957[396] }),
  .ZN({ S10671 })
);
OAI21_X1 #() 
OAI21_X1_527_ (
  .A({ S10671 }),
  .B1({ S25957[396] }),
  .B2({ S10668 }),
  .ZN({ S10672 })
);
OAI21_X1 #() 
OAI21_X1_528_ (
  .A({ S10672 }),
  .B1({ S10665 }),
  .B2({ S10559 }),
  .ZN({ S10674 })
);
NAND3_X1 #() 
NAND3_X1_1085_ (
  .A1({ S10569 }),
  .A2({ S10535 }),
  .A3({ S10538 }),
  .ZN({ S10675 })
);
INV_X1 #() 
INV_X1_314_ (
  .A({ S10675 }),
  .ZN({ S10676 })
);
NOR2_X1 #() 
NOR2_X1_222_ (
  .A1({ S10676 }),
  .A2({ S21 }),
  .ZN({ S10677 })
);
AOI21_X1 #() 
AOI21_X1_587_ (
  .A({ S10677 }),
  .B1({ S10548 }),
  .B2({ S10540 }),
  .ZN({ S10678 })
);
NAND2_X1 #() 
NAND2_X1_944_ (
  .A1({ S10678 }),
  .A2({ S25957[396] }),
  .ZN({ S10679 })
);
NAND2_X1 #() 
NAND2_X1_945_ (
  .A1({ S10679 }),
  .A2({ S10559 }),
  .ZN({ S10680 })
);
AOI22_X1 #() 
AOI22_X1_115_ (
  .A1({ S10527 }),
  .A2({ S25957[394] }),
  .B1({ S8762 }),
  .B2({ S8759 }),
  .ZN({ S10681 })
);
AOI21_X1 #() 
AOI21_X1_588_ (
  .A({ S10542 }),
  .B1({ S10669 }),
  .B2({ S10681 }),
  .ZN({ S10682 })
);
NAND3_X1 #() 
NAND3_X1_1086_ (
  .A1({ S25957[395] }),
  .A2({ S10528 }),
  .A3({ S10535 }),
  .ZN({ S10683 })
);
AOI21_X1 #() 
AOI21_X1_589_ (
  .A({ S25957[396] }),
  .B1({ S10682 }),
  .B2({ S10683 }),
  .ZN({ S10685 })
);
NAND2_X1 #() 
NAND2_X1_946_ (
  .A1({ S10515 }),
  .A2({ S10526 }),
  .ZN({ S10686 })
);
OAI21_X1 #() 
OAI21_X1_529_ (
  .A({ S25957[396] }),
  .B1({ S10568 }),
  .B2({ S21 }),
  .ZN({ S10687 })
);
INV_X1 #() 
INV_X1_315_ (
  .A({ S10687 }),
  .ZN({ S10688 })
);
NAND2_X1 #() 
NAND2_X1_947_ (
  .A1({ S31 }),
  .A2({ S25957[394] }),
  .ZN({ S10689 })
);
NAND2_X1 #() 
NAND2_X1_948_ (
  .A1({ S10689 }),
  .A2({ S21 }),
  .ZN({ S10690 })
);
OAI211_X1 #() 
OAI211_X1_332_ (
  .A({ S10688 }),
  .B({ S10690 }),
  .C1({ S21 }),
  .C2({ S10676 }),
  .ZN({ S10691 })
);
OAI211_X1 #() 
OAI211_X1_333_ (
  .A({ S10691 }),
  .B({ S25957[397] }),
  .C1({ S10564 }),
  .C2({ S10686 }),
  .ZN({ S10692 })
);
OAI211_X1 #() 
OAI211_X1_334_ (
  .A({ S25957[398] }),
  .B({ S10692 }),
  .C1({ S10680 }),
  .C2({ S10685 }),
  .ZN({ S10693 })
);
OAI211_X1 #() 
OAI211_X1_335_ (
  .A({ S10693 }),
  .B({ S25957[399] }),
  .C1({ S25957[398] }),
  .C2({ S10674 }),
  .ZN({ S10694 })
);
AOI22_X1 #() 
AOI22_X1_116_ (
  .A1({ S25957[393] }),
  .A2({ S25957[392] }),
  .B1({ S9037 }),
  .B2({ S9040 }),
  .ZN({ S10696 })
);
OAI21_X1 #() 
OAI21_X1_530_ (
  .A({ S25957[395] }),
  .B1({ S10583 }),
  .B2({ S10696 }),
  .ZN({ S10697 })
);
NAND3_X1 #() 
NAND3_X1_1087_ (
  .A1({ S10697 }),
  .A2({ S25957[396] }),
  .A3({ S10552 }),
  .ZN({ S10698 })
);
NOR2_X1 #() 
NOR2_X1_223_ (
  .A1({ S25957[393] }),
  .A2({ S10529 }),
  .ZN({ S10699 })
);
OAI22_X1 #() 
OAI22_X1_26_ (
  .A1({ S25957[395] }),
  .A2({ S10603 }),
  .B1({ S10615 }),
  .B2({ S10699 }),
  .ZN({ S10700 })
);
OAI21_X1 #() 
OAI21_X1_531_ (
  .A({ S10698 }),
  .B1({ S10700 }),
  .B2({ S25957[396] }),
  .ZN({ S10701 })
);
AOI22_X1 #() 
AOI22_X1_117_ (
  .A1({ S10584 }),
  .A2({ S25957[392] }),
  .B1({ S8762 }),
  .B2({ S8759 }),
  .ZN({ S10702 })
);
AOI211_X1 #() 
AOI211_X1_11_ (
  .A({ S10526 }),
  .B({ S10702 }),
  .C1({ S25957[395] }),
  .C2({ S10603 }),
  .ZN({ S10703 })
);
NAND2_X1 #() 
NAND2_X1_949_ (
  .A1({ S10569 }),
  .A2({ S10541 }),
  .ZN({ S10704 })
);
OAI211_X1 #() 
OAI211_X1_336_ (
  .A({ S25957[395] }),
  .B({ S10526 }),
  .C1({ S10704 }),
  .C2({ S10636 }),
  .ZN({ S10705 })
);
INV_X1 #() 
INV_X1_316_ (
  .A({ S10705 }),
  .ZN({ S10707 })
);
OAI21_X1 #() 
OAI21_X1_532_ (
  .A({ S10559 }),
  .B1({ S10703 }),
  .B2({ S10707 }),
  .ZN({ S10708 })
);
OAI21_X1 #() 
OAI21_X1_533_ (
  .A({ S10708 }),
  .B1({ S10701 }),
  .B2({ S10559 }),
  .ZN({ S10709 })
);
AOI211_X1 #() 
AOI211_X1_12_ (
  .A({ S25957[396] }),
  .B({ S10677 }),
  .C1({ S21 }),
  .C2({ S10545 }),
  .ZN({ S10710 })
);
NAND2_X1 #() 
NAND2_X1_950_ (
  .A1({ S10513 }),
  .A2({ S10546 }),
  .ZN({ S10711 })
);
AOI22_X1 #() 
AOI22_X1_118_ (
  .A1({ S10551 }),
  .A2({ S10609 }),
  .B1({ S10711 }),
  .B2({ S25957[395] }),
  .ZN({ S10712 })
);
NAND2_X1 #() 
NAND2_X1_951_ (
  .A1({ S10569 }),
  .A2({ S25957[393] }),
  .ZN({ S10713 })
);
INV_X1 #() 
INV_X1_317_ (
  .A({ S10713 }),
  .ZN({ S10714 })
);
NAND2_X1 #() 
NAND2_X1_952_ (
  .A1({ S10578 }),
  .A2({ S10526 }),
  .ZN({ S10715 })
);
OAI22_X1 #() 
OAI22_X1_27_ (
  .A1({ S10712 }),
  .A2({ S10526 }),
  .B1({ S10715 }),
  .B2({ S10714 }),
  .ZN({ S10716 })
);
NAND2_X1 #() 
NAND2_X1_953_ (
  .A1({ S10541 }),
  .A2({ S10528 }),
  .ZN({ S10718 })
);
NOR2_X1 #() 
NOR2_X1_224_ (
  .A1({ S10718 }),
  .A2({ S25957[395] }),
  .ZN({ S10719 })
);
OAI21_X1 #() 
OAI21_X1_534_ (
  .A({ S10559 }),
  .B1({ S10719 }),
  .B2({ S10687 }),
  .ZN({ S10720 })
);
OAI221_X1 #() 
OAI221_X1_20_ (
  .A({ S25957[398] }),
  .B1({ S10559 }),
  .B2({ S10716 }),
  .C1({ S10710 }),
  .C2({ S10720 }),
  .ZN({ S10721 })
);
OAI211_X1 #() 
OAI211_X1_337_ (
  .A({ S10721 }),
  .B({ S10598 }),
  .C1({ S25957[398] }),
  .C2({ S10709 }),
  .ZN({ S10722 })
);
NAND2_X1 #() 
NAND2_X1_954_ (
  .A1({ S10694 }),
  .A2({ S10722 }),
  .ZN({ S10723 })
);
NOR2_X1 #() 
NOR2_X1_225_ (
  .A1({ S10723 }),
  .A2({ S25957[598] }),
  .ZN({ S10724 })
);
AND2_X1 #() 
AND2_X1_59_ (
  .A1({ S10723 }),
  .A2({ S25957[598] }),
  .ZN({ S10725 })
);
NOR2_X1 #() 
NOR2_X1_226_ (
  .A1({ S10725 }),
  .A2({ S10724 }),
  .ZN({ S10726 })
);
XNOR2_X1 #() 
XNOR2_X1_32_ (
  .A({ S10726 }),
  .B({ S25957[534] }),
  .ZN({ S25957[278] })
);
NAND2_X1 #() 
NAND2_X1_955_ (
  .A1({ S5065 }),
  .A2({ S5064 }),
  .ZN({ S10728 })
);
NAND2_X1 #() 
NAND2_X1_956_ (
  .A1({ S10538 }),
  .A2({ S10546 }),
  .ZN({ S10729 })
);
AOI22_X1 #() 
AOI22_X1_119_ (
  .A1({ S10561 }),
  .A2({ S10669 }),
  .B1({ S25957[395] }),
  .B2({ S10729 }),
  .ZN({ S10730 })
);
NAND2_X1 #() 
NAND2_X1_957_ (
  .A1({ S10513 }),
  .A2({ S10516 }),
  .ZN({ S10731 })
);
NAND2_X1 #() 
NAND2_X1_958_ (
  .A1({ S10731 }),
  .A2({ S21 }),
  .ZN({ S10732 })
);
NAND4_X1 #() 
NAND4_X1_130_ (
  .A1({ S10546 }),
  .A2({ S25957[394] }),
  .A3({ S8762 }),
  .A4({ S8759 }),
  .ZN({ S10733 })
);
NAND2_X1 #() 
NAND2_X1_959_ (
  .A1({ S10696 }),
  .A2({ S25957[395] }),
  .ZN({ S10734 })
);
NAND3_X1 #() 
NAND3_X1_1088_ (
  .A1({ S10734 }),
  .A2({ S10732 }),
  .A3({ S10733 }),
  .ZN({ S10735 })
);
AND2_X1 #() 
AND2_X1_60_ (
  .A1({ S10735 }),
  .A2({ S10526 }),
  .ZN({ S10736 })
);
AOI211_X1 #() 
AOI211_X1_13_ (
  .A({ S10559 }),
  .B({ S10736 }),
  .C1({ S25957[396] }),
  .C2({ S10730 }),
  .ZN({ S10737 })
);
NAND2_X1 #() 
NAND2_X1_960_ (
  .A1({ S10546 }),
  .A2({ S25957[394] }),
  .ZN({ S10739 })
);
NAND2_X1 #() 
NAND2_X1_961_ (
  .A1({ S10560 }),
  .A2({ S25957[395] }),
  .ZN({ S10740 })
);
AOI21_X1 #() 
AOI21_X1_590_ (
  .A({ S10526 }),
  .B1({ S10740 }),
  .B2({ S10739 }),
  .ZN({ S10741 })
);
NOR3_X1 #() 
NOR3_X1_30_ (
  .A1({ S10634 }),
  .A2({ S10676 }),
  .A3({ S25957[396] }),
  .ZN({ S10742 })
);
OR2_X1 #() 
OR2_X1_14_ (
  .A1({ S10742 }),
  .A2({ S10741 }),
  .ZN({ S10743 })
);
OAI21_X1 #() 
OAI21_X1_535_ (
  .A({ S25957[398] }),
  .B1({ S10743 }),
  .B2({ S25957[397] }),
  .ZN({ S10744 })
);
NAND3_X1 #() 
NAND3_X1_1089_ (
  .A1({ S10575 }),
  .A2({ S21 }),
  .A3({ S10527 }),
  .ZN({ S10745 })
);
OAI211_X1 #() 
OAI211_X1_338_ (
  .A({ S25957[396] }),
  .B({ S10745 }),
  .C1({ S10616 }),
  .C2({ S21 }),
  .ZN({ S10746 })
);
AOI21_X1 #() 
AOI21_X1_591_ (
  .A({ S10518 }),
  .B1({ S10563 }),
  .B2({ S21 }),
  .ZN({ S10747 })
);
AOI21_X1 #() 
AOI21_X1_592_ (
  .A({ S10559 }),
  .B1({ S10747 }),
  .B2({ S10526 }),
  .ZN({ S10748 })
);
INV_X1 #() 
INV_X1_318_ (
  .A({ S10530 }),
  .ZN({ S10750 })
);
OAI21_X1 #() 
OAI21_X1_536_ (
  .A({ S25957[395] }),
  .B1({ S10583 }),
  .B2({ S10750 }),
  .ZN({ S10751 })
);
NAND3_X1 #() 
NAND3_X1_1090_ (
  .A1({ S10751 }),
  .A2({ S10526 }),
  .A3({ S10638 }),
  .ZN({ S10752 })
);
AOI21_X1 #() 
AOI21_X1_593_ (
  .A({ S25957[394] }),
  .B1({ S10547 }),
  .B2({ S10546 }),
  .ZN({ S10753 })
);
NAND2_X1 #() 
NAND2_X1_962_ (
  .A1({ S10753 }),
  .A2({ S25957[395] }),
  .ZN({ S10754 })
);
AOI21_X1 #() 
AOI21_X1_594_ (
  .A({ S25957[393] }),
  .B1({ S25957[392] }),
  .B2({ S10529 }),
  .ZN({ S10755 })
);
NAND2_X1 #() 
NAND2_X1_963_ (
  .A1({ S10755 }),
  .A2({ S21 }),
  .ZN({ S10756 })
);
NAND2_X1 #() 
NAND2_X1_964_ (
  .A1({ S10754 }),
  .A2({ S10756 }),
  .ZN({ S10757 })
);
AOI21_X1 #() 
AOI21_X1_595_ (
  .A({ S25957[397] }),
  .B1({ S10757 }),
  .B2({ S25957[396] }),
  .ZN({ S10758 })
);
AOI22_X1 #() 
AOI22_X1_120_ (
  .A1({ S10758 }),
  .A2({ S10752 }),
  .B1({ S10746 }),
  .B2({ S10748 }),
  .ZN({ S10759 })
);
OAI22_X1 #() 
OAI22_X1_28_ (
  .A1({ S10737 }),
  .A2({ S10744 }),
  .B1({ S10759 }),
  .B2({ S25957[398] }),
  .ZN({ S10761 })
);
INV_X1 #() 
INV_X1_319_ (
  .A({ S10581 }),
  .ZN({ S10762 })
);
NAND2_X1 #() 
NAND2_X1_965_ (
  .A1({ S10562 }),
  .A2({ S10538 }),
  .ZN({ S10763 })
);
NAND2_X1 #() 
NAND2_X1_966_ (
  .A1({ S25957[395] }),
  .A2({ S10569 }),
  .ZN({ S10764 })
);
NAND2_X1 #() 
NAND2_X1_967_ (
  .A1({ S10659 }),
  .A2({ S21 }),
  .ZN({ S10765 })
);
OAI21_X1 #() 
OAI21_X1_537_ (
  .A({ S10765 }),
  .B1({ S10764 }),
  .B2({ S10763 }),
  .ZN({ S10766 })
);
NAND2_X1 #() 
NAND2_X1_968_ (
  .A1({ S10766 }),
  .A2({ S10526 }),
  .ZN({ S10767 })
);
AOI21_X1 #() 
AOI21_X1_596_ (
  .A({ S10513 }),
  .B1({ S25957[395] }),
  .B2({ S25957[393] }),
  .ZN({ S10768 })
);
NOR2_X1 #() 
NOR2_X1_227_ (
  .A1({ S10535 }),
  .A2({ S10528 }),
  .ZN({ S10769 })
);
NOR3_X1 #() 
NOR3_X1_31_ (
  .A1({ S10696 }),
  .A2({ S10769 }),
  .A3({ S25957[395] }),
  .ZN({ S10770 })
);
OAI22_X1 #() 
OAI22_X1_29_ (
  .A1({ S10767 }),
  .A2({ S10768 }),
  .B1({ S10770 }),
  .B2({ S10762 }),
  .ZN({ S10772 })
);
OAI211_X1 #() 
OAI211_X1_339_ (
  .A({ S21 }),
  .B({ S10562 }),
  .C1({ S10579 }),
  .C2({ S25957[394] }),
  .ZN({ S10773 })
);
NAND3_X1 #() 
NAND3_X1_1091_ (
  .A1({ S10612 }),
  .A2({ S25957[395] }),
  .A3({ S10659 }),
  .ZN({ S10774 })
);
NAND3_X1 #() 
NAND3_X1_1092_ (
  .A1({ S10774 }),
  .A2({ S25957[396] }),
  .A3({ S10773 }),
  .ZN({ S10775 })
);
NOR2_X1 #() 
NOR2_X1_228_ (
  .A1({ S21 }),
  .A2({ S25957[392] }),
  .ZN({ S10776 })
);
NAND2_X1 #() 
NAND2_X1_969_ (
  .A1({ S10551 }),
  .A2({ S10546 }),
  .ZN({ S10777 })
);
INV_X1 #() 
INV_X1_320_ (
  .A({ S10777 }),
  .ZN({ S10778 })
);
OAI21_X1 #() 
OAI21_X1_538_ (
  .A({ S10526 }),
  .B1({ S10778 }),
  .B2({ S10776 }),
  .ZN({ S10779 })
);
NAND3_X1 #() 
NAND3_X1_1093_ (
  .A1({ S10779 }),
  .A2({ S10775 }),
  .A3({ S25957[397] }),
  .ZN({ S10780 })
);
OAI211_X1 #() 
OAI211_X1_340_ (
  .A({ S25957[398] }),
  .B({ S10780 }),
  .C1({ S10772 }),
  .C2({ S25957[397] }),
  .ZN({ S10781 })
);
NAND3_X1 #() 
NAND3_X1_1094_ (
  .A1({ S10612 }),
  .A2({ S25957[395] }),
  .A3({ S10585 }),
  .ZN({ S10783 })
);
NAND3_X1 #() 
NAND3_X1_1095_ (
  .A1({ S10545 }),
  .A2({ S21 }),
  .A3({ S10622 }),
  .ZN({ S10784 })
);
NAND3_X1 #() 
NAND3_X1_1096_ (
  .A1({ S10783 }),
  .A2({ S25957[396] }),
  .A3({ S10784 }),
  .ZN({ S10785 })
);
NAND3_X1 #() 
NAND3_X1_1097_ (
  .A1({ S25957[393] }),
  .A2({ S8759 }),
  .A3({ S8762 }),
  .ZN({ S10786 })
);
INV_X1 #() 
INV_X1_321_ (
  .A({ S10625 }),
  .ZN({ S10787 })
);
NOR2_X1 #() 
NOR2_X1_229_ (
  .A1({ S25957[396] }),
  .A2({ S10528 }),
  .ZN({ S10788 })
);
NAND3_X1 #() 
NAND3_X1_1098_ (
  .A1({ S10787 }),
  .A2({ S10786 }),
  .A3({ S10788 }),
  .ZN({ S10789 })
);
NAND3_X1 #() 
NAND3_X1_1099_ (
  .A1({ S10785 }),
  .A2({ S10559 }),
  .A3({ S10789 }),
  .ZN({ S10790 })
);
OAI211_X1 #() 
OAI211_X1_341_ (
  .A({ S10578 }),
  .B({ S10526 }),
  .C1({ S10713 }),
  .C2({ S10539 }),
  .ZN({ S10791 })
);
NAND3_X1 #() 
NAND3_X1_1100_ (
  .A1({ S10734 }),
  .A2({ S25957[396] }),
  .A3({ S10765 }),
  .ZN({ S10792 })
);
AND2_X1 #() 
AND2_X1_61_ (
  .A1({ S10792 }),
  .A2({ S10791 }),
  .ZN({ S10794 })
);
OAI211_X1 #() 
OAI211_X1_342_ (
  .A({ S8507 }),
  .B({ S10790 }),
  .C1({ S10794 }),
  .C2({ S10559 }),
  .ZN({ S10795 })
);
NAND3_X1 #() 
NAND3_X1_1101_ (
  .A1({ S10781 }),
  .A2({ S10598 }),
  .A3({ S10795 }),
  .ZN({ S10796 })
);
OAI211_X1 #() 
OAI211_X1_343_ (
  .A({ S10796 }),
  .B({ S25957[501] }),
  .C1({ S10761 }),
  .C2({ S10598 }),
  .ZN({ S10797 })
);
INV_X1 #() 
INV_X1_322_ (
  .A({ S25957[501] }),
  .ZN({ S10798 })
);
NAND2_X1 #() 
NAND2_X1_970_ (
  .A1({ S10761 }),
  .A2({ S25957[399] }),
  .ZN({ S10799 })
);
NAND2_X1 #() 
NAND2_X1_971_ (
  .A1({ S10781 }),
  .A2({ S10795 }),
  .ZN({ S10800 })
);
NAND2_X1 #() 
NAND2_X1_972_ (
  .A1({ S10800 }),
  .A2({ S10598 }),
  .ZN({ S10801 })
);
NAND3_X1 #() 
NAND3_X1_1102_ (
  .A1({ S10799 }),
  .A2({ S10801 }),
  .A3({ S10798 }),
  .ZN({ S10802 })
);
NAND2_X1 #() 
NAND2_X1_973_ (
  .A1({ S10802 }),
  .A2({ S10797 }),
  .ZN({ S25957[373] })
);
NAND2_X1 #() 
NAND2_X1_974_ (
  .A1({ S25957[373] }),
  .A2({ S10728 }),
  .ZN({ S10804 })
);
INV_X1 #() 
INV_X1_323_ (
  .A({ S10728 }),
  .ZN({ S25957[565] })
);
NAND3_X1 #() 
NAND3_X1_1103_ (
  .A1({ S10802 }),
  .A2({ S10797 }),
  .A3({ S25957[565] }),
  .ZN({ S10805 })
);
NAND3_X1 #() 
NAND3_X1_1104_ (
  .A1({ S10804 }),
  .A2({ S10805 }),
  .A3({ S25957[405] }),
  .ZN({ S10806 })
);
INV_X1 #() 
INV_X1_324_ (
  .A({ S25957[405] }),
  .ZN({ S10807 })
);
NAND2_X1 #() 
NAND2_X1_975_ (
  .A1({ S25957[373] }),
  .A2({ S25957[565] }),
  .ZN({ S10808 })
);
NAND3_X1 #() 
NAND3_X1_1105_ (
  .A1({ S10802 }),
  .A2({ S10797 }),
  .A3({ S10728 }),
  .ZN({ S10809 })
);
NAND3_X1 #() 
NAND3_X1_1106_ (
  .A1({ S10808 }),
  .A2({ S10809 }),
  .A3({ S10807 }),
  .ZN({ S10810 })
);
NAND2_X1 #() 
NAND2_X1_976_ (
  .A1({ S10806 }),
  .A2({ S10810 }),
  .ZN({ S25957[277] })
);
NAND2_X1 #() 
NAND2_X1_977_ (
  .A1({ S7958 }),
  .A2({ S7955 }),
  .ZN({ S10811 })
);
INV_X1 #() 
INV_X1_325_ (
  .A({ S10811 }),
  .ZN({ S25957[436] })
);
NOR2_X1 #() 
NOR2_X1_230_ (
  .A1({ S7957 }),
  .A2({ S7956 }),
  .ZN({ S10813 })
);
INV_X1 #() 
INV_X1_326_ (
  .A({ S10813 }),
  .ZN({ S25957[468] })
);
XNOR2_X1 #() 
XNOR2_X1_33_ (
  .A({ S5122 }),
  .B({ S25957[756] }),
  .ZN({ S25957[628] })
);
NAND2_X1 #() 
NAND2_X1_978_ (
  .A1({ S7913 }),
  .A2({ S7942 }),
  .ZN({ S10814 })
);
XNOR2_X1 #() 
XNOR2_X1_34_ (
  .A({ S10814 }),
  .B({ S25957[628] }),
  .ZN({ S25957[500] })
);
INV_X1 #() 
INV_X1_327_ (
  .A({ S25957[500] }),
  .ZN({ S10815 })
);
AOI21_X1 #() 
AOI21_X1_597_ (
  .A({ S10526 }),
  .B1({ S144 }),
  .B2({ S10529 }),
  .ZN({ S10816 })
);
OAI21_X1 #() 
OAI21_X1_539_ (
  .A({ S10520 }),
  .B1({ S10584 }),
  .B2({ S10690 }),
  .ZN({ S10817 })
);
NAND3_X1 #() 
NAND3_X1_1107_ (
  .A1({ S10590 }),
  .A2({ S21 }),
  .A3({ S10538 }),
  .ZN({ S10818 })
);
AOI21_X1 #() 
AOI21_X1_598_ (
  .A({ S25957[396] }),
  .B1({ S25957[395] }),
  .B2({ S25957[394] }),
  .ZN({ S10820 })
);
AOI21_X1 #() 
AOI21_X1_599_ (
  .A({ S25957[397] }),
  .B1({ S10818 }),
  .B2({ S10820 }),
  .ZN({ S10821 })
);
OAI21_X1 #() 
OAI21_X1_540_ (
  .A({ S10821 }),
  .B1({ S10817 }),
  .B2({ S10526 }),
  .ZN({ S10822 })
);
AOI21_X1 #() 
AOI21_X1_600_ (
  .A({ S10529 }),
  .B1({ S25957[393] }),
  .B2({ S10528 }),
  .ZN({ S10823 })
);
OAI21_X1 #() 
OAI21_X1_541_ (
  .A({ S21 }),
  .B1({ S10753 }),
  .B2({ S10823 }),
  .ZN({ S10824 })
);
NOR2_X1 #() 
NOR2_X1_231_ (
  .A1({ S10589 }),
  .A2({ S21 }),
  .ZN({ S10825 })
);
AOI21_X1 #() 
AOI21_X1_601_ (
  .A({ S25957[396] }),
  .B1({ S10825 }),
  .B2({ S10609 }),
  .ZN({ S10826 })
);
NAND2_X1 #() 
NAND2_X1_979_ (
  .A1({ S10824 }),
  .A2({ S10826 }),
  .ZN({ S10827 })
);
NAND2_X1 #() 
NAND2_X1_980_ (
  .A1({ S10827 }),
  .A2({ S25957[397] }),
  .ZN({ S10828 })
);
OAI21_X1 #() 
OAI21_X1_542_ (
  .A({ S10822 }),
  .B1({ S10828 }),
  .B2({ S10816 }),
  .ZN({ S10829 })
);
NAND2_X1 #() 
NAND2_X1_981_ (
  .A1({ S10739 }),
  .A2({ S21 }),
  .ZN({ S10831 })
);
OAI211_X1 #() 
OAI211_X1_344_ (
  .A({ S10831 }),
  .B({ S25957[396] }),
  .C1({ S10603 }),
  .C2({ S21 }),
  .ZN({ S10832 })
);
OAI221_X1 #() 
OAI221_X1_21_ (
  .A({ S10526 }),
  .B1({ S10627 }),
  .B2({ S10516 }),
  .C1({ S10536 }),
  .C2({ S21 }),
  .ZN({ S10833 })
);
NAND3_X1 #() 
NAND3_X1_1108_ (
  .A1({ S10832 }),
  .A2({ S10833 }),
  .A3({ S25957[397] }),
  .ZN({ S10834 })
);
NAND3_X1 #() 
NAND3_X1_1109_ (
  .A1({ S25957[395] }),
  .A2({ S31 }),
  .A3({ S10513 }),
  .ZN({ S10835 })
);
NAND2_X1 #() 
NAND2_X1_982_ (
  .A1({ S10572 }),
  .A2({ S10835 }),
  .ZN({ S10836 })
);
NAND2_X1 #() 
NAND2_X1_983_ (
  .A1({ S10628 }),
  .A2({ S10669 }),
  .ZN({ S10837 })
);
AOI21_X1 #() 
AOI21_X1_602_ (
  .A({ S10526 }),
  .B1({ S10563 }),
  .B2({ S21 }),
  .ZN({ S10838 })
);
AOI22_X1 #() 
AOI22_X1_121_ (
  .A1({ S10836 }),
  .A2({ S10526 }),
  .B1({ S10837 }),
  .B2({ S10838 }),
  .ZN({ S10839 })
);
OAI211_X1 #() 
OAI211_X1_345_ (
  .A({ S8507 }),
  .B({ S10834 }),
  .C1({ S10839 }),
  .C2({ S25957[397] }),
  .ZN({ S10840 })
);
OAI211_X1 #() 
OAI211_X1_346_ (
  .A({ S10840 }),
  .B({ S10598 }),
  .C1({ S10829 }),
  .C2({ S8507 }),
  .ZN({ S10842 })
);
OAI22_X1 #() 
OAI22_X1_30_ (
  .A1({ S10538 }),
  .A2({ S25957[393] }),
  .B1({ S8765 }),
  .B2({ S8764 }),
  .ZN({ S10843 })
);
NAND2_X1 #() 
NAND2_X1_984_ (
  .A1({ S10581 }),
  .A2({ S10843 }),
  .ZN({ S10844 })
);
NAND3_X1 #() 
NAND3_X1_1110_ (
  .A1({ S10568 }),
  .A2({ S21 }),
  .A3({ S10528 }),
  .ZN({ S10845 })
);
NAND3_X1 #() 
NAND3_X1_1111_ (
  .A1({ S10629 }),
  .A2({ S10526 }),
  .A3({ S10845 }),
  .ZN({ S10846 })
);
NAND3_X1 #() 
NAND3_X1_1112_ (
  .A1({ S10846 }),
  .A2({ S25957[397] }),
  .A3({ S10844 }),
  .ZN({ S10847 })
);
OAI21_X1 #() 
OAI21_X1_543_ (
  .A({ S10838 }),
  .B1({ S10589 }),
  .B2({ S10517 }),
  .ZN({ S10848 })
);
NAND3_X1 #() 
NAND3_X1_1113_ (
  .A1({ S21 }),
  .A2({ S10541 }),
  .A3({ S10538 }),
  .ZN({ S10849 })
);
NAND3_X1 #() 
NAND3_X1_1114_ (
  .A1({ S10623 }),
  .A2({ S10526 }),
  .A3({ S10849 }),
  .ZN({ S10850 })
);
NAND3_X1 #() 
NAND3_X1_1115_ (
  .A1({ S10848 }),
  .A2({ S10559 }),
  .A3({ S10850 }),
  .ZN({ S10851 })
);
NAND3_X1 #() 
NAND3_X1_1116_ (
  .A1({ S10847 }),
  .A2({ S10851 }),
  .A3({ S25957[398] }),
  .ZN({ S10852 })
);
NAND4_X1 #() 
NAND4_X1_131_ (
  .A1({ S10569 }),
  .A2({ S21 }),
  .A3({ S31 }),
  .A4({ S10535 }),
  .ZN({ S10853 })
);
NAND2_X1 #() 
NAND2_X1_985_ (
  .A1({ S10547 }),
  .A2({ S25957[394] }),
  .ZN({ S10854 })
);
NAND3_X1 #() 
NAND3_X1_1117_ (
  .A1({ S10548 }),
  .A2({ S25957[395] }),
  .A3({ S10854 }),
  .ZN({ S10855 })
);
NAND3_X1 #() 
NAND3_X1_1118_ (
  .A1({ S10855 }),
  .A2({ S25957[396] }),
  .A3({ S10853 }),
  .ZN({ S10856 })
);
AOI21_X1 #() 
AOI21_X1_603_ (
  .A({ S25957[395] }),
  .B1({ S10548 }),
  .B2({ S10609 }),
  .ZN({ S10857 })
);
NAND3_X1 #() 
NAND3_X1_1119_ (
  .A1({ S25957[395] }),
  .A2({ S10529 }),
  .A3({ S10547 }),
  .ZN({ S10858 })
);
NAND2_X1 #() 
NAND2_X1_986_ (
  .A1({ S10858 }),
  .A2({ S10740 }),
  .ZN({ S10859 })
);
OAI21_X1 #() 
OAI21_X1_544_ (
  .A({ S10526 }),
  .B1({ S10857 }),
  .B2({ S10859 }),
  .ZN({ S10860 })
);
AOI21_X1 #() 
AOI21_X1_604_ (
  .A({ S10559 }),
  .B1({ S10860 }),
  .B2({ S10856 }),
  .ZN({ S10861 })
);
OAI21_X1 #() 
OAI21_X1_545_ (
  .A({ S21 }),
  .B1({ S10696 }),
  .B2({ S10823 }),
  .ZN({ S10863 })
);
OAI21_X1 #() 
OAI21_X1_546_ (
  .A({ S10863 }),
  .B1({ S10563 }),
  .B2({ S10615 }),
  .ZN({ S10864 })
);
NAND4_X1 #() 
NAND4_X1_132_ (
  .A1({ S10575 }),
  .A2({ S21 }),
  .A3({ S31 }),
  .A4({ S10513 }),
  .ZN({ S10865 })
);
OAI211_X1 #() 
OAI211_X1_347_ (
  .A({ S10516 }),
  .B({ S10529 }),
  .C1({ S8765 }),
  .C2({ S8764 }),
  .ZN({ S10866 })
);
NOR2_X1 #() 
NOR2_X1_232_ (
  .A1({ S10514 }),
  .A2({ S10517 }),
  .ZN({ S10867 })
);
NOR2_X1 #() 
NOR2_X1_233_ (
  .A1({ S10867 }),
  .A2({ S25957[396] }),
  .ZN({ S10868 })
);
NAND3_X1 #() 
NAND3_X1_1120_ (
  .A1({ S10868 }),
  .A2({ S10865 }),
  .A3({ S10866 }),
  .ZN({ S10869 })
);
OAI21_X1 #() 
OAI21_X1_547_ (
  .A({ S10869 }),
  .B1({ S10526 }),
  .B2({ S10864 }),
  .ZN({ S10870 })
);
OAI21_X1 #() 
OAI21_X1_548_ (
  .A({ S8507 }),
  .B1({ S10870 }),
  .B2({ S25957[397] }),
  .ZN({ S10871 })
);
OAI211_X1 #() 
OAI211_X1_348_ (
  .A({ S10852 }),
  .B({ S25957[399] }),
  .C1({ S10871 }),
  .C2({ S10861 }),
  .ZN({ S10872 })
);
NAND3_X1 #() 
NAND3_X1_1121_ (
  .A1({ S10872 }),
  .A2({ S10842 }),
  .A3({ S10815 }),
  .ZN({ S10874 })
);
NAND2_X1 #() 
NAND2_X1_987_ (
  .A1({ S10829 }),
  .A2({ S25957[398] }),
  .ZN({ S10875 })
);
OAI21_X1 #() 
OAI21_X1_549_ (
  .A({ S10834 }),
  .B1({ S10839 }),
  .B2({ S25957[397] }),
  .ZN({ S10876 })
);
NAND2_X1 #() 
NAND2_X1_988_ (
  .A1({ S10876 }),
  .A2({ S8507 }),
  .ZN({ S10877 })
);
NAND3_X1 #() 
NAND3_X1_1122_ (
  .A1({ S10875 }),
  .A2({ S10877 }),
  .A3({ S10598 }),
  .ZN({ S10878 })
);
NAND2_X1 #() 
NAND2_X1_989_ (
  .A1({ S10847 }),
  .A2({ S10851 }),
  .ZN({ S10879 })
);
NAND2_X1 #() 
NAND2_X1_990_ (
  .A1({ S10879 }),
  .A2({ S25957[398] }),
  .ZN({ S10880 })
);
NAND3_X1 #() 
NAND3_X1_1123_ (
  .A1({ S10855 }),
  .A2({ S25957[397] }),
  .A3({ S10853 }),
  .ZN({ S10881 })
);
NAND2_X1 #() 
NAND2_X1_991_ (
  .A1({ S10864 }),
  .A2({ S10559 }),
  .ZN({ S10882 })
);
NAND3_X1 #() 
NAND3_X1_1124_ (
  .A1({ S10882 }),
  .A2({ S25957[396] }),
  .A3({ S10881 }),
  .ZN({ S10883 })
);
NAND2_X1 #() 
NAND2_X1_992_ (
  .A1({ S10546 }),
  .A2({ S10529 }),
  .ZN({ S10885 })
);
NAND3_X1 #() 
NAND3_X1_1125_ (
  .A1({ S25957[394] }),
  .A2({ S25957[393] }),
  .A3({ S10528 }),
  .ZN({ S10886 })
);
AOI21_X1 #() 
AOI21_X1_605_ (
  .A({ S25957[395] }),
  .B1({ S10886 }),
  .B2({ S10885 }),
  .ZN({ S10887 })
);
OAI21_X1 #() 
OAI21_X1_550_ (
  .A({ S10559 }),
  .B1({ S10887 }),
  .B2({ S10867 }),
  .ZN({ S10888 })
);
OAI21_X1 #() 
OAI21_X1_551_ (
  .A({ S25957[397] }),
  .B1({ S10857 }),
  .B2({ S10859 }),
  .ZN({ S10889 })
);
NAND3_X1 #() 
NAND3_X1_1126_ (
  .A1({ S10889 }),
  .A2({ S10526 }),
  .A3({ S10888 }),
  .ZN({ S10890 })
);
NAND3_X1 #() 
NAND3_X1_1127_ (
  .A1({ S10883 }),
  .A2({ S10890 }),
  .A3({ S8507 }),
  .ZN({ S10891 })
);
NAND3_X1 #() 
NAND3_X1_1128_ (
  .A1({ S10891 }),
  .A2({ S10880 }),
  .A3({ S25957[399] }),
  .ZN({ S10892 })
);
NAND3_X1 #() 
NAND3_X1_1129_ (
  .A1({ S10878 }),
  .A2({ S10892 }),
  .A3({ S25957[500] }),
  .ZN({ S10893 })
);
NAND3_X1 #() 
NAND3_X1_1130_ (
  .A1({ S10893 }),
  .A2({ S10874 }),
  .A3({ S25957[468] }),
  .ZN({ S10894 })
);
NAND3_X1 #() 
NAND3_X1_1131_ (
  .A1({ S10872 }),
  .A2({ S10842 }),
  .A3({ S25957[500] }),
  .ZN({ S10896 })
);
NAND3_X1 #() 
NAND3_X1_1132_ (
  .A1({ S10878 }),
  .A2({ S10892 }),
  .A3({ S10815 }),
  .ZN({ S10897 })
);
NAND3_X1 #() 
NAND3_X1_1133_ (
  .A1({ S10897 }),
  .A2({ S10896 }),
  .A3({ S10813 }),
  .ZN({ S10898 })
);
NAND3_X1 #() 
NAND3_X1_1134_ (
  .A1({ S10894 }),
  .A2({ S10898 }),
  .A3({ S5128 }),
  .ZN({ S10899 })
);
NAND3_X1 #() 
NAND3_X1_1135_ (
  .A1({ S10897 }),
  .A2({ S10896 }),
  .A3({ S25957[468] }),
  .ZN({ S10900 })
);
NAND3_X1 #() 
NAND3_X1_1136_ (
  .A1({ S10893 }),
  .A2({ S10874 }),
  .A3({ S10813 }),
  .ZN({ S10901 })
);
NAND3_X1 #() 
NAND3_X1_1137_ (
  .A1({ S10900 }),
  .A2({ S10901 }),
  .A3({ S25957[532] }),
  .ZN({ S10902 })
);
AND2_X1 #() 
AND2_X1_62_ (
  .A1({ S10902 }),
  .A2({ S10899 }),
  .ZN({ S25957[276] })
);
NAND2_X1 #() 
NAND2_X1_993_ (
  .A1({ S8054 }),
  .A2({ S8030 }),
  .ZN({ S25957[499] })
);
NOR2_X1 #() 
NOR2_X1_234_ (
  .A1({ S25957[395] }),
  .A2({ S10584 }),
  .ZN({ S10903 })
);
NAND2_X1 #() 
NAND2_X1_994_ (
  .A1({ S10903 }),
  .A2({ S10545 }),
  .ZN({ S10905 })
);
NAND4_X1 #() 
NAND4_X1_133_ (
  .A1({ S25957[395] }),
  .A2({ S10569 }),
  .A3({ S25957[393] }),
  .A4({ S10538 }),
  .ZN({ S10906 })
);
NAND3_X1 #() 
NAND3_X1_1138_ (
  .A1({ S10905 }),
  .A2({ S10526 }),
  .A3({ S10906 }),
  .ZN({ S10907 })
);
NAND2_X1 #() 
NAND2_X1_995_ (
  .A1({ S10571 }),
  .A2({ S25957[395] }),
  .ZN({ S10908 })
);
NAND2_X1 #() 
NAND2_X1_996_ (
  .A1({ S10675 }),
  .A2({ S21 }),
  .ZN({ S10909 })
);
OAI211_X1 #() 
OAI211_X1_349_ (
  .A({ S10909 }),
  .B({ S25957[396] }),
  .C1({ S10753 }),
  .C2({ S10908 }),
  .ZN({ S10910 })
);
NAND3_X1 #() 
NAND3_X1_1139_ (
  .A1({ S10910 }),
  .A2({ S10907 }),
  .A3({ S25957[397] }),
  .ZN({ S10911 })
);
AOI22_X1 #() 
AOI22_X1_122_ (
  .A1({ S10702 }),
  .A2({ S10612 }),
  .B1({ S10576 }),
  .B2({ S25957[395] }),
  .ZN({ S10912 })
);
AOI21_X1 #() 
AOI21_X1_606_ (
  .A({ S25957[397] }),
  .B1({ S10820 }),
  .B2({ S10711 }),
  .ZN({ S10913 })
);
OAI21_X1 #() 
OAI21_X1_552_ (
  .A({ S10913 }),
  .B1({ S10912 }),
  .B2({ S10526 }),
  .ZN({ S10914 })
);
NAND2_X1 #() 
NAND2_X1_997_ (
  .A1({ S10538 }),
  .A2({ S10535 }),
  .ZN({ S10916 })
);
NOR3_X1 #() 
NOR3_X1_32_ (
  .A1({ S10704 }),
  .A2({ S10916 }),
  .A3({ S21 }),
  .ZN({ S10917 })
);
NOR2_X1 #() 
NOR2_X1_235_ (
  .A1({ S10661 }),
  .A2({ S10729 }),
  .ZN({ S10918 })
);
OAI21_X1 #() 
OAI21_X1_553_ (
  .A({ S10526 }),
  .B1({ S10917 }),
  .B2({ S10918 }),
  .ZN({ S10919 })
);
NAND3_X1 #() 
NAND3_X1_1140_ (
  .A1({ S10886 }),
  .A2({ S21 }),
  .A3({ S10547 }),
  .ZN({ S10920 })
);
AOI21_X1 #() 
AOI21_X1_607_ (
  .A({ S10526 }),
  .B1({ S10663 }),
  .B2({ S25957[395] }),
  .ZN({ S10921 })
);
AOI21_X1 #() 
AOI21_X1_608_ (
  .A({ S10559 }),
  .B1({ S10921 }),
  .B2({ S10920 }),
  .ZN({ S10922 })
);
AOI21_X1 #() 
AOI21_X1_609_ (
  .A({ S8507 }),
  .B1({ S10919 }),
  .B2({ S10922 }),
  .ZN({ S10923 })
);
NAND2_X1 #() 
NAND2_X1_998_ (
  .A1({ S10711 }),
  .A2({ S21 }),
  .ZN({ S10924 })
);
NAND4_X1 #() 
NAND4_X1_134_ (
  .A1({ S25957[395] }),
  .A2({ S25957[394] }),
  .A3({ S10547 }),
  .A4({ S10546 }),
  .ZN({ S10925 })
);
NAND2_X1 #() 
NAND2_X1_999_ (
  .A1({ S10924 }),
  .A2({ S10925 }),
  .ZN({ S10927 })
);
OAI21_X1 #() 
OAI21_X1_554_ (
  .A({ S10526 }),
  .B1({ S10927 }),
  .B2({ S10542 }),
  .ZN({ S10928 })
);
AOI21_X1 #() 
AOI21_X1_610_ (
  .A({ S10526 }),
  .B1({ S10548 }),
  .B2({ S25957[395] }),
  .ZN({ S10929 })
);
AOI21_X1 #() 
AOI21_X1_611_ (
  .A({ S25957[397] }),
  .B1({ S10929 }),
  .B2({ S10849 }),
  .ZN({ S10930 })
);
AOI21_X1 #() 
AOI21_X1_612_ (
  .A({ S25957[398] }),
  .B1({ S10928 }),
  .B2({ S10930 }),
  .ZN({ S10931 })
);
AOI22_X1 #() 
AOI22_X1_123_ (
  .A1({ S10931 }),
  .A2({ S10911 }),
  .B1({ S10923 }),
  .B2({ S10914 }),
  .ZN({ S10932 })
);
OAI21_X1 #() 
OAI21_X1_555_ (
  .A({ S31 }),
  .B1({ S10527 }),
  .B2({ S25957[394] }),
  .ZN({ S10933 })
);
OAI211_X1 #() 
OAI211_X1_350_ (
  .A({ S10773 }),
  .B({ S25957[396] }),
  .C1({ S21 }),
  .C2({ S10933 }),
  .ZN({ S10934 })
);
NAND3_X1 #() 
NAND3_X1_1141_ (
  .A1({ S10734 }),
  .A2({ S10578 }),
  .A3({ S10526 }),
  .ZN({ S10935 })
);
OAI211_X1 #() 
OAI211_X1_351_ (
  .A({ S10934 }),
  .B({ S10559 }),
  .C1({ S10935 }),
  .C2({ S10613 }),
  .ZN({ S10936 })
);
AND2_X1 #() 
AND2_X1_63_ (
  .A1({ S10568 }),
  .A2({ S21 }),
  .ZN({ S10938 })
);
OAI21_X1 #() 
OAI21_X1_556_ (
  .A({ S10788 }),
  .B1({ S10938 }),
  .B2({ S10699 }),
  .ZN({ S10939 })
);
OAI211_X1 #() 
OAI211_X1_352_ (
  .A({ S10908 }),
  .B({ S25957[396] }),
  .C1({ S25957[395] }),
  .C2({ S10633 }),
  .ZN({ S10940 })
);
NAND3_X1 #() 
NAND3_X1_1142_ (
  .A1({ S10940 }),
  .A2({ S10939 }),
  .A3({ S25957[397] }),
  .ZN({ S10941 })
);
NAND3_X1 #() 
NAND3_X1_1143_ (
  .A1({ S10936 }),
  .A2({ S10941 }),
  .A3({ S8507 }),
  .ZN({ S10942 })
);
NAND3_X1 #() 
NAND3_X1_1144_ (
  .A1({ S10568 }),
  .A2({ S21 }),
  .A3({ S10547 }),
  .ZN({ S10943 })
);
NAND3_X1 #() 
NAND3_X1_1145_ (
  .A1({ S10943 }),
  .A2({ S10683 }),
  .A3({ S10526 }),
  .ZN({ S10944 })
);
OAI211_X1 #() 
OAI211_X1_353_ (
  .A({ S25957[397] }),
  .B({ S10944 }),
  .C1({ S10639 }),
  .C2({ S10677 }),
  .ZN({ S10945 })
);
NAND2_X1 #() 
NAND2_X1_1000_ (
  .A1({ S10681 }),
  .A2({ S10669 }),
  .ZN({ S10946 })
);
NAND4_X1 #() 
NAND4_X1_135_ (
  .A1({ S10946 }),
  .A2({ S10858 }),
  .A3({ S10578 }),
  .A4({ S10526 }),
  .ZN({ S10947 })
);
NAND3_X1 #() 
NAND3_X1_1146_ (
  .A1({ S21 }),
  .A2({ S10527 }),
  .A3({ S10513 }),
  .ZN({ S10949 })
);
AOI21_X1 #() 
AOI21_X1_613_ (
  .A({ S25957[397] }),
  .B1({ S25957[396] }),
  .B2({ S10949 }),
  .ZN({ S10950 })
);
NAND2_X1 #() 
NAND2_X1_1001_ (
  .A1({ S10947 }),
  .A2({ S10950 }),
  .ZN({ S10951 })
);
NAND3_X1 #() 
NAND3_X1_1147_ (
  .A1({ S10945 }),
  .A2({ S10951 }),
  .A3({ S25957[398] }),
  .ZN({ S10952 })
);
NAND3_X1 #() 
NAND3_X1_1148_ (
  .A1({ S10952 }),
  .A2({ S10598 }),
  .A3({ S10942 }),
  .ZN({ S10953 })
);
OAI211_X1 #() 
OAI211_X1_354_ (
  .A({ S10953 }),
  .B({ S25957[499] }),
  .C1({ S10932 }),
  .C2({ S10598 }),
  .ZN({ S10954 })
);
INV_X1 #() 
INV_X1_328_ (
  .A({ S25957[499] }),
  .ZN({ S10955 })
);
NAND2_X1 #() 
NAND2_X1_1002_ (
  .A1({ S10928 }),
  .A2({ S10930 }),
  .ZN({ S10956 })
);
AOI21_X1 #() 
AOI21_X1_614_ (
  .A({ S10598 }),
  .B1({ S10956 }),
  .B2({ S10911 }),
  .ZN({ S10957 })
);
AND3_X1 #() 
AND3_X1_45_ (
  .A1({ S10936 }),
  .A2({ S10598 }),
  .A3({ S10941 }),
  .ZN({ S10958 })
);
OAI21_X1 #() 
OAI21_X1_557_ (
  .A({ S8507 }),
  .B1({ S10957 }),
  .B2({ S10958 }),
  .ZN({ S10959 })
);
NOR2_X1 #() 
NOR2_X1_236_ (
  .A1({ S25957[395] }),
  .A2({ S10579 }),
  .ZN({ S10960 })
);
AOI22_X1 #() 
AOI22_X1_124_ (
  .A1({ S10546 }),
  .A2({ S10513 }),
  .B1({ S25957[394] }),
  .B2({ S25957[393] }),
  .ZN({ S10961 })
);
AOI22_X1 #() 
AOI22_X1_125_ (
  .A1({ S10961 }),
  .A2({ S25957[395] }),
  .B1({ S10960 }),
  .B2({ S10718 }),
  .ZN({ S10962 })
);
NAND3_X1 #() 
NAND3_X1_1149_ (
  .A1({ S10920 }),
  .A2({ S25957[396] }),
  .A3({ S10835 }),
  .ZN({ S10963 })
);
OAI211_X1 #() 
OAI211_X1_355_ (
  .A({ S10963 }),
  .B({ S25957[397] }),
  .C1({ S10962 }),
  .C2({ S25957[396] }),
  .ZN({ S10964 })
);
AOI21_X1 #() 
AOI21_X1_615_ (
  .A({ S10598 }),
  .B1({ S10964 }),
  .B2({ S10914 }),
  .ZN({ S10965 })
);
NAND2_X1 #() 
NAND2_X1_1003_ (
  .A1({ S10669 }),
  .A2({ S10513 }),
  .ZN({ S10966 })
);
AOI22_X1 #() 
AOI22_X1_126_ (
  .A1({ S10966 }),
  .A2({ S25957[395] }),
  .B1({ S10681 }),
  .B2({ S10669 }),
  .ZN({ S10967 })
);
INV_X1 #() 
INV_X1_329_ (
  .A({ S10949 }),
  .ZN({ S10968 })
);
AOI21_X1 #() 
AOI21_X1_616_ (
  .A({ S25957[397] }),
  .B1({ S10968 }),
  .B2({ S25957[396] }),
  .ZN({ S10970 })
);
OAI21_X1 #() 
OAI21_X1_558_ (
  .A({ S10970 }),
  .B1({ S10967 }),
  .B2({ S25957[396] }),
  .ZN({ S10971 })
);
AOI21_X1 #() 
AOI21_X1_617_ (
  .A({ S25957[395] }),
  .B1({ S25957[393] }),
  .B2({ S10589 }),
  .ZN({ S10972 })
);
AOI22_X1 #() 
AOI22_X1_127_ (
  .A1({ S10972 }),
  .A2({ S10545 }),
  .B1({ S25957[395] }),
  .B2({ S10675 }),
  .ZN({ S10973 })
);
NAND2_X1 #() 
NAND2_X1_1004_ (
  .A1({ S10943 }),
  .A2({ S10683 }),
  .ZN({ S10974 })
);
NAND2_X1 #() 
NAND2_X1_1005_ (
  .A1({ S10974 }),
  .A2({ S10526 }),
  .ZN({ S10975 })
);
OAI211_X1 #() 
OAI211_X1_356_ (
  .A({ S25957[397] }),
  .B({ S10975 }),
  .C1({ S10973 }),
  .C2({ S10526 }),
  .ZN({ S10976 })
);
AOI21_X1 #() 
AOI21_X1_618_ (
  .A({ S25957[399] }),
  .B1({ S10976 }),
  .B2({ S10971 }),
  .ZN({ S10977 })
);
OAI21_X1 #() 
OAI21_X1_559_ (
  .A({ S25957[398] }),
  .B1({ S10977 }),
  .B2({ S10965 }),
  .ZN({ S10978 })
);
NAND3_X1 #() 
NAND3_X1_1150_ (
  .A1({ S10959 }),
  .A2({ S10978 }),
  .A3({ S10955 }),
  .ZN({ S10979 })
);
AOI21_X1 #() 
AOI21_X1_619_ (
  .A({ S25957[563] }),
  .B1({ S10979 }),
  .B2({ S10954 }),
  .ZN({ S10981 })
);
OAI211_X1 #() 
OAI211_X1_357_ (
  .A({ S10953 }),
  .B({ S10955 }),
  .C1({ S10932 }),
  .C2({ S10598 }),
  .ZN({ S10982 })
);
NAND3_X1 #() 
NAND3_X1_1151_ (
  .A1({ S10959 }),
  .A2({ S10978 }),
  .A3({ S25957[499] }),
  .ZN({ S10983 })
);
AOI21_X1 #() 
AOI21_X1_620_ (
  .A({ S7964 }),
  .B1({ S10983 }),
  .B2({ S10982 }),
  .ZN({ S10984 })
);
OAI21_X1 #() 
OAI21_X1_560_ (
  .A({ S18 }),
  .B1({ S10981 }),
  .B2({ S10984 }),
  .ZN({ S10985 })
);
NAND3_X1 #() 
NAND3_X1_1152_ (
  .A1({ S10983 }),
  .A2({ S10982 }),
  .A3({ S7964 }),
  .ZN({ S10986 })
);
NAND3_X1 #() 
NAND3_X1_1153_ (
  .A1({ S10979 }),
  .A2({ S10954 }),
  .A3({ S25957[563] }),
  .ZN({ S10987 })
);
NAND3_X1 #() 
NAND3_X1_1154_ (
  .A1({ S10986 }),
  .A2({ S10987 }),
  .A3({ S25957[403] }),
  .ZN({ S10988 })
);
NAND2_X1 #() 
NAND2_X1_1006_ (
  .A1({ S10985 }),
  .A2({ S10988 }),
  .ZN({ S32 })
);
OAI21_X1 #() 
OAI21_X1_561_ (
  .A({ S25957[403] }),
  .B1({ S10981 }),
  .B2({ S10984 }),
  .ZN({ S10989 })
);
NAND3_X1 #() 
NAND3_X1_1155_ (
  .A1({ S10986 }),
  .A2({ S10987 }),
  .A3({ S18 }),
  .ZN({ S10991 })
);
NAND2_X1 #() 
NAND2_X1_1007_ (
  .A1({ S10989 }),
  .A2({ S10991 }),
  .ZN({ S25957[275] })
);
NOR2_X1 #() 
NOR2_X1_237_ (
  .A1({ S5283 }),
  .A2({ S5284 }),
  .ZN({ S10992 })
);
NOR2_X1 #() 
NOR2_X1_238_ (
  .A1({ S8121 }),
  .A2({ S8122 }),
  .ZN({ S25957[464] })
);
INV_X1 #() 
INV_X1_330_ (
  .A({ S25957[464] }),
  .ZN({ S10993 })
);
NOR2_X1 #() 
NOR2_X1_239_ (
  .A1({ S10993 }),
  .A2({ S10992 }),
  .ZN({ S10994 })
);
INV_X1 #() 
INV_X1_331_ (
  .A({ S10992 }),
  .ZN({ S25957[560] })
);
NOR2_X1 #() 
NOR2_X1_240_ (
  .A1({ S25957[464] }),
  .A2({ S25957[560] }),
  .ZN({ S10995 })
);
NOR2_X1 #() 
NOR2_X1_241_ (
  .A1({ S10994 }),
  .A2({ S10995 }),
  .ZN({ S25957[432] })
);
INV_X1 #() 
INV_X1_332_ (
  .A({ S25957[432] }),
  .ZN({ S10996 })
);
NAND2_X1 #() 
NAND2_X1_1008_ (
  .A1({ S5279 }),
  .A2({ S5278 }),
  .ZN({ S25957[624] })
);
XNOR2_X1 #() 
XNOR2_X1_35_ (
  .A({ S25957[624] }),
  .B({ S8125 }),
  .ZN({ S25957[592] })
);
NAND4_X1 #() 
NAND4_X1_136_ (
  .A1({ S10568 }),
  .A2({ S25957[395] }),
  .A3({ S10546 }),
  .A4({ S10547 }),
  .ZN({ S10998 })
);
OAI211_X1 #() 
OAI211_X1_358_ (
  .A({ S10526 }),
  .B({ S10998 }),
  .C1({ S10690 }),
  .C2({ S10580 }),
  .ZN({ S10999 })
);
NAND3_X1 #() 
NAND3_X1_1156_ (
  .A1({ S10518 }),
  .A2({ S10569 }),
  .A3({ S10538 }),
  .ZN({ S11000 })
);
NAND3_X1 #() 
NAND3_X1_1157_ (
  .A1({ S10784 }),
  .A2({ S11000 }),
  .A3({ S10526 }),
  .ZN({ S11001 })
);
AOI21_X1 #() 
AOI21_X1_621_ (
  .A({ S10559 }),
  .B1({ S10921 }),
  .B2({ S10777 }),
  .ZN({ S11002 })
);
OAI21_X1 #() 
OAI21_X1_562_ (
  .A({ S21 }),
  .B1({ S10633 }),
  .B2({ S10584 }),
  .ZN({ S11003 })
);
AOI21_X1 #() 
AOI21_X1_622_ (
  .A({ S25957[397] }),
  .B1({ S11003 }),
  .B2({ S10929 }),
  .ZN({ S11004 })
);
AOI22_X1 #() 
AOI22_X1_128_ (
  .A1({ S11004 }),
  .A2({ S10999 }),
  .B1({ S11002 }),
  .B2({ S11001 }),
  .ZN({ S11005 })
);
OAI21_X1 #() 
OAI21_X1_563_ (
  .A({ S25957[396] }),
  .B1({ S10660 }),
  .B2({ S10776 }),
  .ZN({ S11007 })
);
AOI22_X1 #() 
AOI22_X1_129_ (
  .A1({ S10825 }),
  .A2({ S10609 }),
  .B1({ S21 }),
  .B2({ S10731 }),
  .ZN({ S11008 })
);
OAI211_X1 #() 
OAI211_X1_359_ (
  .A({ S10559 }),
  .B({ S11007 }),
  .C1({ S11008 }),
  .C2({ S25957[396] }),
  .ZN({ S11009 })
);
AOI21_X1 #() 
AOI21_X1_623_ (
  .A({ S21 }),
  .B1({ S10545 }),
  .B2({ S10590 }),
  .ZN({ S11010 })
);
NAND3_X1 #() 
NAND3_X1_1158_ (
  .A1({ S10866 }),
  .A2({ S25957[396] }),
  .A3({ S10627 }),
  .ZN({ S11011 })
);
NAND2_X1 #() 
NAND2_X1_1009_ (
  .A1({ S10575 }),
  .A2({ S21 }),
  .ZN({ S11012 })
);
AOI21_X1 #() 
AOI21_X1_624_ (
  .A({ S25957[396] }),
  .B1({ S25957[395] }),
  .B2({ S10584 }),
  .ZN({ S11013 })
);
NAND3_X1 #() 
NAND3_X1_1159_ (
  .A1({ S11013 }),
  .A2({ S10667 }),
  .A3({ S11012 }),
  .ZN({ S11014 })
);
OAI211_X1 #() 
OAI211_X1_360_ (
  .A({ S11014 }),
  .B({ S25957[397] }),
  .C1({ S11010 }),
  .C2({ S11011 }),
  .ZN({ S11015 })
);
NAND3_X1 #() 
NAND3_X1_1160_ (
  .A1({ S11015 }),
  .A2({ S11009 }),
  .A3({ S25957[398] }),
  .ZN({ S11016 })
);
OAI211_X1 #() 
OAI211_X1_361_ (
  .A({ S11016 }),
  .B({ S10598 }),
  .C1({ S11005 }),
  .C2({ S25957[398] }),
  .ZN({ S11018 })
);
OAI21_X1 #() 
OAI21_X1_564_ (
  .A({ S21 }),
  .B1({ S10753 }),
  .B2({ S10550 }),
  .ZN({ S11019 })
);
AOI21_X1 #() 
AOI21_X1_625_ (
  .A({ S10526 }),
  .B1({ S10823 }),
  .B2({ S25957[395] }),
  .ZN({ S11020 })
);
AOI21_X1 #() 
AOI21_X1_626_ (
  .A({ S25957[396] }),
  .B1({ S10628 }),
  .B2({ S10669 }),
  .ZN({ S11021 })
);
AOI22_X1 #() 
AOI22_X1_130_ (
  .A1({ S11021 }),
  .A2({ S11019 }),
  .B1({ S10572 }),
  .B2({ S11020 }),
  .ZN({ S11022 })
);
AOI21_X1 #() 
AOI21_X1_627_ (
  .A({ S10526 }),
  .B1({ S10612 }),
  .B2({ S25957[395] }),
  .ZN({ S11023 })
);
NAND2_X1 #() 
NAND2_X1_1010_ (
  .A1({ S11023 }),
  .A2({ S10853 }),
  .ZN({ S11024 })
);
NAND3_X1 #() 
NAND3_X1_1161_ (
  .A1({ S10767 }),
  .A2({ S10559 }),
  .A3({ S11024 }),
  .ZN({ S11025 })
);
OAI211_X1 #() 
OAI211_X1_362_ (
  .A({ S11025 }),
  .B({ S25957[398] }),
  .C1({ S10559 }),
  .C2({ S11022 }),
  .ZN({ S11026 })
);
NAND2_X1 #() 
NAND2_X1_1011_ (
  .A1({ S25957[395] }),
  .A2({ S10535 }),
  .ZN({ S11027 })
);
OAI211_X1 #() 
OAI211_X1_363_ (
  .A({ S11027 }),
  .B({ S25957[396] }),
  .C1({ S10753 }),
  .C2({ S25957[395] }),
  .ZN({ S11029 })
);
NAND3_X1 #() 
NAND3_X1_1162_ (
  .A1({ S10865 }),
  .A2({ S10683 }),
  .A3({ S10526 }),
  .ZN({ S11030 })
);
AND2_X1 #() 
AND2_X1_64_ (
  .A1({ S11029 }),
  .A2({ S11030 }),
  .ZN({ S11031 })
);
NAND3_X1 #() 
NAND3_X1_1163_ (
  .A1({ S10858 }),
  .A2({ S10740 }),
  .A3({ S10843 }),
  .ZN({ S11032 })
);
NAND2_X1 #() 
NAND2_X1_1012_ (
  .A1({ S11032 }),
  .A2({ S10526 }),
  .ZN({ S11033 })
);
NAND3_X1 #() 
NAND3_X1_1164_ (
  .A1({ S10585 }),
  .A2({ S21 }),
  .A3({ S10538 }),
  .ZN({ S11034 })
);
AOI21_X1 #() 
AOI21_X1_628_ (
  .A({ S10526 }),
  .B1({ S10699 }),
  .B2({ S10528 }),
  .ZN({ S11035 })
);
AOI21_X1 #() 
AOI21_X1_629_ (
  .A({ S10559 }),
  .B1({ S11034 }),
  .B2({ S11035 }),
  .ZN({ S11036 })
);
NAND2_X1 #() 
NAND2_X1_1013_ (
  .A1({ S11033 }),
  .A2({ S11036 }),
  .ZN({ S11037 })
);
OAI211_X1 #() 
OAI211_X1_364_ (
  .A({ S11037 }),
  .B({ S8507 }),
  .C1({ S11031 }),
  .C2({ S25957[397] }),
  .ZN({ S11038 })
);
NAND3_X1 #() 
NAND3_X1_1165_ (
  .A1({ S11026 }),
  .A2({ S25957[399] }),
  .A3({ S11038 }),
  .ZN({ S11040 })
);
AOI21_X1 #() 
AOI21_X1_630_ (
  .A({ S25957[592] }),
  .B1({ S11040 }),
  .B2({ S11018 }),
  .ZN({ S11041 })
);
INV_X1 #() 
INV_X1_333_ (
  .A({ S25957[592] }),
  .ZN({ S11042 })
);
AOI22_X1 #() 
AOI22_X1_131_ (
  .A1({ S10526 }),
  .A2({ S10766 }),
  .B1({ S11023 }),
  .B2({ S10853 }),
  .ZN({ S11043 })
);
AOI22_X1 #() 
AOI22_X1_132_ (
  .A1({ S10528 }),
  .A2({ S10516 }),
  .B1({ S9040 }),
  .B2({ S9037 }),
  .ZN({ S11044 })
);
OAI211_X1 #() 
OAI211_X1_365_ (
  .A({ S25957[396] }),
  .B({ S10733 }),
  .C1({ S10843 }),
  .C2({ S11044 }),
  .ZN({ S11045 })
);
NAND2_X1 #() 
NAND2_X1_1014_ (
  .A1({ S25957[395] }),
  .A2({ S10513 }),
  .ZN({ S11046 })
);
OAI21_X1 #() 
OAI21_X1_565_ (
  .A({ S10526 }),
  .B1({ S11046 }),
  .B2({ S10580 }),
  .ZN({ S11047 })
);
OAI211_X1 #() 
OAI211_X1_366_ (
  .A({ S11045 }),
  .B({ S25957[397] }),
  .C1({ S11047 }),
  .C2({ S10537 }),
  .ZN({ S11048 })
);
OAI211_X1 #() 
OAI211_X1_367_ (
  .A({ S25957[398] }),
  .B({ S11048 }),
  .C1({ S11043 }),
  .C2({ S25957[397] }),
  .ZN({ S11049 })
);
AOI22_X1 #() 
AOI22_X1_133_ (
  .A1({ S11032 }),
  .A2({ S10526 }),
  .B1({ S11034 }),
  .B2({ S11035 }),
  .ZN({ S11051 })
);
NAND3_X1 #() 
NAND3_X1_1166_ (
  .A1({ S11029 }),
  .A2({ S11030 }),
  .A3({ S10559 }),
  .ZN({ S11052 })
);
OAI211_X1 #() 
OAI211_X1_368_ (
  .A({ S11052 }),
  .B({ S8507 }),
  .C1({ S11051 }),
  .C2({ S10559 }),
  .ZN({ S11053 })
);
NAND3_X1 #() 
NAND3_X1_1167_ (
  .A1({ S11049 }),
  .A2({ S11053 }),
  .A3({ S25957[399] }),
  .ZN({ S11054 })
);
NAND3_X1 #() 
NAND3_X1_1168_ (
  .A1({ S10777 }),
  .A2({ S25957[396] }),
  .A3({ S10835 }),
  .ZN({ S11055 })
);
NAND3_X1 #() 
NAND3_X1_1169_ (
  .A1({ S11001 }),
  .A2({ S25957[397] }),
  .A3({ S11055 }),
  .ZN({ S11056 })
);
NAND2_X1 #() 
NAND2_X1_1015_ (
  .A1({ S11003 }),
  .A2({ S10929 }),
  .ZN({ S11057 })
);
NAND3_X1 #() 
NAND3_X1_1170_ (
  .A1({ S11057 }),
  .A2({ S10559 }),
  .A3({ S10999 }),
  .ZN({ S11058 })
);
NAND3_X1 #() 
NAND3_X1_1171_ (
  .A1({ S11058 }),
  .A2({ S11056 }),
  .A3({ S8507 }),
  .ZN({ S11059 })
);
NAND2_X1 #() 
NAND2_X1_1016_ (
  .A1({ S10545 }),
  .A2({ S10590 }),
  .ZN({ S11060 })
);
AOI21_X1 #() 
AOI21_X1_631_ (
  .A({ S11011 }),
  .B1({ S11060 }),
  .B2({ S25957[395] }),
  .ZN({ S11062 })
);
NAND3_X1 #() 
NAND3_X1_1172_ (
  .A1({ S10886 }),
  .A2({ S10885 }),
  .A3({ S25957[395] }),
  .ZN({ S11063 })
);
NAND3_X1 #() 
NAND3_X1_1173_ (
  .A1({ S21 }),
  .A2({ S10528 }),
  .A3({ S10529 }),
  .ZN({ S11064 })
);
AOI21_X1 #() 
AOI21_X1_632_ (
  .A({ S25957[396] }),
  .B1({ S11063 }),
  .B2({ S11064 }),
  .ZN({ S11065 })
);
OAI21_X1 #() 
OAI21_X1_566_ (
  .A({ S25957[397] }),
  .B1({ S11062 }),
  .B2({ S11065 }),
  .ZN({ S11066 })
);
OAI211_X1 #() 
OAI211_X1_369_ (
  .A({ S10732 }),
  .B({ S10526 }),
  .C1({ S10764 }),
  .C2({ S10763 }),
  .ZN({ S11067 })
);
OAI21_X1 #() 
OAI21_X1_567_ (
  .A({ S25957[396] }),
  .B1({ S21 }),
  .B2({ S25957[392] }),
  .ZN({ S11068 })
);
OAI211_X1 #() 
OAI211_X1_370_ (
  .A({ S11067 }),
  .B({ S10559 }),
  .C1({ S10660 }),
  .C2({ S11068 }),
  .ZN({ S11069 })
);
NAND3_X1 #() 
NAND3_X1_1174_ (
  .A1({ S11066 }),
  .A2({ S25957[398] }),
  .A3({ S11069 }),
  .ZN({ S11070 })
);
NAND3_X1 #() 
NAND3_X1_1175_ (
  .A1({ S11070 }),
  .A2({ S11059 }),
  .A3({ S10598 }),
  .ZN({ S11071 })
);
AOI21_X1 #() 
AOI21_X1_633_ (
  .A({ S11042 }),
  .B1({ S11071 }),
  .B2({ S11054 }),
  .ZN({ S11073 })
);
OAI21_X1 #() 
OAI21_X1_568_ (
  .A({ S10996 }),
  .B1({ S11041 }),
  .B2({ S11073 }),
  .ZN({ S11074 })
);
NAND3_X1 #() 
NAND3_X1_1176_ (
  .A1({ S11071 }),
  .A2({ S11054 }),
  .A3({ S11042 }),
  .ZN({ S11075 })
);
NAND3_X1 #() 
NAND3_X1_1177_ (
  .A1({ S11040 }),
  .A2({ S11018 }),
  .A3({ S25957[592] }),
  .ZN({ S11076 })
);
NAND3_X1 #() 
NAND3_X1_1178_ (
  .A1({ S11076 }),
  .A2({ S25957[432] }),
  .A3({ S11075 }),
  .ZN({ S11077 })
);
NAND3_X1 #() 
NAND3_X1_1179_ (
  .A1({ S11074 }),
  .A2({ S25957[400] }),
  .A3({ S11077 }),
  .ZN({ S11078 })
);
NAND3_X1 #() 
NAND3_X1_1180_ (
  .A1({ S8127 }),
  .A2({ S25957[656] }),
  .A3({ S8120 }),
  .ZN({ S11079 })
);
OAI21_X1 #() 
OAI21_X1_569_ (
  .A({ S5282 }),
  .B1({ S8121 }),
  .B2({ S8122 }),
  .ZN({ S11080 })
);
NAND2_X1 #() 
NAND2_X1_1017_ (
  .A1({ S11080 }),
  .A2({ S11079 }),
  .ZN({ S11081 })
);
OAI21_X1 #() 
OAI21_X1_570_ (
  .A({ S25957[432] }),
  .B1({ S11041 }),
  .B2({ S11073 }),
  .ZN({ S11082 })
);
NAND3_X1 #() 
NAND3_X1_1181_ (
  .A1({ S11076 }),
  .A2({ S10996 }),
  .A3({ S11075 }),
  .ZN({ S11084 })
);
NAND3_X1 #() 
NAND3_X1_1182_ (
  .A1({ S11082 }),
  .A2({ S11081 }),
  .A3({ S11084 }),
  .ZN({ S11085 })
);
NAND2_X1 #() 
NAND2_X1_1018_ (
  .A1({ S11078 }),
  .A2({ S11085 }),
  .ZN({ S25957[272] })
);
NOR2_X1 #() 
NOR2_X1_242_ (
  .A1({ S8193 }),
  .A2({ S8198 }),
  .ZN({ S11086 })
);
NAND2_X1 #() 
NAND2_X1_1019_ (
  .A1({ S8129 }),
  .A2({ S8131 }),
  .ZN({ S11087 })
);
NOR3_X1 #() 
NOR3_X1_33_ (
  .A1({ S10611 }),
  .A2({ S10887 }),
  .A3({ S25957[396] }),
  .ZN({ S11088 })
);
AOI21_X1 #() 
AOI21_X1_634_ (
  .A({ S25957[395] }),
  .B1({ S10885 }),
  .B2({ S10535 }),
  .ZN({ S11089 })
);
OAI21_X1 #() 
OAI21_X1_571_ (
  .A({ S10559 }),
  .B1({ S11089 }),
  .B2({ S10687 }),
  .ZN({ S11090 })
);
AOI21_X1 #() 
AOI21_X1_635_ (
  .A({ S21 }),
  .B1({ S10612 }),
  .B2({ S10575 }),
  .ZN({ S11091 })
);
NAND3_X1 #() 
NAND3_X1_1183_ (
  .A1({ S25957[395] }),
  .A2({ S10569 }),
  .A3({ S10541 }),
  .ZN({ S11092 })
);
NAND3_X1 #() 
NAND3_X1_1184_ (
  .A1({ S11092 }),
  .A2({ S10943 }),
  .A3({ S10526 }),
  .ZN({ S11094 })
);
OAI211_X1 #() 
OAI211_X1_371_ (
  .A({ S11094 }),
  .B({ S25957[397] }),
  .C1({ S11091 }),
  .C2({ S10601 }),
  .ZN({ S11095 })
);
OAI211_X1 #() 
OAI211_X1_372_ (
  .A({ S11095 }),
  .B({ S8507 }),
  .C1({ S11088 }),
  .C2({ S11090 }),
  .ZN({ S11096 })
);
NAND3_X1 #() 
NAND3_X1_1185_ (
  .A1({ S21 }),
  .A2({ S10528 }),
  .A3({ S10535 }),
  .ZN({ S11097 })
);
AND3_X1 #() 
AND3_X1_46_ (
  .A1({ S10774 }),
  .A2({ S11097 }),
  .A3({ S25957[396] }),
  .ZN({ S11098 })
);
NAND3_X1 #() 
NAND3_X1_1186_ (
  .A1({ S25957[395] }),
  .A2({ S10527 }),
  .A3({ S10538 }),
  .ZN({ S11099 })
);
OAI211_X1 #() 
OAI211_X1_373_ (
  .A({ S11099 }),
  .B({ S10526 }),
  .C1({ S10949 }),
  .C2({ S10750 }),
  .ZN({ S11100 })
);
NAND2_X1 #() 
NAND2_X1_1020_ (
  .A1({ S11100 }),
  .A2({ S10559 }),
  .ZN({ S11101 })
);
NAND4_X1 #() 
NAND4_X1_137_ (
  .A1({ S10527 }),
  .A2({ S10535 }),
  .A3({ S8759 }),
  .A4({ S8762 }),
  .ZN({ S11102 })
);
NAND3_X1 #() 
NAND3_X1_1187_ (
  .A1({ S10605 }),
  .A2({ S11102 }),
  .A3({ S25957[396] }),
  .ZN({ S11103 })
);
OAI21_X1 #() 
OAI21_X1_572_ (
  .A({ S10526 }),
  .B1({ S10636 }),
  .B2({ S25957[395] }),
  .ZN({ S11105 })
);
OAI211_X1 #() 
OAI211_X1_374_ (
  .A({ S25957[397] }),
  .B({ S11103 }),
  .C1({ S11010 }),
  .C2({ S11105 }),
  .ZN({ S11106 })
);
OAI211_X1 #() 
OAI211_X1_375_ (
  .A({ S11106 }),
  .B({ S25957[398] }),
  .C1({ S11098 }),
  .C2({ S11101 }),
  .ZN({ S11107 })
);
NAND3_X1 #() 
NAND3_X1_1188_ (
  .A1({ S11096 }),
  .A2({ S11107 }),
  .A3({ S25957[399] }),
  .ZN({ S11108 })
);
AOI21_X1 #() 
AOI21_X1_636_ (
  .A({ S10526 }),
  .B1({ S10906 }),
  .B2({ S10845 }),
  .ZN({ S11109 })
);
OAI21_X1 #() 
OAI21_X1_573_ (
  .A({ S25957[397] }),
  .B1({ S11109 }),
  .B2({ S10617 }),
  .ZN({ S11110 })
);
NAND2_X1 #() 
NAND2_X1_1021_ (
  .A1({ S10946 }),
  .A2({ S11013 }),
  .ZN({ S11111 })
);
NAND4_X1 #() 
NAND4_X1_138_ (
  .A1({ S10578 }),
  .A2({ S10849 }),
  .A3({ S25957[396] }),
  .A4({ S10517 }),
  .ZN({ S11112 })
);
NAND3_X1 #() 
NAND3_X1_1189_ (
  .A1({ S11111 }),
  .A2({ S10559 }),
  .A3({ S11112 }),
  .ZN({ S11113 })
);
NAND3_X1 #() 
NAND3_X1_1190_ (
  .A1({ S11110 }),
  .A2({ S11113 }),
  .A3({ S8507 }),
  .ZN({ S11114 })
);
AOI21_X1 #() 
AOI21_X1_637_ (
  .A({ S10570 }),
  .B1({ S30 }),
  .B2({ S10529 }),
  .ZN({ S11116 })
);
OAI21_X1 #() 
OAI21_X1_574_ (
  .A({ S25957[396] }),
  .B1({ S11116 }),
  .B2({ S21 }),
  .ZN({ S11117 })
);
NAND4_X1 #() 
NAND4_X1_139_ (
  .A1({ S10530 }),
  .A2({ S10526 }),
  .A3({ S10517 }),
  .A4({ S10513 }),
  .ZN({ S11118 })
);
AND3_X1 #() 
AND3_X1_47_ (
  .A1({ S10551 }),
  .A2({ S10571 }),
  .A3({ S25957[396] }),
  .ZN({ S11119 })
);
AOI21_X1 #() 
AOI21_X1_638_ (
  .A({ S11119 }),
  .B1({ S11117 }),
  .B2({ S11118 }),
  .ZN({ S11120 })
);
NAND4_X1 #() 
NAND4_X1_140_ (
  .A1({ S10569 }),
  .A2({ S21 }),
  .A3({ S10562 }),
  .A4({ S10538 }),
  .ZN({ S11121 })
);
NAND3_X1 #() 
NAND3_X1_1191_ (
  .A1({ S10925 }),
  .A2({ S11121 }),
  .A3({ S10526 }),
  .ZN({ S11122 })
);
OAI21_X1 #() 
OAI21_X1_575_ (
  .A({ S25957[396] }),
  .B1({ S10531 }),
  .B2({ S10769 }),
  .ZN({ S11123 })
);
OAI211_X1 #() 
OAI211_X1_376_ (
  .A({ S11122 }),
  .B({ S10559 }),
  .C1({ S11123 }),
  .C2({ S11010 }),
  .ZN({ S11124 })
);
OAI211_X1 #() 
OAI211_X1_377_ (
  .A({ S11124 }),
  .B({ S25957[398] }),
  .C1({ S11120 }),
  .C2({ S10559 }),
  .ZN({ S11125 })
);
NAND3_X1 #() 
NAND3_X1_1192_ (
  .A1({ S11125 }),
  .A2({ S10598 }),
  .A3({ S11114 }),
  .ZN({ S11127 })
);
NAND3_X1 #() 
NAND3_X1_1193_ (
  .A1({ S11127 }),
  .A2({ S11108 }),
  .A3({ S11087 }),
  .ZN({ S11128 })
);
INV_X1 #() 
INV_X1_334_ (
  .A({ S11087 }),
  .ZN({ S25957[593] })
);
NOR2_X1 #() 
NOR2_X1_243_ (
  .A1({ S10636 }),
  .A2({ S25957[395] }),
  .ZN({ S11129 })
);
OAI21_X1 #() 
OAI21_X1_576_ (
  .A({ S10526 }),
  .B1({ S11010 }),
  .B2({ S11129 }),
  .ZN({ S11130 })
);
NAND2_X1 #() 
NAND2_X1_1022_ (
  .A1({ S10605 }),
  .A2({ S11102 }),
  .ZN({ S11131 })
);
AOI21_X1 #() 
AOI21_X1_639_ (
  .A({ S10559 }),
  .B1({ S11131 }),
  .B2({ S25957[396] }),
  .ZN({ S11132 })
);
NAND2_X1 #() 
NAND2_X1_1023_ (
  .A1({ S11130 }),
  .A2({ S11132 }),
  .ZN({ S11133 })
);
NAND2_X1 #() 
NAND2_X1_1024_ (
  .A1({ S10774 }),
  .A2({ S11097 }),
  .ZN({ S11134 })
);
NAND2_X1 #() 
NAND2_X1_1025_ (
  .A1({ S11134 }),
  .A2({ S25957[396] }),
  .ZN({ S11135 })
);
OAI21_X1 #() 
OAI21_X1_577_ (
  .A({ S11099 }),
  .B1({ S10949 }),
  .B2({ S10750 }),
  .ZN({ S11137 })
);
AOI21_X1 #() 
AOI21_X1_640_ (
  .A({ S25957[397] }),
  .B1({ S11137 }),
  .B2({ S10526 }),
  .ZN({ S11138 })
);
NAND2_X1 #() 
NAND2_X1_1026_ (
  .A1({ S11135 }),
  .A2({ S11138 }),
  .ZN({ S11139 })
);
NAND3_X1 #() 
NAND3_X1_1194_ (
  .A1({ S11139 }),
  .A2({ S25957[398] }),
  .A3({ S11133 }),
  .ZN({ S11140 })
);
OAI21_X1 #() 
OAI21_X1_578_ (
  .A({ S11094 }),
  .B1({ S11091 }),
  .B2({ S10601 }),
  .ZN({ S11141 })
);
NAND2_X1 #() 
NAND2_X1_1027_ (
  .A1({ S11141 }),
  .A2({ S25957[397] }),
  .ZN({ S11142 })
);
NOR2_X1 #() 
NOR2_X1_244_ (
  .A1({ S10568 }),
  .A2({ S21 }),
  .ZN({ S11143 })
);
OAI21_X1 #() 
OAI21_X1_579_ (
  .A({ S25957[396] }),
  .B1({ S11089 }),
  .B2({ S11143 }),
  .ZN({ S11144 })
);
OAI21_X1 #() 
OAI21_X1_580_ (
  .A({ S10526 }),
  .B1({ S10611 }),
  .B2({ S10887 }),
  .ZN({ S11145 })
);
NAND3_X1 #() 
NAND3_X1_1195_ (
  .A1({ S11145 }),
  .A2({ S10559 }),
  .A3({ S11144 }),
  .ZN({ S11146 })
);
NAND3_X1 #() 
NAND3_X1_1196_ (
  .A1({ S11146 }),
  .A2({ S11142 }),
  .A3({ S8507 }),
  .ZN({ S11148 })
);
NAND3_X1 #() 
NAND3_X1_1197_ (
  .A1({ S11140 }),
  .A2({ S11148 }),
  .A3({ S25957[399] }),
  .ZN({ S11149 })
);
NOR2_X1 #() 
NOR2_X1_245_ (
  .A1({ S10527 }),
  .A2({ S25957[394] }),
  .ZN({ S11150 })
);
OAI21_X1 #() 
OAI21_X1_581_ (
  .A({ S25957[395] }),
  .B1({ S10583 }),
  .B2({ S11150 }),
  .ZN({ S11151 })
);
AOI21_X1 #() 
AOI21_X1_641_ (
  .A({ S25957[396] }),
  .B1({ S10551 }),
  .B2({ S10609 }),
  .ZN({ S11152 })
);
AOI22_X1 #() 
AOI22_X1_134_ (
  .A1({ S10584 }),
  .A2({ S10528 }),
  .B1({ S8762 }),
  .B2({ S8759 }),
  .ZN({ S11153 })
);
NAND3_X1 #() 
NAND3_X1_1198_ (
  .A1({ S25957[394] }),
  .A2({ S25957[393] }),
  .A3({ S25957[392] }),
  .ZN({ S11154 })
);
AOI21_X1 #() 
AOI21_X1_642_ (
  .A({ S10526 }),
  .B1({ S11153 }),
  .B2({ S11154 }),
  .ZN({ S11155 })
);
AOI22_X1 #() 
AOI22_X1_135_ (
  .A1({ S11155 }),
  .A2({ S11151 }),
  .B1({ S11152 }),
  .B2({ S10925 }),
  .ZN({ S11156 })
);
AOI21_X1 #() 
AOI21_X1_643_ (
  .A({ S10526 }),
  .B1({ S10933 }),
  .B2({ S25957[395] }),
  .ZN({ S11157 })
);
INV_X1 #() 
INV_X1_335_ (
  .A({ S11118 }),
  .ZN({ S11159 })
);
AOI21_X1 #() 
AOI21_X1_644_ (
  .A({ S10559 }),
  .B1({ S11035 }),
  .B2({ S10551 }),
  .ZN({ S11160 })
);
OAI21_X1 #() 
OAI21_X1_582_ (
  .A({ S11160 }),
  .B1({ S11157 }),
  .B2({ S11159 }),
  .ZN({ S11161 })
);
OAI211_X1 #() 
OAI211_X1_378_ (
  .A({ S11161 }),
  .B({ S25957[398] }),
  .C1({ S11156 }),
  .C2({ S25957[397] }),
  .ZN({ S11162 })
);
INV_X1 #() 
INV_X1_336_ (
  .A({ S11109 }),
  .ZN({ S11163 })
);
NAND2_X1 #() 
NAND2_X1_1028_ (
  .A1({ S10616 }),
  .A2({ S21 }),
  .ZN({ S11164 })
);
AOI21_X1 #() 
AOI21_X1_645_ (
  .A({ S10559 }),
  .B1({ S11164 }),
  .B2({ S10526 }),
  .ZN({ S11165 })
);
NAND2_X1 #() 
NAND2_X1_1029_ (
  .A1({ S11165 }),
  .A2({ S11163 }),
  .ZN({ S11166 })
);
OAI211_X1 #() 
OAI211_X1_379_ (
  .A({ S10517 }),
  .B({ S10513 }),
  .C1({ S10568 }),
  .C2({ S25957[395] }),
  .ZN({ S11167 })
);
NAND2_X1 #() 
NAND2_X1_1030_ (
  .A1({ S11167 }),
  .A2({ S25957[396] }),
  .ZN({ S11168 })
);
OAI211_X1 #() 
OAI211_X1_380_ (
  .A({ S11168 }),
  .B({ S10559 }),
  .C1({ S10682 }),
  .C2({ S25957[396] }),
  .ZN({ S11170 })
);
NAND3_X1 #() 
NAND3_X1_1199_ (
  .A1({ S11166 }),
  .A2({ S11170 }),
  .A3({ S8507 }),
  .ZN({ S11171 })
);
NAND3_X1 #() 
NAND3_X1_1200_ (
  .A1({ S11162 }),
  .A2({ S11171 }),
  .A3({ S10598 }),
  .ZN({ S11172 })
);
NAND3_X1 #() 
NAND3_X1_1201_ (
  .A1({ S11149 }),
  .A2({ S25957[593] }),
  .A3({ S11172 }),
  .ZN({ S11173 })
);
AOI21_X1 #() 
AOI21_X1_646_ (
  .A({ S11086 }),
  .B1({ S11173 }),
  .B2({ S11128 }),
  .ZN({ S11174 })
);
AND3_X1 #() 
AND3_X1_48_ (
  .A1({ S11173 }),
  .A2({ S11128 }),
  .A3({ S11086 }),
  .ZN({ S11175 })
);
OAI21_X1 #() 
OAI21_X1_583_ (
  .A({ S25957[401] }),
  .B1({ S11175 }),
  .B2({ S11174 }),
  .ZN({ S11176 })
);
AOI21_X1 #() 
AOI21_X1_647_ (
  .A({ S25957[529] }),
  .B1({ S8200 }),
  .B2({ S8201 }),
  .ZN({ S11177 })
);
AND3_X1 #() 
AND3_X1_49_ (
  .A1({ S8201 }),
  .A2({ S8200 }),
  .A3({ S25957[529] }),
  .ZN({ S11178 })
);
NOR2_X1 #() 
NOR2_X1_246_ (
  .A1({ S11178 }),
  .A2({ S11177 }),
  .ZN({ S11179 })
);
INV_X1 #() 
INV_X1_337_ (
  .A({ S11086 }),
  .ZN({ S25957[433] })
);
AND3_X1 #() 
AND3_X1_50_ (
  .A1({ S11127 }),
  .A2({ S11108 }),
  .A3({ S11087 }),
  .ZN({ S11181 })
);
AOI21_X1 #() 
AOI21_X1_648_ (
  .A({ S11087 }),
  .B1({ S11127 }),
  .B2({ S11108 }),
  .ZN({ S11182 })
);
OAI21_X1 #() 
OAI21_X1_584_ (
  .A({ S25957[433] }),
  .B1({ S11181 }),
  .B2({ S11182 }),
  .ZN({ S11183 })
);
NAND3_X1 #() 
NAND3_X1_1202_ (
  .A1({ S11173 }),
  .A2({ S11086 }),
  .A3({ S11128 }),
  .ZN({ S11184 })
);
NAND3_X1 #() 
NAND3_X1_1203_ (
  .A1({ S11183 }),
  .A2({ S11179 }),
  .A3({ S11184 }),
  .ZN({ S11185 })
);
NAND2_X1 #() 
NAND2_X1_1031_ (
  .A1({ S11176 }),
  .A2({ S11185 }),
  .ZN({ S25957[273] })
);
NAND2_X1 #() 
NAND2_X1_1032_ (
  .A1({ S5452 }),
  .A2({ S5453 }),
  .ZN({ S25957[626] })
);
NAND2_X1 #() 
NAND2_X1_1033_ (
  .A1({ S8253 }),
  .A2({ S8226 }),
  .ZN({ S11186 })
);
XOR2_X1 #() 
XOR2_X1_20_ (
  .A({ S11186 }),
  .B({ S25957[626] }),
  .Z({ S11187 })
);
INV_X1 #() 
INV_X1_338_ (
  .A({ S11187 }),
  .ZN({ S25957[498] })
);
NAND3_X1 #() 
NAND3_X1_1204_ (
  .A1({ S25957[395] }),
  .A2({ S10569 }),
  .A3({ S25957[393] }),
  .ZN({ S11189 })
);
NAND3_X1 #() 
NAND3_X1_1205_ (
  .A1({ S10853 }),
  .A2({ S11189 }),
  .A3({ S10526 }),
  .ZN({ S11190 })
);
AOI21_X1 #() 
AOI21_X1_649_ (
  .A({ S21 }),
  .B1({ S10885 }),
  .B2({ S10538 }),
  .ZN({ S11191 })
);
AOI21_X1 #() 
AOI21_X1_650_ (
  .A({ S25957[395] }),
  .B1({ S10854 }),
  .B2({ S10622 }),
  .ZN({ S11192 })
);
OAI21_X1 #() 
OAI21_X1_585_ (
  .A({ S25957[396] }),
  .B1({ S11192 }),
  .B2({ S11191 }),
  .ZN({ S11193 })
);
NAND3_X1 #() 
NAND3_X1_1206_ (
  .A1({ S11193 }),
  .A2({ S10559 }),
  .A3({ S11190 }),
  .ZN({ S11194 })
);
NAND2_X1 #() 
NAND2_X1_1034_ (
  .A1({ S10866 }),
  .A2({ S10786 }),
  .ZN({ S11195 })
);
OAI21_X1 #() 
OAI21_X1_586_ (
  .A({ S25957[396] }),
  .B1({ S11195 }),
  .B2({ S10729 }),
  .ZN({ S11196 })
);
OAI21_X1 #() 
OAI21_X1_587_ (
  .A({ S10526 }),
  .B1({ S10580 }),
  .B2({ S10539 }),
  .ZN({ S11197 })
);
OAI211_X1 #() 
OAI211_X1_381_ (
  .A({ S11196 }),
  .B({ S25957[397] }),
  .C1({ S10549 }),
  .C2({ S11197 }),
  .ZN({ S11199 })
);
NAND3_X1 #() 
NAND3_X1_1207_ (
  .A1({ S11194 }),
  .A2({ S11199 }),
  .A3({ S25957[398] }),
  .ZN({ S11200 })
);
OAI21_X1 #() 
OAI21_X1_588_ (
  .A({ S25957[395] }),
  .B1({ S10696 }),
  .B2({ S10769 }),
  .ZN({ S11201 })
);
AOI21_X1 #() 
AOI21_X1_651_ (
  .A({ S25957[396] }),
  .B1({ S10659 }),
  .B2({ S21 }),
  .ZN({ S11202 })
);
NAND2_X1 #() 
NAND2_X1_1035_ (
  .A1({ S11201 }),
  .A2({ S11202 }),
  .ZN({ S11203 })
);
AOI22_X1 #() 
AOI22_X1_136_ (
  .A1({ S10530 }),
  .A2({ S10628 }),
  .B1({ S10903 }),
  .B2({ S10545 }),
  .ZN({ S11204 })
);
OAI211_X1 #() 
OAI211_X1_382_ (
  .A({ S25957[397] }),
  .B({ S11203 }),
  .C1({ S11204 }),
  .C2({ S10526 }),
  .ZN({ S11205 })
);
AOI21_X1 #() 
AOI21_X1_652_ (
  .A({ S25957[395] }),
  .B1({ S10739 }),
  .B2({ S10622 }),
  .ZN({ S11206 })
);
NOR2_X1 #() 
NOR2_X1_247_ (
  .A1({ S10786 }),
  .A2({ S10589 }),
  .ZN({ S11207 })
);
OAI21_X1 #() 
OAI21_X1_589_ (
  .A({ S25957[396] }),
  .B1({ S11206 }),
  .B2({ S11207 }),
  .ZN({ S11208 })
);
NAND4_X1 #() 
NAND4_X1_141_ (
  .A1({ S10536 }),
  .A2({ S10535 }),
  .A3({ S21 }),
  .A4({ S10526 }),
  .ZN({ S11210 })
);
NAND4_X1 #() 
NAND4_X1_142_ (
  .A1({ S11208 }),
  .A2({ S11210 }),
  .A3({ S10559 }),
  .A4({ S10705 }),
  .ZN({ S11211 })
);
NAND3_X1 #() 
NAND3_X1_1208_ (
  .A1({ S11211 }),
  .A2({ S11205 }),
  .A3({ S8507 }),
  .ZN({ S11212 })
);
NAND3_X1 #() 
NAND3_X1_1209_ (
  .A1({ S11212 }),
  .A2({ S10598 }),
  .A3({ S11200 }),
  .ZN({ S11213 })
);
NAND3_X1 #() 
NAND3_X1_1210_ (
  .A1({ S10536 }),
  .A2({ S25957[395] }),
  .A3({ S10854 }),
  .ZN({ S11214 })
);
NAND3_X1 #() 
NAND3_X1_1211_ (
  .A1({ S11214 }),
  .A2({ S25957[396] }),
  .A3({ S10756 }),
  .ZN({ S11215 })
);
NAND3_X1 #() 
NAND3_X1_1212_ (
  .A1({ S10536 }),
  .A2({ S25957[395] }),
  .A3({ S10739 }),
  .ZN({ S11216 })
);
NAND3_X1 #() 
NAND3_X1_1213_ (
  .A1({ S11216 }),
  .A2({ S10526 }),
  .A3({ S10787 }),
  .ZN({ S11217 })
);
NAND2_X1 #() 
NAND2_X1_1036_ (
  .A1({ S10541 }),
  .A2({ S10538 }),
  .ZN({ S11218 })
);
AOI21_X1 #() 
AOI21_X1_653_ (
  .A({ S10526 }),
  .B1({ S11218 }),
  .B2({ S25957[395] }),
  .ZN({ S11219 })
);
AOI21_X1 #() 
AOI21_X1_654_ (
  .A({ S10559 }),
  .B1({ S11019 }),
  .B2({ S11219 }),
  .ZN({ S11221 })
);
AOI21_X1 #() 
AOI21_X1_655_ (
  .A({ S25957[396] }),
  .B1({ S21 }),
  .B2({ S10584 }),
  .ZN({ S11222 })
);
AOI21_X1 #() 
AOI21_X1_656_ (
  .A({ S25957[397] }),
  .B1({ S11222 }),
  .B2({ S10623 }),
  .ZN({ S11223 })
);
AOI22_X1 #() 
AOI22_X1_137_ (
  .A1({ S11221 }),
  .A2({ S11217 }),
  .B1({ S11223 }),
  .B2({ S11215 }),
  .ZN({ S11224 })
);
OAI21_X1 #() 
OAI21_X1_590_ (
  .A({ S25957[396] }),
  .B1({ S10938 }),
  .B2({ S11207 }),
  .ZN({ S11225 })
);
NAND2_X1 #() 
NAND2_X1_1037_ (
  .A1({ S10655 }),
  .A2({ S10526 }),
  .ZN({ S11226 })
);
NAND3_X1 #() 
NAND3_X1_1214_ (
  .A1({ S11225 }),
  .A2({ S11226 }),
  .A3({ S10559 }),
  .ZN({ S11227 })
);
AOI21_X1 #() 
AOI21_X1_657_ (
  .A({ S25957[396] }),
  .B1({ S10689 }),
  .B2({ S21 }),
  .ZN({ S11228 })
);
OAI211_X1 #() 
OAI211_X1_383_ (
  .A({ S25957[395] }),
  .B({ S10546 }),
  .C1({ S10547 }),
  .C2({ S10529 }),
  .ZN({ S11229 })
);
OAI21_X1 #() 
OAI21_X1_591_ (
  .A({ S25957[396] }),
  .B1({ S21 }),
  .B2({ S10527 }),
  .ZN({ S11230 })
);
NOR2_X1 #() 
NOR2_X1_248_ (
  .A1({ S11230 }),
  .A2({ S10519 }),
  .ZN({ S11232 })
);
AOI22_X1 #() 
AOI22_X1_138_ (
  .A1({ S11232 }),
  .A2({ S10946 }),
  .B1({ S11228 }),
  .B2({ S11229 }),
  .ZN({ S11233 })
);
OAI211_X1 #() 
OAI211_X1_384_ (
  .A({ S11227 }),
  .B({ S8507 }),
  .C1({ S11233 }),
  .C2({ S10559 }),
  .ZN({ S11234 })
);
OAI211_X1 #() 
OAI211_X1_385_ (
  .A({ S11234 }),
  .B({ S25957[399] }),
  .C1({ S11224 }),
  .C2({ S8507 }),
  .ZN({ S11235 })
);
NAND3_X1 #() 
NAND3_X1_1215_ (
  .A1({ S11235 }),
  .A2({ S11213 }),
  .A3({ S25957[498] }),
  .ZN({ S11236 })
);
NAND2_X1 #() 
NAND2_X1_1038_ (
  .A1({ S11221 }),
  .A2({ S11217 }),
  .ZN({ S11237 })
);
NAND2_X1 #() 
NAND2_X1_1039_ (
  .A1({ S11215 }),
  .A2({ S11223 }),
  .ZN({ S11238 })
);
NAND3_X1 #() 
NAND3_X1_1216_ (
  .A1({ S11237 }),
  .A2({ S25957[398] }),
  .A3({ S11238 }),
  .ZN({ S11239 })
);
NAND2_X1 #() 
NAND2_X1_1040_ (
  .A1({ S11228 }),
  .A2({ S11229 }),
  .ZN({ S11240 })
);
NAND2_X1 #() 
NAND2_X1_1041_ (
  .A1({ S11232 }),
  .A2({ S10946 }),
  .ZN({ S11241 })
);
NAND3_X1 #() 
NAND3_X1_1217_ (
  .A1({ S11241 }),
  .A2({ S11240 }),
  .A3({ S25957[397] }),
  .ZN({ S11243 })
);
NAND2_X1 #() 
NAND2_X1_1042_ (
  .A1({ S10568 }),
  .A2({ S21 }),
  .ZN({ S11244 })
);
NAND3_X1 #() 
NAND3_X1_1218_ (
  .A1({ S11189 }),
  .A2({ S25957[396] }),
  .A3({ S11244 }),
  .ZN({ S11245 })
);
OAI211_X1 #() 
OAI211_X1_386_ (
  .A({ S11245 }),
  .B({ S10559 }),
  .C1({ S25957[396] }),
  .C2({ S10655 }),
  .ZN({ S11246 })
);
NAND3_X1 #() 
NAND3_X1_1219_ (
  .A1({ S11243 }),
  .A2({ S11246 }),
  .A3({ S8507 }),
  .ZN({ S11247 })
);
NAND3_X1 #() 
NAND3_X1_1220_ (
  .A1({ S11239 }),
  .A2({ S25957[399] }),
  .A3({ S11247 }),
  .ZN({ S11248 })
);
NAND3_X1 #() 
NAND3_X1_1221_ (
  .A1({ S10560 }),
  .A2({ S21 }),
  .A3({ S10529 }),
  .ZN({ S11249 })
);
NAND3_X1 #() 
NAND3_X1_1222_ (
  .A1({ S11154 }),
  .A2({ S10622 }),
  .A3({ S25957[395] }),
  .ZN({ S11250 })
);
AOI21_X1 #() 
AOI21_X1_658_ (
  .A({ S25957[396] }),
  .B1({ S11250 }),
  .B2({ S11249 }),
  .ZN({ S11251 })
);
NAND3_X1 #() 
NAND3_X1_1223_ (
  .A1({ S10530 }),
  .A2({ S25957[395] }),
  .A3({ S10513 }),
  .ZN({ S11252 })
);
AOI21_X1 #() 
AOI21_X1_659_ (
  .A({ S10526 }),
  .B1({ S10905 }),
  .B2({ S11252 }),
  .ZN({ S11254 })
);
OAI21_X1 #() 
OAI21_X1_592_ (
  .A({ S25957[397] }),
  .B1({ S11254 }),
  .B2({ S11251 }),
  .ZN({ S11255 })
);
AOI21_X1 #() 
AOI21_X1_660_ (
  .A({ S10526 }),
  .B1({ S10863 }),
  .B2({ S11189 }),
  .ZN({ S11256 })
);
OAI21_X1 #() 
OAI21_X1_593_ (
  .A({ S25957[395] }),
  .B1({ S10704 }),
  .B2({ S10636 }),
  .ZN({ S11257 })
);
NAND3_X1 #() 
NAND3_X1_1224_ (
  .A1({ S10536 }),
  .A2({ S21 }),
  .A3({ S10535 }),
  .ZN({ S11258 })
);
AOI21_X1 #() 
AOI21_X1_661_ (
  .A({ S25957[396] }),
  .B1({ S11257 }),
  .B2({ S11258 }),
  .ZN({ S11259 })
);
OAI21_X1 #() 
OAI21_X1_594_ (
  .A({ S10559 }),
  .B1({ S11259 }),
  .B2({ S11256 }),
  .ZN({ S11260 })
);
NAND3_X1 #() 
NAND3_X1_1225_ (
  .A1({ S11260 }),
  .A2({ S8507 }),
  .A3({ S11255 }),
  .ZN({ S11261 })
);
OAI21_X1 #() 
OAI21_X1_595_ (
  .A({ S11196 }),
  .B1({ S10549 }),
  .B2({ S11197 }),
  .ZN({ S11262 })
);
NAND2_X1 #() 
NAND2_X1_1043_ (
  .A1({ S11262 }),
  .A2({ S25957[397] }),
  .ZN({ S11263 })
);
INV_X1 #() 
INV_X1_339_ (
  .A({ S11190 }),
  .ZN({ S11265 })
);
NAND3_X1 #() 
NAND3_X1_1226_ (
  .A1({ S10659 }),
  .A2({ S25957[395] }),
  .A3({ S10513 }),
  .ZN({ S11266 })
);
OAI21_X1 #() 
OAI21_X1_596_ (
  .A({ S21 }),
  .B1({ S10696 }),
  .B2({ S10916 }),
  .ZN({ S11267 })
);
AOI21_X1 #() 
AOI21_X1_662_ (
  .A({ S10526 }),
  .B1({ S11267 }),
  .B2({ S11266 }),
  .ZN({ S11268 })
);
OAI21_X1 #() 
OAI21_X1_597_ (
  .A({ S10559 }),
  .B1({ S11268 }),
  .B2({ S11265 }),
  .ZN({ S11269 })
);
NAND3_X1 #() 
NAND3_X1_1227_ (
  .A1({ S11263 }),
  .A2({ S11269 }),
  .A3({ S25957[398] }),
  .ZN({ S11270 })
);
NAND3_X1 #() 
NAND3_X1_1228_ (
  .A1({ S11261 }),
  .A2({ S11270 }),
  .A3({ S10598 }),
  .ZN({ S11271 })
);
NAND3_X1 #() 
NAND3_X1_1229_ (
  .A1({ S11271 }),
  .A2({ S11187 }),
  .A3({ S11248 }),
  .ZN({ S11272 })
);
AOI21_X1 #() 
AOI21_X1_663_ (
  .A({ S8283 }),
  .B1({ S11272 }),
  .B2({ S11236 }),
  .ZN({ S11273 })
);
NAND3_X1 #() 
NAND3_X1_1230_ (
  .A1({ S11271 }),
  .A2({ S25957[498] }),
  .A3({ S11248 }),
  .ZN({ S11274 })
);
NAND3_X1 #() 
NAND3_X1_1231_ (
  .A1({ S11235 }),
  .A2({ S11213 }),
  .A3({ S11187 }),
  .ZN({ S11276 })
);
AOI21_X1 #() 
AOI21_X1_664_ (
  .A({ S25957[562] }),
  .B1({ S11274 }),
  .B2({ S11276 }),
  .ZN({ S11277 })
);
OAI21_X1 #() 
OAI21_X1_598_ (
  .A({ S25957[402] }),
  .B1({ S11273 }),
  .B2({ S11277 }),
  .ZN({ S11278 })
);
OAI21_X1 #() 
OAI21_X1_599_ (
  .A({ S8281 }),
  .B1({ S8273 }),
  .B2({ S8272 }),
  .ZN({ S11279 })
);
NAND3_X1 #() 
NAND3_X1_1232_ (
  .A1({ S8286 }),
  .A2({ S25957[530] }),
  .A3({ S8287 }),
  .ZN({ S11280 })
);
NAND2_X1 #() 
NAND2_X1_1044_ (
  .A1({ S11279 }),
  .A2({ S11280 }),
  .ZN({ S11281 })
);
NAND3_X1 #() 
NAND3_X1_1233_ (
  .A1({ S11274 }),
  .A2({ S11276 }),
  .A3({ S25957[562] }),
  .ZN({ S11282 })
);
NAND3_X1 #() 
NAND3_X1_1234_ (
  .A1({ S11272 }),
  .A2({ S11236 }),
  .A3({ S8283 }),
  .ZN({ S11283 })
);
NAND3_X1 #() 
NAND3_X1_1235_ (
  .A1({ S11282 }),
  .A2({ S11283 }),
  .A3({ S11281 }),
  .ZN({ S11284 })
);
NAND2_X1 #() 
NAND2_X1_1045_ (
  .A1({ S11278 }),
  .A2({ S11284 }),
  .ZN({ S25957[274] })
);
NAND3_X1 #() 
NAND3_X1_1236_ (
  .A1({ S9613 }),
  .A2({ S5479 }),
  .A3({ S9582 }),
  .ZN({ S11286 })
);
OAI21_X1 #() 
OAI21_X1_600_ (
  .A({ S25957[640] }),
  .B1({ S9579 }),
  .B2({ S9580 }),
  .ZN({ S11287 })
);
AND3_X1 #() 
AND3_X1_51_ (
  .A1({ S9637 }),
  .A2({ S6817 }),
  .A3({ S9656 }),
  .ZN({ S11288 })
);
AOI21_X1 #() 
AOI21_X1_665_ (
  .A({ S6817 }),
  .B1({ S9637 }),
  .B2({ S9656 }),
  .ZN({ S11289 })
);
OAI21_X1 #() 
OAI21_X1_601_ (
  .A({ S25957[641] }),
  .B1({ S11288 }),
  .B2({ S11289 }),
  .ZN({ S11290 })
);
NAND3_X1 #() 
NAND3_X1_1237_ (
  .A1({ S9700 }),
  .A2({ S5464 }),
  .A3({ S9657 }),
  .ZN({ S11291 })
);
NAND4_X1 #() 
NAND4_X1_143_ (
  .A1({ S11287 }),
  .A2({ S11290 }),
  .A3({ S11286 }),
  .A4({ S11291 }),
  .ZN({ S11292 })
);
INV_X1 #() 
INV_X1_340_ (
  .A({ S11292 }),
  .ZN({ S33 })
);
OAI211_X1 #() 
OAI211_X1_387_ (
  .A({ S9581 }),
  .B({ S9614 }),
  .C1({ S9702 }),
  .C2({ S9701 }),
  .ZN({ S34 })
);
INV_X1 #() 
INV_X1_341_ (
  .A({ S25957[389] }),
  .ZN({ S11293 })
);
AOI21_X1 #() 
AOI21_X1_666_ (
  .A({ S5471 }),
  .B1({ S9784 }),
  .B2({ S9785 }),
  .ZN({ S11295 })
);
AND3_X1 #() 
AND3_X1_52_ (
  .A1({ S9784 }),
  .A2({ S5471 }),
  .A3({ S9785 }),
  .ZN({ S11296 })
);
OAI211_X1 #() 
OAI211_X1_388_ (
  .A({ S11290 }),
  .B({ S11291 }),
  .C1({ S11296 }),
  .C2({ S11295 }),
  .ZN({ S11297 })
);
NOR2_X1 #() 
NOR2_X1_249_ (
  .A1({ S11296 }),
  .A2({ S11295 }),
  .ZN({ S11298 })
);
NAND3_X1 #() 
NAND3_X1_1238_ (
  .A1({ S34 }),
  .A2({ S11292 }),
  .A3({ S11298 }),
  .ZN({ S11299 })
);
NAND2_X1 #() 
NAND2_X1_1046_ (
  .A1({ S11287 }),
  .A2({ S11286 }),
  .ZN({ S11300 })
);
NAND2_X1 #() 
NAND2_X1_1047_ (
  .A1({ S25957[386] }),
  .A2({ S11300 }),
  .ZN({ S11301 })
);
NAND2_X1 #() 
NAND2_X1_1048_ (
  .A1({ S24 }),
  .A2({ S11301 }),
  .ZN({ S11302 })
);
INV_X1 #() 
INV_X1_342_ (
  .A({ S11302 }),
  .ZN({ S11303 })
);
NAND3_X1 #() 
NAND3_X1_1239_ (
  .A1({ S11303 }),
  .A2({ S11297 }),
  .A3({ S11299 }),
  .ZN({ S11304 })
);
NOR2_X1 #() 
NOR2_X1_250_ (
  .A1({ S25957[386] }),
  .A2({ S25957[385] }),
  .ZN({ S11306 })
);
AOI21_X1 #() 
AOI21_X1_667_ (
  .A({ S25957[388] }),
  .B1({ S25957[387] }),
  .B2({ S11306 }),
  .ZN({ S11307 })
);
NAND2_X1 #() 
NAND2_X1_1049_ (
  .A1({ S24 }),
  .A2({ S11297 }),
  .ZN({ S11308 })
);
NAND4_X1 #() 
NAND4_X1_144_ (
  .A1({ S9781 }),
  .A2({ S11287 }),
  .A3({ S11286 }),
  .A4({ S9786 }),
  .ZN({ S11309 })
);
INV_X1 #() 
INV_X1_343_ (
  .A({ S11309 }),
  .ZN({ S11310 })
);
OAI211_X1 #() 
OAI211_X1_389_ (
  .A({ S11286 }),
  .B({ S11287 }),
  .C1({ S9702 }),
  .C2({ S9701 }),
  .ZN({ S11311 })
);
NAND4_X1 #() 
NAND4_X1_145_ (
  .A1({ S9581 }),
  .A2({ S11290 }),
  .A3({ S9614 }),
  .A4({ S11291 }),
  .ZN({ S11312 })
);
NAND3_X1 #() 
NAND3_X1_1240_ (
  .A1({ S11311 }),
  .A2({ S11312 }),
  .A3({ S25957[386] }),
  .ZN({ S11313 })
);
NAND3_X1 #() 
NAND3_X1_1241_ (
  .A1({ S11313 }),
  .A2({ S11299 }),
  .A3({ S25957[387] }),
  .ZN({ S11314 })
);
OAI21_X1 #() 
OAI21_X1_602_ (
  .A({ S11314 }),
  .B1({ S11308 }),
  .B2({ S11310 }),
  .ZN({ S11315 })
);
AOI22_X1 #() 
AOI22_X1_139_ (
  .A1({ S11315 }),
  .A2({ S25957[388] }),
  .B1({ S11304 }),
  .B2({ S11307 }),
  .ZN({ S11317 })
);
AOI22_X1 #() 
AOI22_X1_140_ (
  .A1({ S11287 }),
  .A2({ S11286 }),
  .B1({ S11290 }),
  .B2({ S11291 }),
  .ZN({ S11318 })
);
NAND2_X1 #() 
NAND2_X1_1050_ (
  .A1({ S11318 }),
  .A2({ S11298 }),
  .ZN({ S11319 })
);
NAND2_X1 #() 
NAND2_X1_1051_ (
  .A1({ S11319 }),
  .A2({ S24 }),
  .ZN({ S11320 })
);
AOI21_X1 #() 
AOI21_X1_668_ (
  .A({ S25957[388] }),
  .B1({ S11320 }),
  .B2({ S11292 }),
  .ZN({ S11321 })
);
NOR2_X1 #() 
NOR2_X1_251_ (
  .A1({ S11298 }),
  .A2({ S11300 }),
  .ZN({ S11322 })
);
NAND2_X1 #() 
NAND2_X1_1052_ (
  .A1({ S24 }),
  .A2({ S25957[385] }),
  .ZN({ S11323 })
);
NAND2_X1 #() 
NAND2_X1_1053_ (
  .A1({ S11290 }),
  .A2({ S11291 }),
  .ZN({ S11324 })
);
OAI21_X1 #() 
OAI21_X1_603_ (
  .A({ S25957[387] }),
  .B1({ S11322 }),
  .B2({ S11324 }),
  .ZN({ S11325 })
);
OAI21_X1 #() 
OAI21_X1_604_ (
  .A({ S11325 }),
  .B1({ S11322 }),
  .B2({ S11323 }),
  .ZN({ S11326 })
);
AOI21_X1 #() 
AOI21_X1_669_ (
  .A({ S11321 }),
  .B1({ S11326 }),
  .B2({ S25957[388] }),
  .ZN({ S11328 })
);
MUX2_X1 #() 
MUX2_X1_3_ (
  .A({ S11328 }),
  .B({ S11317 }),
  .S({ S11293 }),
  .Z({ S11329 })
);
OAI21_X1 #() 
OAI21_X1_605_ (
  .A({ S5495 }),
  .B1({ S9412 }),
  .B2({ S9411 }),
  .ZN({ S11330 })
);
NAND3_X1 #() 
NAND3_X1_1242_ (
  .A1({ S9405 }),
  .A2({ S9409 }),
  .A3({ S25957[644] }),
  .ZN({ S11331 })
);
NAND2_X1 #() 
NAND2_X1_1054_ (
  .A1({ S11330 }),
  .A2({ S11331 }),
  .ZN({ S11332 })
);
AOI21_X1 #() 
AOI21_X1_670_ (
  .A({ S24 }),
  .B1({ S11324 }),
  .B2({ S25957[386] }),
  .ZN({ S11333 })
);
INV_X1 #() 
INV_X1_344_ (
  .A({ S11333 }),
  .ZN({ S11334 })
);
NAND2_X1 #() 
NAND2_X1_1055_ (
  .A1({ S24 }),
  .A2({ S11312 }),
  .ZN({ S11335 })
);
OAI21_X1 #() 
OAI21_X1_606_ (
  .A({ S11335 }),
  .B1({ S11334 }),
  .B2({ S33 }),
  .ZN({ S11336 })
);
NAND2_X1 #() 
NAND2_X1_1056_ (
  .A1({ S34 }),
  .A2({ S25957[386] }),
  .ZN({ S11337 })
);
AOI22_X1 #() 
AOI22_X1_141_ (
  .A1({ S9614 }),
  .A2({ S9581 }),
  .B1({ S11290 }),
  .B2({ S11291 }),
  .ZN({ S11339 })
);
NAND2_X1 #() 
NAND2_X1_1057_ (
  .A1({ S25957[387] }),
  .A2({ S11339 }),
  .ZN({ S11340 })
);
NAND3_X1 #() 
NAND3_X1_1243_ (
  .A1({ S11340 }),
  .A2({ S11337 }),
  .A3({ S11319 }),
  .ZN({ S11341 })
);
NAND2_X1 #() 
NAND2_X1_1058_ (
  .A1({ S11341 }),
  .A2({ S11332 }),
  .ZN({ S11342 })
);
OAI21_X1 #() 
OAI21_X1_607_ (
  .A({ S11342 }),
  .B1({ S11336 }),
  .B2({ S11332 }),
  .ZN({ S11343 })
);
NAND2_X1 #() 
NAND2_X1_1059_ (
  .A1({ S34 }),
  .A2({ S11292 }),
  .ZN({ S11344 })
);
NAND3_X1 #() 
NAND3_X1_1244_ (
  .A1({ S11298 }),
  .A2({ S25957[384] }),
  .A3({ S25957[385] }),
  .ZN({ S11345 })
);
NAND3_X1 #() 
NAND3_X1_1245_ (
  .A1({ S25957[386] }),
  .A2({ S11300 }),
  .A3({ S11324 }),
  .ZN({ S11346 })
);
NAND2_X1 #() 
NAND2_X1_1060_ (
  .A1({ S11345 }),
  .A2({ S11346 }),
  .ZN({ S11347 })
);
NAND2_X1 #() 
NAND2_X1_1061_ (
  .A1({ S11347 }),
  .A2({ S24 }),
  .ZN({ S11348 })
);
NAND4_X1 #() 
NAND4_X1_146_ (
  .A1({ S9781 }),
  .A2({ S9581 }),
  .A3({ S9614 }),
  .A4({ S9786 }),
  .ZN({ S11350 })
);
NAND2_X1 #() 
NAND2_X1_1062_ (
  .A1({ S25957[387] }),
  .A2({ S11350 }),
  .ZN({ S11351 })
);
OAI21_X1 #() 
OAI21_X1_608_ (
  .A({ S11348 }),
  .B1({ S11344 }),
  .B2({ S11351 }),
  .ZN({ S11352 })
);
INV_X1 #() 
INV_X1_345_ (
  .A({ S11350 }),
  .ZN({ S11353 })
);
NAND4_X1 #() 
NAND4_X1_147_ (
  .A1({ S25957[384] }),
  .A2({ S11324 }),
  .A3({ S9781 }),
  .A4({ S9786 }),
  .ZN({ S11354 })
);
NAND3_X1 #() 
NAND3_X1_1246_ (
  .A1({ S25957[387] }),
  .A2({ S11301 }),
  .A3({ S11354 }),
  .ZN({ S11355 })
);
OAI211_X1 #() 
OAI211_X1_390_ (
  .A({ S11355 }),
  .B({ S25957[388] }),
  .C1({ S11353 }),
  .C2({ S11323 }),
  .ZN({ S11356 })
);
OAI211_X1 #() 
OAI211_X1_391_ (
  .A({ S25957[389] }),
  .B({ S11356 }),
  .C1({ S11352 }),
  .C2({ S25957[388] }),
  .ZN({ S11357 })
);
OAI21_X1 #() 
OAI21_X1_609_ (
  .A({ S11357 }),
  .B1({ S11343 }),
  .B2({ S25957[389] }),
  .ZN({ S11358 })
);
NAND2_X1 #() 
NAND2_X1_1063_ (
  .A1({ S11358 }),
  .A2({ S25957[390] }),
  .ZN({ S11359 })
);
OAI211_X1 #() 
OAI211_X1_392_ (
  .A({ S11359 }),
  .B({ S25957[391] }),
  .C1({ S11329 }),
  .C2({ S25957[390] }),
  .ZN({ S11361 })
);
NAND2_X1 #() 
NAND2_X1_1064_ (
  .A1({ S9184 }),
  .A2({ S9182 }),
  .ZN({ S11362 })
);
NAND3_X1 #() 
NAND3_X1_1247_ (
  .A1({ S11324 }),
  .A2({ S9781 }),
  .A3({ S9786 }),
  .ZN({ S11363 })
);
NAND2_X1 #() 
NAND2_X1_1065_ (
  .A1({ S11363 }),
  .A2({ S11350 }),
  .ZN({ S11364 })
);
NAND2_X1 #() 
NAND2_X1_1066_ (
  .A1({ S11297 }),
  .A2({ S34 }),
  .ZN({ S11365 })
);
AOI21_X1 #() 
AOI21_X1_671_ (
  .A({ S25957[388] }),
  .B1({ S11365 }),
  .B2({ S25957[387] }),
  .ZN({ S11366 })
);
OAI21_X1 #() 
OAI21_X1_610_ (
  .A({ S11366 }),
  .B1({ S11364 }),
  .B2({ S11308 }),
  .ZN({ S11367 })
);
NAND2_X1 #() 
NAND2_X1_1067_ (
  .A1({ S25957[386] }),
  .A2({ S25957[384] }),
  .ZN({ S11368 })
);
NAND2_X1 #() 
NAND2_X1_1068_ (
  .A1({ S25957[387] }),
  .A2({ S11368 }),
  .ZN({ S11369 })
);
OAI22_X1 #() 
OAI22_X1_31_ (
  .A1({ S11369 }),
  .A2({ S11306 }),
  .B1({ S11300 }),
  .B2({ S25957[387] }),
  .ZN({ S11370 })
);
AOI21_X1 #() 
AOI21_X1_672_ (
  .A({ S11293 }),
  .B1({ S11370 }),
  .B2({ S25957[388] }),
  .ZN({ S11372 })
);
NAND2_X1 #() 
NAND2_X1_1069_ (
  .A1({ S11292 }),
  .A2({ S25957[386] }),
  .ZN({ S11373 })
);
NOR2_X1 #() 
NOR2_X1_252_ (
  .A1({ S11313 }),
  .A2({ S25957[387] }),
  .ZN({ S11374 })
);
INV_X1 #() 
INV_X1_346_ (
  .A({ S11374 }),
  .ZN({ S11375 })
);
OAI21_X1 #() 
OAI21_X1_611_ (
  .A({ S11375 }),
  .B1({ S24 }),
  .B2({ S11373 }),
  .ZN({ S11376 })
);
NAND3_X1 #() 
NAND3_X1_1248_ (
  .A1({ S34 }),
  .A2({ S11292 }),
  .A3({ S25957[386] }),
  .ZN({ S11377 })
);
AOI22_X1 #() 
AOI22_X1_142_ (
  .A1({ S33 }),
  .A2({ S11298 }),
  .B1({ S9524 }),
  .B2({ S9515 }),
  .ZN({ S11378 })
);
NAND3_X1 #() 
NAND3_X1_1249_ (
  .A1({ S25957[386] }),
  .A2({ S25957[385] }),
  .A3({ S11300 }),
  .ZN({ S11379 })
);
AOI22_X1 #() 
AOI22_X1_143_ (
  .A1({ S11378 }),
  .A2({ S11377 }),
  .B1({ S25957[387] }),
  .B2({ S11379 }),
  .ZN({ S11380 })
);
NAND2_X1 #() 
NAND2_X1_1070_ (
  .A1({ S11380 }),
  .A2({ S25957[388] }),
  .ZN({ S11381 })
);
OAI21_X1 #() 
OAI21_X1_612_ (
  .A({ S11381 }),
  .B1({ S11376 }),
  .B2({ S25957[388] }),
  .ZN({ S11383 })
);
AOI22_X1 #() 
AOI22_X1_144_ (
  .A1({ S11383 }),
  .A2({ S11293 }),
  .B1({ S11367 }),
  .B2({ S11372 }),
  .ZN({ S11384 })
);
NAND3_X1 #() 
NAND3_X1_1250_ (
  .A1({ S11379 }),
  .A2({ S24 }),
  .A3({ S11350 }),
  .ZN({ S11385 })
);
OAI211_X1 #() 
OAI211_X1_393_ (
  .A({ S11385 }),
  .B({ S25957[388] }),
  .C1({ S11347 }),
  .C2({ S24 }),
  .ZN({ S11386 })
);
INV_X1 #() 
INV_X1_347_ (
  .A({ S11373 }),
  .ZN({ S11387 })
);
OAI21_X1 #() 
OAI21_X1_613_ (
  .A({ S11324 }),
  .B1({ S11295 }),
  .B2({ S11296 }),
  .ZN({ S11388 })
);
NAND4_X1 #() 
NAND4_X1_148_ (
  .A1({ S9781 }),
  .A2({ S9786 }),
  .A3({ S11290 }),
  .A4({ S11291 }),
  .ZN({ S11389 })
);
NAND3_X1 #() 
NAND3_X1_1251_ (
  .A1({ S11388 }),
  .A2({ S11350 }),
  .A3({ S11389 }),
  .ZN({ S11390 })
);
NAND2_X1 #() 
NAND2_X1_1071_ (
  .A1({ S11390 }),
  .A2({ S25957[387] }),
  .ZN({ S11391 })
);
INV_X1 #() 
INV_X1_348_ (
  .A({ S11391 }),
  .ZN({ S11392 })
);
AOI21_X1 #() 
AOI21_X1_673_ (
  .A({ S11392 }),
  .B1({ S11387 }),
  .B2({ S24 }),
  .ZN({ S11394 })
);
OAI21_X1 #() 
OAI21_X1_614_ (
  .A({ S11386 }),
  .B1({ S11394 }),
  .B2({ S25957[388] }),
  .ZN({ S11395 })
);
OAI21_X1 #() 
OAI21_X1_615_ (
  .A({ S25957[390] }),
  .B1({ S11395 }),
  .B2({ S11293 }),
  .ZN({ S11396 })
);
AOI22_X1 #() 
AOI22_X1_145_ (
  .A1({ S11298 }),
  .A2({ S25957[384] }),
  .B1({ S9515 }),
  .B2({ S9524 }),
  .ZN({ S11397 })
);
NAND3_X1 #() 
NAND3_X1_1252_ (
  .A1({ S11311 }),
  .A2({ S11312 }),
  .A3({ S11298 }),
  .ZN({ S11398 })
);
AOI21_X1 #() 
AOI21_X1_674_ (
  .A({ S24 }),
  .B1({ S11398 }),
  .B2({ S11373 }),
  .ZN({ S11399 })
);
AOI21_X1 #() 
AOI21_X1_675_ (
  .A({ S11399 }),
  .B1({ S11397 }),
  .B2({ S11377 }),
  .ZN({ S11400 })
);
NAND3_X1 #() 
NAND3_X1_1253_ (
  .A1({ S25957[387] }),
  .A2({ S11389 }),
  .A3({ S11368 }),
  .ZN({ S11401 })
);
NAND2_X1 #() 
NAND2_X1_1072_ (
  .A1({ S11311 }),
  .A2({ S11298 }),
  .ZN({ S11402 })
);
NAND2_X1 #() 
NAND2_X1_1073_ (
  .A1({ S11402 }),
  .A2({ S11373 }),
  .ZN({ S11403 })
);
AOI21_X1 #() 
AOI21_X1_676_ (
  .A({ S25957[388] }),
  .B1({ S11403 }),
  .B2({ S24 }),
  .ZN({ S11405 })
);
AOI22_X1 #() 
AOI22_X1_146_ (
  .A1({ S11400 }),
  .A2({ S25957[388] }),
  .B1({ S11401 }),
  .B2({ S11405 }),
  .ZN({ S11406 })
);
NOR2_X1 #() 
NOR2_X1_253_ (
  .A1({ S11406 }),
  .A2({ S25957[389] }),
  .ZN({ S11407 })
);
OAI221_X1 #() 
OAI221_X1_22_ (
  .A({ S11362 }),
  .B1({ S11384 }),
  .B2({ S25957[390] }),
  .C1({ S11396 }),
  .C2({ S11407 }),
  .ZN({ S11408 })
);
NAND2_X1 #() 
NAND2_X1_1074_ (
  .A1({ S11408 }),
  .A2({ S11361 }),
  .ZN({ S11409 })
);
NAND2_X1 #() 
NAND2_X1_1075_ (
  .A1({ S11409 }),
  .A2({ S25957[495] }),
  .ZN({ S11410 })
);
NAND3_X1 #() 
NAND3_X1_1254_ (
  .A1({ S11408 }),
  .A2({ S8421 }),
  .A3({ S11361 }),
  .ZN({ S11411 })
);
NAND2_X1 #() 
NAND2_X1_1076_ (
  .A1({ S11410 }),
  .A2({ S11411 }),
  .ZN({ S11412 })
);
NOR2_X1 #() 
NOR2_X1_254_ (
  .A1({ S11412 }),
  .A2({ S5582 }),
  .ZN({ S11413 })
);
INV_X1 #() 
INV_X1_349_ (
  .A({ S11412 }),
  .ZN({ S25957[367] })
);
NOR2_X1 #() 
NOR2_X1_255_ (
  .A1({ S25957[367] }),
  .A2({ S25957[559] }),
  .ZN({ S11415 })
);
OAI21_X1 #() 
OAI21_X1_616_ (
  .A({ S25957[399] }),
  .B1({ S11415 }),
  .B2({ S11413 }),
  .ZN({ S11416 })
);
NOR2_X1 #() 
NOR2_X1_256_ (
  .A1({ S11415 }),
  .A2({ S11413 }),
  .ZN({ S25957[303] })
);
NAND2_X1 #() 
NAND2_X1_1077_ (
  .A1({ S25957[303] }),
  .A2({ S10598 }),
  .ZN({ S11417 })
);
NAND2_X1 #() 
NAND2_X1_1078_ (
  .A1({ S11417 }),
  .A2({ S11416 }),
  .ZN({ S25957[271] })
);
XNOR2_X1 #() 
XNOR2_X1_36_ (
  .A({ S8504 }),
  .B({ S25957[558] }),
  .ZN({ S25957[430] })
);
XOR2_X1 #() 
XOR2_X1_21_ (
  .A({ S8498 }),
  .B({ S25957[622] }),
  .Z({ S25957[494] })
);
AND2_X1 #() 
AND2_X1_65_ (
  .A1({ S9269 }),
  .A2({ S9265 }),
  .ZN({ S11418 })
);
NAND2_X1 #() 
NAND2_X1_1079_ (
  .A1({ S11292 }),
  .A2({ S11298 }),
  .ZN({ S11419 })
);
NOR2_X1 #() 
NOR2_X1_257_ (
  .A1({ S24 }),
  .A2({ S11318 }),
  .ZN({ S11420 })
);
NAND2_X1 #() 
NAND2_X1_1080_ (
  .A1({ S11420 }),
  .A2({ S11419 }),
  .ZN({ S11422 })
);
NAND2_X1 #() 
NAND2_X1_1081_ (
  .A1({ S11311 }),
  .A2({ S25957[386] }),
  .ZN({ S11423 })
);
AOI21_X1 #() 
AOI21_X1_677_ (
  .A({ S24 }),
  .B1({ S11423 }),
  .B2({ S11309 }),
  .ZN({ S11424 })
);
AOI211_X1 #() 
AOI211_X1_14_ (
  .A({ S11332 }),
  .B({ S11424 }),
  .C1({ S11303 }),
  .C2({ S11398 }),
  .ZN({ S11425 })
);
AOI21_X1 #() 
AOI21_X1_678_ (
  .A({ S11425 }),
  .B1({ S11422 }),
  .B2({ S11405 }),
  .ZN({ S11426 })
);
NAND2_X1 #() 
NAND2_X1_1082_ (
  .A1({ S34 }),
  .A2({ S11298 }),
  .ZN({ S11427 })
);
NAND3_X1 #() 
NAND3_X1_1255_ (
  .A1({ S25957[387] }),
  .A2({ S11423 }),
  .A3({ S11427 }),
  .ZN({ S11428 })
);
OAI211_X1 #() 
OAI211_X1_394_ (
  .A({ S11428 }),
  .B({ S25957[388] }),
  .C1({ S25957[387] }),
  .C2({ S11337 }),
  .ZN({ S11429 })
);
OAI21_X1 #() 
OAI21_X1_617_ (
  .A({ S11323 }),
  .B1({ S11334 }),
  .B2({ S33 }),
  .ZN({ S11430 })
);
NAND2_X1 #() 
NAND2_X1_1083_ (
  .A1({ S11430 }),
  .A2({ S11332 }),
  .ZN({ S11431 })
);
AOI21_X1 #() 
AOI21_X1_679_ (
  .A({ S11293 }),
  .B1({ S11431 }),
  .B2({ S11429 }),
  .ZN({ S11433 })
);
AOI21_X1 #() 
AOI21_X1_680_ (
  .A({ S11433 }),
  .B1({ S11426 }),
  .B2({ S11293 }),
  .ZN({ S11434 })
);
NAND4_X1 #() 
NAND4_X1_149_ (
  .A1({ S9515 }),
  .A2({ S25957[386] }),
  .A3({ S25957[385] }),
  .A4({ S9524 }),
  .ZN({ S11435 })
);
NOR2_X1 #() 
NOR2_X1_258_ (
  .A1({ S25957[384] }),
  .A2({ S11324 }),
  .ZN({ S11436 })
);
NAND3_X1 #() 
NAND3_X1_1256_ (
  .A1({ S24 }),
  .A2({ S11436 }),
  .A3({ S11298 }),
  .ZN({ S11437 })
);
NAND2_X1 #() 
NAND2_X1_1084_ (
  .A1({ S11437 }),
  .A2({ S11435 }),
  .ZN({ S11438 })
);
OAI21_X1 #() 
OAI21_X1_618_ (
  .A({ S25957[388] }),
  .B1({ S11438 }),
  .B2({ S11374 }),
  .ZN({ S11439 })
);
OAI21_X1 #() 
OAI21_X1_619_ (
  .A({ S11388 }),
  .B1({ S25957[386] }),
  .B2({ S11312 }),
  .ZN({ S11440 })
);
AOI21_X1 #() 
AOI21_X1_681_ (
  .A({ S25957[388] }),
  .B1({ S11397 }),
  .B2({ S11344 }),
  .ZN({ S11441 })
);
OAI21_X1 #() 
OAI21_X1_620_ (
  .A({ S11441 }),
  .B1({ S24 }),
  .B2({ S11440 }),
  .ZN({ S11442 })
);
NAND3_X1 #() 
NAND3_X1_1257_ (
  .A1({ S11442 }),
  .A2({ S11439 }),
  .A3({ S25957[389] }),
  .ZN({ S11444 })
);
OAI21_X1 #() 
OAI21_X1_621_ (
  .A({ S11309 }),
  .B1({ S11312 }),
  .B2({ S11298 }),
  .ZN({ S11445 })
);
AOI22_X1 #() 
AOI22_X1_147_ (
  .A1({ S11303 }),
  .A2({ S11398 }),
  .B1({ S11445 }),
  .B2({ S25957[387] }),
  .ZN({ S11446 })
);
OAI211_X1 #() 
OAI211_X1_395_ (
  .A({ S11325 }),
  .B({ S25957[388] }),
  .C1({ S25957[387] }),
  .C2({ S11402 }),
  .ZN({ S11447 })
);
OAI211_X1 #() 
OAI211_X1_396_ (
  .A({ S11447 }),
  .B({ S11293 }),
  .C1({ S11446 }),
  .C2({ S25957[388] }),
  .ZN({ S11448 })
);
NAND3_X1 #() 
NAND3_X1_1258_ (
  .A1({ S11444 }),
  .A2({ S11448 }),
  .A3({ S11418 }),
  .ZN({ S11449 })
);
OAI21_X1 #() 
OAI21_X1_622_ (
  .A({ S11449 }),
  .B1({ S11434 }),
  .B2({ S11418 }),
  .ZN({ S11450 })
);
NAND2_X1 #() 
NAND2_X1_1085_ (
  .A1({ S11450 }),
  .A2({ S25957[391] }),
  .ZN({ S11451 })
);
NAND2_X1 #() 
NAND2_X1_1086_ (
  .A1({ S11312 }),
  .A2({ S11298 }),
  .ZN({ S11452 })
);
AOI21_X1 #() 
AOI21_X1_682_ (
  .A({ S24 }),
  .B1({ S11452 }),
  .B2({ S11379 }),
  .ZN({ S11453 })
);
NAND2_X1 #() 
NAND2_X1_1087_ (
  .A1({ S11453 }),
  .A2({ S11332 }),
  .ZN({ S11455 })
);
NOR2_X1 #() 
NOR2_X1_259_ (
  .A1({ S25957[387] }),
  .A2({ S11354 }),
  .ZN({ S11456 })
);
OAI21_X1 #() 
OAI21_X1_623_ (
  .A({ S25957[388] }),
  .B1({ S11392 }),
  .B2({ S11456 }),
  .ZN({ S11457 })
);
AOI21_X1 #() 
AOI21_X1_683_ (
  .A({ S25957[389] }),
  .B1({ S11457 }),
  .B2({ S11455 }),
  .ZN({ S11458 })
);
AOI22_X1 #() 
AOI22_X1_148_ (
  .A1({ S11333 }),
  .A2({ S11389 }),
  .B1({ S24 }),
  .B2({ S11390 }),
  .ZN({ S11459 })
);
NAND2_X1 #() 
NAND2_X1_1088_ (
  .A1({ S25957[387] }),
  .A2({ S11346 }),
  .ZN({ S11460 })
);
NOR2_X1 #() 
NOR2_X1_260_ (
  .A1({ S11460 }),
  .A2({ S33 }),
  .ZN({ S11461 })
);
NOR3_X1 #() 
NOR3_X1_34_ (
  .A1({ S11461 }),
  .A2({ S11397 }),
  .A3({ S11332 }),
  .ZN({ S11462 })
);
AOI211_X1 #() 
AOI211_X1_15_ (
  .A({ S11293 }),
  .B({ S11462 }),
  .C1({ S11332 }),
  .C2({ S11459 }),
  .ZN({ S11463 })
);
NOR2_X1 #() 
NOR2_X1_261_ (
  .A1({ S11463 }),
  .A2({ S11458 }),
  .ZN({ S11464 })
);
AND2_X1 #() 
AND2_X1_66_ (
  .A1({ S11377 }),
  .A2({ S24 }),
  .ZN({ S11466 })
);
NOR3_X1 #() 
NOR3_X1_35_ (
  .A1({ S11466 }),
  .A2({ S11424 }),
  .A3({ S25957[388] }),
  .ZN({ S11467 })
);
NAND3_X1 #() 
NAND3_X1_1259_ (
  .A1({ S25957[386] }),
  .A2({ S25957[385] }),
  .A3({ S25957[384] }),
  .ZN({ S11468 })
);
AOI21_X1 #() 
AOI21_X1_684_ (
  .A({ S25957[387] }),
  .B1({ S11350 }),
  .B2({ S11468 }),
  .ZN({ S11469 })
);
NAND2_X1 #() 
NAND2_X1_1089_ (
  .A1({ S11309 }),
  .A2({ S34 }),
  .ZN({ S11470 })
);
OAI21_X1 #() 
OAI21_X1_624_ (
  .A({ S25957[388] }),
  .B1({ S11470 }),
  .B2({ S24 }),
  .ZN({ S11471 })
);
INV_X1 #() 
INV_X1_350_ (
  .A({ S11323 }),
  .ZN({ S11472 })
);
OAI211_X1 #() 
OAI211_X1_397_ (
  .A({ S11309 }),
  .B({ S11332 }),
  .C1({ S11472 }),
  .C2({ S11420 }),
  .ZN({ S11473 })
);
OAI21_X1 #() 
OAI21_X1_625_ (
  .A({ S11473 }),
  .B1({ S11469 }),
  .B2({ S11471 }),
  .ZN({ S11474 })
);
NAND2_X1 #() 
NAND2_X1_1090_ (
  .A1({ S11474 }),
  .A2({ S25957[389] }),
  .ZN({ S11475 })
);
NAND3_X1 #() 
NAND3_X1_1260_ (
  .A1({ S24 }),
  .A2({ S11300 }),
  .A3({ S11363 }),
  .ZN({ S11477 })
);
INV_X1 #() 
INV_X1_351_ (
  .A({ S11389 }),
  .ZN({ S11478 })
);
NAND2_X1 #() 
NAND2_X1_1091_ (
  .A1({ S25957[387] }),
  .A2({ S11478 }),
  .ZN({ S11479 })
);
NAND3_X1 #() 
NAND3_X1_1261_ (
  .A1({ S11479 }),
  .A2({ S11477 }),
  .A3({ S25957[388] }),
  .ZN({ S11480 })
);
NAND2_X1 #() 
NAND2_X1_1092_ (
  .A1({ S11480 }),
  .A2({ S11293 }),
  .ZN({ S11481 })
);
OAI21_X1 #() 
OAI21_X1_626_ (
  .A({ S11475 }),
  .B1({ S11467 }),
  .B2({ S11481 }),
  .ZN({ S11482 })
);
NAND2_X1 #() 
NAND2_X1_1093_ (
  .A1({ S11482 }),
  .A2({ S25957[390] }),
  .ZN({ S11483 })
);
OAI21_X1 #() 
OAI21_X1_627_ (
  .A({ S11483 }),
  .B1({ S11464 }),
  .B2({ S25957[390] }),
  .ZN({ S11484 })
);
NAND2_X1 #() 
NAND2_X1_1094_ (
  .A1({ S11484 }),
  .A2({ S11362 }),
  .ZN({ S11485 })
);
NAND3_X1 #() 
NAND3_X1_1262_ (
  .A1({ S11485 }),
  .A2({ S11451 }),
  .A3({ S25957[494] }),
  .ZN({ S11486 })
);
INV_X1 #() 
INV_X1_352_ (
  .A({ S25957[494] }),
  .ZN({ S11488 })
);
OAI211_X1 #() 
OAI211_X1_398_ (
  .A({ S11362 }),
  .B({ S11483 }),
  .C1({ S11464 }),
  .C2({ S25957[390] }),
  .ZN({ S11489 })
);
OAI211_X1 #() 
OAI211_X1_399_ (
  .A({ S11489 }),
  .B({ S11488 }),
  .C1({ S11362 }),
  .C2({ S11450 }),
  .ZN({ S11490 })
);
NAND3_X1 #() 
NAND3_X1_1263_ (
  .A1({ S11486 }),
  .A2({ S11490 }),
  .A3({ S25957[462] }),
  .ZN({ S11491 })
);
NAND3_X1 #() 
NAND3_X1_1264_ (
  .A1({ S11485 }),
  .A2({ S11451 }),
  .A3({ S11488 }),
  .ZN({ S11492 })
);
OAI211_X1 #() 
OAI211_X1_400_ (
  .A({ S11489 }),
  .B({ S25957[494] }),
  .C1({ S11362 }),
  .C2({ S11450 }),
  .ZN({ S11493 })
);
NAND3_X1 #() 
NAND3_X1_1265_ (
  .A1({ S11492 }),
  .A2({ S11493 }),
  .A3({ S8504 }),
  .ZN({ S11494 })
);
NAND3_X1 #() 
NAND3_X1_1266_ (
  .A1({ S11491 }),
  .A2({ S11494 }),
  .A3({ S25957[430] }),
  .ZN({ S11495 })
);
INV_X1 #() 
INV_X1_353_ (
  .A({ S25957[430] }),
  .ZN({ S11496 })
);
NAND3_X1 #() 
NAND3_X1_1267_ (
  .A1({ S11492 }),
  .A2({ S11493 }),
  .A3({ S25957[462] }),
  .ZN({ S11497 })
);
NAND3_X1 #() 
NAND3_X1_1268_ (
  .A1({ S11486 }),
  .A2({ S11490 }),
  .A3({ S8504 }),
  .ZN({ S11499 })
);
NAND3_X1 #() 
NAND3_X1_1269_ (
  .A1({ S11497 }),
  .A2({ S11499 }),
  .A3({ S11496 }),
  .ZN({ S11500 })
);
NAND3_X1 #() 
NAND3_X1_1270_ (
  .A1({ S11495 }),
  .A2({ S11500 }),
  .A3({ S8507 }),
  .ZN({ S11501 })
);
NAND3_X1 #() 
NAND3_X1_1271_ (
  .A1({ S11497 }),
  .A2({ S11499 }),
  .A3({ S25957[430] }),
  .ZN({ S11502 })
);
NAND3_X1 #() 
NAND3_X1_1272_ (
  .A1({ S11491 }),
  .A2({ S11494 }),
  .A3({ S11496 }),
  .ZN({ S11503 })
);
NAND3_X1 #() 
NAND3_X1_1273_ (
  .A1({ S11502 }),
  .A2({ S11503 }),
  .A3({ S25957[398] }),
  .ZN({ S11504 })
);
NAND2_X1 #() 
NAND2_X1_1095_ (
  .A1({ S11501 }),
  .A2({ S11504 }),
  .ZN({ S25957[270] })
);
NOR2_X1 #() 
NOR2_X1_262_ (
  .A1({ S8579 }),
  .A2({ S8583 }),
  .ZN({ S11505 })
);
XNOR2_X1 #() 
XNOR2_X1_37_ (
  .A({ S8508 }),
  .B({ S25957[717] }),
  .ZN({ S25957[589] })
);
NAND2_X1 #() 
NAND2_X1_1096_ (
  .A1({ S11363 }),
  .A2({ S11309 }),
  .ZN({ S11506 })
);
NAND2_X1 #() 
NAND2_X1_1097_ (
  .A1({ S11506 }),
  .A2({ S25957[387] }),
  .ZN({ S11508 })
);
NAND2_X1 #() 
NAND2_X1_1098_ (
  .A1({ S11312 }),
  .A2({ S25957[386] }),
  .ZN({ S11509 })
);
NAND2_X1 #() 
NAND2_X1_1099_ (
  .A1({ S11509 }),
  .A2({ S24 }),
  .ZN({ S11510 })
);
NAND3_X1 #() 
NAND3_X1_1274_ (
  .A1({ S11508 }),
  .A2({ S25957[388] }),
  .A3({ S11510 }),
  .ZN({ S11511 })
);
OAI21_X1 #() 
OAI21_X1_628_ (
  .A({ S11332 }),
  .B1({ S11374 }),
  .B2({ S11424 }),
  .ZN({ S11512 })
);
NAND2_X1 #() 
NAND2_X1_1100_ (
  .A1({ S11512 }),
  .A2({ S11511 }),
  .ZN({ S11513 })
);
NAND2_X1 #() 
NAND2_X1_1101_ (
  .A1({ S11513 }),
  .A2({ S11293 }),
  .ZN({ S11514 })
);
AOI21_X1 #() 
AOI21_X1_685_ (
  .A({ S24 }),
  .B1({ S11419 }),
  .B2({ S11509 }),
  .ZN({ S11515 })
);
AOI21_X1 #() 
AOI21_X1_686_ (
  .A({ S25957[387] }),
  .B1({ S11324 }),
  .B2({ S11368 }),
  .ZN({ S11516 })
);
OAI21_X1 #() 
OAI21_X1_629_ (
  .A({ S11332 }),
  .B1({ S11516 }),
  .B2({ S11515 }),
  .ZN({ S11517 })
);
INV_X1 #() 
INV_X1_354_ (
  .A({ S11402 }),
  .ZN({ S11519 })
);
NAND3_X1 #() 
NAND3_X1_1275_ (
  .A1({ S9515 }),
  .A2({ S9524 }),
  .A3({ S11300 }),
  .ZN({ S11520 })
);
OAI221_X1 #() 
OAI221_X1_23_ (
  .A({ S25957[388] }),
  .B1({ S11306 }),
  .B2({ S11520 }),
  .C1({ S11519 }),
  .C2({ S11335 }),
  .ZN({ S11521 })
);
NAND2_X1 #() 
NAND2_X1_1102_ (
  .A1({ S11517 }),
  .A2({ S11521 }),
  .ZN({ S11522 })
);
NAND2_X1 #() 
NAND2_X1_1103_ (
  .A1({ S11522 }),
  .A2({ S25957[389] }),
  .ZN({ S11523 })
);
AOI21_X1 #() 
AOI21_X1_687_ (
  .A({ S11418 }),
  .B1({ S11523 }),
  .B2({ S11514 }),
  .ZN({ S11524 })
);
AOI21_X1 #() 
AOI21_X1_688_ (
  .A({ S25957[386] }),
  .B1({ S11311 }),
  .B2({ S11312 }),
  .ZN({ S11525 })
);
NAND2_X1 #() 
NAND2_X1_1104_ (
  .A1({ S11525 }),
  .A2({ S25957[387] }),
  .ZN({ S11526 })
);
AOI21_X1 #() 
AOI21_X1_689_ (
  .A({ S25957[385] }),
  .B1({ S11298 }),
  .B2({ S25957[384] }),
  .ZN({ S11527 })
);
AOI21_X1 #() 
AOI21_X1_690_ (
  .A({ S11332 }),
  .B1({ S11527 }),
  .B2({ S24 }),
  .ZN({ S11528 })
);
NAND2_X1 #() 
NAND2_X1_1105_ (
  .A1({ S11528 }),
  .A2({ S11526 }),
  .ZN({ S11529 })
);
AOI21_X1 #() 
AOI21_X1_691_ (
  .A({ S24 }),
  .B1({ S11377 }),
  .B2({ S11319 }),
  .ZN({ S11530 })
);
OAI21_X1 #() 
OAI21_X1_630_ (
  .A({ S11332 }),
  .B1({ S11530 }),
  .B2({ S11378 }),
  .ZN({ S11531 })
);
AOI21_X1 #() 
AOI21_X1_692_ (
  .A({ S25957[389] }),
  .B1({ S11531 }),
  .B2({ S11529 }),
  .ZN({ S11532 })
);
INV_X1 #() 
INV_X1_355_ (
  .A({ S11532 }),
  .ZN({ S11533 })
);
OAI21_X1 #() 
OAI21_X1_631_ (
  .A({ S11350 }),
  .B1({ S9526 }),
  .B2({ S9525 }),
  .ZN({ S11534 })
);
OAI221_X1 #() 
OAI221_X1_24_ (
  .A({ S25957[388] }),
  .B1({ S11534 }),
  .B2({ S33 }),
  .C1({ S11403 }),
  .C2({ S24 }),
  .ZN({ S11535 })
);
NAND2_X1 #() 
NAND2_X1_1106_ (
  .A1({ S25957[387] }),
  .A2({ S11324 }),
  .ZN({ S11536 })
);
NAND3_X1 #() 
NAND3_X1_1276_ (
  .A1({ S24 }),
  .A2({ S11363 }),
  .A3({ S11312 }),
  .ZN({ S11537 })
);
NAND3_X1 #() 
NAND3_X1_1277_ (
  .A1({ S11536 }),
  .A2({ S11537 }),
  .A3({ S11332 }),
  .ZN({ S11538 })
);
NAND3_X1 #() 
NAND3_X1_1278_ (
  .A1({ S11535 }),
  .A2({ S25957[389] }),
  .A3({ S11538 }),
  .ZN({ S11540 })
);
AOI21_X1 #() 
AOI21_X1_693_ (
  .A({ S25957[390] }),
  .B1({ S11533 }),
  .B2({ S11540 }),
  .ZN({ S11541 })
);
OR3_X1 #() 
OR3_X1_4_ (
  .A1({ S11541 }),
  .A2({ S11524 }),
  .A3({ S11362 }),
  .ZN({ S11542 })
);
NAND4_X1 #() 
NAND4_X1_150_ (
  .A1({ S11311 }),
  .A2({ S11298 }),
  .A3({ S9515 }),
  .A4({ S9524 }),
  .ZN({ S11543 })
);
NAND2_X1 #() 
NAND2_X1_1107_ (
  .A1({ S11543 }),
  .A2({ S25957[388] }),
  .ZN({ S11544 })
);
NAND3_X1 #() 
NAND3_X1_1279_ (
  .A1({ S11309 }),
  .A2({ S9515 }),
  .A3({ S9524 }),
  .ZN({ S11545 })
);
NOR2_X1 #() 
NOR2_X1_263_ (
  .A1({ S11387 }),
  .A2({ S11545 }),
  .ZN({ S11546 })
);
NAND3_X1 #() 
NAND3_X1_1280_ (
  .A1({ S11301 }),
  .A2({ S11363 }),
  .A3({ S11309 }),
  .ZN({ S11547 })
);
AOI21_X1 #() 
AOI21_X1_694_ (
  .A({ S11546 }),
  .B1({ S24 }),
  .B2({ S11547 }),
  .ZN({ S11548 })
);
NAND2_X1 #() 
NAND2_X1_1108_ (
  .A1({ S11468 }),
  .A2({ S11350 }),
  .ZN({ S11549 })
);
NOR3_X1 #() 
NOR3_X1_36_ (
  .A1({ S11549 }),
  .A2({ S11306 }),
  .A3({ S25957[387] }),
  .ZN({ S11551 })
);
OAI221_X1 #() 
OAI221_X1_25_ (
  .A({ S11293 }),
  .B1({ S11551 }),
  .B2({ S11544 }),
  .C1({ S11548 }),
  .C2({ S25957[388] }),
  .ZN({ S11552 })
);
NAND2_X1 #() 
NAND2_X1_1109_ (
  .A1({ S11436 }),
  .A2({ S11298 }),
  .ZN({ S11553 })
);
NAND3_X1 #() 
NAND3_X1_1281_ (
  .A1({ S11553 }),
  .A2({ S25957[387] }),
  .A3({ S11313 }),
  .ZN({ S11554 })
);
OAI21_X1 #() 
OAI21_X1_632_ (
  .A({ S11554 }),
  .B1({ S25957[387] }),
  .B2({ S11390 }),
  .ZN({ S11555 })
);
INV_X1 #() 
INV_X1_356_ (
  .A({ S11520 }),
  .ZN({ S11556 })
);
NAND3_X1 #() 
NAND3_X1_1282_ (
  .A1({ S24 }),
  .A2({ S11309 }),
  .A3({ S11312 }),
  .ZN({ S11557 })
);
INV_X1 #() 
INV_X1_357_ (
  .A({ S11557 }),
  .ZN({ S11558 })
);
OAI21_X1 #() 
OAI21_X1_633_ (
  .A({ S11332 }),
  .B1({ S11558 }),
  .B2({ S11556 }),
  .ZN({ S11559 })
);
OAI211_X1 #() 
OAI211_X1_401_ (
  .A({ S25957[389] }),
  .B({ S11559 }),
  .C1({ S11555 }),
  .C2({ S11332 }),
  .ZN({ S11560 })
);
NAND3_X1 #() 
NAND3_X1_1283_ (
  .A1({ S11552 }),
  .A2({ S25957[390] }),
  .A3({ S11560 }),
  .ZN({ S11561 })
);
AOI22_X1 #() 
AOI22_X1_149_ (
  .A1({ S11472 }),
  .A2({ S11353 }),
  .B1({ S25957[387] }),
  .B2({ S11419 }),
  .ZN({ S11562 })
);
NAND2_X1 #() 
NAND2_X1_1110_ (
  .A1({ S11309 }),
  .A2({ S25957[385] }),
  .ZN({ S11563 })
);
OAI221_X1 #() 
OAI221_X1_26_ (
  .A({ S11332 }),
  .B1({ S11368 }),
  .B2({ S24 }),
  .C1({ S11302 }),
  .C2({ S11563 }),
  .ZN({ S11564 })
);
OAI211_X1 #() 
OAI211_X1_402_ (
  .A({ S11564 }),
  .B({ S25957[389] }),
  .C1({ S11562 }),
  .C2({ S11332 }),
  .ZN({ S11565 })
);
NAND3_X1 #() 
NAND3_X1_1284_ (
  .A1({ S11377 }),
  .A2({ S11419 }),
  .A3({ S24 }),
  .ZN({ S11566 })
);
INV_X1 #() 
INV_X1_358_ (
  .A({ S11566 }),
  .ZN({ S11567 })
);
AND2_X1 #() 
AND2_X1_67_ (
  .A1({ S11313 }),
  .A2({ S11354 }),
  .ZN({ S11568 })
);
AOI21_X1 #() 
AOI21_X1_695_ (
  .A({ S11567 }),
  .B1({ S25957[387] }),
  .B2({ S11568 }),
  .ZN({ S11569 })
);
OAI211_X1 #() 
OAI211_X1_403_ (
  .A({ S11340 }),
  .B({ S11332 }),
  .C1({ S11368 }),
  .C2({ S11323 }),
  .ZN({ S11570 })
);
OAI211_X1 #() 
OAI211_X1_404_ (
  .A({ S11293 }),
  .B({ S11570 }),
  .C1({ S11569 }),
  .C2({ S11332 }),
  .ZN({ S11571 })
);
NAND2_X1 #() 
NAND2_X1_1111_ (
  .A1({ S11571 }),
  .A2({ S11565 }),
  .ZN({ S11572 })
);
NAND2_X1 #() 
NAND2_X1_1112_ (
  .A1({ S11572 }),
  .A2({ S11418 }),
  .ZN({ S11573 })
);
NAND3_X1 #() 
NAND3_X1_1285_ (
  .A1({ S11573 }),
  .A2({ S11561 }),
  .A3({ S11362 }),
  .ZN({ S11574 })
);
NAND3_X1 #() 
NAND3_X1_1286_ (
  .A1({ S11542 }),
  .A2({ S11574 }),
  .A3({ S25957[589] }),
  .ZN({ S11575 })
);
INV_X1 #() 
INV_X1_359_ (
  .A({ S25957[589] }),
  .ZN({ S11576 })
);
OAI21_X1 #() 
OAI21_X1_634_ (
  .A({ S25957[391] }),
  .B1({ S11541 }),
  .B2({ S11524 }),
  .ZN({ S11577 })
);
NAND2_X1 #() 
NAND2_X1_1113_ (
  .A1({ S11573 }),
  .A2({ S11561 }),
  .ZN({ S11578 })
);
NAND2_X1 #() 
NAND2_X1_1114_ (
  .A1({ S11578 }),
  .A2({ S11362 }),
  .ZN({ S11579 })
);
NAND3_X1 #() 
NAND3_X1_1287_ (
  .A1({ S11579 }),
  .A2({ S11577 }),
  .A3({ S11576 }),
  .ZN({ S11580 })
);
AOI21_X1 #() 
AOI21_X1_696_ (
  .A({ S11505 }),
  .B1({ S11580 }),
  .B2({ S11575 }),
  .ZN({ S11582 })
);
NAND3_X1 #() 
NAND3_X1_1288_ (
  .A1({ S11580 }),
  .A2({ S11505 }),
  .A3({ S11575 }),
  .ZN({ S11583 })
);
INV_X1 #() 
INV_X1_360_ (
  .A({ S11583 }),
  .ZN({ S11584 })
);
OAI21_X1 #() 
OAI21_X1_635_ (
  .A({ S25957[397] }),
  .B1({ S11584 }),
  .B2({ S11582 }),
  .ZN({ S11585 })
);
INV_X1 #() 
INV_X1_361_ (
  .A({ S11505 }),
  .ZN({ S25957[429] })
);
INV_X1 #() 
INV_X1_362_ (
  .A({ S11575 }),
  .ZN({ S11586 })
);
AOI21_X1 #() 
AOI21_X1_697_ (
  .A({ S25957[589] }),
  .B1({ S11542 }),
  .B2({ S11574 }),
  .ZN({ S11587 })
);
OAI21_X1 #() 
OAI21_X1_636_ (
  .A({ S25957[429] }),
  .B1({ S11586 }),
  .B2({ S11587 }),
  .ZN({ S11588 })
);
NAND3_X1 #() 
NAND3_X1_1289_ (
  .A1({ S11588 }),
  .A2({ S10559 }),
  .A3({ S11583 }),
  .ZN({ S11589 })
);
NAND2_X1 #() 
NAND2_X1_1115_ (
  .A1({ S11585 }),
  .A2({ S11589 }),
  .ZN({ S25957[269] })
);
INV_X1 #() 
INV_X1_363_ (
  .A({ S10523 }),
  .ZN({ S25957[428] })
);
NAND2_X1 #() 
NAND2_X1_1116_ (
  .A1({ S5838 }),
  .A2({ S5836 }),
  .ZN({ S25957[620] })
);
XNOR2_X1 #() 
XNOR2_X1_38_ (
  .A({ S25957[620] }),
  .B({ S25957[716] }),
  .ZN({ S11591 })
);
INV_X1 #() 
INV_X1_364_ (
  .A({ S11591 }),
  .ZN({ S25957[588] })
);
NAND2_X1 #() 
NAND2_X1_1117_ (
  .A1({ S11346 }),
  .A2({ S24 }),
  .ZN({ S11592 })
);
INV_X1 #() 
INV_X1_365_ (
  .A({ S11592 }),
  .ZN({ S11593 })
);
NAND3_X1 #() 
NAND3_X1_1290_ (
  .A1({ S24 }),
  .A2({ S11300 }),
  .A3({ S11389 }),
  .ZN({ S11594 })
);
OAI211_X1 #() 
OAI211_X1_405_ (
  .A({ S11332 }),
  .B({ S11594 }),
  .C1({ S11369 }),
  .C2({ S11306 }),
  .ZN({ S11595 })
);
OAI211_X1 #() 
OAI211_X1_406_ (
  .A({ S11595 }),
  .B({ S25957[389] }),
  .C1({ S11544 }),
  .C2({ S11593 }),
  .ZN({ S11596 })
);
INV_X1 #() 
INV_X1_366_ (
  .A({ S11366 }),
  .ZN({ S11597 })
);
AOI22_X1 #() 
AOI22_X1_150_ (
  .A1({ S11368 }),
  .A2({ S11389 }),
  .B1({ S9524 }),
  .B2({ S9515 }),
  .ZN({ S11599 })
);
OAI211_X1 #() 
OAI211_X1_407_ (
  .A({ S25957[388] }),
  .B({ S11537 }),
  .C1({ S11536 }),
  .C2({ S11310 }),
  .ZN({ S11600 })
);
OAI21_X1 #() 
OAI21_X1_637_ (
  .A({ S11600 }),
  .B1({ S11597 }),
  .B2({ S11599 }),
  .ZN({ S11601 })
);
OAI21_X1 #() 
OAI21_X1_638_ (
  .A({ S11596 }),
  .B1({ S11601 }),
  .B2({ S25957[389] }),
  .ZN({ S11602 })
);
NAND2_X1 #() 
NAND2_X1_1118_ (
  .A1({ S11602 }),
  .A2({ S25957[390] }),
  .ZN({ S11603 })
);
AOI21_X1 #() 
AOI21_X1_698_ (
  .A({ S25957[387] }),
  .B1({ S11379 }),
  .B2({ S11452 }),
  .ZN({ S11604 })
);
NOR2_X1 #() 
NOR2_X1_264_ (
  .A1({ S11369 }),
  .A2({ S25957[385] }),
  .ZN({ S11605 })
);
OAI21_X1 #() 
OAI21_X1_639_ (
  .A({ S11332 }),
  .B1({ S11605 }),
  .B2({ S11604 }),
  .ZN({ S11606 })
);
AOI21_X1 #() 
AOI21_X1_699_ (
  .A({ S25957[387] }),
  .B1({ S11419 }),
  .B2({ S11509 }),
  .ZN({ S11607 })
);
AOI21_X1 #() 
AOI21_X1_700_ (
  .A({ S24 }),
  .B1({ S11379 }),
  .B2({ S11363 }),
  .ZN({ S11608 })
);
OAI21_X1 #() 
OAI21_X1_640_ (
  .A({ S25957[388] }),
  .B1({ S11607 }),
  .B2({ S11608 }),
  .ZN({ S11610 })
);
NAND3_X1 #() 
NAND3_X1_1291_ (
  .A1({ S11606 }),
  .A2({ S11610 }),
  .A3({ S11293 }),
  .ZN({ S11611 })
);
AOI21_X1 #() 
AOI21_X1_701_ (
  .A({ S25957[387] }),
  .B1({ S11398 }),
  .B2({ S11373 }),
  .ZN({ S11612 })
);
NAND4_X1 #() 
NAND4_X1_151_ (
  .A1({ S9515 }),
  .A2({ S25957[385] }),
  .A3({ S9524 }),
  .A4({ S11300 }),
  .ZN({ S11613 })
);
NAND2_X1 #() 
NAND2_X1_1119_ (
  .A1({ S11543 }),
  .A2({ S11613 }),
  .ZN({ S11614 })
);
OAI21_X1 #() 
OAI21_X1_641_ (
  .A({ S11332 }),
  .B1({ S11612 }),
  .B2({ S11614 }),
  .ZN({ S11615 })
);
OAI21_X1 #() 
OAI21_X1_642_ (
  .A({ S11339 }),
  .B1({ S25957[387] }),
  .B2({ S25957[386] }),
  .ZN({ S11616 })
);
NAND3_X1 #() 
NAND3_X1_1292_ (
  .A1({ S11616 }),
  .A2({ S25957[388] }),
  .A3({ S11553 }),
  .ZN({ S11617 })
);
NAND3_X1 #() 
NAND3_X1_1293_ (
  .A1({ S11615 }),
  .A2({ S25957[389] }),
  .A3({ S11617 }),
  .ZN({ S11618 })
);
NAND3_X1 #() 
NAND3_X1_1294_ (
  .A1({ S11611 }),
  .A2({ S11618 }),
  .A3({ S11418 }),
  .ZN({ S11619 })
);
NAND3_X1 #() 
NAND3_X1_1295_ (
  .A1({ S11603 }),
  .A2({ S25957[391] }),
  .A3({ S11619 }),
  .ZN({ S11621 })
);
NAND2_X1 #() 
NAND2_X1_1120_ (
  .A1({ S11537 }),
  .A2({ S25957[388] }),
  .ZN({ S11622 })
);
AOI21_X1 #() 
AOI21_X1_702_ (
  .A({ S24 }),
  .B1({ S11301 }),
  .B2({ S11354 }),
  .ZN({ S11623 })
);
NOR2_X1 #() 
NOR2_X1_265_ (
  .A1({ S11622 }),
  .A2({ S11623 }),
  .ZN({ S11624 })
);
NAND2_X1 #() 
NAND2_X1_1121_ (
  .A1({ S11309 }),
  .A2({ S11312 }),
  .ZN({ S11625 })
);
NAND2_X1 #() 
NAND2_X1_1122_ (
  .A1({ S25957[387] }),
  .A2({ S11625 }),
  .ZN({ S11626 })
);
NAND3_X1 #() 
NAND3_X1_1296_ (
  .A1({ S11427 }),
  .A2({ S11346 }),
  .A3({ S24 }),
  .ZN({ S11627 })
);
AOI21_X1 #() 
AOI21_X1_703_ (
  .A({ S25957[388] }),
  .B1({ S11627 }),
  .B2({ S11626 }),
  .ZN({ S11628 })
);
OAI21_X1 #() 
OAI21_X1_643_ (
  .A({ S11293 }),
  .B1({ S11624 }),
  .B2({ S11628 }),
  .ZN({ S11629 })
);
AOI21_X1 #() 
AOI21_X1_704_ (
  .A({ S11332 }),
  .B1({ S11391 }),
  .B2({ S11510 }),
  .ZN({ S11630 })
);
NAND2_X1 #() 
NAND2_X1_1123_ (
  .A1({ S24 }),
  .A2({ S33 }),
  .ZN({ S11632 })
);
AOI21_X1 #() 
AOI21_X1_705_ (
  .A({ S25957[388] }),
  .B1({ S11526 }),
  .B2({ S11632 }),
  .ZN({ S11633 })
);
OAI21_X1 #() 
OAI21_X1_644_ (
  .A({ S25957[389] }),
  .B1({ S11630 }),
  .B2({ S11633 }),
  .ZN({ S11634 })
);
AND2_X1 #() 
AND2_X1_68_ (
  .A1({ S11634 }),
  .A2({ S11629 }),
  .ZN({ S11635 })
);
NAND2_X1 #() 
NAND2_X1_1124_ (
  .A1({ S11363 }),
  .A2({ S11311 }),
  .ZN({ S11636 })
);
OAI211_X1 #() 
OAI211_X1_408_ (
  .A({ S11325 }),
  .B({ S25957[388] }),
  .C1({ S11308 }),
  .C2({ S11636 }),
  .ZN({ S11637 })
);
NAND2_X1 #() 
NAND2_X1_1125_ (
  .A1({ S11419 }),
  .A2({ S11368 }),
  .ZN({ S11638 })
);
INV_X1 #() 
INV_X1_367_ (
  .A({ S11638 }),
  .ZN({ S11639 })
);
AOI21_X1 #() 
AOI21_X1_706_ (
  .A({ S25957[388] }),
  .B1({ S25957[387] }),
  .B2({ S25957[386] }),
  .ZN({ S11640 })
);
OAI21_X1 #() 
OAI21_X1_645_ (
  .A({ S11640 }),
  .B1({ S11639 }),
  .B2({ S25957[387] }),
  .ZN({ S11641 })
);
NAND3_X1 #() 
NAND3_X1_1297_ (
  .A1({ S11637 }),
  .A2({ S11641 }),
  .A3({ S11293 }),
  .ZN({ S11643 })
);
AOI21_X1 #() 
AOI21_X1_707_ (
  .A({ S25957[387] }),
  .B1({ S11299 }),
  .B2({ S11509 }),
  .ZN({ S11644 })
);
OAI21_X1 #() 
OAI21_X1_646_ (
  .A({ S11332 }),
  .B1({ S11387 }),
  .B2({ S11545 }),
  .ZN({ S11645 })
);
INV_X1 #() 
INV_X1_368_ (
  .A({ S145 }),
  .ZN({ S11646 })
);
OAI21_X1 #() 
OAI21_X1_647_ (
  .A({ S25957[388] }),
  .B1({ S11646 }),
  .B2({ S25957[386] }),
  .ZN({ S11647 })
);
OAI211_X1 #() 
OAI211_X1_409_ (
  .A({ S25957[389] }),
  .B({ S11647 }),
  .C1({ S11645 }),
  .C2({ S11644 }),
  .ZN({ S11648 })
);
NAND2_X1 #() 
NAND2_X1_1126_ (
  .A1({ S11643 }),
  .A2({ S11648 }),
  .ZN({ S11649 })
);
NAND2_X1 #() 
NAND2_X1_1127_ (
  .A1({ S11649 }),
  .A2({ S25957[390] }),
  .ZN({ S11650 })
);
OAI211_X1 #() 
OAI211_X1_410_ (
  .A({ S11650 }),
  .B({ S11362 }),
  .C1({ S11635 }),
  .C2({ S25957[390] }),
  .ZN({ S11651 })
);
NAND3_X1 #() 
NAND3_X1_1298_ (
  .A1({ S11651 }),
  .A2({ S11621 }),
  .A3({ S25957[588] }),
  .ZN({ S11652 })
);
INV_X1 #() 
INV_X1_369_ (
  .A({ S11652 }),
  .ZN({ S11654 })
);
AOI21_X1 #() 
AOI21_X1_708_ (
  .A({ S25957[588] }),
  .B1({ S11651 }),
  .B2({ S11621 }),
  .ZN({ S11655 })
);
OAI21_X1 #() 
OAI21_X1_648_ (
  .A({ S10523 }),
  .B1({ S11654 }),
  .B2({ S11655 }),
  .ZN({ S11656 })
);
NAND2_X1 #() 
NAND2_X1_1128_ (
  .A1({ S11651 }),
  .A2({ S11621 }),
  .ZN({ S11657 })
);
NAND2_X1 #() 
NAND2_X1_1129_ (
  .A1({ S11657 }),
  .A2({ S11591 }),
  .ZN({ S11658 })
);
NAND3_X1 #() 
NAND3_X1_1299_ (
  .A1({ S11658 }),
  .A2({ S25957[428] }),
  .A3({ S11652 }),
  .ZN({ S11659 })
);
NAND3_X1 #() 
NAND3_X1_1300_ (
  .A1({ S11656 }),
  .A2({ S11659 }),
  .A3({ S25957[396] }),
  .ZN({ S11660 })
);
OAI21_X1 #() 
OAI21_X1_649_ (
  .A({ S25957[428] }),
  .B1({ S11654 }),
  .B2({ S11655 }),
  .ZN({ S11661 })
);
NAND3_X1 #() 
NAND3_X1_1301_ (
  .A1({ S11658 }),
  .A2({ S10523 }),
  .A3({ S11652 }),
  .ZN({ S11662 })
);
NAND3_X1 #() 
NAND3_X1_1302_ (
  .A1({ S11661 }),
  .A2({ S11662 }),
  .A3({ S10526 }),
  .ZN({ S11663 })
);
NAND2_X1 #() 
NAND2_X1_1130_ (
  .A1({ S11660 }),
  .A2({ S11663 }),
  .ZN({ S25957[268] })
);
NOR2_X1 #() 
NOR2_X1_266_ (
  .A1({ S8755 }),
  .A2({ S8758 }),
  .ZN({ S25957[427] })
);
NOR2_X1 #() 
NOR2_X1_267_ (
  .A1({ S5896 }),
  .A2({ S5897 }),
  .ZN({ S25957[587] })
);
INV_X1 #() 
INV_X1_370_ (
  .A({ S25957[587] }),
  .ZN({ S11665 })
);
NAND3_X1 #() 
NAND3_X1_1303_ (
  .A1({ S11344 }),
  .A2({ S24 }),
  .A3({ S11301 }),
  .ZN({ S11666 })
);
NAND3_X1 #() 
NAND3_X1_1304_ (
  .A1({ S25957[387] }),
  .A2({ S11423 }),
  .A3({ S11452 }),
  .ZN({ S11667 })
);
AND2_X1 #() 
AND2_X1_69_ (
  .A1({ S11667 }),
  .A2({ S11666 }),
  .ZN({ S11668 })
);
NAND2_X1 #() 
NAND2_X1_1131_ (
  .A1({ S11379 }),
  .A2({ S24 }),
  .ZN({ S11669 })
);
AOI21_X1 #() 
AOI21_X1_709_ (
  .A({ S11332 }),
  .B1({ S25957[387] }),
  .B2({ S11625 }),
  .ZN({ S11670 })
);
OAI21_X1 #() 
OAI21_X1_650_ (
  .A({ S11670 }),
  .B1({ S11339 }),
  .B2({ S11669 }),
  .ZN({ S11671 })
);
OAI211_X1 #() 
OAI211_X1_411_ (
  .A({ S25957[389] }),
  .B({ S11671 }),
  .C1({ S11668 }),
  .C2({ S25957[388] }),
  .ZN({ S11673 })
);
NAND3_X1 #() 
NAND3_X1_1305_ (
  .A1({ S11640 }),
  .A2({ S34 }),
  .A3({ S11309 }),
  .ZN({ S11674 })
);
OAI21_X1 #() 
OAI21_X1_651_ (
  .A({ S25957[387] }),
  .B1({ S11353 }),
  .B2({ S11324 }),
  .ZN({ S11675 })
);
NAND3_X1 #() 
NAND3_X1_1306_ (
  .A1({ S11313 }),
  .A2({ S24 }),
  .A3({ S11354 }),
  .ZN({ S11676 })
);
AND2_X1 #() 
AND2_X1_70_ (
  .A1({ S11676 }),
  .A2({ S11675 }),
  .ZN({ S11677 })
);
OAI211_X1 #() 
OAI211_X1_412_ (
  .A({ S11293 }),
  .B({ S11674 }),
  .C1({ S11677 }),
  .C2({ S11332 }),
  .ZN({ S11678 })
);
NAND3_X1 #() 
NAND3_X1_1307_ (
  .A1({ S11678 }),
  .A2({ S11673 }),
  .A3({ S25957[390] }),
  .ZN({ S11679 })
);
OAI21_X1 #() 
OAI21_X1_652_ (
  .A({ S11309 }),
  .B1({ S11339 }),
  .B2({ S11298 }),
  .ZN({ S11680 })
);
NAND2_X1 #() 
NAND2_X1_1132_ (
  .A1({ S11680 }),
  .A2({ S24 }),
  .ZN({ S11681 })
);
OAI211_X1 #() 
OAI211_X1_413_ (
  .A({ S11681 }),
  .B({ S25957[388] }),
  .C1({ S11525 }),
  .C2({ S11460 }),
  .ZN({ S11682 })
);
NAND2_X1 #() 
NAND2_X1_1133_ (
  .A1({ S11297 }),
  .A2({ S11312 }),
  .ZN({ S11684 })
);
NAND3_X1 #() 
NAND3_X1_1308_ (
  .A1({ S11684 }),
  .A2({ S25957[387] }),
  .A3({ S11301 }),
  .ZN({ S11685 })
);
NAND3_X1 #() 
NAND3_X1_1309_ (
  .A1({ S11377 }),
  .A2({ S24 }),
  .A3({ S11363 }),
  .ZN({ S11686 })
);
NAND3_X1 #() 
NAND3_X1_1310_ (
  .A1({ S11685 }),
  .A2({ S11686 }),
  .A3({ S11332 }),
  .ZN({ S11687 })
);
NAND3_X1 #() 
NAND3_X1_1311_ (
  .A1({ S11682 }),
  .A2({ S11687 }),
  .A3({ S25957[389] }),
  .ZN({ S11688 })
);
NAND3_X1 #() 
NAND3_X1_1312_ (
  .A1({ S24 }),
  .A2({ S11301 }),
  .A3({ S11363 }),
  .ZN({ S11689 })
);
NAND2_X1 #() 
NAND2_X1_1134_ (
  .A1({ S11398 }),
  .A2({ S25957[387] }),
  .ZN({ S11690 })
);
NAND3_X1 #() 
NAND3_X1_1313_ (
  .A1({ S11690 }),
  .A2({ S25957[388] }),
  .A3({ S11689 }),
  .ZN({ S11691 })
);
NAND2_X1 #() 
NAND2_X1_1135_ (
  .A1({ S11313 }),
  .A2({ S11363 }),
  .ZN({ S11692 })
);
AOI22_X1 #() 
AOI22_X1_151_ (
  .A1({ S11692 }),
  .A2({ S25957[387] }),
  .B1({ S11397 }),
  .B2({ S34 }),
  .ZN({ S11693 })
);
OAI211_X1 #() 
OAI211_X1_414_ (
  .A({ S11293 }),
  .B({ S11691 }),
  .C1({ S11693 }),
  .C2({ S25957[388] }),
  .ZN({ S11695 })
);
NAND3_X1 #() 
NAND3_X1_1314_ (
  .A1({ S11695 }),
  .A2({ S11688 }),
  .A3({ S11418 }),
  .ZN({ S11696 })
);
NAND3_X1 #() 
NAND3_X1_1315_ (
  .A1({ S11679 }),
  .A2({ S11696 }),
  .A3({ S25957[391] }),
  .ZN({ S11697 })
);
NAND2_X1 #() 
NAND2_X1_1136_ (
  .A1({ S11403 }),
  .A2({ S24 }),
  .ZN({ S11698 })
);
NAND2_X1 #() 
NAND2_X1_1137_ (
  .A1({ S11698 }),
  .A2({ S11332 }),
  .ZN({ S11699 })
);
NAND3_X1 #() 
NAND3_X1_1316_ (
  .A1({ S24 }),
  .A2({ S11368 }),
  .A3({ S11292 }),
  .ZN({ S11700 })
);
OR2_X1 #() 
OR2_X1_15_ (
  .A1({ S11700 }),
  .A2({ S11332 }),
  .ZN({ S11701 })
);
OAI211_X1 #() 
OAI211_X1_415_ (
  .A({ S11293 }),
  .B({ S11701 }),
  .C1({ S11699 }),
  .C2({ S11623 }),
  .ZN({ S11702 })
);
OAI211_X1 #() 
OAI211_X1_416_ (
  .A({ S11332 }),
  .B({ S11435 }),
  .C1({ S11556 }),
  .C2({ S11365 }),
  .ZN({ S11703 })
);
AOI22_X1 #() 
AOI22_X1_152_ (
  .A1({ S11378 }),
  .A2({ S11377 }),
  .B1({ S11680 }),
  .B2({ S25957[387] }),
  .ZN({ S11704 })
);
OAI211_X1 #() 
OAI211_X1_417_ (
  .A({ S25957[389] }),
  .B({ S11703 }),
  .C1({ S11704 }),
  .C2({ S11332 }),
  .ZN({ S11706 })
);
NAND3_X1 #() 
NAND3_X1_1317_ (
  .A1({ S11702 }),
  .A2({ S11706 }),
  .A3({ S25957[390] }),
  .ZN({ S11707 })
);
NAND3_X1 #() 
NAND3_X1_1318_ (
  .A1({ S11354 }),
  .A2({ S24 }),
  .A3({ S11297 }),
  .ZN({ S11708 })
);
OAI21_X1 #() 
OAI21_X1_653_ (
  .A({ S34 }),
  .B1({ S11292 }),
  .B2({ S25957[386] }),
  .ZN({ S11709 })
);
NAND2_X1 #() 
NAND2_X1_1138_ (
  .A1({ S11709 }),
  .A2({ S25957[387] }),
  .ZN({ S11710 })
);
NAND3_X1 #() 
NAND3_X1_1319_ (
  .A1({ S11710 }),
  .A2({ S11708 }),
  .A3({ S25957[388] }),
  .ZN({ S11711 })
);
AOI22_X1 #() 
AOI22_X1_153_ (
  .A1({ S11638 }),
  .A2({ S25957[387] }),
  .B1({ S11397 }),
  .B2({ S11377 }),
  .ZN({ S11712 })
);
OAI211_X1 #() 
OAI211_X1_418_ (
  .A({ S11293 }),
  .B({ S11711 }),
  .C1({ S11712 }),
  .C2({ S25957[388] }),
  .ZN({ S11713 })
);
OAI221_X1 #() 
OAI221_X1_27_ (
  .A({ S25957[388] }),
  .B1({ S11520 }),
  .B2({ S11388 }),
  .C1({ S11313 }),
  .C2({ S25957[387] }),
  .ZN({ S11714 })
);
NAND2_X1 #() 
NAND2_X1_1139_ (
  .A1({ S11389 }),
  .A2({ S25957[384] }),
  .ZN({ S11715 })
);
OAI21_X1 #() 
OAI21_X1_654_ (
  .A({ S11332 }),
  .B1({ S11333 }),
  .B2({ S11715 }),
  .ZN({ S11717 })
);
NAND3_X1 #() 
NAND3_X1_1320_ (
  .A1({ S11717 }),
  .A2({ S11714 }),
  .A3({ S25957[389] }),
  .ZN({ S11718 })
);
NAND3_X1 #() 
NAND3_X1_1321_ (
  .A1({ S11713 }),
  .A2({ S11418 }),
  .A3({ S11718 }),
  .ZN({ S11719 })
);
NAND3_X1 #() 
NAND3_X1_1322_ (
  .A1({ S11707 }),
  .A2({ S11719 }),
  .A3({ S11362 }),
  .ZN({ S11720 })
);
AND3_X1 #() 
AND3_X1_53_ (
  .A1({ S11697 }),
  .A2({ S11720 }),
  .A3({ S11665 }),
  .ZN({ S11721 })
);
AOI21_X1 #() 
AOI21_X1_710_ (
  .A({ S11665 }),
  .B1({ S11697 }),
  .B2({ S11720 }),
  .ZN({ S11722 })
);
OAI21_X1 #() 
OAI21_X1_655_ (
  .A({ S25957[427] }),
  .B1({ S11721 }),
  .B2({ S11722 }),
  .ZN({ S11723 })
);
INV_X1 #() 
INV_X1_371_ (
  .A({ S25957[427] }),
  .ZN({ S11724 })
);
NAND3_X1 #() 
NAND3_X1_1323_ (
  .A1({ S11697 }),
  .A2({ S11720 }),
  .A3({ S11665 }),
  .ZN({ S11725 })
);
NAND2_X1 #() 
NAND2_X1_1140_ (
  .A1({ S11697 }),
  .A2({ S11720 }),
  .ZN({ S11726 })
);
NAND2_X1 #() 
NAND2_X1_1141_ (
  .A1({ S11726 }),
  .A2({ S25957[587] }),
  .ZN({ S11728 })
);
NAND3_X1 #() 
NAND3_X1_1324_ (
  .A1({ S11728 }),
  .A2({ S11724 }),
  .A3({ S11725 }),
  .ZN({ S11729 })
);
NAND3_X1 #() 
NAND3_X1_1325_ (
  .A1({ S11723 }),
  .A2({ S11729 }),
  .A3({ S21 }),
  .ZN({ S11730 })
);
NAND3_X1 #() 
NAND3_X1_1326_ (
  .A1({ S11728 }),
  .A2({ S25957[427] }),
  .A3({ S11725 }),
  .ZN({ S11731 })
);
OAI21_X1 #() 
OAI21_X1_656_ (
  .A({ S11724 }),
  .B1({ S11721 }),
  .B2({ S11722 }),
  .ZN({ S11732 })
);
NAND3_X1 #() 
NAND3_X1_1327_ (
  .A1({ S11732 }),
  .A2({ S11731 }),
  .A3({ S25957[395] }),
  .ZN({ S11733 })
);
NAND2_X1 #() 
NAND2_X1_1142_ (
  .A1({ S11730 }),
  .A2({ S11733 }),
  .ZN({ S35 })
);
NAND3_X1 #() 
NAND3_X1_1328_ (
  .A1({ S11732 }),
  .A2({ S11731 }),
  .A3({ S21 }),
  .ZN({ S11734 })
);
NAND3_X1 #() 
NAND3_X1_1329_ (
  .A1({ S11723 }),
  .A2({ S11729 }),
  .A3({ S25957[395] }),
  .ZN({ S11735 })
);
NAND2_X1 #() 
NAND2_X1_1143_ (
  .A1({ S11734 }),
  .A2({ S11735 }),
  .ZN({ S25957[267] })
);
NOR2_X1 #() 
NOR2_X1_268_ (
  .A1({ S8833 }),
  .A2({ S8810 }),
  .ZN({ S25957[456] })
);
INV_X1 #() 
INV_X1_372_ (
  .A({ S25957[456] }),
  .ZN({ S11737 })
);
NAND4_X1 #() 
NAND4_X1_152_ (
  .A1({ S8786 }),
  .A2({ S8809 }),
  .A3({ S5957 }),
  .A4({ S6002 }),
  .ZN({ S11738 })
);
NAND2_X1 #() 
NAND2_X1_1144_ (
  .A1({ S5957 }),
  .A2({ S6002 }),
  .ZN({ S25957[616] })
);
NAND3_X1 #() 
NAND3_X1_1330_ (
  .A1({ S8818 }),
  .A2({ S8832 }),
  .A3({ S25957[616] }),
  .ZN({ S11739 })
);
NAND2_X1 #() 
NAND2_X1_1145_ (
  .A1({ S11738 }),
  .A2({ S11739 }),
  .ZN({ S25957[488] })
);
INV_X1 #() 
INV_X1_373_ (
  .A({ S25957[488] }),
  .ZN({ S11740 })
);
NAND3_X1 #() 
NAND3_X1_1331_ (
  .A1({ S11563 }),
  .A2({ S24 }),
  .A3({ S11354 }),
  .ZN({ S11741 })
);
NAND3_X1 #() 
NAND3_X1_1332_ (
  .A1({ S11355 }),
  .A2({ S11741 }),
  .A3({ S11332 }),
  .ZN({ S11742 })
);
AOI22_X1 #() 
AOI22_X1_154_ (
  .A1({ S25957[385] }),
  .A2({ S11300 }),
  .B1({ S9781 }),
  .B2({ S9786 }),
  .ZN({ S11743 })
);
NAND2_X1 #() 
NAND2_X1_1146_ (
  .A1({ S11743 }),
  .A2({ S25957[387] }),
  .ZN({ S11745 })
);
AND2_X1 #() 
AND2_X1_71_ (
  .A1({ S11627 }),
  .A2({ S11745 }),
  .ZN({ S11746 })
);
OAI211_X1 #() 
OAI211_X1_419_ (
  .A({ S25957[389] }),
  .B({ S11742 }),
  .C1({ S11746 }),
  .C2({ S11332 }),
  .ZN({ S11747 })
);
AOI21_X1 #() 
AOI21_X1_711_ (
  .A({ S25957[387] }),
  .B1({ S11423 }),
  .B2({ S11452 }),
  .ZN({ S11748 })
);
NOR2_X1 #() 
NOR2_X1_269_ (
  .A1({ S11313 }),
  .A2({ S24 }),
  .ZN({ S11749 })
);
OAI21_X1 #() 
OAI21_X1_657_ (
  .A({ S25957[388] }),
  .B1({ S11748 }),
  .B2({ S11749 }),
  .ZN({ S11750 })
);
AOI21_X1 #() 
AOI21_X1_712_ (
  .A({ S25957[387] }),
  .B1({ S11298 }),
  .B2({ S11436 }),
  .ZN({ S11751 })
);
OAI21_X1 #() 
OAI21_X1_658_ (
  .A({ S11332 }),
  .B1({ S11546 }),
  .B2({ S11751 }),
  .ZN({ S11752 })
);
NAND3_X1 #() 
NAND3_X1_1333_ (
  .A1({ S11752 }),
  .A2({ S11750 }),
  .A3({ S11293 }),
  .ZN({ S11753 })
);
NAND3_X1 #() 
NAND3_X1_1334_ (
  .A1({ S11753 }),
  .A2({ S11747 }),
  .A3({ S25957[390] }),
  .ZN({ S11754 })
);
OAI21_X1 #() 
OAI21_X1_659_ (
  .A({ S11332 }),
  .B1({ S11593 }),
  .B2({ S11614 }),
  .ZN({ S11756 })
);
NAND3_X1 #() 
NAND3_X1_1335_ (
  .A1({ S24 }),
  .A2({ S11300 }),
  .A3({ S11297 }),
  .ZN({ S11757 })
);
NAND2_X1 #() 
NAND2_X1_1147_ (
  .A1({ S11460 }),
  .A2({ S11700 }),
  .ZN({ S11758 })
);
NAND3_X1 #() 
NAND3_X1_1336_ (
  .A1({ S11758 }),
  .A2({ S25957[388] }),
  .A3({ S11757 }),
  .ZN({ S11759 })
);
NAND3_X1 #() 
NAND3_X1_1337_ (
  .A1({ S11759 }),
  .A2({ S11756 }),
  .A3({ S25957[389] }),
  .ZN({ S11760 })
);
AOI22_X1 #() 
AOI22_X1_155_ (
  .A1({ S11556 }),
  .A2({ S11297 }),
  .B1({ S11445 }),
  .B2({ S24 }),
  .ZN({ S11761 })
);
OAI211_X1 #() 
OAI211_X1_420_ (
  .A({ S25957[388] }),
  .B({ S11435 }),
  .C1({ S11299 }),
  .C2({ S25957[387] }),
  .ZN({ S11762 })
);
OAI211_X1 #() 
OAI211_X1_421_ (
  .A({ S11293 }),
  .B({ S11762 }),
  .C1({ S11761 }),
  .C2({ S25957[388] }),
  .ZN({ S11763 })
);
NAND3_X1 #() 
NAND3_X1_1338_ (
  .A1({ S11760 }),
  .A2({ S11418 }),
  .A3({ S11763 }),
  .ZN({ S11764 })
);
NAND3_X1 #() 
NAND3_X1_1339_ (
  .A1({ S11754 }),
  .A2({ S11764 }),
  .A3({ S25957[391] }),
  .ZN({ S11765 })
);
NAND3_X1 #() 
NAND3_X1_1340_ (
  .A1({ S11566 }),
  .A2({ S11428 }),
  .A3({ S11332 }),
  .ZN({ S11767 })
);
AOI21_X1 #() 
AOI21_X1_713_ (
  .A({ S11293 }),
  .B1({ S11670 }),
  .B2({ S11557 }),
  .ZN({ S11768 })
);
NAND3_X1 #() 
NAND3_X1_1341_ (
  .A1({ S11377 }),
  .A2({ S25957[387] }),
  .A3({ S11427 }),
  .ZN({ S11769 })
);
AOI22_X1 #() 
AOI22_X1_156_ (
  .A1({ S9781 }),
  .A2({ S9786 }),
  .B1({ S11287 }),
  .B2({ S11286 }),
  .ZN({ S11770 })
);
OAI211_X1 #() 
OAI211_X1_422_ (
  .A({ S11324 }),
  .B({ S24 }),
  .C1({ S11310 }),
  .C2({ S11770 }),
  .ZN({ S11771 })
);
NAND3_X1 #() 
NAND3_X1_1342_ (
  .A1({ S11769 }),
  .A2({ S11771 }),
  .A3({ S11332 }),
  .ZN({ S11772 })
);
AOI21_X1 #() 
AOI21_X1_714_ (
  .A({ S11298 }),
  .B1({ S34 }),
  .B2({ S11292 }),
  .ZN({ S11773 })
);
OAI21_X1 #() 
OAI21_X1_660_ (
  .A({ S24 }),
  .B1({ S11773 }),
  .B2({ S11306 }),
  .ZN({ S11774 })
);
AOI21_X1 #() 
AOI21_X1_715_ (
  .A({ S11332 }),
  .B1({ S11398 }),
  .B2({ S25957[387] }),
  .ZN({ S11775 })
);
AOI21_X1 #() 
AOI21_X1_716_ (
  .A({ S25957[389] }),
  .B1({ S11774 }),
  .B2({ S11775 }),
  .ZN({ S11776 })
);
AOI22_X1 #() 
AOI22_X1_157_ (
  .A1({ S11776 }),
  .A2({ S11772 }),
  .B1({ S11768 }),
  .B2({ S11767 }),
  .ZN({ S11778 })
);
NAND4_X1 #() 
NAND4_X1_153_ (
  .A1({ S11363 }),
  .A2({ S34 }),
  .A3({ S9524 }),
  .A4({ S9515 }),
  .ZN({ S11779 })
);
NAND3_X1 #() 
NAND3_X1_1343_ (
  .A1({ S24 }),
  .A2({ S11301 }),
  .A3({ S11312 }),
  .ZN({ S11780 })
);
OAI211_X1 #() 
OAI211_X1_423_ (
  .A({ S25957[388] }),
  .B({ S11780 }),
  .C1({ S11549 }),
  .C2({ S11779 }),
  .ZN({ S11781 })
);
NAND2_X1 #() 
NAND2_X1_1148_ (
  .A1({ S25957[387] }),
  .A2({ S11306 }),
  .ZN({ S11782 })
);
NAND2_X1 #() 
NAND2_X1_1149_ (
  .A1({ S11445 }),
  .A2({ S25957[387] }),
  .ZN({ S11783 })
);
AOI21_X1 #() 
AOI21_X1_717_ (
  .A({ S25957[388] }),
  .B1({ S24 }),
  .B2({ S11350 }),
  .ZN({ S11784 })
);
NAND3_X1 #() 
NAND3_X1_1344_ (
  .A1({ S11784 }),
  .A2({ S11783 }),
  .A3({ S11782 }),
  .ZN({ S11785 })
);
NAND3_X1 #() 
NAND3_X1_1345_ (
  .A1({ S11785 }),
  .A2({ S11781 }),
  .A3({ S25957[389] }),
  .ZN({ S11786 })
);
NAND4_X1 #() 
NAND4_X1_154_ (
  .A1({ S11553 }),
  .A2({ S11520 }),
  .A3({ S25957[388] }),
  .A4({ S11388 }),
  .ZN({ S11787 })
);
OAI21_X1 #() 
OAI21_X1_661_ (
  .A({ S11787 }),
  .B1({ S11645 }),
  .B2({ S11516 }),
  .ZN({ S11789 })
);
NAND2_X1 #() 
NAND2_X1_1150_ (
  .A1({ S11789 }),
  .A2({ S11293 }),
  .ZN({ S11790 })
);
NAND3_X1 #() 
NAND3_X1_1346_ (
  .A1({ S11790 }),
  .A2({ S25957[390] }),
  .A3({ S11786 }),
  .ZN({ S11791 })
);
OAI211_X1 #() 
OAI211_X1_424_ (
  .A({ S11791 }),
  .B({ S11362 }),
  .C1({ S25957[390] }),
  .C2({ S11778 }),
  .ZN({ S11792 })
);
NAND3_X1 #() 
NAND3_X1_1347_ (
  .A1({ S11792 }),
  .A2({ S11765 }),
  .A3({ S11740 }),
  .ZN({ S11793 })
);
OAI211_X1 #() 
OAI211_X1_425_ (
  .A({ S11787 }),
  .B({ S11293 }),
  .C1({ S11645 }),
  .C2({ S11516 }),
  .ZN({ S11794 })
);
NAND3_X1 #() 
NAND3_X1_1348_ (
  .A1({ S11377 }),
  .A2({ S25957[387] }),
  .A3({ S11345 }),
  .ZN({ S11795 })
);
AOI21_X1 #() 
AOI21_X1_718_ (
  .A({ S11332 }),
  .B1({ S11795 }),
  .B2({ S11477 }),
  .ZN({ S11796 })
);
NAND2_X1 #() 
NAND2_X1_1151_ (
  .A1({ S11534 }),
  .A2({ S11332 }),
  .ZN({ S11797 })
);
NOR2_X1 #() 
NOR2_X1_270_ (
  .A1({ S11453 }),
  .A2({ S11797 }),
  .ZN({ S11798 })
);
OAI21_X1 #() 
OAI21_X1_662_ (
  .A({ S25957[389] }),
  .B1({ S11796 }),
  .B2({ S11798 }),
  .ZN({ S11800 })
);
AOI21_X1 #() 
AOI21_X1_719_ (
  .A({ S25957[391] }),
  .B1({ S11800 }),
  .B2({ S11794 }),
  .ZN({ S11801 })
);
AND3_X1 #() 
AND3_X1_54_ (
  .A1({ S11355 }),
  .A2({ S11741 }),
  .A3({ S11332 }),
  .ZN({ S11802 })
);
AOI21_X1 #() 
AOI21_X1_720_ (
  .A({ S11332 }),
  .B1({ S11627 }),
  .B2({ S11745 }),
  .ZN({ S11803 })
);
OAI21_X1 #() 
OAI21_X1_663_ (
  .A({ S25957[389] }),
  .B1({ S11802 }),
  .B2({ S11803 }),
  .ZN({ S11804 })
);
AOI22_X1 #() 
AOI22_X1_158_ (
  .A1({ S11368 }),
  .A2({ S11389 }),
  .B1({ S25957[385] }),
  .B2({ S25957[384] }),
  .ZN({ S11805 })
);
NAND2_X1 #() 
NAND2_X1_1152_ (
  .A1({ S11773 }),
  .A2({ S25957[387] }),
  .ZN({ S11806 })
);
OAI211_X1 #() 
OAI211_X1_426_ (
  .A({ S11806 }),
  .B({ S25957[388] }),
  .C1({ S25957[387] }),
  .C2({ S11805 }),
  .ZN({ S11807 })
);
NAND2_X1 #() 
NAND2_X1_1153_ (
  .A1({ S11549 }),
  .A2({ S11323 }),
  .ZN({ S11808 })
);
AOI21_X1 #() 
AOI21_X1_721_ (
  .A({ S25957[389] }),
  .B1({ S11808 }),
  .B2({ S11784 }),
  .ZN({ S11809 })
);
NAND2_X1 #() 
NAND2_X1_1154_ (
  .A1({ S11809 }),
  .A2({ S11807 }),
  .ZN({ S11811 })
);
AOI21_X1 #() 
AOI21_X1_722_ (
  .A({ S11362 }),
  .B1({ S11804 }),
  .B2({ S11811 }),
  .ZN({ S11812 })
);
OAI21_X1 #() 
OAI21_X1_664_ (
  .A({ S25957[390] }),
  .B1({ S11812 }),
  .B2({ S11801 }),
  .ZN({ S11813 })
);
NAND2_X1 #() 
NAND2_X1_1155_ (
  .A1({ S11768 }),
  .A2({ S11767 }),
  .ZN({ S11814 })
);
NAND2_X1 #() 
NAND2_X1_1156_ (
  .A1({ S11774 }),
  .A2({ S11775 }),
  .ZN({ S11815 })
);
NAND3_X1 #() 
NAND3_X1_1349_ (
  .A1({ S11815 }),
  .A2({ S11772 }),
  .A3({ S11293 }),
  .ZN({ S11816 })
);
AOI21_X1 #() 
AOI21_X1_723_ (
  .A({ S25957[391] }),
  .B1({ S11816 }),
  .B2({ S11814 }),
  .ZN({ S11817 })
);
NAND2_X1 #() 
NAND2_X1_1157_ (
  .A1({ S25957[387] }),
  .A2({ S11297 }),
  .ZN({ S11818 })
);
OAI211_X1 #() 
OAI211_X1_427_ (
  .A({ S11818 }),
  .B({ S11293 }),
  .C1({ S25957[387] }),
  .C2({ S11525 }),
  .ZN({ S11819 })
);
AOI22_X1 #() 
AOI22_X1_159_ (
  .A1({ S11770 }),
  .A2({ S25957[385] }),
  .B1({ S11339 }),
  .B2({ S11298 }),
  .ZN({ S11820 })
);
OAI211_X1 #() 
OAI211_X1_428_ (
  .A({ S25957[389] }),
  .B({ S11460 }),
  .C1({ S11820 }),
  .C2({ S25957[387] }),
  .ZN({ S11822 })
);
AOI21_X1 #() 
AOI21_X1_724_ (
  .A({ S11332 }),
  .B1({ S11822 }),
  .B2({ S11819 }),
  .ZN({ S11823 })
);
NAND4_X1 #() 
NAND4_X1_155_ (
  .A1({ S11592 }),
  .A2({ S25957[389] }),
  .A3({ S11543 }),
  .A4({ S11613 }),
  .ZN({ S11824 })
);
NAND3_X1 #() 
NAND3_X1_1350_ (
  .A1({ S11368 }),
  .A2({ S34 }),
  .A3({ S11350 }),
  .ZN({ S11825 })
);
NAND4_X1 #() 
NAND4_X1_156_ (
  .A1({ S11297 }),
  .A2({ S11300 }),
  .A3({ S9524 }),
  .A4({ S9515 }),
  .ZN({ S11826 })
);
OAI211_X1 #() 
OAI211_X1_429_ (
  .A({ S11293 }),
  .B({ S11826 }),
  .C1({ S11825 }),
  .C2({ S25957[387] }),
  .ZN({ S11827 })
);
AOI21_X1 #() 
AOI21_X1_725_ (
  .A({ S25957[388] }),
  .B1({ S11827 }),
  .B2({ S11824 }),
  .ZN({ S11828 })
);
NOR3_X1 #() 
NOR3_X1_37_ (
  .A1({ S11823 }),
  .A2({ S11828 }),
  .A3({ S11362 }),
  .ZN({ S11829 })
);
OAI21_X1 #() 
OAI21_X1_665_ (
  .A({ S11418 }),
  .B1({ S11829 }),
  .B2({ S11817 }),
  .ZN({ S11830 })
);
NAND3_X1 #() 
NAND3_X1_1351_ (
  .A1({ S11813 }),
  .A2({ S11830 }),
  .A3({ S25957[488] }),
  .ZN({ S11831 })
);
NAND3_X1 #() 
NAND3_X1_1352_ (
  .A1({ S11831 }),
  .A2({ S11737 }),
  .A3({ S11793 }),
  .ZN({ S11833 })
);
NAND3_X1 #() 
NAND3_X1_1353_ (
  .A1({ S11792 }),
  .A2({ S11765 }),
  .A3({ S25957[488] }),
  .ZN({ S11834 })
);
NAND3_X1 #() 
NAND3_X1_1354_ (
  .A1({ S11813 }),
  .A2({ S11830 }),
  .A3({ S11740 }),
  .ZN({ S11835 })
);
NAND3_X1 #() 
NAND3_X1_1355_ (
  .A1({ S11835 }),
  .A2({ S25957[456] }),
  .A3({ S11834 }),
  .ZN({ S11836 })
);
AOI21_X1 #() 
AOI21_X1_726_ (
  .A({ S7576 }),
  .B1({ S11833 }),
  .B2({ S11836 }),
  .ZN({ S11837 })
);
NAND3_X1 #() 
NAND3_X1_1356_ (
  .A1({ S11831 }),
  .A2({ S25957[456] }),
  .A3({ S11793 }),
  .ZN({ S11838 })
);
NAND3_X1 #() 
NAND3_X1_1357_ (
  .A1({ S11835 }),
  .A2({ S11737 }),
  .A3({ S11834 }),
  .ZN({ S11839 })
);
AOI21_X1 #() 
AOI21_X1_727_ (
  .A({ S25957[520] }),
  .B1({ S11838 }),
  .B2({ S11839 }),
  .ZN({ S11840 })
);
NOR2_X1 #() 
NOR2_X1_271_ (
  .A1({ S11837 }),
  .A2({ S11840 }),
  .ZN({ S25957[264] })
);
NAND3_X1 #() 
NAND3_X1_1358_ (
  .A1({ S11377 }),
  .A2({ S25957[387] }),
  .A3({ S11309 }),
  .ZN({ S11841 })
);
AOI21_X1 #() 
AOI21_X1_728_ (
  .A({ S11332 }),
  .B1({ S11841 }),
  .B2({ S11385 }),
  .ZN({ S11843 })
);
NAND3_X1 #() 
NAND3_X1_1359_ (
  .A1({ S24 }),
  .A2({ S34 }),
  .A3({ S11297 }),
  .ZN({ S11844 })
);
AND3_X1 #() 
AND3_X1_55_ (
  .A1({ S11508 }),
  .A2({ S11332 }),
  .A3({ S11844 }),
  .ZN({ S11845 })
);
OAI21_X1 #() 
OAI21_X1_666_ (
  .A({ S25957[389] }),
  .B1({ S11845 }),
  .B2({ S11843 }),
  .ZN({ S11846 })
);
OAI211_X1 #() 
OAI211_X1_430_ (
  .A({ S11479 }),
  .B({ S25957[388] }),
  .C1({ S11440 }),
  .C2({ S25957[387] }),
  .ZN({ S11847 })
);
INV_X1 #() 
INV_X1_374_ (
  .A({ S11553 }),
  .ZN({ S11848 })
);
OAI21_X1 #() 
OAI21_X1_667_ (
  .A({ S11332 }),
  .B1({ S11848 }),
  .B2({ S11510 }),
  .ZN({ S11849 })
);
OAI211_X1 #() 
OAI211_X1_431_ (
  .A({ S11293 }),
  .B({ S11847 }),
  .C1({ S11849 }),
  .C2({ S11399 }),
  .ZN({ S11850 })
);
NAND3_X1 #() 
NAND3_X1_1360_ (
  .A1({ S11846 }),
  .A2({ S11418 }),
  .A3({ S11850 }),
  .ZN({ S11851 })
);
AOI21_X1 #() 
AOI21_X1_729_ (
  .A({ S24 }),
  .B1({ S11377 }),
  .B2({ S11345 }),
  .ZN({ S11852 })
);
NAND2_X1 #() 
NAND2_X1_1158_ (
  .A1({ S11669 }),
  .A2({ S11332 }),
  .ZN({ S11854 })
);
NAND2_X1 #() 
NAND2_X1_1159_ (
  .A1({ S11373 }),
  .A2({ S24 }),
  .ZN({ S11855 })
);
NAND3_X1 #() 
NAND3_X1_1361_ (
  .A1({ S11675 }),
  .A2({ S25957[388] }),
  .A3({ S11855 }),
  .ZN({ S11856 })
);
OAI211_X1 #() 
OAI211_X1_432_ (
  .A({ S11856 }),
  .B({ S25957[389] }),
  .C1({ S11852 }),
  .C2({ S11854 }),
  .ZN({ S11857 })
);
NAND3_X1 #() 
NAND3_X1_1362_ (
  .A1({ S11554 }),
  .A2({ S25957[388] }),
  .A3({ S11757 }),
  .ZN({ S11858 })
);
NAND2_X1 #() 
NAND2_X1_1160_ (
  .A1({ S11368 }),
  .A2({ S11292 }),
  .ZN({ S11859 })
);
OAI21_X1 #() 
OAI21_X1_668_ (
  .A({ S25957[387] }),
  .B1({ S11353 }),
  .B2({ S11339 }),
  .ZN({ S11860 })
);
OAI211_X1 #() 
OAI211_X1_433_ (
  .A({ S11860 }),
  .B({ S11332 }),
  .C1({ S11320 }),
  .C2({ S11859 }),
  .ZN({ S11861 })
);
NAND3_X1 #() 
NAND3_X1_1363_ (
  .A1({ S11858 }),
  .A2({ S11861 }),
  .A3({ S11293 }),
  .ZN({ S11862 })
);
NAND3_X1 #() 
NAND3_X1_1364_ (
  .A1({ S11862 }),
  .A2({ S11857 }),
  .A3({ S25957[390] }),
  .ZN({ S11863 })
);
NAND3_X1 #() 
NAND3_X1_1365_ (
  .A1({ S11851 }),
  .A2({ S11863 }),
  .A3({ S25957[391] }),
  .ZN({ S11865 })
);
NAND3_X1 #() 
NAND3_X1_1366_ (
  .A1({ S11325 }),
  .A2({ S11689 }),
  .A3({ S25957[388] }),
  .ZN({ S11866 })
);
OAI211_X1 #() 
OAI211_X1_434_ (
  .A({ S11782 }),
  .B({ S11332 }),
  .C1({ S11390 }),
  .C2({ S11302 }),
  .ZN({ S11867 })
);
NAND3_X1 #() 
NAND3_X1_1367_ (
  .A1({ S11866 }),
  .A2({ S11867 }),
  .A3({ S11293 }),
  .ZN({ S11868 })
);
AOI21_X1 #() 
AOI21_X1_730_ (
  .A({ S11332 }),
  .B1({ S11685 }),
  .B2({ S11594 }),
  .ZN({ S11869 })
);
OAI21_X1 #() 
OAI21_X1_669_ (
  .A({ S25957[389] }),
  .B1({ S11869 }),
  .B2({ S11405 }),
  .ZN({ S11870 })
);
NAND3_X1 #() 
NAND3_X1_1368_ (
  .A1({ S11870 }),
  .A2({ S11418 }),
  .A3({ S11868 }),
  .ZN({ S11871 })
);
NAND2_X1 #() 
NAND2_X1_1161_ (
  .A1({ S11710 }),
  .A2({ S25957[388] }),
  .ZN({ S11872 })
);
NOR2_X1 #() 
NOR2_X1_272_ (
  .A1({ S11592 }),
  .A2({ S11310 }),
  .ZN({ S11873 })
);
NAND4_X1 #() 
NAND4_X1_157_ (
  .A1({ S11536 }),
  .A2({ S11319 }),
  .A3({ S11332 }),
  .A4({ S11368 }),
  .ZN({ S11874 })
);
OAI211_X1 #() 
OAI211_X1_435_ (
  .A({ S11874 }),
  .B({ S25957[389] }),
  .C1({ S11872 }),
  .C2({ S11873 }),
  .ZN({ S11876 })
);
NAND3_X1 #() 
NAND3_X1_1369_ (
  .A1({ S11319 }),
  .A2({ S11468 }),
  .A3({ S24 }),
  .ZN({ S11877 })
);
OAI211_X1 #() 
OAI211_X1_436_ (
  .A({ S11877 }),
  .B({ S25957[388] }),
  .C1({ S11549 }),
  .C2({ S11779 }),
  .ZN({ S11878 })
);
OAI211_X1 #() 
OAI211_X1_437_ (
  .A({ S11806 }),
  .B({ S11332 }),
  .C1({ S11310 }),
  .C2({ S11855 }),
  .ZN({ S11879 })
);
NAND3_X1 #() 
NAND3_X1_1370_ (
  .A1({ S11879 }),
  .A2({ S11878 }),
  .A3({ S11293 }),
  .ZN({ S11880 })
);
NAND3_X1 #() 
NAND3_X1_1371_ (
  .A1({ S11880 }),
  .A2({ S25957[390] }),
  .A3({ S11876 }),
  .ZN({ S11881 })
);
NAND3_X1 #() 
NAND3_X1_1372_ (
  .A1({ S11871 }),
  .A2({ S11881 }),
  .A3({ S11362 }),
  .ZN({ S11882 })
);
AND3_X1 #() 
AND3_X1_56_ (
  .A1({ S11865 }),
  .A2({ S11882 }),
  .A3({ S25957[585] }),
  .ZN({ S11883 })
);
AOI21_X1 #() 
AOI21_X1_731_ (
  .A({ S25957[585] }),
  .B1({ S11865 }),
  .B2({ S11882 }),
  .ZN({ S11884 })
);
OAI21_X1 #() 
OAI21_X1_670_ (
  .A({ S25957[521] }),
  .B1({ S11883 }),
  .B2({ S11884 }),
  .ZN({ S11885 })
);
NAND3_X1 #() 
NAND3_X1_1373_ (
  .A1({ S11865 }),
  .A2({ S11882 }),
  .A3({ S25957[585] }),
  .ZN({ S11887 })
);
NAND2_X1 #() 
NAND2_X1_1162_ (
  .A1({ S11865 }),
  .A2({ S11882 }),
  .ZN({ S11888 })
);
NAND2_X1 #() 
NAND2_X1_1163_ (
  .A1({ S11888 }),
  .A2({ S8934 }),
  .ZN({ S11889 })
);
NAND3_X1 #() 
NAND3_X1_1374_ (
  .A1({ S11889 }),
  .A2({ S11887 }),
  .A3({ S7588 }),
  .ZN({ S11890 })
);
NAND2_X1 #() 
NAND2_X1_1164_ (
  .A1({ S11885 }),
  .A2({ S11890 }),
  .ZN({ S25957[265] })
);
NAND2_X1 #() 
NAND2_X1_1165_ (
  .A1({ S6179 }),
  .A2({ S6178 }),
  .ZN({ S11891 })
);
NAND2_X1 #() 
NAND2_X1_1166_ (
  .A1({ S9035 }),
  .A2({ S9033 }),
  .ZN({ S25957[490] })
);
NOR2_X1 #() 
NOR2_X1_273_ (
  .A1({ S11684 }),
  .A2({ S24 }),
  .ZN({ S11892 })
);
OAI21_X1 #() 
OAI21_X1_671_ (
  .A({ S11332 }),
  .B1({ S11748 }),
  .B2({ S11892 }),
  .ZN({ S11893 })
);
NAND4_X1 #() 
NAND4_X1_158_ (
  .A1({ S11301 }),
  .A2({ S11363 }),
  .A3({ S9524 }),
  .A4({ S9515 }),
  .ZN({ S11894 })
);
NAND3_X1 #() 
NAND3_X1_1375_ (
  .A1({ S11423 }),
  .A2({ S11419 }),
  .A3({ S24 }),
  .ZN({ S11896 })
);
OAI211_X1 #() 
OAI211_X1_438_ (
  .A({ S11896 }),
  .B({ S25957[388] }),
  .C1({ S11894 }),
  .C2({ S11310 }),
  .ZN({ S11897 })
);
NAND3_X1 #() 
NAND3_X1_1376_ (
  .A1({ S11893 }),
  .A2({ S11293 }),
  .A3({ S11897 }),
  .ZN({ S11898 })
);
AOI21_X1 #() 
AOI21_X1_732_ (
  .A({ S24 }),
  .B1({ S11377 }),
  .B2({ S11398 }),
  .ZN({ S11899 })
);
OAI21_X1 #() 
OAI21_X1_672_ (
  .A({ S11332 }),
  .B1({ S25957[387] }),
  .B2({ S11715 }),
  .ZN({ S11900 })
);
NAND3_X1 #() 
NAND3_X1_1377_ (
  .A1({ S25957[387] }),
  .A2({ S11363 }),
  .A3({ S11311 }),
  .ZN({ S11901 })
);
AND2_X1 #() 
AND2_X1_72_ (
  .A1({ S11901 }),
  .A2({ S11700 }),
  .ZN({ S11902 })
);
OAI22_X1 #() 
OAI22_X1_32_ (
  .A1({ S11902 }),
  .A2({ S11332 }),
  .B1({ S11899 }),
  .B2({ S11900 }),
  .ZN({ S11903 })
);
OAI211_X1 #() 
OAI211_X1_439_ (
  .A({ S11898 }),
  .B({ S25957[390] }),
  .C1({ S11903 }),
  .C2({ S11293 }),
  .ZN({ S11904 })
);
NAND3_X1 #() 
NAND3_X1_1378_ (
  .A1({ S25957[387] }),
  .A2({ S11419 }),
  .A3({ S11468 }),
  .ZN({ S11905 })
);
NAND3_X1 #() 
NAND3_X1_1379_ (
  .A1({ S11905 }),
  .A2({ S11332 }),
  .A3({ S11437 }),
  .ZN({ S11907 })
);
NAND3_X1 #() 
NAND3_X1_1380_ (
  .A1({ S11319 }),
  .A2({ S25957[387] }),
  .A3({ S11368 }),
  .ZN({ S11908 })
);
NAND3_X1 #() 
NAND3_X1_1381_ (
  .A1({ S11686 }),
  .A2({ S11908 }),
  .A3({ S25957[388] }),
  .ZN({ S11909 })
);
NAND3_X1 #() 
NAND3_X1_1382_ (
  .A1({ S11909 }),
  .A2({ S11907 }),
  .A3({ S25957[389] }),
  .ZN({ S11910 })
);
NAND4_X1 #() 
NAND4_X1_159_ (
  .A1({ S11783 }),
  .A2({ S11741 }),
  .A3({ S11332 }),
  .A4({ S11782 }),
  .ZN({ S11911 })
);
OAI21_X1 #() 
OAI21_X1_673_ (
  .A({ S24 }),
  .B1({ S11364 }),
  .B2({ S11743 }),
  .ZN({ S11912 })
);
NAND4_X1 #() 
NAND4_X1_160_ (
  .A1({ S11309 }),
  .A2({ S9515 }),
  .A3({ S25957[385] }),
  .A4({ S9524 }),
  .ZN({ S11913 })
);
NAND3_X1 #() 
NAND3_X1_1383_ (
  .A1({ S11912 }),
  .A2({ S25957[388] }),
  .A3({ S11913 }),
  .ZN({ S11914 })
);
NAND3_X1 #() 
NAND3_X1_1384_ (
  .A1({ S11914 }),
  .A2({ S11911 }),
  .A3({ S11293 }),
  .ZN({ S11915 })
);
NAND2_X1 #() 
NAND2_X1_1167_ (
  .A1({ S11915 }),
  .A2({ S11910 }),
  .ZN({ S11916 })
);
NAND2_X1 #() 
NAND2_X1_1168_ (
  .A1({ S11916 }),
  .A2({ S11418 }),
  .ZN({ S11918 })
);
NAND3_X1 #() 
NAND3_X1_1385_ (
  .A1({ S11918 }),
  .A2({ S11904 }),
  .A3({ S11362 }),
  .ZN({ S11919 })
);
NAND2_X1 #() 
NAND2_X1_1169_ (
  .A1({ S11306 }),
  .A2({ S24 }),
  .ZN({ S11920 })
);
NAND3_X1 #() 
NAND3_X1_1386_ (
  .A1({ S11299 }),
  .A2({ S25957[387] }),
  .A3({ S11423 }),
  .ZN({ S11921 })
);
AOI22_X1 #() 
AOI22_X1_160_ (
  .A1({ S11366 }),
  .A2({ S11920 }),
  .B1({ S11528 }),
  .B2({ S11921 }),
  .ZN({ S11922 })
);
NAND3_X1 #() 
NAND3_X1_1387_ (
  .A1({ S11299 }),
  .A2({ S25957[387] }),
  .A3({ S11509 }),
  .ZN({ S11923 })
);
NAND3_X1 #() 
NAND3_X1_1388_ (
  .A1({ S11923 }),
  .A2({ S11332 }),
  .A3({ S11308 }),
  .ZN({ S11924 })
);
NAND2_X1 #() 
NAND2_X1_1170_ (
  .A1({ S11741 }),
  .A2({ S11894 }),
  .ZN({ S11925 })
);
AOI21_X1 #() 
AOI21_X1_733_ (
  .A({ S11293 }),
  .B1({ S11925 }),
  .B2({ S25957[388] }),
  .ZN({ S11926 })
);
AOI22_X1 #() 
AOI22_X1_161_ (
  .A1({ S11293 }),
  .A2({ S11922 }),
  .B1({ S11926 }),
  .B2({ S11924 }),
  .ZN({ S11927 })
);
NAND4_X1 #() 
NAND4_X1_161_ (
  .A1({ S11363 }),
  .A2({ S25957[384] }),
  .A3({ S9524 }),
  .A4({ S9515 }),
  .ZN({ S11929 })
);
OAI211_X1 #() 
OAI211_X1_440_ (
  .A({ S25957[388] }),
  .B({ S11929 }),
  .C1({ S11390 }),
  .C2({ S11302 }),
  .ZN({ S11930 })
);
OAI22_X1 #() 
OAI22_X1_33_ (
  .A1({ S11318 }),
  .A2({ S11298 }),
  .B1({ S9526 }),
  .B2({ S9525 }),
  .ZN({ S11931 })
);
OAI21_X1 #() 
OAI21_X1_674_ (
  .A({ S11312 }),
  .B1({ S11311 }),
  .B2({ S11298 }),
  .ZN({ S11932 })
);
OAI211_X1 #() 
OAI211_X1_441_ (
  .A({ S11931 }),
  .B({ S11332 }),
  .C1({ S11932 }),
  .C2({ S24 }),
  .ZN({ S11933 })
);
NAND3_X1 #() 
NAND3_X1_1389_ (
  .A1({ S11930 }),
  .A2({ S25957[389] }),
  .A3({ S11933 }),
  .ZN({ S11934 })
);
OAI211_X1 #() 
OAI211_X1_442_ (
  .A({ S11913 }),
  .B({ S25957[388] }),
  .C1({ S25957[387] }),
  .C2({ S11478 }),
  .ZN({ S11935 })
);
OAI211_X1 #() 
OAI211_X1_443_ (
  .A({ S11935 }),
  .B({ S11293 }),
  .C1({ S11438 }),
  .C2({ S25957[388] }),
  .ZN({ S11936 })
);
NAND2_X1 #() 
NAND2_X1_1171_ (
  .A1({ S11934 }),
  .A2({ S11936 }),
  .ZN({ S11937 })
);
NAND2_X1 #() 
NAND2_X1_1172_ (
  .A1({ S11937 }),
  .A2({ S11418 }),
  .ZN({ S11938 })
);
OAI211_X1 #() 
OAI211_X1_444_ (
  .A({ S11938 }),
  .B({ S25957[391] }),
  .C1({ S11927 }),
  .C2({ S11418 }),
  .ZN({ S11940 })
);
NAND3_X1 #() 
NAND3_X1_1390_ (
  .A1({ S11919 }),
  .A2({ S11940 }),
  .A3({ S25957[490] }),
  .ZN({ S11941 })
);
INV_X1 #() 
INV_X1_375_ (
  .A({ S25957[490] }),
  .ZN({ S11942 })
);
NAND3_X1 #() 
NAND3_X1_1391_ (
  .A1({ S11418 }),
  .A2({ S11934 }),
  .A3({ S11936 }),
  .ZN({ S11943 })
);
NAND2_X1 #() 
NAND2_X1_1173_ (
  .A1({ S11926 }),
  .A2({ S11924 }),
  .ZN({ S11944 })
);
NAND2_X1 #() 
NAND2_X1_1174_ (
  .A1({ S11366 }),
  .A2({ S11920 }),
  .ZN({ S11945 })
);
NAND2_X1 #() 
NAND2_X1_1175_ (
  .A1({ S11528 }),
  .A2({ S11921 }),
  .ZN({ S11946 })
);
NAND3_X1 #() 
NAND3_X1_1392_ (
  .A1({ S11945 }),
  .A2({ S11946 }),
  .A3({ S11293 }),
  .ZN({ S11947 })
);
NAND3_X1 #() 
NAND3_X1_1393_ (
  .A1({ S11944 }),
  .A2({ S11947 }),
  .A3({ S25957[390] }),
  .ZN({ S11948 })
);
NAND3_X1 #() 
NAND3_X1_1394_ (
  .A1({ S11948 }),
  .A2({ S25957[391] }),
  .A3({ S11943 }),
  .ZN({ S11949 })
);
NOR2_X1 #() 
NOR2_X1_274_ (
  .A1({ S11899 }),
  .A2({ S11900 }),
  .ZN({ S11951 })
);
AOI21_X1 #() 
AOI21_X1_734_ (
  .A({ S11332 }),
  .B1({ S11901 }),
  .B2({ S11700 }),
  .ZN({ S11952 })
);
OAI21_X1 #() 
OAI21_X1_675_ (
  .A({ S25957[389] }),
  .B1({ S11951 }),
  .B2({ S11952 }),
  .ZN({ S11953 })
);
NAND2_X1 #() 
NAND2_X1_1176_ (
  .A1({ S11547 }),
  .A2({ S25957[387] }),
  .ZN({ S11954 })
);
AOI22_X1 #() 
AOI22_X1_162_ (
  .A1({ S25957[384] }),
  .A2({ S11324 }),
  .B1({ S9786 }),
  .B2({ S9781 }),
  .ZN({ S11955 })
);
OAI21_X1 #() 
OAI21_X1_676_ (
  .A({ S24 }),
  .B1({ S11364 }),
  .B2({ S11955 }),
  .ZN({ S11956 })
);
NAND3_X1 #() 
NAND3_X1_1395_ (
  .A1({ S11956 }),
  .A2({ S11954 }),
  .A3({ S25957[388] }),
  .ZN({ S11957 })
);
NAND2_X1 #() 
NAND2_X1_1177_ (
  .A1({ S25957[387] }),
  .A2({ S11563 }),
  .ZN({ S11958 })
);
OAI211_X1 #() 
OAI211_X1_445_ (
  .A({ S11332 }),
  .B({ S11958 }),
  .C1({ S11805 }),
  .C2({ S25957[387] }),
  .ZN({ S11959 })
);
NAND3_X1 #() 
NAND3_X1_1396_ (
  .A1({ S11957 }),
  .A2({ S11293 }),
  .A3({ S11959 }),
  .ZN({ S11960 })
);
AOI21_X1 #() 
AOI21_X1_735_ (
  .A({ S11418 }),
  .B1({ S11953 }),
  .B2({ S11960 }),
  .ZN({ S11962 })
);
AOI21_X1 #() 
AOI21_X1_736_ (
  .A({ S25957[390] }),
  .B1({ S11915 }),
  .B2({ S11910 }),
  .ZN({ S11963 })
);
OAI21_X1 #() 
OAI21_X1_677_ (
  .A({ S11362 }),
  .B1({ S11962 }),
  .B2({ S11963 }),
  .ZN({ S11964 })
);
NAND3_X1 #() 
NAND3_X1_1397_ (
  .A1({ S11964 }),
  .A2({ S11942 }),
  .A3({ S11949 }),
  .ZN({ S11965 })
);
AOI21_X1 #() 
AOI21_X1_737_ (
  .A({ S11891 }),
  .B1({ S11941 }),
  .B2({ S11965 }),
  .ZN({ S11966 })
);
INV_X1 #() 
INV_X1_376_ (
  .A({ S11891 }),
  .ZN({ S25957[554] })
);
NAND3_X1 #() 
NAND3_X1_1398_ (
  .A1({ S11964 }),
  .A2({ S25957[490] }),
  .A3({ S11949 }),
  .ZN({ S11967 })
);
NAND3_X1 #() 
NAND3_X1_1399_ (
  .A1({ S11919 }),
  .A2({ S11940 }),
  .A3({ S11942 }),
  .ZN({ S11968 })
);
AOI21_X1 #() 
AOI21_X1_738_ (
  .A({ S25957[554] }),
  .B1({ S11968 }),
  .B2({ S11967 }),
  .ZN({ S11969 })
);
OAI21_X1 #() 
OAI21_X1_678_ (
  .A({ S25957[394] }),
  .B1({ S11966 }),
  .B2({ S11969 }),
  .ZN({ S11970 })
);
NAND3_X1 #() 
NAND3_X1_1400_ (
  .A1({ S11968 }),
  .A2({ S11967 }),
  .A3({ S25957[554] }),
  .ZN({ S11972 })
);
NAND3_X1 #() 
NAND3_X1_1401_ (
  .A1({ S11941 }),
  .A2({ S11965 }),
  .A3({ S11891 }),
  .ZN({ S11973 })
);
NAND3_X1 #() 
NAND3_X1_1402_ (
  .A1({ S11972 }),
  .A2({ S11973 }),
  .A3({ S10529 }),
  .ZN({ S11974 })
);
NAND2_X1 #() 
NAND2_X1_1178_ (
  .A1({ S11970 }),
  .A2({ S11974 }),
  .ZN({ S25957[266] })
);
AOI21_X1 #() 
AOI21_X1_739_ (
  .A({ S7386 }),
  .B1({ S10343 }),
  .B2({ S10344 }),
  .ZN({ S11975 })
);
AND3_X1 #() 
AND3_X1_57_ (
  .A1({ S10343 }),
  .A2({ S10344 }),
  .A3({ S7386 }),
  .ZN({ S11976 })
);
OAI21_X1 #() 
OAI21_X1_679_ (
  .A({ S25957[409] }),
  .B1({ S11975 }),
  .B2({ S11976 }),
  .ZN({ S11977 })
);
INV_X1 #() 
INV_X1_377_ (
  .A({ S11977 }),
  .ZN({ S36 })
);
NAND4_X1 #() 
NAND4_X1_162_ (
  .A1({ S10342 }),
  .A2({ S10345 }),
  .A3({ S10403 }),
  .A4({ S10406 }),
  .ZN({ S37 })
);
NOR2_X1 #() 
NOR2_X1_275_ (
  .A1({ S9178 }),
  .A2({ S9176 }),
  .ZN({ S25957[455] })
);
XOR2_X1 #() 
XOR2_X1_22_ (
  .A({ S6326 }),
  .B({ S25957[743] }),
  .Z({ S25957[615] })
);
NAND2_X1 #() 
NAND2_X1_1179_ (
  .A1({ S9127 }),
  .A2({ S9175 }),
  .ZN({ S11979 })
);
XOR2_X1 #() 
XOR2_X1_23_ (
  .A({ S11979 }),
  .B({ S25957[615] }),
  .Z({ S25957[487] })
);
INV_X1 #() 
INV_X1_378_ (
  .A({ S25957[487] }),
  .ZN({ S11980 })
);
NAND2_X1 #() 
NAND2_X1_1180_ (
  .A1({ S10005 }),
  .A2({ S10008 }),
  .ZN({ S11981 })
);
NAND3_X1 #() 
NAND3_X1_1403_ (
  .A1({ S10153 }),
  .A2({ S10155 }),
  .A3({ S9063 }),
  .ZN({ S11982 })
);
NAND3_X1 #() 
NAND3_X1_1404_ (
  .A1({ S10158 }),
  .A2({ S10157 }),
  .A3({ S25957[540] }),
  .ZN({ S11983 })
);
NAND2_X1 #() 
NAND2_X1_1181_ (
  .A1({ S11982 }),
  .A2({ S11983 }),
  .ZN({ S11984 })
);
NAND3_X1 #() 
NAND3_X1_1405_ (
  .A1({ S10405 }),
  .A2({ S10404 }),
  .A3({ S25957[537] }),
  .ZN({ S11985 })
);
NAND3_X1 #() 
NAND3_X1_1406_ (
  .A1({ S10397 }),
  .A2({ S10402 }),
  .A3({ S9169 }),
  .ZN({ S11986 })
);
NAND3_X1 #() 
NAND3_X1_1407_ (
  .A1({ S10498 }),
  .A2({ S9051 }),
  .A3({ S10502 }),
  .ZN({ S11988 })
);
NAND3_X1 #() 
NAND3_X1_1408_ (
  .A1({ S10505 }),
  .A2({ S25957[538] }),
  .A3({ S10506 }),
  .ZN({ S11989 })
);
NAND4_X1 #() 
NAND4_X1_163_ (
  .A1({ S11988 }),
  .A2({ S11989 }),
  .A3({ S11985 }),
  .A4({ S11986 }),
  .ZN({ S11990 })
);
AOI22_X1 #() 
AOI22_X1_163_ (
  .A1({ S11988 }),
  .A2({ S11989 }),
  .B1({ S11986 }),
  .B2({ S11985 }),
  .ZN({ S11991 })
);
NAND2_X1 #() 
NAND2_X1_1182_ (
  .A1({ S11991 }),
  .A2({ S25957[408] }),
  .ZN({ S11992 })
);
NAND2_X1 #() 
NAND2_X1_1183_ (
  .A1({ S11992 }),
  .A2({ S11990 }),
  .ZN({ S11993 })
);
NAND2_X1 #() 
NAND2_X1_1184_ (
  .A1({ S11993 }),
  .A2({ S25957[411] }),
  .ZN({ S11994 })
);
NAND4_X1 #() 
NAND4_X1_164_ (
  .A1({ S10342 }),
  .A2({ S10345 }),
  .A3({ S11988 }),
  .A4({ S11989 }),
  .ZN({ S11995 })
);
NAND4_X1 #() 
NAND4_X1_165_ (
  .A1({ S11988 }),
  .A2({ S11989 }),
  .A3({ S10403 }),
  .A4({ S10406 }),
  .ZN({ S11996 })
);
NAND3_X1 #() 
NAND3_X1_1409_ (
  .A1({ S11995 }),
  .A2({ S28 }),
  .A3({ S11996 }),
  .ZN({ S11997 })
);
AND3_X1 #() 
AND3_X1_58_ (
  .A1({ S11994 }),
  .A2({ S11984 }),
  .A3({ S11997 }),
  .ZN({ S11999 })
);
NAND2_X1 #() 
NAND2_X1_1185_ (
  .A1({ S11988 }),
  .A2({ S11989 }),
  .ZN({ S12000 })
);
NAND3_X1 #() 
NAND3_X1_1410_ (
  .A1({ S25957[408] }),
  .A2({ S25957[409] }),
  .A3({ S12000 }),
  .ZN({ S12001 })
);
OAI21_X1 #() 
OAI21_X1_680_ (
  .A({ S25957[411] }),
  .B1({ S11996 }),
  .B2({ S25957[408] }),
  .ZN({ S12002 })
);
INV_X1 #() 
INV_X1_379_ (
  .A({ S12002 }),
  .ZN({ S12003 })
);
NOR2_X1 #() 
NOR2_X1_276_ (
  .A1({ S11990 }),
  .A2({ S25957[408] }),
  .ZN({ S12004 })
);
NAND4_X1 #() 
NAND4_X1_166_ (
  .A1({ S10342 }),
  .A2({ S10345 }),
  .A3({ S10503 }),
  .A4({ S10507 }),
  .ZN({ S12005 })
);
NAND2_X1 #() 
NAND2_X1_1186_ (
  .A1({ S12005 }),
  .A2({ S28 }),
  .ZN({ S12006 })
);
NOR2_X1 #() 
NOR2_X1_277_ (
  .A1({ S12006 }),
  .A2({ S12004 }),
  .ZN({ S12007 })
);
AOI211_X1 #() 
AOI211_X1_16_ (
  .A({ S11984 }),
  .B({ S12007 }),
  .C1({ S12001 }),
  .C2({ S12003 }),
  .ZN({ S12008 })
);
OAI21_X1 #() 
OAI21_X1_681_ (
  .A({ S25957[413] }),
  .B1({ S12008 }),
  .B2({ S11999 }),
  .ZN({ S12010 })
);
NAND4_X1 #() 
NAND4_X1_167_ (
  .A1({ S10503 }),
  .A2({ S10507 }),
  .A3({ S11985 }),
  .A4({ S11986 }),
  .ZN({ S12011 })
);
NOR2_X1 #() 
NOR2_X1_278_ (
  .A1({ S11976 }),
  .A2({ S11975 }),
  .ZN({ S12012 })
);
OAI21_X1 #() 
OAI21_X1_682_ (
  .A({ S25957[411] }),
  .B1({ S12012 }),
  .B2({ S12000 }),
  .ZN({ S12013 })
);
INV_X1 #() 
INV_X1_380_ (
  .A({ S12013 }),
  .ZN({ S12014 })
);
NAND3_X1 #() 
NAND3_X1_1411_ (
  .A1({ S12011 }),
  .A2({ S11996 }),
  .A3({ S25957[408] }),
  .ZN({ S12015 })
);
AOI21_X1 #() 
AOI21_X1_740_ (
  .A({ S25957[412] }),
  .B1({ S12015 }),
  .B2({ S28 }),
  .ZN({ S12016 })
);
INV_X1 #() 
INV_X1_381_ (
  .A({ S12016 }),
  .ZN({ S12017 })
);
AOI21_X1 #() 
AOI21_X1_741_ (
  .A({ S12017 }),
  .B1({ S12014 }),
  .B2({ S12011 }),
  .ZN({ S12018 })
);
AND4_X1 #() 
AND4_X1_4_ (
  .A1({ S10342 }),
  .A2({ S10503 }),
  .A3({ S10507 }),
  .A4({ S10345 }),
  .ZN({ S12019 })
);
AOI21_X1 #() 
AOI21_X1_742_ (
  .A({ S12000 }),
  .B1({ S11977 }),
  .B2({ S37 }),
  .ZN({ S12021 })
);
OAI21_X1 #() 
OAI21_X1_683_ (
  .A({ S28 }),
  .B1({ S12021 }),
  .B2({ S12019 }),
  .ZN({ S12022 })
);
INV_X1 #() 
INV_X1_382_ (
  .A({ S12022 }),
  .ZN({ S12023 })
);
NAND2_X1 #() 
NAND2_X1_1187_ (
  .A1({ S11977 }),
  .A2({ S25957[410] }),
  .ZN({ S12024 })
);
NAND2_X1 #() 
NAND2_X1_1188_ (
  .A1({ S11985 }),
  .A2({ S11986 }),
  .ZN({ S12025 })
);
OAI21_X1 #() 
OAI21_X1_684_ (
  .A({ S12025 }),
  .B1({ S11975 }),
  .B2({ S11976 }),
  .ZN({ S12026 })
);
NAND4_X1 #() 
NAND4_X1_168_ (
  .A1({ S10342 }),
  .A2({ S10345 }),
  .A3({ S11985 }),
  .A4({ S11986 }),
  .ZN({ S12027 })
);
NAND3_X1 #() 
NAND3_X1_1412_ (
  .A1({ S12026 }),
  .A2({ S12000 }),
  .A3({ S12027 }),
  .ZN({ S12028 })
);
AOI21_X1 #() 
AOI21_X1_743_ (
  .A({ S28 }),
  .B1({ S12028 }),
  .B2({ S12024 }),
  .ZN({ S12029 })
);
NOR3_X1 #() 
NOR3_X1_38_ (
  .A1({ S12023 }),
  .A2({ S12029 }),
  .A3({ S11984 }),
  .ZN({ S12030 })
);
OR3_X1 #() 
OR3_X1_5_ (
  .A1({ S12030 }),
  .A2({ S12018 }),
  .A3({ S25957[413] }),
  .ZN({ S12032 })
);
AOI21_X1 #() 
AOI21_X1_744_ (
  .A({ S11981 }),
  .B1({ S12032 }),
  .B2({ S12010 }),
  .ZN({ S12033 })
);
AND2_X1 #() 
AND2_X1_73_ (
  .A1({ S10091 }),
  .A2({ S10088 }),
  .ZN({ S12034 })
);
NAND4_X1 #() 
NAND4_X1_169_ (
  .A1({ S10503 }),
  .A2({ S10507 }),
  .A3({ S10403 }),
  .A4({ S10406 }),
  .ZN({ S12035 })
);
NAND2_X1 #() 
NAND2_X1_1189_ (
  .A1({ S12005 }),
  .A2({ S12035 }),
  .ZN({ S12036 })
);
NAND2_X1 #() 
NAND2_X1_1190_ (
  .A1({ S28 }),
  .A2({ S11990 }),
  .ZN({ S12037 })
);
NAND3_X1 #() 
NAND3_X1_1413_ (
  .A1({ S12026 }),
  .A2({ S25957[411] }),
  .A3({ S12011 }),
  .ZN({ S12038 })
);
OAI21_X1 #() 
OAI21_X1_685_ (
  .A({ S12038 }),
  .B1({ S12036 }),
  .B2({ S12037 }),
  .ZN({ S12039 })
);
NAND2_X1 #() 
NAND2_X1_1191_ (
  .A1({ S28 }),
  .A2({ S25957[408] }),
  .ZN({ S12040 })
);
NAND2_X1 #() 
NAND2_X1_1192_ (
  .A1({ S12014 }),
  .A2({ S12035 }),
  .ZN({ S12041 })
);
AND3_X1 #() 
AND3_X1_59_ (
  .A1({ S12041 }),
  .A2({ S12040 }),
  .A3({ S25957[412] }),
  .ZN({ S12043 })
);
AOI211_X1 #() 
AOI211_X1_17_ (
  .A({ S12034 }),
  .B({ S12043 }),
  .C1({ S11984 }),
  .C2({ S12039 }),
  .ZN({ S12044 })
);
NAND3_X1 #() 
NAND3_X1_1414_ (
  .A1({ S11977 }),
  .A2({ S25957[410] }),
  .A3({ S37 }),
  .ZN({ S12045 })
);
AOI22_X1 #() 
AOI22_X1_164_ (
  .A1({ S10342 }),
  .A2({ S10345 }),
  .B1({ S11989 }),
  .B2({ S11988 }),
  .ZN({ S12046 })
);
AOI21_X1 #() 
AOI21_X1_745_ (
  .A({ S25957[411] }),
  .B1({ S12046 }),
  .B2({ S25957[409] }),
  .ZN({ S12047 })
);
AOI21_X1 #() 
AOI21_X1_746_ (
  .A({ S11984 }),
  .B1({ S12047 }),
  .B2({ S12045 }),
  .ZN({ S12048 })
);
OAI21_X1 #() 
OAI21_X1_686_ (
  .A({ S12048 }),
  .B1({ S28 }),
  .B2({ S12004 }),
  .ZN({ S12049 })
);
NAND4_X1 #() 
NAND4_X1_170_ (
  .A1({ S12026 }),
  .A2({ S12027 }),
  .A3({ S28 }),
  .A4({ S25957[410] }),
  .ZN({ S12050 })
);
NAND2_X1 #() 
NAND2_X1_1193_ (
  .A1({ S25957[411] }),
  .A2({ S25957[410] }),
  .ZN({ S12051 })
);
OAI211_X1 #() 
OAI211_X1_446_ (
  .A({ S12050 }),
  .B({ S11984 }),
  .C1({ S36 }),
  .C2({ S12051 }),
  .ZN({ S12052 })
);
AND3_X1 #() 
AND3_X1_60_ (
  .A1({ S12049 }),
  .A2({ S12034 }),
  .A3({ S12052 }),
  .ZN({ S12054 })
);
NOR3_X1 #() 
NOR3_X1_39_ (
  .A1({ S12044 }),
  .A2({ S12054 }),
  .A3({ S25957[414] }),
  .ZN({ S12055 })
);
OAI21_X1 #() 
OAI21_X1_687_ (
  .A({ S9910 }),
  .B1({ S12055 }),
  .B2({ S12033 }),
  .ZN({ S12056 })
);
NAND2_X1 #() 
NAND2_X1_1194_ (
  .A1({ S12005 }),
  .A2({ S12011 }),
  .ZN({ S12057 })
);
AOI21_X1 #() 
AOI21_X1_747_ (
  .A({ S11984 }),
  .B1({ S12057 }),
  .B2({ S25957[411] }),
  .ZN({ S12058 })
);
OAI211_X1 #() 
OAI211_X1_447_ (
  .A({ S25957[410] }),
  .B({ S25957[409] }),
  .C1({ S10251 }),
  .C2({ S10250 }),
  .ZN({ S12059 })
);
AOI22_X1 #() 
AOI22_X1_165_ (
  .A1({ S10342 }),
  .A2({ S10345 }),
  .B1({ S10507 }),
  .B2({ S10503 }),
  .ZN({ S12060 })
);
NAND2_X1 #() 
NAND2_X1_1195_ (
  .A1({ S12060 }),
  .A2({ S25957[411] }),
  .ZN({ S12061 })
);
NAND3_X1 #() 
NAND3_X1_1415_ (
  .A1({ S28 }),
  .A2({ S25957[408] }),
  .A3({ S25957[409] }),
  .ZN({ S12062 })
);
NAND4_X1 #() 
NAND4_X1_171_ (
  .A1({ S12058 }),
  .A2({ S12059 }),
  .A3({ S12061 }),
  .A4({ S12062 }),
  .ZN({ S12063 })
);
NAND2_X1 #() 
NAND2_X1_1196_ (
  .A1({ S12026 }),
  .A2({ S12027 }),
  .ZN({ S12065 })
);
NAND3_X1 #() 
NAND3_X1_1416_ (
  .A1({ S12065 }),
  .A2({ S25957[411] }),
  .A3({ S12005 }),
  .ZN({ S12066 })
);
OAI211_X1 #() 
OAI211_X1_448_ (
  .A({ S28 }),
  .B({ S11990 }),
  .C1({ S12012 }),
  .C2({ S12000 }),
  .ZN({ S12067 })
);
OAI211_X1 #() 
OAI211_X1_449_ (
  .A({ S12066 }),
  .B({ S11984 }),
  .C1({ S12036 }),
  .C2({ S12067 }),
  .ZN({ S12068 })
);
NAND3_X1 #() 
NAND3_X1_1417_ (
  .A1({ S12068 }),
  .A2({ S12063 }),
  .A3({ S25957[413] }),
  .ZN({ S12069 })
);
INV_X1 #() 
INV_X1_383_ (
  .A({ S12027 }),
  .ZN({ S12070 })
);
NOR2_X1 #() 
NOR2_X1_279_ (
  .A1({ S12070 }),
  .A2({ S25957[411] }),
  .ZN({ S12071 })
);
NAND2_X1 #() 
NAND2_X1_1197_ (
  .A1({ S25957[411] }),
  .A2({ S11996 }),
  .ZN({ S12072 })
);
NOR2_X1 #() 
NOR2_X1_280_ (
  .A1({ S36 }),
  .A2({ S12072 }),
  .ZN({ S12073 })
);
OAI21_X1 #() 
OAI21_X1_688_ (
  .A({ S25957[412] }),
  .B1({ S12073 }),
  .B2({ S12071 }),
  .ZN({ S12074 })
);
NAND2_X1 #() 
NAND2_X1_1198_ (
  .A1({ S37 }),
  .A2({ S25957[410] }),
  .ZN({ S12076 })
);
NAND2_X1 #() 
NAND2_X1_1199_ (
  .A1({ S11991 }),
  .A2({ S12012 }),
  .ZN({ S12077 })
);
NOR2_X1 #() 
NOR2_X1_281_ (
  .A1({ S12026 }),
  .A2({ S28 }),
  .ZN({ S12078 })
);
NOR2_X1 #() 
NOR2_X1_282_ (
  .A1({ S12078 }),
  .A2({ S25957[412] }),
  .ZN({ S12079 })
);
NAND3_X1 #() 
NAND3_X1_1418_ (
  .A1({ S12079 }),
  .A2({ S12076 }),
  .A3({ S12077 }),
  .ZN({ S12080 })
);
AND2_X1 #() 
AND2_X1_74_ (
  .A1({ S12080 }),
  .A2({ S12074 }),
  .ZN({ S12081 })
);
OAI21_X1 #() 
OAI21_X1_689_ (
  .A({ S12069 }),
  .B1({ S12081 }),
  .B2({ S25957[413] }),
  .ZN({ S12082 })
);
NAND2_X1 #() 
NAND2_X1_1200_ (
  .A1({ S11991 }),
  .A2({ S25957[411] }),
  .ZN({ S12083 })
);
NAND4_X1 #() 
NAND4_X1_172_ (
  .A1({ S12015 }),
  .A2({ S12027 }),
  .A3({ S28 }),
  .A4({ S11995 }),
  .ZN({ S12084 })
);
AOI21_X1 #() 
AOI21_X1_748_ (
  .A({ S25957[412] }),
  .B1({ S12084 }),
  .B2({ S12083 }),
  .ZN({ S12085 })
);
NAND3_X1 #() 
NAND3_X1_1419_ (
  .A1({ S12026 }),
  .A2({ S25957[410] }),
  .A3({ S12027 }),
  .ZN({ S12087 })
);
NAND3_X1 #() 
NAND3_X1_1420_ (
  .A1({ S11977 }),
  .A2({ S12000 }),
  .A3({ S37 }),
  .ZN({ S12088 })
);
NAND3_X1 #() 
NAND3_X1_1421_ (
  .A1({ S12087 }),
  .A2({ S12088 }),
  .A3({ S25957[411] }),
  .ZN({ S12089 })
);
OAI211_X1 #() 
OAI211_X1_450_ (
  .A({ S10503 }),
  .B({ S10507 }),
  .C1({ S11976 }),
  .C2({ S11975 }),
  .ZN({ S12090 })
);
NAND2_X1 #() 
NAND2_X1_1201_ (
  .A1({ S12090 }),
  .A2({ S28 }),
  .ZN({ S12091 })
);
INV_X1 #() 
INV_X1_384_ (
  .A({ S12091 }),
  .ZN({ S12092 })
);
NAND2_X1 #() 
NAND2_X1_1202_ (
  .A1({ S12092 }),
  .A2({ S11990 }),
  .ZN({ S12093 })
);
NAND2_X1 #() 
NAND2_X1_1203_ (
  .A1({ S12093 }),
  .A2({ S12089 }),
  .ZN({ S12094 })
);
OAI21_X1 #() 
OAI21_X1_690_ (
  .A({ S12034 }),
  .B1({ S12094 }),
  .B2({ S11984 }),
  .ZN({ S12095 })
);
OAI21_X1 #() 
OAI21_X1_691_ (
  .A({ S25957[411] }),
  .B1({ S12060 }),
  .B2({ S12025 }),
  .ZN({ S12096 })
);
NAND2_X1 #() 
NAND2_X1_1204_ (
  .A1({ S25957[408] }),
  .A2({ S25957[410] }),
  .ZN({ S12098 })
);
AOI22_X1 #() 
AOI22_X1_166_ (
  .A1({ S10245 }),
  .A2({ S10249 }),
  .B1({ S10406 }),
  .B2({ S10403 }),
  .ZN({ S12099 })
);
NAND2_X1 #() 
NAND2_X1_1205_ (
  .A1({ S12098 }),
  .A2({ S12099 }),
  .ZN({ S12100 })
);
AOI21_X1 #() 
AOI21_X1_749_ (
  .A({ S11984 }),
  .B1({ S12096 }),
  .B2({ S12100 }),
  .ZN({ S12101 })
);
OAI21_X1 #() 
OAI21_X1_692_ (
  .A({ S28 }),
  .B1({ S12035 }),
  .B2({ S25957[408] }),
  .ZN({ S12102 })
);
AOI21_X1 #() 
AOI21_X1_750_ (
  .A({ S25957[412] }),
  .B1({ S12102 }),
  .B2({ S11977 }),
  .ZN({ S12103 })
);
OAI21_X1 #() 
OAI21_X1_693_ (
  .A({ S25957[413] }),
  .B1({ S12101 }),
  .B2({ S12103 }),
  .ZN({ S12104 })
);
OAI211_X1 #() 
OAI211_X1_451_ (
  .A({ S11981 }),
  .B({ S12104 }),
  .C1({ S12095 }),
  .C2({ S12085 }),
  .ZN({ S12105 })
);
OAI211_X1 #() 
OAI211_X1_452_ (
  .A({ S12105 }),
  .B({ S25957[415] }),
  .C1({ S12082 }),
  .C2({ S11981 }),
  .ZN({ S12106 })
);
NAND3_X1 #() 
NAND3_X1_1422_ (
  .A1({ S12056 }),
  .A2({ S11980 }),
  .A3({ S12106 }),
  .ZN({ S12107 })
);
NAND2_X1 #() 
NAND2_X1_1206_ (
  .A1({ S12056 }),
  .A2({ S12106 }),
  .ZN({ S12109 })
);
NAND2_X1 #() 
NAND2_X1_1207_ (
  .A1({ S12109 }),
  .A2({ S25957[487] }),
  .ZN({ S12110 })
);
NAND2_X1 #() 
NAND2_X1_1208_ (
  .A1({ S12110 }),
  .A2({ S12107 }),
  .ZN({ S25957[359] })
);
NAND2_X1 #() 
NAND2_X1_1209_ (
  .A1({ S25957[359] }),
  .A2({ S25957[455] }),
  .ZN({ S12111 })
);
INV_X1 #() 
INV_X1_385_ (
  .A({ S25957[455] }),
  .ZN({ S12112 })
);
NAND3_X1 #() 
NAND3_X1_1423_ (
  .A1({ S12110 }),
  .A2({ S12107 }),
  .A3({ S12112 }),
  .ZN({ S12113 })
);
NAND3_X1 #() 
NAND3_X1_1424_ (
  .A1({ S12111 }),
  .A2({ S12113 }),
  .A3({ S25957[423] }),
  .ZN({ S12114 })
);
INV_X1 #() 
INV_X1_386_ (
  .A({ S12114 }),
  .ZN({ S12115 })
);
AOI21_X1 #() 
AOI21_X1_751_ (
  .A({ S25957[423] }),
  .B1({ S12111 }),
  .B2({ S12113 }),
  .ZN({ S12116 })
);
OAI21_X1 #() 
OAI21_X1_694_ (
  .A({ S11362 }),
  .B1({ S12115 }),
  .B2({ S12116 }),
  .ZN({ S12117 })
);
INV_X1 #() 
INV_X1_387_ (
  .A({ S12116 }),
  .ZN({ S12119 })
);
NAND3_X1 #() 
NAND3_X1_1425_ (
  .A1({ S12119 }),
  .A2({ S25957[391] }),
  .A3({ S12114 }),
  .ZN({ S12120 })
);
NAND2_X1 #() 
NAND2_X1_1210_ (
  .A1({ S12117 }),
  .A2({ S12120 }),
  .ZN({ S12121 })
);
INV_X1 #() 
INV_X1_388_ (
  .A({ S12121 }),
  .ZN({ S25957[263] })
);
XOR2_X1 #() 
XOR2_X1_24_ (
  .A({ S25957[486] }),
  .B({ S25957[582] }),
  .Z({ S25957[454] })
);
AOI21_X1 #() 
AOI21_X1_752_ (
  .A({ S28 }),
  .B1({ S12076 }),
  .B2({ S12001 }),
  .ZN({ S12122 })
);
NAND2_X1 #() 
NAND2_X1_1211_ (
  .A1({ S12001 }),
  .A2({ S28 }),
  .ZN({ S12123 })
);
NAND2_X1 #() 
NAND2_X1_1212_ (
  .A1({ S12012 }),
  .A2({ S12011 }),
  .ZN({ S12124 })
);
INV_X1 #() 
INV_X1_389_ (
  .A({ S12124 }),
  .ZN({ S12125 })
);
NAND3_X1 #() 
NAND3_X1_1426_ (
  .A1({ S25957[408] }),
  .A2({ S12025 }),
  .A3({ S25957[410] }),
  .ZN({ S12126 })
);
NAND3_X1 #() 
NAND3_X1_1427_ (
  .A1({ S12126 }),
  .A2({ S25957[411] }),
  .A3({ S12005 }),
  .ZN({ S12128 })
);
OAI211_X1 #() 
OAI211_X1_453_ (
  .A({ S12128 }),
  .B({ S25957[412] }),
  .C1({ S12123 }),
  .C2({ S12125 }),
  .ZN({ S12129 })
);
OAI211_X1 #() 
OAI211_X1_454_ (
  .A({ S12129 }),
  .B({ S12034 }),
  .C1({ S12017 }),
  .C2({ S12122 }),
  .ZN({ S12130 })
);
INV_X1 #() 
INV_X1_390_ (
  .A({ S12130 }),
  .ZN({ S12131 })
);
OAI21_X1 #() 
OAI21_X1_695_ (
  .A({ S11984 }),
  .B1({ S12073 }),
  .B2({ S12099 }),
  .ZN({ S12132 })
);
NAND4_X1 #() 
NAND4_X1_173_ (
  .A1({ S12090 }),
  .A2({ S11995 }),
  .A3({ S25957[411] }),
  .A4({ S12025 }),
  .ZN({ S12133 })
);
OAI211_X1 #() 
OAI211_X1_455_ (
  .A({ S12133 }),
  .B({ S25957[412] }),
  .C1({ S25957[411] }),
  .C2({ S12076 }),
  .ZN({ S12134 })
);
AOI21_X1 #() 
AOI21_X1_753_ (
  .A({ S12034 }),
  .B1({ S12132 }),
  .B2({ S12134 }),
  .ZN({ S12135 })
);
OAI21_X1 #() 
OAI21_X1_696_ (
  .A({ S25957[414] }),
  .B1({ S12131 }),
  .B2({ S12135 }),
  .ZN({ S12136 })
);
INV_X1 #() 
INV_X1_391_ (
  .A({ S12065 }),
  .ZN({ S12137 })
);
INV_X1 #() 
INV_X1_392_ (
  .A({ S11996 }),
  .ZN({ S12139 })
);
NOR2_X1 #() 
NOR2_X1_283_ (
  .A1({ S12139 }),
  .A2({ S28 }),
  .ZN({ S12140 })
);
NAND4_X1 #() 
NAND4_X1_174_ (
  .A1({ S12000 }),
  .A2({ S25957[409] }),
  .A3({ S10345 }),
  .A4({ S10342 }),
  .ZN({ S12141 })
);
AOI22_X1 #() 
AOI22_X1_167_ (
  .A1({ S12092 }),
  .A2({ S12137 }),
  .B1({ S12140 }),
  .B2({ S12141 }),
  .ZN({ S12142 })
);
NOR2_X1 #() 
NOR2_X1_284_ (
  .A1({ S28 }),
  .A2({ S11990 }),
  .ZN({ S12143 })
);
NOR2_X1 #() 
NOR2_X1_285_ (
  .A1({ S12143 }),
  .A2({ S11984 }),
  .ZN({ S12144 })
);
OAI211_X1 #() 
OAI211_X1_456_ (
  .A({ S12144 }),
  .B({ S12050 }),
  .C1({ S12141 }),
  .C2({ S25957[411] }),
  .ZN({ S12145 })
);
OAI21_X1 #() 
OAI21_X1_697_ (
  .A({ S12145 }),
  .B1({ S12142 }),
  .B2({ S25957[412] }),
  .ZN({ S12146 })
);
INV_X1 #() 
INV_X1_393_ (
  .A({ S12096 }),
  .ZN({ S12147 })
);
AOI21_X1 #() 
AOI21_X1_754_ (
  .A({ S12147 }),
  .B1({ S12057 }),
  .B2({ S28 }),
  .ZN({ S12148 })
);
NAND2_X1 #() 
NAND2_X1_1213_ (
  .A1({ S12004 }),
  .A2({ S25957[411] }),
  .ZN({ S12150 })
);
AOI21_X1 #() 
AOI21_X1_755_ (
  .A({ S25957[412] }),
  .B1({ S12046 }),
  .B2({ S25957[411] }),
  .ZN({ S12151 })
);
OAI211_X1 #() 
OAI211_X1_457_ (
  .A({ S12150 }),
  .B({ S12151 }),
  .C1({ S12123 }),
  .C2({ S12125 }),
  .ZN({ S12152 })
);
OAI211_X1 #() 
OAI211_X1_458_ (
  .A({ S12034 }),
  .B({ S12152 }),
  .C1({ S12148 }),
  .C2({ S11984 }),
  .ZN({ S12153 })
);
OAI21_X1 #() 
OAI21_X1_698_ (
  .A({ S12153 }),
  .B1({ S12146 }),
  .B2({ S12034 }),
  .ZN({ S12154 })
);
NAND2_X1 #() 
NAND2_X1_1214_ (
  .A1({ S12154 }),
  .A2({ S11981 }),
  .ZN({ S12155 })
);
NAND2_X1 #() 
NAND2_X1_1215_ (
  .A1({ S12155 }),
  .A2({ S12136 }),
  .ZN({ S12156 })
);
NAND2_X1 #() 
NAND2_X1_1216_ (
  .A1({ S12156 }),
  .A2({ S25957[415] }),
  .ZN({ S12157 })
);
OAI211_X1 #() 
OAI211_X1_459_ (
  .A({ S25957[412] }),
  .B({ S12091 }),
  .C1({ S12002 }),
  .C2({ S36 }),
  .ZN({ S12158 })
);
INV_X1 #() 
INV_X1_394_ (
  .A({ S12011 }),
  .ZN({ S12159 })
);
NAND3_X1 #() 
NAND3_X1_1428_ (
  .A1({ S11992 }),
  .A2({ S28 }),
  .A3({ S11990 }),
  .ZN({ S12161 })
);
OAI211_X1 #() 
OAI211_X1_460_ (
  .A({ S12161 }),
  .B({ S11984 }),
  .C1({ S12159 }),
  .C2({ S12072 }),
  .ZN({ S12162 })
);
NAND3_X1 #() 
NAND3_X1_1429_ (
  .A1({ S12162 }),
  .A2({ S25957[413] }),
  .A3({ S12158 }),
  .ZN({ S12163 })
);
NAND2_X1 #() 
NAND2_X1_1217_ (
  .A1({ S12090 }),
  .A2({ S12035 }),
  .ZN({ S12164 })
);
OAI21_X1 #() 
OAI21_X1_699_ (
  .A({ S25957[411] }),
  .B1({ S12164 }),
  .B2({ S12004 }),
  .ZN({ S12165 })
);
OR2_X1 #() 
OR2_X1_16_ (
  .A1({ S12165 }),
  .A2({ S25957[412] }),
  .ZN({ S12166 })
);
AOI21_X1 #() 
AOI21_X1_756_ (
  .A({ S11984 }),
  .B1({ S11992 }),
  .B2({ S28 }),
  .ZN({ S12167 })
);
NAND2_X1 #() 
NAND2_X1_1218_ (
  .A1({ S11994 }),
  .A2({ S12167 }),
  .ZN({ S12168 })
);
AOI21_X1 #() 
AOI21_X1_757_ (
  .A({ S25957[413] }),
  .B1({ S12166 }),
  .B2({ S12168 }),
  .ZN({ S12169 })
);
NOR2_X1 #() 
NOR2_X1_286_ (
  .A1({ S12169 }),
  .A2({ S25957[414] }),
  .ZN({ S12170 })
);
AOI21_X1 #() 
AOI21_X1_758_ (
  .A({ S12000 }),
  .B1({ S12026 }),
  .B2({ S12027 }),
  .ZN({ S12172 })
);
AND2_X1 #() 
AND2_X1_75_ (
  .A1({ S12128 }),
  .A2({ S11984 }),
  .ZN({ S12173 })
);
OAI21_X1 #() 
OAI21_X1_700_ (
  .A({ S12173 }),
  .B1({ S25957[411] }),
  .B2({ S12172 }),
  .ZN({ S12174 })
);
NAND2_X1 #() 
NAND2_X1_1219_ (
  .A1({ S12090 }),
  .A2({ S37 }),
  .ZN({ S12175 })
);
NAND3_X1 #() 
NAND3_X1_1430_ (
  .A1({ S12024 }),
  .A2({ S28 }),
  .A3({ S12090 }),
  .ZN({ S12176 })
);
OAI211_X1 #() 
OAI211_X1_461_ (
  .A({ S12176 }),
  .B({ S25957[412] }),
  .C1({ S28 }),
  .C2({ S12175 }),
  .ZN({ S12177 })
);
NAND2_X1 #() 
NAND2_X1_1220_ (
  .A1({ S12099 }),
  .A2({ S12090 }),
  .ZN({ S12178 })
);
OAI21_X1 #() 
OAI21_X1_701_ (
  .A({ S12178 }),
  .B1({ S12175 }),
  .B2({ S28 }),
  .ZN({ S12179 })
);
NAND2_X1 #() 
NAND2_X1_1221_ (
  .A1({ S12179 }),
  .A2({ S11984 }),
  .ZN({ S12180 })
);
NAND2_X1 #() 
NAND2_X1_1222_ (
  .A1({ S12177 }),
  .A2({ S12180 }),
  .ZN({ S12181 })
);
NAND2_X1 #() 
NAND2_X1_1223_ (
  .A1({ S12012 }),
  .A2({ S12035 }),
  .ZN({ S12183 })
);
AOI21_X1 #() 
AOI21_X1_759_ (
  .A({ S11984 }),
  .B1({ S12159 }),
  .B2({ S25957[411] }),
  .ZN({ S12184 })
);
OAI21_X1 #() 
OAI21_X1_702_ (
  .A({ S12184 }),
  .B1({ S25957[411] }),
  .B2({ S12183 }),
  .ZN({ S12185 })
);
AND2_X1 #() 
AND2_X1_76_ (
  .A1({ S12185 }),
  .A2({ S12034 }),
  .ZN({ S12186 })
);
AOI22_X1 #() 
AOI22_X1_168_ (
  .A1({ S12181 }),
  .A2({ S25957[413] }),
  .B1({ S12186 }),
  .B2({ S12174 }),
  .ZN({ S12187 })
);
AOI22_X1 #() 
AOI22_X1_169_ (
  .A1({ S12187 }),
  .A2({ S25957[414] }),
  .B1({ S12163 }),
  .B2({ S12170 }),
  .ZN({ S12188 })
);
NAND2_X1 #() 
NAND2_X1_1224_ (
  .A1({ S12188 }),
  .A2({ S9910 }),
  .ZN({ S12189 })
);
NAND2_X1 #() 
NAND2_X1_1225_ (
  .A1({ S12189 }),
  .A2({ S12157 }),
  .ZN({ S12190 })
);
NAND2_X1 #() 
NAND2_X1_1226_ (
  .A1({ S12190 }),
  .A2({ S25957[486] }),
  .ZN({ S12191 })
);
OR2_X1 #() 
OR2_X1_17_ (
  .A1({ S12190 }),
  .A2({ S25957[486] }),
  .ZN({ S12192 })
);
NAND2_X1 #() 
NAND2_X1_1227_ (
  .A1({ S12192 }),
  .A2({ S12191 }),
  .ZN({ S25957[358] })
);
NAND2_X1 #() 
NAND2_X1_1228_ (
  .A1({ S25957[358] }),
  .A2({ S25957[454] }),
  .ZN({ S12194 })
);
INV_X1 #() 
INV_X1_395_ (
  .A({ S25957[454] }),
  .ZN({ S12195 })
);
NAND3_X1 #() 
NAND3_X1_1431_ (
  .A1({ S12192 }),
  .A2({ S12195 }),
  .A3({ S12191 }),
  .ZN({ S12196 })
);
NAND3_X1 #() 
NAND3_X1_1432_ (
  .A1({ S12194 }),
  .A2({ S12196 }),
  .A3({ S25957[518] }),
  .ZN({ S12197 })
);
NAND2_X1 #() 
NAND2_X1_1229_ (
  .A1({ S12194 }),
  .A2({ S12196 }),
  .ZN({ S12198 })
);
NAND2_X1 #() 
NAND2_X1_1230_ (
  .A1({ S12198 }),
  .A2({ S6416 }),
  .ZN({ S12199 })
);
AND2_X1 #() 
AND2_X1_77_ (
  .A1({ S12199 }),
  .A2({ S12197 }),
  .ZN({ S25957[262] })
);
NOR2_X1 #() 
NOR2_X1_287_ (
  .A1({ S9336 }),
  .A2({ S9334 }),
  .ZN({ S12200 })
);
INV_X1 #() 
INV_X1_396_ (
  .A({ S12200 }),
  .ZN({ S25957[453] })
);
NAND2_X1 #() 
NAND2_X1_1231_ (
  .A1({ S6496 }),
  .A2({ S6497 }),
  .ZN({ S25957[613] })
);
NAND2_X1 #() 
NAND2_X1_1232_ (
  .A1({ S9297 }),
  .A2({ S9333 }),
  .ZN({ S12202 })
);
XNOR2_X1 #() 
XNOR2_X1_39_ (
  .A({ S12202 }),
  .B({ S25957[613] }),
  .ZN({ S25957[485] })
);
INV_X1 #() 
INV_X1_397_ (
  .A({ S25957[485] }),
  .ZN({ S12203 })
);
NAND2_X1 #() 
NAND2_X1_1233_ (
  .A1({ S11977 }),
  .A2({ S12000 }),
  .ZN({ S12204 })
);
NAND2_X1 #() 
NAND2_X1_1234_ (
  .A1({ S12027 }),
  .A2({ S25957[410] }),
  .ZN({ S12205 })
);
AOI21_X1 #() 
AOI21_X1_760_ (
  .A({ S28 }),
  .B1({ S12204 }),
  .B2({ S12205 }),
  .ZN({ S12206 })
);
NAND3_X1 #() 
NAND3_X1_1433_ (
  .A1({ S37 }),
  .A2({ S28 }),
  .A3({ S12035 }),
  .ZN({ S12207 })
);
INV_X1 #() 
INV_X1_398_ (
  .A({ S12207 }),
  .ZN({ S12208 })
);
NOR3_X1 #() 
NOR3_X1_40_ (
  .A1({ S12206 }),
  .A2({ S12208 }),
  .A3({ S25957[412] }),
  .ZN({ S12209 })
);
NOR2_X1 #() 
NOR2_X1_288_ (
  .A1({ S28 }),
  .A2({ S25957[408] }),
  .ZN({ S12211 })
);
AOI21_X1 #() 
AOI21_X1_761_ (
  .A({ S12057 }),
  .B1({ S12040 }),
  .B2({ S12037 }),
  .ZN({ S12212 })
);
AOI21_X1 #() 
AOI21_X1_762_ (
  .A({ S12212 }),
  .B1({ S12211 }),
  .B2({ S12035 }),
  .ZN({ S12213 })
);
OAI21_X1 #() 
OAI21_X1_703_ (
  .A({ S25957[413] }),
  .B1({ S12213 }),
  .B2({ S11984 }),
  .ZN({ S12214 })
);
OAI211_X1 #() 
OAI211_X1_462_ (
  .A({ S12205 }),
  .B({ S25957[412] }),
  .C1({ S28 }),
  .C2({ S12027 }),
  .ZN({ S12215 })
);
NAND2_X1 #() 
NAND2_X1_1235_ (
  .A1({ S12173 }),
  .A2({ S12050 }),
  .ZN({ S12216 })
);
NAND3_X1 #() 
NAND3_X1_1434_ (
  .A1({ S12216 }),
  .A2({ S12034 }),
  .A3({ S12215 }),
  .ZN({ S12217 })
);
OAI211_X1 #() 
OAI211_X1_463_ (
  .A({ S25957[414] }),
  .B({ S12217 }),
  .C1({ S12214 }),
  .C2({ S12209 }),
  .ZN({ S12218 })
);
NAND2_X1 #() 
NAND2_X1_1236_ (
  .A1({ S12045 }),
  .A2({ S12077 }),
  .ZN({ S12219 })
);
AOI211_X1 #() 
AOI211_X1_18_ (
  .A({ S12047 }),
  .B({ S25957[412] }),
  .C1({ S12219 }),
  .C2({ S25957[411] }),
  .ZN({ S12220 })
);
NOR2_X1 #() 
NOR2_X1_289_ (
  .A1({ S12088 }),
  .A2({ S28 }),
  .ZN({ S12222 })
);
AOI21_X1 #() 
AOI21_X1_763_ (
  .A({ S12222 }),
  .B1({ S12092 }),
  .B2({ S12025 }),
  .ZN({ S12223 })
);
OAI21_X1 #() 
OAI21_X1_704_ (
  .A({ S12034 }),
  .B1({ S12223 }),
  .B2({ S11984 }),
  .ZN({ S12224 })
);
NAND2_X1 #() 
NAND2_X1_1237_ (
  .A1({ S12071 }),
  .A2({ S12035 }),
  .ZN({ S12225 })
);
NOR2_X1 #() 
NOR2_X1_290_ (
  .A1({ S28 }),
  .A2({ S25957[409] }),
  .ZN({ S12226 })
);
NOR2_X1 #() 
NOR2_X1_291_ (
  .A1({ S12226 }),
  .A2({ S25957[412] }),
  .ZN({ S12227 })
);
NAND2_X1 #() 
NAND2_X1_1238_ (
  .A1({ S12225 }),
  .A2({ S12227 }),
  .ZN({ S12228 })
);
OAI221_X1 #() 
OAI221_X1_28_ (
  .A({ S25957[412] }),
  .B1({ S12015 }),
  .B2({ S28 }),
  .C1({ S12006 }),
  .C2({ S36 }),
  .ZN({ S12229 })
);
NAND3_X1 #() 
NAND3_X1_1435_ (
  .A1({ S12228 }),
  .A2({ S12229 }),
  .A3({ S25957[413] }),
  .ZN({ S12230 })
);
OAI211_X1 #() 
OAI211_X1_464_ (
  .A({ S12230 }),
  .B({ S11981 }),
  .C1({ S12220 }),
  .C2({ S12224 }),
  .ZN({ S12231 })
);
NAND3_X1 #() 
NAND3_X1_1436_ (
  .A1({ S12231 }),
  .A2({ S25957[415] }),
  .A3({ S12218 }),
  .ZN({ S12233 })
);
NAND4_X1 #() 
NAND4_X1_175_ (
  .A1({ S12090 }),
  .A2({ S11995 }),
  .A3({ S25957[411] }),
  .A4({ S11996 }),
  .ZN({ S12234 })
);
INV_X1 #() 
INV_X1_399_ (
  .A({ S11995 }),
  .ZN({ S12235 })
);
NOR2_X1 #() 
NOR2_X1_292_ (
  .A1({ S12164 }),
  .A2({ S12235 }),
  .ZN({ S12236 })
);
OAI21_X1 #() 
OAI21_X1_705_ (
  .A({ S12234 }),
  .B1({ S12236 }),
  .B2({ S25957[411] }),
  .ZN({ S12237 })
);
NAND3_X1 #() 
NAND3_X1_1437_ (
  .A1({ S25957[408] }),
  .A2({ S25957[409] }),
  .A3({ S25957[410] }),
  .ZN({ S12238 })
);
NAND3_X1 #() 
NAND3_X1_1438_ (
  .A1({ S12204 }),
  .A2({ S28 }),
  .A3({ S12238 }),
  .ZN({ S12239 })
);
AOI22_X1 #() 
AOI22_X1_170_ (
  .A1({ S12237 }),
  .A2({ S11984 }),
  .B1({ S12239 }),
  .B2({ S12058 }),
  .ZN({ S12240 })
);
NAND3_X1 #() 
NAND3_X1_1439_ (
  .A1({ S12027 }),
  .A2({ S25957[411] }),
  .A3({ S12000 }),
  .ZN({ S12241 })
);
NAND4_X1 #() 
NAND4_X1_176_ (
  .A1({ S11977 }),
  .A2({ S37 }),
  .A3({ S25957[411] }),
  .A4({ S25957[410] }),
  .ZN({ S12242 })
);
NAND2_X1 #() 
NAND2_X1_1239_ (
  .A1({ S11993 }),
  .A2({ S28 }),
  .ZN({ S12244 })
);
NAND4_X1 #() 
NAND4_X1_177_ (
  .A1({ S12244 }),
  .A2({ S12242 }),
  .A3({ S12241 }),
  .A4({ S25957[412] }),
  .ZN({ S12245 })
);
INV_X1 #() 
INV_X1_400_ (
  .A({ S12211 }),
  .ZN({ S12246 })
);
OAI21_X1 #() 
OAI21_X1_706_ (
  .A({ S12246 }),
  .B1({ S12091 }),
  .B2({ S12070 }),
  .ZN({ S12247 })
);
AOI21_X1 #() 
AOI21_X1_764_ (
  .A({ S12034 }),
  .B1({ S12247 }),
  .B2({ S11984 }),
  .ZN({ S12248 })
);
AOI22_X1 #() 
AOI22_X1_171_ (
  .A1({ S12240 }),
  .A2({ S12034 }),
  .B1({ S12245 }),
  .B2({ S12248 }),
  .ZN({ S12249 })
);
NAND2_X1 #() 
NAND2_X1_1240_ (
  .A1({ S12036 }),
  .A2({ S25957[411] }),
  .ZN({ S12250 })
);
NAND2_X1 #() 
NAND2_X1_1241_ (
  .A1({ S12141 }),
  .A2({ S28 }),
  .ZN({ S12251 })
);
NAND3_X1 #() 
NAND3_X1_1440_ (
  .A1({ S12250 }),
  .A2({ S25957[412] }),
  .A3({ S12251 }),
  .ZN({ S12252 })
);
OAI211_X1 #() 
OAI211_X1_465_ (
  .A({ S11984 }),
  .B({ S12061 }),
  .C1({ S12178 }),
  .C2({ S12235 }),
  .ZN({ S12253 })
);
AOI21_X1 #() 
AOI21_X1_765_ (
  .A({ S12034 }),
  .B1({ S12252 }),
  .B2({ S12253 }),
  .ZN({ S12255 })
);
NAND2_X1 #() 
NAND2_X1_1242_ (
  .A1({ S12026 }),
  .A2({ S12000 }),
  .ZN({ S12256 })
);
AOI21_X1 #() 
AOI21_X1_766_ (
  .A({ S28 }),
  .B1({ S12045 }),
  .B2({ S12256 }),
  .ZN({ S12257 })
);
AND3_X1 #() 
AND3_X1_61_ (
  .A1({ S12045 }),
  .A2({ S28 }),
  .A3({ S12204 }),
  .ZN({ S12258 })
);
NOR3_X1 #() 
NOR3_X1_41_ (
  .A1({ S12258 }),
  .A2({ S12257 }),
  .A3({ S11984 }),
  .ZN({ S12259 })
);
INV_X1 #() 
INV_X1_401_ (
  .A({ S12238 }),
  .ZN({ S12260 })
);
AOI21_X1 #() 
AOI21_X1_767_ (
  .A({ S12078 }),
  .B1({ S28 }),
  .B2({ S12260 }),
  .ZN({ S12261 })
);
OAI21_X1 #() 
OAI21_X1_707_ (
  .A({ S12034 }),
  .B1({ S12261 }),
  .B2({ S25957[412] }),
  .ZN({ S12262 })
);
NOR2_X1 #() 
NOR2_X1_293_ (
  .A1({ S12259 }),
  .A2({ S12262 }),
  .ZN({ S12263 })
);
OAI21_X1 #() 
OAI21_X1_708_ (
  .A({ S11981 }),
  .B1({ S12263 }),
  .B2({ S12255 }),
  .ZN({ S12264 })
);
OAI21_X1 #() 
OAI21_X1_709_ (
  .A({ S12264 }),
  .B1({ S11981 }),
  .B2({ S12249 }),
  .ZN({ S12266 })
);
OR2_X1 #() 
OR2_X1_18_ (
  .A1({ S12266 }),
  .A2({ S25957[415] }),
  .ZN({ S12267 })
);
NAND3_X1 #() 
NAND3_X1_1441_ (
  .A1({ S12267 }),
  .A2({ S12203 }),
  .A3({ S12233 }),
  .ZN({ S12268 })
);
NAND2_X1 #() 
NAND2_X1_1243_ (
  .A1({ S12231 }),
  .A2({ S12218 }),
  .ZN({ S12269 })
);
NAND2_X1 #() 
NAND2_X1_1244_ (
  .A1({ S12269 }),
  .A2({ S25957[415] }),
  .ZN({ S12270 })
);
NAND2_X1 #() 
NAND2_X1_1245_ (
  .A1({ S12266 }),
  .A2({ S9910 }),
  .ZN({ S12271 })
);
NAND3_X1 #() 
NAND3_X1_1442_ (
  .A1({ S12271 }),
  .A2({ S12270 }),
  .A3({ S25957[485] }),
  .ZN({ S12272 })
);
NAND3_X1 #() 
NAND3_X1_1443_ (
  .A1({ S12268 }),
  .A2({ S25957[453] }),
  .A3({ S12272 }),
  .ZN({ S12273 })
);
NAND3_X1 #() 
NAND3_X1_1444_ (
  .A1({ S12267 }),
  .A2({ S25957[485] }),
  .A3({ S12233 }),
  .ZN({ S12274 })
);
NAND3_X1 #() 
NAND3_X1_1445_ (
  .A1({ S12271 }),
  .A2({ S12270 }),
  .A3({ S12203 }),
  .ZN({ S12275 })
);
NAND3_X1 #() 
NAND3_X1_1446_ (
  .A1({ S12274 }),
  .A2({ S12200 }),
  .A3({ S12275 }),
  .ZN({ S12277 })
);
NAND3_X1 #() 
NAND3_X1_1447_ (
  .A1({ S12273 }),
  .A2({ S12277 }),
  .A3({ S8295 }),
  .ZN({ S12278 })
);
NAND2_X1 #() 
NAND2_X1_1246_ (
  .A1({ S12268 }),
  .A2({ S12272 }),
  .ZN({ S25957[357] })
);
NAND2_X1 #() 
NAND2_X1_1247_ (
  .A1({ S25957[357] }),
  .A2({ S25957[453] }),
  .ZN({ S12279 })
);
NAND3_X1 #() 
NAND3_X1_1448_ (
  .A1({ S12268 }),
  .A2({ S12200 }),
  .A3({ S12272 }),
  .ZN({ S12280 })
);
NAND3_X1 #() 
NAND3_X1_1449_ (
  .A1({ S12279 }),
  .A2({ S12280 }),
  .A3({ S25957[517] }),
  .ZN({ S12281 })
);
AND2_X1 #() 
AND2_X1_78_ (
  .A1({ S12281 }),
  .A2({ S12278 }),
  .ZN({ S25957[261] })
);
INV_X1 #() 
INV_X1_402_ (
  .A({ S25957[548] }),
  .ZN({ S12282 })
);
NOR2_X1 #() 
NOR2_X1_294_ (
  .A1({ S9412 }),
  .A2({ S9411 }),
  .ZN({ S25957[452] })
);
XNOR2_X1 #() 
XNOR2_X1_40_ (
  .A({ S25957[452] }),
  .B({ S12282 }),
  .ZN({ S25957[420] })
);
NAND2_X1 #() 
NAND2_X1_1248_ (
  .A1({ S3840 }),
  .A2({ S3839 }),
  .ZN({ S25957[740] })
);
XNOR2_X1 #() 
XNOR2_X1_41_ (
  .A({ S6573 }),
  .B({ S25957[740] }),
  .ZN({ S25957[612] })
);
NAND3_X1 #() 
NAND3_X1_1450_ (
  .A1({ S9403 }),
  .A2({ S25957[612] }),
  .A3({ S9376 }),
  .ZN({ S12284 })
);
INV_X1 #() 
INV_X1_403_ (
  .A({ S25957[612] }),
  .ZN({ S12285 })
);
NAND3_X1 #() 
NAND3_X1_1451_ (
  .A1({ S9406 }),
  .A2({ S12285 }),
  .A3({ S9408 }),
  .ZN({ S12286 })
);
NAND2_X1 #() 
NAND2_X1_1249_ (
  .A1({ S12284 }),
  .A2({ S12286 }),
  .ZN({ S12287 })
);
NAND3_X1 #() 
NAND3_X1_1452_ (
  .A1({ S11995 }),
  .A2({ S28 }),
  .A3({ S12035 }),
  .ZN({ S12288 })
);
NAND3_X1 #() 
NAND3_X1_1453_ (
  .A1({ S12038 }),
  .A2({ S11984 }),
  .A3({ S12288 }),
  .ZN({ S12289 })
);
NAND2_X1 #() 
NAND2_X1_1250_ (
  .A1({ S12090 }),
  .A2({ S12025 }),
  .ZN({ S12290 })
);
OAI211_X1 #() 
OAI211_X1_466_ (
  .A({ S12225 }),
  .B({ S25957[412] }),
  .C1({ S28 }),
  .C2({ S12290 }),
  .ZN({ S12291 })
);
NAND3_X1 #() 
NAND3_X1_1454_ (
  .A1({ S12291 }),
  .A2({ S12034 }),
  .A3({ S12289 }),
  .ZN({ S12293 })
);
NAND3_X1 #() 
NAND3_X1_1455_ (
  .A1({ S28 }),
  .A2({ S12012 }),
  .A3({ S12011 }),
  .ZN({ S12294 })
);
NAND3_X1 #() 
NAND3_X1_1456_ (
  .A1({ S12041 }),
  .A2({ S11984 }),
  .A3({ S12294 }),
  .ZN({ S12295 })
);
OAI21_X1 #() 
OAI21_X1_710_ (
  .A({ S28 }),
  .B1({ S11996 }),
  .B2({ S25957[408] }),
  .ZN({ S12296 })
);
AOI21_X1 #() 
AOI21_X1_768_ (
  .A({ S12034 }),
  .B1({ S12058 }),
  .B2({ S12296 }),
  .ZN({ S12297 })
);
NAND2_X1 #() 
NAND2_X1_1251_ (
  .A1({ S12295 }),
  .A2({ S12297 }),
  .ZN({ S12298 })
);
NAND3_X1 #() 
NAND3_X1_1457_ (
  .A1({ S12293 }),
  .A2({ S25957[414] }),
  .A3({ S12298 }),
  .ZN({ S12299 })
);
AOI21_X1 #() 
AOI21_X1_769_ (
  .A({ S25957[411] }),
  .B1({ S12204 }),
  .B2({ S12205 }),
  .ZN({ S12300 })
);
NAND3_X1 #() 
NAND3_X1_1458_ (
  .A1({ S12150 }),
  .A2({ S25957[412] }),
  .A3({ S12083 }),
  .ZN({ S12301 })
);
NOR3_X1 #() 
NOR3_X1_42_ (
  .A1({ S12060 }),
  .A2({ S28 }),
  .A3({ S25957[409] }),
  .ZN({ S12302 })
);
AOI21_X1 #() 
AOI21_X1_770_ (
  .A({ S12000 }),
  .B1({ S12012 }),
  .B2({ S25957[409] }),
  .ZN({ S12304 })
);
OAI21_X1 #() 
OAI21_X1_711_ (
  .A({ S11984 }),
  .B1({ S12251 }),
  .B2({ S12304 }),
  .ZN({ S12305 })
);
OAI221_X1 #() 
OAI221_X1_29_ (
  .A({ S12034 }),
  .B1({ S12305 }),
  .B2({ S12302 }),
  .C1({ S12300 }),
  .C2({ S12301 }),
  .ZN({ S12306 })
);
AOI21_X1 #() 
AOI21_X1_771_ (
  .A({ S25957[411] }),
  .B1({ S12028 }),
  .B2({ S12024 }),
  .ZN({ S12307 })
);
NAND4_X1 #() 
NAND4_X1_178_ (
  .A1({ S25957[410] }),
  .A2({ S25957[409] }),
  .A3({ S10345 }),
  .A4({ S10342 }),
  .ZN({ S12308 })
);
AOI21_X1 #() 
AOI21_X1_772_ (
  .A({ S28 }),
  .B1({ S12256 }),
  .B2({ S12308 }),
  .ZN({ S12309 })
);
OR2_X1 #() 
OR2_X1_19_ (
  .A1({ S12309 }),
  .A2({ S25957[412] }),
  .ZN({ S12310 })
);
NAND2_X1 #() 
NAND2_X1_1252_ (
  .A1({ S12126 }),
  .A2({ S12141 }),
  .ZN({ S12311 })
);
OAI21_X1 #() 
OAI21_X1_712_ (
  .A({ S25957[412] }),
  .B1({ S12311 }),
  .B2({ S12078 }),
  .ZN({ S12312 })
);
OAI211_X1 #() 
OAI211_X1_467_ (
  .A({ S25957[413] }),
  .B({ S12312 }),
  .C1({ S12310 }),
  .C2({ S12307 }),
  .ZN({ S12313 })
);
NAND3_X1 #() 
NAND3_X1_1459_ (
  .A1({ S12313 }),
  .A2({ S12306 }),
  .A3({ S11981 }),
  .ZN({ S12315 })
);
NAND3_X1 #() 
NAND3_X1_1460_ (
  .A1({ S12315 }),
  .A2({ S12299 }),
  .A3({ S25957[415] }),
  .ZN({ S12316 })
);
INV_X1 #() 
INV_X1_404_ (
  .A({ S12316 }),
  .ZN({ S12317 })
);
AOI21_X1 #() 
AOI21_X1_773_ (
  .A({ S11984 }),
  .B1({ S146 }),
  .B2({ S12000 }),
  .ZN({ S12318 })
);
NAND2_X1 #() 
NAND2_X1_1253_ (
  .A1({ S12304 }),
  .A2({ S28 }),
  .ZN({ S12319 })
);
AOI21_X1 #() 
AOI21_X1_774_ (
  .A({ S25957[410] }),
  .B1({ S12026 }),
  .B2({ S12027 }),
  .ZN({ S12320 })
);
NAND2_X1 #() 
NAND2_X1_1254_ (
  .A1({ S12320 }),
  .A2({ S28 }),
  .ZN({ S12321 })
);
NAND4_X1 #() 
NAND4_X1_179_ (
  .A1({ S12321 }),
  .A2({ S12234 }),
  .A3({ S12319 }),
  .A4({ S11984 }),
  .ZN({ S12322 })
);
NAND2_X1 #() 
NAND2_X1_1255_ (
  .A1({ S12322 }),
  .A2({ S25957[413] }),
  .ZN({ S12323 })
);
NAND2_X1 #() 
NAND2_X1_1256_ (
  .A1({ S12204 }),
  .A2({ S12098 }),
  .ZN({ S12324 })
);
NAND2_X1 #() 
NAND2_X1_1257_ (
  .A1({ S12324 }),
  .A2({ S28 }),
  .ZN({ S12326 })
);
INV_X1 #() 
INV_X1_405_ (
  .A({ S12326 }),
  .ZN({ S12327 })
);
NAND2_X1 #() 
NAND2_X1_1258_ (
  .A1({ S12051 }),
  .A2({ S11984 }),
  .ZN({ S12328 })
);
OAI211_X1 #() 
OAI211_X1_468_ (
  .A({ S12096 }),
  .B({ S25957[412] }),
  .C1({ S12067 }),
  .C2({ S11991 }),
  .ZN({ S12329 })
);
OAI211_X1 #() 
OAI211_X1_469_ (
  .A({ S12329 }),
  .B({ S12034 }),
  .C1({ S12327 }),
  .C2({ S12328 }),
  .ZN({ S12330 })
);
OAI21_X1 #() 
OAI21_X1_713_ (
  .A({ S12330 }),
  .B1({ S12323 }),
  .B2({ S12318 }),
  .ZN({ S12331 })
);
NAND2_X1 #() 
NAND2_X1_1259_ (
  .A1({ S12331 }),
  .A2({ S25957[414] }),
  .ZN({ S12332 })
);
OAI211_X1 #() 
OAI211_X1_470_ (
  .A({ S37 }),
  .B({ S25957[411] }),
  .C1({ S12012 }),
  .C2({ S12000 }),
  .ZN({ S12333 })
);
INV_X1 #() 
INV_X1_406_ (
  .A({ S12333 }),
  .ZN({ S12334 })
);
AOI21_X1 #() 
AOI21_X1_775_ (
  .A({ S25957[411] }),
  .B1({ S12076 }),
  .B2({ S12077 }),
  .ZN({ S12335 })
);
OAI21_X1 #() 
OAI21_X1_714_ (
  .A({ S11984 }),
  .B1({ S12335 }),
  .B2({ S12334 }),
  .ZN({ S12337 })
);
NAND2_X1 #() 
NAND2_X1_1260_ (
  .A1({ S12014 }),
  .A2({ S12256 }),
  .ZN({ S12338 })
);
NAND3_X1 #() 
NAND3_X1_1461_ (
  .A1({ S12338 }),
  .A2({ S12225 }),
  .A3({ S25957[412] }),
  .ZN({ S12339 })
);
NAND3_X1 #() 
NAND3_X1_1462_ (
  .A1({ S12339 }),
  .A2({ S12337 }),
  .A3({ S12034 }),
  .ZN({ S12340 })
);
NAND3_X1 #() 
NAND3_X1_1463_ (
  .A1({ S11994 }),
  .A2({ S25957[412] }),
  .A3({ S12319 }),
  .ZN({ S12341 })
);
INV_X1 #() 
INV_X1_407_ (
  .A({ S12062 }),
  .ZN({ S12342 })
);
OAI21_X1 #() 
OAI21_X1_715_ (
  .A({ S11984 }),
  .B1({ S12222 }),
  .B2({ S12342 }),
  .ZN({ S12343 })
);
NAND3_X1 #() 
NAND3_X1_1464_ (
  .A1({ S12341 }),
  .A2({ S12343 }),
  .A3({ S25957[413] }),
  .ZN({ S12344 })
);
AND2_X1 #() 
AND2_X1_79_ (
  .A1({ S12344 }),
  .A2({ S11981 }),
  .ZN({ S12345 })
);
NAND2_X1 #() 
NAND2_X1_1261_ (
  .A1({ S12345 }),
  .A2({ S12340 }),
  .ZN({ S12346 })
);
AOI21_X1 #() 
AOI21_X1_776_ (
  .A({ S25957[415] }),
  .B1({ S12346 }),
  .B2({ S12332 }),
  .ZN({ S12348 })
);
OAI21_X1 #() 
OAI21_X1_716_ (
  .A({ S12287 }),
  .B1({ S12348 }),
  .B2({ S12317 }),
  .ZN({ S12349 })
);
INV_X1 #() 
INV_X1_408_ (
  .A({ S12287 }),
  .ZN({ S25957[484] })
);
AOI22_X1 #() 
AOI22_X1_172_ (
  .A1({ S12340 }),
  .A2({ S12345 }),
  .B1({ S12331 }),
  .B2({ S25957[414] }),
  .ZN({ S12350 })
);
OAI211_X1 #() 
OAI211_X1_471_ (
  .A({ S25957[484] }),
  .B({ S12316 }),
  .C1({ S12350 }),
  .C2({ S25957[415] }),
  .ZN({ S12351 })
);
AOI21_X1 #() 
AOI21_X1_777_ (
  .A({ S25957[548] }),
  .B1({ S12349 }),
  .B2({ S12351 }),
  .ZN({ S12352 })
);
OAI211_X1 #() 
OAI211_X1_472_ (
  .A({ S12287 }),
  .B({ S12316 }),
  .C1({ S12350 }),
  .C2({ S25957[415] }),
  .ZN({ S12353 })
);
OAI21_X1 #() 
OAI21_X1_717_ (
  .A({ S25957[484] }),
  .B1({ S12348 }),
  .B2({ S12317 }),
  .ZN({ S12354 })
);
AOI21_X1 #() 
AOI21_X1_778_ (
  .A({ S12282 }),
  .B1({ S12354 }),
  .B2({ S12353 }),
  .ZN({ S12355 })
);
OAI21_X1 #() 
OAI21_X1_718_ (
  .A({ S25957[388] }),
  .B1({ S12352 }),
  .B2({ S12355 }),
  .ZN({ S12356 })
);
NAND3_X1 #() 
NAND3_X1_1465_ (
  .A1({ S12354 }),
  .A2({ S12353 }),
  .A3({ S12282 }),
  .ZN({ S12358 })
);
NAND2_X1 #() 
NAND2_X1_1262_ (
  .A1({ S12354 }),
  .A2({ S12353 }),
  .ZN({ S25957[356] })
);
NAND2_X1 #() 
NAND2_X1_1263_ (
  .A1({ S25957[356] }),
  .A2({ S25957[548] }),
  .ZN({ S12359 })
);
NAND3_X1 #() 
NAND3_X1_1466_ (
  .A1({ S12359 }),
  .A2({ S11332 }),
  .A3({ S12358 }),
  .ZN({ S12360 })
);
NAND2_X1 #() 
NAND2_X1_1264_ (
  .A1({ S12360 }),
  .A2({ S12356 }),
  .ZN({ S25957[260] })
);
NAND2_X1 #() 
NAND2_X1_1265_ (
  .A1({ S9509 }),
  .A2({ S9514 }),
  .ZN({ S12361 })
);
INV_X1 #() 
INV_X1_409_ (
  .A({ S25957[579] }),
  .ZN({ S12362 })
);
NAND3_X1 #() 
NAND3_X1_1467_ (
  .A1({ S11977 }),
  .A2({ S25957[411] }),
  .A3({ S11990 }),
  .ZN({ S12363 })
);
NAND3_X1 #() 
NAND3_X1_1468_ (
  .A1({ S12087 }),
  .A2({ S28 }),
  .A3({ S11992 }),
  .ZN({ S12364 })
);
AOI21_X1 #() 
AOI21_X1_779_ (
  .A({ S11984 }),
  .B1({ S12364 }),
  .B2({ S12363 }),
  .ZN({ S12365 })
);
OAI21_X1 #() 
OAI21_X1_719_ (
  .A({ S12034 }),
  .B1({ S12328 }),
  .B2({ S12175 }),
  .ZN({ S12367 })
);
NOR2_X1 #() 
NOR2_X1_295_ (
  .A1({ S12365 }),
  .A2({ S12367 }),
  .ZN({ S12368 })
);
OAI211_X1 #() 
OAI211_X1_473_ (
  .A({ S11977 }),
  .B({ S28 }),
  .C1({ S25957[408] }),
  .C2({ S12035 }),
  .ZN({ S12369 })
);
OAI211_X1 #() 
OAI211_X1_474_ (
  .A({ S12369 }),
  .B({ S11984 }),
  .C1({ S12311 }),
  .C2({ S28 }),
  .ZN({ S12370 })
);
NAND3_X1 #() 
NAND3_X1_1469_ (
  .A1({ S12308 }),
  .A2({ S28 }),
  .A3({ S12026 }),
  .ZN({ S12371 })
);
NAND3_X1 #() 
NAND3_X1_1470_ (
  .A1({ S12371 }),
  .A2({ S12333 }),
  .A3({ S25957[412] }),
  .ZN({ S12372 })
);
AND3_X1 #() 
AND3_X1_62_ (
  .A1({ S12370 }),
  .A2({ S25957[413] }),
  .A3({ S12372 }),
  .ZN({ S12373 })
);
OAI21_X1 #() 
OAI21_X1_720_ (
  .A({ S25957[414] }),
  .B1({ S12368 }),
  .B2({ S12373 }),
  .ZN({ S12374 })
);
AND3_X1 #() 
AND3_X1_63_ (
  .A1({ S12045 }),
  .A2({ S12035 }),
  .A3({ S28 }),
  .ZN({ S12375 })
);
OAI211_X1 #() 
OAI211_X1_475_ (
  .A({ S12005 }),
  .B({ S28 }),
  .C1({ S12012 }),
  .C2({ S11996 }),
  .ZN({ S12376 })
);
OAI211_X1 #() 
OAI211_X1_476_ (
  .A({ S25957[412] }),
  .B({ S12376 }),
  .C1({ S12320 }),
  .C2({ S12002 }),
  .ZN({ S12378 })
);
NAND4_X1 #() 
NAND4_X1_180_ (
  .A1({ S12090 }),
  .A2({ S11995 }),
  .A3({ S25957[411] }),
  .A4({ S25957[409] }),
  .ZN({ S12379 })
);
NAND2_X1 #() 
NAND2_X1_1266_ (
  .A1({ S12379 }),
  .A2({ S11984 }),
  .ZN({ S12380 })
);
OAI21_X1 #() 
OAI21_X1_721_ (
  .A({ S12378 }),
  .B1({ S12375 }),
  .B2({ S12380 }),
  .ZN({ S12381 })
);
NAND2_X1 #() 
NAND2_X1_1267_ (
  .A1({ S12381 }),
  .A2({ S25957[413] }),
  .ZN({ S12382 })
);
NAND3_X1 #() 
NAND3_X1_1471_ (
  .A1({ S12087 }),
  .A2({ S25957[411] }),
  .A3({ S12035 }),
  .ZN({ S12383 })
);
AOI21_X1 #() 
AOI21_X1_780_ (
  .A({ S25957[412] }),
  .B1({ S12175 }),
  .B2({ S28 }),
  .ZN({ S12384 })
);
NAND2_X1 #() 
NAND2_X1_1268_ (
  .A1({ S12383 }),
  .A2({ S12384 }),
  .ZN({ S12385 })
);
AOI21_X1 #() 
AOI21_X1_781_ (
  .A({ S25957[410] }),
  .B1({ S11977 }),
  .B2({ S37 }),
  .ZN({ S12386 })
);
OAI211_X1 #() 
OAI211_X1_477_ (
  .A({ S25957[412] }),
  .B({ S12288 }),
  .C1({ S12386 }),
  .C2({ S28 }),
  .ZN({ S12387 })
);
NAND2_X1 #() 
NAND2_X1_1269_ (
  .A1({ S12385 }),
  .A2({ S12387 }),
  .ZN({ S12389 })
);
NAND2_X1 #() 
NAND2_X1_1270_ (
  .A1({ S12389 }),
  .A2({ S12034 }),
  .ZN({ S12390 })
);
NAND3_X1 #() 
NAND3_X1_1472_ (
  .A1({ S12390 }),
  .A2({ S12382 }),
  .A3({ S11981 }),
  .ZN({ S12391 })
);
NAND3_X1 #() 
NAND3_X1_1473_ (
  .A1({ S12391 }),
  .A2({ S12374 }),
  .A3({ S25957[415] }),
  .ZN({ S12392 })
);
OAI211_X1 #() 
OAI211_X1_478_ (
  .A({ S25957[412] }),
  .B({ S12128 }),
  .C1({ S12123 }),
  .C2({ S12172 }),
  .ZN({ S12393 })
);
NAND3_X1 #() 
NAND3_X1_1474_ (
  .A1({ S12026 }),
  .A2({ S28 }),
  .A3({ S12011 }),
  .ZN({ S12394 })
);
AOI21_X1 #() 
AOI21_X1_782_ (
  .A({ S25957[412] }),
  .B1({ S12211 }),
  .B2({ S11990 }),
  .ZN({ S12395 })
);
AOI21_X1 #() 
AOI21_X1_783_ (
  .A({ S12034 }),
  .B1({ S12395 }),
  .B2({ S12394 }),
  .ZN({ S12396 })
);
NAND2_X1 #() 
NAND2_X1_1271_ (
  .A1({ S12396 }),
  .A2({ S12393 }),
  .ZN({ S12397 })
);
OAI21_X1 #() 
OAI21_X1_722_ (
  .A({ S28 }),
  .B1({ S11991 }),
  .B2({ S12012 }),
  .ZN({ S12398 })
);
NOR2_X1 #() 
NOR2_X1_296_ (
  .A1({ S12398 }),
  .A2({ S11984 }),
  .ZN({ S12400 })
);
AOI21_X1 #() 
AOI21_X1_784_ (
  .A({ S12400 }),
  .B1({ S12338 }),
  .B2({ S12016 }),
  .ZN({ S12401 })
);
OAI211_X1 #() 
OAI211_X1_479_ (
  .A({ S12397 }),
  .B({ S25957[414] }),
  .C1({ S25957[413] }),
  .C2({ S12401 }),
  .ZN({ S12402 })
);
NAND4_X1 #() 
NAND4_X1_181_ (
  .A1({ S12098 }),
  .A2({ S12026 }),
  .A3({ S25957[411] }),
  .A4({ S12027 }),
  .ZN({ S12403 })
);
NAND2_X1 #() 
NAND2_X1_1272_ (
  .A1({ S12161 }),
  .A2({ S12403 }),
  .ZN({ S12404 })
);
NAND2_X1 #() 
NAND2_X1_1273_ (
  .A1({ S12404 }),
  .A2({ S25957[412] }),
  .ZN({ S12405 })
);
NAND2_X1 #() 
NAND2_X1_1274_ (
  .A1({ S12324 }),
  .A2({ S25957[411] }),
  .ZN({ S12406 })
);
NAND3_X1 #() 
NAND3_X1_1475_ (
  .A1({ S12406 }),
  .A2({ S12022 }),
  .A3({ S11984 }),
  .ZN({ S12407 })
);
NAND3_X1 #() 
NAND3_X1_1476_ (
  .A1({ S12407 }),
  .A2({ S12034 }),
  .A3({ S12405 }),
  .ZN({ S12408 })
);
AOI21_X1 #() 
AOI21_X1_785_ (
  .A({ S12000 }),
  .B1({ S12062 }),
  .B2({ S37 }),
  .ZN({ S12409 })
);
NAND3_X1 #() 
NAND3_X1_1477_ (
  .A1({ S28 }),
  .A2({ S12011 }),
  .A3({ S25957[408] }),
  .ZN({ S12411 })
);
OAI211_X1 #() 
OAI211_X1_480_ (
  .A({ S12411 }),
  .B({ S11984 }),
  .C1({ S12126 }),
  .C2({ S28 }),
  .ZN({ S12412 })
);
OAI21_X1 #() 
OAI21_X1_723_ (
  .A({ S12412 }),
  .B1({ S12409 }),
  .B2({ S11984 }),
  .ZN({ S12413 })
);
AOI21_X1 #() 
AOI21_X1_786_ (
  .A({ S25957[414] }),
  .B1({ S12413 }),
  .B2({ S25957[413] }),
  .ZN({ S12414 })
);
NAND2_X1 #() 
NAND2_X1_1275_ (
  .A1({ S12408 }),
  .A2({ S12414 }),
  .ZN({ S12415 })
);
NAND3_X1 #() 
NAND3_X1_1478_ (
  .A1({ S12415 }),
  .A2({ S12402 }),
  .A3({ S9910 }),
  .ZN({ S12416 })
);
NAND3_X1 #() 
NAND3_X1_1479_ (
  .A1({ S12392 }),
  .A2({ S12362 }),
  .A3({ S12416 }),
  .ZN({ S12417 })
);
NAND3_X1 #() 
NAND3_X1_1480_ (
  .A1({ S12370 }),
  .A2({ S12372 }),
  .A3({ S25957[413] }),
  .ZN({ S12418 })
);
OAI211_X1 #() 
OAI211_X1_481_ (
  .A({ S12418 }),
  .B({ S25957[414] }),
  .C1({ S12365 }),
  .C2({ S12367 }),
  .ZN({ S12419 })
);
NAND3_X1 #() 
NAND3_X1_1481_ (
  .A1({ S12385 }),
  .A2({ S12387 }),
  .A3({ S12034 }),
  .ZN({ S12420 })
);
OAI211_X1 #() 
OAI211_X1_482_ (
  .A({ S12420 }),
  .B({ S11981 }),
  .C1({ S12381 }),
  .C2({ S12034 }),
  .ZN({ S12422 })
);
NAND3_X1 #() 
NAND3_X1_1482_ (
  .A1({ S12422 }),
  .A2({ S12419 }),
  .A3({ S25957[415] }),
  .ZN({ S12423 })
);
INV_X1 #() 
INV_X1_410_ (
  .A({ S12338 }),
  .ZN({ S12424 })
);
NOR2_X1 #() 
NOR2_X1_297_ (
  .A1({ S12400 }),
  .A2({ S25957[413] }),
  .ZN({ S12425 })
);
OAI21_X1 #() 
OAI21_X1_724_ (
  .A({ S12425 }),
  .B1({ S12424 }),
  .B2({ S12017 }),
  .ZN({ S12426 })
);
AOI22_X1 #() 
AOI22_X1_173_ (
  .A1({ S12048 }),
  .A2({ S12128 }),
  .B1({ S12395 }),
  .B2({ S12394 }),
  .ZN({ S12427 })
);
OAI211_X1 #() 
OAI211_X1_483_ (
  .A({ S12426 }),
  .B({ S25957[414] }),
  .C1({ S12427 }),
  .C2({ S12034 }),
  .ZN({ S12428 })
);
AOI21_X1 #() 
AOI21_X1_787_ (
  .A({ S25957[412] }),
  .B1({ S12406 }),
  .B2({ S12022 }),
  .ZN({ S12429 })
);
NAND3_X1 #() 
NAND3_X1_1483_ (
  .A1({ S12161 }),
  .A2({ S25957[412] }),
  .A3({ S12403 }),
  .ZN({ S12430 })
);
NAND2_X1 #() 
NAND2_X1_1276_ (
  .A1({ S12430 }),
  .A2({ S12034 }),
  .ZN({ S12431 })
);
OAI211_X1 #() 
OAI211_X1_484_ (
  .A({ S12412 }),
  .B({ S25957[413] }),
  .C1({ S12409 }),
  .C2({ S11984 }),
  .ZN({ S12433 })
);
OAI211_X1 #() 
OAI211_X1_485_ (
  .A({ S11981 }),
  .B({ S12433 }),
  .C1({ S12429 }),
  .C2({ S12431 }),
  .ZN({ S12434 })
);
NAND3_X1 #() 
NAND3_X1_1484_ (
  .A1({ S12428 }),
  .A2({ S12434 }),
  .A3({ S9910 }),
  .ZN({ S12435 })
);
NAND3_X1 #() 
NAND3_X1_1485_ (
  .A1({ S12435 }),
  .A2({ S12423 }),
  .A3({ S25957[579] }),
  .ZN({ S12436 })
);
AOI21_X1 #() 
AOI21_X1_788_ (
  .A({ S12361 }),
  .B1({ S12417 }),
  .B2({ S12436 }),
  .ZN({ S12437 })
);
AND3_X1 #() 
AND3_X1_64_ (
  .A1({ S12417 }),
  .A2({ S12361 }),
  .A3({ S12436 }),
  .ZN({ S12438 })
);
OAI21_X1 #() 
OAI21_X1_725_ (
  .A({ S24 }),
  .B1({ S12438 }),
  .B2({ S12437 }),
  .ZN({ S12439 })
);
INV_X1 #() 
INV_X1_411_ (
  .A({ S12361 }),
  .ZN({ S25957[419] })
);
AOI21_X1 #() 
AOI21_X1_789_ (
  .A({ S25957[579] }),
  .B1({ S12435 }),
  .B2({ S12423 }),
  .ZN({ S12440 })
);
INV_X1 #() 
INV_X1_412_ (
  .A({ S12436 }),
  .ZN({ S12441 })
);
OAI21_X1 #() 
OAI21_X1_726_ (
  .A({ S25957[419] }),
  .B1({ S12441 }),
  .B2({ S12440 }),
  .ZN({ S12443 })
);
NAND3_X1 #() 
NAND3_X1_1486_ (
  .A1({ S12417 }),
  .A2({ S12361 }),
  .A3({ S12436 }),
  .ZN({ S12444 })
);
NAND3_X1 #() 
NAND3_X1_1487_ (
  .A1({ S12443 }),
  .A2({ S25957[387] }),
  .A3({ S12444 }),
  .ZN({ S12445 })
);
NAND2_X1 #() 
NAND2_X1_1277_ (
  .A1({ S12439 }),
  .A2({ S12445 }),
  .ZN({ S38 })
);
NAND3_X1 #() 
NAND3_X1_1488_ (
  .A1({ S12443 }),
  .A2({ S24 }),
  .A3({ S12444 }),
  .ZN({ S12446 })
);
OAI21_X1 #() 
OAI21_X1_727_ (
  .A({ S25957[387] }),
  .B1({ S12438 }),
  .B2({ S12437 }),
  .ZN({ S12447 })
);
NAND2_X1 #() 
NAND2_X1_1278_ (
  .A1({ S12447 }),
  .A2({ S12446 }),
  .ZN({ S25957[259] })
);
NAND2_X1 #() 
NAND2_X1_1279_ (
  .A1({ S6752 }),
  .A2({ S6748 }),
  .ZN({ S25957[544] })
);
NOR2_X1 #() 
NOR2_X1_298_ (
  .A1({ S9579 }),
  .A2({ S9580 }),
  .ZN({ S12448 })
);
XNOR2_X1 #() 
XNOR2_X1_42_ (
  .A({ S12448 }),
  .B({ S25957[544] }),
  .ZN({ S25957[416] })
);
INV_X1 #() 
INV_X1_413_ (
  .A({ S12448 }),
  .ZN({ S25957[448] })
);
NAND2_X1 #() 
NAND2_X1_1280_ (
  .A1({ S6755 }),
  .A2({ S6757 }),
  .ZN({ S12450 })
);
NAND3_X1 #() 
NAND3_X1_1489_ (
  .A1({ S9578 }),
  .A2({ S9549 }),
  .A3({ S12450 }),
  .ZN({ S12451 })
);
INV_X1 #() 
INV_X1_414_ (
  .A({ S12450 }),
  .ZN({ S25957[608] })
);
NAND3_X1 #() 
NAND3_X1_1490_ (
  .A1({ S9587 }),
  .A2({ S9612 }),
  .A3({ S25957[608] }),
  .ZN({ S12452 })
);
NAND2_X1 #() 
NAND2_X1_1281_ (
  .A1({ S12452 }),
  .A2({ S12451 }),
  .ZN({ S25957[480] })
);
NAND3_X1 #() 
NAND3_X1_1491_ (
  .A1({ S12012 }),
  .A2({ S12025 }),
  .A3({ S25957[410] }),
  .ZN({ S12453 })
);
AOI21_X1 #() 
AOI21_X1_790_ (
  .A({ S28 }),
  .B1({ S12453 }),
  .B2({ S12005 }),
  .ZN({ S12454 })
);
AOI21_X1 #() 
AOI21_X1_791_ (
  .A({ S25957[411] }),
  .B1({ S12308 }),
  .B2({ S12090 }),
  .ZN({ S12455 })
);
OAI21_X1 #() 
OAI21_X1_728_ (
  .A({ S11984 }),
  .B1({ S12454 }),
  .B2({ S12455 }),
  .ZN({ S12456 })
);
NAND2_X1 #() 
NAND2_X1_1282_ (
  .A1({ S12321 }),
  .A2({ S12144 }),
  .ZN({ S12458 })
);
AOI21_X1 #() 
AOI21_X1_792_ (
  .A({ S25957[413] }),
  .B1({ S12456 }),
  .B2({ S12458 }),
  .ZN({ S12459 })
);
NAND3_X1 #() 
NAND3_X1_1492_ (
  .A1({ S28 }),
  .A2({ S12012 }),
  .A3({ S11990 }),
  .ZN({ S12460 })
);
NAND2_X1 #() 
NAND2_X1_1283_ (
  .A1({ S12398 }),
  .A2({ S12002 }),
  .ZN({ S12461 })
);
AOI21_X1 #() 
AOI21_X1_793_ (
  .A({ S11984 }),
  .B1({ S12461 }),
  .B2({ S12460 }),
  .ZN({ S12462 })
);
NAND2_X1 #() 
NAND2_X1_1284_ (
  .A1({ S12296 }),
  .A2({ S11984 }),
  .ZN({ S12463 })
);
OAI21_X1 #() 
OAI21_X1_729_ (
  .A({ S25957[413] }),
  .B1({ S12309 }),
  .B2({ S12463 }),
  .ZN({ S12464 })
);
OAI21_X1 #() 
OAI21_X1_730_ (
  .A({ S11981 }),
  .B1({ S12464 }),
  .B2({ S12462 }),
  .ZN({ S12465 })
);
AOI21_X1 #() 
AOI21_X1_794_ (
  .A({ S25957[411] }),
  .B1({ S12015 }),
  .B2({ S12027 }),
  .ZN({ S12466 })
);
OAI21_X1 #() 
OAI21_X1_731_ (
  .A({ S11984 }),
  .B1({ S12013 }),
  .B2({ S12057 }),
  .ZN({ S12467 })
);
NOR2_X1 #() 
NOR2_X1_299_ (
  .A1({ S12467 }),
  .A2({ S12466 }),
  .ZN({ S12469 })
);
OAI21_X1 #() 
OAI21_X1_732_ (
  .A({ S25957[412] }),
  .B1({ S12205 }),
  .B2({ S28 }),
  .ZN({ S12470 })
);
OAI21_X1 #() 
OAI21_X1_733_ (
  .A({ S25957[413] }),
  .B1({ S12335 }),
  .B2({ S12470 }),
  .ZN({ S12471 })
);
NAND3_X1 #() 
NAND3_X1_1493_ (
  .A1({ S12234 }),
  .A2({ S12251 }),
  .A3({ S11984 }),
  .ZN({ S12472 })
);
NAND4_X1 #() 
NAND4_X1_182_ (
  .A1({ S12026 }),
  .A2({ S12027 }),
  .A3({ S25957[411] }),
  .A4({ S25957[410] }),
  .ZN({ S12473 })
);
AOI21_X1 #() 
AOI21_X1_795_ (
  .A({ S11984 }),
  .B1({ S11991 }),
  .B2({ S28 }),
  .ZN({ S12474 })
);
NAND3_X1 #() 
NAND3_X1_1494_ (
  .A1({ S12473 }),
  .A2({ S12376 }),
  .A3({ S12474 }),
  .ZN({ S12475 })
);
NAND3_X1 #() 
NAND3_X1_1495_ (
  .A1({ S12475 }),
  .A2({ S12472 }),
  .A3({ S12034 }),
  .ZN({ S12476 })
);
OAI211_X1 #() 
OAI211_X1_486_ (
  .A({ S12476 }),
  .B({ S25957[414] }),
  .C1({ S12471 }),
  .C2({ S12469 }),
  .ZN({ S12477 })
);
OAI211_X1 #() 
OAI211_X1_487_ (
  .A({ S12477 }),
  .B({ S25957[415] }),
  .C1({ S12465 }),
  .C2({ S12459 }),
  .ZN({ S12478 })
);
OAI211_X1 #() 
OAI211_X1_488_ (
  .A({ S12333 }),
  .B({ S25957[412] }),
  .C1({ S12070 }),
  .C2({ S12091 }),
  .ZN({ S12480 })
);
NAND2_X1 #() 
NAND2_X1_1285_ (
  .A1({ S12133 }),
  .A2({ S11984 }),
  .ZN({ S12481 })
);
OAI211_X1 #() 
OAI211_X1_489_ (
  .A({ S25957[413] }),
  .B({ S12480 }),
  .C1({ S12258 }),
  .C2({ S12481 }),
  .ZN({ S12482 })
);
OAI211_X1 #() 
OAI211_X1_490_ (
  .A({ S12050 }),
  .B({ S12474 }),
  .C1({ S12386 }),
  .C2({ S28 }),
  .ZN({ S12483 })
);
NAND4_X1 #() 
NAND4_X1_183_ (
  .A1({ S12026 }),
  .A2({ S12090 }),
  .A3({ S25957[411] }),
  .A4({ S12027 }),
  .ZN({ S12484 })
);
OAI211_X1 #() 
OAI211_X1_491_ (
  .A({ S12484 }),
  .B({ S11984 }),
  .C1({ S12057 }),
  .C2({ S12067 }),
  .ZN({ S12485 })
);
NAND3_X1 #() 
NAND3_X1_1496_ (
  .A1({ S12485 }),
  .A2({ S12483 }),
  .A3({ S12034 }),
  .ZN({ S12486 })
);
NAND3_X1 #() 
NAND3_X1_1497_ (
  .A1({ S12482 }),
  .A2({ S12486 }),
  .A3({ S11981 }),
  .ZN({ S12487 })
);
AOI21_X1 #() 
AOI21_X1_796_ (
  .A({ S25957[412] }),
  .B1({ S12005 }),
  .B2({ S28 }),
  .ZN({ S12488 })
);
AOI21_X1 #() 
AOI21_X1_797_ (
  .A({ S28 }),
  .B1({ S11977 }),
  .B2({ S12000 }),
  .ZN({ S12489 })
);
AOI21_X1 #() 
AOI21_X1_798_ (
  .A({ S11984 }),
  .B1({ S12489 }),
  .B2({ S12087 }),
  .ZN({ S12491 })
);
NAND2_X1 #() 
NAND2_X1_1286_ (
  .A1({ S12183 }),
  .A2({ S28 }),
  .ZN({ S12492 })
);
AOI22_X1 #() 
AOI22_X1_174_ (
  .A1({ S12491 }),
  .A2({ S12492 }),
  .B1({ S12165 }),
  .B2({ S12488 }),
  .ZN({ S12493 })
);
NAND3_X1 #() 
NAND3_X1_1498_ (
  .A1({ S12234 }),
  .A2({ S11984 }),
  .A3({ S12207 }),
  .ZN({ S12494 })
);
NAND4_X1 #() 
NAND4_X1_184_ (
  .A1({ S12246 }),
  .A2({ S12141 }),
  .A3({ S25957[412] }),
  .A4({ S11996 }),
  .ZN({ S12495 })
);
NAND3_X1 #() 
NAND3_X1_1499_ (
  .A1({ S12495 }),
  .A2({ S12034 }),
  .A3({ S12494 }),
  .ZN({ S12496 })
);
OAI211_X1 #() 
OAI211_X1_492_ (
  .A({ S25957[414] }),
  .B({ S12496 }),
  .C1({ S12493 }),
  .C2({ S12034 }),
  .ZN({ S12497 })
);
NAND3_X1 #() 
NAND3_X1_1500_ (
  .A1({ S12497 }),
  .A2({ S9910 }),
  .A3({ S12487 }),
  .ZN({ S12498 })
);
NAND3_X1 #() 
NAND3_X1_1501_ (
  .A1({ S12498 }),
  .A2({ S12478 }),
  .A3({ S25957[480] }),
  .ZN({ S12499 })
);
INV_X1 #() 
INV_X1_415_ (
  .A({ S25957[480] }),
  .ZN({ S12500 })
);
NAND2_X1 #() 
NAND2_X1_1287_ (
  .A1({ S12498 }),
  .A2({ S12478 }),
  .ZN({ S12502 })
);
NAND2_X1 #() 
NAND2_X1_1288_ (
  .A1({ S12502 }),
  .A2({ S12500 }),
  .ZN({ S12503 })
);
NAND3_X1 #() 
NAND3_X1_1502_ (
  .A1({ S12503 }),
  .A2({ S25957[448] }),
  .A3({ S12499 }),
  .ZN({ S12504 })
);
NAND2_X1 #() 
NAND2_X1_1289_ (
  .A1({ S12502 }),
  .A2({ S25957[480] }),
  .ZN({ S12505 })
);
NAND3_X1 #() 
NAND3_X1_1503_ (
  .A1({ S12498 }),
  .A2({ S12478 }),
  .A3({ S12500 }),
  .ZN({ S12506 })
);
NAND3_X1 #() 
NAND3_X1_1504_ (
  .A1({ S12505 }),
  .A2({ S12448 }),
  .A3({ S12506 }),
  .ZN({ S12507 })
);
NAND3_X1 #() 
NAND3_X1_1505_ (
  .A1({ S12504 }),
  .A2({ S12507 }),
  .A3({ S25957[416] }),
  .ZN({ S12508 })
);
INV_X1 #() 
INV_X1_416_ (
  .A({ S25957[416] }),
  .ZN({ S12509 })
);
NAND3_X1 #() 
NAND3_X1_1506_ (
  .A1({ S12505 }),
  .A2({ S25957[448] }),
  .A3({ S12506 }),
  .ZN({ S12510 })
);
NAND3_X1 #() 
NAND3_X1_1507_ (
  .A1({ S12503 }),
  .A2({ S12448 }),
  .A3({ S12499 }),
  .ZN({ S12511 })
);
NAND3_X1 #() 
NAND3_X1_1508_ (
  .A1({ S12510 }),
  .A2({ S12511 }),
  .A3({ S12509 }),
  .ZN({ S12513 })
);
NAND3_X1 #() 
NAND3_X1_1509_ (
  .A1({ S12508 }),
  .A2({ S12513 }),
  .A3({ S11300 }),
  .ZN({ S12514 })
);
NAND3_X1 #() 
NAND3_X1_1510_ (
  .A1({ S12510 }),
  .A2({ S12511 }),
  .A3({ S25957[416] }),
  .ZN({ S12515 })
);
NAND3_X1 #() 
NAND3_X1_1511_ (
  .A1({ S12504 }),
  .A2({ S12507 }),
  .A3({ S12509 }),
  .ZN({ S12516 })
);
NAND3_X1 #() 
NAND3_X1_1512_ (
  .A1({ S12515 }),
  .A2({ S12516 }),
  .A3({ S25957[384] }),
  .ZN({ S12517 })
);
NAND2_X1 #() 
NAND2_X1_1290_ (
  .A1({ S12514 }),
  .A2({ S12517 }),
  .ZN({ S25957[256] })
);
NOR2_X1 #() 
NOR2_X1_300_ (
  .A1({ S11288 }),
  .A2({ S11289 }),
  .ZN({ S12518 })
);
INV_X1 #() 
INV_X1_417_ (
  .A({ S12518 }),
  .ZN({ S25957[449] })
);
NAND2_X1 #() 
NAND2_X1_1291_ (
  .A1({ S6819 }),
  .A2({ S6818 }),
  .ZN({ S25957[609] })
);
NAND2_X1 #() 
NAND2_X1_1292_ (
  .A1({ S9637 }),
  .A2({ S9656 }),
  .ZN({ S12519 })
);
OR2_X1 #() 
OR2_X1_20_ (
  .A1({ S12519 }),
  .A2({ S25957[609] }),
  .ZN({ S12521 })
);
NAND2_X1 #() 
NAND2_X1_1293_ (
  .A1({ S12519 }),
  .A2({ S25957[609] }),
  .ZN({ S12522 })
);
NAND2_X1 #() 
NAND2_X1_1294_ (
  .A1({ S12521 }),
  .A2({ S12522 }),
  .ZN({ S25957[481] })
);
AOI21_X1 #() 
AOI21_X1_799_ (
  .A({ S28 }),
  .B1({ S12087 }),
  .B2({ S12005 }),
  .ZN({ S12523 })
);
OAI21_X1 #() 
OAI21_X1_734_ (
  .A({ S25957[412] }),
  .B1({ S12523 }),
  .B2({ S12007 }),
  .ZN({ S12524 })
);
INV_X1 #() 
INV_X1_418_ (
  .A({ S37 }),
  .ZN({ S12525 })
);
OAI211_X1 #() 
OAI211_X1_493_ (
  .A({ S12241 }),
  .B({ S11984 }),
  .C1({ S12525 }),
  .C2({ S12037 }),
  .ZN({ S12526 })
);
AOI21_X1 #() 
AOI21_X1_800_ (
  .A({ S12034 }),
  .B1({ S12524 }),
  .B2({ S12526 }),
  .ZN({ S12527 })
);
NAND3_X1 #() 
NAND3_X1_1513_ (
  .A1({ S12141 }),
  .A2({ S28 }),
  .A3({ S11996 }),
  .ZN({ S12528 })
);
AOI21_X1 #() 
AOI21_X1_801_ (
  .A({ S25957[413] }),
  .B1({ S12184 }),
  .B2({ S12528 }),
  .ZN({ S12529 })
);
OAI21_X1 #() 
OAI21_X1_735_ (
  .A({ S12529 }),
  .B1({ S12029 }),
  .B2({ S12305 }),
  .ZN({ S12531 })
);
NAND2_X1 #() 
NAND2_X1_1295_ (
  .A1({ S12531 }),
  .A2({ S11981 }),
  .ZN({ S12532 })
);
NAND4_X1 #() 
NAND4_X1_185_ (
  .A1({ S12242 }),
  .A2({ S12241 }),
  .A3({ S25957[412] }),
  .A4({ S12460 }),
  .ZN({ S12533 })
);
AOI22_X1 #() 
AOI22_X1_175_ (
  .A1({ S12000 }),
  .A2({ S12025 }),
  .B1({ S10342 }),
  .B2({ S10345 }),
  .ZN({ S12534 })
);
NAND3_X1 #() 
NAND3_X1_1514_ (
  .A1({ S11977 }),
  .A2({ S25957[411] }),
  .A3({ S11995 }),
  .ZN({ S12535 })
);
OAI211_X1 #() 
OAI211_X1_494_ (
  .A({ S12535 }),
  .B({ S11984 }),
  .C1({ S12102 }),
  .C2({ S12534 }),
  .ZN({ S12536 })
);
NAND3_X1 #() 
NAND3_X1_1515_ (
  .A1({ S12533 }),
  .A2({ S12536 }),
  .A3({ S12034 }),
  .ZN({ S12537 })
);
NAND3_X1 #() 
NAND3_X1_1516_ (
  .A1({ S12005 }),
  .A2({ S25957[411] }),
  .A3({ S12035 }),
  .ZN({ S12538 })
);
NOR2_X1 #() 
NOR2_X1_301_ (
  .A1({ S12021 }),
  .A2({ S12538 }),
  .ZN({ S12539 })
);
NAND3_X1 #() 
NAND3_X1_1517_ (
  .A1({ S12363 }),
  .A2({ S25957[412] }),
  .A3({ S11997 }),
  .ZN({ S12540 })
);
NAND3_X1 #() 
NAND3_X1_1518_ (
  .A1({ S12037 }),
  .A2({ S12040 }),
  .A3({ S11984 }),
  .ZN({ S12542 })
);
OAI211_X1 #() 
OAI211_X1_495_ (
  .A({ S12540 }),
  .B({ S25957[413] }),
  .C1({ S12539 }),
  .C2({ S12542 }),
  .ZN({ S12543 })
);
NAND3_X1 #() 
NAND3_X1_1519_ (
  .A1({ S12543 }),
  .A2({ S12537 }),
  .A3({ S25957[414] }),
  .ZN({ S12544 })
);
OAI211_X1 #() 
OAI211_X1_496_ (
  .A({ S12544 }),
  .B({ S25957[415] }),
  .C1({ S12527 }),
  .C2({ S12532 }),
  .ZN({ S12545 })
);
OAI21_X1 #() 
OAI21_X1_736_ (
  .A({ S25957[412] }),
  .B1({ S12021 }),
  .B2({ S12538 }),
  .ZN({ S12546 })
);
NOR2_X1 #() 
NOR2_X1_302_ (
  .A1({ S12260 }),
  .A2({ S12102 }),
  .ZN({ S12547 })
);
NAND3_X1 #() 
NAND3_X1_1520_ (
  .A1({ S12176 }),
  .A2({ S11984 }),
  .A3({ S12473 }),
  .ZN({ S12548 })
);
OAI211_X1 #() 
OAI211_X1_497_ (
  .A({ S12548 }),
  .B({ S12034 }),
  .C1({ S12546 }),
  .C2({ S12547 }),
  .ZN({ S12549 })
);
NAND3_X1 #() 
NAND3_X1_1521_ (
  .A1({ S12453 }),
  .A2({ S28 }),
  .A3({ S12090 }),
  .ZN({ S12550 })
);
NAND3_X1 #() 
NAND3_X1_1522_ (
  .A1({ S12550 }),
  .A2({ S25957[412] }),
  .A3({ S12403 }),
  .ZN({ S12551 })
);
AOI21_X1 #() 
AOI21_X1_802_ (
  .A({ S12060 }),
  .B1({ S11991 }),
  .B2({ S12012 }),
  .ZN({ S12553 })
);
AOI21_X1 #() 
AOI21_X1_803_ (
  .A({ S12034 }),
  .B1({ S12227 }),
  .B2({ S12553 }),
  .ZN({ S12554 })
);
AOI21_X1 #() 
AOI21_X1_804_ (
  .A({ S11981 }),
  .B1({ S12554 }),
  .B2({ S12551 }),
  .ZN({ S12555 })
);
NAND2_X1 #() 
NAND2_X1_1296_ (
  .A1({ S12549 }),
  .A2({ S12555 }),
  .ZN({ S12556 })
);
AOI21_X1 #() 
AOI21_X1_805_ (
  .A({ S11984 }),
  .B1({ S12379 }),
  .B2({ S12294 }),
  .ZN({ S12557 })
);
OAI21_X1 #() 
OAI21_X1_737_ (
  .A({ S25957[413] }),
  .B1({ S12557 }),
  .B2({ S12016 }),
  .ZN({ S12558 })
);
NAND3_X1 #() 
NAND3_X1_1523_ (
  .A1({ S12096 }),
  .A2({ S25957[412] }),
  .A3({ S12288 }),
  .ZN({ S12559 })
);
NAND4_X1 #() 
NAND4_X1_186_ (
  .A1({ S28 }),
  .A2({ S12011 }),
  .A3({ S11996 }),
  .A4({ S25957[408] }),
  .ZN({ S12560 })
);
NAND3_X1 #() 
NAND3_X1_1524_ (
  .A1({ S12560 }),
  .A2({ S11984 }),
  .A3({ S12083 }),
  .ZN({ S12561 })
);
NAND3_X1 #() 
NAND3_X1_1525_ (
  .A1({ S12559 }),
  .A2({ S12034 }),
  .A3({ S12561 }),
  .ZN({ S12562 })
);
NAND3_X1 #() 
NAND3_X1_1526_ (
  .A1({ S12558 }),
  .A2({ S12562 }),
  .A3({ S11981 }),
  .ZN({ S12564 })
);
NAND3_X1 #() 
NAND3_X1_1527_ (
  .A1({ S12556 }),
  .A2({ S9910 }),
  .A3({ S12564 }),
  .ZN({ S12565 })
);
NAND3_X1 #() 
NAND3_X1_1528_ (
  .A1({ S12545 }),
  .A2({ S12565 }),
  .A3({ S25957[481] }),
  .ZN({ S12566 })
);
INV_X1 #() 
INV_X1_419_ (
  .A({ S25957[481] }),
  .ZN({ S12567 })
);
NAND2_X1 #() 
NAND2_X1_1297_ (
  .A1({ S12545 }),
  .A2({ S12565 }),
  .ZN({ S12568 })
);
NAND2_X1 #() 
NAND2_X1_1298_ (
  .A1({ S12568 }),
  .A2({ S12567 }),
  .ZN({ S12569 })
);
NAND3_X1 #() 
NAND3_X1_1529_ (
  .A1({ S12569 }),
  .A2({ S25957[449] }),
  .A3({ S12566 }),
  .ZN({ S12570 })
);
NAND2_X1 #() 
NAND2_X1_1299_ (
  .A1({ S12568 }),
  .A2({ S25957[481] }),
  .ZN({ S12571 })
);
NAND3_X1 #() 
NAND3_X1_1530_ (
  .A1({ S12545 }),
  .A2({ S12565 }),
  .A3({ S12567 }),
  .ZN({ S12572 })
);
NAND3_X1 #() 
NAND3_X1_1531_ (
  .A1({ S12571 }),
  .A2({ S12518 }),
  .A3({ S12572 }),
  .ZN({ S12573 })
);
NAND3_X1 #() 
NAND3_X1_1532_ (
  .A1({ S12570 }),
  .A2({ S12573 }),
  .A3({ S25957[513] }),
  .ZN({ S12575 })
);
NAND3_X1 #() 
NAND3_X1_1533_ (
  .A1({ S12571 }),
  .A2({ S25957[449] }),
  .A3({ S12572 }),
  .ZN({ S12576 })
);
NAND3_X1 #() 
NAND3_X1_1534_ (
  .A1({ S12569 }),
  .A2({ S12518 }),
  .A3({ S12566 }),
  .ZN({ S12577 })
);
NAND3_X1 #() 
NAND3_X1_1535_ (
  .A1({ S12576 }),
  .A2({ S12577 }),
  .A3({ S8341 }),
  .ZN({ S12578 })
);
AND2_X1 #() 
AND2_X1_80_ (
  .A1({ S12578 }),
  .A2({ S12575 }),
  .ZN({ S25957[257] })
);
NAND2_X1 #() 
NAND2_X1_1300_ (
  .A1({ S6887 }),
  .A2({ S6901 }),
  .ZN({ S25957[546] })
);
NOR2_X1 #() 
NOR2_X1_303_ (
  .A1({ S9780 }),
  .A2({ S9756 }),
  .ZN({ S25957[450] })
);
AND2_X1 #() 
AND2_X1_81_ (
  .A1({ S25957[450] }),
  .A2({ S25957[546] }),
  .ZN({ S12579 })
);
NOR2_X1 #() 
NOR2_X1_304_ (
  .A1({ S25957[450] }),
  .A2({ S25957[546] }),
  .ZN({ S12580 })
);
NOR2_X1 #() 
NOR2_X1_305_ (
  .A1({ S12579 }),
  .A2({ S12580 }),
  .ZN({ S25957[418] })
);
NAND2_X1 #() 
NAND2_X1_1301_ (
  .A1({ S4108 }),
  .A2({ S4129 }),
  .ZN({ S12582 })
);
XNOR2_X1 #() 
XNOR2_X1_43_ (
  .A({ S12582 }),
  .B({ S25957[866] }),
  .ZN({ S12583 })
);
INV_X1 #() 
INV_X1_420_ (
  .A({ S12583 }),
  .ZN({ S25957[738] })
);
NAND2_X1 #() 
NAND2_X1_1302_ (
  .A1({ S6884 }),
  .A2({ S6857 }),
  .ZN({ S12584 })
);
XNOR2_X1 #() 
XNOR2_X1_44_ (
  .A({ S12584 }),
  .B({ S25957[738] }),
  .ZN({ S25957[610] })
);
NAND2_X1 #() 
NAND2_X1_1303_ (
  .A1({ S9755 }),
  .A2({ S9727 }),
  .ZN({ S12585 })
);
NAND2_X1 #() 
NAND2_X1_1304_ (
  .A1({ S12585 }),
  .A2({ S25957[610] }),
  .ZN({ S12586 })
);
OR2_X1 #() 
OR2_X1_21_ (
  .A1({ S12585 }),
  .A2({ S25957[610] }),
  .ZN({ S12587 })
);
NAND2_X1 #() 
NAND2_X1_1305_ (
  .A1({ S12587 }),
  .A2({ S12586 }),
  .ZN({ S12588 })
);
INV_X1 #() 
INV_X1_421_ (
  .A({ S12588 }),
  .ZN({ S25957[482] })
);
NAND3_X1 #() 
NAND3_X1_1536_ (
  .A1({ S12088 }),
  .A2({ S25957[411] }),
  .A3({ S12205 }),
  .ZN({ S12590 })
);
NAND3_X1 #() 
NAND3_X1_1537_ (
  .A1({ S12590 }),
  .A2({ S11984 }),
  .A3({ S12037 }),
  .ZN({ S12591 })
);
NAND3_X1 #() 
NAND3_X1_1538_ (
  .A1({ S12290 }),
  .A2({ S28 }),
  .A3({ S12001 }),
  .ZN({ S12592 })
);
NAND2_X1 #() 
NAND2_X1_1306_ (
  .A1({ S11995 }),
  .A2({ S12035 }),
  .ZN({ S12593 })
);
AOI21_X1 #() 
AOI21_X1_806_ (
  .A({ S11984 }),
  .B1({ S12593 }),
  .B2({ S25957[411] }),
  .ZN({ S12594 })
);
AOI21_X1 #() 
AOI21_X1_807_ (
  .A({ S12034 }),
  .B1({ S12594 }),
  .B2({ S12592 }),
  .ZN({ S12595 })
);
NAND2_X1 #() 
NAND2_X1_1307_ (
  .A1({ S12595 }),
  .A2({ S12591 }),
  .ZN({ S12596 })
);
OAI211_X1 #() 
OAI211_X1_498_ (
  .A({ S12038 }),
  .B({ S11984 }),
  .C1({ S25957[411] }),
  .C2({ S12035 }),
  .ZN({ S12597 })
);
NAND2_X1 #() 
NAND2_X1_1308_ (
  .A1({ S37 }),
  .A2({ S11996 }),
  .ZN({ S12598 })
);
AOI21_X1 #() 
AOI21_X1_808_ (
  .A({ S11984 }),
  .B1({ S12598 }),
  .B2({ S28 }),
  .ZN({ S12599 })
);
NAND4_X1 #() 
NAND4_X1_187_ (
  .A1({ S12015 }),
  .A2({ S12027 }),
  .A3({ S25957[411] }),
  .A4({ S11995 }),
  .ZN({ S12601 })
);
AOI21_X1 #() 
AOI21_X1_809_ (
  .A({ S25957[413] }),
  .B1({ S12601 }),
  .B2({ S12599 }),
  .ZN({ S12602 })
);
NAND2_X1 #() 
NAND2_X1_1309_ (
  .A1({ S12602 }),
  .A2({ S12597 }),
  .ZN({ S12603 })
);
NAND3_X1 #() 
NAND3_X1_1539_ (
  .A1({ S12596 }),
  .A2({ S12603 }),
  .A3({ S25957[414] }),
  .ZN({ S12604 })
);
NAND2_X1 #() 
NAND2_X1_1310_ (
  .A1({ S12534 }),
  .A2({ S25957[411] }),
  .ZN({ S12605 })
);
NAND3_X1 #() 
NAND3_X1_1540_ (
  .A1({ S12605 }),
  .A2({ S12560 }),
  .A3({ S25957[412] }),
  .ZN({ S12606 })
);
OAI211_X1 #() 
OAI211_X1_499_ (
  .A({ S12027 }),
  .B({ S25957[411] }),
  .C1({ S12012 }),
  .C2({ S11996 }),
  .ZN({ S12607 })
);
NAND3_X1 #() 
NAND3_X1_1541_ (
  .A1({ S12607 }),
  .A2({ S12067 }),
  .A3({ S11984 }),
  .ZN({ S12608 })
);
NAND3_X1 #() 
NAND3_X1_1542_ (
  .A1({ S12606 }),
  .A2({ S12608 }),
  .A3({ S25957[413] }),
  .ZN({ S12609 })
);
INV_X1 #() 
INV_X1_422_ (
  .A({ S12143 }),
  .ZN({ S12610 })
);
AOI21_X1 #() 
AOI21_X1_810_ (
  .A({ S25957[412] }),
  .B1({ S12019 }),
  .B2({ S12099 }),
  .ZN({ S12612 })
);
NAND2_X1 #() 
NAND2_X1_1311_ (
  .A1({ S12612 }),
  .A2({ S12610 }),
  .ZN({ S12613 })
);
NAND2_X1 #() 
NAND2_X1_1312_ (
  .A1({ S28 }),
  .A2({ S12011 }),
  .ZN({ S12614 })
);
NAND3_X1 #() 
NAND3_X1_1543_ (
  .A1({ S12090 }),
  .A2({ S25957[411] }),
  .A3({ S25957[409] }),
  .ZN({ S12615 })
);
NAND3_X1 #() 
NAND3_X1_1544_ (
  .A1({ S12615 }),
  .A2({ S25957[412] }),
  .A3({ S12614 }),
  .ZN({ S12616 })
);
NAND3_X1 #() 
NAND3_X1_1545_ (
  .A1({ S12613 }),
  .A2({ S12616 }),
  .A3({ S12034 }),
  .ZN({ S12617 })
);
NAND3_X1 #() 
NAND3_X1_1546_ (
  .A1({ S12609 }),
  .A2({ S12617 }),
  .A3({ S11981 }),
  .ZN({ S12618 })
);
NAND3_X1 #() 
NAND3_X1_1547_ (
  .A1({ S12604 }),
  .A2({ S25957[415] }),
  .A3({ S12618 }),
  .ZN({ S12619 })
);
NAND4_X1 #() 
NAND4_X1_188_ (
  .A1({ S12308 }),
  .A2({ S12090 }),
  .A3({ S12035 }),
  .A4({ S25957[411] }),
  .ZN({ S12620 })
);
AOI21_X1 #() 
AOI21_X1_811_ (
  .A({ S25957[412] }),
  .B1({ S12592 }),
  .B2({ S12620 }),
  .ZN({ S12621 })
);
NAND2_X1 #() 
NAND2_X1_1313_ (
  .A1({ S12046 }),
  .A2({ S25957[411] }),
  .ZN({ S12623 })
);
OAI211_X1 #() 
OAI211_X1_500_ (
  .A({ S12623 }),
  .B({ S25957[412] }),
  .C1({ S28 }),
  .C2({ S12183 }),
  .ZN({ S12624 })
);
NOR2_X1 #() 
NOR2_X1_306_ (
  .A1({ S12375 }),
  .A2({ S12624 }),
  .ZN({ S12625 })
);
NAND4_X1 #() 
NAND4_X1_189_ (
  .A1({ S12238 }),
  .A2({ S12005 }),
  .A3({ S12035 }),
  .A4({ S25957[411] }),
  .ZN({ S12626 })
);
NAND2_X1 #() 
NAND2_X1_1314_ (
  .A1({ S12626 }),
  .A2({ S12612 }),
  .ZN({ S12627 })
);
NAND2_X1 #() 
NAND2_X1_1315_ (
  .A1({ S12627 }),
  .A2({ S25957[413] }),
  .ZN({ S12628 })
);
NAND2_X1 #() 
NAND2_X1_1316_ (
  .A1({ S12615 }),
  .A2({ S25957[412] }),
  .ZN({ S12629 })
);
OAI21_X1 #() 
OAI21_X1_738_ (
  .A({ S12034 }),
  .B1({ S12300 }),
  .B2({ S12629 }),
  .ZN({ S12630 })
);
OAI22_X1 #() 
OAI22_X1_34_ (
  .A1({ S12625 }),
  .A2({ S12628 }),
  .B1({ S12630 }),
  .B2({ S12621 }),
  .ZN({ S12631 })
);
AND2_X1 #() 
AND2_X1_82_ (
  .A1({ S12411 }),
  .A2({ S11984 }),
  .ZN({ S12632 })
);
OAI211_X1 #() 
OAI211_X1_501_ (
  .A({ S25957[411] }),
  .B({ S12035 }),
  .C1({ S12012 }),
  .C2({ S11996 }),
  .ZN({ S12634 })
);
NAND2_X1 #() 
NAND2_X1_1317_ (
  .A1({ S12634 }),
  .A2({ S12398 }),
  .ZN({ S12635 })
);
AOI22_X1 #() 
AOI22_X1_176_ (
  .A1({ S12089 }),
  .A2({ S12632 }),
  .B1({ S12635 }),
  .B2({ S25957[412] }),
  .ZN({ S12636 })
);
OAI21_X1 #() 
OAI21_X1_739_ (
  .A({ S12025 }),
  .B1({ S25957[411] }),
  .B2({ S12000 }),
  .ZN({ S12637 })
);
NAND3_X1 #() 
NAND3_X1_1548_ (
  .A1({ S12376 }),
  .A2({ S12151 }),
  .A3({ S12637 }),
  .ZN({ S12638 })
);
AOI21_X1 #() 
AOI21_X1_812_ (
  .A({ S28 }),
  .B1({ S12124 }),
  .B2({ S12090 }),
  .ZN({ S12639 })
);
OAI211_X1 #() 
OAI211_X1_502_ (
  .A({ S25957[412] }),
  .B({ S12059 }),
  .C1({ S12534 }),
  .C2({ S25957[411] }),
  .ZN({ S12640 })
);
OAI211_X1 #() 
OAI211_X1_503_ (
  .A({ S12638 }),
  .B({ S12034 }),
  .C1({ S12639 }),
  .C2({ S12640 }),
  .ZN({ S12641 })
);
OAI211_X1 #() 
OAI211_X1_504_ (
  .A({ S12641 }),
  .B({ S25957[414] }),
  .C1({ S12636 }),
  .C2({ S12034 }),
  .ZN({ S12642 })
);
OAI211_X1 #() 
OAI211_X1_505_ (
  .A({ S12642 }),
  .B({ S9910 }),
  .C1({ S12631 }),
  .C2({ S25957[414] }),
  .ZN({ S12643 })
);
NAND3_X1 #() 
NAND3_X1_1549_ (
  .A1({ S12643 }),
  .A2({ S12619 }),
  .A3({ S25957[482] }),
  .ZN({ S12645 })
);
NAND2_X1 #() 
NAND2_X1_1318_ (
  .A1({ S12089 }),
  .A2({ S12632 }),
  .ZN({ S12646 })
);
NAND2_X1 #() 
NAND2_X1_1319_ (
  .A1({ S12635 }),
  .A2({ S25957[412] }),
  .ZN({ S12647 })
);
AOI21_X1 #() 
AOI21_X1_813_ (
  .A({ S12034 }),
  .B1({ S12646 }),
  .B2({ S12647 }),
  .ZN({ S12648 })
);
NOR2_X1 #() 
NOR2_X1_307_ (
  .A1({ S12640 }),
  .A2({ S12639 }),
  .ZN({ S12649 })
);
NAND2_X1 #() 
NAND2_X1_1320_ (
  .A1({ S12638 }),
  .A2({ S12034 }),
  .ZN({ S12650 })
);
NOR2_X1 #() 
NOR2_X1_308_ (
  .A1({ S12650 }),
  .A2({ S12649 }),
  .ZN({ S12651 })
);
OAI21_X1 #() 
OAI21_X1_740_ (
  .A({ S25957[414] }),
  .B1({ S12648 }),
  .B2({ S12651 }),
  .ZN({ S12652 })
);
NAND2_X1 #() 
NAND2_X1_1321_ (
  .A1({ S12631 }),
  .A2({ S11981 }),
  .ZN({ S12653 })
);
NAND3_X1 #() 
NAND3_X1_1550_ (
  .A1({ S12653 }),
  .A2({ S12652 }),
  .A3({ S9910 }),
  .ZN({ S12654 })
);
AOI22_X1 #() 
AOI22_X1_177_ (
  .A1({ S12595 }),
  .A2({ S12591 }),
  .B1({ S12602 }),
  .B2({ S12597 }),
  .ZN({ S12656 })
);
NAND2_X1 #() 
NAND2_X1_1322_ (
  .A1({ S12609 }),
  .A2({ S12617 }),
  .ZN({ S12657 })
);
NAND2_X1 #() 
NAND2_X1_1323_ (
  .A1({ S12657 }),
  .A2({ S11981 }),
  .ZN({ S12658 })
);
OAI211_X1 #() 
OAI211_X1_506_ (
  .A({ S12658 }),
  .B({ S25957[415] }),
  .C1({ S12656 }),
  .C2({ S11981 }),
  .ZN({ S12659 })
);
NAND3_X1 #() 
NAND3_X1_1551_ (
  .A1({ S12654 }),
  .A2({ S12588 }),
  .A3({ S12659 }),
  .ZN({ S12660 })
);
NAND3_X1 #() 
NAND3_X1_1552_ (
  .A1({ S12660 }),
  .A2({ S25957[450] }),
  .A3({ S12645 }),
  .ZN({ S12661 })
);
INV_X1 #() 
INV_X1_423_ (
  .A({ S25957[450] }),
  .ZN({ S12662 })
);
NAND3_X1 #() 
NAND3_X1_1553_ (
  .A1({ S12643 }),
  .A2({ S12619 }),
  .A3({ S12588 }),
  .ZN({ S12663 })
);
NAND3_X1 #() 
NAND3_X1_1554_ (
  .A1({ S12654 }),
  .A2({ S25957[482] }),
  .A3({ S12659 }),
  .ZN({ S12664 })
);
NAND3_X1 #() 
NAND3_X1_1555_ (
  .A1({ S12664 }),
  .A2({ S12662 }),
  .A3({ S12663 }),
  .ZN({ S12665 })
);
NAND3_X1 #() 
NAND3_X1_1556_ (
  .A1({ S12661 }),
  .A2({ S12665 }),
  .A3({ S25957[418] }),
  .ZN({ S12667 })
);
INV_X1 #() 
INV_X1_424_ (
  .A({ S25957[418] }),
  .ZN({ S12668 })
);
NAND3_X1 #() 
NAND3_X1_1557_ (
  .A1({ S12660 }),
  .A2({ S12662 }),
  .A3({ S12645 }),
  .ZN({ S12669 })
);
NAND3_X1 #() 
NAND3_X1_1558_ (
  .A1({ S12664 }),
  .A2({ S25957[450] }),
  .A3({ S12663 }),
  .ZN({ S12670 })
);
NAND3_X1 #() 
NAND3_X1_1559_ (
  .A1({ S12669 }),
  .A2({ S12670 }),
  .A3({ S12668 }),
  .ZN({ S12671 })
);
NAND3_X1 #() 
NAND3_X1_1560_ (
  .A1({ S12667 }),
  .A2({ S12671 }),
  .A3({ S11298 }),
  .ZN({ S12672 })
);
NAND3_X1 #() 
NAND3_X1_1561_ (
  .A1({ S12661 }),
  .A2({ S12665 }),
  .A3({ S12668 }),
  .ZN({ S12673 })
);
NAND3_X1 #() 
NAND3_X1_1562_ (
  .A1({ S12669 }),
  .A2({ S12670 }),
  .A3({ S25957[418] }),
  .ZN({ S12674 })
);
NAND3_X1 #() 
NAND3_X1_1563_ (
  .A1({ S12673 }),
  .A2({ S12674 }),
  .A3({ S25957[386] }),
  .ZN({ S12675 })
);
NAND2_X1 #() 
NAND2_X1_1324_ (
  .A1({ S12672 }),
  .A2({ S12675 }),
  .ZN({ S25957[258] })
);
OAI21_X1 #() 
OAI21_X1_741_ (
  .A({ S25957[400] }),
  .B1({ S11178 }),
  .B2({ S11177 }),
  .ZN({ S12677 })
);
INV_X1 #() 
INV_X1_425_ (
  .A({ S12677 }),
  .ZN({ S39 })
);
NAND3_X1 #() 
NAND3_X1_1564_ (
  .A1({ S8199 }),
  .A2({ S11081 }),
  .A3({ S8202 }),
  .ZN({ S40 })
);
XNOR2_X1 #() 
XNOR2_X1_45_ (
  .A({ S7025 }),
  .B({ S25957[767] }),
  .ZN({ S25957[639] })
);
XNOR2_X1 #() 
XNOR2_X1_46_ (
  .A({ S9899 }),
  .B({ S25957[639] }),
  .ZN({ S12678 })
);
NAND3_X1 #() 
NAND3_X1_1565_ (
  .A1({ S11279 }),
  .A2({ S25957[400] }),
  .A3({ S11280 }),
  .ZN({ S12679 })
);
AOI21_X1 #() 
AOI21_X1_814_ (
  .A({ S11179 }),
  .B1({ S8064 }),
  .B2({ S8067 }),
  .ZN({ S12680 })
);
NAND2_X1 #() 
NAND2_X1_1325_ (
  .A1({ S12680 }),
  .A2({ S12679 }),
  .ZN({ S12681 })
);
NAND3_X1 #() 
NAND3_X1_1566_ (
  .A1({ S7961 }),
  .A2({ S5128 }),
  .A3({ S7962 }),
  .ZN({ S12682 })
);
NAND3_X1 #() 
NAND3_X1_1567_ (
  .A1({ S7958 }),
  .A2({ S25957[532] }),
  .A3({ S7955 }),
  .ZN({ S12683 })
);
NAND2_X1 #() 
NAND2_X1_1326_ (
  .A1({ S12682 }),
  .A2({ S12683 }),
  .ZN({ S12685 })
);
AOI22_X1 #() 
AOI22_X1_178_ (
  .A1({ S8068 }),
  .A2({ S8069 }),
  .B1({ S12679 }),
  .B2({ S25957[401] }),
  .ZN({ S12686 })
);
NOR2_X1 #() 
NOR2_X1_309_ (
  .A1({ S12686 }),
  .A2({ S12685 }),
  .ZN({ S12687 })
);
NAND2_X1 #() 
NAND2_X1_1327_ (
  .A1({ S12687 }),
  .A2({ S12681 }),
  .ZN({ S12688 })
);
NAND3_X1 #() 
NAND3_X1_1568_ (
  .A1({ S8274 }),
  .A2({ S11081 }),
  .A3({ S8288 }),
  .ZN({ S12689 })
);
AOI21_X1 #() 
AOI21_X1_815_ (
  .A({ S25957[404] }),
  .B1({ S18 }),
  .B2({ S12689 }),
  .ZN({ S12690 })
);
NAND3_X1 #() 
NAND3_X1_1569_ (
  .A1({ S8064 }),
  .A2({ S8067 }),
  .A3({ S11081 }),
  .ZN({ S12691 })
);
INV_X1 #() 
INV_X1_426_ (
  .A({ S12691 }),
  .ZN({ S12692 })
);
OAI21_X1 #() 
OAI21_X1_742_ (
  .A({ S12690 }),
  .B1({ S12692 }),
  .B2({ S11179 }),
  .ZN({ S12693 })
);
NAND3_X1 #() 
NAND3_X1_1570_ (
  .A1({ S12688 }),
  .A2({ S12693 }),
  .A3({ S25957[405] }),
  .ZN({ S12694 })
);
NAND3_X1 #() 
NAND3_X1_1571_ (
  .A1({ S12677 }),
  .A2({ S40 }),
  .A3({ S25957[402] }),
  .ZN({ S12696 })
);
OAI21_X1 #() 
OAI21_X1_743_ (
  .A({ S11081 }),
  .B1({ S11178 }),
  .B2({ S11177 }),
  .ZN({ S12697 })
);
NAND3_X1 #() 
NAND3_X1_1572_ (
  .A1({ S8199 }),
  .A2({ S25957[400] }),
  .A3({ S8202 }),
  .ZN({ S12698 })
);
NAND3_X1 #() 
NAND3_X1_1573_ (
  .A1({ S12697 }),
  .A2({ S12698 }),
  .A3({ S11281 }),
  .ZN({ S12699 })
);
NAND3_X1 #() 
NAND3_X1_1574_ (
  .A1({ S25957[403] }),
  .A2({ S12696 }),
  .A3({ S12699 }),
  .ZN({ S12700 })
);
NAND4_X1 #() 
NAND4_X1_190_ (
  .A1({ S8274 }),
  .A2({ S8199 }),
  .A3({ S8288 }),
  .A4({ S8202 }),
  .ZN({ S12701 })
);
NAND3_X1 #() 
NAND3_X1_1575_ (
  .A1({ S8064 }),
  .A2({ S8067 }),
  .A3({ S12701 }),
  .ZN({ S12702 })
);
AOI21_X1 #() 
AOI21_X1_816_ (
  .A({ S25957[402] }),
  .B1({ S12697 }),
  .B2({ S12698 }),
  .ZN({ S12703 })
);
NAND2_X1 #() 
NAND2_X1_1328_ (
  .A1({ S12698 }),
  .A2({ S25957[402] }),
  .ZN({ S12704 })
);
INV_X1 #() 
INV_X1_427_ (
  .A({ S12704 }),
  .ZN({ S12705 })
);
OAI21_X1 #() 
OAI21_X1_744_ (
  .A({ S18 }),
  .B1({ S12703 }),
  .B2({ S12705 }),
  .ZN({ S12707 })
);
AOI21_X1 #() 
AOI21_X1_817_ (
  .A({ S25957[404] }),
  .B1({ S12707 }),
  .B2({ S12702 }),
  .ZN({ S12708 })
);
NAND4_X1 #() 
NAND4_X1_191_ (
  .A1({ S11279 }),
  .A2({ S8199 }),
  .A3({ S11280 }),
  .A4({ S8202 }),
  .ZN({ S12709 })
);
NAND3_X1 #() 
NAND3_X1_1576_ (
  .A1({ S8068 }),
  .A2({ S8069 }),
  .A3({ S12689 }),
  .ZN({ S12710 })
);
INV_X1 #() 
INV_X1_428_ (
  .A({ S12710 }),
  .ZN({ S12711 })
);
AOI21_X1 #() 
AOI21_X1_818_ (
  .A({ S12685 }),
  .B1({ S12711 }),
  .B2({ S12709 }),
  .ZN({ S12712 })
);
AOI21_X1 #() 
AOI21_X1_819_ (
  .A({ S12708 }),
  .B1({ S12700 }),
  .B2({ S12712 }),
  .ZN({ S12713 })
);
OAI21_X1 #() 
OAI21_X1_745_ (
  .A({ S12694 }),
  .B1({ S12713 }),
  .B2({ S25957[405] }),
  .ZN({ S12714 })
);
NAND3_X1 #() 
NAND3_X1_1577_ (
  .A1({ S12677 }),
  .A2({ S12679 }),
  .A3({ S12689 }),
  .ZN({ S12715 })
);
AOI21_X1 #() 
AOI21_X1_820_ (
  .A({ S12685 }),
  .B1({ S25957[403] }),
  .B2({ S12715 }),
  .ZN({ S12716 })
);
OAI21_X1 #() 
OAI21_X1_746_ (
  .A({ S12716 }),
  .B1({ S11179 }),
  .B2({ S12710 }),
  .ZN({ S12718 })
);
NAND3_X1 #() 
NAND3_X1_1578_ (
  .A1({ S8064 }),
  .A2({ S8067 }),
  .A3({ S11179 }),
  .ZN({ S12719 })
);
INV_X1 #() 
INV_X1_429_ (
  .A({ S12719 }),
  .ZN({ S12720 })
);
NAND2_X1 #() 
NAND2_X1_1329_ (
  .A1({ S12689 }),
  .A2({ S40 }),
  .ZN({ S12721 })
);
INV_X1 #() 
INV_X1_430_ (
  .A({ S12721 }),
  .ZN({ S12722 })
);
OAI21_X1 #() 
OAI21_X1_747_ (
  .A({ S12722 }),
  .B1({ S12720 }),
  .B2({ S12692 }),
  .ZN({ S12723 })
);
AOI21_X1 #() 
AOI21_X1_821_ (
  .A({ S11081 }),
  .B1({ S11279 }),
  .B2({ S11280 }),
  .ZN({ S12724 })
);
NAND2_X1 #() 
NAND2_X1_1330_ (
  .A1({ S12724 }),
  .A2({ S25957[401] }),
  .ZN({ S12725 })
);
AOI21_X1 #() 
AOI21_X1_822_ (
  .A({ S25957[400] }),
  .B1({ S8274 }),
  .B2({ S8288 }),
  .ZN({ S12726 })
);
NAND2_X1 #() 
NAND2_X1_1331_ (
  .A1({ S12726 }),
  .A2({ S11179 }),
  .ZN({ S12727 })
);
NAND2_X1 #() 
NAND2_X1_1332_ (
  .A1({ S12725 }),
  .A2({ S12727 }),
  .ZN({ S12729 })
);
INV_X1 #() 
INV_X1_431_ (
  .A({ S12729 }),
  .ZN({ S12730 })
);
OAI21_X1 #() 
OAI21_X1_748_ (
  .A({ S12723 }),
  .B1({ S25957[403] }),
  .B2({ S12730 }),
  .ZN({ S12731 })
);
OAI211_X1 #() 
OAI211_X1_507_ (
  .A({ S25957[405] }),
  .B({ S12718 }),
  .C1({ S12731 }),
  .C2({ S25957[404] }),
  .ZN({ S12732 })
);
NAND2_X1 #() 
NAND2_X1_1333_ (
  .A1({ S40 }),
  .A2({ S11281 }),
  .ZN({ S12733 })
);
NAND2_X1 #() 
NAND2_X1_1334_ (
  .A1({ S12727 }),
  .A2({ S12733 }),
  .ZN({ S12734 })
);
INV_X1 #() 
INV_X1_432_ (
  .A({ S12698 }),
  .ZN({ S12735 })
);
NAND2_X1 #() 
NAND2_X1_1335_ (
  .A1({ S25957[403] }),
  .A2({ S12735 }),
  .ZN({ S12736 })
);
AOI21_X1 #() 
AOI21_X1_823_ (
  .A({ S25957[404] }),
  .B1({ S12736 }),
  .B2({ S12734 }),
  .ZN({ S12737 })
);
AOI21_X1 #() 
AOI21_X1_824_ (
  .A({ S25957[400] }),
  .B1({ S8199 }),
  .B2({ S8202 }),
  .ZN({ S12738 })
);
NAND3_X1 #() 
NAND3_X1_1579_ (
  .A1({ S25957[403] }),
  .A2({ S12677 }),
  .A3({ S12709 }),
  .ZN({ S12740 })
);
OAI211_X1 #() 
OAI211_X1_508_ (
  .A({ S12740 }),
  .B({ S25957[404] }),
  .C1({ S25957[403] }),
  .C2({ S12738 }),
  .ZN({ S12741 })
);
NAND2_X1 #() 
NAND2_X1_1336_ (
  .A1({ S12741 }),
  .A2({ S10807 }),
  .ZN({ S12742 })
);
OAI21_X1 #() 
OAI21_X1_749_ (
  .A({ S12732 }),
  .B1({ S12737 }),
  .B2({ S12742 }),
  .ZN({ S12743 })
);
MUX2_X1 #() 
MUX2_X1_4_ (
  .A({ S12714 }),
  .B({ S12743 }),
  .S({ S25957[406] }),
  .Z({ S12744 })
);
NAND2_X1 #() 
NAND2_X1_1337_ (
  .A1({ S12744 }),
  .A2({ S25957[407] }),
  .ZN({ S12745 })
);
NOR2_X1 #() 
NOR2_X1_310_ (
  .A1({ S12729 }),
  .A2({ S18 }),
  .ZN({ S12746 })
);
OAI21_X1 #() 
OAI21_X1_750_ (
  .A({ S11081 }),
  .B1({ S11281 }),
  .B2({ S25957[401] }),
  .ZN({ S12747 })
);
NAND2_X1 #() 
NAND2_X1_1338_ (
  .A1({ S18 }),
  .A2({ S12747 }),
  .ZN({ S12748 })
);
NAND2_X1 #() 
NAND2_X1_1339_ (
  .A1({ S12748 }),
  .A2({ S25957[404] }),
  .ZN({ S12749 })
);
OAI211_X1 #() 
OAI211_X1_509_ (
  .A({ S11279 }),
  .B({ S11280 }),
  .C1({ S11178 }),
  .C2({ S11177 }),
  .ZN({ S12751 })
);
NAND2_X1 #() 
NAND2_X1_1340_ (
  .A1({ S12724 }),
  .A2({ S11179 }),
  .ZN({ S12752 })
);
NAND2_X1 #() 
NAND2_X1_1341_ (
  .A1({ S12752 }),
  .A2({ S12751 }),
  .ZN({ S12753 })
);
NAND2_X1 #() 
NAND2_X1_1342_ (
  .A1({ S12753 }),
  .A2({ S25957[403] }),
  .ZN({ S12754 })
);
NAND2_X1 #() 
NAND2_X1_1343_ (
  .A1({ S12677 }),
  .A2({ S25957[402] }),
  .ZN({ S12755 })
);
NAND3_X1 #() 
NAND3_X1_1580_ (
  .A1({ S12755 }),
  .A2({ S8068 }),
  .A3({ S8069 }),
  .ZN({ S12756 })
);
NAND3_X1 #() 
NAND3_X1_1581_ (
  .A1({ S12754 }),
  .A2({ S12685 }),
  .A3({ S12756 }),
  .ZN({ S12757 })
);
OAI21_X1 #() 
OAI21_X1_751_ (
  .A({ S12757 }),
  .B1({ S12746 }),
  .B2({ S12749 }),
  .ZN({ S12758 })
);
AOI22_X1 #() 
AOI22_X1_179_ (
  .A1({ S12699 }),
  .A2({ S12755 }),
  .B1({ S8069 }),
  .B2({ S8068 }),
  .ZN({ S12759 })
);
INV_X1 #() 
INV_X1_433_ (
  .A({ S12759 }),
  .ZN({ S12760 })
);
NAND3_X1 #() 
NAND3_X1_1582_ (
  .A1({ S8274 }),
  .A2({ S25957[400] }),
  .A3({ S8288 }),
  .ZN({ S12762 })
);
NAND3_X1 #() 
NAND3_X1_1583_ (
  .A1({ S18 }),
  .A2({ S12762 }),
  .A3({ S12696 }),
  .ZN({ S12763 })
);
NAND3_X1 #() 
NAND3_X1_1584_ (
  .A1({ S12760 }),
  .A2({ S25957[404] }),
  .A3({ S12763 }),
  .ZN({ S12764 })
);
OAI211_X1 #() 
OAI211_X1_510_ (
  .A({ S8274 }),
  .B({ S8288 }),
  .C1({ S11178 }),
  .C2({ S11177 }),
  .ZN({ S12765 })
);
NAND4_X1 #() 
NAND4_X1_192_ (
  .A1({ S8064 }),
  .A2({ S8067 }),
  .A3({ S12765 }),
  .A4({ S12679 }),
  .ZN({ S12766 })
);
NAND3_X1 #() 
NAND3_X1_1585_ (
  .A1({ S12765 }),
  .A2({ S12709 }),
  .A3({ S25957[400] }),
  .ZN({ S12767 })
);
AOI21_X1 #() 
AOI21_X1_825_ (
  .A({ S25957[404] }),
  .B1({ S18 }),
  .B2({ S12767 }),
  .ZN({ S12768 })
);
AOI21_X1 #() 
AOI21_X1_826_ (
  .A({ S25957[405] }),
  .B1({ S12768 }),
  .B2({ S12766 }),
  .ZN({ S12769 })
);
AOI22_X1 #() 
AOI22_X1_180_ (
  .A1({ S12758 }),
  .A2({ S25957[405] }),
  .B1({ S12764 }),
  .B2({ S12769 }),
  .ZN({ S12770 })
);
NAND3_X1 #() 
NAND3_X1_1586_ (
  .A1({ S11279 }),
  .A2({ S11081 }),
  .A3({ S11280 }),
  .ZN({ S12771 })
);
NOR2_X1 #() 
NOR2_X1_311_ (
  .A1({ S12771 }),
  .A2({ S11179 }),
  .ZN({ S12773 })
);
NAND3_X1 #() 
NAND3_X1_1587_ (
  .A1({ S25957[402] }),
  .A2({ S25957[401] }),
  .A3({ S25957[400] }),
  .ZN({ S12774 })
);
NAND2_X1 #() 
NAND2_X1_1344_ (
  .A1({ S12679 }),
  .A2({ S11179 }),
  .ZN({ S12775 })
);
NAND3_X1 #() 
NAND3_X1_1588_ (
  .A1({ S12774 }),
  .A2({ S12775 }),
  .A3({ S12689 }),
  .ZN({ S12776 })
);
AOI21_X1 #() 
AOI21_X1_827_ (
  .A({ S12685 }),
  .B1({ S12776 }),
  .B2({ S18 }),
  .ZN({ S12777 })
);
OAI21_X1 #() 
OAI21_X1_752_ (
  .A({ S12777 }),
  .B1({ S18 }),
  .B2({ S12773 }),
  .ZN({ S12778 })
);
NAND3_X1 #() 
NAND3_X1_1589_ (
  .A1({ S12697 }),
  .A2({ S12698 }),
  .A3({ S25957[402] }),
  .ZN({ S12779 })
);
NOR2_X1 #() 
NOR2_X1_312_ (
  .A1({ S25957[403] }),
  .A2({ S12779 }),
  .ZN({ S12780 })
);
OAI21_X1 #() 
OAI21_X1_753_ (
  .A({ S12685 }),
  .B1({ S18 }),
  .B2({ S12755 }),
  .ZN({ S12781 })
);
OAI21_X1 #() 
OAI21_X1_754_ (
  .A({ S12778 }),
  .B1({ S12780 }),
  .B2({ S12781 }),
  .ZN({ S12782 })
);
NAND4_X1 #() 
NAND4_X1_193_ (
  .A1({ S8064 }),
  .A2({ S8067 }),
  .A3({ S12679 }),
  .A4({ S12701 }),
  .ZN({ S12783 })
);
OAI21_X1 #() 
OAI21_X1_755_ (
  .A({ S12783 }),
  .B1({ S25957[403] }),
  .B2({ S11081 }),
  .ZN({ S12784 })
);
NOR2_X1 #() 
NOR2_X1_313_ (
  .A1({ S12784 }),
  .A2({ S12685 }),
  .ZN({ S12785 })
);
NAND2_X1 #() 
NAND2_X1_1345_ (
  .A1({ S12701 }),
  .A2({ S12689 }),
  .ZN({ S12786 })
);
NAND3_X1 #() 
NAND3_X1_1590_ (
  .A1({ S8068 }),
  .A2({ S8069 }),
  .A3({ S12751 }),
  .ZN({ S12787 })
);
NAND4_X1 #() 
NAND4_X1_194_ (
  .A1({ S8064 }),
  .A2({ S8067 }),
  .A3({ S12765 }),
  .A4({ S12698 }),
  .ZN({ S12788 })
);
OAI21_X1 #() 
OAI21_X1_756_ (
  .A({ S12788 }),
  .B1({ S12787 }),
  .B2({ S12786 }),
  .ZN({ S12789 })
);
AOI21_X1 #() 
AOI21_X1_828_ (
  .A({ S12785 }),
  .B1({ S12685 }),
  .B2({ S12789 }),
  .ZN({ S12790 })
);
AOI21_X1 #() 
AOI21_X1_829_ (
  .A({ S25957[406] }),
  .B1({ S12790 }),
  .B2({ S25957[405] }),
  .ZN({ S12791 })
);
OAI21_X1 #() 
OAI21_X1_757_ (
  .A({ S12791 }),
  .B1({ S25957[405] }),
  .B2({ S12782 }),
  .ZN({ S12792 })
);
OAI21_X1 #() 
OAI21_X1_758_ (
  .A({ S12792 }),
  .B1({ S12770 }),
  .B2({ S7784 }),
  .ZN({ S12794 })
);
NAND2_X1 #() 
NAND2_X1_1346_ (
  .A1({ S12794 }),
  .A2({ S7707 }),
  .ZN({ S12795 })
);
NAND2_X1 #() 
NAND2_X1_1347_ (
  .A1({ S12745 }),
  .A2({ S12795 }),
  .ZN({ S12796 })
);
NAND2_X1 #() 
NAND2_X1_1348_ (
  .A1({ S12796 }),
  .A2({ S12678 }),
  .ZN({ S12797 })
);
INV_X1 #() 
INV_X1_434_ (
  .A({ S12678 }),
  .ZN({ S25957[511] })
);
NAND3_X1 #() 
NAND3_X1_1591_ (
  .A1({ S12745 }),
  .A2({ S25957[511] }),
  .A3({ S12795 }),
  .ZN({ S12798 })
);
NAND3_X1 #() 
NAND3_X1_1592_ (
  .A1({ S12797 }),
  .A2({ S25957[575] }),
  .A3({ S12798 }),
  .ZN({ S12799 })
);
NAND2_X1 #() 
NAND2_X1_1349_ (
  .A1({ S12797 }),
  .A2({ S12798 }),
  .ZN({ S25957[383] })
);
NAND2_X1 #() 
NAND2_X1_1350_ (
  .A1({ S25957[383] }),
  .A2({ S9903 }),
  .ZN({ S12800 })
);
NAND3_X1 #() 
NAND3_X1_1593_ (
  .A1({ S12800 }),
  .A2({ S9910 }),
  .A3({ S12799 }),
  .ZN({ S12801 })
);
NAND2_X1 #() 
NAND2_X1_1351_ (
  .A1({ S12800 }),
  .A2({ S12799 }),
  .ZN({ S25957[319] })
);
NAND2_X1 #() 
NAND2_X1_1352_ (
  .A1({ S25957[319] }),
  .A2({ S25957[415] }),
  .ZN({ S12803 })
);
AND2_X1 #() 
AND2_X1_83_ (
  .A1({ S12803 }),
  .A2({ S12801 }),
  .ZN({ S25957[287] })
);
NAND2_X1 #() 
NAND2_X1_1353_ (
  .A1({ S12697 }),
  .A2({ S12679 }),
  .ZN({ S12804 })
);
INV_X1 #() 
INV_X1_435_ (
  .A({ S12804 }),
  .ZN({ S12805 })
);
NAND4_X1 #() 
NAND4_X1_195_ (
  .A1({ S12755 }),
  .A2({ S12762 }),
  .A3({ S8068 }),
  .A4({ S8069 }),
  .ZN({ S12806 })
);
OAI211_X1 #() 
OAI211_X1_511_ (
  .A({ S12806 }),
  .B({ S25957[404] }),
  .C1({ S18 }),
  .C2({ S12805 }),
  .ZN({ S12807 })
);
OAI211_X1 #() 
OAI211_X1_512_ (
  .A({ S12685 }),
  .B({ S12804 }),
  .C1({ S25957[403] }),
  .C2({ S25957[401] }),
  .ZN({ S12808 })
);
NAND3_X1 #() 
NAND3_X1_1594_ (
  .A1({ S12807 }),
  .A2({ S25957[405] }),
  .A3({ S12808 }),
  .ZN({ S12809 })
);
NAND2_X1 #() 
NAND2_X1_1354_ (
  .A1({ S12704 }),
  .A2({ S12762 }),
  .ZN({ S12810 })
);
NAND2_X1 #() 
NAND2_X1_1355_ (
  .A1({ S12810 }),
  .A2({ S25957[403] }),
  .ZN({ S12812 })
);
NAND2_X1 #() 
NAND2_X1_1356_ (
  .A1({ S12812 }),
  .A2({ S12685 }),
  .ZN({ S12813 })
);
AOI21_X1 #() 
AOI21_X1_830_ (
  .A({ S12813 }),
  .B1({ S12696 }),
  .B2({ S18 }),
  .ZN({ S12814 })
);
NAND2_X1 #() 
NAND2_X1_1357_ (
  .A1({ S12701 }),
  .A2({ S11081 }),
  .ZN({ S12815 })
);
INV_X1 #() 
INV_X1_436_ (
  .A({ S12815 }),
  .ZN({ S12816 })
);
OAI21_X1 #() 
OAI21_X1_759_ (
  .A({ S25957[404] }),
  .B1({ S18 }),
  .B2({ S12765 }),
  .ZN({ S12817 })
);
AOI21_X1 #() 
AOI21_X1_831_ (
  .A({ S12817 }),
  .B1({ S12816 }),
  .B2({ S18 }),
  .ZN({ S12818 })
);
OAI21_X1 #() 
OAI21_X1_760_ (
  .A({ S10807 }),
  .B1({ S12814 }),
  .B2({ S12818 }),
  .ZN({ S12819 })
);
NAND3_X1 #() 
NAND3_X1_1595_ (
  .A1({ S12819 }),
  .A2({ S25957[406] }),
  .A3({ S12809 }),
  .ZN({ S12820 })
);
INV_X1 #() 
INV_X1_437_ (
  .A({ S12751 }),
  .ZN({ S12821 })
);
NAND2_X1 #() 
NAND2_X1_1358_ (
  .A1({ S12753 }),
  .A2({ S18 }),
  .ZN({ S12823 })
);
OAI21_X1 #() 
OAI21_X1_761_ (
  .A({ S12823 }),
  .B1({ S12821 }),
  .B2({ S12702 }),
  .ZN({ S12824 })
);
NOR2_X1 #() 
NOR2_X1_314_ (
  .A1({ S25957[403] }),
  .A2({ S12724 }),
  .ZN({ S12825 })
);
OAI21_X1 #() 
OAI21_X1_762_ (
  .A({ S12677 }),
  .B1({ S40 }),
  .B2({ S11281 }),
  .ZN({ S12826 })
);
NOR2_X1 #() 
NOR2_X1_315_ (
  .A1({ S18 }),
  .A2({ S12826 }),
  .ZN({ S12827 })
);
OAI21_X1 #() 
OAI21_X1_763_ (
  .A({ S25957[404] }),
  .B1({ S12825 }),
  .B2({ S12827 }),
  .ZN({ S12828 })
);
OAI211_X1 #() 
OAI211_X1_513_ (
  .A({ S12828 }),
  .B({ S25957[405] }),
  .C1({ S12824 }),
  .C2({ S25957[404] }),
  .ZN({ S12829 })
);
OAI211_X1 #() 
OAI211_X1_514_ (
  .A({ S12701 }),
  .B({ S12762 }),
  .C1({ S12771 }),
  .C2({ S11179 }),
  .ZN({ S12830 })
);
NAND2_X1 #() 
NAND2_X1_1359_ (
  .A1({ S12830 }),
  .A2({ S25957[403] }),
  .ZN({ S12831 })
);
NAND2_X1 #() 
NAND2_X1_1360_ (
  .A1({ S18 }),
  .A2({ S12752 }),
  .ZN({ S12832 })
);
NAND3_X1 #() 
NAND3_X1_1596_ (
  .A1({ S12754 }),
  .A2({ S25957[404] }),
  .A3({ S12832 }),
  .ZN({ S12834 })
);
OAI211_X1 #() 
OAI211_X1_515_ (
  .A({ S12834 }),
  .B({ S10807 }),
  .C1({ S25957[404] }),
  .C2({ S12831 }),
  .ZN({ S12835 })
);
NAND3_X1 #() 
NAND3_X1_1597_ (
  .A1({ S12829 }),
  .A2({ S12835 }),
  .A3({ S7784 }),
  .ZN({ S12836 })
);
AOI21_X1 #() 
AOI21_X1_832_ (
  .A({ S25957[407] }),
  .B1({ S12820 }),
  .B2({ S12836 }),
  .ZN({ S12837 })
);
NAND3_X1 #() 
NAND3_X1_1598_ (
  .A1({ S12821 }),
  .A2({ S8064 }),
  .A3({ S8067 }),
  .ZN({ S12838 })
);
NOR2_X1 #() 
NOR2_X1_316_ (
  .A1({ S12689 }),
  .A2({ S11179 }),
  .ZN({ S12839 })
);
NAND3_X1 #() 
NAND3_X1_1599_ (
  .A1({ S12839 }),
  .A2({ S8068 }),
  .A3({ S8069 }),
  .ZN({ S12840 })
);
NAND2_X1 #() 
NAND2_X1_1361_ (
  .A1({ S12840 }),
  .A2({ S12838 }),
  .ZN({ S12841 })
);
OAI21_X1 #() 
OAI21_X1_764_ (
  .A({ S25957[404] }),
  .B1({ S12841 }),
  .B2({ S12780 }),
  .ZN({ S12842 })
);
OAI21_X1 #() 
OAI21_X1_765_ (
  .A({ S40 }),
  .B1({ S12679 }),
  .B2({ S11179 }),
  .ZN({ S12843 })
);
NAND2_X1 #() 
NAND2_X1_1362_ (
  .A1({ S18 }),
  .A2({ S12843 }),
  .ZN({ S12845 })
);
NAND2_X1 #() 
NAND2_X1_1363_ (
  .A1({ S12697 }),
  .A2({ S11281 }),
  .ZN({ S12846 })
);
NAND2_X1 #() 
NAND2_X1_1364_ (
  .A1({ S12846 }),
  .A2({ S12751 }),
  .ZN({ S12847 })
);
NAND2_X1 #() 
NAND2_X1_1365_ (
  .A1({ S12847 }),
  .A2({ S25957[403] }),
  .ZN({ S12848 })
);
NAND3_X1 #() 
NAND3_X1_1600_ (
  .A1({ S12848 }),
  .A2({ S12685 }),
  .A3({ S12845 }),
  .ZN({ S12849 })
);
NAND3_X1 #() 
NAND3_X1_1601_ (
  .A1({ S12842 }),
  .A2({ S25957[405] }),
  .A3({ S12849 }),
  .ZN({ S12850 })
);
NAND2_X1 #() 
NAND2_X1_1366_ (
  .A1({ S12698 }),
  .A2({ S11281 }),
  .ZN({ S12851 })
);
OAI21_X1 #() 
OAI21_X1_766_ (
  .A({ S12687 }),
  .B1({ S25957[403] }),
  .B2({ S12851 }),
  .ZN({ S12852 })
);
NAND3_X1 #() 
NAND3_X1_1602_ (
  .A1({ S12677 }),
  .A2({ S40 }),
  .A3({ S11281 }),
  .ZN({ S12853 })
);
AOI21_X1 #() 
AOI21_X1_833_ (
  .A({ S25957[403] }),
  .B1({ S12679 }),
  .B2({ S12853 }),
  .ZN({ S12854 })
);
AOI21_X1 #() 
AOI21_X1_834_ (
  .A({ S11081 }),
  .B1({ S8274 }),
  .B2({ S8288 }),
  .ZN({ S12856 })
);
NOR3_X1 #() 
NOR3_X1_43_ (
  .A1({ S18 }),
  .A2({ S12856 }),
  .A3({ S12721 }),
  .ZN({ S12857 })
);
OAI21_X1 #() 
OAI21_X1_767_ (
  .A({ S12685 }),
  .B1({ S12854 }),
  .B2({ S12857 }),
  .ZN({ S12858 })
);
NAND3_X1 #() 
NAND3_X1_1603_ (
  .A1({ S12858 }),
  .A2({ S12852 }),
  .A3({ S10807 }),
  .ZN({ S12859 })
);
NAND3_X1 #() 
NAND3_X1_1604_ (
  .A1({ S12859 }),
  .A2({ S7784 }),
  .A3({ S12850 }),
  .ZN({ S12860 })
);
NAND2_X1 #() 
NAND2_X1_1367_ (
  .A1({ S40 }),
  .A2({ S25957[402] }),
  .ZN({ S12861 })
);
NAND4_X1 #() 
NAND4_X1_196_ (
  .A1({ S12704 }),
  .A2({ S12733 }),
  .A3({ S8064 }),
  .A4({ S8067 }),
  .ZN({ S12862 })
);
OAI21_X1 #() 
OAI21_X1_768_ (
  .A({ S12862 }),
  .B1({ S25957[403] }),
  .B2({ S12861 }),
  .ZN({ S12863 })
);
INV_X1 #() 
INV_X1_438_ (
  .A({ S12740 }),
  .ZN({ S12864 })
);
OAI21_X1 #() 
OAI21_X1_769_ (
  .A({ S12685 }),
  .B1({ S12864 }),
  .B2({ S12680 }),
  .ZN({ S12865 })
);
OAI211_X1 #() 
OAI211_X1_516_ (
  .A({ S12865 }),
  .B({ S25957[405] }),
  .C1({ S12685 }),
  .C2({ S12863 }),
  .ZN({ S12867 })
);
INV_X1 #() 
INV_X1_439_ (
  .A({ S12812 }),
  .ZN({ S12868 })
);
NOR3_X1 #() 
NOR3_X1_44_ (
  .A1({ S12868 }),
  .A2({ S12854 }),
  .A3({ S12685 }),
  .ZN({ S12869 })
);
INV_X1 #() 
INV_X1_440_ (
  .A({ S12702 }),
  .ZN({ S12870 })
);
NAND2_X1 #() 
NAND2_X1_1368_ (
  .A1({ S18 }),
  .A2({ S12767 }),
  .ZN({ S12871 })
);
NAND2_X1 #() 
NAND2_X1_1369_ (
  .A1({ S12871 }),
  .A2({ S12685 }),
  .ZN({ S12872 })
);
AOI21_X1 #() 
AOI21_X1_835_ (
  .A({ S12872 }),
  .B1({ S12722 }),
  .B2({ S12870 }),
  .ZN({ S12873 })
);
OAI21_X1 #() 
OAI21_X1_770_ (
  .A({ S10807 }),
  .B1({ S12873 }),
  .B2({ S12869 }),
  .ZN({ S12874 })
);
NAND3_X1 #() 
NAND3_X1_1605_ (
  .A1({ S12874 }),
  .A2({ S25957[406] }),
  .A3({ S12867 }),
  .ZN({ S12875 })
);
AOI21_X1 #() 
AOI21_X1_836_ (
  .A({ S7707 }),
  .B1({ S12875 }),
  .B2({ S12860 }),
  .ZN({ S12876 })
);
NOR2_X1 #() 
NOR2_X1_317_ (
  .A1({ S12876 }),
  .A2({ S12837 }),
  .ZN({ S12877 })
);
NAND2_X1 #() 
NAND2_X1_1370_ (
  .A1({ S12877 }),
  .A2({ S25957[510] }),
  .ZN({ S12878 })
);
OAI211_X1 #() 
OAI211_X1_517_ (
  .A({ S9989 }),
  .B({ S9992 }),
  .C1({ S12876 }),
  .C2({ S12837 }),
  .ZN({ S12879 })
);
NAND2_X1 #() 
NAND2_X1_1371_ (
  .A1({ S12878 }),
  .A2({ S12879 }),
  .ZN({ S12880 })
);
NOR2_X1 #() 
NOR2_X1_318_ (
  .A1({ S12880 }),
  .A2({ S9998 }),
  .ZN({ S12881 })
);
AOI21_X1 #() 
AOI21_X1_837_ (
  .A({ S25957[574] }),
  .B1({ S12878 }),
  .B2({ S12879 }),
  .ZN({ S12882 })
);
OAI21_X1 #() 
OAI21_X1_771_ (
  .A({ S25957[414] }),
  .B1({ S12881 }),
  .B2({ S12882 }),
  .ZN({ S12883 })
);
INV_X1 #() 
INV_X1_441_ (
  .A({ S12880 }),
  .ZN({ S25957[382] })
);
NAND2_X1 #() 
NAND2_X1_1372_ (
  .A1({ S25957[382] }),
  .A2({ S25957[574] }),
  .ZN({ S12884 })
);
INV_X1 #() 
INV_X1_442_ (
  .A({ S12882 }),
  .ZN({ S12885 })
);
NAND3_X1 #() 
NAND3_X1_1606_ (
  .A1({ S12884 }),
  .A2({ S11981 }),
  .A3({ S12885 }),
  .ZN({ S12887 })
);
NAND2_X1 #() 
NAND2_X1_1373_ (
  .A1({ S12887 }),
  .A2({ S12883 }),
  .ZN({ S25957[286] })
);
NAND2_X1 #() 
NAND2_X1_1374_ (
  .A1({ S7197 }),
  .A2({ S7200 }),
  .ZN({ S25957[573] })
);
INV_X1 #() 
INV_X1_443_ (
  .A({ S25957[573] }),
  .ZN({ S12888 })
);
NOR2_X1 #() 
NOR2_X1_319_ (
  .A1({ S12762 }),
  .A2({ S11179 }),
  .ZN({ S12889 })
);
NOR2_X1 #() 
NOR2_X1_320_ (
  .A1({ S25957[403] }),
  .A2({ S12889 }),
  .ZN({ S12890 })
);
NAND3_X1 #() 
NAND3_X1_1607_ (
  .A1({ S11179 }),
  .A2({ S11281 }),
  .A3({ S11081 }),
  .ZN({ S12891 })
);
AOI21_X1 #() 
AOI21_X1_838_ (
  .A({ S18 }),
  .B1({ S12891 }),
  .B2({ S12696 }),
  .ZN({ S12892 })
);
NOR3_X1 #() 
NOR3_X1_45_ (
  .A1({ S12892 }),
  .A2({ S12890 }),
  .A3({ S25957[404] }),
  .ZN({ S12893 })
);
OAI21_X1 #() 
OAI21_X1_772_ (
  .A({ S18 }),
  .B1({ S12726 }),
  .B2({ S12735 }),
  .ZN({ S12894 })
);
OAI211_X1 #() 
OAI211_X1_518_ (
  .A({ S12894 }),
  .B({ S25957[404] }),
  .C1({ S18 }),
  .C2({ S12767 }),
  .ZN({ S12896 })
);
NAND4_X1 #() 
NAND4_X1_197_ (
  .A1({ S8068 }),
  .A2({ S8069 }),
  .A3({ S12701 }),
  .A4({ S12697 }),
  .ZN({ S12897 })
);
NAND3_X1 #() 
NAND3_X1_1608_ (
  .A1({ S12897 }),
  .A2({ S12685 }),
  .A3({ S12719 }),
  .ZN({ S12898 })
);
NAND3_X1 #() 
NAND3_X1_1609_ (
  .A1({ S12896 }),
  .A2({ S25957[405] }),
  .A3({ S12898 }),
  .ZN({ S12899 })
);
NAND2_X1 #() 
NAND2_X1_1375_ (
  .A1({ S25957[403] }),
  .A2({ S12703 }),
  .ZN({ S12900 })
);
NAND2_X1 #() 
NAND2_X1_1376_ (
  .A1({ S12709 }),
  .A2({ S40 }),
  .ZN({ S12901 })
);
NAND3_X1 #() 
NAND3_X1_1610_ (
  .A1({ S12901 }),
  .A2({ S8068 }),
  .A3({ S8069 }),
  .ZN({ S12902 })
);
NAND2_X1 #() 
NAND2_X1_1377_ (
  .A1({ S12900 }),
  .A2({ S12902 }),
  .ZN({ S12903 })
);
NAND2_X1 #() 
NAND2_X1_1378_ (
  .A1({ S12903 }),
  .A2({ S25957[404] }),
  .ZN({ S12904 })
);
NAND2_X1 #() 
NAND2_X1_1379_ (
  .A1({ S12904 }),
  .A2({ S10807 }),
  .ZN({ S12905 })
);
OAI211_X1 #() 
OAI211_X1_519_ (
  .A({ S12899 }),
  .B({ S7784 }),
  .C1({ S12905 }),
  .C2({ S12893 }),
  .ZN({ S12907 })
);
NAND2_X1 #() 
NAND2_X1_1380_ (
  .A1({ S12709 }),
  .A2({ S12679 }),
  .ZN({ S12908 })
);
NAND2_X1 #() 
NAND2_X1_1381_ (
  .A1({ S18 }),
  .A2({ S12908 }),
  .ZN({ S12909 })
);
NAND2_X1 #() 
NAND2_X1_1382_ (
  .A1({ S25957[403] }),
  .A2({ S12846 }),
  .ZN({ S12910 })
);
NAND3_X1 #() 
NAND3_X1_1611_ (
  .A1({ S12909 }),
  .A2({ S12910 }),
  .A3({ S25957[404] }),
  .ZN({ S12911 })
);
OAI21_X1 #() 
OAI21_X1_773_ (
  .A({ S12911 }),
  .B1({ S12813 }),
  .B2({ S12780 }),
  .ZN({ S12912 })
);
INV_X1 #() 
INV_X1_444_ (
  .A({ S12775 }),
  .ZN({ S12913 })
);
NAND3_X1 #() 
NAND3_X1_1612_ (
  .A1({ S12679 }),
  .A2({ S12689 }),
  .A3({ S25957[401] }),
  .ZN({ S12914 })
);
NAND2_X1 #() 
NAND2_X1_1383_ (
  .A1({ S25957[403] }),
  .A2({ S12914 }),
  .ZN({ S12915 })
);
OAI211_X1 #() 
OAI211_X1_520_ (
  .A({ S12915 }),
  .B({ S12685 }),
  .C1({ S25957[403] }),
  .C2({ S12913 }),
  .ZN({ S12916 })
);
NAND2_X1 #() 
NAND2_X1_1384_ (
  .A1({ S12697 }),
  .A2({ S25957[402] }),
  .ZN({ S12918 })
);
NAND3_X1 #() 
NAND3_X1_1613_ (
  .A1({ S18 }),
  .A2({ S12918 }),
  .A3({ S12698 }),
  .ZN({ S12919 })
);
OAI211_X1 #() 
OAI211_X1_521_ (
  .A({ S12919 }),
  .B({ S25957[404] }),
  .C1({ S18 }),
  .C2({ S12816 }),
  .ZN({ S12920 })
);
NAND3_X1 #() 
NAND3_X1_1614_ (
  .A1({ S12920 }),
  .A2({ S12916 }),
  .A3({ S25957[405] }),
  .ZN({ S12921 })
);
OAI211_X1 #() 
OAI211_X1_522_ (
  .A({ S12921 }),
  .B({ S25957[406] }),
  .C1({ S12912 }),
  .C2({ S25957[405] }),
  .ZN({ S12922 })
);
NAND3_X1 #() 
NAND3_X1_1615_ (
  .A1({ S12907 }),
  .A2({ S12922 }),
  .A3({ S25957[407] }),
  .ZN({ S12923 })
);
NAND2_X1 #() 
NAND2_X1_1385_ (
  .A1({ S18 }),
  .A2({ S12826 }),
  .ZN({ S12924 })
);
NAND2_X1 #() 
NAND2_X1_1386_ (
  .A1({ S12779 }),
  .A2({ S12752 }),
  .ZN({ S12925 })
);
OAI211_X1 #() 
OAI211_X1_523_ (
  .A({ S12924 }),
  .B({ S25957[404] }),
  .C1({ S18 }),
  .C2({ S12925 }),
  .ZN({ S12926 })
);
INV_X1 #() 
INV_X1_445_ (
  .A({ S12774 }),
  .ZN({ S12927 })
);
AOI22_X1 #() 
AOI22_X1_181_ (
  .A1({ S12720 }),
  .A2({ S25957[400] }),
  .B1({ S18 }),
  .B2({ S12927 }),
  .ZN({ S12929 })
);
OAI211_X1 #() 
OAI211_X1_524_ (
  .A({ S10807 }),
  .B({ S12926 }),
  .C1({ S12929 }),
  .C2({ S25957[404] }),
  .ZN({ S12930 })
);
NAND3_X1 #() 
NAND3_X1_1616_ (
  .A1({ S12709 }),
  .A2({ S12771 }),
  .A3({ S12762 }),
  .ZN({ S12931 })
);
NOR2_X1 #() 
NOR2_X1_321_ (
  .A1({ S18 }),
  .A2({ S12931 }),
  .ZN({ S12932 })
);
NOR3_X1 #() 
NOR3_X1_46_ (
  .A1({ S25957[403] }),
  .A2({ S12839 }),
  .A3({ S12856 }),
  .ZN({ S12933 })
);
OAI21_X1 #() 
OAI21_X1_774_ (
  .A({ S12685 }),
  .B1({ S12933 }),
  .B2({ S12932 }),
  .ZN({ S12934 })
);
NAND2_X1 #() 
NAND2_X1_1387_ (
  .A1({ S12677 }),
  .A2({ S11281 }),
  .ZN({ S12935 })
);
NAND3_X1 #() 
NAND3_X1_1617_ (
  .A1({ S18 }),
  .A2({ S12935 }),
  .A3({ S12774 }),
  .ZN({ S12936 })
);
NAND4_X1 #() 
NAND4_X1_198_ (
  .A1({ S8064 }),
  .A2({ S8067 }),
  .A3({ S11281 }),
  .A4({ S12698 }),
  .ZN({ S12937 })
);
AND2_X1 #() 
AND2_X1_84_ (
  .A1({ S12937 }),
  .A2({ S25957[404] }),
  .ZN({ S12938 })
);
AOI21_X1 #() 
AOI21_X1_839_ (
  .A({ S25957[405] }),
  .B1({ S12938 }),
  .B2({ S12936 }),
  .ZN({ S12940 })
);
NAND2_X1 #() 
NAND2_X1_1388_ (
  .A1({ S25957[403] }),
  .A2({ S12779 }),
  .ZN({ S12941 })
);
OAI211_X1 #() 
OAI211_X1_525_ (
  .A({ S12823 }),
  .B({ S25957[404] }),
  .C1({ S12839 }),
  .C2({ S12941 }),
  .ZN({ S12942 })
);
NAND2_X1 #() 
NAND2_X1_1389_ (
  .A1({ S12679 }),
  .A2({ S40 }),
  .ZN({ S12943 })
);
NAND3_X1 #() 
NAND3_X1_1618_ (
  .A1({ S12943 }),
  .A2({ S8068 }),
  .A3({ S8069 }),
  .ZN({ S12944 })
);
NAND2_X1 #() 
NAND2_X1_1390_ (
  .A1({ S12944 }),
  .A2({ S12691 }),
  .ZN({ S12945 })
);
AOI21_X1 #() 
AOI21_X1_840_ (
  .A({ S10807 }),
  .B1({ S12945 }),
  .B2({ S12685 }),
  .ZN({ S12946 })
);
AOI22_X1 #() 
AOI22_X1_182_ (
  .A1({ S12940 }),
  .A2({ S12934 }),
  .B1({ S12942 }),
  .B2({ S12946 }),
  .ZN({ S12947 })
);
NOR2_X1 #() 
NOR2_X1_322_ (
  .A1({ S18 }),
  .A2({ S12679 }),
  .ZN({ S12948 })
);
AOI21_X1 #() 
AOI21_X1_841_ (
  .A({ S11179 }),
  .B1({ S12679 }),
  .B2({ S12689 }),
  .ZN({ S12949 })
);
AND2_X1 #() 
AND2_X1_85_ (
  .A1({ S18 }),
  .A2({ S12949 }),
  .ZN({ S12951 })
);
OAI21_X1 #() 
OAI21_X1_775_ (
  .A({ S12685 }),
  .B1({ S12951 }),
  .B2({ S12948 }),
  .ZN({ S12952 })
);
AOI21_X1 #() 
AOI21_X1_842_ (
  .A({ S12685 }),
  .B1({ S18 }),
  .B2({ S12839 }),
  .ZN({ S12953 })
);
NAND2_X1 #() 
NAND2_X1_1391_ (
  .A1({ S25957[403] }),
  .A2({ S12935 }),
  .ZN({ S12954 })
);
AOI21_X1 #() 
AOI21_X1_843_ (
  .A({ S10807 }),
  .B1({ S12953 }),
  .B2({ S12954 }),
  .ZN({ S12955 })
);
AOI21_X1 #() 
AOI21_X1_844_ (
  .A({ S25957[406] }),
  .B1({ S12955 }),
  .B2({ S12952 }),
  .ZN({ S12956 })
);
AOI22_X1 #() 
AOI22_X1_183_ (
  .A1({ S12947 }),
  .A2({ S25957[406] }),
  .B1({ S12956 }),
  .B2({ S12930 }),
  .ZN({ S12957 })
);
OAI211_X1 #() 
OAI211_X1_526_ (
  .A({ S12923 }),
  .B({ S25957[509] }),
  .C1({ S25957[407] }),
  .C2({ S12957 }),
  .ZN({ S12958 })
);
INV_X1 #() 
INV_X1_446_ (
  .A({ S25957[509] }),
  .ZN({ S12959 })
);
AND3_X1 #() 
AND3_X1_65_ (
  .A1({ S12907 }),
  .A2({ S12922 }),
  .A3({ S25957[407] }),
  .ZN({ S12960 })
);
NOR2_X1 #() 
NOR2_X1_323_ (
  .A1({ S12957 }),
  .A2({ S25957[407] }),
  .ZN({ S12962 })
);
OAI21_X1 #() 
OAI21_X1_776_ (
  .A({ S12959 }),
  .B1({ S12962 }),
  .B2({ S12960 }),
  .ZN({ S12963 })
);
NAND3_X1 #() 
NAND3_X1_1619_ (
  .A1({ S12963 }),
  .A2({ S12888 }),
  .A3({ S12958 }),
  .ZN({ S12964 })
);
OAI211_X1 #() 
OAI211_X1_527_ (
  .A({ S12923 }),
  .B({ S12959 }),
  .C1({ S25957[407] }),
  .C2({ S12957 }),
  .ZN({ S12965 })
);
OAI21_X1 #() 
OAI21_X1_777_ (
  .A({ S25957[509] }),
  .B1({ S12962 }),
  .B2({ S12960 }),
  .ZN({ S12966 })
);
NAND3_X1 #() 
NAND3_X1_1620_ (
  .A1({ S12966 }),
  .A2({ S25957[573] }),
  .A3({ S12965 }),
  .ZN({ S12967 })
);
NAND3_X1 #() 
NAND3_X1_1621_ (
  .A1({ S12964 }),
  .A2({ S12967 }),
  .A3({ S25957[413] }),
  .ZN({ S12968 })
);
NAND2_X1 #() 
NAND2_X1_1392_ (
  .A1({ S12964 }),
  .A2({ S12967 }),
  .ZN({ S25957[317] })
);
NAND2_X1 #() 
NAND2_X1_1393_ (
  .A1({ S25957[317] }),
  .A2({ S12034 }),
  .ZN({ S12969 })
);
NAND2_X1 #() 
NAND2_X1_1394_ (
  .A1({ S12969 }),
  .A2({ S12968 }),
  .ZN({ S25957[285] })
);
NAND2_X1 #() 
NAND2_X1_1395_ (
  .A1({ S10153 }),
  .A2({ S10155 }),
  .ZN({ S25957[444] })
);
XNOR2_X1 #() 
XNOR2_X1_47_ (
  .A({ S7263 }),
  .B({ S25957[764] }),
  .ZN({ S25957[636] })
);
NAND2_X1 #() 
NAND2_X1_1396_ (
  .A1({ S10148 }),
  .A2({ S10120 }),
  .ZN({ S12971 })
);
XNOR2_X1 #() 
XNOR2_X1_48_ (
  .A({ S12971 }),
  .B({ S25957[636] }),
  .ZN({ S25957[508] })
);
INV_X1 #() 
INV_X1_447_ (
  .A({ S25957[508] }),
  .ZN({ S12972 })
);
AND2_X1 #() 
AND2_X1_86_ (
  .A1({ S12699 }),
  .A2({ S12755 }),
  .ZN({ S12973 })
);
NAND4_X1 #() 
NAND4_X1_199_ (
  .A1({ S12918 }),
  .A2({ S12698 }),
  .A3({ S8064 }),
  .A4({ S8067 }),
  .ZN({ S12974 })
);
OAI211_X1 #() 
OAI211_X1_528_ (
  .A({ S25957[405] }),
  .B({ S12974 }),
  .C1({ S12973 }),
  .C2({ S25957[403] }),
  .ZN({ S12975 })
);
NAND2_X1 #() 
NAND2_X1_1397_ (
  .A1({ S12830 }),
  .A2({ S18 }),
  .ZN({ S12976 })
);
OAI211_X1 #() 
OAI211_X1_529_ (
  .A({ S12976 }),
  .B({ S10807 }),
  .C1({ S18 }),
  .C2({ S12775 }),
  .ZN({ S12977 })
);
AOI21_X1 #() 
AOI21_X1_845_ (
  .A({ S25957[404] }),
  .B1({ S12975 }),
  .B2({ S12977 }),
  .ZN({ S12979 })
);
OAI21_X1 #() 
OAI21_X1_778_ (
  .A({ S12698 }),
  .B1({ S12697 }),
  .B2({ S25957[402] }),
  .ZN({ S12980 })
);
NAND3_X1 #() 
NAND3_X1_1622_ (
  .A1({ S12701 }),
  .A2({ S12677 }),
  .A3({ S12771 }),
  .ZN({ S12981 })
);
NAND2_X1 #() 
NAND2_X1_1398_ (
  .A1({ S18 }),
  .A2({ S12981 }),
  .ZN({ S12982 })
);
OAI211_X1 #() 
OAI211_X1_530_ (
  .A({ S12982 }),
  .B({ S25957[405] }),
  .C1({ S18 }),
  .C2({ S12980 }),
  .ZN({ S12983 })
);
NAND2_X1 #() 
NAND2_X1_1399_ (
  .A1({ S18 }),
  .A2({ S12914 }),
  .ZN({ S12984 })
);
NAND3_X1 #() 
NAND3_X1_1623_ (
  .A1({ S25957[403] }),
  .A2({ S12918 }),
  .A3({ S12765 }),
  .ZN({ S12985 })
);
NAND3_X1 #() 
NAND3_X1_1624_ (
  .A1({ S12985 }),
  .A2({ S10807 }),
  .A3({ S12984 }),
  .ZN({ S12986 })
);
AOI21_X1 #() 
AOI21_X1_846_ (
  .A({ S12685 }),
  .B1({ S12983 }),
  .B2({ S12986 }),
  .ZN({ S12987 })
);
OAI21_X1 #() 
OAI21_X1_779_ (
  .A({ S7784 }),
  .B1({ S12979 }),
  .B2({ S12987 }),
  .ZN({ S12988 })
);
NAND3_X1 #() 
NAND3_X1_1625_ (
  .A1({ S12727 }),
  .A2({ S8068 }),
  .A3({ S8069 }),
  .ZN({ S12990 })
);
NAND2_X1 #() 
NAND2_X1_1400_ (
  .A1({ S12990 }),
  .A2({ S12937 }),
  .ZN({ S12991 })
);
AOI21_X1 #() 
AOI21_X1_847_ (
  .A({ S25957[400] }),
  .B1({ S11281 }),
  .B2({ S25957[401] }),
  .ZN({ S12992 })
);
NAND3_X1 #() 
NAND3_X1_1626_ (
  .A1({ S12992 }),
  .A2({ S8068 }),
  .A3({ S8069 }),
  .ZN({ S12993 })
);
NAND3_X1 #() 
NAND3_X1_1627_ (
  .A1({ S12993 }),
  .A2({ S12685 }),
  .A3({ S12783 }),
  .ZN({ S12994 })
);
OAI211_X1 #() 
OAI211_X1_531_ (
  .A({ S12994 }),
  .B({ S25957[405] }),
  .C1({ S12991 }),
  .C2({ S12685 }),
  .ZN({ S12995 })
);
OAI211_X1 #() 
OAI211_X1_532_ (
  .A({ S12897 }),
  .B({ S25957[404] }),
  .C1({ S12719 }),
  .C2({ S12724 }),
  .ZN({ S12996 })
);
NAND4_X1 #() 
NAND4_X1_200_ (
  .A1({ S8068 }),
  .A2({ S8069 }),
  .A3({ S12701 }),
  .A4({ S12771 }),
  .ZN({ S12997 })
);
NAND3_X1 #() 
NAND3_X1_1628_ (
  .A1({ S12788 }),
  .A2({ S12997 }),
  .A3({ S12685 }),
  .ZN({ S12998 })
);
NAND3_X1 #() 
NAND3_X1_1629_ (
  .A1({ S12996 }),
  .A2({ S10807 }),
  .A3({ S12998 }),
  .ZN({ S12999 })
);
NAND3_X1 #() 
NAND3_X1_1630_ (
  .A1({ S12995 }),
  .A2({ S12999 }),
  .A3({ S25957[406] }),
  .ZN({ S13001 })
);
NAND3_X1 #() 
NAND3_X1_1631_ (
  .A1({ S12988 }),
  .A2({ S13001 }),
  .A3({ S25957[407] }),
  .ZN({ S13002 })
);
NAND2_X1 #() 
NAND2_X1_1401_ (
  .A1({ S18 }),
  .A2({ S39 }),
  .ZN({ S13003 })
);
AOI21_X1 #() 
AOI21_X1_848_ (
  .A({ S25957[404] }),
  .B1({ S12900 }),
  .B2({ S13003 }),
  .ZN({ S13004 })
);
AND3_X1 #() 
AND3_X1_66_ (
  .A1({ S12754 }),
  .A2({ S12909 }),
  .A3({ S25957[404] }),
  .ZN({ S13005 })
);
OAI21_X1 #() 
OAI21_X1_780_ (
  .A({ S25957[405] }),
  .B1({ S13005 }),
  .B2({ S13004 }),
  .ZN({ S13006 })
);
INV_X1 #() 
INV_X1_448_ (
  .A({ S12897 }),
  .ZN({ S13007 })
);
NOR2_X1 #() 
NOR2_X1_324_ (
  .A1({ S18 }),
  .A2({ S12715 }),
  .ZN({ S13008 })
);
OAI21_X1 #() 
OAI21_X1_781_ (
  .A({ S25957[404] }),
  .B1({ S13007 }),
  .B2({ S13008 }),
  .ZN({ S13009 })
);
NAND4_X1 #() 
NAND4_X1_201_ (
  .A1({ S12727 }),
  .A2({ S12733 }),
  .A3({ S8068 }),
  .A4({ S8069 }),
  .ZN({ S13010 })
);
NAND4_X1 #() 
NAND4_X1_202_ (
  .A1({ S8064 }),
  .A2({ S8067 }),
  .A3({ S40 }),
  .A4({ S12679 }),
  .ZN({ S13012 })
);
NAND3_X1 #() 
NAND3_X1_1632_ (
  .A1({ S13010 }),
  .A2({ S12685 }),
  .A3({ S13012 }),
  .ZN({ S13013 })
);
NAND3_X1 #() 
NAND3_X1_1633_ (
  .A1({ S13009 }),
  .A2({ S10807 }),
  .A3({ S13013 }),
  .ZN({ S13014 })
);
NAND3_X1 #() 
NAND3_X1_1634_ (
  .A1({ S13006 }),
  .A2({ S7784 }),
  .A3({ S13014 }),
  .ZN({ S13015 })
);
AOI21_X1 #() 
AOI21_X1_849_ (
  .A({ S25957[403] }),
  .B1({ S12918 }),
  .B2({ S12853 }),
  .ZN({ S13016 })
);
NOR3_X1 #() 
NOR3_X1_47_ (
  .A1({ S13016 }),
  .A2({ S12932 }),
  .A3({ S25957[404] }),
  .ZN({ S13017 })
);
AND2_X1 #() 
AND2_X1_87_ (
  .A1({ S11281 }),
  .A2({ S147 }),
  .ZN({ S13018 })
);
OAI21_X1 #() 
OAI21_X1_782_ (
  .A({ S25957[405] }),
  .B1({ S12685 }),
  .B2({ S13018 }),
  .ZN({ S13019 })
);
INV_X1 #() 
INV_X1_449_ (
  .A({ S12701 }),
  .ZN({ S13020 })
);
OAI211_X1 #() 
OAI211_X1_533_ (
  .A({ S8064 }),
  .B({ S8067 }),
  .C1({ S12856 }),
  .C2({ S11179 }),
  .ZN({ S13021 })
);
NAND3_X1 #() 
NAND3_X1_1635_ (
  .A1({ S12861 }),
  .A2({ S8068 }),
  .A3({ S8069 }),
  .ZN({ S13023 })
);
OAI211_X1 #() 
OAI211_X1_534_ (
  .A({ S13021 }),
  .B({ S25957[404] }),
  .C1({ S13023 }),
  .C2({ S13020 }),
  .ZN({ S13024 })
);
AOI22_X1 #() 
AOI22_X1_184_ (
  .A1({ S12935 }),
  .A2({ S12679 }),
  .B1({ S8064 }),
  .B2({ S8067 }),
  .ZN({ S13025 })
);
NAND2_X1 #() 
NAND2_X1_1402_ (
  .A1({ S25957[403] }),
  .A2({ S25957[402] }),
  .ZN({ S13026 })
);
NAND2_X1 #() 
NAND2_X1_1403_ (
  .A1({ S13026 }),
  .A2({ S12685 }),
  .ZN({ S13027 })
);
OAI211_X1 #() 
OAI211_X1_535_ (
  .A({ S13024 }),
  .B({ S10807 }),
  .C1({ S13027 }),
  .C2({ S13025 }),
  .ZN({ S13028 })
);
OAI211_X1 #() 
OAI211_X1_536_ (
  .A({ S13028 }),
  .B({ S25957[406] }),
  .C1({ S13017 }),
  .C2({ S13019 }),
  .ZN({ S13029 })
);
NAND3_X1 #() 
NAND3_X1_1636_ (
  .A1({ S13015 }),
  .A2({ S7707 }),
  .A3({ S13029 }),
  .ZN({ S13030 })
);
NAND3_X1 #() 
NAND3_X1_1637_ (
  .A1({ S13030 }),
  .A2({ S13002 }),
  .A3({ S12972 }),
  .ZN({ S13031 })
);
OAI21_X1 #() 
OAI21_X1_783_ (
  .A({ S13021 }),
  .B1({ S13023 }),
  .B2({ S13020 }),
  .ZN({ S13032 })
);
NAND2_X1 #() 
NAND2_X1_1404_ (
  .A1({ S13032 }),
  .A2({ S25957[404] }),
  .ZN({ S13034 })
);
NOR2_X1 #() 
NOR2_X1_325_ (
  .A1({ S18 }),
  .A2({ S11281 }),
  .ZN({ S13035 })
);
OAI21_X1 #() 
OAI21_X1_784_ (
  .A({ S12685 }),
  .B1({ S13035 }),
  .B2({ S13025 }),
  .ZN({ S13036 })
);
NAND3_X1 #() 
NAND3_X1_1638_ (
  .A1({ S13034 }),
  .A2({ S10807 }),
  .A3({ S13036 }),
  .ZN({ S13037 })
);
OAI21_X1 #() 
OAI21_X1_785_ (
  .A({ S12685 }),
  .B1({ S13016 }),
  .B2({ S12932 }),
  .ZN({ S13038 })
);
AOI21_X1 #() 
AOI21_X1_850_ (
  .A({ S10807 }),
  .B1({ S25957[404] }),
  .B2({ S13018 }),
  .ZN({ S13039 })
);
NAND2_X1 #() 
NAND2_X1_1405_ (
  .A1({ S13038 }),
  .A2({ S13039 }),
  .ZN({ S13040 })
);
NAND3_X1 #() 
NAND3_X1_1639_ (
  .A1({ S13037 }),
  .A2({ S13040 }),
  .A3({ S25957[406] }),
  .ZN({ S13041 })
);
NAND2_X1 #() 
NAND2_X1_1406_ (
  .A1({ S12900 }),
  .A2({ S13003 }),
  .ZN({ S13042 })
);
NAND2_X1 #() 
NAND2_X1_1407_ (
  .A1({ S13042 }),
  .A2({ S12685 }),
  .ZN({ S13043 })
);
NAND3_X1 #() 
NAND3_X1_1640_ (
  .A1({ S12754 }),
  .A2({ S25957[404] }),
  .A3({ S12909 }),
  .ZN({ S13045 })
);
NAND3_X1 #() 
NAND3_X1_1641_ (
  .A1({ S13043 }),
  .A2({ S25957[405] }),
  .A3({ S13045 }),
  .ZN({ S13046 })
);
OAI211_X1 #() 
OAI211_X1_537_ (
  .A({ S12897 }),
  .B({ S25957[404] }),
  .C1({ S18 }),
  .C2({ S12715 }),
  .ZN({ S13047 })
);
NAND2_X1 #() 
NAND2_X1_1408_ (
  .A1({ S13010 }),
  .A2({ S13012 }),
  .ZN({ S13048 })
);
NAND2_X1 #() 
NAND2_X1_1409_ (
  .A1({ S13048 }),
  .A2({ S12685 }),
  .ZN({ S13049 })
);
NAND3_X1 #() 
NAND3_X1_1642_ (
  .A1({ S13049 }),
  .A2({ S13047 }),
  .A3({ S10807 }),
  .ZN({ S13050 })
);
NAND3_X1 #() 
NAND3_X1_1643_ (
  .A1({ S13046 }),
  .A2({ S13050 }),
  .A3({ S7784 }),
  .ZN({ S13051 })
);
NAND3_X1 #() 
NAND3_X1_1644_ (
  .A1({ S13041 }),
  .A2({ S13051 }),
  .A3({ S7707 }),
  .ZN({ S13052 })
);
NAND2_X1 #() 
NAND2_X1_1410_ (
  .A1({ S12995 }),
  .A2({ S12999 }),
  .ZN({ S13053 })
);
NAND2_X1 #() 
NAND2_X1_1411_ (
  .A1({ S13053 }),
  .A2({ S25957[406] }),
  .ZN({ S13054 })
);
NAND2_X1 #() 
NAND2_X1_1412_ (
  .A1({ S25957[403] }),
  .A2({ S12699 }),
  .ZN({ S13056 })
);
NAND4_X1 #() 
NAND4_X1_203_ (
  .A1({ S12846 }),
  .A2({ S12704 }),
  .A3({ S8068 }),
  .A4({ S8069 }),
  .ZN({ S13057 })
);
OAI21_X1 #() 
OAI21_X1_786_ (
  .A({ S13057 }),
  .B1({ S13056 }),
  .B2({ S12705 }),
  .ZN({ S13058 })
);
AOI22_X1 #() 
AOI22_X1_185_ (
  .A1({ S12699 }),
  .A2({ S12755 }),
  .B1({ S8067 }),
  .B2({ S8064 }),
  .ZN({ S13059 })
);
NAND3_X1 #() 
NAND3_X1_1645_ (
  .A1({ S25957[402] }),
  .A2({ S25957[401] }),
  .A3({ S11081 }),
  .ZN({ S13060 })
);
AOI22_X1 #() 
AOI22_X1_186_ (
  .A1({ S13060 }),
  .A2({ S12851 }),
  .B1({ S8068 }),
  .B2({ S8069 }),
  .ZN({ S13061 })
);
OAI21_X1 #() 
OAI21_X1_787_ (
  .A({ S12685 }),
  .B1({ S13059 }),
  .B2({ S13061 }),
  .ZN({ S13062 })
);
OAI211_X1 #() 
OAI211_X1_538_ (
  .A({ S13062 }),
  .B({ S25957[405] }),
  .C1({ S13058 }),
  .C2({ S12685 }),
  .ZN({ S13063 })
);
NAND2_X1 #() 
NAND2_X1_1413_ (
  .A1({ S12985 }),
  .A2({ S12984 }),
  .ZN({ S13064 })
);
NAND2_X1 #() 
NAND2_X1_1414_ (
  .A1({ S13064 }),
  .A2({ S25957[404] }),
  .ZN({ S13065 })
);
AOI22_X1 #() 
AOI22_X1_187_ (
  .A1({ S12846 }),
  .A2({ S13060 }),
  .B1({ S8064 }),
  .B2({ S8067 }),
  .ZN({ S13067 })
);
NOR2_X1 #() 
NOR2_X1_326_ (
  .A1({ S18 }),
  .A2({ S12775 }),
  .ZN({ S13068 })
);
OAI21_X1 #() 
OAI21_X1_788_ (
  .A({ S12685 }),
  .B1({ S13068 }),
  .B2({ S13067 }),
  .ZN({ S13069 })
);
NAND3_X1 #() 
NAND3_X1_1646_ (
  .A1({ S13065 }),
  .A2({ S10807 }),
  .A3({ S13069 }),
  .ZN({ S13070 })
);
NAND3_X1 #() 
NAND3_X1_1647_ (
  .A1({ S13070 }),
  .A2({ S13063 }),
  .A3({ S7784 }),
  .ZN({ S13071 })
);
NAND3_X1 #() 
NAND3_X1_1648_ (
  .A1({ S13071 }),
  .A2({ S13054 }),
  .A3({ S25957[407] }),
  .ZN({ S13072 })
);
NAND3_X1 #() 
NAND3_X1_1649_ (
  .A1({ S13072 }),
  .A2({ S13052 }),
  .A3({ S25957[508] }),
  .ZN({ S13073 })
);
NAND3_X1 #() 
NAND3_X1_1650_ (
  .A1({ S13031 }),
  .A2({ S13073 }),
  .A3({ S25957[572] }),
  .ZN({ S13074 })
);
NAND3_X1 #() 
NAND3_X1_1651_ (
  .A1({ S13030 }),
  .A2({ S13002 }),
  .A3({ S25957[508] }),
  .ZN({ S13075 })
);
NAND3_X1 #() 
NAND3_X1_1652_ (
  .A1({ S13072 }),
  .A2({ S13052 }),
  .A3({ S12972 }),
  .ZN({ S13076 })
);
NAND3_X1 #() 
NAND3_X1_1653_ (
  .A1({ S13075 }),
  .A2({ S13076 }),
  .A3({ S10092 }),
  .ZN({ S13078 })
);
NAND3_X1 #() 
NAND3_X1_1654_ (
  .A1({ S13074 }),
  .A2({ S13078 }),
  .A3({ S25957[412] }),
  .ZN({ S13079 })
);
NAND3_X1 #() 
NAND3_X1_1655_ (
  .A1({ S13075 }),
  .A2({ S13076 }),
  .A3({ S25957[572] }),
  .ZN({ S13080 })
);
NAND3_X1 #() 
NAND3_X1_1656_ (
  .A1({ S13031 }),
  .A2({ S13073 }),
  .A3({ S10092 }),
  .ZN({ S13081 })
);
NAND3_X1 #() 
NAND3_X1_1657_ (
  .A1({ S13080 }),
  .A2({ S13081 }),
  .A3({ S11984 }),
  .ZN({ S13082 })
);
NAND2_X1 #() 
NAND2_X1_1415_ (
  .A1({ S13079 }),
  .A2({ S13082 }),
  .ZN({ S25957[284] })
);
INV_X1 #() 
INV_X1_450_ (
  .A({ S12765 }),
  .ZN({ S13083 })
);
OAI21_X1 #() 
OAI21_X1_789_ (
  .A({ S12709 }),
  .B1({ S25957[403] }),
  .B2({ S13083 }),
  .ZN({ S13084 })
);
NAND3_X1 #() 
NAND3_X1_1658_ (
  .A1({ S13084 }),
  .A2({ S12685 }),
  .A3({ S25957[400] }),
  .ZN({ S13085 })
);
INV_X1 #() 
INV_X1_451_ (
  .A({ S40 }),
  .ZN({ S13086 })
);
NOR2_X1 #() 
NOR2_X1_327_ (
  .A1({ S25957[403] }),
  .A2({ S12677 }),
  .ZN({ S13088 })
);
OAI211_X1 #() 
OAI211_X1_539_ (
  .A({ S25957[404] }),
  .B({ S25957[402] }),
  .C1({ S13088 }),
  .C2({ S13086 }),
  .ZN({ S13089 })
);
NAND3_X1 #() 
NAND3_X1_1659_ (
  .A1({ S13089 }),
  .A2({ S25957[405] }),
  .A3({ S13085 }),
  .ZN({ S13090 })
);
OAI21_X1 #() 
OAI21_X1_790_ (
  .A({ S40 }),
  .B1({ S12677 }),
  .B2({ S25957[402] }),
  .ZN({ S13091 })
);
OAI211_X1 #() 
OAI211_X1_540_ (
  .A({ S12823 }),
  .B({ S25957[404] }),
  .C1({ S18 }),
  .C2({ S13091 }),
  .ZN({ S13092 })
);
NAND3_X1 #() 
NAND3_X1_1660_ (
  .A1({ S25957[403] }),
  .A2({ S12771 }),
  .A3({ S12725 }),
  .ZN({ S13093 })
);
NAND3_X1 #() 
NAND3_X1_1661_ (
  .A1({ S12763 }),
  .A2({ S13093 }),
  .A3({ S12685 }),
  .ZN({ S13094 })
);
NAND3_X1 #() 
NAND3_X1_1662_ (
  .A1({ S13092 }),
  .A2({ S13094 }),
  .A3({ S10807 }),
  .ZN({ S13095 })
);
AND2_X1 #() 
AND2_X1_88_ (
  .A1({ S13095 }),
  .A2({ S13090 }),
  .ZN({ S13096 })
);
NAND4_X1 #() 
NAND4_X1_204_ (
  .A1({ S8068 }),
  .A2({ S8069 }),
  .A3({ S12677 }),
  .A4({ S12679 }),
  .ZN({ S13097 })
);
INV_X1 #() 
INV_X1_452_ (
  .A({ S13097 }),
  .ZN({ S13099 })
);
NAND2_X1 #() 
NAND2_X1_1416_ (
  .A1({ S13099 }),
  .A2({ S25957[404] }),
  .ZN({ S13100 })
);
OAI211_X1 #() 
OAI211_X1_541_ (
  .A({ S13100 }),
  .B({ S10807 }),
  .C1({ S12872 }),
  .C2({ S13008 }),
  .ZN({ S13101 })
);
AOI22_X1 #() 
AOI22_X1_188_ (
  .A1({ S12890 }),
  .A2({ S12696 }),
  .B1({ S25957[403] }),
  .B2({ S12810 }),
  .ZN({ S13102 })
);
NAND4_X1 #() 
NAND4_X1_205_ (
  .A1({ S8068 }),
  .A2({ S8069 }),
  .A3({ S12765 }),
  .A4({ S12698 }),
  .ZN({ S13103 })
);
NAND3_X1 #() 
NAND3_X1_1663_ (
  .A1({ S12721 }),
  .A2({ S8064 }),
  .A3({ S8067 }),
  .ZN({ S13104 })
);
NAND2_X1 #() 
NAND2_X1_1417_ (
  .A1({ S13104 }),
  .A2({ S13103 }),
  .ZN({ S13105 })
);
NAND2_X1 #() 
NAND2_X1_1418_ (
  .A1({ S13105 }),
  .A2({ S12685 }),
  .ZN({ S13106 })
);
OAI211_X1 #() 
OAI211_X1_542_ (
  .A({ S13106 }),
  .B({ S25957[405] }),
  .C1({ S13102 }),
  .C2({ S12685 }),
  .ZN({ S13107 })
);
NAND3_X1 #() 
NAND3_X1_1664_ (
  .A1({ S13107 }),
  .A2({ S13101 }),
  .A3({ S25957[406] }),
  .ZN({ S13108 })
);
OAI211_X1 #() 
OAI211_X1_543_ (
  .A({ S7707 }),
  .B({ S13108 }),
  .C1({ S13096 }),
  .C2({ S25957[406] }),
  .ZN({ S13110 })
);
NAND4_X1 #() 
NAND4_X1_206_ (
  .A1({ S8064 }),
  .A2({ S8067 }),
  .A3({ S12751 }),
  .A4({ S12677 }),
  .ZN({ S13111 })
);
OAI211_X1 #() 
OAI211_X1_544_ (
  .A({ S25957[404] }),
  .B({ S13111 }),
  .C1({ S12925 }),
  .C2({ S25957[403] }),
  .ZN({ S13112 })
);
NAND2_X1 #() 
NAND2_X1_1419_ (
  .A1({ S18 }),
  .A2({ S12804 }),
  .ZN({ S13113 })
);
AOI21_X1 #() 
AOI21_X1_851_ (
  .A({ S25957[404] }),
  .B1({ S25957[403] }),
  .B2({ S12839 }),
  .ZN({ S13114 })
);
AOI21_X1 #() 
AOI21_X1_852_ (
  .A({ S25957[405] }),
  .B1({ S13114 }),
  .B2({ S13113 }),
  .ZN({ S13115 })
);
INV_X1 #() 
INV_X1_453_ (
  .A({ S13012 }),
  .ZN({ S13116 })
);
NOR3_X1 #() 
NOR3_X1_48_ (
  .A1({ S25957[403] }),
  .A2({ S12773 }),
  .A3({ S12735 }),
  .ZN({ S13117 })
);
OAI21_X1 #() 
OAI21_X1_791_ (
  .A({ S25957[404] }),
  .B1({ S13117 }),
  .B2({ S13116 }),
  .ZN({ S13118 })
);
NAND3_X1 #() 
NAND3_X1_1665_ (
  .A1({ S18 }),
  .A2({ S12698 }),
  .A3({ S12815 }),
  .ZN({ S13119 })
);
NOR2_X1 #() 
NOR2_X1_328_ (
  .A1({ S18 }),
  .A2({ S12981 }),
  .ZN({ S13121 })
);
NOR2_X1 #() 
NOR2_X1_329_ (
  .A1({ S13121 }),
  .A2({ S25957[404] }),
  .ZN({ S13122 })
);
AOI21_X1 #() 
AOI21_X1_853_ (
  .A({ S10807 }),
  .B1({ S13122 }),
  .B2({ S13119 }),
  .ZN({ S13123 })
);
AOI22_X1 #() 
AOI22_X1_189_ (
  .A1({ S13123 }),
  .A2({ S13118 }),
  .B1({ S13115 }),
  .B2({ S13112 }),
  .ZN({ S13124 })
);
NAND3_X1 #() 
NAND3_X1_1666_ (
  .A1({ S13056 }),
  .A2({ S25957[404] }),
  .A3({ S12997 }),
  .ZN({ S13125 })
);
NOR2_X1 #() 
NOR2_X1_330_ (
  .A1({ S12805 }),
  .A2({ S25957[403] }),
  .ZN({ S13126 })
);
AOI22_X1 #() 
AOI22_X1_190_ (
  .A1({ S12774 }),
  .A2({ S12775 }),
  .B1({ S8068 }),
  .B2({ S8069 }),
  .ZN({ S13127 })
);
OAI21_X1 #() 
OAI21_X1_792_ (
  .A({ S12685 }),
  .B1({ S13126 }),
  .B2({ S13127 }),
  .ZN({ S13128 })
);
NAND2_X1 #() 
NAND2_X1_1420_ (
  .A1({ S13128 }),
  .A2({ S13125 }),
  .ZN({ S13129 })
);
NAND2_X1 #() 
NAND2_X1_1421_ (
  .A1({ S12810 }),
  .A2({ S18 }),
  .ZN({ S13130 })
);
NAND3_X1 #() 
NAND3_X1_1667_ (
  .A1({ S25957[403] }),
  .A2({ S12853 }),
  .A3({ S12727 }),
  .ZN({ S13132 })
);
NAND2_X1 #() 
NAND2_X1_1422_ (
  .A1({ S13132 }),
  .A2({ S13130 }),
  .ZN({ S13133 })
);
NAND3_X1 #() 
NAND3_X1_1668_ (
  .A1({ S18 }),
  .A2({ S12701 }),
  .A3({ S12696 }),
  .ZN({ S13134 })
);
NAND2_X1 #() 
NAND2_X1_1423_ (
  .A1({ S25957[403] }),
  .A2({ S12949 }),
  .ZN({ S13135 })
);
NAND3_X1 #() 
NAND3_X1_1669_ (
  .A1({ S13134 }),
  .A2({ S13135 }),
  .A3({ S12685 }),
  .ZN({ S13136 })
);
OAI211_X1 #() 
OAI211_X1_545_ (
  .A({ S13136 }),
  .B({ S25957[405] }),
  .C1({ S13133 }),
  .C2({ S12685 }),
  .ZN({ S13137 })
);
OAI211_X1 #() 
OAI211_X1_546_ (
  .A({ S13137 }),
  .B({ S7784 }),
  .C1({ S13129 }),
  .C2({ S25957[405] }),
  .ZN({ S13138 })
);
OAI211_X1 #() 
OAI211_X1_547_ (
  .A({ S13138 }),
  .B({ S25957[407] }),
  .C1({ S13124 }),
  .C2({ S7784 }),
  .ZN({ S13139 })
);
NAND3_X1 #() 
NAND3_X1_1670_ (
  .A1({ S13110 }),
  .A2({ S25957[795] }),
  .A3({ S13139 }),
  .ZN({ S13140 })
);
NAND2_X1 #() 
NAND2_X1_1424_ (
  .A1({ S13115 }),
  .A2({ S13112 }),
  .ZN({ S13141 })
);
OAI211_X1 #() 
OAI211_X1_548_ (
  .A({ S13119 }),
  .B({ S12685 }),
  .C1({ S18 }),
  .C2({ S12981 }),
  .ZN({ S13143 })
);
NAND3_X1 #() 
NAND3_X1_1671_ (
  .A1({ S13118 }),
  .A2({ S25957[405] }),
  .A3({ S13143 }),
  .ZN({ S13144 })
);
AOI21_X1 #() 
AOI21_X1_854_ (
  .A({ S7784 }),
  .B1({ S13144 }),
  .B2({ S13141 }),
  .ZN({ S13145 })
);
NAND3_X1 #() 
NAND3_X1_1672_ (
  .A1({ S13128 }),
  .A2({ S13125 }),
  .A3({ S10807 }),
  .ZN({ S13146 })
);
AND3_X1 #() 
AND3_X1_67_ (
  .A1({ S13146 }),
  .A2({ S13137 }),
  .A3({ S7784 }),
  .ZN({ S13147 })
);
OAI21_X1 #() 
OAI21_X1_793_ (
  .A({ S25957[407] }),
  .B1({ S13147 }),
  .B2({ S13145 }),
  .ZN({ S13148 })
);
NAND2_X1 #() 
NAND2_X1_1425_ (
  .A1({ S12777 }),
  .A2({ S12812 }),
  .ZN({ S13149 })
);
NAND3_X1 #() 
NAND3_X1_1673_ (
  .A1({ S13104 }),
  .A2({ S13103 }),
  .A3({ S12685 }),
  .ZN({ S13150 })
);
NAND3_X1 #() 
NAND3_X1_1674_ (
  .A1({ S13149 }),
  .A2({ S13150 }),
  .A3({ S25957[405] }),
  .ZN({ S13151 })
);
OAI21_X1 #() 
OAI21_X1_794_ (
  .A({ S13100 }),
  .B1({ S12872 }),
  .B2({ S13008 }),
  .ZN({ S13152 })
);
NAND2_X1 #() 
NAND2_X1_1426_ (
  .A1({ S13152 }),
  .A2({ S10807 }),
  .ZN({ S13154 })
);
AOI21_X1 #() 
AOI21_X1_855_ (
  .A({ S7784 }),
  .B1({ S13154 }),
  .B2({ S13151 }),
  .ZN({ S13155 })
);
AOI21_X1 #() 
AOI21_X1_856_ (
  .A({ S25957[406] }),
  .B1({ S13095 }),
  .B2({ S13090 }),
  .ZN({ S13156 })
);
OAI21_X1 #() 
OAI21_X1_795_ (
  .A({ S7707 }),
  .B1({ S13155 }),
  .B2({ S13156 }),
  .ZN({ S13157 })
);
NAND3_X1 #() 
NAND3_X1_1675_ (
  .A1({ S13148 }),
  .A2({ S13157 }),
  .A3({ S107 }),
  .ZN({ S13158 })
);
AND2_X1 #() 
AND2_X1_89_ (
  .A1({ S13158 }),
  .A2({ S13140 }),
  .ZN({ S41 })
);
NAND2_X1 #() 
NAND2_X1_1427_ (
  .A1({ S13158 }),
  .A2({ S13140 }),
  .ZN({ S25957[283] })
);
XNOR2_X1 #() 
XNOR2_X1_49_ (
  .A({ S25957[632] }),
  .B({ S25957[728] }),
  .ZN({ S13159 })
);
INV_X1 #() 
INV_X1_454_ (
  .A({ S13159 }),
  .ZN({ S25957[600] })
);
OAI211_X1 #() 
OAI211_X1_549_ (
  .A({ S8064 }),
  .B({ S8067 }),
  .C1({ S40 }),
  .C2({ S11281 }),
  .ZN({ S13160 })
);
AOI22_X1 #() 
AOI22_X1_191_ (
  .A1({ S12724 }),
  .A2({ S11179 }),
  .B1({ S12738 }),
  .B2({ S25957[402] }),
  .ZN({ S13162 })
);
OAI211_X1 #() 
OAI211_X1_550_ (
  .A({ S13160 }),
  .B({ S25957[404] }),
  .C1({ S13162 }),
  .C2({ S25957[403] }),
  .ZN({ S13163 })
);
NAND3_X1 #() 
NAND3_X1_1676_ (
  .A1({ S12974 }),
  .A2({ S12990 }),
  .A3({ S12685 }),
  .ZN({ S13164 })
);
NAND3_X1 #() 
NAND3_X1_1677_ (
  .A1({ S13163 }),
  .A2({ S13164 }),
  .A3({ S25957[405] }),
  .ZN({ S13165 })
);
NAND4_X1 #() 
NAND4_X1_207_ (
  .A1({ S12918 }),
  .A2({ S12689 }),
  .A3({ S8068 }),
  .A4({ S8069 }),
  .ZN({ S13166 })
);
NAND3_X1 #() 
NAND3_X1_1678_ (
  .A1({ S13166 }),
  .A2({ S12685 }),
  .A3({ S13104 }),
  .ZN({ S13167 })
);
NAND3_X1 #() 
NAND3_X1_1679_ (
  .A1({ S8064 }),
  .A2({ S8067 }),
  .A3({ S12751 }),
  .ZN({ S13168 })
);
OAI211_X1 #() 
OAI211_X1_551_ (
  .A({ S13168 }),
  .B({ S25957[404] }),
  .C1({ S25957[403] }),
  .C2({ S12703 }),
  .ZN({ S13169 })
);
NAND3_X1 #() 
NAND3_X1_1680_ (
  .A1({ S13167 }),
  .A2({ S13169 }),
  .A3({ S10807 }),
  .ZN({ S13170 })
);
NAND3_X1 #() 
NAND3_X1_1681_ (
  .A1({ S13165 }),
  .A2({ S7784 }),
  .A3({ S13170 }),
  .ZN({ S13171 })
);
NAND2_X1 #() 
NAND2_X1_1428_ (
  .A1({ S12762 }),
  .A2({ S25957[401] }),
  .ZN({ S13173 })
);
NAND4_X1 #() 
NAND4_X1_208_ (
  .A1({ S12752 }),
  .A2({ S13173 }),
  .A3({ S8068 }),
  .A4({ S8069 }),
  .ZN({ S13174 })
);
AOI21_X1 #() 
AOI21_X1_857_ (
  .A({ S25957[404] }),
  .B1({ S25957[403] }),
  .B2({ S12715 }),
  .ZN({ S13175 })
);
NAND3_X1 #() 
NAND3_X1_1682_ (
  .A1({ S12908 }),
  .A2({ S8064 }),
  .A3({ S8067 }),
  .ZN({ S13176 })
);
NAND2_X1 #() 
NAND2_X1_1429_ (
  .A1({ S13010 }),
  .A2({ S13176 }),
  .ZN({ S13177 })
);
AOI22_X1 #() 
AOI22_X1_192_ (
  .A1({ S13177 }),
  .A2({ S25957[404] }),
  .B1({ S13175 }),
  .B2({ S13174 }),
  .ZN({ S13178 })
);
NAND4_X1 #() 
NAND4_X1_209_ (
  .A1({ S12908 }),
  .A2({ S12698 }),
  .A3({ S8064 }),
  .A4({ S8067 }),
  .ZN({ S13179 })
);
NAND3_X1 #() 
NAND3_X1_1683_ (
  .A1({ S13179 }),
  .A2({ S12982 }),
  .A3({ S25957[404] }),
  .ZN({ S13180 })
);
OAI211_X1 #() 
OAI211_X1_552_ (
  .A({ S12685 }),
  .B({ S12710 }),
  .C1({ S12680 }),
  .C2({ S12931 }),
  .ZN({ S13181 })
);
NAND3_X1 #() 
NAND3_X1_1684_ (
  .A1({ S13180 }),
  .A2({ S13181 }),
  .A3({ S10807 }),
  .ZN({ S13182 })
);
OAI211_X1 #() 
OAI211_X1_553_ (
  .A({ S13182 }),
  .B({ S25957[406] }),
  .C1({ S13178 }),
  .C2({ S10807 }),
  .ZN({ S13184 })
);
NAND3_X1 #() 
NAND3_X1_1685_ (
  .A1({ S13184 }),
  .A2({ S25957[407] }),
  .A3({ S13171 }),
  .ZN({ S13185 })
);
NAND3_X1 #() 
NAND3_X1_1686_ (
  .A1({ S12944 }),
  .A2({ S13012 }),
  .A3({ S25957[404] }),
  .ZN({ S13186 })
);
NAND3_X1 #() 
NAND3_X1_1687_ (
  .A1({ S12924 }),
  .A2({ S12862 }),
  .A3({ S12685 }),
  .ZN({ S13187 })
);
NAND3_X1 #() 
NAND3_X1_1688_ (
  .A1({ S13187 }),
  .A2({ S25957[405] }),
  .A3({ S13186 }),
  .ZN({ S13188 })
);
NAND4_X1 #() 
NAND4_X1_210_ (
  .A1({ S12861 }),
  .A2({ S12851 }),
  .A3({ S8068 }),
  .A4({ S8069 }),
  .ZN({ S13189 })
);
NAND2_X1 #() 
NAND2_X1_1430_ (
  .A1({ S25957[403] }),
  .A2({ S12843 }),
  .ZN({ S13190 })
);
NAND3_X1 #() 
NAND3_X1_1689_ (
  .A1({ S13190 }),
  .A2({ S13189 }),
  .A3({ S12685 }),
  .ZN({ S13191 })
);
OAI211_X1 #() 
OAI211_X1_554_ (
  .A({ S12701 }),
  .B({ S40 }),
  .C1({ S12677 }),
  .C2({ S11281 }),
  .ZN({ S13192 })
);
NAND2_X1 #() 
NAND2_X1_1431_ (
  .A1({ S13192 }),
  .A2({ S18 }),
  .ZN({ S13193 })
);
NAND3_X1 #() 
NAND3_X1_1690_ (
  .A1({ S13193 }),
  .A2({ S13056 }),
  .A3({ S25957[404] }),
  .ZN({ S13195 })
);
NAND3_X1 #() 
NAND3_X1_1691_ (
  .A1({ S13195 }),
  .A2({ S13191 }),
  .A3({ S10807 }),
  .ZN({ S13196 })
);
NAND3_X1 #() 
NAND3_X1_1692_ (
  .A1({ S13196 }),
  .A2({ S13188 }),
  .A3({ S7784 }),
  .ZN({ S13197 })
);
NAND3_X1 #() 
NAND3_X1_1693_ (
  .A1({ S25957[403] }),
  .A2({ S12931 }),
  .A3({ S12775 }),
  .ZN({ S13198 })
);
AOI21_X1 #() 
AOI21_X1_858_ (
  .A({ S12685 }),
  .B1({ S18 }),
  .B2({ S12815 }),
  .ZN({ S13199 })
);
AOI22_X1 #() 
AOI22_X1_193_ (
  .A1({ S12690 }),
  .A2({ S12831 }),
  .B1({ S13199 }),
  .B2({ S13198 }),
  .ZN({ S13200 })
);
OAI21_X1 #() 
OAI21_X1_796_ (
  .A({ S12685 }),
  .B1({ S12913 }),
  .B2({ S25957[403] }),
  .ZN({ S13201 })
);
NAND3_X1 #() 
NAND3_X1_1694_ (
  .A1({ S12847 }),
  .A2({ S12691 }),
  .A3({ S25957[404] }),
  .ZN({ S13202 })
);
OAI211_X1 #() 
OAI211_X1_555_ (
  .A({ S13202 }),
  .B({ S10807 }),
  .C1({ S13201 }),
  .C2({ S12932 }),
  .ZN({ S13203 })
);
OAI211_X1 #() 
OAI211_X1_556_ (
  .A({ S25957[406] }),
  .B({ S13203 }),
  .C1({ S13200 }),
  .C2({ S10807 }),
  .ZN({ S13204 })
);
NAND3_X1 #() 
NAND3_X1_1695_ (
  .A1({ S13204 }),
  .A2({ S7707 }),
  .A3({ S13197 }),
  .ZN({ S13206 })
);
AND3_X1 #() 
AND3_X1_68_ (
  .A1({ S13185 }),
  .A2({ S13206 }),
  .A3({ S25957[600] }),
  .ZN({ S13207 })
);
AOI21_X1 #() 
AOI21_X1_859_ (
  .A({ S25957[600] }),
  .B1({ S13185 }),
  .B2({ S13206 }),
  .ZN({ S13208 })
);
OAI21_X1 #() 
OAI21_X1_797_ (
  .A({ S25957[536] }),
  .B1({ S13207 }),
  .B2({ S13208 }),
  .ZN({ S13209 })
);
NAND3_X1 #() 
NAND3_X1_1696_ (
  .A1({ S13185 }),
  .A2({ S13206 }),
  .A3({ S25957[600] }),
  .ZN({ S13210 })
);
NAND3_X1 #() 
NAND3_X1_1697_ (
  .A1({ S13165 }),
  .A2({ S25957[407] }),
  .A3({ S13170 }),
  .ZN({ S13211 })
);
NAND3_X1 #() 
NAND3_X1_1698_ (
  .A1({ S13196 }),
  .A2({ S13188 }),
  .A3({ S7707 }),
  .ZN({ S13212 })
);
NAND2_X1 #() 
NAND2_X1_1432_ (
  .A1({ S13212 }),
  .A2({ S13211 }),
  .ZN({ S13213 })
);
NAND2_X1 #() 
NAND2_X1_1433_ (
  .A1({ S13213 }),
  .A2({ S7784 }),
  .ZN({ S13214 })
);
NAND2_X1 #() 
NAND2_X1_1434_ (
  .A1({ S13175 }),
  .A2({ S13174 }),
  .ZN({ S13215 })
);
NAND2_X1 #() 
NAND2_X1_1435_ (
  .A1({ S13177 }),
  .A2({ S25957[404] }),
  .ZN({ S13217 })
);
NAND3_X1 #() 
NAND3_X1_1699_ (
  .A1({ S13217 }),
  .A2({ S25957[405] }),
  .A3({ S13215 }),
  .ZN({ S13218 })
);
NAND3_X1 #() 
NAND3_X1_1700_ (
  .A1({ S12941 }),
  .A2({ S13057 }),
  .A3({ S25957[404] }),
  .ZN({ S13219 })
);
AOI22_X1 #() 
AOI22_X1_194_ (
  .A1({ S8064 }),
  .A2({ S8067 }),
  .B1({ S12738 }),
  .B2({ S11281 }),
  .ZN({ S13220 })
);
OAI21_X1 #() 
OAI21_X1_798_ (
  .A({ S12685 }),
  .B1({ S12932 }),
  .B2({ S13220 }),
  .ZN({ S13221 })
);
NAND3_X1 #() 
NAND3_X1_1701_ (
  .A1({ S13221 }),
  .A2({ S10807 }),
  .A3({ S13219 }),
  .ZN({ S13222 })
);
AOI21_X1 #() 
AOI21_X1_860_ (
  .A({ S7707 }),
  .B1({ S13218 }),
  .B2({ S13222 }),
  .ZN({ S13223 })
);
NAND2_X1 #() 
NAND2_X1_1436_ (
  .A1({ S12738 }),
  .A2({ S11281 }),
  .ZN({ S13224 })
);
NAND3_X1 #() 
NAND3_X1_1702_ (
  .A1({ S12691 }),
  .A2({ S12709 }),
  .A3({ S13224 }),
  .ZN({ S13225 })
);
NAND2_X1 #() 
NAND2_X1_1437_ (
  .A1({ S13225 }),
  .A2({ S25957[404] }),
  .ZN({ S13226 })
);
AOI22_X1 #() 
AOI22_X1_195_ (
  .A1({ S8064 }),
  .A2({ S8067 }),
  .B1({ S12679 }),
  .B2({ S11179 }),
  .ZN({ S13228 })
);
OAI21_X1 #() 
OAI21_X1_799_ (
  .A({ S12685 }),
  .B1({ S12932 }),
  .B2({ S13228 }),
  .ZN({ S13229 })
);
NAND3_X1 #() 
NAND3_X1_1703_ (
  .A1({ S13229 }),
  .A2({ S13226 }),
  .A3({ S10807 }),
  .ZN({ S13230 })
);
NAND4_X1 #() 
NAND4_X1_211_ (
  .A1({ S8068 }),
  .A2({ S8069 }),
  .A3({ S12697 }),
  .A4({ S12771 }),
  .ZN({ S13231 })
);
OAI211_X1 #() 
OAI211_X1_557_ (
  .A({ S25957[404] }),
  .B({ S13231 }),
  .C1({ S12776 }),
  .C2({ S18 }),
  .ZN({ S13232 })
);
NAND2_X1 #() 
NAND2_X1_1438_ (
  .A1({ S12690 }),
  .A2({ S12831 }),
  .ZN({ S13233 })
);
NAND3_X1 #() 
NAND3_X1_1704_ (
  .A1({ S13233 }),
  .A2({ S13232 }),
  .A3({ S25957[405] }),
  .ZN({ S13234 })
);
AOI21_X1 #() 
AOI21_X1_861_ (
  .A({ S25957[407] }),
  .B1({ S13230 }),
  .B2({ S13234 }),
  .ZN({ S13235 })
);
OAI21_X1 #() 
OAI21_X1_800_ (
  .A({ S25957[406] }),
  .B1({ S13223 }),
  .B2({ S13235 }),
  .ZN({ S13236 })
);
NAND3_X1 #() 
NAND3_X1_1705_ (
  .A1({ S13236 }),
  .A2({ S13159 }),
  .A3({ S13214 }),
  .ZN({ S13237 })
);
NAND3_X1 #() 
NAND3_X1_1706_ (
  .A1({ S13237 }),
  .A2({ S7386 }),
  .A3({ S13210 }),
  .ZN({ S13239 })
);
NAND2_X1 #() 
NAND2_X1_1439_ (
  .A1({ S13209 }),
  .A2({ S13239 }),
  .ZN({ S25957[280] })
);
NAND2_X1 #() 
NAND2_X1_1440_ (
  .A1({ S7459 }),
  .A2({ S7463 }),
  .ZN({ S13240 })
);
INV_X1 #() 
INV_X1_455_ (
  .A({ S13173 }),
  .ZN({ S13241 })
);
AOI21_X1 #() 
AOI21_X1_862_ (
  .A({ S12726 }),
  .B1({ S8068 }),
  .B2({ S8069 }),
  .ZN({ S13242 })
);
AOI22_X1 #() 
AOI22_X1_196_ (
  .A1({ S13242 }),
  .A2({ S13241 }),
  .B1({ S18 }),
  .B2({ S12992 }),
  .ZN({ S13243 })
);
OAI21_X1 #() 
OAI21_X1_801_ (
  .A({ S12872 }),
  .B1({ S13243 }),
  .B2({ S12685 }),
  .ZN({ S13244 })
);
AOI22_X1 #() 
AOI22_X1_197_ (
  .A1({ S12698 }),
  .A2({ S12679 }),
  .B1({ S11179 }),
  .B2({ S25957[402] }),
  .ZN({ S13245 })
);
OAI211_X1 #() 
OAI211_X1_558_ (
  .A({ S12685 }),
  .B({ S12702 }),
  .C1({ S13245 }),
  .C2({ S25957[403] }),
  .ZN({ S13246 })
);
AOI22_X1 #() 
AOI22_X1_198_ (
  .A1({ S8064 }),
  .A2({ S8067 }),
  .B1({ S12765 }),
  .B2({ S12679 }),
  .ZN({ S13247 })
);
NOR2_X1 #() 
NOR2_X1_331_ (
  .A1({ S25957[405] }),
  .A2({ S12685 }),
  .ZN({ S13249 })
);
OAI21_X1 #() 
OAI21_X1_802_ (
  .A({ S13249 }),
  .B1({ S13247 }),
  .B2({ S12686 }),
  .ZN({ S13250 })
);
NAND3_X1 #() 
NAND3_X1_1707_ (
  .A1({ S13250 }),
  .A2({ S7707 }),
  .A3({ S13246 }),
  .ZN({ S13251 })
);
AOI21_X1 #() 
AOI21_X1_863_ (
  .A({ S13251 }),
  .B1({ S13244 }),
  .B2({ S25957[405] }),
  .ZN({ S13252 })
);
NOR2_X1 #() 
NOR2_X1_332_ (
  .A1({ S18 }),
  .A2({ S12765 }),
  .ZN({ S13253 })
);
AOI22_X1 #() 
AOI22_X1_199_ (
  .A1({ S12846 }),
  .A2({ S12751 }),
  .B1({ S8064 }),
  .B2({ S8067 }),
  .ZN({ S13254 })
);
OAI21_X1 #() 
OAI21_X1_803_ (
  .A({ S25957[404] }),
  .B1({ S13253 }),
  .B2({ S13254 }),
  .ZN({ S13255 })
);
OAI21_X1 #() 
OAI21_X1_804_ (
  .A({ S12685 }),
  .B1({ S12759 }),
  .B2({ S13067 }),
  .ZN({ S13256 })
);
NAND3_X1 #() 
NAND3_X1_1708_ (
  .A1({ S13256 }),
  .A2({ S13255 }),
  .A3({ S10807 }),
  .ZN({ S13257 })
);
AOI21_X1 #() 
AOI21_X1_864_ (
  .A({ S12724 }),
  .B1({ S8068 }),
  .B2({ S8069 }),
  .ZN({ S13258 })
);
AOI22_X1 #() 
AOI22_X1_200_ (
  .A1({ S13258 }),
  .A2({ S12696 }),
  .B1({ S18 }),
  .B2({ S12747 }),
  .ZN({ S13260 })
);
AOI22_X1 #() 
AOI22_X1_201_ (
  .A1({ S8068 }),
  .A2({ S8069 }),
  .B1({ S12697 }),
  .B2({ S11281 }),
  .ZN({ S13261 })
);
AOI22_X1 #() 
AOI22_X1_202_ (
  .A1({ S8064 }),
  .A2({ S8067 }),
  .B1({ S12751 }),
  .B2({ S40 }),
  .ZN({ S13262 })
);
OAI21_X1 #() 
OAI21_X1_805_ (
  .A({ S12685 }),
  .B1({ S13262 }),
  .B2({ S13261 }),
  .ZN({ S13263 })
);
OAI211_X1 #() 
OAI211_X1_559_ (
  .A({ S13263 }),
  .B({ S25957[405] }),
  .C1({ S13260 }),
  .C2({ S12685 }),
  .ZN({ S13264 })
);
AOI21_X1 #() 
AOI21_X1_865_ (
  .A({ S7707 }),
  .B1({ S13257 }),
  .B2({ S13264 }),
  .ZN({ S13265 })
);
OAI21_X1 #() 
OAI21_X1_806_ (
  .A({ S7784 }),
  .B1({ S13265 }),
  .B2({ S13252 }),
  .ZN({ S13266 })
);
INV_X1 #() 
INV_X1_456_ (
  .A({ S12891 }),
  .ZN({ S13267 })
);
NAND4_X1 #() 
NAND4_X1_212_ (
  .A1({ S8064 }),
  .A2({ S8067 }),
  .A3({ S12677 }),
  .A4({ S12771 }),
  .ZN({ S13268 })
);
OAI211_X1 #() 
OAI211_X1_560_ (
  .A({ S12685 }),
  .B({ S13268 }),
  .C1({ S13097 }),
  .C2({ S13267 }),
  .ZN({ S13269 })
);
NAND3_X1 #() 
NAND3_X1_1709_ (
  .A1({ S25957[403] }),
  .A2({ S13224 }),
  .A3({ S12779 }),
  .ZN({ S13271 })
);
AOI21_X1 #() 
AOI21_X1_866_ (
  .A({ S12685 }),
  .B1({ S18 }),
  .B2({ S12721 }),
  .ZN({ S13272 })
);
NAND2_X1 #() 
NAND2_X1_1441_ (
  .A1({ S13272 }),
  .A2({ S13271 }),
  .ZN({ S13273 })
);
NAND3_X1 #() 
NAND3_X1_1710_ (
  .A1({ S13273 }),
  .A2({ S13269 }),
  .A3({ S10807 }),
  .ZN({ S13274 })
);
AOI21_X1 #() 
AOI21_X1_867_ (
  .A({ S18 }),
  .B1({ S12696 }),
  .B2({ S12725 }),
  .ZN({ S13275 })
);
NAND3_X1 #() 
NAND3_X1_1711_ (
  .A1({ S12756 }),
  .A2({ S13111 }),
  .A3({ S25957[404] }),
  .ZN({ S13276 })
);
OAI21_X1 #() 
OAI21_X1_807_ (
  .A({ S12685 }),
  .B1({ S25957[403] }),
  .B2({ S12773 }),
  .ZN({ S13277 })
);
OAI211_X1 #() 
OAI211_X1_561_ (
  .A({ S13276 }),
  .B({ S25957[405] }),
  .C1({ S13275 }),
  .C2({ S13277 }),
  .ZN({ S13278 })
);
NAND3_X1 #() 
NAND3_X1_1712_ (
  .A1({ S13274 }),
  .A2({ S13278 }),
  .A3({ S25957[407] }),
  .ZN({ S13279 })
);
NAND4_X1 #() 
NAND4_X1_213_ (
  .A1({ S12719 }),
  .A2({ S12891 }),
  .A3({ S12685 }),
  .A4({ S12679 }),
  .ZN({ S13280 })
);
NAND2_X1 #() 
NAND2_X1_1442_ (
  .A1({ S25957[403] }),
  .A2({ S13091 }),
  .ZN({ S13282 })
);
NAND4_X1 #() 
NAND4_X1_214_ (
  .A1({ S12727 }),
  .A2({ S12762 }),
  .A3({ S8069 }),
  .A4({ S8068 }),
  .ZN({ S13283 })
);
NAND3_X1 #() 
NAND3_X1_1713_ (
  .A1({ S13282 }),
  .A2({ S13283 }),
  .A3({ S25957[404] }),
  .ZN({ S13284 })
);
NAND3_X1 #() 
NAND3_X1_1714_ (
  .A1({ S13284 }),
  .A2({ S25957[405] }),
  .A3({ S13280 }),
  .ZN({ S13285 })
);
NAND4_X1 #() 
NAND4_X1_215_ (
  .A1({ S12891 }),
  .A2({ S12774 }),
  .A3({ S8068 }),
  .A4({ S8069 }),
  .ZN({ S13286 })
);
NAND3_X1 #() 
NAND3_X1_1715_ (
  .A1({ S13198 }),
  .A2({ S25957[404] }),
  .A3({ S13286 }),
  .ZN({ S13287 })
);
NAND3_X1 #() 
NAND3_X1_1716_ (
  .A1({ S13179 }),
  .A2({ S12806 }),
  .A3({ S12685 }),
  .ZN({ S13288 })
);
NAND3_X1 #() 
NAND3_X1_1717_ (
  .A1({ S13287 }),
  .A2({ S13288 }),
  .A3({ S10807 }),
  .ZN({ S13289 })
);
NAND3_X1 #() 
NAND3_X1_1718_ (
  .A1({ S13289 }),
  .A2({ S13285 }),
  .A3({ S7707 }),
  .ZN({ S13290 })
);
NAND2_X1 #() 
NAND2_X1_1443_ (
  .A1({ S13290 }),
  .A2({ S13279 }),
  .ZN({ S13291 })
);
NAND2_X1 #() 
NAND2_X1_1444_ (
  .A1({ S13291 }),
  .A2({ S25957[406] }),
  .ZN({ S13293 })
);
AOI21_X1 #() 
AOI21_X1_868_ (
  .A({ S13240 }),
  .B1({ S13266 }),
  .B2({ S13293 }),
  .ZN({ S13294 })
);
INV_X1 #() 
INV_X1_457_ (
  .A({ S13240 }),
  .ZN({ S25957[601] })
);
NAND3_X1 #() 
NAND3_X1_1719_ (
  .A1({ S13274 }),
  .A2({ S13278 }),
  .A3({ S25957[406] }),
  .ZN({ S13295 })
);
NOR3_X1 #() 
NOR3_X1_49_ (
  .A1({ S12759 }),
  .A2({ S13067 }),
  .A3({ S25957[404] }),
  .ZN({ S13296 })
);
OAI21_X1 #() 
OAI21_X1_808_ (
  .A({ S10807 }),
  .B1({ S12817 }),
  .B2({ S13254 }),
  .ZN({ S13297 })
);
NAND3_X1 #() 
NAND3_X1_1720_ (
  .A1({ S12910 }),
  .A2({ S13103 }),
  .A3({ S12685 }),
  .ZN({ S13298 })
);
NAND3_X1 #() 
NAND3_X1_1721_ (
  .A1({ S25957[403] }),
  .A2({ S12762 }),
  .A3({ S12696 }),
  .ZN({ S13299 })
);
INV_X1 #() 
INV_X1_458_ (
  .A({ S13299 }),
  .ZN({ S13300 })
);
OAI211_X1 #() 
OAI211_X1_562_ (
  .A({ S25957[405] }),
  .B({ S13298 }),
  .C1({ S13300 }),
  .C2({ S12749 }),
  .ZN({ S13301 })
);
OAI211_X1 #() 
OAI211_X1_563_ (
  .A({ S13301 }),
  .B({ S7784 }),
  .C1({ S13297 }),
  .C2({ S13296 }),
  .ZN({ S13303 })
);
NAND3_X1 #() 
NAND3_X1_1722_ (
  .A1({ S13303 }),
  .A2({ S25957[407] }),
  .A3({ S13295 }),
  .ZN({ S13304 })
);
AOI21_X1 #() 
AOI21_X1_869_ (
  .A({ S7784 }),
  .B1({ S13289 }),
  .B2({ S13285 }),
  .ZN({ S13305 })
);
AOI21_X1 #() 
AOI21_X1_870_ (
  .A({ S12685 }),
  .B1({ S13135 }),
  .B2({ S12993 }),
  .ZN({ S13306 })
);
OAI21_X1 #() 
OAI21_X1_809_ (
  .A({ S25957[405] }),
  .B1({ S13306 }),
  .B2({ S12768 }),
  .ZN({ S13307 })
);
NAND3_X1 #() 
NAND3_X1_1723_ (
  .A1({ S13020 }),
  .A2({ S8064 }),
  .A3({ S8067 }),
  .ZN({ S13308 })
);
NAND2_X1 #() 
NAND2_X1_1445_ (
  .A1({ S12679 }),
  .A2({ S12698 }),
  .ZN({ S13309 })
);
NAND4_X1 #() 
NAND4_X1_216_ (
  .A1({ S13309 }),
  .A2({ S8068 }),
  .A3({ S12709 }),
  .A4({ S8069 }),
  .ZN({ S13310 })
);
AOI21_X1 #() 
AOI21_X1_871_ (
  .A({ S25957[404] }),
  .B1({ S13310 }),
  .B2({ S13308 }),
  .ZN({ S13311 })
);
AOI21_X1 #() 
AOI21_X1_872_ (
  .A({ S12685 }),
  .B1({ S13021 }),
  .B2({ S12997 }),
  .ZN({ S13312 })
);
OAI21_X1 #() 
OAI21_X1_810_ (
  .A({ S10807 }),
  .B1({ S13311 }),
  .B2({ S13312 }),
  .ZN({ S13314 })
);
AOI21_X1 #() 
AOI21_X1_873_ (
  .A({ S25957[406] }),
  .B1({ S13307 }),
  .B2({ S13314 }),
  .ZN({ S13315 })
);
OAI21_X1 #() 
OAI21_X1_811_ (
  .A({ S7707 }),
  .B1({ S13315 }),
  .B2({ S13305 }),
  .ZN({ S13316 })
);
AOI21_X1 #() 
AOI21_X1_874_ (
  .A({ S25957[601] }),
  .B1({ S13316 }),
  .B2({ S13304 }),
  .ZN({ S13317 })
);
OAI21_X1 #() 
OAI21_X1_812_ (
  .A({ S25957[537] }),
  .B1({ S13294 }),
  .B2({ S13317 }),
  .ZN({ S13318 })
);
NAND3_X1 #() 
NAND3_X1_1724_ (
  .A1({ S13316 }),
  .A2({ S13304 }),
  .A3({ S25957[601] }),
  .ZN({ S13319 })
);
NAND3_X1 #() 
NAND3_X1_1725_ (
  .A1({ S13266 }),
  .A2({ S13293 }),
  .A3({ S13240 }),
  .ZN({ S13320 })
);
NAND3_X1 #() 
NAND3_X1_1726_ (
  .A1({ S13320 }),
  .A2({ S13319 }),
  .A3({ S9169 }),
  .ZN({ S13321 })
);
NAND2_X1 #() 
NAND2_X1_1446_ (
  .A1({ S13318 }),
  .A2({ S13321 }),
  .ZN({ S25957[281] })
);
OAI21_X1 #() 
OAI21_X1_813_ (
  .A({ S12697 }),
  .B1({ S12698 }),
  .B2({ S11281 }),
  .ZN({ S13322 })
);
OAI21_X1 #() 
OAI21_X1_814_ (
  .A({ S13023 }),
  .B1({ S18 }),
  .B2({ S13322 }),
  .ZN({ S13324 })
);
NAND2_X1 #() 
NAND2_X1_1447_ (
  .A1({ S12701 }),
  .A2({ S25957[400] }),
  .ZN({ S13325 })
);
AOI21_X1 #() 
AOI21_X1_875_ (
  .A({ S12685 }),
  .B1({ S25957[403] }),
  .B2({ S13325 }),
  .ZN({ S13326 })
);
AOI22_X1 #() 
AOI22_X1_203_ (
  .A1({ S13324 }),
  .A2({ S12685 }),
  .B1({ S13326 }),
  .B2({ S12871 }),
  .ZN({ S13327 })
);
NAND3_X1 #() 
NAND3_X1_1727_ (
  .A1({ S12840 }),
  .A2({ S12838 }),
  .A3({ S12685 }),
  .ZN({ S13328 })
);
NAND4_X1 #() 
NAND4_X1_217_ (
  .A1({ S8064 }),
  .A2({ S8067 }),
  .A3({ S25957[401] }),
  .A4({ S12762 }),
  .ZN({ S13329 })
);
OAI211_X1 #() 
OAI211_X1_564_ (
  .A({ S13329 }),
  .B({ S25957[404] }),
  .C1({ S25957[403] }),
  .C2({ S13083 }),
  .ZN({ S13330 })
);
NAND3_X1 #() 
NAND3_X1_1728_ (
  .A1({ S13330 }),
  .A2({ S13328 }),
  .A3({ S10807 }),
  .ZN({ S13331 })
);
OAI211_X1 #() 
OAI211_X1_565_ (
  .A({ S7784 }),
  .B({ S13331 }),
  .C1({ S13327 }),
  .C2({ S10807 }),
  .ZN({ S13332 })
);
OAI21_X1 #() 
OAI21_X1_815_ (
  .A({ S18 }),
  .B1({ S12703 }),
  .B2({ S12821 }),
  .ZN({ S13333 })
);
NAND3_X1 #() 
NAND3_X1_1729_ (
  .A1({ S13333 }),
  .A2({ S25957[404] }),
  .A3({ S12766 }),
  .ZN({ S13335 })
);
NAND2_X1 #() 
NAND2_X1_1448_ (
  .A1({ S12853 }),
  .A2({ S12918 }),
  .ZN({ S13336 })
);
OAI211_X1 #() 
OAI211_X1_566_ (
  .A({ S12787 }),
  .B({ S12685 }),
  .C1({ S13336 }),
  .C2({ S18 }),
  .ZN({ S13337 })
);
NAND3_X1 #() 
NAND3_X1_1730_ (
  .A1({ S13335 }),
  .A2({ S25957[405] }),
  .A3({ S13337 }),
  .ZN({ S13338 })
);
NAND4_X1 #() 
NAND4_X1_218_ (
  .A1({ S12853 }),
  .A2({ S12704 }),
  .A3({ S8064 }),
  .A4({ S8067 }),
  .ZN({ S13339 })
);
NAND3_X1 #() 
NAND3_X1_1731_ (
  .A1({ S13339 }),
  .A2({ S25957[404] }),
  .A3({ S12902 }),
  .ZN({ S13340 })
);
OAI211_X1 #() 
OAI211_X1_567_ (
  .A({ S12788 }),
  .B({ S12685 }),
  .C1({ S25957[403] }),
  .C2({ S12701 }),
  .ZN({ S13341 })
);
NAND3_X1 #() 
NAND3_X1_1732_ (
  .A1({ S13340 }),
  .A2({ S13341 }),
  .A3({ S10807 }),
  .ZN({ S13342 })
);
NAND3_X1 #() 
NAND3_X1_1733_ (
  .A1({ S13338 }),
  .A2({ S25957[406] }),
  .A3({ S13342 }),
  .ZN({ S13343 })
);
NAND3_X1 #() 
NAND3_X1_1734_ (
  .A1({ S13332 }),
  .A2({ S13343 }),
  .A3({ S25957[407] }),
  .ZN({ S13344 })
);
NAND4_X1 #() 
NAND4_X1_219_ (
  .A1({ S8068 }),
  .A2({ S8069 }),
  .A3({ S12679 }),
  .A4({ S12698 }),
  .ZN({ S13346 })
);
AOI21_X1 #() 
AOI21_X1_876_ (
  .A({ S25957[404] }),
  .B1({ S12700 }),
  .B2({ S13346 }),
  .ZN({ S13347 })
);
NAND4_X1 #() 
NAND4_X1_220_ (
  .A1({ S8064 }),
  .A2({ S8067 }),
  .A3({ S12701 }),
  .A4({ S12698 }),
  .ZN({ S13348 })
);
AOI21_X1 #() 
AOI21_X1_877_ (
  .A({ S12685 }),
  .B1({ S13097 }),
  .B2({ S13348 }),
  .ZN({ S13349 })
);
NOR3_X1 #() 
NOR3_X1_50_ (
  .A1({ S13347 }),
  .A2({ S13349 }),
  .A3({ S10807 }),
  .ZN({ S13350 })
);
NAND3_X1 #() 
NAND3_X1_1735_ (
  .A1({ S13057 }),
  .A2({ S12685 }),
  .A3({ S13329 }),
  .ZN({ S13351 })
);
NAND4_X1 #() 
NAND4_X1_221_ (
  .A1({ S12935 }),
  .A2({ S12704 }),
  .A3({ S8068 }),
  .A4({ S8069 }),
  .ZN({ S13352 })
);
NAND4_X1 #() 
NAND4_X1_222_ (
  .A1({ S12846 }),
  .A2({ S12771 }),
  .A3({ S8064 }),
  .A4({ S8067 }),
  .ZN({ S13353 })
);
NAND3_X1 #() 
NAND3_X1_1736_ (
  .A1({ S13352 }),
  .A2({ S13353 }),
  .A3({ S25957[404] }),
  .ZN({ S13354 })
);
NAND3_X1 #() 
NAND3_X1_1737_ (
  .A1({ S13354 }),
  .A2({ S13351 }),
  .A3({ S10807 }),
  .ZN({ S13355 })
);
NAND2_X1 #() 
NAND2_X1_1449_ (
  .A1({ S13355 }),
  .A2({ S25957[406] }),
  .ZN({ S13357 })
);
NOR2_X1 #() 
NOR2_X1_333_ (
  .A1({ S13357 }),
  .A2({ S13350 }),
  .ZN({ S13358 })
);
NAND3_X1 #() 
NAND3_X1_1738_ (
  .A1({ S12831 }),
  .A2({ S12685 }),
  .A3({ S13174 }),
  .ZN({ S13359 })
);
NAND3_X1 #() 
NAND3_X1_1739_ (
  .A1({ S12984 }),
  .A2({ S25957[404] }),
  .A3({ S13329 }),
  .ZN({ S13360 })
);
NAND3_X1 #() 
NAND3_X1_1740_ (
  .A1({ S13359 }),
  .A2({ S13360 }),
  .A3({ S10807 }),
  .ZN({ S13361 })
);
NAND4_X1 #() 
NAND4_X1_223_ (
  .A1({ S12891 }),
  .A2({ S12679 }),
  .A3({ S8067 }),
  .A4({ S8064 }),
  .ZN({ S13362 })
);
NAND3_X1 #() 
NAND3_X1_1741_ (
  .A1({ S13134 }),
  .A2({ S25957[404] }),
  .A3({ S13362 }),
  .ZN({ S13363 })
);
INV_X1 #() 
INV_X1_459_ (
  .A({ S12931 }),
  .ZN({ S13364 })
);
OAI211_X1 #() 
OAI211_X1_568_ (
  .A({ S12840 }),
  .B({ S12685 }),
  .C1({ S13364 }),
  .C2({ S12702 }),
  .ZN({ S13365 })
);
NAND3_X1 #() 
NAND3_X1_1742_ (
  .A1({ S13363 }),
  .A2({ S13365 }),
  .A3({ S25957[405] }),
  .ZN({ S13366 })
);
AOI21_X1 #() 
AOI21_X1_878_ (
  .A({ S25957[406] }),
  .B1({ S13366 }),
  .B2({ S13361 }),
  .ZN({ S13368 })
);
OAI21_X1 #() 
OAI21_X1_816_ (
  .A({ S7707 }),
  .B1({ S13358 }),
  .B2({ S13368 }),
  .ZN({ S13369 })
);
AOI21_X1 #() 
AOI21_X1_879_ (
  .A({ S25957[794] }),
  .B1({ S13369 }),
  .B2({ S13344 }),
  .ZN({ S13370 })
);
AND3_X1 #() 
AND3_X1_69_ (
  .A1({ S13332 }),
  .A2({ S13343 }),
  .A3({ S25957[407] }),
  .ZN({ S13371 })
);
NAND2_X1 #() 
NAND2_X1_1450_ (
  .A1({ S12701 }),
  .A2({ S12762 }),
  .ZN({ S13372 })
);
AOI22_X1 #() 
AOI22_X1_204_ (
  .A1({ S13372 }),
  .A2({ S12698 }),
  .B1({ S8068 }),
  .B2({ S8069 }),
  .ZN({ S13373 })
);
INV_X1 #() 
INV_X1_460_ (
  .A({ S13309 }),
  .ZN({ S13374 })
);
AOI22_X1 #() 
AOI22_X1_205_ (
  .A1({ S13373 }),
  .A2({ S12696 }),
  .B1({ S18 }),
  .B2({ S13374 }),
  .ZN({ S13375 })
);
NAND2_X1 #() 
NAND2_X1_1451_ (
  .A1({ S13097 }),
  .A2({ S13348 }),
  .ZN({ S13376 })
);
NAND2_X1 #() 
NAND2_X1_1452_ (
  .A1({ S13376 }),
  .A2({ S25957[404] }),
  .ZN({ S13377 })
);
OAI211_X1 #() 
OAI211_X1_569_ (
  .A({ S25957[405] }),
  .B({ S13377 }),
  .C1({ S13375 }),
  .C2({ S25957[404] }),
  .ZN({ S13379 })
);
NAND3_X1 #() 
NAND3_X1_1743_ (
  .A1({ S13379 }),
  .A2({ S25957[406] }),
  .A3({ S13355 }),
  .ZN({ S13380 })
);
NAND2_X1 #() 
NAND2_X1_1453_ (
  .A1({ S13366 }),
  .A2({ S13361 }),
  .ZN({ S13381 })
);
NAND2_X1 #() 
NAND2_X1_1454_ (
  .A1({ S13381 }),
  .A2({ S7784 }),
  .ZN({ S13382 })
);
AOI21_X1 #() 
AOI21_X1_880_ (
  .A({ S25957[407] }),
  .B1({ S13382 }),
  .B2({ S13380 }),
  .ZN({ S13383 })
);
NOR3_X1 #() 
NOR3_X1_51_ (
  .A1({ S13383 }),
  .A2({ S13371 }),
  .A3({ S3488 }),
  .ZN({ S13384 })
);
NOR2_X1 #() 
NOR2_X1_334_ (
  .A1({ S13384 }),
  .A2({ S13370 }),
  .ZN({ S25957[282] })
);
NAND3_X1 #() 
NAND3_X1_1744_ (
  .A1({ S11838 }),
  .A2({ S11839 }),
  .A3({ S25957[520] }),
  .ZN({ S13385 })
);
NAND3_X1 #() 
NAND3_X1_1745_ (
  .A1({ S11833 }),
  .A2({ S11836 }),
  .A3({ S7576 }),
  .ZN({ S13386 })
);
AND3_X1 #() 
AND3_X1_70_ (
  .A1({ S13385 }),
  .A2({ S13386 }),
  .A3({ S25957[265] }),
  .ZN({ S42 })
);
OAI21_X1 #() 
OAI21_X1_817_ (
  .A({ S7588 }),
  .B1({ S11883 }),
  .B2({ S11884 }),
  .ZN({ S13388 })
);
NAND3_X1 #() 
NAND3_X1_1746_ (
  .A1({ S11889 }),
  .A2({ S11887 }),
  .A3({ S25957[521] }),
  .ZN({ S13389 })
);
NAND2_X1 #() 
NAND2_X1_1455_ (
  .A1({ S13388 }),
  .A2({ S13389 }),
  .ZN({ S13390 })
);
OAI21_X1 #() 
OAI21_X1_818_ (
  .A({ S13390 }),
  .B1({ S11837 }),
  .B2({ S11840 }),
  .ZN({ S43 })
);
NAND2_X1 #() 
NAND2_X1_1456_ (
  .A1({ S7688 }),
  .A2({ S7693 }),
  .ZN({ S25957[503] })
);
XNOR2_X1 #() 
XNOR2_X1_50_ (
  .A({ S10644 }),
  .B({ S25957[503] }),
  .ZN({ S25957[375] })
);
AND2_X1 #() 
AND2_X1_90_ (
  .A1({ S11504 }),
  .A2({ S11501 }),
  .ZN({ S13391 })
);
OAI21_X1 #() 
OAI21_X1_819_ (
  .A({ S10559 }),
  .B1({ S11584 }),
  .B2({ S11582 }),
  .ZN({ S13392 })
);
NAND3_X1 #() 
NAND3_X1_1747_ (
  .A1({ S11588 }),
  .A2({ S25957[397] }),
  .A3({ S11583 }),
  .ZN({ S13393 })
);
NAND2_X1 #() 
NAND2_X1_1457_ (
  .A1({ S13392 }),
  .A2({ S13393 }),
  .ZN({ S13394 })
);
NAND3_X1 #() 
NAND3_X1_1748_ (
  .A1({ S11970 }),
  .A2({ S25957[265] }),
  .A3({ S11974 }),
  .ZN({ S13396 })
);
AOI21_X1 #() 
AOI21_X1_881_ (
  .A({ S25957[265] }),
  .B1({ S13386 }),
  .B2({ S13385 }),
  .ZN({ S13397 })
);
NAND2_X1 #() 
NAND2_X1_1458_ (
  .A1({ S13397 }),
  .A2({ S25957[266] }),
  .ZN({ S13398 })
);
NAND4_X1 #() 
NAND4_X1_224_ (
  .A1({ S11734 }),
  .A2({ S11735 }),
  .A3({ S13385 }),
  .A4({ S13386 }),
  .ZN({ S13399 })
);
OAI211_X1 #() 
OAI211_X1_570_ (
  .A({ S13398 }),
  .B({ S13396 }),
  .C1({ S25957[266] }),
  .C2({ S13399 }),
  .ZN({ S13400 })
);
NAND3_X1 #() 
NAND3_X1_1749_ (
  .A1({ S11970 }),
  .A2({ S13390 }),
  .A3({ S11974 }),
  .ZN({ S13401 })
);
OAI21_X1 #() 
OAI21_X1_820_ (
  .A({ S25957[265] }),
  .B1({ S11837 }),
  .B2({ S11840 }),
  .ZN({ S13402 })
);
AOI21_X1 #() 
AOI21_X1_882_ (
  .A({ S35 }),
  .B1({ S13402 }),
  .B2({ S13401 }),
  .ZN({ S13403 })
);
AOI21_X1 #() 
AOI21_X1_883_ (
  .A({ S13390 }),
  .B1({ S13386 }),
  .B2({ S13385 }),
  .ZN({ S13404 })
);
NOR2_X1 #() 
NOR2_X1_335_ (
  .A1({ S13404 }),
  .A2({ S25957[267] }),
  .ZN({ S13405 })
);
INV_X1 #() 
INV_X1_461_ (
  .A({ S13405 }),
  .ZN({ S13407 })
);
NAND2_X1 #() 
NAND2_X1_1459_ (
  .A1({ S13407 }),
  .A2({ S25957[268] }),
  .ZN({ S13408 })
);
OAI221_X1 #() 
OAI221_X1_30_ (
  .A({ S13394 }),
  .B1({ S13403 }),
  .B2({ S13408 }),
  .C1({ S13400 }),
  .C2({ S25957[268] }),
  .ZN({ S13409 })
);
NAND3_X1 #() 
NAND3_X1_1750_ (
  .A1({ S11656 }),
  .A2({ S11659 }),
  .A3({ S10526 }),
  .ZN({ S13410 })
);
NAND3_X1 #() 
NAND3_X1_1751_ (
  .A1({ S11661 }),
  .A2({ S11662 }),
  .A3({ S25957[396] }),
  .ZN({ S13411 })
);
NAND2_X1 #() 
NAND2_X1_1460_ (
  .A1({ S13410 }),
  .A2({ S13411 }),
  .ZN({ S13412 })
);
NAND2_X1 #() 
NAND2_X1_1461_ (
  .A1({ S43 }),
  .A2({ S25957[266] }),
  .ZN({ S13413 })
);
OAI21_X1 #() 
OAI21_X1_821_ (
  .A({ S10529 }),
  .B1({ S11966 }),
  .B2({ S11969 }),
  .ZN({ S13414 })
);
NAND3_X1 #() 
NAND3_X1_1752_ (
  .A1({ S11972 }),
  .A2({ S11973 }),
  .A3({ S25957[394] }),
  .ZN({ S13415 })
);
NAND2_X1 #() 
NAND2_X1_1462_ (
  .A1({ S13414 }),
  .A2({ S13415 }),
  .ZN({ S13416 })
);
NAND3_X1 #() 
NAND3_X1_1753_ (
  .A1({ S13385 }),
  .A2({ S13386 }),
  .A3({ S25957[265] }),
  .ZN({ S13418 })
);
NAND2_X1 #() 
NAND2_X1_1463_ (
  .A1({ S13416 }),
  .A2({ S13418 }),
  .ZN({ S13419 })
);
NAND3_X1 #() 
NAND3_X1_1754_ (
  .A1({ S13413 }),
  .A2({ S35 }),
  .A3({ S13419 }),
  .ZN({ S13420 })
);
NAND2_X1 #() 
NAND2_X1_1464_ (
  .A1({ S13396 }),
  .A2({ S25957[267] }),
  .ZN({ S13421 })
);
NAND2_X1 #() 
NAND2_X1_1465_ (
  .A1({ S43 }),
  .A2({ S13418 }),
  .ZN({ S13422 })
);
OAI211_X1 #() 
OAI211_X1_571_ (
  .A({ S13420 }),
  .B({ S13412 }),
  .C1({ S13421 }),
  .C2({ S13422 }),
  .ZN({ S13423 })
);
NAND2_X1 #() 
NAND2_X1_1466_ (
  .A1({ S13385 }),
  .A2({ S13386 }),
  .ZN({ S13424 })
);
NAND3_X1 #() 
NAND3_X1_1755_ (
  .A1({ S13424 }),
  .A2({ S13414 }),
  .A3({ S13415 }),
  .ZN({ S13425 })
);
AND3_X1 #() 
AND3_X1_71_ (
  .A1({ S13385 }),
  .A2({ S13386 }),
  .A3({ S13390 }),
  .ZN({ S13426 })
);
NAND2_X1 #() 
NAND2_X1_1467_ (
  .A1({ S13426 }),
  .A2({ S13416 }),
  .ZN({ S13427 })
);
NAND3_X1 #() 
NAND3_X1_1756_ (
  .A1({ S13427 }),
  .A2({ S25957[267] }),
  .A3({ S13425 }),
  .ZN({ S13429 })
);
AOI21_X1 #() 
AOI21_X1_884_ (
  .A({ S25957[267] }),
  .B1({ S13416 }),
  .B2({ S13424 }),
  .ZN({ S13430 })
);
INV_X1 #() 
INV_X1_462_ (
  .A({ S13430 }),
  .ZN({ S13431 })
);
OAI211_X1 #() 
OAI211_X1_572_ (
  .A({ S13429 }),
  .B({ S25957[268] }),
  .C1({ S13431 }),
  .C2({ S13390 }),
  .ZN({ S13432 })
);
NAND3_X1 #() 
NAND3_X1_1757_ (
  .A1({ S13423 }),
  .A2({ S13432 }),
  .A3({ S25957[269] }),
  .ZN({ S13433 })
);
AOI21_X1 #() 
AOI21_X1_885_ (
  .A({ S13391 }),
  .B1({ S13409 }),
  .B2({ S13433 }),
  .ZN({ S13434 })
);
NAND3_X1 #() 
NAND3_X1_1758_ (
  .A1({ S13414 }),
  .A2({ S25957[265] }),
  .A3({ S13415 }),
  .ZN({ S13435 })
);
NAND3_X1 #() 
NAND3_X1_1759_ (
  .A1({ S43 }),
  .A2({ S25957[266] }),
  .A3({ S13418 }),
  .ZN({ S13436 })
);
NAND3_X1 #() 
NAND3_X1_1760_ (
  .A1({ S13385 }),
  .A2({ S13386 }),
  .A3({ S13390 }),
  .ZN({ S13437 })
);
NAND3_X1 #() 
NAND3_X1_1761_ (
  .A1({ S13402 }),
  .A2({ S13416 }),
  .A3({ S13437 }),
  .ZN({ S13438 })
);
AOI21_X1 #() 
AOI21_X1_886_ (
  .A({ S35 }),
  .B1({ S13438 }),
  .B2({ S13436 }),
  .ZN({ S13440 })
);
AOI21_X1 #() 
AOI21_X1_887_ (
  .A({ S25957[267] }),
  .B1({ S25957[264] }),
  .B2({ S13416 }),
  .ZN({ S13441 })
);
AOI21_X1 #() 
AOI21_X1_888_ (
  .A({ S13440 }),
  .B1({ S13435 }),
  .B2({ S13441 }),
  .ZN({ S13442 })
);
NOR2_X1 #() 
NOR2_X1_336_ (
  .A1({ S13426 }),
  .A2({ S13416 }),
  .ZN({ S13443 })
);
NOR2_X1 #() 
NOR2_X1_337_ (
  .A1({ S13419 }),
  .A2({ S13397 }),
  .ZN({ S13444 })
);
NOR3_X1 #() 
NOR3_X1_52_ (
  .A1({ S13444 }),
  .A2({ S13443 }),
  .A3({ S25957[267] }),
  .ZN({ S13445 })
);
OAI21_X1 #() 
OAI21_X1_822_ (
  .A({ S13412 }),
  .B1({ S13401 }),
  .B2({ S35 }),
  .ZN({ S13446 })
);
OAI22_X1 #() 
OAI22_X1_35_ (
  .A1({ S13442 }),
  .A2({ S13412 }),
  .B1({ S13445 }),
  .B2({ S13446 }),
  .ZN({ S13447 })
);
NAND4_X1 #() 
NAND4_X1_225_ (
  .A1({ S13414 }),
  .A2({ S13415 }),
  .A3({ S13385 }),
  .A4({ S13386 }),
  .ZN({ S13448 })
);
NAND2_X1 #() 
NAND2_X1_1468_ (
  .A1({ S35 }),
  .A2({ S25957[265] }),
  .ZN({ S13449 })
);
INV_X1 #() 
INV_X1_463_ (
  .A({ S13449 }),
  .ZN({ S13451 })
);
NAND2_X1 #() 
NAND2_X1_1469_ (
  .A1({ S25957[267] }),
  .A2({ S13390 }),
  .ZN({ S13452 })
);
OAI211_X1 #() 
OAI211_X1_573_ (
  .A({ S13452 }),
  .B({ S25957[268] }),
  .C1({ S35 }),
  .C2({ S13448 }),
  .ZN({ S13453 })
);
AOI21_X1 #() 
AOI21_X1_889_ (
  .A({ S13453 }),
  .B1({ S13451 }),
  .B2({ S13448 }),
  .ZN({ S13454 })
);
NAND3_X1 #() 
NAND3_X1_1762_ (
  .A1({ S13424 }),
  .A2({ S11970 }),
  .A3({ S11974 }),
  .ZN({ S13455 })
);
AOI21_X1 #() 
AOI21_X1_890_ (
  .A({ S25957[268] }),
  .B1({ S13455 }),
  .B2({ S35 }),
  .ZN({ S13456 })
);
NAND2_X1 #() 
NAND2_X1_1470_ (
  .A1({ S25957[267] }),
  .A2({ S13424 }),
  .ZN({ S13457 })
);
NAND2_X1 #() 
NAND2_X1_1471_ (
  .A1({ S13457 }),
  .A2({ S25957[265] }),
  .ZN({ S13458 })
);
AND2_X1 #() 
AND2_X1_91_ (
  .A1({ S13456 }),
  .A2({ S13458 }),
  .ZN({ S13459 })
);
NOR3_X1 #() 
NOR3_X1_53_ (
  .A1({ S13454 }),
  .A2({ S13459 }),
  .A3({ S13394 }),
  .ZN({ S13460 })
);
AOI21_X1 #() 
AOI21_X1_891_ (
  .A({ S13460 }),
  .B1({ S13447 }),
  .B2({ S13394 }),
  .ZN({ S13462 })
);
NOR2_X1 #() 
NOR2_X1_338_ (
  .A1({ S13462 }),
  .A2({ S25957[270] }),
  .ZN({ S13463 })
);
OAI21_X1 #() 
OAI21_X1_823_ (
  .A({ S25957[271] }),
  .B1({ S13463 }),
  .B2({ S13434 }),
  .ZN({ S13464 })
);
INV_X1 #() 
INV_X1_464_ (
  .A({ S25957[271] }),
  .ZN({ S13465 })
);
NAND3_X1 #() 
NAND3_X1_1763_ (
  .A1({ S13396 }),
  .A2({ S25957[267] }),
  .A3({ S13437 }),
  .ZN({ S13466 })
);
INV_X1 #() 
INV_X1_465_ (
  .A({ S13466 }),
  .ZN({ S13467 })
);
NAND2_X1 #() 
NAND2_X1_1472_ (
  .A1({ S13435 }),
  .A2({ S35 }),
  .ZN({ S13468 })
);
INV_X1 #() 
INV_X1_466_ (
  .A({ S13468 }),
  .ZN({ S13469 })
);
AOI21_X1 #() 
AOI21_X1_892_ (
  .A({ S13467 }),
  .B1({ S13419 }),
  .B2({ S13469 }),
  .ZN({ S13470 })
);
AOI21_X1 #() 
AOI21_X1_893_ (
  .A({ S35 }),
  .B1({ S25957[264] }),
  .B2({ S25957[266] }),
  .ZN({ S13471 })
);
NAND2_X1 #() 
NAND2_X1_1473_ (
  .A1({ S13471 }),
  .A2({ S13401 }),
  .ZN({ S13473 })
);
NAND3_X1 #() 
NAND3_X1_1764_ (
  .A1({ S13473 }),
  .A2({ S25957[268] }),
  .A3({ S13399 }),
  .ZN({ S13474 })
);
OAI211_X1 #() 
OAI211_X1_574_ (
  .A({ S25957[269] }),
  .B({ S13474 }),
  .C1({ S13470 }),
  .C2({ S25957[268] }),
  .ZN({ S13475 })
);
AOI21_X1 #() 
AOI21_X1_894_ (
  .A({ S35 }),
  .B1({ S25957[266] }),
  .B2({ S13418 }),
  .ZN({ S13476 })
);
AOI21_X1 #() 
AOI21_X1_895_ (
  .A({ S25957[267] }),
  .B1({ S13422 }),
  .B2({ S25957[266] }),
  .ZN({ S13477 })
);
OAI21_X1 #() 
OAI21_X1_824_ (
  .A({ S13412 }),
  .B1({ S13477 }),
  .B2({ S13476 }),
  .ZN({ S13478 })
);
AOI21_X1 #() 
AOI21_X1_896_ (
  .A({ S25957[267] }),
  .B1({ S42 }),
  .B2({ S13416 }),
  .ZN({ S13479 })
);
AND2_X1 #() 
AND2_X1_92_ (
  .A1({ S13479 }),
  .A2({ S13436 }),
  .ZN({ S13480 })
);
NOR2_X1 #() 
NOR2_X1_339_ (
  .A1({ S13435 }),
  .A2({ S25957[264] }),
  .ZN({ S13481 })
);
OAI21_X1 #() 
OAI21_X1_825_ (
  .A({ S25957[268] }),
  .B1({ S13481 }),
  .B2({ S35 }),
  .ZN({ S13482 })
);
OAI211_X1 #() 
OAI211_X1_575_ (
  .A({ S13478 }),
  .B({ S13394 }),
  .C1({ S13480 }),
  .C2({ S13482 }),
  .ZN({ S13484 })
);
NAND3_X1 #() 
NAND3_X1_1765_ (
  .A1({ S13484 }),
  .A2({ S13475 }),
  .A3({ S13391 }),
  .ZN({ S13485 })
);
NAND2_X1 #() 
NAND2_X1_1474_ (
  .A1({ S25957[266] }),
  .A2({ S13418 }),
  .ZN({ S13486 })
);
NAND2_X1 #() 
NAND2_X1_1475_ (
  .A1({ S13438 }),
  .A2({ S13486 }),
  .ZN({ S13487 })
);
NAND2_X1 #() 
NAND2_X1_1476_ (
  .A1({ S13487 }),
  .A2({ S25957[267] }),
  .ZN({ S13488 })
);
NAND2_X1 #() 
NAND2_X1_1477_ (
  .A1({ S13441 }),
  .A2({ S13436 }),
  .ZN({ S13489 })
);
NAND3_X1 #() 
NAND3_X1_1766_ (
  .A1({ S13488 }),
  .A2({ S25957[268] }),
  .A3({ S13489 }),
  .ZN({ S13490 })
);
NAND2_X1 #() 
NAND2_X1_1478_ (
  .A1({ S13471 }),
  .A2({ S13396 }),
  .ZN({ S13491 })
);
NAND2_X1 #() 
NAND2_X1_1479_ (
  .A1({ S13416 }),
  .A2({ S13437 }),
  .ZN({ S13492 })
);
NAND2_X1 #() 
NAND2_X1_1480_ (
  .A1({ S13486 }),
  .A2({ S13492 }),
  .ZN({ S13493 })
);
AOI21_X1 #() 
AOI21_X1_897_ (
  .A({ S25957[268] }),
  .B1({ S13493 }),
  .B2({ S35 }),
  .ZN({ S13495 })
);
AOI21_X1 #() 
AOI21_X1_898_ (
  .A({ S25957[269] }),
  .B1({ S13495 }),
  .B2({ S13491 }),
  .ZN({ S13496 })
);
INV_X1 #() 
INV_X1_467_ (
  .A({ S13455 }),
  .ZN({ S13497 })
);
NAND2_X1 #() 
NAND2_X1_1481_ (
  .A1({ S13404 }),
  .A2({ S25957[266] }),
  .ZN({ S13498 })
);
NAND2_X1 #() 
NAND2_X1_1482_ (
  .A1({ S13498 }),
  .A2({ S35 }),
  .ZN({ S13499 })
);
OAI21_X1 #() 
OAI21_X1_826_ (
  .A({ S25957[268] }),
  .B1({ S13499 }),
  .B2({ S13497 }),
  .ZN({ S13500 })
);
NOR2_X1 #() 
NOR2_X1_340_ (
  .A1({ S25957[266] }),
  .A2({ S13418 }),
  .ZN({ S13501 })
);
NAND2_X1 #() 
NAND2_X1_1483_ (
  .A1({ S13398 }),
  .A2({ S25957[267] }),
  .ZN({ S13502 })
);
NOR2_X1 #() 
NOR2_X1_341_ (
  .A1({ S13502 }),
  .A2({ S13501 }),
  .ZN({ S13503 })
);
NAND3_X1 #() 
NAND3_X1_1767_ (
  .A1({ S13414 }),
  .A2({ S13390 }),
  .A3({ S13415 }),
  .ZN({ S13504 })
);
NAND3_X1 #() 
NAND3_X1_1768_ (
  .A1({ S13492 }),
  .A2({ S25957[267] }),
  .A3({ S13504 }),
  .ZN({ S13506 })
);
AOI21_X1 #() 
AOI21_X1_899_ (
  .A({ S25957[267] }),
  .B1({ S25957[266] }),
  .B2({ S13418 }),
  .ZN({ S13507 })
);
INV_X1 #() 
INV_X1_468_ (
  .A({ S13507 }),
  .ZN({ S13508 })
);
NAND3_X1 #() 
NAND3_X1_1769_ (
  .A1({ S13508 }),
  .A2({ S13506 }),
  .A3({ S13412 }),
  .ZN({ S13509 })
);
OAI21_X1 #() 
OAI21_X1_827_ (
  .A({ S13509 }),
  .B1({ S13500 }),
  .B2({ S13503 }),
  .ZN({ S13510 })
);
AOI22_X1 #() 
AOI22_X1_206_ (
  .A1({ S13510 }),
  .A2({ S25957[269] }),
  .B1({ S13496 }),
  .B2({ S13490 }),
  .ZN({ S13511 })
);
OAI21_X1 #() 
OAI21_X1_828_ (
  .A({ S13485 }),
  .B1({ S13511 }),
  .B2({ S13391 }),
  .ZN({ S13512 })
);
NAND2_X1 #() 
NAND2_X1_1484_ (
  .A1({ S13512 }),
  .A2({ S13465 }),
  .ZN({ S13513 })
);
NAND2_X1 #() 
NAND2_X1_1485_ (
  .A1({ S13464 }),
  .A2({ S13513 }),
  .ZN({ S13514 })
);
NAND2_X1 #() 
NAND2_X1_1486_ (
  .A1({ S13514 }),
  .A2({ S25957[375] }),
  .ZN({ S13515 })
);
INV_X1 #() 
INV_X1_469_ (
  .A({ S25957[375] }),
  .ZN({ S13517 })
);
NAND3_X1 #() 
NAND3_X1_1770_ (
  .A1({ S13464 }),
  .A2({ S13517 }),
  .A3({ S13513 }),
  .ZN({ S13518 })
);
NAND2_X1 #() 
NAND2_X1_1487_ (
  .A1({ S13515 }),
  .A2({ S13518 }),
  .ZN({ S25957[247] })
);
INV_X1 #() 
INV_X1_470_ (
  .A({ S25957[247] }),
  .ZN({ S13519 })
);
NAND2_X1 #() 
NAND2_X1_1488_ (
  .A1({ S13519 }),
  .A2({ S25957[343] }),
  .ZN({ S13520 })
);
NAND2_X1 #() 
NAND2_X1_1489_ (
  .A1({ S25957[247] }),
  .A2({ S10648 }),
  .ZN({ S13521 })
);
NAND2_X1 #() 
NAND2_X1_1490_ (
  .A1({ S13520 }),
  .A2({ S13521 }),
  .ZN({ S25957[215] })
);
INV_X1 #() 
INV_X1_471_ (
  .A({ S25957[215] }),
  .ZN({ S13522 })
);
NAND2_X1 #() 
NAND2_X1_1491_ (
  .A1({ S13522 }),
  .A2({ S7707 }),
  .ZN({ S13523 })
);
NAND2_X1 #() 
NAND2_X1_1492_ (
  .A1({ S25957[215] }),
  .A2({ S25957[407] }),
  .ZN({ S13524 })
);
NAND2_X1 #() 
NAND2_X1_1493_ (
  .A1({ S13523 }),
  .A2({ S13524 }),
  .ZN({ S13526 })
);
INV_X1 #() 
INV_X1_472_ (
  .A({ S13526 }),
  .ZN({ S25957[151] })
);
XNOR2_X1 #() 
XNOR2_X1_51_ (
  .A({ S7777 }),
  .B({ S25957[630] }),
  .ZN({ S25957[502] })
);
XNOR2_X1 #() 
XNOR2_X1_52_ (
  .A({ S10723 }),
  .B({ S25957[502] }),
  .ZN({ S25957[374] })
);
INV_X1 #() 
INV_X1_473_ (
  .A({ S25957[374] }),
  .ZN({ S13527 })
);
INV_X1 #() 
INV_X1_474_ (
  .A({ S13422 }),
  .ZN({ S13528 })
);
NAND2_X1 #() 
NAND2_X1_1494_ (
  .A1({ S13404 }),
  .A2({ S13416 }),
  .ZN({ S13529 })
);
NAND3_X1 #() 
NAND3_X1_1771_ (
  .A1({ S13529 }),
  .A2({ S25957[267] }),
  .A3({ S13504 }),
  .ZN({ S13530 })
);
NAND2_X1 #() 
NAND2_X1_1495_ (
  .A1({ S13396 }),
  .A2({ S35 }),
  .ZN({ S13531 })
);
OAI21_X1 #() 
OAI21_X1_829_ (
  .A({ S13530 }),
  .B1({ S13528 }),
  .B2({ S13531 }),
  .ZN({ S13532 })
);
NAND2_X1 #() 
NAND2_X1_1496_ (
  .A1({ S13532 }),
  .A2({ S13412 }),
  .ZN({ S13534 })
);
NAND2_X1 #() 
NAND2_X1_1497_ (
  .A1({ S13443 }),
  .A2({ S13405 }),
  .ZN({ S13535 })
);
NAND3_X1 #() 
NAND3_X1_1772_ (
  .A1({ S25957[266] }),
  .A2({ S25957[267] }),
  .A3({ S25957[265] }),
  .ZN({ S13536 })
);
NAND4_X1 #() 
NAND4_X1_226_ (
  .A1({ S11970 }),
  .A2({ S11734 }),
  .A3({ S11735 }),
  .A4({ S11974 }),
  .ZN({ S13537 })
);
INV_X1 #() 
INV_X1_475_ (
  .A({ S13537 }),
  .ZN({ S13538 })
);
NAND2_X1 #() 
NAND2_X1_1498_ (
  .A1({ S13538 }),
  .A2({ S13404 }),
  .ZN({ S13539 })
);
NAND4_X1 #() 
NAND4_X1_227_ (
  .A1({ S13535 }),
  .A2({ S13539 }),
  .A3({ S25957[268] }),
  .A4({ S13536 }),
  .ZN({ S13540 })
);
NAND3_X1 #() 
NAND3_X1_1773_ (
  .A1({ S13534 }),
  .A2({ S25957[269] }),
  .A3({ S13540 }),
  .ZN({ S13541 })
);
INV_X1 #() 
INV_X1_476_ (
  .A({ S13492 }),
  .ZN({ S13542 })
);
NAND2_X1 #() 
NAND2_X1_1499_ (
  .A1({ S13402 }),
  .A2({ S25957[266] }),
  .ZN({ S13543 })
);
NAND3_X1 #() 
NAND3_X1_1774_ (
  .A1({ S13543 }),
  .A2({ S25957[267] }),
  .A3({ S13401 }),
  .ZN({ S13545 })
);
OAI211_X1 #() 
OAI211_X1_576_ (
  .A({ S13545 }),
  .B({ S25957[268] }),
  .C1({ S25957[267] }),
  .C2({ S13542 }),
  .ZN({ S13546 })
);
NAND4_X1 #() 
NAND4_X1_228_ (
  .A1({ S11970 }),
  .A2({ S11974 }),
  .A3({ S13385 }),
  .A4({ S13386 }),
  .ZN({ S13547 })
);
NAND2_X1 #() 
NAND2_X1_1500_ (
  .A1({ S13547 }),
  .A2({ S13402 }),
  .ZN({ S13548 })
);
NAND3_X1 #() 
NAND3_X1_1775_ (
  .A1({ S13548 }),
  .A2({ S25957[267] }),
  .A3({ S13455 }),
  .ZN({ S13549 })
);
NAND2_X1 #() 
NAND2_X1_1501_ (
  .A1({ S13537 }),
  .A2({ S13399 }),
  .ZN({ S13550 })
);
NAND2_X1 #() 
NAND2_X1_1502_ (
  .A1({ S13438 }),
  .A2({ S13550 }),
  .ZN({ S13551 })
);
NAND3_X1 #() 
NAND3_X1_1776_ (
  .A1({ S13549 }),
  .A2({ S13551 }),
  .A3({ S13412 }),
  .ZN({ S13552 })
);
NAND3_X1 #() 
NAND3_X1_1777_ (
  .A1({ S13546 }),
  .A2({ S13552 }),
  .A3({ S13394 }),
  .ZN({ S13553 })
);
NAND3_X1 #() 
NAND3_X1_1778_ (
  .A1({ S13541 }),
  .A2({ S25957[271] }),
  .A3({ S13553 }),
  .ZN({ S13554 })
);
INV_X1 #() 
INV_X1_477_ (
  .A({ S13504 }),
  .ZN({ S13556 })
);
OAI211_X1 #() 
OAI211_X1_577_ (
  .A({ S13435 }),
  .B({ S35 }),
  .C1({ S25957[266] }),
  .C2({ S13437 }),
  .ZN({ S13557 })
);
OAI211_X1 #() 
OAI211_X1_578_ (
  .A({ S13557 }),
  .B({ S13412 }),
  .C1({ S13556 }),
  .C2({ S13421 }),
  .ZN({ S13558 })
);
INV_X1 #() 
INV_X1_478_ (
  .A({ S13547 }),
  .ZN({ S13559 })
);
AOI21_X1 #() 
AOI21_X1_900_ (
  .A({ S35 }),
  .B1({ S13416 }),
  .B2({ S13424 }),
  .ZN({ S13560 })
);
AOI22_X1 #() 
AOI22_X1_207_ (
  .A1({ S13560 }),
  .A2({ S13422 }),
  .B1({ S13559 }),
  .B2({ S35 }),
  .ZN({ S13561 })
);
OAI211_X1 #() 
OAI211_X1_579_ (
  .A({ S13558 }),
  .B({ S25957[269] }),
  .C1({ S13561 }),
  .C2({ S13412 }),
  .ZN({ S13562 })
);
NOR2_X1 #() 
NOR2_X1_342_ (
  .A1({ S13404 }),
  .A2({ S25957[266] }),
  .ZN({ S13563 })
);
OAI21_X1 #() 
OAI21_X1_830_ (
  .A({ S25957[267] }),
  .B1({ S13481 }),
  .B2({ S13563 }),
  .ZN({ S13564 })
);
AOI22_X1 #() 
AOI22_X1_208_ (
  .A1({ S13564 }),
  .A2({ S13412 }),
  .B1({ S35 }),
  .B2({ S13427 }),
  .ZN({ S13565 })
);
OAI211_X1 #() 
OAI211_X1_580_ (
  .A({ S13565 }),
  .B({ S13394 }),
  .C1({ S13412 }),
  .C2({ S13506 }),
  .ZN({ S13567 })
);
NAND3_X1 #() 
NAND3_X1_1779_ (
  .A1({ S13567 }),
  .A2({ S13465 }),
  .A3({ S13562 }),
  .ZN({ S13568 })
);
NAND2_X1 #() 
NAND2_X1_1503_ (
  .A1({ S13568 }),
  .A2({ S13554 }),
  .ZN({ S13569 })
);
NAND2_X1 #() 
NAND2_X1_1504_ (
  .A1({ S13569 }),
  .A2({ S13391 }),
  .ZN({ S13570 })
);
AOI21_X1 #() 
AOI21_X1_901_ (
  .A({ S35 }),
  .B1({ S13397 }),
  .B2({ S25957[266] }),
  .ZN({ S13571 })
);
NAND2_X1 #() 
NAND2_X1_1505_ (
  .A1({ S13571 }),
  .A2({ S13419 }),
  .ZN({ S13572 })
);
OAI21_X1 #() 
OAI21_X1_831_ (
  .A({ S25957[267] }),
  .B1({ S13416 }),
  .B2({ S13437 }),
  .ZN({ S13573 })
);
OAI21_X1 #() 
OAI21_X1_832_ (
  .A({ S25957[268] }),
  .B1({ S13573 }),
  .B2({ S13497 }),
  .ZN({ S13574 })
);
INV_X1 #() 
INV_X1_479_ (
  .A({ S13574 }),
  .ZN({ S13575 })
);
AOI22_X1 #() 
AOI22_X1_209_ (
  .A1({ S13575 }),
  .A2({ S13551 }),
  .B1({ S13495 }),
  .B2({ S13572 }),
  .ZN({ S13576 })
);
OAI21_X1 #() 
OAI21_X1_833_ (
  .A({ S13412 }),
  .B1({ S13403 }),
  .B2({ S13451 }),
  .ZN({ S13578 })
);
AOI21_X1 #() 
AOI21_X1_902_ (
  .A({ S25957[265] }),
  .B1({ S11735 }),
  .B2({ S11734 }),
  .ZN({ S13579 })
);
NAND3_X1 #() 
NAND3_X1_1780_ (
  .A1({ S13425 }),
  .A2({ S13547 }),
  .A3({ S13579 }),
  .ZN({ S13580 })
);
OAI21_X1 #() 
OAI21_X1_834_ (
  .A({ S13580 }),
  .B1({ S25957[267] }),
  .B2({ S13413 }),
  .ZN({ S13581 })
);
OAI21_X1 #() 
OAI21_X1_835_ (
  .A({ S13578 }),
  .B1({ S13581 }),
  .B2({ S13412 }),
  .ZN({ S13582 })
);
AND2_X1 #() 
AND2_X1_93_ (
  .A1({ S13582 }),
  .A2({ S25957[269] }),
  .ZN({ S13583 })
);
AOI211_X1 #() 
AOI211_X1_19_ (
  .A({ S13465 }),
  .B({ S13583 }),
  .C1({ S13394 }),
  .C2({ S13576 }),
  .ZN({ S13584 })
);
NAND2_X1 #() 
NAND2_X1_1506_ (
  .A1({ S13448 }),
  .A2({ S13402 }),
  .ZN({ S13585 })
);
NAND3_X1 #() 
NAND3_X1_1781_ (
  .A1({ S13486 }),
  .A2({ S35 }),
  .A3({ S13547 }),
  .ZN({ S13586 })
);
NAND2_X1 #() 
NAND2_X1_1507_ (
  .A1({ S13586 }),
  .A2({ S25957[268] }),
  .ZN({ S13587 })
);
AOI21_X1 #() 
AOI21_X1_903_ (
  .A({ S13587 }),
  .B1({ S13585 }),
  .B2({ S25957[267] }),
  .ZN({ S13589 })
);
NOR2_X1 #() 
NOR2_X1_343_ (
  .A1({ S13448 }),
  .A2({ S35 }),
  .ZN({ S13590 })
);
INV_X1 #() 
INV_X1_480_ (
  .A({ S13590 }),
  .ZN({ S13591 })
);
NAND2_X1 #() 
NAND2_X1_1508_ (
  .A1({ S13547 }),
  .A2({ S25957[265] }),
  .ZN({ S13592 })
);
AOI21_X1 #() 
AOI21_X1_904_ (
  .A({ S25957[268] }),
  .B1({ S13591 }),
  .B2({ S13592 }),
  .ZN({ S13593 })
);
OAI21_X1 #() 
OAI21_X1_836_ (
  .A({ S25957[269] }),
  .B1({ S13589 }),
  .B2({ S13593 }),
  .ZN({ S13594 })
);
NAND2_X1 #() 
NAND2_X1_1509_ (
  .A1({ S13401 }),
  .A2({ S13424 }),
  .ZN({ S13595 })
);
NAND2_X1 #() 
NAND2_X1_1510_ (
  .A1({ S13595 }),
  .A2({ S35 }),
  .ZN({ S13596 })
);
AOI21_X1 #() 
AOI21_X1_905_ (
  .A({ S13412 }),
  .B1({ S13596 }),
  .B2({ S13421 }),
  .ZN({ S13597 })
);
NAND2_X1 #() 
NAND2_X1_1511_ (
  .A1({ S13436 }),
  .A2({ S35 }),
  .ZN({ S13598 })
);
NAND2_X1 #() 
NAND2_X1_1512_ (
  .A1({ S13426 }),
  .A2({ S25957[266] }),
  .ZN({ S13600 })
);
AOI21_X1 #() 
AOI21_X1_906_ (
  .A({ S25957[268] }),
  .B1({ S13560 }),
  .B2({ S13600 }),
  .ZN({ S13601 })
);
AOI21_X1 #() 
AOI21_X1_907_ (
  .A({ S13597 }),
  .B1({ S13601 }),
  .B2({ S13598 }),
  .ZN({ S13602 })
);
NAND2_X1 #() 
NAND2_X1_1513_ (
  .A1({ S13602 }),
  .A2({ S13394 }),
  .ZN({ S13603 })
);
AND3_X1 #() 
AND3_X1_72_ (
  .A1({ S13594 }),
  .A2({ S13465 }),
  .A3({ S13603 }),
  .ZN({ S13604 })
);
OAI21_X1 #() 
OAI21_X1_837_ (
  .A({ S25957[270] }),
  .B1({ S13584 }),
  .B2({ S13604 }),
  .ZN({ S13605 })
);
NAND2_X1 #() 
NAND2_X1_1514_ (
  .A1({ S13605 }),
  .A2({ S13570 }),
  .ZN({ S13606 })
);
NAND2_X1 #() 
NAND2_X1_1515_ (
  .A1({ S13606 }),
  .A2({ S13527 }),
  .ZN({ S13607 })
);
NAND3_X1 #() 
NAND3_X1_1782_ (
  .A1({ S13605 }),
  .A2({ S25957[374] }),
  .A3({ S13570 }),
  .ZN({ S13608 })
);
AOI21_X1 #() 
AOI21_X1_908_ (
  .A({ S10726 }),
  .B1({ S13607 }),
  .B2({ S13608 }),
  .ZN({ S13609 })
);
INV_X1 #() 
INV_X1_481_ (
  .A({ S13609 }),
  .ZN({ S13611 })
);
NAND3_X1 #() 
NAND3_X1_1783_ (
  .A1({ S13607 }),
  .A2({ S10726 }),
  .A3({ S13608 }),
  .ZN({ S13612 })
);
AOI21_X1 #() 
AOI21_X1_909_ (
  .A({ S25957[406] }),
  .B1({ S13611 }),
  .B2({ S13612 }),
  .ZN({ S13613 })
);
INV_X1 #() 
INV_X1_482_ (
  .A({ S13612 }),
  .ZN({ S13614 })
);
NOR3_X1 #() 
NOR3_X1_54_ (
  .A1({ S13614 }),
  .A2({ S13609 }),
  .A3({ S7784 }),
  .ZN({ S13615 })
);
NOR2_X1 #() 
NOR2_X1_344_ (
  .A1({ S13613 }),
  .A2({ S13615 }),
  .ZN({ S25957[150] })
);
NAND2_X1 #() 
NAND2_X1_1516_ (
  .A1({ S7867 }),
  .A2({ S7869 }),
  .ZN({ S13616 })
);
INV_X1 #() 
INV_X1_483_ (
  .A({ S13616 }),
  .ZN({ S25957[469] })
);
INV_X1 #() 
INV_X1_484_ (
  .A({ S13448 }),
  .ZN({ S13617 })
);
OAI21_X1 #() 
OAI21_X1_838_ (
  .A({ S13593 }),
  .B1({ S13617 }),
  .B2({ S13538 }),
  .ZN({ S13618 })
);
NAND2_X1 #() 
NAND2_X1_1517_ (
  .A1({ S13419 }),
  .A2({ S25957[267] }),
  .ZN({ S13619 })
);
NAND3_X1 #() 
NAND3_X1_1784_ (
  .A1({ S13539 }),
  .A2({ S25957[268] }),
  .A3({ S13619 }),
  .ZN({ S13620 })
);
NAND3_X1 #() 
NAND3_X1_1785_ (
  .A1({ S13618 }),
  .A2({ S25957[269] }),
  .A3({ S13620 }),
  .ZN({ S13621 })
);
NAND2_X1 #() 
NAND2_X1_1518_ (
  .A1({ S13436 }),
  .A2({ S13492 }),
  .ZN({ S13622 })
);
NAND2_X1 #() 
NAND2_X1_1519_ (
  .A1({ S13622 }),
  .A2({ S25957[267] }),
  .ZN({ S13623 })
);
NAND4_X1 #() 
NAND4_X1_229_ (
  .A1({ S13455 }),
  .A2({ S13437 }),
  .A3({ S35 }),
  .A4({ S13402 }),
  .ZN({ S13624 })
);
NAND3_X1 #() 
NAND3_X1_1786_ (
  .A1({ S13623 }),
  .A2({ S25957[268] }),
  .A3({ S13624 }),
  .ZN({ S13625 })
);
AOI22_X1 #() 
AOI22_X1_210_ (
  .A1({ S13451 }),
  .A2({ S13617 }),
  .B1({ S25957[267] }),
  .B2({ S13426 }),
  .ZN({ S13626 })
);
OAI211_X1 #() 
OAI211_X1_581_ (
  .A({ S13625 }),
  .B({ S13394 }),
  .C1({ S25957[268] }),
  .C2({ S13626 }),
  .ZN({ S13627 })
);
NAND2_X1 #() 
NAND2_X1_1520_ (
  .A1({ S13621 }),
  .A2({ S13627 }),
  .ZN({ S13628 })
);
NAND2_X1 #() 
NAND2_X1_1521_ (
  .A1({ S13628 }),
  .A2({ S13391 }),
  .ZN({ S13630 })
);
NAND3_X1 #() 
NAND3_X1_1787_ (
  .A1({ S13492 }),
  .A2({ S35 }),
  .A3({ S13504 }),
  .ZN({ S13631 })
);
NAND3_X1 #() 
NAND3_X1_1788_ (
  .A1({ S13402 }),
  .A2({ S25957[266] }),
  .A3({ S13437 }),
  .ZN({ S13632 })
);
NAND3_X1 #() 
NAND3_X1_1789_ (
  .A1({ S13632 }),
  .A2({ S25957[267] }),
  .A3({ S13529 }),
  .ZN({ S13633 })
);
NAND3_X1 #() 
NAND3_X1_1790_ (
  .A1({ S13633 }),
  .A2({ S25957[268] }),
  .A3({ S13631 }),
  .ZN({ S13634 })
);
NAND2_X1 #() 
NAND2_X1_1522_ (
  .A1({ S13405 }),
  .A2({ S13547 }),
  .ZN({ S13635 })
);
AND2_X1 #() 
AND2_X1_94_ (
  .A1({ S13635 }),
  .A2({ S13457 }),
  .ZN({ S13636 })
);
OAI21_X1 #() 
OAI21_X1_839_ (
  .A({ S13634 }),
  .B1({ S13636 }),
  .B2({ S25957[268] }),
  .ZN({ S13637 })
);
NAND2_X1 #() 
NAND2_X1_1523_ (
  .A1({ S13476 }),
  .A2({ S13547 }),
  .ZN({ S13638 })
);
NAND3_X1 #() 
NAND3_X1_1791_ (
  .A1({ S13529 }),
  .A2({ S35 }),
  .A3({ S13448 }),
  .ZN({ S13639 })
);
AOI21_X1 #() 
AOI21_X1_910_ (
  .A({ S25957[268] }),
  .B1({ S13638 }),
  .B2({ S13639 }),
  .ZN({ S13641 })
);
AOI21_X1 #() 
AOI21_X1_911_ (
  .A({ S25957[265] }),
  .B1({ S13414 }),
  .B2({ S13415 }),
  .ZN({ S13642 })
);
AOI21_X1 #() 
AOI21_X1_912_ (
  .A({ S13642 }),
  .B1({ S13486 }),
  .B2({ S13547 }),
  .ZN({ S13643 })
);
NAND3_X1 #() 
NAND3_X1_1792_ (
  .A1({ S13416 }),
  .A2({ S25957[267] }),
  .A3({ S13437 }),
  .ZN({ S13644 })
);
NAND2_X1 #() 
NAND2_X1_1524_ (
  .A1({ S13644 }),
  .A2({ S25957[268] }),
  .ZN({ S13645 })
);
AOI21_X1 #() 
AOI21_X1_913_ (
  .A({ S13645 }),
  .B1({ S13643 }),
  .B2({ S35 }),
  .ZN({ S13646 })
);
OR2_X1 #() 
OR2_X1_22_ (
  .A1({ S13646 }),
  .A2({ S25957[269] }),
  .ZN({ S13647 })
);
OAI22_X1 #() 
OAI22_X1_36_ (
  .A1({ S13647 }),
  .A2({ S13641 }),
  .B1({ S13637 }),
  .B2({ S13394 }),
  .ZN({ S13648 })
);
NAND2_X1 #() 
NAND2_X1_1525_ (
  .A1({ S13648 }),
  .A2({ S25957[270] }),
  .ZN({ S13649 })
);
NAND3_X1 #() 
NAND3_X1_1793_ (
  .A1({ S13630 }),
  .A2({ S13649 }),
  .A3({ S13465 }),
  .ZN({ S13650 })
);
NAND2_X1 #() 
NAND2_X1_1526_ (
  .A1({ S13405 }),
  .A2({ S13401 }),
  .ZN({ S13652 })
);
NOR2_X1 #() 
NOR2_X1_345_ (
  .A1({ S25957[268] }),
  .A2({ S13579 }),
  .ZN({ S13653 })
);
NAND3_X1 #() 
NAND3_X1_1794_ (
  .A1({ S13486 }),
  .A2({ S13492 }),
  .A3({ S25957[267] }),
  .ZN({ S13654 })
);
AOI21_X1 #() 
AOI21_X1_914_ (
  .A({ S13412 }),
  .B1({ S13430 }),
  .B2({ S13418 }),
  .ZN({ S13655 })
);
AOI22_X1 #() 
AOI22_X1_211_ (
  .A1({ S13655 }),
  .A2({ S13654 }),
  .B1({ S13653 }),
  .B2({ S13652 }),
  .ZN({ S13656 })
);
NAND2_X1 #() 
NAND2_X1_1527_ (
  .A1({ S13397 }),
  .A2({ S13416 }),
  .ZN({ S13657 })
);
NAND2_X1 #() 
NAND2_X1_1528_ (
  .A1({ S13436 }),
  .A2({ S13657 }),
  .ZN({ S13658 })
);
AOI21_X1 #() 
AOI21_X1_915_ (
  .A({ S13479 }),
  .B1({ S13658 }),
  .B2({ S25957[267] }),
  .ZN({ S13659 })
);
NAND2_X1 #() 
NAND2_X1_1529_ (
  .A1({ S13659 }),
  .A2({ S13412 }),
  .ZN({ S13660 })
);
NAND3_X1 #() 
NAND3_X1_1795_ (
  .A1({ S43 }),
  .A2({ S13416 }),
  .A3({ S13418 }),
  .ZN({ S13661 })
);
NAND2_X1 #() 
NAND2_X1_1530_ (
  .A1({ S13441 }),
  .A2({ S13390 }),
  .ZN({ S13663 })
);
OAI21_X1 #() 
OAI21_X1_840_ (
  .A({ S13663 }),
  .B1({ S35 }),
  .B2({ S13661 }),
  .ZN({ S13664 })
);
AOI21_X1 #() 
AOI21_X1_916_ (
  .A({ S25957[269] }),
  .B1({ S13664 }),
  .B2({ S25957[268] }),
  .ZN({ S13665 })
);
AOI22_X1 #() 
AOI22_X1_212_ (
  .A1({ S13665 }),
  .A2({ S13660 }),
  .B1({ S13656 }),
  .B2({ S25957[269] }),
  .ZN({ S13666 })
);
NAND2_X1 #() 
NAND2_X1_1531_ (
  .A1({ S13666 }),
  .A2({ S13391 }),
  .ZN({ S13667 })
);
NAND2_X1 #() 
NAND2_X1_1532_ (
  .A1({ S13402 }),
  .A2({ S13416 }),
  .ZN({ S13668 })
);
NAND2_X1 #() 
NAND2_X1_1533_ (
  .A1({ S13404 }),
  .A2({ S35 }),
  .ZN({ S13669 })
);
AOI21_X1 #() 
AOI21_X1_917_ (
  .A({ S13412 }),
  .B1({ S13668 }),
  .B2({ S13669 }),
  .ZN({ S13670 })
);
AOI21_X1 #() 
AOI21_X1_918_ (
  .A({ S13670 }),
  .B1({ S13601 }),
  .B2({ S13535 }),
  .ZN({ S13671 })
);
OAI221_X1 #() 
OAI221_X1_31_ (
  .A({ S25957[268] }),
  .B1({ S13457 }),
  .B2({ S13642 }),
  .C1({ S13542 }),
  .C2({ S13407 }),
  .ZN({ S13672 })
);
NAND3_X1 #() 
NAND3_X1_1796_ (
  .A1({ S13435 }),
  .A2({ S25957[267] }),
  .A3({ S13418 }),
  .ZN({ S13674 })
);
INV_X1 #() 
INV_X1_485_ (
  .A({ S13674 }),
  .ZN({ S13675 })
);
NAND2_X1 #() 
NAND2_X1_1534_ (
  .A1({ S13449 }),
  .A2({ S13448 }),
  .ZN({ S13676 })
);
OAI21_X1 #() 
OAI21_X1_841_ (
  .A({ S13412 }),
  .B1({ S13675 }),
  .B2({ S13676 }),
  .ZN({ S13677 })
);
NAND2_X1 #() 
NAND2_X1_1535_ (
  .A1({ S13672 }),
  .A2({ S13677 }),
  .ZN({ S13678 })
);
MUX2_X1 #() 
MUX2_X1_5_ (
  .A({ S13671 }),
  .B({ S13678 }),
  .S({ S25957[269] }),
  .Z({ S13679 })
);
OAI21_X1 #() 
OAI21_X1_842_ (
  .A({ S13667 }),
  .B1({ S13679 }),
  .B2({ S13391 }),
  .ZN({ S13680 })
);
OR2_X1 #() 
OR2_X1_23_ (
  .A1({ S13680 }),
  .A2({ S13465 }),
  .ZN({ S13681 })
);
NAND3_X1 #() 
NAND3_X1_1797_ (
  .A1({ S13681 }),
  .A2({ S25957[469] }),
  .A3({ S13650 }),
  .ZN({ S13682 })
);
NAND2_X1 #() 
NAND2_X1_1536_ (
  .A1({ S13681 }),
  .A2({ S13650 }),
  .ZN({ S13683 })
);
NAND2_X1 #() 
NAND2_X1_1537_ (
  .A1({ S13683 }),
  .A2({ S13616 }),
  .ZN({ S13685 })
);
AOI21_X1 #() 
AOI21_X1_919_ (
  .A({ S10807 }),
  .B1({ S13685 }),
  .B2({ S13682 }),
  .ZN({ S13686 })
);
AND3_X1 #() 
AND3_X1_73_ (
  .A1({ S13685 }),
  .A2({ S13682 }),
  .A3({ S10807 }),
  .ZN({ S13687 })
);
NOR2_X1 #() 
NOR2_X1_346_ (
  .A1({ S13687 }),
  .A2({ S13686 }),
  .ZN({ S13688 })
);
INV_X1 #() 
INV_X1_486_ (
  .A({ S13688 }),
  .ZN({ S25957[149] })
);
NAND2_X1 #() 
NAND2_X1_1538_ (
  .A1({ S10894 }),
  .A2({ S10898 }),
  .ZN({ S25957[340] })
);
XNOR2_X1 #() 
XNOR2_X1_53_ (
  .A({ S25957[340] }),
  .B({ S10811 }),
  .ZN({ S25957[308] })
);
NAND2_X1 #() 
NAND2_X1_1539_ (
  .A1({ S10893 }),
  .A2({ S10874 }),
  .ZN({ S25957[372] })
);
INV_X1 #() 
INV_X1_487_ (
  .A({ S25957[372] }),
  .ZN({ S13689 })
);
NOR2_X1 #() 
NOR2_X1_347_ (
  .A1({ S13396 }),
  .A2({ S25957[264] }),
  .ZN({ S13690 })
);
AOI21_X1 #() 
AOI21_X1_920_ (
  .A({ S13437 }),
  .B1({ S13416 }),
  .B2({ S35 }),
  .ZN({ S13692 })
);
OAI21_X1 #() 
OAI21_X1_843_ (
  .A({ S25957[268] }),
  .B1({ S13692 }),
  .B2({ S13690 }),
  .ZN({ S13693 })
);
AOI21_X1 #() 
AOI21_X1_921_ (
  .A({ S25957[267] }),
  .B1({ S13438 }),
  .B2({ S13486 }),
  .ZN({ S13694 })
);
NAND2_X1 #() 
NAND2_X1_1540_ (
  .A1({ S13404 }),
  .A2({ S25957[267] }),
  .ZN({ S13695 })
);
NAND3_X1 #() 
NAND3_X1_1798_ (
  .A1({ S13644 }),
  .A2({ S13695 }),
  .A3({ S13412 }),
  .ZN({ S13696 })
);
OAI21_X1 #() 
OAI21_X1_844_ (
  .A({ S13693 }),
  .B1({ S13694 }),
  .B2({ S13696 }),
  .ZN({ S13697 })
);
NOR2_X1 #() 
NOR2_X1_348_ (
  .A1({ S13617 }),
  .A2({ S13452 }),
  .ZN({ S13698 })
);
INV_X1 #() 
INV_X1_488_ (
  .A({ S13698 }),
  .ZN({ S13699 })
);
NAND2_X1 #() 
NAND2_X1_1541_ (
  .A1({ S13668 }),
  .A2({ S13498 }),
  .ZN({ S13700 })
);
NAND2_X1 #() 
NAND2_X1_1542_ (
  .A1({ S13700 }),
  .A2({ S35 }),
  .ZN({ S13701 })
);
NAND3_X1 #() 
NAND3_X1_1799_ (
  .A1({ S13701 }),
  .A2({ S13699 }),
  .A3({ S13412 }),
  .ZN({ S13702 })
);
NAND4_X1 #() 
NAND4_X1_230_ (
  .A1({ S13396 }),
  .A2({ S13504 }),
  .A3({ S25957[267] }),
  .A4({ S13418 }),
  .ZN({ S13703 })
);
OAI211_X1 #() 
OAI211_X1_582_ (
  .A({ S25957[268] }),
  .B({ S13703 }),
  .C1({ S13499 }),
  .C2({ S13501 }),
  .ZN({ S13704 })
);
NAND3_X1 #() 
NAND3_X1_1800_ (
  .A1({ S13702 }),
  .A2({ S13394 }),
  .A3({ S13704 }),
  .ZN({ S13705 })
);
OAI211_X1 #() 
OAI211_X1_583_ (
  .A({ S13705 }),
  .B({ S13391 }),
  .C1({ S13394 }),
  .C2({ S13697 }),
  .ZN({ S13706 })
);
NAND2_X1 #() 
NAND2_X1_1543_ (
  .A1({ S13398 }),
  .A2({ S35 }),
  .ZN({ S13707 })
);
NAND3_X1 #() 
NAND3_X1_1801_ (
  .A1({ S13707 }),
  .A2({ S25957[268] }),
  .A3({ S13644 }),
  .ZN({ S13708 })
);
NAND3_X1 #() 
NAND3_X1_1802_ (
  .A1({ S13396 }),
  .A2({ S35 }),
  .A3({ S13424 }),
  .ZN({ S13709 })
);
NAND3_X1 #() 
NAND3_X1_1803_ (
  .A1({ S13473 }),
  .A2({ S13412 }),
  .A3({ S13709 }),
  .ZN({ S13710 })
);
NAND3_X1 #() 
NAND3_X1_1804_ (
  .A1({ S13710 }),
  .A2({ S13708 }),
  .A3({ S25957[269] }),
  .ZN({ S13711 })
);
NAND2_X1 #() 
NAND2_X1_1544_ (
  .A1({ S13425 }),
  .A2({ S13401 }),
  .ZN({ S13713 })
);
OAI211_X1 #() 
OAI211_X1_584_ (
  .A({ S13412 }),
  .B({ S13466 }),
  .C1({ S13713 }),
  .C2({ S25957[267] }),
  .ZN({ S13714 })
);
AOI21_X1 #() 
AOI21_X1_922_ (
  .A({ S13412 }),
  .B1({ S13405 }),
  .B2({ S13401 }),
  .ZN({ S13715 })
);
OAI21_X1 #() 
OAI21_X1_845_ (
  .A({ S13715 }),
  .B1({ S13559 }),
  .B2({ S13452 }),
  .ZN({ S13716 })
);
NAND3_X1 #() 
NAND3_X1_1805_ (
  .A1({ S13716 }),
  .A2({ S13394 }),
  .A3({ S13714 }),
  .ZN({ S13717 })
);
NAND3_X1 #() 
NAND3_X1_1806_ (
  .A1({ S13717 }),
  .A2({ S25957[270] }),
  .A3({ S13711 }),
  .ZN({ S13718 })
);
NAND3_X1 #() 
NAND3_X1_1807_ (
  .A1({ S13706 }),
  .A2({ S25957[271] }),
  .A3({ S13718 }),
  .ZN({ S13719 })
);
OAI21_X1 #() 
OAI21_X1_846_ (
  .A({ S13396 }),
  .B1({ S43 }),
  .B2({ S13416 }),
  .ZN({ S13720 })
);
NAND2_X1 #() 
NAND2_X1_1545_ (
  .A1({ S13547 }),
  .A2({ S35 }),
  .ZN({ S13721 })
);
NAND3_X1 #() 
NAND3_X1_1808_ (
  .A1({ S13448 }),
  .A2({ S43 }),
  .A3({ S25957[267] }),
  .ZN({ S13722 })
);
OAI21_X1 #() 
OAI21_X1_847_ (
  .A({ S13722 }),
  .B1({ S13720 }),
  .B2({ S13721 }),
  .ZN({ S13724 })
);
NAND2_X1 #() 
NAND2_X1_1546_ (
  .A1({ S13724 }),
  .A2({ S13412 }),
  .ZN({ S13725 })
);
NAND2_X1 #() 
NAND2_X1_1547_ (
  .A1({ S13401 }),
  .A2({ S25957[264] }),
  .ZN({ S13726 })
);
NAND2_X1 #() 
NAND2_X1_1548_ (
  .A1({ S13560 }),
  .A2({ S13726 }),
  .ZN({ S13727 })
);
AOI21_X1 #() 
AOI21_X1_923_ (
  .A({ S25957[269] }),
  .B1({ S13715 }),
  .B2({ S13727 }),
  .ZN({ S13728 })
);
NAND2_X1 #() 
NAND2_X1_1549_ (
  .A1({ S13725 }),
  .A2({ S13728 }),
  .ZN({ S13729 })
);
AOI22_X1 #() 
AOI22_X1_213_ (
  .A1({ S13444 }),
  .A2({ S25957[267] }),
  .B1({ S13451 }),
  .B2({ S25957[264] }),
  .ZN({ S13730 })
);
OAI211_X1 #() 
OAI211_X1_585_ (
  .A({ S13506 }),
  .B({ S25957[268] }),
  .C1({ S25957[267] }),
  .C2({ S13543 }),
  .ZN({ S13731 })
);
OAI211_X1 #() 
OAI211_X1_586_ (
  .A({ S13731 }),
  .B({ S25957[269] }),
  .C1({ S13730 }),
  .C2({ S25957[268] }),
  .ZN({ S13732 })
);
AND2_X1 #() 
AND2_X1_95_ (
  .A1({ S13732 }),
  .A2({ S13729 }),
  .ZN({ S13733 })
);
OAI211_X1 #() 
OAI211_X1_587_ (
  .A({ S35 }),
  .B({ S13401 }),
  .C1({ S13397 }),
  .C2({ S13416 }),
  .ZN({ S13734 })
);
INV_X1 #() 
INV_X1_489_ (
  .A({ S13734 }),
  .ZN({ S13735 })
);
NAND2_X1 #() 
NAND2_X1_1550_ (
  .A1({ S42 }),
  .A2({ S13416 }),
  .ZN({ S13736 })
);
NAND3_X1 #() 
NAND3_X1_1809_ (
  .A1({ S13736 }),
  .A2({ S35 }),
  .A3({ S13425 }),
  .ZN({ S13737 })
);
NOR2_X1 #() 
NOR2_X1_349_ (
  .A1({ S13416 }),
  .A2({ S35 }),
  .ZN({ S13738 })
);
NOR2_X1 #() 
NOR2_X1_350_ (
  .A1({ S13738 }),
  .A2({ S25957[268] }),
  .ZN({ S13739 })
);
NAND2_X1 #() 
NAND2_X1_1551_ (
  .A1({ S13737 }),
  .A2({ S13739 }),
  .ZN({ S13740 })
);
OAI211_X1 #() 
OAI211_X1_588_ (
  .A({ S13740 }),
  .B({ S13394 }),
  .C1({ S13453 }),
  .C2({ S13735 }),
  .ZN({ S13741 })
);
AOI21_X1 #() 
AOI21_X1_924_ (
  .A({ S25957[267] }),
  .B1({ S13661 }),
  .B2({ S13543 }),
  .ZN({ S13742 })
);
INV_X1 #() 
INV_X1_490_ (
  .A({ S148 }),
  .ZN({ S13743 })
);
OAI21_X1 #() 
OAI21_X1_848_ (
  .A({ S25957[268] }),
  .B1({ S13743 }),
  .B2({ S25957[266] }),
  .ZN({ S13745 })
);
NAND2_X1 #() 
NAND2_X1_1552_ (
  .A1({ S13638 }),
  .A2({ S13412 }),
  .ZN({ S13746 })
);
OAI211_X1 #() 
OAI211_X1_589_ (
  .A({ S25957[269] }),
  .B({ S13745 }),
  .C1({ S13746 }),
  .C2({ S13742 }),
  .ZN({ S13747 })
);
NAND3_X1 #() 
NAND3_X1_1810_ (
  .A1({ S13747 }),
  .A2({ S13741 }),
  .A3({ S25957[270] }),
  .ZN({ S13748 })
);
OAI211_X1 #() 
OAI211_X1_590_ (
  .A({ S13465 }),
  .B({ S13748 }),
  .C1({ S13733 }),
  .C2({ S25957[270] }),
  .ZN({ S13749 })
);
NAND3_X1 #() 
NAND3_X1_1811_ (
  .A1({ S13749 }),
  .A2({ S13719 }),
  .A3({ S13689 }),
  .ZN({ S13750 })
);
AOI21_X1 #() 
AOI21_X1_925_ (
  .A({ S25957[271] }),
  .B1({ S13732 }),
  .B2({ S13729 }),
  .ZN({ S13751 })
);
OAI21_X1 #() 
OAI21_X1_849_ (
  .A({ S13703 }),
  .B1({ S13499 }),
  .B2({ S13501 }),
  .ZN({ S13752 })
);
NAND2_X1 #() 
NAND2_X1_1553_ (
  .A1({ S13752 }),
  .A2({ S25957[268] }),
  .ZN({ S13753 })
);
AOI21_X1 #() 
AOI21_X1_926_ (
  .A({ S25957[267] }),
  .B1({ S13668 }),
  .B2({ S13498 }),
  .ZN({ S13754 })
);
OAI21_X1 #() 
OAI21_X1_850_ (
  .A({ S13412 }),
  .B1({ S13754 }),
  .B2({ S13698 }),
  .ZN({ S13756 })
);
NAND3_X1 #() 
NAND3_X1_1812_ (
  .A1({ S13753 }),
  .A2({ S13756 }),
  .A3({ S13394 }),
  .ZN({ S13757 })
);
NAND2_X1 #() 
NAND2_X1_1554_ (
  .A1({ S13697 }),
  .A2({ S25957[269] }),
  .ZN({ S13758 })
);
AOI21_X1 #() 
AOI21_X1_927_ (
  .A({ S13465 }),
  .B1({ S13757 }),
  .B2({ S13758 }),
  .ZN({ S13759 })
);
OAI21_X1 #() 
OAI21_X1_851_ (
  .A({ S13391 }),
  .B1({ S13759 }),
  .B2({ S13751 }),
  .ZN({ S13760 })
);
NAND3_X1 #() 
NAND3_X1_1813_ (
  .A1({ S13717 }),
  .A2({ S25957[271] }),
  .A3({ S13711 }),
  .ZN({ S13761 })
);
NAND3_X1 #() 
NAND3_X1_1814_ (
  .A1({ S13747 }),
  .A2({ S13741 }),
  .A3({ S13465 }),
  .ZN({ S13762 })
);
NAND2_X1 #() 
NAND2_X1_1555_ (
  .A1({ S13761 }),
  .A2({ S13762 }),
  .ZN({ S13763 })
);
NAND2_X1 #() 
NAND2_X1_1556_ (
  .A1({ S13763 }),
  .A2({ S25957[270] }),
  .ZN({ S13764 })
);
NAND3_X1 #() 
NAND3_X1_1815_ (
  .A1({ S13764 }),
  .A2({ S13760 }),
  .A3({ S25957[372] }),
  .ZN({ S13765 })
);
AOI21_X1 #() 
AOI21_X1_928_ (
  .A({ S10811 }),
  .B1({ S13765 }),
  .B2({ S13750 }),
  .ZN({ S13767 })
);
NAND3_X1 #() 
NAND3_X1_1816_ (
  .A1({ S13749 }),
  .A2({ S13719 }),
  .A3({ S25957[372] }),
  .ZN({ S13768 })
);
NAND3_X1 #() 
NAND3_X1_1817_ (
  .A1({ S13764 }),
  .A2({ S13760 }),
  .A3({ S13689 }),
  .ZN({ S13769 })
);
AOI21_X1 #() 
AOI21_X1_929_ (
  .A({ S25957[436] }),
  .B1({ S13769 }),
  .B2({ S13768 }),
  .ZN({ S13770 })
);
OAI21_X1 #() 
OAI21_X1_852_ (
  .A({ S25957[276] }),
  .B1({ S13767 }),
  .B2({ S13770 }),
  .ZN({ S13771 })
);
NAND2_X1 #() 
NAND2_X1_1557_ (
  .A1({ S10899 }),
  .A2({ S10902 }),
  .ZN({ S13772 })
);
NAND3_X1 #() 
NAND3_X1_1818_ (
  .A1({ S13769 }),
  .A2({ S13768 }),
  .A3({ S25957[436] }),
  .ZN({ S13773 })
);
NAND3_X1 #() 
NAND3_X1_1819_ (
  .A1({ S13765 }),
  .A2({ S13750 }),
  .A3({ S10811 }),
  .ZN({ S13774 })
);
NAND3_X1 #() 
NAND3_X1_1820_ (
  .A1({ S13773 }),
  .A2({ S13774 }),
  .A3({ S13772 }),
  .ZN({ S13775 })
);
NAND2_X1 #() 
NAND2_X1_1558_ (
  .A1({ S13771 }),
  .A2({ S13775 }),
  .ZN({ S25957[148] })
);
NOR2_X1 #() 
NOR2_X1_351_ (
  .A1({ S10981 }),
  .A2({ S10984 }),
  .ZN({ S25957[307] })
);
INV_X1 #() 
INV_X1_491_ (
  .A({ S25957[307] }),
  .ZN({ S13777 })
);
NAND2_X1 #() 
NAND2_X1_1559_ (
  .A1({ S8055 }),
  .A2({ S8058 }),
  .ZN({ S25957[467] })
);
NAND2_X1 #() 
NAND2_X1_1560_ (
  .A1({ S10979 }),
  .A2({ S10954 }),
  .ZN({ S13778 })
);
XOR2_X1 #() 
XOR2_X1_25_ (
  .A({ S13778 }),
  .B({ S25957[467] }),
  .Z({ S13779 })
);
INV_X1 #() 
INV_X1_492_ (
  .A({ S13778 }),
  .ZN({ S25957[371] })
);
NAND3_X1 #() 
NAND3_X1_1821_ (
  .A1({ S13436 }),
  .A2({ S35 }),
  .A3({ S13401 }),
  .ZN({ S13780 })
);
AOI21_X1 #() 
AOI21_X1_930_ (
  .A({ S35 }),
  .B1({ S13402 }),
  .B2({ S13435 }),
  .ZN({ S13781 })
);
AOI21_X1 #() 
AOI21_X1_931_ (
  .A({ S25957[268] }),
  .B1({ S13781 }),
  .B2({ S13425 }),
  .ZN({ S13782 })
);
NAND2_X1 #() 
NAND2_X1_1561_ (
  .A1({ S13571 }),
  .A2({ S13661 }),
  .ZN({ S13783 })
);
AOI21_X1 #() 
AOI21_X1_932_ (
  .A({ S13412 }),
  .B1({ S13430 }),
  .B2({ S13600 }),
  .ZN({ S13785 })
);
AOI22_X1 #() 
AOI22_X1_214_ (
  .A1({ S13782 }),
  .A2({ S13780 }),
  .B1({ S13785 }),
  .B2({ S13783 }),
  .ZN({ S13786 })
);
NAND3_X1 #() 
NAND3_X1_1822_ (
  .A1({ S13422 }),
  .A2({ S25957[267] }),
  .A3({ S13416 }),
  .ZN({ S13787 })
);
NAND2_X1 #() 
NAND2_X1_1562_ (
  .A1({ S13713 }),
  .A2({ S35 }),
  .ZN({ S13788 })
);
NAND3_X1 #() 
NAND3_X1_1823_ (
  .A1({ S13788 }),
  .A2({ S13787 }),
  .A3({ S25957[268] }),
  .ZN({ S13789 })
);
NAND2_X1 #() 
NAND2_X1_1563_ (
  .A1({ S13585 }),
  .A2({ S35 }),
  .ZN({ S13790 })
);
NOR2_X1 #() 
NOR2_X1_352_ (
  .A1({ S13416 }),
  .A2({ S13418 }),
  .ZN({ S13791 })
);
AOI21_X1 #() 
AOI21_X1_933_ (
  .A({ S25957[265] }),
  .B1({ S25957[264] }),
  .B2({ S25957[266] }),
  .ZN({ S13792 })
);
OAI21_X1 #() 
OAI21_X1_853_ (
  .A({ S25957[267] }),
  .B1({ S13792 }),
  .B2({ S13791 }),
  .ZN({ S13793 })
);
NAND3_X1 #() 
NAND3_X1_1824_ (
  .A1({ S13793 }),
  .A2({ S13412 }),
  .A3({ S13790 }),
  .ZN({ S13794 })
);
NAND3_X1 #() 
NAND3_X1_1825_ (
  .A1({ S13794 }),
  .A2({ S13394 }),
  .A3({ S13789 }),
  .ZN({ S13796 })
);
OAI211_X1 #() 
OAI211_X1_591_ (
  .A({ S13796 }),
  .B({ S13391 }),
  .C1({ S13394 }),
  .C2({ S13786 }),
  .ZN({ S13797 })
);
NAND4_X1 #() 
NAND4_X1_231_ (
  .A1({ S13425 }),
  .A2({ S35 }),
  .A3({ S13402 }),
  .A4({ S13437 }),
  .ZN({ S13798 })
);
NAND2_X1 #() 
NAND2_X1_1564_ (
  .A1({ S25957[266] }),
  .A2({ S13437 }),
  .ZN({ S13799 })
);
NAND3_X1 #() 
NAND3_X1_1826_ (
  .A1({ S13668 }),
  .A2({ S25957[267] }),
  .A3({ S13799 }),
  .ZN({ S13800 })
);
AOI21_X1 #() 
AOI21_X1_934_ (
  .A({ S25957[268] }),
  .B1({ S13800 }),
  .B2({ S13798 }),
  .ZN({ S13801 })
);
OAI211_X1 #() 
OAI211_X1_592_ (
  .A({ S35 }),
  .B({ S13437 }),
  .C1({ S13435 }),
  .C2({ S25957[264] }),
  .ZN({ S13802 })
);
NAND3_X1 #() 
NAND3_X1_1827_ (
  .A1({ S13802 }),
  .A2({ S25957[268] }),
  .A3({ S13722 }),
  .ZN({ S13803 })
);
NAND2_X1 #() 
NAND2_X1_1565_ (
  .A1({ S13803 }),
  .A2({ S25957[269] }),
  .ZN({ S13804 })
);
NOR2_X1 #() 
NOR2_X1_353_ (
  .A1({ S13804 }),
  .A2({ S13801 }),
  .ZN({ S13805 })
);
NAND3_X1 #() 
NAND3_X1_1828_ (
  .A1({ S13632 }),
  .A2({ S35 }),
  .A3({ S13427 }),
  .ZN({ S13807 })
);
NAND2_X1 #() 
NAND2_X1_1566_ (
  .A1({ S13807 }),
  .A2({ S13674 }),
  .ZN({ S13808 })
);
NAND2_X1 #() 
NAND2_X1_1567_ (
  .A1({ S25957[266] }),
  .A2({ S25957[267] }),
  .ZN({ S13809 })
);
NAND4_X1 #() 
NAND4_X1_232_ (
  .A1({ S13809 }),
  .A2({ S13412 }),
  .A3({ S13547 }),
  .A4({ S43 }),
  .ZN({ S13810 })
);
NAND2_X1 #() 
NAND2_X1_1568_ (
  .A1({ S13810 }),
  .A2({ S13394 }),
  .ZN({ S13811 })
);
AOI21_X1 #() 
AOI21_X1_935_ (
  .A({ S13811 }),
  .B1({ S13808 }),
  .B2({ S25957[268] }),
  .ZN({ S13812 })
);
OAI21_X1 #() 
OAI21_X1_854_ (
  .A({ S25957[270] }),
  .B1({ S13805 }),
  .B2({ S13812 }),
  .ZN({ S13813 })
);
NAND3_X1 #() 
NAND3_X1_1829_ (
  .A1({ S13797 }),
  .A2({ S25957[271] }),
  .A3({ S13813 }),
  .ZN({ S13814 })
);
NAND3_X1 #() 
NAND3_X1_1830_ (
  .A1({ S13736 }),
  .A2({ S25957[267] }),
  .A3({ S13425 }),
  .ZN({ S13815 })
);
AOI21_X1 #() 
AOI21_X1_936_ (
  .A({ S25957[268] }),
  .B1({ S13489 }),
  .B2({ S13815 }),
  .ZN({ S13816 })
);
OAI211_X1 #() 
OAI211_X1_593_ (
  .A({ S43 }),
  .B({ S25957[267] }),
  .C1({ S25957[266] }),
  .C2({ S13418 }),
  .ZN({ S13818 })
);
AOI21_X1 #() 
AOI21_X1_937_ (
  .A({ S13412 }),
  .B1({ S13631 }),
  .B2({ S13818 }),
  .ZN({ S13819 })
);
OAI21_X1 #() 
OAI21_X1_855_ (
  .A({ S13394 }),
  .B1({ S13816 }),
  .B2({ S13819 }),
  .ZN({ S13820 })
);
NAND4_X1 #() 
NAND4_X1_233_ (
  .A1({ S13573 }),
  .A2({ S13396 }),
  .A3({ S25957[264] }),
  .A4({ S13412 }),
  .ZN({ S13821 })
);
AOI21_X1 #() 
AOI21_X1_938_ (
  .A({ S13571 }),
  .B1({ S13632 }),
  .B2({ S35 }),
  .ZN({ S13822 })
);
NAND2_X1 #() 
NAND2_X1_1569_ (
  .A1({ S13822 }),
  .A2({ S25957[268] }),
  .ZN({ S13823 })
);
NAND3_X1 #() 
NAND3_X1_1831_ (
  .A1({ S13823 }),
  .A2({ S25957[269] }),
  .A3({ S13821 }),
  .ZN({ S13824 })
);
NAND3_X1 #() 
NAND3_X1_1832_ (
  .A1({ S13820 }),
  .A2({ S13824 }),
  .A3({ S13391 }),
  .ZN({ S13825 })
);
NAND3_X1 #() 
NAND3_X1_1833_ (
  .A1({ S13396 }),
  .A2({ S35 }),
  .A3({ S13437 }),
  .ZN({ S13826 })
);
NAND3_X1 #() 
NAND3_X1_1834_ (
  .A1({ S13435 }),
  .A2({ S25957[267] }),
  .A3({ S13424 }),
  .ZN({ S13827 })
);
NAND3_X1 #() 
NAND3_X1_1835_ (
  .A1({ S13826 }),
  .A2({ S13827 }),
  .A3({ S13412 }),
  .ZN({ S13829 })
);
OAI211_X1 #() 
OAI211_X1_594_ (
  .A({ S25957[269] }),
  .B({ S13829 }),
  .C1({ S13480 }),
  .C2({ S13574 }),
  .ZN({ S13830 })
);
NAND3_X1 #() 
NAND3_X1_1836_ (
  .A1({ S13448 }),
  .A2({ S35 }),
  .A3({ S13418 }),
  .ZN({ S13831 })
);
NOR2_X1 #() 
NOR2_X1_354_ (
  .A1({ S13831 }),
  .A2({ S13412 }),
  .ZN({ S13832 })
);
AOI21_X1 #() 
AOI21_X1_939_ (
  .A({ S13832 }),
  .B1({ S13495 }),
  .B2({ S13727 }),
  .ZN({ S13833 })
);
OAI211_X1 #() 
OAI211_X1_595_ (
  .A({ S13830 }),
  .B({ S25957[270] }),
  .C1({ S13833 }),
  .C2({ S25957[269] }),
  .ZN({ S13834 })
);
NAND3_X1 #() 
NAND3_X1_1837_ (
  .A1({ S13825 }),
  .A2({ S13834 }),
  .A3({ S13465 }),
  .ZN({ S13835 })
);
NAND3_X1 #() 
NAND3_X1_1838_ (
  .A1({ S13814 }),
  .A2({ S25957[371] }),
  .A3({ S13835 }),
  .ZN({ S13836 })
);
NAND2_X1 #() 
NAND2_X1_1570_ (
  .A1({ S13800 }),
  .A2({ S13798 }),
  .ZN({ S13837 })
);
NAND2_X1 #() 
NAND2_X1_1571_ (
  .A1({ S13837 }),
  .A2({ S13412 }),
  .ZN({ S13838 })
);
NAND3_X1 #() 
NAND3_X1_1839_ (
  .A1({ S13838 }),
  .A2({ S25957[269] }),
  .A3({ S13803 }),
  .ZN({ S13840 })
);
AOI21_X1 #() 
AOI21_X1_940_ (
  .A({ S13675 }),
  .B1({ S13622 }),
  .B2({ S35 }),
  .ZN({ S13841 })
);
INV_X1 #() 
INV_X1_493_ (
  .A({ S13811 }),
  .ZN({ S13842 })
);
OAI21_X1 #() 
OAI21_X1_856_ (
  .A({ S13842 }),
  .B1({ S13841 }),
  .B2({ S13412 }),
  .ZN({ S13843 })
);
NAND3_X1 #() 
NAND3_X1_1840_ (
  .A1({ S13840 }),
  .A2({ S13843 }),
  .A3({ S25957[270] }),
  .ZN({ S13844 })
);
NAND4_X1 #() 
NAND4_X1_234_ (
  .A1({ S13425 }),
  .A2({ S13547 }),
  .A3({ S25957[267] }),
  .A4({ S25957[265] }),
  .ZN({ S13845 })
);
NAND3_X1 #() 
NAND3_X1_1841_ (
  .A1({ S13780 }),
  .A2({ S13412 }),
  .A3({ S13845 }),
  .ZN({ S13846 })
);
NAND2_X1 #() 
NAND2_X1_1572_ (
  .A1({ S13785 }),
  .A2({ S13783 }),
  .ZN({ S13847 })
);
NAND3_X1 #() 
NAND3_X1_1842_ (
  .A1({ S13847 }),
  .A2({ S13846 }),
  .A3({ S25957[269] }),
  .ZN({ S13848 })
);
NOR2_X1 #() 
NOR2_X1_355_ (
  .A1({ S13721 }),
  .A2({ S13397 }),
  .ZN({ S13849 })
);
NAND2_X1 #() 
NAND2_X1_1573_ (
  .A1({ S42 }),
  .A2({ S25957[266] }),
  .ZN({ S13851 })
);
NAND2_X1 #() 
NAND2_X1_1574_ (
  .A1({ S13448 }),
  .A2({ S13390 }),
  .ZN({ S13852 })
);
AOI21_X1 #() 
AOI21_X1_941_ (
  .A({ S35 }),
  .B1({ S13852 }),
  .B2({ S13851 }),
  .ZN({ S13853 })
);
OAI21_X1 #() 
OAI21_X1_857_ (
  .A({ S13412 }),
  .B1({ S13853 }),
  .B2({ S13849 }),
  .ZN({ S13854 })
);
NAND2_X1 #() 
NAND2_X1_1575_ (
  .A1({ S13438 }),
  .A2({ S25957[267] }),
  .ZN({ S13855 })
);
AOI21_X1 #() 
AOI21_X1_942_ (
  .A({ S13412 }),
  .B1({ S13550 }),
  .B2({ S13401 }),
  .ZN({ S13856 })
);
AOI21_X1 #() 
AOI21_X1_943_ (
  .A({ S25957[269] }),
  .B1({ S13856 }),
  .B2({ S13855 }),
  .ZN({ S13857 })
);
NAND2_X1 #() 
NAND2_X1_1576_ (
  .A1({ S13857 }),
  .A2({ S13854 }),
  .ZN({ S13858 })
);
NAND3_X1 #() 
NAND3_X1_1843_ (
  .A1({ S13858 }),
  .A2({ S13848 }),
  .A3({ S13391 }),
  .ZN({ S13859 })
);
NAND3_X1 #() 
NAND3_X1_1844_ (
  .A1({ S13844 }),
  .A2({ S13859 }),
  .A3({ S25957[271] }),
  .ZN({ S13860 })
);
AOI22_X1 #() 
AOI22_X1_215_ (
  .A1({ S13479 }),
  .A2({ S13436 }),
  .B1({ S13560 }),
  .B2({ S13600 }),
  .ZN({ S13862 })
);
AOI21_X1 #() 
AOI21_X1_944_ (
  .A({ S25957[267] }),
  .B1({ S43 }),
  .B2({ S13435 }),
  .ZN({ S13863 })
);
INV_X1 #() 
INV_X1_494_ (
  .A({ S13827 }),
  .ZN({ S13864 })
);
OAI21_X1 #() 
OAI21_X1_858_ (
  .A({ S13412 }),
  .B1({ S13864 }),
  .B2({ S13863 }),
  .ZN({ S13865 })
);
OAI211_X1 #() 
OAI211_X1_596_ (
  .A({ S13865 }),
  .B({ S25957[269] }),
  .C1({ S13862 }),
  .C2({ S13412 }),
  .ZN({ S13866 })
);
NAND2_X1 #() 
NAND2_X1_1577_ (
  .A1({ S13492 }),
  .A2({ S13448 }),
  .ZN({ S13867 })
);
AOI22_X1 #() 
AOI22_X1_216_ (
  .A1({ S13867 }),
  .A2({ S25957[267] }),
  .B1({ S13507 }),
  .B2({ S13492 }),
  .ZN({ S13868 })
);
AOI21_X1 #() 
AOI21_X1_945_ (
  .A({ S25957[267] }),
  .B1({ S13401 }),
  .B2({ S25957[264] }),
  .ZN({ S13869 })
);
AOI21_X1 #() 
AOI21_X1_946_ (
  .A({ S25957[269] }),
  .B1({ S25957[268] }),
  .B2({ S13869 }),
  .ZN({ S13870 })
);
OAI21_X1 #() 
OAI21_X1_859_ (
  .A({ S13870 }),
  .B1({ S13868 }),
  .B2({ S25957[268] }),
  .ZN({ S13871 })
);
NAND3_X1 #() 
NAND3_X1_1845_ (
  .A1({ S13866 }),
  .A2({ S13871 }),
  .A3({ S25957[270] }),
  .ZN({ S13873 })
);
AOI21_X1 #() 
AOI21_X1_947_ (
  .A({ S35 }),
  .B1({ S13426 }),
  .B2({ S25957[266] }),
  .ZN({ S13874 })
);
OAI21_X1 #() 
OAI21_X1_860_ (
  .A({ S25957[264] }),
  .B1({ S25957[266] }),
  .B2({ S13390 }),
  .ZN({ S13875 })
);
OAI21_X1 #() 
OAI21_X1_861_ (
  .A({ S13412 }),
  .B1({ S13874 }),
  .B2({ S13875 }),
  .ZN({ S13876 })
);
OAI211_X1 #() 
OAI211_X1_597_ (
  .A({ S25957[269] }),
  .B({ S13876 }),
  .C1({ S13822 }),
  .C2({ S13412 }),
  .ZN({ S13877 })
);
OAI21_X1 #() 
OAI21_X1_862_ (
  .A({ S43 }),
  .B1({ S25957[266] }),
  .B2({ S13418 }),
  .ZN({ S13878 })
);
AND2_X1 #() 
AND2_X1_96_ (
  .A1({ S13878 }),
  .A2({ S25957[267] }),
  .ZN({ S13879 })
);
NAND2_X1 #() 
NAND2_X1_1578_ (
  .A1({ S13557 }),
  .A2({ S25957[268] }),
  .ZN({ S13880 })
);
OAI21_X1 #() 
OAI21_X1_863_ (
  .A({ S13394 }),
  .B1({ S13879 }),
  .B2({ S13880 }),
  .ZN({ S13881 })
);
OAI211_X1 #() 
OAI211_X1_598_ (
  .A({ S13877 }),
  .B({ S13391 }),
  .C1({ S13816 }),
  .C2({ S13881 }),
  .ZN({ S13882 })
);
NAND3_X1 #() 
NAND3_X1_1846_ (
  .A1({ S13882 }),
  .A2({ S13873 }),
  .A3({ S13465 }),
  .ZN({ S13884 })
);
NAND3_X1 #() 
NAND3_X1_1847_ (
  .A1({ S13860 }),
  .A2({ S13884 }),
  .A3({ S13778 }),
  .ZN({ S13885 })
);
NAND3_X1 #() 
NAND3_X1_1848_ (
  .A1({ S13836 }),
  .A2({ S13885 }),
  .A3({ S13779 }),
  .ZN({ S13886 })
);
INV_X1 #() 
INV_X1_495_ (
  .A({ S13779 }),
  .ZN({ S25957[339] })
);
NAND3_X1 #() 
NAND3_X1_1849_ (
  .A1({ S13814 }),
  .A2({ S13778 }),
  .A3({ S13835 }),
  .ZN({ S13887 })
);
NAND3_X1 #() 
NAND3_X1_1850_ (
  .A1({ S13860 }),
  .A2({ S13884 }),
  .A3({ S25957[371] }),
  .ZN({ S13888 })
);
NAND3_X1 #() 
NAND3_X1_1851_ (
  .A1({ S13887 }),
  .A2({ S13888 }),
  .A3({ S25957[339] }),
  .ZN({ S13889 })
);
AOI21_X1 #() 
AOI21_X1_948_ (
  .A({ S13777 }),
  .B1({ S13886 }),
  .B2({ S13889 }),
  .ZN({ S13890 })
);
NAND3_X1 #() 
NAND3_X1_1852_ (
  .A1({ S13836 }),
  .A2({ S13885 }),
  .A3({ S25957[339] }),
  .ZN({ S13891 })
);
NAND3_X1 #() 
NAND3_X1_1853_ (
  .A1({ S13887 }),
  .A2({ S13888 }),
  .A3({ S13779 }),
  .ZN({ S13892 })
);
AOI21_X1 #() 
AOI21_X1_949_ (
  .A({ S25957[307] }),
  .B1({ S13891 }),
  .B2({ S13892 }),
  .ZN({ S13894 })
);
OAI21_X1 #() 
OAI21_X1_864_ (
  .A({ S32 }),
  .B1({ S13890 }),
  .B2({ S13894 }),
  .ZN({ S13895 })
);
NAND3_X1 #() 
NAND3_X1_1854_ (
  .A1({ S13891 }),
  .A2({ S13892 }),
  .A3({ S25957[307] }),
  .ZN({ S13896 })
);
NAND3_X1 #() 
NAND3_X1_1855_ (
  .A1({ S13886 }),
  .A2({ S13889 }),
  .A3({ S13777 }),
  .ZN({ S13897 })
);
NAND3_X1 #() 
NAND3_X1_1856_ (
  .A1({ S13896 }),
  .A2({ S13897 }),
  .A3({ S25957[275] }),
  .ZN({ S13898 })
);
NAND2_X1 #() 
NAND2_X1_1579_ (
  .A1({ S13895 }),
  .A2({ S13898 }),
  .ZN({ S44 })
);
OAI21_X1 #() 
OAI21_X1_865_ (
  .A({ S25957[275] }),
  .B1({ S13890 }),
  .B2({ S13894 }),
  .ZN({ S13899 })
);
NAND3_X1 #() 
NAND3_X1_1857_ (
  .A1({ S13896 }),
  .A2({ S13897 }),
  .A3({ S32 }),
  .ZN({ S13900 })
);
NAND2_X1 #() 
NAND2_X1_1580_ (
  .A1({ S13899 }),
  .A2({ S13900 }),
  .ZN({ S25957[147] })
);
NAND3_X1 #() 
NAND3_X1_1858_ (
  .A1({ S13592 }),
  .A2({ S13427 }),
  .A3({ S35 }),
  .ZN({ S13901 })
);
AOI21_X1 #() 
AOI21_X1_950_ (
  .A({ S25957[268] }),
  .B1({ S13867 }),
  .B2({ S25957[267] }),
  .ZN({ S13903 })
);
OAI22_X1 #() 
OAI22_X1_37_ (
  .A1({ S13720 }),
  .A2({ S13721 }),
  .B1({ S13543 }),
  .B2({ S35 }),
  .ZN({ S13904 })
);
AOI22_X1 #() 
AOI22_X1_217_ (
  .A1({ S13903 }),
  .A2({ S13901 }),
  .B1({ S13904 }),
  .B2({ S25957[268] }),
  .ZN({ S13905 })
);
OAI21_X1 #() 
OAI21_X1_866_ (
  .A({ S35 }),
  .B1({ S13443 }),
  .B2({ S13563 }),
  .ZN({ S13906 })
);
AOI21_X1 #() 
AOI21_X1_951_ (
  .A({ S13412 }),
  .B1({ S13422 }),
  .B2({ S13738 }),
  .ZN({ S13907 })
);
NAND2_X1 #() 
NAND2_X1_1581_ (
  .A1({ S13906 }),
  .A2({ S13907 }),
  .ZN({ S13908 })
);
NAND3_X1 #() 
NAND3_X1_1859_ (
  .A1({ S13486 }),
  .A2({ S13449 }),
  .A3({ S13547 }),
  .ZN({ S13909 })
);
AOI21_X1 #() 
AOI21_X1_952_ (
  .A({ S25957[269] }),
  .B1({ S13456 }),
  .B2({ S13909 }),
  .ZN({ S13910 })
);
NAND2_X1 #() 
NAND2_X1_1582_ (
  .A1({ S13908 }),
  .A2({ S13910 }),
  .ZN({ S13911 })
);
OAI211_X1 #() 
OAI211_X1_599_ (
  .A({ S13911 }),
  .B({ S25957[270] }),
  .C1({ S13905 }),
  .C2({ S13394 }),
  .ZN({ S13912 })
);
NAND3_X1 #() 
NAND3_X1_1860_ (
  .A1({ S13502 }),
  .A2({ S25957[268] }),
  .A3({ S13831 }),
  .ZN({ S13914 })
);
NAND4_X1 #() 
NAND4_X1_235_ (
  .A1({ S13707 }),
  .A2({ S13695 }),
  .A3({ S13644 }),
  .A4({ S13412 }),
  .ZN({ S13915 })
);
NAND3_X1 #() 
NAND3_X1_1861_ (
  .A1({ S13435 }),
  .A2({ S35 }),
  .A3({ S13424 }),
  .ZN({ S13916 })
);
OR2_X1 #() 
OR2_X1_24_ (
  .A1({ S13916 }),
  .A2({ S13412 }),
  .ZN({ S13917 })
);
NAND4_X1 #() 
NAND4_X1_236_ (
  .A1({ S13915 }),
  .A2({ S13914 }),
  .A3({ S13917 }),
  .A4({ S25957[269] }),
  .ZN({ S13918 })
);
OAI21_X1 #() 
OAI21_X1_867_ (
  .A({ S13536 }),
  .B1({ S13422 }),
  .B2({ S13537 }),
  .ZN({ S13919 })
);
NAND2_X1 #() 
NAND2_X1_1583_ (
  .A1({ S13919 }),
  .A2({ S25957[268] }),
  .ZN({ S13920 })
);
NAND4_X1 #() 
NAND4_X1_237_ (
  .A1({ S13455 }),
  .A2({ S13448 }),
  .A3({ S43 }),
  .A4({ S35 }),
  .ZN({ S13921 })
);
NAND3_X1 #() 
NAND3_X1_1862_ (
  .A1({ S13921 }),
  .A2({ S13412 }),
  .A3({ S13827 }),
  .ZN({ S13922 })
);
NAND3_X1 #() 
NAND3_X1_1863_ (
  .A1({ S13920 }),
  .A2({ S13394 }),
  .A3({ S13922 }),
  .ZN({ S13923 })
);
NAND3_X1 #() 
NAND3_X1_1864_ (
  .A1({ S13923 }),
  .A2({ S13918 }),
  .A3({ S13391 }),
  .ZN({ S13925 })
);
NAND3_X1 #() 
NAND3_X1_1865_ (
  .A1({ S13912 }),
  .A2({ S25957[271] }),
  .A3({ S13925 }),
  .ZN({ S13926 })
);
NAND3_X1 #() 
NAND3_X1_1866_ (
  .A1({ S13635 }),
  .A2({ S25957[268] }),
  .A3({ S13722 }),
  .ZN({ S13927 })
);
NAND3_X1 #() 
NAND3_X1_1867_ (
  .A1({ S13624 }),
  .A2({ S13412 }),
  .A3({ S13580 }),
  .ZN({ S13928 })
);
NAND3_X1 #() 
NAND3_X1_1868_ (
  .A1({ S13927 }),
  .A2({ S13928 }),
  .A3({ S25957[269] }),
  .ZN({ S13929 })
);
OAI21_X1 #() 
OAI21_X1_868_ (
  .A({ S35 }),
  .B1({ S13792 }),
  .B2({ S13791 }),
  .ZN({ S13930 })
);
AOI21_X1 #() 
AOI21_X1_953_ (
  .A({ S13412 }),
  .B1({ S13930 }),
  .B2({ S13855 }),
  .ZN({ S13931 })
);
NAND4_X1 #() 
NAND4_X1_238_ (
  .A1({ S13402 }),
  .A2({ S13396 }),
  .A3({ S25957[267] }),
  .A4({ S13437 }),
  .ZN({ S13932 })
);
NAND3_X1 #() 
NAND3_X1_1869_ (
  .A1({ S13413 }),
  .A2({ S35 }),
  .A3({ S13492 }),
  .ZN({ S13933 })
);
AOI21_X1 #() 
AOI21_X1_954_ (
  .A({ S25957[268] }),
  .B1({ S13933 }),
  .B2({ S13932 }),
  .ZN({ S13934 })
);
OAI21_X1 #() 
OAI21_X1_869_ (
  .A({ S13394 }),
  .B1({ S13931 }),
  .B2({ S13934 }),
  .ZN({ S13936 })
);
NAND3_X1 #() 
NAND3_X1_1870_ (
  .A1({ S13936 }),
  .A2({ S13391 }),
  .A3({ S13929 }),
  .ZN({ S13937 })
);
NAND4_X1 #() 
NAND4_X1_239_ (
  .A1({ S13851 }),
  .A2({ S13419 }),
  .A3({ S43 }),
  .A4({ S25957[267] }),
  .ZN({ S13938 })
);
AOI21_X1 #() 
AOI21_X1_955_ (
  .A({ S13412 }),
  .B1({ S13595 }),
  .B2({ S35 }),
  .ZN({ S13939 })
);
AOI22_X1 #() 
AOI22_X1_218_ (
  .A1({ S13564 }),
  .A2({ S13456 }),
  .B1({ S13938 }),
  .B2({ S13939 }),
  .ZN({ S13940 })
);
OAI211_X1 #() 
OAI211_X1_600_ (
  .A({ S13638 }),
  .B({ S13412 }),
  .C1({ S25957[267] }),
  .C2({ S13792 }),
  .ZN({ S13941 })
);
AOI21_X1 #() 
AOI21_X1_956_ (
  .A({ S13424 }),
  .B1({ S25957[266] }),
  .B2({ S13390 }),
  .ZN({ S13942 })
);
OAI211_X1 #() 
OAI211_X1_601_ (
  .A({ S35 }),
  .B({ S13435 }),
  .C1({ S13404 }),
  .C2({ S25957[266] }),
  .ZN({ S13943 })
);
OAI211_X1 #() 
OAI211_X1_602_ (
  .A({ S13943 }),
  .B({ S25957[268] }),
  .C1({ S35 }),
  .C2({ S13942 }),
  .ZN({ S13944 })
);
NAND3_X1 #() 
NAND3_X1_1871_ (
  .A1({ S13941 }),
  .A2({ S13394 }),
  .A3({ S13944 }),
  .ZN({ S13945 })
);
OAI211_X1 #() 
OAI211_X1_603_ (
  .A({ S13945 }),
  .B({ S25957[270] }),
  .C1({ S13940 }),
  .C2({ S13394 }),
  .ZN({ S13947 })
);
NAND3_X1 #() 
NAND3_X1_1872_ (
  .A1({ S13937 }),
  .A2({ S13947 }),
  .A3({ S13465 }),
  .ZN({ S13948 })
);
NAND3_X1 #() 
NAND3_X1_1873_ (
  .A1({ S13948 }),
  .A2({ S13926 }),
  .A3({ S10993 }),
  .ZN({ S13949 })
);
NAND3_X1 #() 
NAND3_X1_1874_ (
  .A1({ S13901 }),
  .A2({ S13429 }),
  .A3({ S13412 }),
  .ZN({ S13950 })
);
NAND2_X1 #() 
NAND2_X1_1584_ (
  .A1({ S13904 }),
  .A2({ S25957[268] }),
  .ZN({ S13951 })
);
AOI21_X1 #() 
AOI21_X1_957_ (
  .A({ S13394 }),
  .B1({ S13951 }),
  .B2({ S13950 }),
  .ZN({ S13952 })
);
AND2_X1 #() 
AND2_X1_97_ (
  .A1({ S13908 }),
  .A2({ S13910 }),
  .ZN({ S13953 })
);
OAI21_X1 #() 
OAI21_X1_870_ (
  .A({ S25957[270] }),
  .B1({ S13952 }),
  .B2({ S13953 }),
  .ZN({ S13954 })
);
NAND2_X1 #() 
NAND2_X1_1585_ (
  .A1({ S13923 }),
  .A2({ S13918 }),
  .ZN({ S13955 })
);
NAND2_X1 #() 
NAND2_X1_1586_ (
  .A1({ S13955 }),
  .A2({ S13391 }),
  .ZN({ S13956 })
);
NAND3_X1 #() 
NAND3_X1_1875_ (
  .A1({ S13954 }),
  .A2({ S25957[271] }),
  .A3({ S13956 }),
  .ZN({ S13958 })
);
AOI21_X1 #() 
AOI21_X1_958_ (
  .A({ S35 }),
  .B1({ S13422 }),
  .B2({ S13416 }),
  .ZN({ S13959 })
);
AOI21_X1 #() 
AOI21_X1_959_ (
  .A({ S25957[267] }),
  .B1({ S13852 }),
  .B2({ S13851 }),
  .ZN({ S13960 })
);
OAI21_X1 #() 
OAI21_X1_871_ (
  .A({ S25957[268] }),
  .B1({ S13960 }),
  .B2({ S13959 }),
  .ZN({ S13961 })
);
OAI21_X1 #() 
OAI21_X1_872_ (
  .A({ S35 }),
  .B1({ S13397 }),
  .B2({ S13416 }),
  .ZN({ S13962 })
);
OAI21_X1 #() 
OAI21_X1_873_ (
  .A({ S13932 }),
  .B1({ S13542 }),
  .B2({ S13962 }),
  .ZN({ S13963 })
);
NAND2_X1 #() 
NAND2_X1_1587_ (
  .A1({ S13963 }),
  .A2({ S13412 }),
  .ZN({ S13964 })
);
NAND3_X1 #() 
NAND3_X1_1876_ (
  .A1({ S13961 }),
  .A2({ S13964 }),
  .A3({ S13391 }),
  .ZN({ S13965 })
);
AOI22_X1 #() 
AOI22_X1_219_ (
  .A1({ S13476 }),
  .A2({ S13547 }),
  .B1({ S13852 }),
  .B2({ S35 }),
  .ZN({ S13966 })
);
NAND3_X1 #() 
NAND3_X1_1877_ (
  .A1({ S13529 }),
  .A2({ S35 }),
  .A3({ S13504 }),
  .ZN({ S13967 })
);
NAND2_X1 #() 
NAND2_X1_1588_ (
  .A1({ S13476 }),
  .A2({ S13455 }),
  .ZN({ S13969 })
);
NAND3_X1 #() 
NAND3_X1_1878_ (
  .A1({ S13969 }),
  .A2({ S25957[268] }),
  .A3({ S13967 }),
  .ZN({ S13970 })
);
OAI211_X1 #() 
OAI211_X1_604_ (
  .A({ S13970 }),
  .B({ S25957[270] }),
  .C1({ S25957[268] }),
  .C2({ S13966 }),
  .ZN({ S13971 })
);
AOI21_X1 #() 
AOI21_X1_960_ (
  .A({ S25957[269] }),
  .B1({ S13965 }),
  .B2({ S13971 }),
  .ZN({ S13972 })
);
NAND2_X1 #() 
NAND2_X1_1589_ (
  .A1({ S13927 }),
  .A2({ S13928 }),
  .ZN({ S13973 })
);
NAND2_X1 #() 
NAND2_X1_1590_ (
  .A1({ S13973 }),
  .A2({ S13391 }),
  .ZN({ S13974 })
);
NAND2_X1 #() 
NAND2_X1_1591_ (
  .A1({ S13938 }),
  .A2({ S13939 }),
  .ZN({ S13975 })
);
NAND2_X1 #() 
NAND2_X1_1592_ (
  .A1({ S13564 }),
  .A2({ S13456 }),
  .ZN({ S13976 })
);
NAND3_X1 #() 
NAND3_X1_1879_ (
  .A1({ S13976 }),
  .A2({ S25957[270] }),
  .A3({ S13975 }),
  .ZN({ S13977 })
);
AOI21_X1 #() 
AOI21_X1_961_ (
  .A({ S13394 }),
  .B1({ S13974 }),
  .B2({ S13977 }),
  .ZN({ S13978 })
);
OAI21_X1 #() 
OAI21_X1_874_ (
  .A({ S13465 }),
  .B1({ S13972 }),
  .B2({ S13978 }),
  .ZN({ S13980 })
);
NAND3_X1 #() 
NAND3_X1_1880_ (
  .A1({ S13980 }),
  .A2({ S13958 }),
  .A3({ S25957[464] }),
  .ZN({ S13981 })
);
AOI21_X1 #() 
AOI21_X1_962_ (
  .A({ S11081 }),
  .B1({ S13981 }),
  .B2({ S13949 }),
  .ZN({ S13982 })
);
AND3_X1 #() 
AND3_X1_74_ (
  .A1({ S13981 }),
  .A2({ S13949 }),
  .A3({ S11081 }),
  .ZN({ S13983 })
);
NOR2_X1 #() 
NOR2_X1_356_ (
  .A1({ S13983 }),
  .A2({ S13982 }),
  .ZN({ S25957[144] })
);
NAND2_X1 #() 
NAND2_X1_1593_ (
  .A1({ S8192 }),
  .A2({ S8178 }),
  .ZN({ S25957[497] })
);
XNOR2_X1 #() 
XNOR2_X1_54_ (
  .A({ S25957[497] }),
  .B({ S11087 }),
  .ZN({ S25957[465] })
);
INV_X1 #() 
INV_X1_496_ (
  .A({ S25957[465] }),
  .ZN({ S13984 })
);
NAND3_X1 #() 
NAND3_X1_1881_ (
  .A1({ S13508 }),
  .A2({ S25957[268] }),
  .A3({ S13674 }),
  .ZN({ S13985 })
);
NAND3_X1 #() 
NAND3_X1_1882_ (
  .A1({ S13938 }),
  .A2({ S13412 }),
  .A3({ S13499 }),
  .ZN({ S13986 })
);
NAND3_X1 #() 
NAND3_X1_1883_ (
  .A1({ S13986 }),
  .A2({ S25957[269] }),
  .A3({ S13985 }),
  .ZN({ S13988 })
);
NAND3_X1 #() 
NAND3_X1_1884_ (
  .A1({ S13633 }),
  .A2({ S25957[268] }),
  .A3({ S13916 }),
  .ZN({ S13989 })
);
NAND2_X1 #() 
NAND2_X1_1594_ (
  .A1({ S13869 }),
  .A2({ S13657 }),
  .ZN({ S13990 })
);
NAND3_X1 #() 
NAND3_X1_1885_ (
  .A1({ S13425 }),
  .A2({ S25957[267] }),
  .A3({ S13418 }),
  .ZN({ S13991 })
);
NAND3_X1 #() 
NAND3_X1_1886_ (
  .A1({ S13990 }),
  .A2({ S13412 }),
  .A3({ S13991 }),
  .ZN({ S13992 })
);
NAND3_X1 #() 
NAND3_X1_1887_ (
  .A1({ S13989 }),
  .A2({ S13992 }),
  .A3({ S13394 }),
  .ZN({ S13993 })
);
NAND3_X1 #() 
NAND3_X1_1888_ (
  .A1({ S13993 }),
  .A2({ S13988 }),
  .A3({ S25957[270] }),
  .ZN({ S13994 })
);
AOI21_X1 #() 
AOI21_X1_963_ (
  .A({ S25957[268] }),
  .B1({ S13700 }),
  .B2({ S35 }),
  .ZN({ S13995 })
);
NAND2_X1 #() 
NAND2_X1_1595_ (
  .A1({ S13995 }),
  .A2({ S13488 }),
  .ZN({ S13996 })
);
NOR2_X1 #() 
NOR2_X1_357_ (
  .A1({ S13396 }),
  .A2({ S35 }),
  .ZN({ S13997 })
);
NOR2_X1 #() 
NOR2_X1_358_ (
  .A1({ S13997 }),
  .A2({ S13412 }),
  .ZN({ S13999 })
);
AOI21_X1 #() 
AOI21_X1_964_ (
  .A({ S25957[269] }),
  .B1({ S13999 }),
  .B2({ S13967 }),
  .ZN({ S14000 })
);
NAND2_X1 #() 
NAND2_X1_1596_ (
  .A1({ S13996 }),
  .A2({ S14000 }),
  .ZN({ S14001 })
);
NAND3_X1 #() 
NAND3_X1_1889_ (
  .A1({ S13739 }),
  .A2({ S13695 }),
  .A3({ S13826 }),
  .ZN({ S14002 })
);
AOI21_X1 #() 
AOI21_X1_965_ (
  .A({ S35 }),
  .B1({ S13632 }),
  .B2({ S13455 }),
  .ZN({ S14003 })
);
OAI211_X1 #() 
OAI211_X1_605_ (
  .A({ S14002 }),
  .B({ S25957[269] }),
  .C1({ S13500 }),
  .C2({ S14003 }),
  .ZN({ S14004 })
);
NAND3_X1 #() 
NAND3_X1_1890_ (
  .A1({ S14001 }),
  .A2({ S13391 }),
  .A3({ S14004 }),
  .ZN({ S14005 })
);
NAND3_X1 #() 
NAND3_X1_1891_ (
  .A1({ S14005 }),
  .A2({ S25957[271] }),
  .A3({ S13994 }),
  .ZN({ S14006 })
);
AOI21_X1 #() 
AOI21_X1_966_ (
  .A({ S13412 }),
  .B1({ S13845 }),
  .B2({ S13709 }),
  .ZN({ S14007 })
);
OAI21_X1 #() 
OAI21_X1_875_ (
  .A({ S25957[269] }),
  .B1({ S14007 }),
  .B2({ S13495 }),
  .ZN({ S14008 })
);
AOI21_X1 #() 
AOI21_X1_967_ (
  .A({ S13642 }),
  .B1({ S13399 }),
  .B2({ S13537 }),
  .ZN({ S14010 })
);
NOR2_X1 #() 
NOR2_X1_359_ (
  .A1({ S13493 }),
  .A2({ S25957[267] }),
  .ZN({ S14011 })
);
OAI221_X1 #() 
OAI221_X1_32_ (
  .A({ S13394 }),
  .B1({ S13453 }),
  .B2({ S14010 }),
  .C1({ S14011 }),
  .C2({ S13446 }),
  .ZN({ S14012 })
);
NAND3_X1 #() 
NAND3_X1_1892_ (
  .A1({ S14012 }),
  .A2({ S14008 }),
  .A3({ S13391 }),
  .ZN({ S14013 })
);
OAI211_X1 #() 
OAI211_X1_606_ (
  .A({ S13586 }),
  .B({ S13412 }),
  .C1({ S13528 }),
  .C2({ S13809 }),
  .ZN({ S14014 })
);
NAND3_X1 #() 
NAND3_X1_1893_ (
  .A1({ S13851 }),
  .A2({ S13657 }),
  .A3({ S35 }),
  .ZN({ S14015 })
);
NAND3_X1 #() 
NAND3_X1_1894_ (
  .A1({ S13938 }),
  .A2({ S25957[268] }),
  .A3({ S14015 }),
  .ZN({ S14016 })
);
NAND3_X1 #() 
NAND3_X1_1895_ (
  .A1({ S14016 }),
  .A2({ S14014 }),
  .A3({ S13394 }),
  .ZN({ S14017 })
);
NAND3_X1 #() 
NAND3_X1_1896_ (
  .A1({ S13653 }),
  .A2({ S13448 }),
  .A3({ S13657 }),
  .ZN({ S14018 })
);
INV_X1 #() 
INV_X1_497_ (
  .A({ S13398 }),
  .ZN({ S14019 })
);
OAI21_X1 #() 
OAI21_X1_876_ (
  .A({ S25957[268] }),
  .B1({ S14019 }),
  .B2({ S13721 }),
  .ZN({ S14021 })
);
OAI211_X1 #() 
OAI211_X1_607_ (
  .A({ S25957[269] }),
  .B({ S14018 }),
  .C1({ S14021 }),
  .C2({ S13879 }),
  .ZN({ S14022 })
);
NAND3_X1 #() 
NAND3_X1_1897_ (
  .A1({ S14017 }),
  .A2({ S14022 }),
  .A3({ S25957[270] }),
  .ZN({ S14023 })
);
NAND3_X1 #() 
NAND3_X1_1898_ (
  .A1({ S14013 }),
  .A2({ S14023 }),
  .A3({ S13465 }),
  .ZN({ S14024 })
);
AND3_X1 #() 
AND3_X1_75_ (
  .A1({ S14006 }),
  .A2({ S14024 }),
  .A3({ S13984 }),
  .ZN({ S14025 })
);
AOI21_X1 #() 
AOI21_X1_968_ (
  .A({ S13984 }),
  .B1({ S14006 }),
  .B2({ S14024 }),
  .ZN({ S14026 })
);
OAI21_X1 #() 
OAI21_X1_877_ (
  .A({ S11179 }),
  .B1({ S14025 }),
  .B2({ S14026 }),
  .ZN({ S14027 })
);
NAND3_X1 #() 
NAND3_X1_1899_ (
  .A1({ S14006 }),
  .A2({ S14024 }),
  .A3({ S13984 }),
  .ZN({ S14028 })
);
NAND2_X1 #() 
NAND2_X1_1597_ (
  .A1({ S13989 }),
  .A2({ S13992 }),
  .ZN({ S14029 })
);
NAND2_X1 #() 
NAND2_X1_1598_ (
  .A1({ S14029 }),
  .A2({ S13394 }),
  .ZN({ S14030 })
);
OAI21_X1 #() 
OAI21_X1_878_ (
  .A({ S25957[268] }),
  .B1({ S13675 }),
  .B2({ S13507 }),
  .ZN({ S14032 })
);
INV_X1 #() 
INV_X1_498_ (
  .A({ S13499 }),
  .ZN({ S14033 })
);
AOI21_X1 #() 
AOI21_X1_969_ (
  .A({ S35 }),
  .B1({ S13436 }),
  .B2({ S13736 }),
  .ZN({ S14034 })
);
OAI21_X1 #() 
OAI21_X1_879_ (
  .A({ S13412 }),
  .B1({ S14034 }),
  .B2({ S14033 }),
  .ZN({ S14035 })
);
NAND3_X1 #() 
NAND3_X1_1900_ (
  .A1({ S14035 }),
  .A2({ S25957[269] }),
  .A3({ S14032 }),
  .ZN({ S14036 })
);
NAND3_X1 #() 
NAND3_X1_1901_ (
  .A1({ S14030 }),
  .A2({ S25957[270] }),
  .A3({ S14036 }),
  .ZN({ S14037 })
);
AOI22_X1 #() 
AOI22_X1_220_ (
  .A1({ S13995 }),
  .A2({ S13488 }),
  .B1({ S13967 }),
  .B2({ S13999 }),
  .ZN({ S14038 })
);
OAI21_X1 #() 
OAI21_X1_880_ (
  .A({ S13424 }),
  .B1({ S13416 }),
  .B2({ S25957[265] }),
  .ZN({ S14039 })
);
AOI21_X1 #() 
AOI21_X1_970_ (
  .A({ S35 }),
  .B1({ S25957[264] }),
  .B2({ S13416 }),
  .ZN({ S14040 })
);
AOI22_X1 #() 
AOI22_X1_221_ (
  .A1({ S14040 }),
  .A2({ S13436 }),
  .B1({ S14039 }),
  .B2({ S35 }),
  .ZN({ S14041 })
);
OAI21_X1 #() 
OAI21_X1_881_ (
  .A({ S13826 }),
  .B1({ S13563 }),
  .B2({ S35 }),
  .ZN({ S14043 })
);
NAND2_X1 #() 
NAND2_X1_1599_ (
  .A1({ S14043 }),
  .A2({ S13412 }),
  .ZN({ S14044 })
);
OAI211_X1 #() 
OAI211_X1_608_ (
  .A({ S14044 }),
  .B({ S25957[269] }),
  .C1({ S14041 }),
  .C2({ S13412 }),
  .ZN({ S14045 })
);
OAI211_X1 #() 
OAI211_X1_609_ (
  .A({ S14045 }),
  .B({ S13391 }),
  .C1({ S14038 }),
  .C2({ S25957[269] }),
  .ZN({ S14046 })
);
NAND3_X1 #() 
NAND3_X1_1902_ (
  .A1({ S14037 }),
  .A2({ S14046 }),
  .A3({ S25957[271] }),
  .ZN({ S14047 })
);
AOI22_X1 #() 
AOI22_X1_222_ (
  .A1({ S13878 }),
  .A2({ S25957[267] }),
  .B1({ S13441 }),
  .B2({ S13398 }),
  .ZN({ S14048 })
);
NAND3_X1 #() 
NAND3_X1_1903_ (
  .A1({ S13657 }),
  .A2({ S13452 }),
  .A3({ S13448 }),
  .ZN({ S14049 })
);
NAND2_X1 #() 
NAND2_X1_1600_ (
  .A1({ S14049 }),
  .A2({ S13412 }),
  .ZN({ S14050 })
);
OAI211_X1 #() 
OAI211_X1_610_ (
  .A({ S14050 }),
  .B({ S25957[269] }),
  .C1({ S14048 }),
  .C2({ S13412 }),
  .ZN({ S14051 })
);
NAND2_X1 #() 
NAND2_X1_1601_ (
  .A1({ S43 }),
  .A2({ S13416 }),
  .ZN({ S14052 })
);
AOI21_X1 #() 
AOI21_X1_971_ (
  .A({ S25957[267] }),
  .B1({ S14052 }),
  .B2({ S13486 }),
  .ZN({ S14054 })
);
OAI21_X1 #() 
OAI21_X1_882_ (
  .A({ S25957[268] }),
  .B1({ S14034 }),
  .B2({ S14054 }),
  .ZN({ S14055 })
);
OAI21_X1 #() 
OAI21_X1_883_ (
  .A({ S13586 }),
  .B1({ S35 }),
  .B2({ S13632 }),
  .ZN({ S14056 })
);
NAND2_X1 #() 
NAND2_X1_1602_ (
  .A1({ S14056 }),
  .A2({ S13412 }),
  .ZN({ S14057 })
);
NAND3_X1 #() 
NAND3_X1_1904_ (
  .A1({ S14055 }),
  .A2({ S14057 }),
  .A3({ S13394 }),
  .ZN({ S14058 })
);
NAND3_X1 #() 
NAND3_X1_1905_ (
  .A1({ S14058 }),
  .A2({ S25957[270] }),
  .A3({ S14051 }),
  .ZN({ S14059 })
);
INV_X1 #() 
INV_X1_499_ (
  .A({ S13495 }),
  .ZN({ S14060 })
);
INV_X1 #() 
INV_X1_500_ (
  .A({ S14007 }),
  .ZN({ S14061 })
);
NAND3_X1 #() 
NAND3_X1_1906_ (
  .A1({ S14061 }),
  .A2({ S14060 }),
  .A3({ S25957[269] }),
  .ZN({ S14062 })
);
NOR2_X1 #() 
NOR2_X1_360_ (
  .A1({ S13453 }),
  .A2({ S14010 }),
  .ZN({ S14063 })
);
AOI21_X1 #() 
AOI21_X1_972_ (
  .A({ S13446 }),
  .B1({ S13492 }),
  .B2({ S13507 }),
  .ZN({ S14065 })
);
OAI21_X1 #() 
OAI21_X1_884_ (
  .A({ S13394 }),
  .B1({ S14065 }),
  .B2({ S14063 }),
  .ZN({ S14066 })
);
NAND3_X1 #() 
NAND3_X1_1907_ (
  .A1({ S14062 }),
  .A2({ S14066 }),
  .A3({ S13391 }),
  .ZN({ S14067 })
);
NAND3_X1 #() 
NAND3_X1_1908_ (
  .A1({ S14059 }),
  .A2({ S13465 }),
  .A3({ S14067 }),
  .ZN({ S14068 })
);
NAND3_X1 #() 
NAND3_X1_1909_ (
  .A1({ S14047 }),
  .A2({ S14068 }),
  .A3({ S25957[465] }),
  .ZN({ S14069 })
);
NAND3_X1 #() 
NAND3_X1_1910_ (
  .A1({ S14069 }),
  .A2({ S25957[401] }),
  .A3({ S14028 }),
  .ZN({ S14070 })
);
NAND2_X1 #() 
NAND2_X1_1603_ (
  .A1({ S14027 }),
  .A2({ S14070 }),
  .ZN({ S25957[145] })
);
NOR2_X1 #() 
NOR2_X1_361_ (
  .A1({ S8284 }),
  .A2({ S8285 }),
  .ZN({ S25957[466] })
);
NAND3_X1 #() 
NAND3_X1_1911_ (
  .A1({ S13564 }),
  .A2({ S13412 }),
  .A3({ S13901 }),
  .ZN({ S14071 })
);
NAND3_X1 #() 
NAND3_X1_1912_ (
  .A1({ S13547 }),
  .A2({ S25957[267] }),
  .A3({ S25957[265] }),
  .ZN({ S14072 })
);
OAI211_X1 #() 
OAI211_X1_611_ (
  .A({ S25957[268] }),
  .B({ S14072 }),
  .C1({ S13499 }),
  .C2({ S13501 }),
  .ZN({ S14074 })
);
NAND3_X1 #() 
NAND3_X1_1913_ (
  .A1({ S14071 }),
  .A2({ S13394 }),
  .A3({ S14074 }),
  .ZN({ S14075 })
);
OAI211_X1 #() 
OAI211_X1_612_ (
  .A({ S13539 }),
  .B({ S13412 }),
  .C1({ S13619 }),
  .C2({ S13791 }),
  .ZN({ S14076 })
);
NAND2_X1 #() 
NAND2_X1_1604_ (
  .A1({ S13471 }),
  .A2({ S13657 }),
  .ZN({ S14077 })
);
NAND3_X1 #() 
NAND3_X1_1914_ (
  .A1({ S13780 }),
  .A2({ S14077 }),
  .A3({ S25957[268] }),
  .ZN({ S14078 })
);
NAND3_X1 #() 
NAND3_X1_1915_ (
  .A1({ S14078 }),
  .A2({ S14076 }),
  .A3({ S25957[269] }),
  .ZN({ S14079 })
);
NAND2_X1 #() 
NAND2_X1_1605_ (
  .A1({ S14075 }),
  .A2({ S14079 }),
  .ZN({ S14080 })
);
NAND2_X1 #() 
NAND2_X1_1606_ (
  .A1({ S14080 }),
  .A2({ S13391 }),
  .ZN({ S14081 })
);
OAI21_X1 #() 
OAI21_X1_885_ (
  .A({ S13412 }),
  .B1({ S13531 }),
  .B2({ S13424 }),
  .ZN({ S14082 })
);
NOR3_X1 #() 
NOR3_X1_55_ (
  .A1({ S13642 }),
  .A2({ S13426 }),
  .A3({ S35 }),
  .ZN({ S14083 })
);
OAI21_X1 #() 
OAI21_X1_886_ (
  .A({ S25957[268] }),
  .B1({ S14083 }),
  .B2({ S13869 }),
  .ZN({ S14085 })
);
OAI211_X1 #() 
OAI211_X1_613_ (
  .A({ S14085 }),
  .B({ S25957[269] }),
  .C1({ S13440 }),
  .C2({ S14082 }),
  .ZN({ S14086 })
);
NAND2_X1 #() 
NAND2_X1_1607_ (
  .A1({ S13419 }),
  .A2({ S13799 }),
  .ZN({ S14087 })
);
AOI22_X1 #() 
AOI22_X1_223_ (
  .A1({ S14087 }),
  .A2({ S35 }),
  .B1({ S13471 }),
  .B2({ S13529 }),
  .ZN({ S14088 })
);
NAND3_X1 #() 
NAND3_X1_1916_ (
  .A1({ S13668 }),
  .A2({ S35 }),
  .A3({ S13799 }),
  .ZN({ S14089 })
);
NAND3_X1 #() 
NAND3_X1_1917_ (
  .A1({ S14089 }),
  .A2({ S13412 }),
  .A3({ S14072 }),
  .ZN({ S14090 })
);
OAI211_X1 #() 
OAI211_X1_614_ (
  .A({ S14090 }),
  .B({ S13394 }),
  .C1({ S14088 }),
  .C2({ S13412 }),
  .ZN({ S14091 })
);
NAND3_X1 #() 
NAND3_X1_1918_ (
  .A1({ S14091 }),
  .A2({ S14086 }),
  .A3({ S25957[270] }),
  .ZN({ S14092 })
);
NAND3_X1 #() 
NAND3_X1_1919_ (
  .A1({ S14081 }),
  .A2({ S13465 }),
  .A3({ S14092 }),
  .ZN({ S14093 })
);
AOI22_X1 #() 
AOI22_X1_224_ (
  .A1({ S13469 }),
  .A2({ S13448 }),
  .B1({ S13874 }),
  .B2({ S13402 }),
  .ZN({ S14094 })
);
NAND2_X1 #() 
NAND2_X1_1608_ (
  .A1({ S13493 }),
  .A2({ S35 }),
  .ZN({ S14096 })
);
AOI21_X1 #() 
AOI21_X1_973_ (
  .A({ S13412 }),
  .B1({ S13726 }),
  .B2({ S25957[267] }),
  .ZN({ S14097 })
);
NAND2_X1 #() 
NAND2_X1_1609_ (
  .A1({ S14096 }),
  .A2({ S14097 }),
  .ZN({ S14098 })
);
OAI21_X1 #() 
OAI21_X1_887_ (
  .A({ S14098 }),
  .B1({ S14094 }),
  .B2({ S25957[268] }),
  .ZN({ S14099 })
);
NAND3_X1 #() 
NAND3_X1_1920_ (
  .A1({ S14072 }),
  .A2({ S25957[268] }),
  .A3({ S13531 }),
  .ZN({ S14100 })
);
OAI211_X1 #() 
OAI211_X1_615_ (
  .A({ S13536 }),
  .B({ S13412 }),
  .C1({ S13455 }),
  .C2({ S13449 }),
  .ZN({ S14101 })
);
NAND2_X1 #() 
NAND2_X1_1610_ (
  .A1({ S14100 }),
  .A2({ S14101 }),
  .ZN({ S14102 })
);
AOI21_X1 #() 
AOI21_X1_974_ (
  .A({ S25957[270] }),
  .B1({ S14102 }),
  .B2({ S13394 }),
  .ZN({ S14103 })
);
OAI21_X1 #() 
OAI21_X1_888_ (
  .A({ S14103 }),
  .B1({ S14099 }),
  .B2({ S13394 }),
  .ZN({ S14104 })
);
NAND3_X1 #() 
NAND3_X1_1921_ (
  .A1({ S13661 }),
  .A2({ S25957[267] }),
  .A3({ S13799 }),
  .ZN({ S14105 })
);
NAND3_X1 #() 
NAND3_X1_1922_ (
  .A1({ S14105 }),
  .A2({ S13663 }),
  .A3({ S25957[268] }),
  .ZN({ S14107 })
);
OAI211_X1 #() 
OAI211_X1_616_ (
  .A({ S13466 }),
  .B({ S13412 }),
  .C1({ S25957[267] }),
  .C2({ S13401 }),
  .ZN({ S14108 })
);
AND2_X1 #() 
AND2_X1_98_ (
  .A1({ S14108 }),
  .A2({ S13394 }),
  .ZN({ S14109 })
);
AND2_X1 #() 
AND2_X1_99_ (
  .A1({ S13592 }),
  .A2({ S13427 }),
  .ZN({ S14110 })
);
OAI211_X1 #() 
OAI211_X1_617_ (
  .A({ S25957[268] }),
  .B({ S13491 }),
  .C1({ S14110 }),
  .C2({ S25957[267] }),
  .ZN({ S14111 })
);
NAND3_X1 #() 
NAND3_X1_1923_ (
  .A1({ S13661 }),
  .A2({ S25957[267] }),
  .A3({ S13543 }),
  .ZN({ S14112 })
);
NOR2_X1 #() 
NOR2_X1_362_ (
  .A1({ S13469 }),
  .A2({ S25957[268] }),
  .ZN({ S14113 })
);
AOI21_X1 #() 
AOI21_X1_975_ (
  .A({ S13394 }),
  .B1({ S14113 }),
  .B2({ S14112 }),
  .ZN({ S14114 })
);
AOI22_X1 #() 
AOI22_X1_225_ (
  .A1({ S14111 }),
  .A2({ S14114 }),
  .B1({ S14109 }),
  .B2({ S14107 }),
  .ZN({ S14115 })
);
OAI211_X1 #() 
OAI211_X1_618_ (
  .A({ S14104 }),
  .B({ S25957[271] }),
  .C1({ S14115 }),
  .C2({ S13391 }),
  .ZN({ S14116 })
);
NAND3_X1 #() 
NAND3_X1_1924_ (
  .A1({ S14093 }),
  .A2({ S14116 }),
  .A3({ S25957[466] }),
  .ZN({ S14118 })
);
INV_X1 #() 
INV_X1_501_ (
  .A({ S25957[466] }),
  .ZN({ S14119 })
);
NAND3_X1 #() 
NAND3_X1_1925_ (
  .A1({ S14100 }),
  .A2({ S14101 }),
  .A3({ S13394 }),
  .ZN({ S14120 })
);
NAND2_X1 #() 
NAND2_X1_1611_ (
  .A1({ S13507 }),
  .A2({ S13492 }),
  .ZN({ S14121 })
);
OAI211_X1 #() 
OAI211_X1_619_ (
  .A({ S14121 }),
  .B({ S25957[268] }),
  .C1({ S35 }),
  .C2({ S13726 }),
  .ZN({ S14122 })
);
OAI211_X1 #() 
OAI211_X1_620_ (
  .A({ S13962 }),
  .B({ S13412 }),
  .C1({ S13573 }),
  .C2({ S13404 }),
  .ZN({ S14123 })
);
NAND3_X1 #() 
NAND3_X1_1926_ (
  .A1({ S14122 }),
  .A2({ S25957[269] }),
  .A3({ S14123 }),
  .ZN({ S14124 })
);
AOI21_X1 #() 
AOI21_X1_976_ (
  .A({ S25957[270] }),
  .B1({ S14124 }),
  .B2({ S14120 }),
  .ZN({ S14125 })
);
NAND2_X1 #() 
NAND2_X1_1612_ (
  .A1({ S14109 }),
  .A2({ S14107 }),
  .ZN({ S14126 })
);
NAND2_X1 #() 
NAND2_X1_1613_ (
  .A1({ S14111 }),
  .A2({ S14114 }),
  .ZN({ S14127 })
);
AOI21_X1 #() 
AOI21_X1_977_ (
  .A({ S13391 }),
  .B1({ S14127 }),
  .B2({ S14126 }),
  .ZN({ S14129 })
);
OAI21_X1 #() 
OAI21_X1_889_ (
  .A({ S25957[271] }),
  .B1({ S14129 }),
  .B2({ S14125 }),
  .ZN({ S14130 })
);
AOI21_X1 #() 
AOI21_X1_978_ (
  .A({ S25957[270] }),
  .B1({ S14075 }),
  .B2({ S14079 }),
  .ZN({ S14131 })
);
AND3_X1 #() 
AND3_X1_76_ (
  .A1({ S14091 }),
  .A2({ S14086 }),
  .A3({ S25957[270] }),
  .ZN({ S14132 })
);
OAI21_X1 #() 
OAI21_X1_890_ (
  .A({ S13465 }),
  .B1({ S14132 }),
  .B2({ S14131 }),
  .ZN({ S14133 })
);
NAND3_X1 #() 
NAND3_X1_1927_ (
  .A1({ S14133 }),
  .A2({ S14130 }),
  .A3({ S14119 }),
  .ZN({ S14134 })
);
AOI21_X1 #() 
AOI21_X1_979_ (
  .A({ S11281 }),
  .B1({ S14134 }),
  .B2({ S14118 }),
  .ZN({ S14135 })
);
AND3_X1 #() 
AND3_X1_77_ (
  .A1({ S14134 }),
  .A2({ S14118 }),
  .A3({ S11281 }),
  .ZN({ S14136 })
);
NOR2_X1 #() 
NOR2_X1_363_ (
  .A1({ S14136 }),
  .A2({ S14135 }),
  .ZN({ S25957[146] })
);
NAND3_X1 #() 
NAND3_X1_1928_ (
  .A1({ S12515 }),
  .A2({ S12516 }),
  .A3({ S11300 }),
  .ZN({ S14137 })
);
NAND3_X1 #() 
NAND3_X1_1929_ (
  .A1({ S12508 }),
  .A2({ S12513 }),
  .A3({ S25957[384] }),
  .ZN({ S14139 })
);
NAND3_X1 #() 
NAND3_X1_1930_ (
  .A1({ S25957[257] }),
  .A2({ S14137 }),
  .A3({ S14139 }),
  .ZN({ S14140 })
);
INV_X1 #() 
INV_X1_502_ (
  .A({ S14140 }),
  .ZN({ S45 })
);
NAND2_X1 #() 
NAND2_X1_1614_ (
  .A1({ S12575 }),
  .A2({ S12578 }),
  .ZN({ S14141 })
);
NAND3_X1 #() 
NAND3_X1_1931_ (
  .A1({ S12514 }),
  .A2({ S12517 }),
  .A3({ S14141 }),
  .ZN({ S46 })
);
NOR2_X1 #() 
NOR2_X1_364_ (
  .A1({ S8423 }),
  .A2({ S8422 }),
  .ZN({ S25957[431] })
);
INV_X1 #() 
INV_X1_503_ (
  .A({ S25957[262] }),
  .ZN({ S14142 })
);
OAI21_X1 #() 
OAI21_X1_891_ (
  .A({ S11332 }),
  .B1({ S12352 }),
  .B2({ S12355 }),
  .ZN({ S14143 })
);
NAND3_X1 #() 
NAND3_X1_1932_ (
  .A1({ S12359 }),
  .A2({ S25957[388] }),
  .A3({ S12358 }),
  .ZN({ S14144 })
);
NAND2_X1 #() 
NAND2_X1_1615_ (
  .A1({ S14144 }),
  .A2({ S14143 }),
  .ZN({ S14145 })
);
NAND4_X1 #() 
NAND4_X1_240_ (
  .A1({ S12514 }),
  .A2({ S12517 }),
  .A3({ S12672 }),
  .A4({ S12675 }),
  .ZN({ S14147 })
);
NAND3_X1 #() 
NAND3_X1_1933_ (
  .A1({ S12673 }),
  .A2({ S12674 }),
  .A3({ S11298 }),
  .ZN({ S14148 })
);
NAND3_X1 #() 
NAND3_X1_1934_ (
  .A1({ S12667 }),
  .A2({ S12671 }),
  .A3({ S25957[386] }),
  .ZN({ S14149 })
);
NAND4_X1 #() 
NAND4_X1_241_ (
  .A1({ S14137 }),
  .A2({ S14139 }),
  .A3({ S14148 }),
  .A4({ S14149 }),
  .ZN({ S14150 })
);
NAND3_X1 #() 
NAND3_X1_1935_ (
  .A1({ S25957[257] }),
  .A2({ S12672 }),
  .A3({ S12675 }),
  .ZN({ S14151 })
);
NAND3_X1 #() 
NAND3_X1_1936_ (
  .A1({ S14147 }),
  .A2({ S14150 }),
  .A3({ S14151 }),
  .ZN({ S14152 })
);
NAND2_X1 #() 
NAND2_X1_1616_ (
  .A1({ S14152 }),
  .A2({ S25957[259] }),
  .ZN({ S14153 })
);
NAND2_X1 #() 
NAND2_X1_1617_ (
  .A1({ S14148 }),
  .A2({ S14149 }),
  .ZN({ S14154 })
);
NAND2_X1 #() 
NAND2_X1_1618_ (
  .A1({ S14140 }),
  .A2({ S14154 }),
  .ZN({ S14155 })
);
NAND3_X1 #() 
NAND3_X1_1937_ (
  .A1({ S25957[257] }),
  .A2({ S12514 }),
  .A3({ S12517 }),
  .ZN({ S14156 })
);
NAND3_X1 #() 
NAND3_X1_1938_ (
  .A1({ S14137 }),
  .A2({ S14139 }),
  .A3({ S14141 }),
  .ZN({ S14158 })
);
NAND2_X1 #() 
NAND2_X1_1619_ (
  .A1({ S14156 }),
  .A2({ S14158 }),
  .ZN({ S14159 })
);
AOI21_X1 #() 
AOI21_X1_980_ (
  .A({ S14141 }),
  .B1({ S14148 }),
  .B2({ S14149 }),
  .ZN({ S14160 })
);
NOR2_X1 #() 
NOR2_X1_365_ (
  .A1({ S14160 }),
  .A2({ S38 }),
  .ZN({ S14161 })
);
NAND3_X1 #() 
NAND3_X1_1939_ (
  .A1({ S25957[257] }),
  .A2({ S14148 }),
  .A3({ S14149 }),
  .ZN({ S14162 })
);
NAND3_X1 #() 
NAND3_X1_1940_ (
  .A1({ S14150 }),
  .A2({ S14162 }),
  .A3({ S38 }),
  .ZN({ S14163 })
);
INV_X1 #() 
INV_X1_504_ (
  .A({ S14163 }),
  .ZN({ S14164 })
);
AOI22_X1 #() 
AOI22_X1_226_ (
  .A1({ S14164 }),
  .A2({ S14155 }),
  .B1({ S14159 }),
  .B2({ S14161 }),
  .ZN({ S14165 })
);
NAND2_X1 #() 
NAND2_X1_1620_ (
  .A1({ S14147 }),
  .A2({ S25957[257] }),
  .ZN({ S14166 })
);
INV_X1 #() 
INV_X1_505_ (
  .A({ S14166 }),
  .ZN({ S14167 })
);
AOI21_X1 #() 
AOI21_X1_981_ (
  .A({ S14145 }),
  .B1({ S14167 }),
  .B2({ S38 }),
  .ZN({ S14169 })
);
AOI22_X1 #() 
AOI22_X1_227_ (
  .A1({ S14165 }),
  .A2({ S14145 }),
  .B1({ S14169 }),
  .B2({ S14153 }),
  .ZN({ S14170 })
);
NAND2_X1 #() 
NAND2_X1_1621_ (
  .A1({ S14156 }),
  .A2({ S38 }),
  .ZN({ S14171 })
);
INV_X1 #() 
INV_X1_506_ (
  .A({ S14171 }),
  .ZN({ S14172 })
);
NAND3_X1 #() 
NAND3_X1_1941_ (
  .A1({ S12672 }),
  .A2({ S12675 }),
  .A3({ S14141 }),
  .ZN({ S14173 })
);
AOI21_X1 #() 
AOI21_X1_982_ (
  .A({ S38 }),
  .B1({ S14156 }),
  .B2({ S14173 }),
  .ZN({ S14174 })
);
OAI21_X1 #() 
OAI21_X1_892_ (
  .A({ S25957[260] }),
  .B1({ S14172 }),
  .B2({ S14174 }),
  .ZN({ S14175 })
);
NAND3_X1 #() 
NAND3_X1_1942_ (
  .A1({ S14148 }),
  .A2({ S14149 }),
  .A3({ S14141 }),
  .ZN({ S14176 })
);
OAI21_X1 #() 
OAI21_X1_893_ (
  .A({ S25957[259] }),
  .B1({ S14176 }),
  .B2({ S25957[256] }),
  .ZN({ S14177 })
);
NAND4_X1 #() 
NAND4_X1_242_ (
  .A1({ S14137 }),
  .A2({ S14139 }),
  .A3({ S12672 }),
  .A4({ S12675 }),
  .ZN({ S14178 })
);
NAND2_X1 #() 
NAND2_X1_1622_ (
  .A1({ S14178 }),
  .A2({ S14151 }),
  .ZN({ S14180 })
);
OAI21_X1 #() 
OAI21_X1_894_ (
  .A({ S38 }),
  .B1({ S14176 }),
  .B2({ S25957[256] }),
  .ZN({ S14181 })
);
OAI221_X1 #() 
OAI221_X1_33_ (
  .A({ S14145 }),
  .B1({ S14177 }),
  .B2({ S14160 }),
  .C1({ S14180 }),
  .C2({ S14181 }),
  .ZN({ S14182 })
);
AOI21_X1 #() 
AOI21_X1_983_ (
  .A({ S25957[261] }),
  .B1({ S14182 }),
  .B2({ S14175 }),
  .ZN({ S14183 })
);
AOI21_X1 #() 
AOI21_X1_984_ (
  .A({ S14183 }),
  .B1({ S14170 }),
  .B2({ S25957[261] }),
  .ZN({ S14184 })
);
NOR2_X1 #() 
NOR2_X1_366_ (
  .A1({ S14184 }),
  .A2({ S14142 }),
  .ZN({ S14185 })
);
INV_X1 #() 
INV_X1_507_ (
  .A({ S25957[261] }),
  .ZN({ S14186 })
);
NAND3_X1 #() 
NAND3_X1_1943_ (
  .A1({ S14156 }),
  .A2({ S14158 }),
  .A3({ S14154 }),
  .ZN({ S14187 })
);
NAND3_X1 #() 
NAND3_X1_1944_ (
  .A1({ S25957[256] }),
  .A2({ S25957[258] }),
  .A3({ S14141 }),
  .ZN({ S14188 })
);
AOI21_X1 #() 
AOI21_X1_985_ (
  .A({ S25957[259] }),
  .B1({ S14187 }),
  .B2({ S14188 }),
  .ZN({ S14189 })
);
NAND2_X1 #() 
NAND2_X1_1623_ (
  .A1({ S25957[259] }),
  .A2({ S14141 }),
  .ZN({ S14191 })
);
NOR2_X1 #() 
NOR2_X1_367_ (
  .A1({ S14191 }),
  .A2({ S25957[258] }),
  .ZN({ S14192 })
);
NOR3_X1 #() 
NOR3_X1_56_ (
  .A1({ S14189 }),
  .A2({ S14192 }),
  .A3({ S25957[260] }),
  .ZN({ S14193 })
);
NAND2_X1 #() 
NAND2_X1_1624_ (
  .A1({ S14147 }),
  .A2({ S38 }),
  .ZN({ S14194 })
);
INV_X1 #() 
INV_X1_508_ (
  .A({ S14194 }),
  .ZN({ S14195 })
);
NAND2_X1 #() 
NAND2_X1_1625_ (
  .A1({ S14137 }),
  .A2({ S14139 }),
  .ZN({ S14196 })
);
NAND3_X1 #() 
NAND3_X1_1945_ (
  .A1({ S14196 }),
  .A2({ S25957[258] }),
  .A3({ S25957[257] }),
  .ZN({ S14197 })
);
NAND4_X1 #() 
NAND4_X1_243_ (
  .A1({ S14187 }),
  .A2({ S14188 }),
  .A3({ S25957[259] }),
  .A4({ S14197 }),
  .ZN({ S14198 })
);
INV_X1 #() 
INV_X1_509_ (
  .A({ S14198 }),
  .ZN({ S14199 })
);
AOI211_X1 #() 
AOI211_X1_20_ (
  .A({ S14145 }),
  .B({ S14199 }),
  .C1({ S14176 }),
  .C2({ S14195 }),
  .ZN({ S14200 })
);
OAI21_X1 #() 
OAI21_X1_895_ (
  .A({ S14186 }),
  .B1({ S14200 }),
  .B2({ S14193 }),
  .ZN({ S14202 })
);
AOI21_X1 #() 
AOI21_X1_986_ (
  .A({ S38 }),
  .B1({ S14150 }),
  .B2({ S25957[257] }),
  .ZN({ S14203 })
);
INV_X1 #() 
INV_X1_510_ (
  .A({ S14150 }),
  .ZN({ S14204 })
);
NOR2_X1 #() 
NOR2_X1_368_ (
  .A1({ S25957[259] }),
  .A2({ S14141 }),
  .ZN({ S14205 })
);
INV_X1 #() 
INV_X1_511_ (
  .A({ S14205 }),
  .ZN({ S14206 })
);
OAI21_X1 #() 
OAI21_X1_896_ (
  .A({ S25957[260] }),
  .B1({ S14204 }),
  .B2({ S14206 }),
  .ZN({ S14207 })
);
AOI21_X1 #() 
AOI21_X1_987_ (
  .A({ S25957[260] }),
  .B1({ S14147 }),
  .B2({ S38 }),
  .ZN({ S14208 })
);
AOI21_X1 #() 
AOI21_X1_988_ (
  .A({ S38 }),
  .B1({ S14137 }),
  .B2({ S14139 }),
  .ZN({ S14209 })
);
OAI21_X1 #() 
OAI21_X1_897_ (
  .A({ S14208 }),
  .B1({ S14141 }),
  .B2({ S14209 }),
  .ZN({ S14210 })
);
OAI211_X1 #() 
OAI211_X1_621_ (
  .A({ S14210 }),
  .B({ S25957[261] }),
  .C1({ S14203 }),
  .C2({ S14207 }),
  .ZN({ S14211 })
);
AOI21_X1 #() 
AOI21_X1_989_ (
  .A({ S25957[262] }),
  .B1({ S14202 }),
  .B2({ S14211 }),
  .ZN({ S14213 })
);
OAI21_X1 #() 
OAI21_X1_898_ (
  .A({ S25957[263] }),
  .B1({ S14213 }),
  .B2({ S14185 }),
  .ZN({ S14214 })
);
NAND3_X1 #() 
NAND3_X1_1946_ (
  .A1({ S25957[256] }),
  .A2({ S14154 }),
  .A3({ S25957[257] }),
  .ZN({ S14215 })
);
INV_X1 #() 
INV_X1_512_ (
  .A({ S14177 }),
  .ZN({ S14216 })
);
INV_X1 #() 
INV_X1_513_ (
  .A({ S14197 }),
  .ZN({ S14217 })
);
OAI21_X1 #() 
OAI21_X1_899_ (
  .A({ S25957[260] }),
  .B1({ S14217 }),
  .B2({ S14194 }),
  .ZN({ S14218 })
);
AOI21_X1 #() 
AOI21_X1_990_ (
  .A({ S14218 }),
  .B1({ S14216 }),
  .B2({ S14215 }),
  .ZN({ S14219 })
);
NAND2_X1 #() 
NAND2_X1_1626_ (
  .A1({ S14158 }),
  .A2({ S14154 }),
  .ZN({ S14220 })
);
NAND2_X1 #() 
NAND2_X1_1627_ (
  .A1({ S14220 }),
  .A2({ S14176 }),
  .ZN({ S14221 })
);
INV_X1 #() 
INV_X1_514_ (
  .A({ S14221 }),
  .ZN({ S14222 })
);
NAND2_X1 #() 
NAND2_X1_1628_ (
  .A1({ S14222 }),
  .A2({ S25957[259] }),
  .ZN({ S14224 })
);
NAND3_X1 #() 
NAND3_X1_1947_ (
  .A1({ S38 }),
  .A2({ S12672 }),
  .A3({ S12675 }),
  .ZN({ S14225 })
);
NAND2_X1 #() 
NAND2_X1_1629_ (
  .A1({ S14205 }),
  .A2({ S25957[256] }),
  .ZN({ S14226 })
);
NAND2_X1 #() 
NAND2_X1_1630_ (
  .A1({ S14226 }),
  .A2({ S14225 }),
  .ZN({ S14227 })
);
NOR2_X1 #() 
NOR2_X1_369_ (
  .A1({ S14227 }),
  .A2({ S25957[260] }),
  .ZN({ S14228 })
);
AOI21_X1 #() 
AOI21_X1_991_ (
  .A({ S14219 }),
  .B1({ S14224 }),
  .B2({ S14228 }),
  .ZN({ S14229 })
);
NAND3_X1 #() 
NAND3_X1_1948_ (
  .A1({ S14156 }),
  .A2({ S14158 }),
  .A3({ S25957[258] }),
  .ZN({ S14230 })
);
AOI21_X1 #() 
AOI21_X1_992_ (
  .A({ S25957[259] }),
  .B1({ S14230 }),
  .B2({ S14147 }),
  .ZN({ S14231 })
);
NAND2_X1 #() 
NAND2_X1_1631_ (
  .A1({ S14140 }),
  .A2({ S25957[258] }),
  .ZN({ S14232 })
);
AOI21_X1 #() 
AOI21_X1_993_ (
  .A({ S38 }),
  .B1({ S14187 }),
  .B2({ S14232 }),
  .ZN({ S14233 })
);
NOR3_X1 #() 
NOR3_X1_57_ (
  .A1({ S14231 }),
  .A2({ S14233 }),
  .A3({ S14145 }),
  .ZN({ S14235 })
);
NAND2_X1 #() 
NAND2_X1_1632_ (
  .A1({ S14150 }),
  .A2({ S25957[259] }),
  .ZN({ S14236 })
);
NOR2_X1 #() 
NOR2_X1_370_ (
  .A1({ S14236 }),
  .A2({ S14160 }),
  .ZN({ S14237 })
);
AOI21_X1 #() 
AOI21_X1_994_ (
  .A({ S25957[259] }),
  .B1({ S14232 }),
  .B2({ S14220 }),
  .ZN({ S14238 })
);
NOR2_X1 #() 
NOR2_X1_371_ (
  .A1({ S14238 }),
  .A2({ S25957[260] }),
  .ZN({ S14239 })
);
INV_X1 #() 
INV_X1_515_ (
  .A({ S14239 }),
  .ZN({ S14240 })
);
OAI21_X1 #() 
OAI21_X1_900_ (
  .A({ S14186 }),
  .B1({ S14240 }),
  .B2({ S14237 }),
  .ZN({ S14241 })
);
OAI22_X1 #() 
OAI22_X1_38_ (
  .A1({ S14229 }),
  .A2({ S14186 }),
  .B1({ S14241 }),
  .B2({ S14235 }),
  .ZN({ S14242 })
);
NAND2_X1 #() 
NAND2_X1_1633_ (
  .A1({ S14242 }),
  .A2({ S25957[262] }),
  .ZN({ S14243 })
);
AOI21_X1 #() 
AOI21_X1_995_ (
  .A({ S38 }),
  .B1({ S14140 }),
  .B2({ S25957[258] }),
  .ZN({ S14244 })
);
INV_X1 #() 
INV_X1_516_ (
  .A({ S14230 }),
  .ZN({ S14246 })
);
NOR2_X1 #() 
NOR2_X1_372_ (
  .A1({ S14246 }),
  .A2({ S25957[259] }),
  .ZN({ S14247 })
);
NOR2_X1 #() 
NOR2_X1_373_ (
  .A1({ S14247 }),
  .A2({ S14244 }),
  .ZN({ S14248 })
);
NOR2_X1 #() 
NOR2_X1_374_ (
  .A1({ S14248 }),
  .A2({ S25957[260] }),
  .ZN({ S14249 })
);
NAND2_X1 #() 
NAND2_X1_1634_ (
  .A1({ S14197 }),
  .A2({ S25957[259] }),
  .ZN({ S14250 })
);
AOI21_X1 #() 
AOI21_X1_996_ (
  .A({ S25957[259] }),
  .B1({ S14230 }),
  .B2({ S14155 }),
  .ZN({ S14251 })
);
NOR2_X1 #() 
NOR2_X1_375_ (
  .A1({ S14251 }),
  .A2({ S14145 }),
  .ZN({ S14252 })
);
AOI211_X1 #() 
AOI211_X1_21_ (
  .A({ S25957[261] }),
  .B({ S14249 }),
  .C1({ S14250 }),
  .C2({ S14252 }),
  .ZN({ S14253 })
);
NAND2_X1 #() 
NAND2_X1_1635_ (
  .A1({ S14162 }),
  .A2({ S38 }),
  .ZN({ S14254 })
);
INV_X1 #() 
INV_X1_517_ (
  .A({ S14254 }),
  .ZN({ S14255 })
);
AOI22_X1 #() 
AOI22_X1_228_ (
  .A1({ S14255 }),
  .A2({ S14155 }),
  .B1({ S14161 }),
  .B2({ S14158 }),
  .ZN({ S14257 })
);
NAND2_X1 #() 
NAND2_X1_1636_ (
  .A1({ S25957[256] }),
  .A2({ S38 }),
  .ZN({ S14258 })
);
NAND3_X1 #() 
NAND3_X1_1949_ (
  .A1({ S14150 }),
  .A2({ S25957[259] }),
  .A3({ S14173 }),
  .ZN({ S14259 })
);
NAND3_X1 #() 
NAND3_X1_1950_ (
  .A1({ S14259 }),
  .A2({ S25957[260] }),
  .A3({ S14258 }),
  .ZN({ S14260 })
);
OAI21_X1 #() 
OAI21_X1_901_ (
  .A({ S14260 }),
  .B1({ S14257 }),
  .B2({ S25957[260] }),
  .ZN({ S14261 })
);
OAI21_X1 #() 
OAI21_X1_902_ (
  .A({ S14142 }),
  .B1({ S14261 }),
  .B2({ S14186 }),
  .ZN({ S14262 })
);
OAI21_X1 #() 
OAI21_X1_903_ (
  .A({ S14243 }),
  .B1({ S14253 }),
  .B2({ S14262 }),
  .ZN({ S14263 })
);
NAND2_X1 #() 
NAND2_X1_1637_ (
  .A1({ S14263 }),
  .A2({ S12121 }),
  .ZN({ S14264 })
);
NAND2_X1 #() 
NAND2_X1_1638_ (
  .A1({ S14264 }),
  .A2({ S14214 }),
  .ZN({ S14265 })
);
NAND2_X1 #() 
NAND2_X1_1639_ (
  .A1({ S14265 }),
  .A2({ S25957[367] }),
  .ZN({ S14266 })
);
NAND3_X1 #() 
NAND3_X1_1951_ (
  .A1({ S14264 }),
  .A2({ S11412 }),
  .A3({ S14214 }),
  .ZN({ S14268 })
);
NAND2_X1 #() 
NAND2_X1_1640_ (
  .A1({ S14266 }),
  .A2({ S14268 }),
  .ZN({ S25957[239] })
);
NOR2_X1 #() 
NOR2_X1_376_ (
  .A1({ S25957[239] }),
  .A2({ S25957[431] }),
  .ZN({ S14269 })
);
AND2_X1 #() 
AND2_X1_100_ (
  .A1({ S25957[239] }),
  .A2({ S25957[431] }),
  .ZN({ S14270 })
);
NOR2_X1 #() 
NOR2_X1_377_ (
  .A1({ S14270 }),
  .A2({ S14269 }),
  .ZN({ S25957[175] })
);
XNOR2_X1 #() 
XNOR2_X1_55_ (
  .A({ S25957[175] }),
  .B({ S25957[271] }),
  .ZN({ S14271 })
);
INV_X1 #() 
INV_X1_518_ (
  .A({ S14271 }),
  .ZN({ S25957[143] })
);
NOR3_X1 #() 
NOR3_X1_58_ (
  .A1({ S14174 }),
  .A2({ S14205 }),
  .A3({ S25957[260] }),
  .ZN({ S14272 })
);
INV_X1 #() 
INV_X1_519_ (
  .A({ S46 }),
  .ZN({ S14273 })
);
NAND2_X1 #() 
NAND2_X1_1641_ (
  .A1({ S14155 }),
  .A2({ S25957[259] }),
  .ZN({ S14274 })
);
NOR2_X1 #() 
NOR2_X1_378_ (
  .A1({ S14274 }),
  .A2({ S14273 }),
  .ZN({ S14276 })
);
INV_X1 #() 
INV_X1_520_ (
  .A({ S14187 }),
  .ZN({ S14277 })
);
NAND4_X1 #() 
NAND4_X1_244_ (
  .A1({ S12514 }),
  .A2({ S12517 }),
  .A3({ S14148 }),
  .A4({ S14149 }),
  .ZN({ S14278 })
);
NAND2_X1 #() 
NAND2_X1_1642_ (
  .A1({ S14278 }),
  .A2({ S38 }),
  .ZN({ S14279 })
);
NOR2_X1 #() 
NOR2_X1_379_ (
  .A1({ S14277 }),
  .A2({ S14279 }),
  .ZN({ S14280 })
);
INV_X1 #() 
INV_X1_521_ (
  .A({ S14147 }),
  .ZN({ S14281 })
);
NAND2_X1 #() 
NAND2_X1_1643_ (
  .A1({ S14188 }),
  .A2({ S25957[259] }),
  .ZN({ S14282 })
);
NOR2_X1 #() 
NOR2_X1_380_ (
  .A1({ S14282 }),
  .A2({ S14281 }),
  .ZN({ S14283 })
);
INV_X1 #() 
INV_X1_522_ (
  .A({ S14283 }),
  .ZN({ S14284 })
);
NAND2_X1 #() 
NAND2_X1_1644_ (
  .A1({ S14284 }),
  .A2({ S25957[260] }),
  .ZN({ S14285 })
);
OAI22_X1 #() 
OAI22_X1_39_ (
  .A1({ S14285 }),
  .A2({ S14280 }),
  .B1({ S14240 }),
  .B2({ S14276 }),
  .ZN({ S14287 })
);
OAI21_X1 #() 
OAI21_X1_904_ (
  .A({ S25957[260] }),
  .B1({ S14151 }),
  .B2({ S38 }),
  .ZN({ S14288 })
);
INV_X1 #() 
INV_X1_523_ (
  .A({ S14288 }),
  .ZN({ S14289 })
);
NAND2_X1 #() 
NAND2_X1_1645_ (
  .A1({ S14289 }),
  .A2({ S14163 }),
  .ZN({ S14290 })
);
OAI21_X1 #() 
OAI21_X1_905_ (
  .A({ S25957[261] }),
  .B1({ S14290 }),
  .B2({ S14283 }),
  .ZN({ S14291 })
);
OAI22_X1 #() 
OAI22_X1_40_ (
  .A1({ S14287 }),
  .A2({ S25957[261] }),
  .B1({ S14272 }),
  .B2({ S14291 }),
  .ZN({ S14292 })
);
INV_X1 #() 
INV_X1_524_ (
  .A({ S14280 }),
  .ZN({ S14293 })
);
INV_X1 #() 
INV_X1_525_ (
  .A({ S14178 }),
  .ZN({ S14294 })
);
OAI21_X1 #() 
OAI21_X1_906_ (
  .A({ S25957[259] }),
  .B1({ S14217 }),
  .B2({ S14294 }),
  .ZN({ S14295 })
);
AOI21_X1 #() 
AOI21_X1_997_ (
  .A({ S25957[260] }),
  .B1({ S14293 }),
  .B2({ S14295 }),
  .ZN({ S14296 })
);
INV_X1 #() 
INV_X1_526_ (
  .A({ S14203 }),
  .ZN({ S14298 })
);
INV_X1 #() 
INV_X1_527_ (
  .A({ S14225 }),
  .ZN({ S14299 })
);
AOI21_X1 #() 
AOI21_X1_998_ (
  .A({ S14145 }),
  .B1({ S14299 }),
  .B2({ S14158 }),
  .ZN({ S14300 })
);
AND2_X1 #() 
AND2_X1_101_ (
  .A1({ S14298 }),
  .A2({ S14300 }),
  .ZN({ S14301 })
);
OAI21_X1 #() 
OAI21_X1_907_ (
  .A({ S14186 }),
  .B1({ S14296 }),
  .B2({ S14301 }),
  .ZN({ S14302 })
);
AOI21_X1 #() 
AOI21_X1_999_ (
  .A({ S14141 }),
  .B1({ S12672 }),
  .B2({ S12675 }),
  .ZN({ S14303 })
);
NAND3_X1 #() 
NAND3_X1_1952_ (
  .A1({ S14178 }),
  .A2({ S25957[259] }),
  .A3({ S14173 }),
  .ZN({ S14304 })
);
NAND2_X1 #() 
NAND2_X1_1646_ (
  .A1({ S14303 }),
  .A2({ S25957[256] }),
  .ZN({ S14305 })
);
NAND3_X1 #() 
NAND3_X1_1953_ (
  .A1({ S14305 }),
  .A2({ S38 }),
  .A3({ S46 }),
  .ZN({ S14306 })
);
OAI211_X1 #() 
OAI211_X1_622_ (
  .A({ S14306 }),
  .B({ S14145 }),
  .C1({ S14303 }),
  .C2({ S14304 }),
  .ZN({ S14307 })
);
NAND2_X1 #() 
NAND2_X1_1647_ (
  .A1({ S14303 }),
  .A2({ S25957[259] }),
  .ZN({ S14309 })
);
NAND2_X1 #() 
NAND2_X1_1648_ (
  .A1({ S14281 }),
  .A2({ S14205 }),
  .ZN({ S14310 })
);
NAND2_X1 #() 
NAND2_X1_1649_ (
  .A1({ S14310 }),
  .A2({ S14309 }),
  .ZN({ S14311 })
);
NOR2_X1 #() 
NOR2_X1_381_ (
  .A1({ S14230 }),
  .A2({ S25957[259] }),
  .ZN({ S14312 })
);
INV_X1 #() 
INV_X1_528_ (
  .A({ S14312 }),
  .ZN({ S14313 })
);
NAND2_X1 #() 
NAND2_X1_1650_ (
  .A1({ S14313 }),
  .A2({ S25957[260] }),
  .ZN({ S14314 })
);
OAI211_X1 #() 
OAI211_X1_623_ (
  .A({ S25957[261] }),
  .B({ S14307 }),
  .C1({ S14314 }),
  .C2({ S14311 }),
  .ZN({ S14315 })
);
AOI21_X1 #() 
AOI21_X1_1000_ (
  .A({ S25957[262] }),
  .B1({ S14302 }),
  .B2({ S14315 }),
  .ZN({ S14316 })
);
AOI21_X1 #() 
AOI21_X1_1001_ (
  .A({ S14316 }),
  .B1({ S14292 }),
  .B2({ S25957[262] }),
  .ZN({ S14317 })
);
NAND2_X1 #() 
NAND2_X1_1651_ (
  .A1({ S14161 }),
  .A2({ S14176 }),
  .ZN({ S14318 })
);
NAND2_X1 #() 
NAND2_X1_1652_ (
  .A1({ S14221 }),
  .A2({ S38 }),
  .ZN({ S14320 })
);
AOI21_X1 #() 
AOI21_X1_1002_ (
  .A({ S25957[260] }),
  .B1({ S14320 }),
  .B2({ S14318 }),
  .ZN({ S14321 })
);
NOR3_X1 #() 
NOR3_X1_59_ (
  .A1({ S14159 }),
  .A2({ S14281 }),
  .A3({ S38 }),
  .ZN({ S14322 })
);
AOI211_X1 #() 
AOI211_X1_22_ (
  .A({ S14145 }),
  .B({ S14322 }),
  .C1({ S38 }),
  .C2({ S14294 }),
  .ZN({ S14323 })
);
OAI21_X1 #() 
OAI21_X1_908_ (
  .A({ S25957[261] }),
  .B1({ S14323 }),
  .B2({ S14321 }),
  .ZN({ S14324 })
);
NOR2_X1 #() 
NOR2_X1_382_ (
  .A1({ S14222 }),
  .A2({ S38 }),
  .ZN({ S14325 })
);
NAND2_X1 #() 
NAND2_X1_1653_ (
  .A1({ S14156 }),
  .A2({ S14154 }),
  .ZN({ S14326 })
);
AOI21_X1 #() 
AOI21_X1_1003_ (
  .A({ S38 }),
  .B1({ S14326 }),
  .B2({ S14197 }),
  .ZN({ S14327 })
);
NAND2_X1 #() 
NAND2_X1_1654_ (
  .A1({ S38 }),
  .A2({ S14141 }),
  .ZN({ S14328 })
);
OAI21_X1 #() 
OAI21_X1_909_ (
  .A({ S25957[260] }),
  .B1({ S14178 }),
  .B2({ S14328 }),
  .ZN({ S14329 })
);
OAI221_X1 #() 
OAI221_X1_34_ (
  .A({ S14186 }),
  .B1({ S25957[260] }),
  .B2({ S14327 }),
  .C1({ S14325 }),
  .C2({ S14329 }),
  .ZN({ S14331 })
);
NAND3_X1 #() 
NAND3_X1_1954_ (
  .A1({ S14324 }),
  .A2({ S14142 }),
  .A3({ S14331 }),
  .ZN({ S14332 })
);
NAND2_X1 #() 
NAND2_X1_1655_ (
  .A1({ S14173 }),
  .A2({ S38 }),
  .ZN({ S14333 })
);
INV_X1 #() 
INV_X1_529_ (
  .A({ S14333 }),
  .ZN({ S14334 })
);
NAND2_X1 #() 
NAND2_X1_1656_ (
  .A1({ S14334 }),
  .A2({ S14196 }),
  .ZN({ S14335 })
);
NAND3_X1 #() 
NAND3_X1_1955_ (
  .A1({ S14197 }),
  .A2({ S14188 }),
  .A3({ S38 }),
  .ZN({ S14336 })
);
NOR2_X1 #() 
NOR2_X1_383_ (
  .A1({ S14283 }),
  .A2({ S25957[260] }),
  .ZN({ S14337 })
);
AOI22_X1 #() 
AOI22_X1_229_ (
  .A1({ S14337 }),
  .A2({ S14336 }),
  .B1({ S14335 }),
  .B2({ S14289 }),
  .ZN({ S14338 })
);
NAND2_X1 #() 
NAND2_X1_1657_ (
  .A1({ S14150 }),
  .A2({ S14156 }),
  .ZN({ S14339 })
);
NAND2_X1 #() 
NAND2_X1_1658_ (
  .A1({ S14339 }),
  .A2({ S25957[259] }),
  .ZN({ S14340 })
);
NAND3_X1 #() 
NAND3_X1_1956_ (
  .A1({ S14232 }),
  .A2({ S38 }),
  .A3({ S14178 }),
  .ZN({ S14342 })
);
NAND3_X1 #() 
NAND3_X1_1957_ (
  .A1({ S14342 }),
  .A2({ S14340 }),
  .A3({ S25957[260] }),
  .ZN({ S14343 })
);
NOR2_X1 #() 
NOR2_X1_384_ (
  .A1({ S14150 }),
  .A2({ S38 }),
  .ZN({ S14344 })
);
INV_X1 #() 
INV_X1_530_ (
  .A({ S14344 }),
  .ZN({ S14345 })
);
NAND2_X1 #() 
NAND2_X1_1659_ (
  .A1({ S14178 }),
  .A2({ S25957[257] }),
  .ZN({ S14346 })
);
AOI21_X1 #() 
AOI21_X1_1004_ (
  .A({ S25957[260] }),
  .B1({ S14345 }),
  .B2({ S14346 }),
  .ZN({ S14347 })
);
INV_X1 #() 
INV_X1_531_ (
  .A({ S14347 }),
  .ZN({ S14348 })
);
AOI21_X1 #() 
AOI21_X1_1005_ (
  .A({ S14186 }),
  .B1({ S14348 }),
  .B2({ S14343 }),
  .ZN({ S14349 })
);
AOI21_X1 #() 
AOI21_X1_1006_ (
  .A({ S14349 }),
  .B1({ S14338 }),
  .B2({ S14186 }),
  .ZN({ S14350 })
);
NAND2_X1 #() 
NAND2_X1_1660_ (
  .A1({ S14350 }),
  .A2({ S25957[262] }),
  .ZN({ S14351 })
);
NAND3_X1 #() 
NAND3_X1_1958_ (
  .A1({ S14332 }),
  .A2({ S14351 }),
  .A3({ S12121 }),
  .ZN({ S14353 })
);
OAI21_X1 #() 
OAI21_X1_910_ (
  .A({ S14353 }),
  .B1({ S14317 }),
  .B2({ S12121 }),
  .ZN({ S14354 })
);
NOR2_X1 #() 
NOR2_X1_385_ (
  .A1({ S14354 }),
  .A2({ S8504 }),
  .ZN({ S14355 })
);
NAND2_X1 #() 
NAND2_X1_1661_ (
  .A1({ S14354 }),
  .A2({ S8504 }),
  .ZN({ S14356 })
);
INV_X1 #() 
INV_X1_532_ (
  .A({ S14356 }),
  .ZN({ S14357 })
);
NOR2_X1 #() 
NOR2_X1_386_ (
  .A1({ S14357 }),
  .A2({ S14355 }),
  .ZN({ S25957[206] })
);
NAND2_X1 #() 
NAND2_X1_1662_ (
  .A1({ S25957[206] }),
  .A2({ S25957[398] }),
  .ZN({ S14358 })
);
INV_X1 #() 
INV_X1_533_ (
  .A({ S25957[206] }),
  .ZN({ S14359 })
);
NAND2_X1 #() 
NAND2_X1_1663_ (
  .A1({ S14359 }),
  .A2({ S8507 }),
  .ZN({ S14360 })
);
NAND2_X1 #() 
NAND2_X1_1664_ (
  .A1({ S14360 }),
  .A2({ S14358 }),
  .ZN({ S14361 })
);
INV_X1 #() 
INV_X1_534_ (
  .A({ S14361 }),
  .ZN({ S25957[142] })
);
NOR2_X1 #() 
NOR2_X1_387_ (
  .A1({ S11586 }),
  .A2({ S11587 }),
  .ZN({ S14363 })
);
INV_X1 #() 
INV_X1_535_ (
  .A({ S14363 }),
  .ZN({ S25957[333] })
);
NAND2_X1 #() 
NAND2_X1_1665_ (
  .A1({ S8577 }),
  .A2({ S8578 }),
  .ZN({ S25957[493] })
);
NAND2_X1 #() 
NAND2_X1_1666_ (
  .A1({ S11579 }),
  .A2({ S11577 }),
  .ZN({ S14364 })
);
XOR2_X1 #() 
XOR2_X1_26_ (
  .A({ S14364 }),
  .B({ S25957[493] }),
  .Z({ S14365 })
);
INV_X1 #() 
INV_X1_536_ (
  .A({ S14365 }),
  .ZN({ S25957[365] })
);
INV_X1 #() 
INV_X1_537_ (
  .A({ S14304 }),
  .ZN({ S14366 })
);
OAI21_X1 #() 
OAI21_X1_911_ (
  .A({ S25957[260] }),
  .B1({ S14171 }),
  .B2({ S14154 }),
  .ZN({ S14367 })
);
NAND2_X1 #() 
NAND2_X1_1667_ (
  .A1({ S14337 }),
  .A2({ S14313 }),
  .ZN({ S14368 })
);
OAI21_X1 #() 
OAI21_X1_912_ (
  .A({ S14368 }),
  .B1({ S14366 }),
  .B2({ S14367 }),
  .ZN({ S14370 })
);
INV_X1 #() 
INV_X1_538_ (
  .A({ S14278 }),
  .ZN({ S14371 })
);
NAND2_X1 #() 
NAND2_X1_1668_ (
  .A1({ S14205 }),
  .A2({ S25957[258] }),
  .ZN({ S14372 })
);
NAND2_X1 #() 
NAND2_X1_1669_ (
  .A1({ S14156 }),
  .A2({ S25957[259] }),
  .ZN({ S14373 })
);
OAI221_X1 #() 
OAI221_X1_35_ (
  .A({ S14300 }),
  .B1({ S14373 }),
  .B2({ S14371 }),
  .C1({ S25957[256] }),
  .C2({ S14372 }),
  .ZN({ S14374 })
);
NAND3_X1 #() 
NAND3_X1_1959_ (
  .A1({ S14140 }),
  .A2({ S14162 }),
  .A3({ S25957[259] }),
  .ZN({ S14375 })
);
NAND4_X1 #() 
NAND4_X1_245_ (
  .A1({ S14375 }),
  .A2({ S14206 }),
  .A3({ S14150 }),
  .A4({ S14145 }),
  .ZN({ S14376 })
);
AOI21_X1 #() 
AOI21_X1_1007_ (
  .A({ S14186 }),
  .B1({ S14374 }),
  .B2({ S14376 }),
  .ZN({ S14377 })
);
AOI21_X1 #() 
AOI21_X1_1008_ (
  .A({ S14377 }),
  .B1({ S14370 }),
  .B2({ S14186 }),
  .ZN({ S14378 })
);
NOR2_X1 #() 
NOR2_X1_388_ (
  .A1({ S14378 }),
  .A2({ S12121 }),
  .ZN({ S14379 })
);
NAND2_X1 #() 
NAND2_X1_1670_ (
  .A1({ S14160 }),
  .A2({ S14196 }),
  .ZN({ S14381 })
);
NAND2_X1 #() 
NAND2_X1_1671_ (
  .A1({ S14381 }),
  .A2({ S25957[259] }),
  .ZN({ S14382 })
);
OAI22_X1 #() 
OAI22_X1_41_ (
  .A1({ S14246 }),
  .A2({ S14382 }),
  .B1({ S14221 }),
  .B2({ S25957[259] }),
  .ZN({ S14383 })
);
NAND2_X1 #() 
NAND2_X1_1672_ (
  .A1({ S14383 }),
  .A2({ S25957[260] }),
  .ZN({ S14384 })
);
NAND3_X1 #() 
NAND3_X1_1960_ (
  .A1({ S14178 }),
  .A2({ S14156 }),
  .A3({ S38 }),
  .ZN({ S14385 })
);
OAI21_X1 #() 
OAI21_X1_913_ (
  .A({ S14385 }),
  .B1({ S38 }),
  .B2({ S25957[256] }),
  .ZN({ S14386 })
);
OAI211_X1 #() 
OAI211_X1_624_ (
  .A({ S14384 }),
  .B({ S25957[261] }),
  .C1({ S25957[260] }),
  .C2({ S14386 }),
  .ZN({ S14387 })
);
NAND4_X1 #() 
NAND4_X1_246_ (
  .A1({ S14178 }),
  .A2({ S14278 }),
  .A3({ S25957[259] }),
  .A4({ S14176 }),
  .ZN({ S14388 })
);
NAND3_X1 #() 
NAND3_X1_1961_ (
  .A1({ S14381 }),
  .A2({ S38 }),
  .A3({ S14150 }),
  .ZN({ S14389 })
);
NAND2_X1 #() 
NAND2_X1_1673_ (
  .A1({ S14389 }),
  .A2({ S14388 }),
  .ZN({ S14390 })
);
NAND2_X1 #() 
NAND2_X1_1674_ (
  .A1({ S14390 }),
  .A2({ S14145 }),
  .ZN({ S14392 })
);
INV_X1 #() 
INV_X1_539_ (
  .A({ S14392 }),
  .ZN({ S14393 })
);
NAND2_X1 #() 
NAND2_X1_1675_ (
  .A1({ S14232 }),
  .A2({ S14215 }),
  .ZN({ S14394 })
);
NAND3_X1 #() 
NAND3_X1_1962_ (
  .A1({ S14158 }),
  .A2({ S25957[259] }),
  .A3({ S14154 }),
  .ZN({ S14395 })
);
INV_X1 #() 
INV_X1_540_ (
  .A({ S14395 }),
  .ZN({ S14396 })
);
AOI211_X1 #() 
AOI211_X1_23_ (
  .A({ S14145 }),
  .B({ S14396 }),
  .C1({ S38 }),
  .C2({ S14394 }),
  .ZN({ S14397 })
);
OAI21_X1 #() 
OAI21_X1_914_ (
  .A({ S14186 }),
  .B1({ S14393 }),
  .B2({ S14397 }),
  .ZN({ S14398 })
);
NAND2_X1 #() 
NAND2_X1_1676_ (
  .A1({ S14398 }),
  .A2({ S14387 }),
  .ZN({ S14399 })
);
NOR2_X1 #() 
NOR2_X1_389_ (
  .A1({ S14399 }),
  .A2({ S25957[263] }),
  .ZN({ S14400 })
);
OAI21_X1 #() 
OAI21_X1_915_ (
  .A({ S25957[262] }),
  .B1({ S14379 }),
  .B2({ S14400 }),
  .ZN({ S14401 })
);
NAND2_X1 #() 
NAND2_X1_1677_ (
  .A1({ S14197 }),
  .A2({ S14188 }),
  .ZN({ S14403 })
);
NOR2_X1 #() 
NOR2_X1_390_ (
  .A1({ S14173 }),
  .A2({ S25957[256] }),
  .ZN({ S14404 })
);
INV_X1 #() 
INV_X1_541_ (
  .A({ S14404 }),
  .ZN({ S14405 })
);
NAND2_X1 #() 
NAND2_X1_1678_ (
  .A1({ S14405 }),
  .A2({ S25957[259] }),
  .ZN({ S14406 })
);
NOR2_X1 #() 
NOR2_X1_391_ (
  .A1({ S14140 }),
  .A2({ S25957[258] }),
  .ZN({ S14407 })
);
AOI21_X1 #() 
AOI21_X1_1009_ (
  .A({ S25957[260] }),
  .B1({ S14407 }),
  .B2({ S38 }),
  .ZN({ S14408 })
);
OAI21_X1 #() 
OAI21_X1_916_ (
  .A({ S14408 }),
  .B1({ S14406 }),
  .B2({ S14403 }),
  .ZN({ S14409 })
);
NOR2_X1 #() 
NOR2_X1_392_ (
  .A1({ S14155 }),
  .A2({ S14273 }),
  .ZN({ S14410 })
);
NAND2_X1 #() 
NAND2_X1_1679_ (
  .A1({ S14410 }),
  .A2({ S25957[259] }),
  .ZN({ S14411 })
);
INV_X1 #() 
INV_X1_542_ (
  .A({ S14328 }),
  .ZN({ S14412 })
);
AOI21_X1 #() 
AOI21_X1_1010_ (
  .A({ S14145 }),
  .B1({ S14412 }),
  .B2({ S14178 }),
  .ZN({ S14414 })
);
AOI21_X1 #() 
AOI21_X1_1011_ (
  .A({ S25957[261] }),
  .B1({ S14411 }),
  .B2({ S14414 }),
  .ZN({ S14415 })
);
NAND2_X1 #() 
NAND2_X1_1680_ (
  .A1({ S14278 }),
  .A2({ S25957[259] }),
  .ZN({ S14416 })
);
OAI221_X1 #() 
OAI221_X1_36_ (
  .A({ S25957[260] }),
  .B1({ S14194 }),
  .B2({ S45 }),
  .C1({ S14221 }),
  .C2({ S14416 }),
  .ZN({ S14417 })
);
AOI21_X1 #() 
AOI21_X1_1012_ (
  .A({ S25957[259] }),
  .B1({ S14140 }),
  .B2({ S14176 }),
  .ZN({ S14418 })
);
NAND2_X1 #() 
NAND2_X1_1681_ (
  .A1({ S14145 }),
  .A2({ S14191 }),
  .ZN({ S14419 })
);
OAI21_X1 #() 
OAI21_X1_917_ (
  .A({ S14417 }),
  .B1({ S14418 }),
  .B2({ S14419 }),
  .ZN({ S14420 })
);
AOI22_X1 #() 
AOI22_X1_230_ (
  .A1({ S14420 }),
  .A2({ S25957[261] }),
  .B1({ S14409 }),
  .B2({ S14415 }),
  .ZN({ S14421 })
);
NOR2_X1 #() 
NOR2_X1_393_ (
  .A1({ S14421 }),
  .A2({ S12121 }),
  .ZN({ S14422 })
);
NAND3_X1 #() 
NAND3_X1_1963_ (
  .A1({ S14274 }),
  .A2({ S14310 }),
  .A3({ S25957[260] }),
  .ZN({ S14423 })
);
INV_X1 #() 
INV_X1_543_ (
  .A({ S14279 }),
  .ZN({ S14425 })
);
OAI21_X1 #() 
OAI21_X1_918_ (
  .A({ S14347 }),
  .B1({ S14344 }),
  .B2({ S14425 }),
  .ZN({ S14426 })
);
NAND3_X1 #() 
NAND3_X1_1964_ (
  .A1({ S14426 }),
  .A2({ S25957[261] }),
  .A3({ S14423 }),
  .ZN({ S14427 })
);
NAND3_X1 #() 
NAND3_X1_1965_ (
  .A1({ S25957[256] }),
  .A2({ S14154 }),
  .A3({ S14141 }),
  .ZN({ S14428 })
);
NAND2_X1 #() 
NAND2_X1_1682_ (
  .A1({ S14230 }),
  .A2({ S14428 }),
  .ZN({ S14429 })
);
NAND4_X1 #() 
NAND4_X1_247_ (
  .A1({ S14147 }),
  .A2({ S14156 }),
  .A3({ S14158 }),
  .A4({ S38 }),
  .ZN({ S14430 })
);
OAI21_X1 #() 
OAI21_X1_919_ (
  .A({ S14430 }),
  .B1({ S14429 }),
  .B2({ S38 }),
  .ZN({ S14431 })
);
NOR2_X1 #() 
NOR2_X1_394_ (
  .A1({ S25957[257] }),
  .A2({ S38 }),
  .ZN({ S14432 })
);
NAND2_X1 #() 
NAND2_X1_1683_ (
  .A1({ S14432 }),
  .A2({ S25957[256] }),
  .ZN({ S14433 })
);
OAI21_X1 #() 
OAI21_X1_920_ (
  .A({ S14433 }),
  .B1({ S14226 }),
  .B2({ S14154 }),
  .ZN({ S14434 })
);
AOI21_X1 #() 
AOI21_X1_1013_ (
  .A({ S25957[261] }),
  .B1({ S14434 }),
  .B2({ S14145 }),
  .ZN({ S14436 })
);
OAI21_X1 #() 
OAI21_X1_921_ (
  .A({ S14436 }),
  .B1({ S14431 }),
  .B2({ S14145 }),
  .ZN({ S14437 })
);
AOI21_X1 #() 
AOI21_X1_1014_ (
  .A({ S25957[263] }),
  .B1({ S14427 }),
  .B2({ S14437 }),
  .ZN({ S14438 })
);
OAI21_X1 #() 
OAI21_X1_922_ (
  .A({ S14142 }),
  .B1({ S14422 }),
  .B2({ S14438 }),
  .ZN({ S14439 })
);
NAND3_X1 #() 
NAND3_X1_1966_ (
  .A1({ S14401 }),
  .A2({ S25957[365] }),
  .A3({ S14439 }),
  .ZN({ S14440 })
);
OR2_X1 #() 
OR2_X1_25_ (
  .A1({ S14421 }),
  .A2({ S25957[262] }),
  .ZN({ S14441 })
);
OAI211_X1 #() 
OAI211_X1_625_ (
  .A({ S14441 }),
  .B({ S25957[263] }),
  .C1({ S14142 }),
  .C2({ S14378 }),
  .ZN({ S14442 })
);
NAND2_X1 #() 
NAND2_X1_1684_ (
  .A1({ S14427 }),
  .A2({ S14437 }),
  .ZN({ S14443 })
);
AOI21_X1 #() 
AOI21_X1_1015_ (
  .A({ S25957[263] }),
  .B1({ S14443 }),
  .B2({ S14142 }),
  .ZN({ S14444 })
);
OAI21_X1 #() 
OAI21_X1_923_ (
  .A({ S14444 }),
  .B1({ S14399 }),
  .B2({ S14142 }),
  .ZN({ S14445 })
);
NAND3_X1 #() 
NAND3_X1_1967_ (
  .A1({ S14442 }),
  .A2({ S14365 }),
  .A3({ S14445 }),
  .ZN({ S14447 })
);
NAND2_X1 #() 
NAND2_X1_1685_ (
  .A1({ S14440 }),
  .A2({ S14447 }),
  .ZN({ S25957[237] })
);
INV_X1 #() 
INV_X1_544_ (
  .A({ S25957[237] }),
  .ZN({ S14448 })
);
NAND2_X1 #() 
NAND2_X1_1686_ (
  .A1({ S14448 }),
  .A2({ S25957[333] }),
  .ZN({ S14449 })
);
NAND2_X1 #() 
NAND2_X1_1687_ (
  .A1({ S25957[237] }),
  .A2({ S14363 }),
  .ZN({ S14450 })
);
NAND2_X1 #() 
NAND2_X1_1688_ (
  .A1({ S14449 }),
  .A2({ S14450 }),
  .ZN({ S25957[205] })
);
NAND2_X1 #() 
NAND2_X1_1689_ (
  .A1({ S25957[205] }),
  .A2({ S25957[397] }),
  .ZN({ S14451 })
);
NAND3_X1 #() 
NAND3_X1_1968_ (
  .A1({ S14449 }),
  .A2({ S14450 }),
  .A3({ S10559 }),
  .ZN({ S14452 })
);
AND2_X1 #() 
AND2_X1_102_ (
  .A1({ S14451 }),
  .A2({ S14452 }),
  .ZN({ S25957[141] })
);
NAND2_X1 #() 
NAND2_X1_1690_ (
  .A1({ S11656 }),
  .A2({ S11659 }),
  .ZN({ S25957[300] })
);
NOR2_X1 #() 
NOR2_X1_395_ (
  .A1({ S11654 }),
  .A2({ S11655 }),
  .ZN({ S14454 })
);
INV_X1 #() 
INV_X1_545_ (
  .A({ S14454 }),
  .ZN({ S25957[332] })
);
XNOR2_X1 #() 
XNOR2_X1_56_ (
  .A({ S8655 }),
  .B({ S25957[620] }),
  .ZN({ S25957[492] })
);
XOR2_X1 #() 
XOR2_X1_27_ (
  .A({ S11657 }),
  .B({ S25957[492] }),
  .Z({ S25957[364] })
);
INV_X1 #() 
INV_X1_546_ (
  .A({ S25957[364] }),
  .ZN({ S14455 })
);
NAND3_X1 #() 
NAND3_X1_1969_ (
  .A1({ S14181 }),
  .A2({ S14395 }),
  .A3({ S25957[260] }),
  .ZN({ S14456 })
);
NOR2_X1 #() 
NOR2_X1_396_ (
  .A1({ S14160 }),
  .A2({ S25957[259] }),
  .ZN({ S14457 })
);
NAND2_X1 #() 
NAND2_X1_1691_ (
  .A1({ S14457 }),
  .A2({ S14196 }),
  .ZN({ S14458 })
);
NAND3_X1 #() 
NAND3_X1_1970_ (
  .A1({ S14458 }),
  .A2({ S14145 }),
  .A3({ S14259 }),
  .ZN({ S14459 })
);
NAND3_X1 #() 
NAND3_X1_1971_ (
  .A1({ S14459 }),
  .A2({ S14456 }),
  .A3({ S25957[261] }),
  .ZN({ S14460 })
);
AOI21_X1 #() 
AOI21_X1_1016_ (
  .A({ S25957[260] }),
  .B1({ S14161 }),
  .B2({ S14158 }),
  .ZN({ S14462 })
);
OAI21_X1 #() 
OAI21_X1_924_ (
  .A({ S14462 }),
  .B1({ S14371 }),
  .B2({ S14333 }),
  .ZN({ S14463 })
);
NOR2_X1 #() 
NOR2_X1_397_ (
  .A1({ S14418 }),
  .A2({ S14145 }),
  .ZN({ S14464 })
);
OAI21_X1 #() 
OAI21_X1_925_ (
  .A({ S14464 }),
  .B1({ S14294 }),
  .B2({ S14191 }),
  .ZN({ S14465 })
);
NAND3_X1 #() 
NAND3_X1_1972_ (
  .A1({ S14465 }),
  .A2({ S14463 }),
  .A3({ S14186 }),
  .ZN({ S14466 })
);
NAND2_X1 #() 
NAND2_X1_1692_ (
  .A1({ S14460 }),
  .A2({ S14466 }),
  .ZN({ S14467 })
);
NAND2_X1 #() 
NAND2_X1_1693_ (
  .A1({ S14467 }),
  .A2({ S25957[262] }),
  .ZN({ S14468 })
);
NOR2_X1 #() 
NOR2_X1_398_ (
  .A1({ S14236 }),
  .A2({ S25957[257] }),
  .ZN({ S14469 })
);
AOI21_X1 #() 
AOI21_X1_1017_ (
  .A({ S25957[259] }),
  .B1({ S14326 }),
  .B2({ S14197 }),
  .ZN({ S14470 })
);
OR2_X1 #() 
OR2_X1_26_ (
  .A1({ S14470 }),
  .A2({ S25957[260] }),
  .ZN({ S14471 })
);
NAND2_X1 #() 
NAND2_X1_1694_ (
  .A1({ S14151 }),
  .A2({ S14176 }),
  .ZN({ S14473 })
);
OAI21_X1 #() 
OAI21_X1_926_ (
  .A({ S38 }),
  .B1({ S14166 }),
  .B2({ S14204 }),
  .ZN({ S14474 })
);
OAI21_X1 #() 
OAI21_X1_927_ (
  .A({ S14474 }),
  .B1({ S14236 }),
  .B2({ S14473 }),
  .ZN({ S14475 })
);
OAI22_X1 #() 
OAI22_X1_42_ (
  .A1({ S14471 }),
  .A2({ S14469 }),
  .B1({ S14475 }),
  .B2({ S14145 }),
  .ZN({ S14476 })
);
INV_X1 #() 
INV_X1_547_ (
  .A({ S14158 }),
  .ZN({ S14477 })
);
AOI22_X1 #() 
AOI22_X1_231_ (
  .A1({ S14477 }),
  .A2({ S14225 }),
  .B1({ S14196 }),
  .B2({ S14160 }),
  .ZN({ S14478 })
);
AOI21_X1 #() 
AOI21_X1_1018_ (
  .A({ S25957[259] }),
  .B1({ S14187 }),
  .B2({ S14232 }),
  .ZN({ S14479 })
);
NAND4_X1 #() 
NAND4_X1_248_ (
  .A1({ S14196 }),
  .A2({ S25957[258] }),
  .A3({ S25957[259] }),
  .A4({ S25957[257] }),
  .ZN({ S14480 })
);
NAND3_X1 #() 
NAND3_X1_1973_ (
  .A1({ S14395 }),
  .A2({ S14480 }),
  .A3({ S14145 }),
  .ZN({ S14481 })
);
OAI221_X1 #() 
OAI221_X1_37_ (
  .A({ S25957[261] }),
  .B1({ S14478 }),
  .B2({ S14145 }),
  .C1({ S14479 }),
  .C2({ S14481 }),
  .ZN({ S14482 })
);
OAI21_X1 #() 
OAI21_X1_928_ (
  .A({ S14482 }),
  .B1({ S14476 }),
  .B2({ S25957[261] }),
  .ZN({ S14484 })
);
NAND2_X1 #() 
NAND2_X1_1695_ (
  .A1({ S14484 }),
  .A2({ S14142 }),
  .ZN({ S14485 })
);
NAND2_X1 #() 
NAND2_X1_1696_ (
  .A1({ S14485 }),
  .A2({ S14468 }),
  .ZN({ S14486 })
);
NAND2_X1 #() 
NAND2_X1_1697_ (
  .A1({ S14486 }),
  .A2({ S25957[263] }),
  .ZN({ S14487 })
);
INV_X1 #() 
INV_X1_548_ (
  .A({ S14224 }),
  .ZN({ S14488 })
);
AND2_X1 #() 
AND2_X1_103_ (
  .A1({ S14411 }),
  .A2({ S14226 }),
  .ZN({ S14489 })
);
OAI22_X1 #() 
OAI22_X1_43_ (
  .A1({ S14489 }),
  .A2({ S25957[260] }),
  .B1({ S14488 }),
  .B2({ S14367 }),
  .ZN({ S14490 })
);
NAND2_X1 #() 
NAND2_X1_1698_ (
  .A1({ S14490 }),
  .A2({ S25957[261] }),
  .ZN({ S14491 })
);
INV_X1 #() 
INV_X1_549_ (
  .A({ S14180 }),
  .ZN({ S14492 })
);
INV_X1 #() 
INV_X1_550_ (
  .A({ S14181 }),
  .ZN({ S14493 })
);
NAND3_X1 #() 
NAND3_X1_1974_ (
  .A1({ S14150 }),
  .A2({ S25957[259] }),
  .A3({ S46 }),
  .ZN({ S14494 })
);
INV_X1 #() 
INV_X1_551_ (
  .A({ S14494 }),
  .ZN({ S14495 })
);
AOI21_X1 #() 
AOI21_X1_1019_ (
  .A({ S14495 }),
  .B1({ S14493 }),
  .B2({ S14492 }),
  .ZN({ S14496 })
);
OAI21_X1 #() 
OAI21_X1_929_ (
  .A({ S14464 }),
  .B1({ S38 }),
  .B2({ S14152 }),
  .ZN({ S14497 })
);
OAI21_X1 #() 
OAI21_X1_930_ (
  .A({ S14497 }),
  .B1({ S14496 }),
  .B2({ S25957[260] }),
  .ZN({ S14498 })
);
NAND2_X1 #() 
NAND2_X1_1699_ (
  .A1({ S14498 }),
  .A2({ S14186 }),
  .ZN({ S14499 })
);
AOI21_X1 #() 
AOI21_X1_1020_ (
  .A({ S25957[262] }),
  .B1({ S14491 }),
  .B2({ S14499 }),
  .ZN({ S14500 })
);
NAND3_X1 #() 
NAND3_X1_1975_ (
  .A1({ S14473 }),
  .A2({ S38 }),
  .A3({ S14150 }),
  .ZN({ S14501 })
);
AOI21_X1 #() 
AOI21_X1_1021_ (
  .A({ S14145 }),
  .B1({ S14298 }),
  .B2({ S14501 }),
  .ZN({ S14502 })
);
NAND2_X1 #() 
NAND2_X1_1700_ (
  .A1({ S25957[258] }),
  .A2({ S25957[259] }),
  .ZN({ S14503 })
);
NAND2_X1 #() 
NAND2_X1_1701_ (
  .A1({ S14279 }),
  .A2({ S14503 }),
  .ZN({ S14505 })
);
AND2_X1 #() 
AND2_X1_104_ (
  .A1({ S14408 }),
  .A2({ S14505 }),
  .ZN({ S14506 })
);
OAI21_X1 #() 
OAI21_X1_931_ (
  .A({ S14186 }),
  .B1({ S14502 }),
  .B2({ S14506 }),
  .ZN({ S14507 })
);
NAND2_X1 #() 
NAND2_X1_1702_ (
  .A1({ S14187 }),
  .A2({ S14197 }),
  .ZN({ S14508 })
);
OAI211_X1 #() 
OAI211_X1_626_ (
  .A({ S14145 }),
  .B({ S14388 }),
  .C1({ S14508 }),
  .C2({ S25957[259] }),
  .ZN({ S14509 })
);
INV_X1 #() 
INV_X1_552_ (
  .A({ S149 }),
  .ZN({ S14510 })
);
OAI21_X1 #() 
OAI21_X1_932_ (
  .A({ S25957[260] }),
  .B1({ S14510 }),
  .B2({ S25957[258] }),
  .ZN({ S14511 })
);
NAND3_X1 #() 
NAND3_X1_1976_ (
  .A1({ S14509 }),
  .A2({ S25957[261] }),
  .A3({ S14511 }),
  .ZN({ S14512 })
);
AOI21_X1 #() 
AOI21_X1_1022_ (
  .A({ S14142 }),
  .B1({ S14507 }),
  .B2({ S14512 }),
  .ZN({ S14513 })
);
OAI21_X1 #() 
OAI21_X1_933_ (
  .A({ S12121 }),
  .B1({ S14500 }),
  .B2({ S14513 }),
  .ZN({ S14514 })
);
NAND3_X1 #() 
NAND3_X1_1977_ (
  .A1({ S14487 }),
  .A2({ S14514 }),
  .A3({ S14455 }),
  .ZN({ S14516 })
);
NAND3_X1 #() 
NAND3_X1_1978_ (
  .A1({ S14485 }),
  .A2({ S14468 }),
  .A3({ S25957[263] }),
  .ZN({ S14517 })
);
OR3_X1 #() 
OR3_X1_6_ (
  .A1({ S14500 }),
  .A2({ S14513 }),
  .A3({ S25957[263] }),
  .ZN({ S14518 })
);
NAND3_X1 #() 
NAND3_X1_1979_ (
  .A1({ S14518 }),
  .A2({ S25957[364] }),
  .A3({ S14517 }),
  .ZN({ S14519 })
);
NAND3_X1 #() 
NAND3_X1_1980_ (
  .A1({ S14519 }),
  .A2({ S25957[332] }),
  .A3({ S14516 }),
  .ZN({ S14520 })
);
NAND3_X1 #() 
NAND3_X1_1981_ (
  .A1({ S14518 }),
  .A2({ S14455 }),
  .A3({ S14517 }),
  .ZN({ S14521 })
);
NAND3_X1 #() 
NAND3_X1_1982_ (
  .A1({ S14487 }),
  .A2({ S14514 }),
  .A3({ S25957[364] }),
  .ZN({ S14522 })
);
NAND3_X1 #() 
NAND3_X1_1983_ (
  .A1({ S14521 }),
  .A2({ S14454 }),
  .A3({ S14522 }),
  .ZN({ S14523 })
);
NAND3_X1 #() 
NAND3_X1_1984_ (
  .A1({ S14520 }),
  .A2({ S14523 }),
  .A3({ S25957[396] }),
  .ZN({ S14524 })
);
NAND3_X1 #() 
NAND3_X1_1985_ (
  .A1({ S14521 }),
  .A2({ S25957[332] }),
  .A3({ S14522 }),
  .ZN({ S14525 })
);
NAND3_X1 #() 
NAND3_X1_1986_ (
  .A1({ S14519 }),
  .A2({ S14454 }),
  .A3({ S14516 }),
  .ZN({ S14527 })
);
NAND3_X1 #() 
NAND3_X1_1987_ (
  .A1({ S14525 }),
  .A2({ S14527 }),
  .A3({ S10526 }),
  .ZN({ S14528 })
);
NAND2_X1 #() 
NAND2_X1_1703_ (
  .A1({ S14524 }),
  .A2({ S14528 }),
  .ZN({ S25957[140] })
);
NAND2_X1 #() 
NAND2_X1_1704_ (
  .A1({ S8754 }),
  .A2({ S8747 }),
  .ZN({ S25957[491] })
);
XNOR2_X1 #() 
XNOR2_X1_57_ (
  .A({ S25957[491] }),
  .B({ S11665 }),
  .ZN({ S25957[459] })
);
INV_X1 #() 
INV_X1_553_ (
  .A({ S25957[459] }),
  .ZN({ S14529 })
);
AOI22_X1 #() 
AOI22_X1_232_ (
  .A1({ S14247 }),
  .A2({ S14428 }),
  .B1({ S25957[259] }),
  .B2({ S14166 }),
  .ZN({ S14530 })
);
NAND3_X1 #() 
NAND3_X1_1988_ (
  .A1({ S14339 }),
  .A2({ S14145 }),
  .A3({ S14503 }),
  .ZN({ S14531 })
);
OAI211_X1 #() 
OAI211_X1_627_ (
  .A({ S14186 }),
  .B({ S14531 }),
  .C1({ S14530 }),
  .C2({ S14145 }),
  .ZN({ S14532 })
);
AOI21_X1 #() 
AOI21_X1_1023_ (
  .A({ S14303 }),
  .B1({ S14150 }),
  .B2({ S14156 }),
  .ZN({ S14533 })
);
NAND2_X1 #() 
NAND2_X1_1705_ (
  .A1({ S14533 }),
  .A2({ S25957[259] }),
  .ZN({ S14535 })
);
OAI21_X1 #() 
OAI21_X1_934_ (
  .A({ S14535 }),
  .B1({ S14159 }),
  .B2({ S14279 }),
  .ZN({ S14536 })
);
NAND2_X1 #() 
NAND2_X1_1706_ (
  .A1({ S14536 }),
  .A2({ S14145 }),
  .ZN({ S14537 })
);
NAND3_X1 #() 
NAND3_X1_1989_ (
  .A1({ S14197 }),
  .A2({ S38 }),
  .A3({ S14158 }),
  .ZN({ S14538 })
);
NOR2_X1 #() 
NOR2_X1_399_ (
  .A1({ S14495 }),
  .A2({ S14145 }),
  .ZN({ S14539 })
);
AOI21_X1 #() 
AOI21_X1_1024_ (
  .A({ S14186 }),
  .B1({ S14539 }),
  .B2({ S14538 }),
  .ZN({ S14540 })
);
AOI21_X1 #() 
AOI21_X1_1025_ (
  .A({ S14142 }),
  .B1({ S14537 }),
  .B2({ S14540 }),
  .ZN({ S14541 })
);
NAND2_X1 #() 
NAND2_X1_1707_ (
  .A1({ S14532 }),
  .A2({ S14541 }),
  .ZN({ S14542 })
);
NAND2_X1 #() 
NAND2_X1_1708_ (
  .A1({ S14156 }),
  .A2({ S14162 }),
  .ZN({ S14543 })
);
NAND3_X1 #() 
NAND3_X1_1990_ (
  .A1({ S14543 }),
  .A2({ S25957[259] }),
  .A3({ S14278 }),
  .ZN({ S14544 })
);
NAND3_X1 #() 
NAND3_X1_1991_ (
  .A1({ S14334 }),
  .A2({ S14197 }),
  .A3({ S14188 }),
  .ZN({ S14546 })
);
NAND3_X1 #() 
NAND3_X1_1992_ (
  .A1({ S14546 }),
  .A2({ S14145 }),
  .A3({ S14544 }),
  .ZN({ S14547 })
);
AOI21_X1 #() 
AOI21_X1_1026_ (
  .A({ S14145 }),
  .B1({ S14195 }),
  .B2({ S14188 }),
  .ZN({ S14548 })
);
OAI21_X1 #() 
OAI21_X1_935_ (
  .A({ S14548 }),
  .B1({ S14177 }),
  .B2({ S14410 }),
  .ZN({ S14549 })
);
NAND3_X1 #() 
NAND3_X1_1993_ (
  .A1({ S14549 }),
  .A2({ S25957[261] }),
  .A3({ S14547 }),
  .ZN({ S14550 })
);
NAND2_X1 #() 
NAND2_X1_1709_ (
  .A1({ S14304 }),
  .A2({ S14433 }),
  .ZN({ S14551 })
);
NAND2_X1 #() 
NAND2_X1_1710_ (
  .A1({ S14339 }),
  .A2({ S38 }),
  .ZN({ S14552 })
);
NAND4_X1 #() 
NAND4_X1_249_ (
  .A1({ S14156 }),
  .A2({ S14158 }),
  .A3({ S25957[259] }),
  .A4({ S25957[258] }),
  .ZN({ S14553 })
);
NAND2_X1 #() 
NAND2_X1_1711_ (
  .A1({ S14552 }),
  .A2({ S14553 }),
  .ZN({ S14554 })
);
OAI21_X1 #() 
OAI21_X1_936_ (
  .A({ S14145 }),
  .B1({ S14554 }),
  .B2({ S14192 }),
  .ZN({ S14555 })
);
OAI21_X1 #() 
OAI21_X1_937_ (
  .A({ S25957[260] }),
  .B1({ S14371 }),
  .B2({ S14333 }),
  .ZN({ S14557 })
);
OAI21_X1 #() 
OAI21_X1_938_ (
  .A({ S14555 }),
  .B1({ S14551 }),
  .B2({ S14557 }),
  .ZN({ S14558 })
);
OAI211_X1 #() 
OAI211_X1_628_ (
  .A({ S14142 }),
  .B({ S14550 }),
  .C1({ S14558 }),
  .C2({ S25957[261] }),
  .ZN({ S14559 })
);
NAND2_X1 #() 
NAND2_X1_1712_ (
  .A1({ S14559 }),
  .A2({ S14542 }),
  .ZN({ S14560 })
);
NAND2_X1 #() 
NAND2_X1_1713_ (
  .A1({ S14560 }),
  .A2({ S25957[263] }),
  .ZN({ S14561 })
);
NAND2_X1 #() 
NAND2_X1_1714_ (
  .A1({ S14457 }),
  .A2({ S14158 }),
  .ZN({ S14562 })
);
AOI21_X1 #() 
AOI21_X1_1027_ (
  .A({ S25957[260] }),
  .B1({ S14209 }),
  .B2({ S14162 }),
  .ZN({ S14563 })
);
AOI22_X1 #() 
AOI22_X1_233_ (
  .A1({ S14252 }),
  .A2({ S14284 }),
  .B1({ S14563 }),
  .B2({ S14562 }),
  .ZN({ S14564 })
);
NAND4_X1 #() 
NAND4_X1_250_ (
  .A1({ S14151 }),
  .A2({ S14176 }),
  .A3({ S25957[256] }),
  .A4({ S38 }),
  .ZN({ S14565 })
);
AOI21_X1 #() 
AOI21_X1_1028_ (
  .A({ S25957[260] }),
  .B1({ S14153 }),
  .B2({ S14565 }),
  .ZN({ S14566 })
);
NAND3_X1 #() 
NAND3_X1_1994_ (
  .A1({ S14150 }),
  .A2({ S14140 }),
  .A3({ S38 }),
  .ZN({ S14568 })
);
OAI21_X1 #() 
OAI21_X1_939_ (
  .A({ S14186 }),
  .B1({ S14568 }),
  .B2({ S14145 }),
  .ZN({ S14569 })
);
OAI22_X1 #() 
OAI22_X1_44_ (
  .A1({ S14564 }),
  .A2({ S14186 }),
  .B1({ S14566 }),
  .B2({ S14569 }),
  .ZN({ S14570 })
);
OAI21_X1 #() 
OAI21_X1_940_ (
  .A({ S25957[256] }),
  .B1({ S25957[258] }),
  .B2({ S14141 }),
  .ZN({ S14571 })
);
AOI21_X1 #() 
AOI21_X1_1029_ (
  .A({ S25957[260] }),
  .B1({ S14571 }),
  .B2({ S38 }),
  .ZN({ S14572 })
);
NAND2_X1 #() 
NAND2_X1_1715_ (
  .A1({ S14572 }),
  .A2({ S14282 }),
  .ZN({ S14573 })
);
NAND2_X1 #() 
NAND2_X1_1716_ (
  .A1({ S14177 }),
  .A2({ S25957[260] }),
  .ZN({ S14574 })
);
OAI21_X1 #() 
OAI21_X1_941_ (
  .A({ S14573 }),
  .B1({ S14247 }),
  .B2({ S14574 }),
  .ZN({ S14575 })
);
NAND2_X1 #() 
NAND2_X1_1717_ (
  .A1({ S14575 }),
  .A2({ S25957[261] }),
  .ZN({ S14576 })
);
NOR2_X1 #() 
NOR2_X1_400_ (
  .A1({ S14407 }),
  .A2({ S14416 }),
  .ZN({ S14577 })
);
OAI21_X1 #() 
OAI21_X1_942_ (
  .A({ S14145 }),
  .B1({ S14231 }),
  .B2({ S14577 }),
  .ZN({ S14579 })
);
NAND4_X1 #() 
NAND4_X1_251_ (
  .A1({ S14150 }),
  .A2({ S14156 }),
  .A3({ S14158 }),
  .A4({ S25957[259] }),
  .ZN({ S14580 })
);
NAND2_X1 #() 
NAND2_X1_1718_ (
  .A1({ S14320 }),
  .A2({ S14580 }),
  .ZN({ S14581 })
);
OAI211_X1 #() 
OAI211_X1_629_ (
  .A({ S14579 }),
  .B({ S14186 }),
  .C1({ S14145 }),
  .C2({ S14581 }),
  .ZN({ S14582 })
);
NAND3_X1 #() 
NAND3_X1_1995_ (
  .A1({ S14582 }),
  .A2({ S14576 }),
  .A3({ S14142 }),
  .ZN({ S14583 })
);
OAI21_X1 #() 
OAI21_X1_943_ (
  .A({ S14583 }),
  .B1({ S14570 }),
  .B2({ S14142 }),
  .ZN({ S14584 })
);
NAND2_X1 #() 
NAND2_X1_1719_ (
  .A1({ S14584 }),
  .A2({ S12121 }),
  .ZN({ S14585 })
);
NAND3_X1 #() 
NAND3_X1_1996_ (
  .A1({ S14561 }),
  .A2({ S14585 }),
  .A3({ S14529 }),
  .ZN({ S14586 })
);
NAND3_X1 #() 
NAND3_X1_1997_ (
  .A1({ S14559 }),
  .A2({ S14542 }),
  .A3({ S25957[263] }),
  .ZN({ S14587 })
);
OAI211_X1 #() 
OAI211_X1_630_ (
  .A({ S14587 }),
  .B({ S25957[459] }),
  .C1({ S14584 }),
  .C2({ S25957[263] }),
  .ZN({ S14588 })
);
AOI21_X1 #() 
AOI21_X1_1030_ (
  .A({ S25957[395] }),
  .B1({ S14586 }),
  .B2({ S14588 }),
  .ZN({ S14590 })
);
AND3_X1 #() 
AND3_X1_78_ (
  .A1({ S14586 }),
  .A2({ S25957[395] }),
  .A3({ S14588 }),
  .ZN({ S14591 })
);
NOR2_X1 #() 
NOR2_X1_401_ (
  .A1({ S14591 }),
  .A2({ S14590 }),
  .ZN({ S47 })
);
INV_X1 #() 
INV_X1_554_ (
  .A({ S47 }),
  .ZN({ S25957[139] })
);
NAND2_X1 #() 
NAND2_X1_1720_ (
  .A1({ S8834 }),
  .A2({ S8838 }),
  .ZN({ S25957[424] })
);
NAND2_X1 #() 
NAND2_X1_1721_ (
  .A1({ S11838 }),
  .A2({ S11839 }),
  .ZN({ S14592 })
);
XNOR2_X1 #() 
XNOR2_X1_58_ (
  .A({ S14592 }),
  .B({ S25957[424] }),
  .ZN({ S25957[296] })
);
NAND2_X1 #() 
NAND2_X1_1722_ (
  .A1({ S11835 }),
  .A2({ S11834 }),
  .ZN({ S25957[360] })
);
INV_X1 #() 
INV_X1_555_ (
  .A({ S25957[360] }),
  .ZN({ S14593 })
);
NAND3_X1 #() 
NAND3_X1_1998_ (
  .A1({ S14156 }),
  .A2({ S25957[259] }),
  .A3({ S25957[258] }),
  .ZN({ S14594 })
);
OAI21_X1 #() 
OAI21_X1_944_ (
  .A({ S14594 }),
  .B1({ S14181 }),
  .B2({ S14180 }),
  .ZN({ S14596 })
);
NAND3_X1 #() 
NAND3_X1_1999_ (
  .A1({ S14346 }),
  .A2({ S38 }),
  .A3({ S14428 }),
  .ZN({ S14597 })
);
AOI21_X1 #() 
AOI21_X1_1031_ (
  .A({ S25957[260] }),
  .B1({ S14152 }),
  .B2({ S25957[259] }),
  .ZN({ S14598 })
);
AOI22_X1 #() 
AOI22_X1_234_ (
  .A1({ S14597 }),
  .A2({ S14598 }),
  .B1({ S14596 }),
  .B2({ S25957[260] }),
  .ZN({ S14599 })
);
OAI21_X1 #() 
OAI21_X1_945_ (
  .A({ S14553 }),
  .B1({ S14533 }),
  .B2({ S25957[259] }),
  .ZN({ S14600 })
);
NAND3_X1 #() 
NAND3_X1_2000_ (
  .A1({ S14232 }),
  .A2({ S14178 }),
  .A3({ S14206 }),
  .ZN({ S14601 })
);
NAND2_X1 #() 
NAND2_X1_1723_ (
  .A1({ S14601 }),
  .A2({ S14208 }),
  .ZN({ S14602 })
);
OAI211_X1 #() 
OAI211_X1_631_ (
  .A({ S14186 }),
  .B({ S14602 }),
  .C1({ S14600 }),
  .C2({ S14145 }),
  .ZN({ S14603 })
);
OAI211_X1 #() 
OAI211_X1_632_ (
  .A({ S25957[262] }),
  .B({ S14603 }),
  .C1({ S14599 }),
  .C2({ S14186 }),
  .ZN({ S14604 })
);
AOI21_X1 #() 
AOI21_X1_1032_ (
  .A({ S25957[256] }),
  .B1({ S14225 }),
  .B2({ S14328 }),
  .ZN({ S14605 })
);
AOI21_X1 #() 
AOI21_X1_1033_ (
  .A({ S14605 }),
  .B1({ S14568 }),
  .B2({ S14177 }),
  .ZN({ S14607 })
);
NAND4_X1 #() 
NAND4_X1_252_ (
  .A1({ S14181 }),
  .A2({ S14395 }),
  .A3({ S14480 }),
  .A4({ S14145 }),
  .ZN({ S14608 })
);
OAI211_X1 #() 
OAI211_X1_633_ (
  .A({ S25957[261] }),
  .B({ S14608 }),
  .C1({ S14607 }),
  .C2({ S14145 }),
  .ZN({ S14609 })
);
INV_X1 #() 
INV_X1_556_ (
  .A({ S14309 }),
  .ZN({ S14610 })
);
AOI21_X1 #() 
AOI21_X1_1034_ (
  .A({ S14225 }),
  .B1({ S14156 }),
  .B2({ S14158 }),
  .ZN({ S14611 })
);
OAI21_X1 #() 
OAI21_X1_946_ (
  .A({ S25957[260] }),
  .B1({ S14610 }),
  .B2({ S14611 }),
  .ZN({ S14612 })
);
NAND4_X1 #() 
NAND4_X1_253_ (
  .A1({ S14147 }),
  .A2({ S14150 }),
  .A3({ S38 }),
  .A4({ S46 }),
  .ZN({ S14613 })
);
AOI21_X1 #() 
AOI21_X1_1035_ (
  .A({ S25957[261] }),
  .B1({ S14563 }),
  .B2({ S14613 }),
  .ZN({ S14614 })
);
AOI21_X1 #() 
AOI21_X1_1036_ (
  .A({ S25957[262] }),
  .B1({ S14614 }),
  .B2({ S14612 }),
  .ZN({ S14615 })
);
AOI21_X1 #() 
AOI21_X1_1037_ (
  .A({ S12121 }),
  .B1({ S14615 }),
  .B2({ S14609 }),
  .ZN({ S14616 })
);
NAND2_X1 #() 
NAND2_X1_1724_ (
  .A1({ S14604 }),
  .A2({ S14616 }),
  .ZN({ S14618 })
);
NAND4_X1 #() 
NAND4_X1_254_ (
  .A1({ S14215 }),
  .A2({ S14197 }),
  .A3({ S14188 }),
  .A4({ S25957[259] }),
  .ZN({ S14619 })
);
AOI21_X1 #() 
AOI21_X1_1038_ (
  .A({ S14145 }),
  .B1({ S14619 }),
  .B2({ S14335 }),
  .ZN({ S14620 })
);
NAND2_X1 #() 
NAND2_X1_1725_ (
  .A1({ S14194 }),
  .A2({ S14145 }),
  .ZN({ S14621 })
);
NOR2_X1 #() 
NOR2_X1_402_ (
  .A1({ S14327 }),
  .A2({ S14621 }),
  .ZN({ S14622 })
);
OAI21_X1 #() 
OAI21_X1_947_ (
  .A({ S25957[261] }),
  .B1({ S14620 }),
  .B2({ S14622 }),
  .ZN({ S14623 })
);
NAND3_X1 #() 
NAND3_X1_2001_ (
  .A1({ S46 }),
  .A2({ S14173 }),
  .A3({ S38 }),
  .ZN({ S14624 })
);
NAND3_X1 #() 
NAND3_X1_2002_ (
  .A1({ S14388 }),
  .A2({ S14145 }),
  .A3({ S14624 }),
  .ZN({ S14625 })
);
OAI21_X1 #() 
OAI21_X1_948_ (
  .A({ S14196 }),
  .B1({ S14160 }),
  .B2({ S25957[259] }),
  .ZN({ S14626 })
);
AND2_X1 #() 
AND2_X1_105_ (
  .A1({ S25957[260] }),
  .A2({ S14176 }),
  .ZN({ S14627 })
);
AOI21_X1 #() 
AOI21_X1_1039_ (
  .A({ S25957[261] }),
  .B1({ S14627 }),
  .B2({ S14626 }),
  .ZN({ S14629 })
);
NAND2_X1 #() 
NAND2_X1_1726_ (
  .A1({ S14629 }),
  .A2({ S14625 }),
  .ZN({ S14630 })
);
NAND3_X1 #() 
NAND3_X1_2003_ (
  .A1({ S14623 }),
  .A2({ S25957[262] }),
  .A3({ S14630 }),
  .ZN({ S14631 })
);
INV_X1 #() 
INV_X1_557_ (
  .A({ S14428 }),
  .ZN({ S14632 })
);
NAND3_X1 #() 
NAND3_X1_2004_ (
  .A1({ S14305 }),
  .A2({ S25957[259] }),
  .A3({ S46 }),
  .ZN({ S14633 })
);
OAI211_X1 #() 
OAI211_X1_634_ (
  .A({ S14633 }),
  .B({ S14145 }),
  .C1({ S14632 }),
  .C2({ S14181 }),
  .ZN({ S14634 })
);
NAND2_X1 #() 
NAND2_X1_1727_ (
  .A1({ S14150 }),
  .A2({ S14141 }),
  .ZN({ S14635 })
);
AOI21_X1 #() 
AOI21_X1_1040_ (
  .A({ S25957[259] }),
  .B1({ S14635 }),
  .B2({ S14305 }),
  .ZN({ S14636 })
);
OAI21_X1 #() 
OAI21_X1_949_ (
  .A({ S25957[260] }),
  .B1({ S14636 }),
  .B2({ S14551 }),
  .ZN({ S14637 })
);
AOI21_X1 #() 
AOI21_X1_1041_ (
  .A({ S25957[261] }),
  .B1({ S14637 }),
  .B2({ S14634 }),
  .ZN({ S14638 })
);
NAND3_X1 #() 
NAND3_X1_2005_ (
  .A1({ S14385 }),
  .A2({ S14494 }),
  .A3({ S25957[260] }),
  .ZN({ S14640 })
);
NAND3_X1 #() 
NAND3_X1_2006_ (
  .A1({ S14178 }),
  .A2({ S14278 }),
  .A3({ S14432 }),
  .ZN({ S14641 })
);
NAND3_X1 #() 
NAND3_X1_2007_ (
  .A1({ S14430 }),
  .A2({ S14641 }),
  .A3({ S14145 }),
  .ZN({ S14642 })
);
NAND3_X1 #() 
NAND3_X1_2008_ (
  .A1({ S14642 }),
  .A2({ S14640 }),
  .A3({ S25957[261] }),
  .ZN({ S14643 })
);
NAND2_X1 #() 
NAND2_X1_1728_ (
  .A1({ S14643 }),
  .A2({ S14142 }),
  .ZN({ S14644 })
);
OAI211_X1 #() 
OAI211_X1_635_ (
  .A({ S14631 }),
  .B({ S12121 }),
  .C1({ S14638 }),
  .C2({ S14644 }),
  .ZN({ S14645 })
);
NAND3_X1 #() 
NAND3_X1_2009_ (
  .A1({ S14645 }),
  .A2({ S14593 }),
  .A3({ S14618 }),
  .ZN({ S14646 })
);
AND2_X1 #() 
AND2_X1_106_ (
  .A1({ S14604 }),
  .A2({ S14616 }),
  .ZN({ S14647 })
);
NOR2_X1 #() 
NOR2_X1_403_ (
  .A1({ S14333 }),
  .A2({ S25957[256] }),
  .ZN({ S14648 })
);
AOI21_X1 #() 
AOI21_X1_1042_ (
  .A({ S38 }),
  .B1({ S14230 }),
  .B2({ S14155 }),
  .ZN({ S14649 })
);
OAI21_X1 #() 
OAI21_X1_950_ (
  .A({ S25957[260] }),
  .B1({ S14649 }),
  .B2({ S14648 }),
  .ZN({ S14651 })
);
INV_X1 #() 
INV_X1_558_ (
  .A({ S14327 }),
  .ZN({ S14652 })
);
NAND2_X1 #() 
NAND2_X1_1729_ (
  .A1({ S14652 }),
  .A2({ S14208 }),
  .ZN({ S14653 })
);
NAND2_X1 #() 
NAND2_X1_1730_ (
  .A1({ S14651 }),
  .A2({ S14653 }),
  .ZN({ S14654 })
);
NAND2_X1 #() 
NAND2_X1_1731_ (
  .A1({ S14630 }),
  .A2({ S25957[262] }),
  .ZN({ S14655 })
);
AOI21_X1 #() 
AOI21_X1_1043_ (
  .A({ S14655 }),
  .B1({ S14654 }),
  .B2({ S25957[261] }),
  .ZN({ S14656 })
);
OAI21_X1 #() 
OAI21_X1_951_ (
  .A({ S12121 }),
  .B1({ S14638 }),
  .B2({ S14644 }),
  .ZN({ S14657 })
);
NOR2_X1 #() 
NOR2_X1_404_ (
  .A1({ S14657 }),
  .A2({ S14656 }),
  .ZN({ S14658 })
);
OAI21_X1 #() 
OAI21_X1_952_ (
  .A({ S25957[360] }),
  .B1({ S14658 }),
  .B2({ S14647 }),
  .ZN({ S14659 })
);
AOI21_X1 #() 
AOI21_X1_1044_ (
  .A({ S14592 }),
  .B1({ S14659 }),
  .B2({ S14646 }),
  .ZN({ S14660 })
);
INV_X1 #() 
INV_X1_559_ (
  .A({ S14592 }),
  .ZN({ S25957[328] })
);
NAND3_X1 #() 
NAND3_X1_2010_ (
  .A1({ S14645 }),
  .A2({ S25957[360] }),
  .A3({ S14618 }),
  .ZN({ S14662 })
);
OAI21_X1 #() 
OAI21_X1_953_ (
  .A({ S14593 }),
  .B1({ S14658 }),
  .B2({ S14647 }),
  .ZN({ S14663 })
);
AOI21_X1 #() 
AOI21_X1_1045_ (
  .A({ S25957[328] }),
  .B1({ S14663 }),
  .B2({ S14662 }),
  .ZN({ S14664 })
);
OAI21_X1 #() 
OAI21_X1_954_ (
  .A({ S25957[296] }),
  .B1({ S14660 }),
  .B2({ S14664 }),
  .ZN({ S14665 })
);
INV_X1 #() 
INV_X1_560_ (
  .A({ S25957[296] }),
  .ZN({ S14666 })
);
NAND3_X1 #() 
NAND3_X1_2011_ (
  .A1({ S14663 }),
  .A2({ S14662 }),
  .A3({ S25957[328] }),
  .ZN({ S14667 })
);
NAND3_X1 #() 
NAND3_X1_2012_ (
  .A1({ S14659 }),
  .A2({ S14646 }),
  .A3({ S14592 }),
  .ZN({ S14668 })
);
NAND3_X1 #() 
NAND3_X1_2013_ (
  .A1({ S14667 }),
  .A2({ S14668 }),
  .A3({ S14666 }),
  .ZN({ S14669 })
);
NAND3_X1 #() 
NAND3_X1_2014_ (
  .A1({ S14665 }),
  .A2({ S25957[264] }),
  .A3({ S14669 }),
  .ZN({ S14670 })
);
NAND3_X1 #() 
NAND3_X1_2015_ (
  .A1({ S14667 }),
  .A2({ S14668 }),
  .A3({ S25957[296] }),
  .ZN({ S14672 })
);
OAI21_X1 #() 
OAI21_X1_955_ (
  .A({ S14666 }),
  .B1({ S14660 }),
  .B2({ S14664 }),
  .ZN({ S14673 })
);
NAND3_X1 #() 
NAND3_X1_2016_ (
  .A1({ S14673 }),
  .A2({ S13424 }),
  .A3({ S14672 }),
  .ZN({ S14674 })
);
NAND2_X1 #() 
NAND2_X1_1732_ (
  .A1({ S14670 }),
  .A2({ S14674 }),
  .ZN({ S25957[136] })
);
NOR2_X1 #() 
NOR2_X1_405_ (
  .A1({ S11883 }),
  .A2({ S11884 }),
  .ZN({ S25957[329] })
);
NAND2_X1 #() 
NAND2_X1_1733_ (
  .A1({ S8936 }),
  .A2({ S8935 }),
  .ZN({ S25957[489] })
);
XNOR2_X1 #() 
XNOR2_X1_59_ (
  .A({ S11888 }),
  .B({ S25957[489] }),
  .ZN({ S25957[361] })
);
NAND3_X1 #() 
NAND3_X1_2017_ (
  .A1({ S14375 }),
  .A2({ S14225 }),
  .A3({ S14226 }),
  .ZN({ S14675 })
);
AOI21_X1 #() 
AOI21_X1_1046_ (
  .A({ S25957[260] }),
  .B1({ S14371 }),
  .B2({ S14205 }),
  .ZN({ S14676 })
);
AOI22_X1 #() 
AOI22_X1_235_ (
  .A1({ S14676 }),
  .A2({ S14619 }),
  .B1({ S14675 }),
  .B2({ S25957[260] }),
  .ZN({ S14677 })
);
INV_X1 #() 
INV_X1_561_ (
  .A({ S14605 }),
  .ZN({ S14679 })
);
OAI211_X1 #() 
OAI211_X1_636_ (
  .A({ S25957[260] }),
  .B({ S14679 }),
  .C1({ S14246 }),
  .C2({ S14382 }),
  .ZN({ S14680 })
);
NAND3_X1 #() 
NAND3_X1_2018_ (
  .A1({ S14278 }),
  .A2({ S14140 }),
  .A3({ S25957[259] }),
  .ZN({ S14681 })
);
OAI211_X1 #() 
OAI211_X1_637_ (
  .A({ S14145 }),
  .B({ S14681 }),
  .C1({ S14568 }),
  .C2({ S14404 }),
  .ZN({ S14682 })
);
NAND3_X1 #() 
NAND3_X1_2019_ (
  .A1({ S14680 }),
  .A2({ S14186 }),
  .A3({ S14682 }),
  .ZN({ S14683 })
);
OAI211_X1 #() 
OAI211_X1_638_ (
  .A({ S14683 }),
  .B({ S25957[262] }),
  .C1({ S14186 }),
  .C2({ S14677 }),
  .ZN({ S14684 })
);
NOR2_X1 #() 
NOR2_X1_406_ (
  .A1({ S14471 }),
  .A2({ S14233 }),
  .ZN({ S14685 })
);
AOI21_X1 #() 
AOI21_X1_1047_ (
  .A({ S38 }),
  .B1({ S14230 }),
  .B2({ S14147 }),
  .ZN({ S14686 })
);
NAND3_X1 #() 
NAND3_X1_2020_ (
  .A1({ S14562 }),
  .A2({ S14145 }),
  .A3({ S14304 }),
  .ZN({ S14687 })
);
OAI211_X1 #() 
OAI211_X1_639_ (
  .A({ S14687 }),
  .B({ S25957[261] }),
  .C1({ S14218 }),
  .C2({ S14686 }),
  .ZN({ S14688 })
);
AOI21_X1 #() 
AOI21_X1_1048_ (
  .A({ S25957[259] }),
  .B1({ S14326 }),
  .B2({ S14162 }),
  .ZN({ S14690 })
);
OAI21_X1 #() 
OAI21_X1_956_ (
  .A({ S14186 }),
  .B1({ S14690 }),
  .B2({ S14288 }),
  .ZN({ S14691 })
);
OAI211_X1 #() 
OAI211_X1_640_ (
  .A({ S14142 }),
  .B({ S14688 }),
  .C1({ S14685 }),
  .C2({ S14691 }),
  .ZN({ S14692 })
);
NAND3_X1 #() 
NAND3_X1_2021_ (
  .A1({ S14692 }),
  .A2({ S14684 }),
  .A3({ S25957[263] }),
  .ZN({ S14693 })
);
OAI211_X1 #() 
OAI211_X1_641_ (
  .A({ S14580 }),
  .B({ S25957[260] }),
  .C1({ S14181 }),
  .C2({ S14294 }),
  .ZN({ S14694 })
);
NAND4_X1 #() 
NAND4_X1_255_ (
  .A1({ S14405 }),
  .A2({ S14191 }),
  .A3({ S14150 }),
  .A4({ S14145 }),
  .ZN({ S14695 })
);
NAND3_X1 #() 
NAND3_X1_2022_ (
  .A1({ S14694 }),
  .A2({ S14695 }),
  .A3({ S25957[261] }),
  .ZN({ S14696 })
);
NAND2_X1 #() 
NAND2_X1_1734_ (
  .A1({ S14492 }),
  .A2({ S14227 }),
  .ZN({ S14697 })
);
AOI21_X1 #() 
AOI21_X1_1049_ (
  .A({ S14145 }),
  .B1({ S14697 }),
  .B2({ S14619 }),
  .ZN({ S14698 })
);
NAND3_X1 #() 
NAND3_X1_2023_ (
  .A1({ S14342 }),
  .A2({ S14145 }),
  .A3({ S14553 }),
  .ZN({ S14699 })
);
NAND2_X1 #() 
NAND2_X1_1735_ (
  .A1({ S14699 }),
  .A2({ S14186 }),
  .ZN({ S14701 })
);
OAI21_X1 #() 
OAI21_X1_957_ (
  .A({ S14696 }),
  .B1({ S14698 }),
  .B2({ S14701 }),
  .ZN({ S14702 })
);
AOI21_X1 #() 
AOI21_X1_1050_ (
  .A({ S14145 }),
  .B1({ S14544 }),
  .B2({ S14458 }),
  .ZN({ S14703 })
);
OAI21_X1 #() 
OAI21_X1_958_ (
  .A({ S25957[261] }),
  .B1({ S14703 }),
  .B2({ S14239 }),
  .ZN({ S14704 })
);
NOR2_X1 #() 
NOR2_X1_407_ (
  .A1({ S14371 }),
  .A2({ S14333 }),
  .ZN({ S14705 })
);
OAI21_X1 #() 
OAI21_X1_959_ (
  .A({ S25957[260] }),
  .B1({ S14705 }),
  .B2({ S14203 }),
  .ZN({ S14706 })
);
INV_X1 #() 
INV_X1_562_ (
  .A({ S14565 }),
  .ZN({ S14707 })
);
OAI21_X1 #() 
OAI21_X1_960_ (
  .A({ S14145 }),
  .B1({ S14707 }),
  .B2({ S14192 }),
  .ZN({ S14708 })
);
NAND2_X1 #() 
NAND2_X1_1736_ (
  .A1({ S14708 }),
  .A2({ S14706 }),
  .ZN({ S14709 })
);
NAND2_X1 #() 
NAND2_X1_1737_ (
  .A1({ S14709 }),
  .A2({ S14186 }),
  .ZN({ S14710 })
);
NAND3_X1 #() 
NAND3_X1_2024_ (
  .A1({ S14710 }),
  .A2({ S14142 }),
  .A3({ S14704 }),
  .ZN({ S14712 })
);
OAI211_X1 #() 
OAI211_X1_642_ (
  .A({ S14712 }),
  .B({ S12121 }),
  .C1({ S14142 }),
  .C2({ S14702 }),
  .ZN({ S14713 })
);
NAND3_X1 #() 
NAND3_X1_2025_ (
  .A1({ S14713 }),
  .A2({ S14693 }),
  .A3({ S25957[361] }),
  .ZN({ S14714 })
);
INV_X1 #() 
INV_X1_563_ (
  .A({ S25957[361] }),
  .ZN({ S14715 })
);
NAND2_X1 #() 
NAND2_X1_1738_ (
  .A1({ S14702 }),
  .A2({ S25957[262] }),
  .ZN({ S14716 })
);
OAI21_X1 #() 
OAI21_X1_961_ (
  .A({ S25957[261] }),
  .B1({ S14238 }),
  .B2({ S25957[260] }),
  .ZN({ S14717 })
);
OAI221_X1 #() 
OAI221_X1_38_ (
  .A({ S14142 }),
  .B1({ S14717 }),
  .B2({ S14703 }),
  .C1({ S14709 }),
  .C2({ S25957[261] }),
  .ZN({ S14718 })
);
NAND3_X1 #() 
NAND3_X1_2026_ (
  .A1({ S14716 }),
  .A2({ S14718 }),
  .A3({ S12121 }),
  .ZN({ S14719 })
);
OAI21_X1 #() 
OAI21_X1_962_ (
  .A({ S14683 }),
  .B1({ S14186 }),
  .B2({ S14677 }),
  .ZN({ S14720 })
);
NAND2_X1 #() 
NAND2_X1_1739_ (
  .A1({ S14720 }),
  .A2({ S25957[262] }),
  .ZN({ S14721 })
);
OAI21_X1 #() 
OAI21_X1_963_ (
  .A({ S14687 }),
  .B1({ S14218 }),
  .B2({ S14686 }),
  .ZN({ S14723 })
);
NAND2_X1 #() 
NAND2_X1_1740_ (
  .A1({ S14723 }),
  .A2({ S25957[261] }),
  .ZN({ S14724 })
);
NOR2_X1 #() 
NOR2_X1_408_ (
  .A1({ S14151 }),
  .A2({ S38 }),
  .ZN({ S14725 })
);
OAI21_X1 #() 
OAI21_X1_964_ (
  .A({ S25957[260] }),
  .B1({ S14690 }),
  .B2({ S14725 }),
  .ZN({ S14726 })
);
OAI21_X1 #() 
OAI21_X1_965_ (
  .A({ S14145 }),
  .B1({ S14233 }),
  .B2({ S14470 }),
  .ZN({ S14727 })
);
NAND3_X1 #() 
NAND3_X1_2027_ (
  .A1({ S14727 }),
  .A2({ S14726 }),
  .A3({ S14186 }),
  .ZN({ S14728 })
);
NAND3_X1 #() 
NAND3_X1_2028_ (
  .A1({ S14724 }),
  .A2({ S14142 }),
  .A3({ S14728 }),
  .ZN({ S14729 })
);
NAND3_X1 #() 
NAND3_X1_2029_ (
  .A1({ S14721 }),
  .A2({ S25957[263] }),
  .A3({ S14729 }),
  .ZN({ S14730 })
);
NAND3_X1 #() 
NAND3_X1_2030_ (
  .A1({ S14730 }),
  .A2({ S14719 }),
  .A3({ S14715 }),
  .ZN({ S14731 })
);
NAND3_X1 #() 
NAND3_X1_2031_ (
  .A1({ S14731 }),
  .A2({ S14714 }),
  .A3({ S25957[329] }),
  .ZN({ S14732 })
);
INV_X1 #() 
INV_X1_564_ (
  .A({ S25957[329] }),
  .ZN({ S14734 })
);
NAND3_X1 #() 
NAND3_X1_2032_ (
  .A1({ S14713 }),
  .A2({ S14693 }),
  .A3({ S14715 }),
  .ZN({ S14735 })
);
NAND3_X1 #() 
NAND3_X1_2033_ (
  .A1({ S14730 }),
  .A2({ S14719 }),
  .A3({ S25957[361] }),
  .ZN({ S14736 })
);
NAND3_X1 #() 
NAND3_X1_2034_ (
  .A1({ S14736 }),
  .A2({ S14735 }),
  .A3({ S14734 }),
  .ZN({ S14737 })
);
NAND3_X1 #() 
NAND3_X1_2035_ (
  .A1({ S14732 }),
  .A2({ S14737 }),
  .A3({ S10516 }),
  .ZN({ S14738 })
);
NAND3_X1 #() 
NAND3_X1_2036_ (
  .A1({ S14731 }),
  .A2({ S14714 }),
  .A3({ S14734 }),
  .ZN({ S14739 })
);
NAND3_X1 #() 
NAND3_X1_2037_ (
  .A1({ S14736 }),
  .A2({ S14735 }),
  .A3({ S25957[329] }),
  .ZN({ S14740 })
);
NAND3_X1 #() 
NAND3_X1_2038_ (
  .A1({ S14739 }),
  .A2({ S14740 }),
  .A3({ S25957[393] }),
  .ZN({ S14741 })
);
NAND2_X1 #() 
NAND2_X1_1741_ (
  .A1({ S14738 }),
  .A2({ S14741 }),
  .ZN({ S25957[137] })
);
NAND2_X1 #() 
NAND2_X1_1742_ (
  .A1({ S9038 }),
  .A2({ S9039 }),
  .ZN({ S25957[458] })
);
XNOR2_X1 #() 
XNOR2_X1_60_ (
  .A({ S25957[458] }),
  .B({ S25957[554] }),
  .ZN({ S14743 })
);
NAND2_X1 #() 
NAND2_X1_1743_ (
  .A1({ S11968 }),
  .A2({ S11967 }),
  .ZN({ S14744 })
);
INV_X1 #() 
INV_X1_565_ (
  .A({ S14744 }),
  .ZN({ S25957[362] })
);
INV_X1 #() 
INV_X1_566_ (
  .A({ S14188 }),
  .ZN({ S14745 })
);
OAI211_X1 #() 
OAI211_X1_643_ (
  .A({ S14163 }),
  .B({ S14145 }),
  .C1({ S14745 }),
  .C2({ S14373 }),
  .ZN({ S14746 })
);
NAND3_X1 #() 
NAND3_X1_2039_ (
  .A1({ S14173 }),
  .A2({ S25957[256] }),
  .A3({ S25957[259] }),
  .ZN({ S14747 })
);
NAND3_X1 #() 
NAND3_X1_2040_ (
  .A1({ S14565 }),
  .A2({ S25957[260] }),
  .A3({ S14747 }),
  .ZN({ S14748 })
);
NAND3_X1 #() 
NAND3_X1_2041_ (
  .A1({ S14746 }),
  .A2({ S14748 }),
  .A3({ S25957[261] }),
  .ZN({ S14749 })
);
NOR2_X1 #() 
NOR2_X1_409_ (
  .A1({ S14346 }),
  .A2({ S38 }),
  .ZN({ S14750 })
);
OAI211_X1 #() 
OAI211_X1_644_ (
  .A({ S14309 }),
  .B({ S14145 }),
  .C1({ S14206 }),
  .C2({ S14147 }),
  .ZN({ S14751 })
);
OAI21_X1 #() 
OAI21_X1_966_ (
  .A({ S25957[260] }),
  .B1({ S14160 }),
  .B2({ S25957[259] }),
  .ZN({ S14753 })
);
OAI211_X1 #() 
OAI211_X1_645_ (
  .A({ S14751 }),
  .B({ S14186 }),
  .C1({ S14750 }),
  .C2({ S14753 }),
  .ZN({ S14754 })
);
NAND3_X1 #() 
NAND3_X1_2042_ (
  .A1({ S14749 }),
  .A2({ S14142 }),
  .A3({ S14754 }),
  .ZN({ S14755 })
);
NAND2_X1 #() 
NAND2_X1_1744_ (
  .A1({ S14508 }),
  .A2({ S25957[259] }),
  .ZN({ S14756 })
);
NAND3_X1 #() 
NAND3_X1_2043_ (
  .A1({ S14756 }),
  .A2({ S14145 }),
  .A3({ S14254 }),
  .ZN({ S14757 })
);
OAI21_X1 #() 
OAI21_X1_967_ (
  .A({ S38 }),
  .B1({ S14632 }),
  .B2({ S14543 }),
  .ZN({ S14758 })
);
AOI21_X1 #() 
AOI21_X1_1051_ (
  .A({ S14145 }),
  .B1({ S14161 }),
  .B2({ S14150 }),
  .ZN({ S14759 })
);
AOI21_X1 #() 
AOI21_X1_1052_ (
  .A({ S14186 }),
  .B1({ S14758 }),
  .B2({ S14759 }),
  .ZN({ S14760 })
);
NAND2_X1 #() 
NAND2_X1_1745_ (
  .A1({ S14760 }),
  .A2({ S14757 }),
  .ZN({ S14761 })
);
NAND2_X1 #() 
NAND2_X1_1746_ (
  .A1({ S14412 }),
  .A2({ S14154 }),
  .ZN({ S14762 })
);
NAND2_X1 #() 
NAND2_X1_1747_ (
  .A1({ S14462 }),
  .A2({ S14762 }),
  .ZN({ S14764 })
);
NAND2_X1 #() 
NAND2_X1_1748_ (
  .A1({ S14187 }),
  .A2({ S14188 }),
  .ZN({ S14765 })
);
NAND2_X1 #() 
NAND2_X1_1749_ (
  .A1({ S14765 }),
  .A2({ S25957[259] }),
  .ZN({ S14766 })
);
NAND2_X1 #() 
NAND2_X1_1750_ (
  .A1({ S14766 }),
  .A2({ S14414 }),
  .ZN({ S14767 })
);
NAND3_X1 #() 
NAND3_X1_2044_ (
  .A1({ S14767 }),
  .A2({ S14764 }),
  .A3({ S14186 }),
  .ZN({ S14768 })
);
NAND3_X1 #() 
NAND3_X1_2045_ (
  .A1({ S14761 }),
  .A2({ S14768 }),
  .A3({ S25957[262] }),
  .ZN({ S14769 })
);
NAND3_X1 #() 
NAND3_X1_2046_ (
  .A1({ S14769 }),
  .A2({ S25957[263] }),
  .A3({ S14755 }),
  .ZN({ S14770 })
);
OAI211_X1 #() 
OAI211_X1_646_ (
  .A({ S14150 }),
  .B({ S25957[259] }),
  .C1({ S14156 }),
  .C2({ S25957[258] }),
  .ZN({ S14771 })
);
NAND3_X1 #() 
NAND3_X1_2047_ (
  .A1({ S14771 }),
  .A2({ S14568 }),
  .A3({ S14372 }),
  .ZN({ S14772 })
);
NAND2_X1 #() 
NAND2_X1_1751_ (
  .A1({ S14533 }),
  .A2({ S38 }),
  .ZN({ S14773 })
);
AOI21_X1 #() 
AOI21_X1_1053_ (
  .A({ S25957[260] }),
  .B1({ S14543 }),
  .B2({ S25957[259] }),
  .ZN({ S14775 })
);
AOI22_X1 #() 
AOI22_X1_236_ (
  .A1({ S14772 }),
  .A2({ S25957[260] }),
  .B1({ S14773 }),
  .B2({ S14775 }),
  .ZN({ S14776 })
);
NAND2_X1 #() 
NAND2_X1_1752_ (
  .A1({ S14333 }),
  .A2({ S14191 }),
  .ZN({ S14777 })
);
AND3_X1 #() 
AND3_X1_79_ (
  .A1({ S14278 }),
  .A2({ S25957[260] }),
  .A3({ S14156 }),
  .ZN({ S14778 })
);
AOI22_X1 #() 
AOI22_X1_237_ (
  .A1({ S14198 }),
  .A2({ S14572 }),
  .B1({ S14778 }),
  .B2({ S14777 }),
  .ZN({ S14779 })
);
NAND2_X1 #() 
NAND2_X1_1753_ (
  .A1({ S14779 }),
  .A2({ S25957[261] }),
  .ZN({ S14780 })
);
OAI211_X1 #() 
OAI211_X1_647_ (
  .A({ S14780 }),
  .B({ S25957[262] }),
  .C1({ S25957[261] }),
  .C2({ S14776 }),
  .ZN({ S14781 })
);
NAND3_X1 #() 
NAND3_X1_2048_ (
  .A1({ S14155 }),
  .A2({ S14305 }),
  .A3({ S25957[259] }),
  .ZN({ S14782 })
);
NAND3_X1 #() 
NAND3_X1_2049_ (
  .A1({ S14782 }),
  .A2({ S14145 }),
  .A3({ S14310 }),
  .ZN({ S14783 })
);
OAI211_X1 #() 
OAI211_X1_648_ (
  .A({ S14150 }),
  .B({ S25957[259] }),
  .C1({ S25957[256] }),
  .C2({ S14173 }),
  .ZN({ S14784 })
);
NAND3_X1 #() 
NAND3_X1_2050_ (
  .A1({ S14546 }),
  .A2({ S25957[260] }),
  .A3({ S14784 }),
  .ZN({ S14786 })
);
NAND3_X1 #() 
NAND3_X1_2051_ (
  .A1({ S14786 }),
  .A2({ S14783 }),
  .A3({ S25957[261] }),
  .ZN({ S14787 })
);
NAND3_X1 #() 
NAND3_X1_2052_ (
  .A1({ S14652 }),
  .A2({ S14145 }),
  .A3({ S14597 }),
  .ZN({ S14788 })
);
AOI21_X1 #() 
AOI21_X1_1054_ (
  .A({ S14145 }),
  .B1({ S14543 }),
  .B2({ S25957[259] }),
  .ZN({ S14789 })
);
AOI21_X1 #() 
AOI21_X1_1055_ (
  .A({ S25957[261] }),
  .B1({ S14474 }),
  .B2({ S14789 }),
  .ZN({ S14790 })
);
NAND2_X1 #() 
NAND2_X1_1754_ (
  .A1({ S14788 }),
  .A2({ S14790 }),
  .ZN({ S14791 })
);
NAND3_X1 #() 
NAND3_X1_2053_ (
  .A1({ S14791 }),
  .A2({ S14787 }),
  .A3({ S14142 }),
  .ZN({ S14792 })
);
NAND3_X1 #() 
NAND3_X1_2054_ (
  .A1({ S14781 }),
  .A2({ S12121 }),
  .A3({ S14792 }),
  .ZN({ S14793 })
);
NAND3_X1 #() 
NAND3_X1_2055_ (
  .A1({ S14793 }),
  .A2({ S14770 }),
  .A3({ S25957[362] }),
  .ZN({ S14794 })
);
AOI22_X1 #() 
AOI22_X1_238_ (
  .A1({ S14766 }),
  .A2({ S14414 }),
  .B1({ S14462 }),
  .B2({ S14762 }),
  .ZN({ S14795 })
);
AOI22_X1 #() 
AOI22_X1_239_ (
  .A1({ S14795 }),
  .A2({ S14186 }),
  .B1({ S14760 }),
  .B2({ S14757 }),
  .ZN({ S14797 })
);
NAND2_X1 #() 
NAND2_X1_1755_ (
  .A1({ S14749 }),
  .A2({ S14754 }),
  .ZN({ S14798 })
);
NAND2_X1 #() 
NAND2_X1_1756_ (
  .A1({ S14798 }),
  .A2({ S14142 }),
  .ZN({ S14799 })
);
OAI211_X1 #() 
OAI211_X1_649_ (
  .A({ S14799 }),
  .B({ S25957[263] }),
  .C1({ S14797 }),
  .C2({ S14142 }),
  .ZN({ S14800 })
);
NAND2_X1 #() 
NAND2_X1_1757_ (
  .A1({ S14772 }),
  .A2({ S25957[260] }),
  .ZN({ S14801 })
);
NAND2_X1 #() 
NAND2_X1_1758_ (
  .A1({ S14773 }),
  .A2({ S14775 }),
  .ZN({ S14802 })
);
AOI21_X1 #() 
AOI21_X1_1056_ (
  .A({ S25957[261] }),
  .B1({ S14801 }),
  .B2({ S14802 }),
  .ZN({ S14803 })
);
NAND2_X1 #() 
NAND2_X1_1759_ (
  .A1({ S14198 }),
  .A2({ S14572 }),
  .ZN({ S14804 })
);
NAND2_X1 #() 
NAND2_X1_1760_ (
  .A1({ S14778 }),
  .A2({ S14777 }),
  .ZN({ S14805 })
);
AND3_X1 #() 
AND3_X1_80_ (
  .A1({ S14804 }),
  .A2({ S25957[261] }),
  .A3({ S14805 }),
  .ZN({ S14806 })
);
OAI21_X1 #() 
OAI21_X1_968_ (
  .A({ S25957[262] }),
  .B1({ S14806 }),
  .B2({ S14803 }),
  .ZN({ S14808 })
);
NAND2_X1 #() 
NAND2_X1_1761_ (
  .A1({ S14791 }),
  .A2({ S14787 }),
  .ZN({ S14809 })
);
NAND2_X1 #() 
NAND2_X1_1762_ (
  .A1({ S14809 }),
  .A2({ S14142 }),
  .ZN({ S14810 })
);
NAND3_X1 #() 
NAND3_X1_2056_ (
  .A1({ S14810 }),
  .A2({ S14808 }),
  .A3({ S12121 }),
  .ZN({ S14811 })
);
NAND3_X1 #() 
NAND3_X1_2057_ (
  .A1({ S14811 }),
  .A2({ S14744 }),
  .A3({ S14800 }),
  .ZN({ S14812 })
);
AOI21_X1 #() 
AOI21_X1_1057_ (
  .A({ S14743 }),
  .B1({ S14812 }),
  .B2({ S14794 }),
  .ZN({ S14813 })
);
INV_X1 #() 
INV_X1_567_ (
  .A({ S14743 }),
  .ZN({ S25957[426] })
);
NAND3_X1 #() 
NAND3_X1_2058_ (
  .A1({ S14793 }),
  .A2({ S14770 }),
  .A3({ S14744 }),
  .ZN({ S14814 })
);
NAND3_X1 #() 
NAND3_X1_2059_ (
  .A1({ S14811 }),
  .A2({ S25957[362] }),
  .A3({ S14800 }),
  .ZN({ S14815 })
);
AOI21_X1 #() 
AOI21_X1_1058_ (
  .A({ S25957[426] }),
  .B1({ S14815 }),
  .B2({ S14814 }),
  .ZN({ S14816 })
);
OAI21_X1 #() 
OAI21_X1_969_ (
  .A({ S13416 }),
  .B1({ S14813 }),
  .B2({ S14816 }),
  .ZN({ S14818 })
);
NAND3_X1 #() 
NAND3_X1_2060_ (
  .A1({ S14815 }),
  .A2({ S25957[426] }),
  .A3({ S14814 }),
  .ZN({ S14819 })
);
NAND3_X1 #() 
NAND3_X1_2061_ (
  .A1({ S14812 }),
  .A2({ S14743 }),
  .A3({ S14794 }),
  .ZN({ S14820 })
);
NAND3_X1 #() 
NAND3_X1_2062_ (
  .A1({ S14819 }),
  .A2({ S14820 }),
  .A3({ S25957[266] }),
  .ZN({ S14821 })
);
NAND2_X1 #() 
NAND2_X1_1763_ (
  .A1({ S14818 }),
  .A2({ S14821 }),
  .ZN({ S25957[138] })
);
AOI22_X1 #() 
AOI22_X1_240_ (
  .A1({ S13318 }),
  .A2({ S13321 }),
  .B1({ S13209 }),
  .B2({ S13239 }),
  .ZN({ S48 })
);
NAND4_X1 #() 
NAND4_X1_256_ (
  .A1({ S13318 }),
  .A2({ S13209 }),
  .A3({ S13239 }),
  .A4({ S13321 }),
  .ZN({ S49 })
);
NOR2_X1 #() 
NOR2_X1_410_ (
  .A1({ S12115 }),
  .A2({ S12116 }),
  .ZN({ S25957[295] })
);
NAND2_X1 #() 
NAND2_X1_1764_ (
  .A1({ S12803 }),
  .A2({ S12801 }),
  .ZN({ S14822 })
);
INV_X1 #() 
INV_X1_568_ (
  .A({ S25957[286] }),
  .ZN({ S14823 })
);
AOI21_X1 #() 
AOI21_X1_1059_ (
  .A({ S7386 }),
  .B1({ S13237 }),
  .B2({ S13210 }),
  .ZN({ S14825 })
);
NOR3_X1 #() 
NOR3_X1_60_ (
  .A1({ S13207 }),
  .A2({ S13208 }),
  .A3({ S25957[536] }),
  .ZN({ S14826 })
);
OAI21_X1 #() 
OAI21_X1_970_ (
  .A({ S25957[282] }),
  .B1({ S14826 }),
  .B2({ S14825 }),
  .ZN({ S14827 })
);
AOI21_X1 #() 
AOI21_X1_1060_ (
  .A({ S9169 }),
  .B1({ S13320 }),
  .B2({ S13319 }),
  .ZN({ S14828 })
);
AND3_X1 #() 
AND3_X1_81_ (
  .A1({ S13320 }),
  .A2({ S13319 }),
  .A3({ S9169 }),
  .ZN({ S14829 })
);
OAI21_X1 #() 
OAI21_X1_971_ (
  .A({ S25957[282] }),
  .B1({ S14829 }),
  .B2({ S14828 }),
  .ZN({ S14830 })
);
NAND2_X1 #() 
NAND2_X1_1765_ (
  .A1({ S14830 }),
  .A2({ S14827 }),
  .ZN({ S14831 })
);
OAI21_X1 #() 
OAI21_X1_972_ (
  .A({ S3488 }),
  .B1({ S13383 }),
  .B2({ S13371 }),
  .ZN({ S14832 })
);
NAND3_X1 #() 
NAND3_X1_2063_ (
  .A1({ S13369 }),
  .A2({ S25957[794] }),
  .A3({ S13344 }),
  .ZN({ S14833 })
);
NAND2_X1 #() 
NAND2_X1_1766_ (
  .A1({ S14832 }),
  .A2({ S14833 }),
  .ZN({ S14834 })
);
NAND3_X1 #() 
NAND3_X1_2064_ (
  .A1({ S13318 }),
  .A2({ S13321 }),
  .A3({ S14834 }),
  .ZN({ S14836 })
);
NAND3_X1 #() 
NAND3_X1_2065_ (
  .A1({ S14834 }),
  .A2({ S13209 }),
  .A3({ S13239 }),
  .ZN({ S14837 })
);
NAND2_X1 #() 
NAND2_X1_1767_ (
  .A1({ S14836 }),
  .A2({ S14837 }),
  .ZN({ S14838 })
);
NOR2_X1 #() 
NOR2_X1_411_ (
  .A1({ S14831 }),
  .A2({ S14838 }),
  .ZN({ S14839 })
);
NOR2_X1 #() 
NOR2_X1_412_ (
  .A1({ S14839 }),
  .A2({ S41 }),
  .ZN({ S14840 })
);
NOR2_X1 #() 
NOR2_X1_413_ (
  .A1({ S14829 }),
  .A2({ S14828 }),
  .ZN({ S14841 })
);
NAND4_X1 #() 
NAND4_X1_257_ (
  .A1({ S13209 }),
  .A2({ S13239 }),
  .A3({ S14832 }),
  .A4({ S14833 }),
  .ZN({ S14842 })
);
OAI211_X1 #() 
OAI211_X1_650_ (
  .A({ S41 }),
  .B({ S14837 }),
  .C1({ S14841 }),
  .C2({ S14842 }),
  .ZN({ S14843 })
);
NAND2_X1 #() 
NAND2_X1_1768_ (
  .A1({ S14843 }),
  .A2({ S25957[284] }),
  .ZN({ S14844 })
);
NAND3_X1 #() 
NAND3_X1_2066_ (
  .A1({ S25957[282] }),
  .A2({ S13318 }),
  .A3({ S13321 }),
  .ZN({ S14845 })
);
INV_X1 #() 
INV_X1_569_ (
  .A({ S14845 }),
  .ZN({ S14847 })
);
NAND2_X1 #() 
NAND2_X1_1769_ (
  .A1({ S14842 }),
  .A2({ S41 }),
  .ZN({ S14848 })
);
NOR2_X1 #() 
NOR2_X1_414_ (
  .A1({ S14847 }),
  .A2({ S14848 }),
  .ZN({ S14849 })
);
NAND3_X1 #() 
NAND3_X1_2067_ (
  .A1({ S13074 }),
  .A2({ S13078 }),
  .A3({ S11984 }),
  .ZN({ S14850 })
);
NAND3_X1 #() 
NAND3_X1_2068_ (
  .A1({ S13080 }),
  .A2({ S13081 }),
  .A3({ S25957[412] }),
  .ZN({ S14851 })
);
NAND2_X1 #() 
NAND2_X1_1770_ (
  .A1({ S14850 }),
  .A2({ S14851 }),
  .ZN({ S14852 })
);
OAI21_X1 #() 
OAI21_X1_973_ (
  .A({ S14834 }),
  .B1({ S14829 }),
  .B2({ S14828 }),
  .ZN({ S14853 })
);
OAI21_X1 #() 
OAI21_X1_974_ (
  .A({ S14834 }),
  .B1({ S14826 }),
  .B2({ S14825 }),
  .ZN({ S14854 })
);
NAND2_X1 #() 
NAND2_X1_1771_ (
  .A1({ S14854 }),
  .A2({ S14841 }),
  .ZN({ S14855 })
);
NAND3_X1 #() 
NAND3_X1_2069_ (
  .A1({ S14855 }),
  .A2({ S25957[283] }),
  .A3({ S14853 }),
  .ZN({ S14856 })
);
NAND2_X1 #() 
NAND2_X1_1772_ (
  .A1({ S14856 }),
  .A2({ S14852 }),
  .ZN({ S14858 })
);
OAI22_X1 #() 
OAI22_X1_45_ (
  .A1({ S14840 }),
  .A2({ S14844 }),
  .B1({ S14858 }),
  .B2({ S14849 }),
  .ZN({ S14859 })
);
NAND2_X1 #() 
NAND2_X1_1773_ (
  .A1({ S14845 }),
  .A2({ S14842 }),
  .ZN({ S14860 })
);
INV_X1 #() 
INV_X1_570_ (
  .A({ S14860 }),
  .ZN({ S14861 })
);
OAI211_X1 #() 
OAI211_X1_651_ (
  .A({ S13318 }),
  .B({ S13321 }),
  .C1({ S14826 }),
  .C2({ S14825 }),
  .ZN({ S14862 })
);
NAND2_X1 #() 
NAND2_X1_1774_ (
  .A1({ S14854 }),
  .A2({ S14836 }),
  .ZN({ S14863 })
);
NAND2_X1 #() 
NAND2_X1_1775_ (
  .A1({ S14863 }),
  .A2({ S14862 }),
  .ZN({ S14864 })
);
AOI21_X1 #() 
AOI21_X1_1061_ (
  .A({ S41 }),
  .B1({ S14864 }),
  .B2({ S14861 }),
  .ZN({ S14865 })
);
OAI211_X1 #() 
OAI211_X1_652_ (
  .A({ S13209 }),
  .B({ S13239 }),
  .C1({ S14829 }),
  .C2({ S14828 }),
  .ZN({ S14866 })
);
NAND3_X1 #() 
NAND3_X1_2070_ (
  .A1({ S14866 }),
  .A2({ S14862 }),
  .A3({ S25957[282] }),
  .ZN({ S14867 })
);
AOI21_X1 #() 
AOI21_X1_1062_ (
  .A({ S25957[283] }),
  .B1({ S14867 }),
  .B2({ S14837 }),
  .ZN({ S14869 })
);
OR3_X1 #() 
OR3_X1_7_ (
  .A1({ S14865 }),
  .A2({ S14869 }),
  .A3({ S14852 }),
  .ZN({ S14870 })
);
AOI21_X1 #() 
AOI21_X1_1063_ (
  .A({ S41 }),
  .B1({ S25957[280] }),
  .B2({ S25957[282] }),
  .ZN({ S14871 })
);
NAND2_X1 #() 
NAND2_X1_1776_ (
  .A1({ S14871 }),
  .A2({ S14853 }),
  .ZN({ S14872 })
);
NAND4_X1 #() 
NAND4_X1_258_ (
  .A1({ S14853 }),
  .A2({ S14845 }),
  .A3({ S14842 }),
  .A4({ S14837 }),
  .ZN({ S14873 })
);
AOI21_X1 #() 
AOI21_X1_1064_ (
  .A({ S25957[284] }),
  .B1({ S14873 }),
  .B2({ S41 }),
  .ZN({ S14874 })
);
AOI21_X1 #() 
AOI21_X1_1065_ (
  .A({ S25957[285] }),
  .B1({ S14874 }),
  .B2({ S14872 }),
  .ZN({ S14875 })
);
AOI22_X1 #() 
AOI22_X1_241_ (
  .A1({ S14870 }),
  .A2({ S14875 }),
  .B1({ S14859 }),
  .B2({ S25957[285] }),
  .ZN({ S14876 })
);
NOR2_X1 #() 
NOR2_X1_415_ (
  .A1({ S14861 }),
  .A2({ S41 }),
  .ZN({ S14877 })
);
AOI22_X1 #() 
AOI22_X1_242_ (
  .A1({ S14845 }),
  .A2({ S14827 }),
  .B1({ S14841 }),
  .B2({ S25957[280] }),
  .ZN({ S14878 })
);
NAND2_X1 #() 
NAND2_X1_1777_ (
  .A1({ S14878 }),
  .A2({ S41 }),
  .ZN({ S14880 })
);
NAND2_X1 #() 
NAND2_X1_1778_ (
  .A1({ S14880 }),
  .A2({ S14852 }),
  .ZN({ S14881 })
);
NAND2_X1 #() 
NAND2_X1_1779_ (
  .A1({ S48 }),
  .A2({ S14834 }),
  .ZN({ S14882 })
);
INV_X1 #() 
INV_X1_571_ (
  .A({ S14882 }),
  .ZN({ S14883 })
);
NAND2_X1 #() 
NAND2_X1_1780_ (
  .A1({ S49 }),
  .A2({ S25957[282] }),
  .ZN({ S14884 })
);
OAI21_X1 #() 
OAI21_X1_975_ (
  .A({ S41 }),
  .B1({ S14884 }),
  .B2({ S48 }),
  .ZN({ S14885 })
);
NOR2_X1 #() 
NOR2_X1_416_ (
  .A1({ S14885 }),
  .A2({ S14883 }),
  .ZN({ S14886 })
);
NOR2_X1 #() 
NOR2_X1_417_ (
  .A1({ S14841 }),
  .A2({ S14842 }),
  .ZN({ S14887 })
);
OAI21_X1 #() 
OAI21_X1_976_ (
  .A({ S25957[284] }),
  .B1({ S14887 }),
  .B2({ S41 }),
  .ZN({ S14888 })
);
OAI22_X1 #() 
OAI22_X1_46_ (
  .A1({ S14881 }),
  .A2({ S14877 }),
  .B1({ S14886 }),
  .B2({ S14888 }),
  .ZN({ S14889 })
);
NAND2_X1 #() 
NAND2_X1_1781_ (
  .A1({ S25957[280] }),
  .A2({ S41 }),
  .ZN({ S14891 })
);
NAND2_X1 #() 
NAND2_X1_1782_ (
  .A1({ S14871 }),
  .A2({ S14836 }),
  .ZN({ S14892 })
);
NAND3_X1 #() 
NAND3_X1_2071_ (
  .A1({ S14892 }),
  .A2({ S25957[284] }),
  .A3({ S14891 }),
  .ZN({ S14893 })
);
INV_X1 #() 
INV_X1_572_ (
  .A({ S14838 }),
  .ZN({ S14894 })
);
AOI21_X1 #() 
AOI21_X1_1066_ (
  .A({ S14834 }),
  .B1({ S13318 }),
  .B2({ S13321 }),
  .ZN({ S14895 })
);
NOR2_X1 #() 
NOR2_X1_418_ (
  .A1({ S14895 }),
  .A2({ S25957[283] }),
  .ZN({ S14896 })
);
AOI21_X1 #() 
AOI21_X1_1067_ (
  .A({ S25957[282] }),
  .B1({ S13321 }),
  .B2({ S13318 }),
  .ZN({ S14897 })
);
NOR2_X1 #() 
NOR2_X1_419_ (
  .A1({ S14897 }),
  .A2({ S41 }),
  .ZN({ S14898 })
);
AOI22_X1 #() 
AOI22_X1_243_ (
  .A1({ S14898 }),
  .A2({ S14862 }),
  .B1({ S14894 }),
  .B2({ S14896 }),
  .ZN({ S14899 })
);
OAI211_X1 #() 
OAI211_X1_653_ (
  .A({ S25957[285] }),
  .B({ S14893 }),
  .C1({ S14899 }),
  .C2({ S25957[284] }),
  .ZN({ S14900 })
);
OAI211_X1 #() 
OAI211_X1_654_ (
  .A({ S14823 }),
  .B({ S14900 }),
  .C1({ S14889 }),
  .C2({ S25957[285] }),
  .ZN({ S14902 })
);
OAI211_X1 #() 
OAI211_X1_655_ (
  .A({ S14902 }),
  .B({ S14822 }),
  .C1({ S14876 }),
  .C2({ S14823 }),
  .ZN({ S14903 })
);
INV_X1 #() 
INV_X1_573_ (
  .A({ S14842 }),
  .ZN({ S14904 })
);
NAND2_X1 #() 
NAND2_X1_1783_ (
  .A1({ S14904 }),
  .A2({ S25957[281] }),
  .ZN({ S14905 })
);
AOI21_X1 #() 
AOI21_X1_1068_ (
  .A({ S41 }),
  .B1({ S14905 }),
  .B2({ S14862 }),
  .ZN({ S14906 })
);
AOI211_X1 #() 
AOI211_X1_24_ (
  .A({ S25957[284] }),
  .B({ S14906 }),
  .C1({ S41 }),
  .C2({ S14839 }),
  .ZN({ S14907 })
);
NAND2_X1 #() 
NAND2_X1_1784_ (
  .A1({ S14862 }),
  .A2({ S14834 }),
  .ZN({ S14908 })
);
OAI21_X1 #() 
OAI21_X1_977_ (
  .A({ S25957[284] }),
  .B1({ S14908 }),
  .B2({ S41 }),
  .ZN({ S14909 })
);
AOI21_X1 #() 
AOI21_X1_1069_ (
  .A({ S25957[283] }),
  .B1({ S13318 }),
  .B2({ S13321 }),
  .ZN({ S14910 })
);
INV_X1 #() 
INV_X1_574_ (
  .A({ S25957[280] }),
  .ZN({ S14911 })
);
NAND2_X1 #() 
NAND2_X1_1785_ (
  .A1({ S25957[282] }),
  .A2({ S25957[283] }),
  .ZN({ S14913 })
);
NOR2_X1 #() 
NOR2_X1_420_ (
  .A1({ S14911 }),
  .A2({ S14913 }),
  .ZN({ S14914 })
);
AOI211_X1 #() 
AOI211_X1_25_ (
  .A({ S14914 }),
  .B({ S14909 }),
  .C1({ S14910 }),
  .C2({ S14837 }),
  .ZN({ S14915 })
);
OAI21_X1 #() 
OAI21_X1_978_ (
  .A({ S25957[285] }),
  .B1({ S14907 }),
  .B2({ S14915 }),
  .ZN({ S14916 })
);
NAND2_X1 #() 
NAND2_X1_1786_ (
  .A1({ S25957[317] }),
  .A2({ S25957[413] }),
  .ZN({ S14917 })
);
NAND3_X1 #() 
NAND3_X1_2072_ (
  .A1({ S12964 }),
  .A2({ S12967 }),
  .A3({ S12034 }),
  .ZN({ S14918 })
);
NAND2_X1 #() 
NAND2_X1_1787_ (
  .A1({ S14917 }),
  .A2({ S14918 }),
  .ZN({ S14919 })
);
INV_X1 #() 
INV_X1_575_ (
  .A({ S14866 }),
  .ZN({ S14920 })
);
NOR2_X1 #() 
NOR2_X1_421_ (
  .A1({ S14920 }),
  .A2({ S25957[283] }),
  .ZN({ S14921 })
);
AOI21_X1 #() 
AOI21_X1_1070_ (
  .A({ S41 }),
  .B1({ S14866 }),
  .B2({ S14836 }),
  .ZN({ S14922 })
);
OAI21_X1 #() 
OAI21_X1_979_ (
  .A({ S25957[284] }),
  .B1({ S14921 }),
  .B2({ S14922 }),
  .ZN({ S14924 })
);
OAI211_X1 #() 
OAI211_X1_656_ (
  .A({ S14853 }),
  .B({ S14854 }),
  .C1({ S14845 }),
  .C2({ S25957[280] }),
  .ZN({ S14925 })
);
NOR2_X1 #() 
NOR2_X1_422_ (
  .A1({ S25957[281] }),
  .A2({ S41 }),
  .ZN({ S14926 })
);
AOI21_X1 #() 
AOI21_X1_1071_ (
  .A({ S25957[284] }),
  .B1({ S25957[280] }),
  .B2({ S14926 }),
  .ZN({ S14927 })
);
NAND2_X1 #() 
NAND2_X1_1788_ (
  .A1({ S14927 }),
  .A2({ S14925 }),
  .ZN({ S14928 })
);
NAND3_X1 #() 
NAND3_X1_2073_ (
  .A1({ S14924 }),
  .A2({ S14919 }),
  .A3({ S14928 }),
  .ZN({ S14929 })
);
NAND3_X1 #() 
NAND3_X1_2074_ (
  .A1({ S14916 }),
  .A2({ S25957[286] }),
  .A3({ S14929 }),
  .ZN({ S14930 })
);
AOI21_X1 #() 
AOI21_X1_1072_ (
  .A({ S41 }),
  .B1({ S14838 }),
  .B2({ S49 }),
  .ZN({ S14931 })
);
AOI21_X1 #() 
AOI21_X1_1073_ (
  .A({ S25957[283] }),
  .B1({ S25957[280] }),
  .B2({ S14834 }),
  .ZN({ S14932 })
);
AOI22_X1 #() 
AOI22_X1_244_ (
  .A1({ S14931 }),
  .A2({ S14867 }),
  .B1({ S14830 }),
  .B2({ S14932 }),
  .ZN({ S14933 })
);
OAI22_X1 #() 
OAI22_X1_47_ (
  .A1({ S14829 }),
  .A2({ S14828 }),
  .B1({ S14826 }),
  .B2({ S14825 }),
  .ZN({ S14935 })
);
NAND3_X1 #() 
NAND3_X1_2075_ (
  .A1({ S14935 }),
  .A2({ S14834 }),
  .A3({ S49 }),
  .ZN({ S14936 })
);
INV_X1 #() 
INV_X1_576_ (
  .A({ S14848 }),
  .ZN({ S14937 })
);
NAND3_X1 #() 
NAND3_X1_2076_ (
  .A1({ S14936 }),
  .A2({ S14937 }),
  .A3({ S14830 }),
  .ZN({ S14938 })
);
AND3_X1 #() 
AND3_X1_82_ (
  .A1({ S13318 }),
  .A2({ S13321 }),
  .A3({ S14834 }),
  .ZN({ S14939 })
);
NAND2_X1 #() 
NAND2_X1_1789_ (
  .A1({ S14939 }),
  .A2({ S25957[283] }),
  .ZN({ S14940 })
);
NAND3_X1 #() 
NAND3_X1_2077_ (
  .A1({ S14938 }),
  .A2({ S14852 }),
  .A3({ S14940 }),
  .ZN({ S14941 })
);
OAI21_X1 #() 
OAI21_X1_980_ (
  .A({ S14941 }),
  .B1({ S14933 }),
  .B2({ S14852 }),
  .ZN({ S14942 })
);
AOI21_X1 #() 
AOI21_X1_1074_ (
  .A({ S14834 }),
  .B1({ S13239 }),
  .B2({ S13209 }),
  .ZN({ S14943 })
);
NAND2_X1 #() 
NAND2_X1_1790_ (
  .A1({ S25957[281] }),
  .A2({ S41 }),
  .ZN({ S14944 })
);
NOR2_X1 #() 
NOR2_X1_423_ (
  .A1({ S14914 }),
  .A2({ S14926 }),
  .ZN({ S14946 })
);
OAI21_X1 #() 
OAI21_X1_981_ (
  .A({ S14946 }),
  .B1({ S14943 }),
  .B2({ S14944 }),
  .ZN({ S14947 })
);
OAI21_X1 #() 
OAI21_X1_982_ (
  .A({ S41 }),
  .B1({ S14837 }),
  .B2({ S25957[281] }),
  .ZN({ S14948 })
);
AOI21_X1 #() 
AOI21_X1_1075_ (
  .A({ S25957[284] }),
  .B1({ S14948 }),
  .B2({ S14935 }),
  .ZN({ S14949 })
);
AOI21_X1 #() 
AOI21_X1_1076_ (
  .A({ S14949 }),
  .B1({ S14947 }),
  .B2({ S25957[284] }),
  .ZN({ S14950 })
);
AOI21_X1 #() 
AOI21_X1_1077_ (
  .A({ S25957[286] }),
  .B1({ S14950 }),
  .B2({ S25957[285] }),
  .ZN({ S14951 })
);
OAI21_X1 #() 
OAI21_X1_983_ (
  .A({ S14951 }),
  .B1({ S25957[285] }),
  .B2({ S14942 }),
  .ZN({ S14952 })
);
NAND3_X1 #() 
NAND3_X1_2078_ (
  .A1({ S14930 }),
  .A2({ S25957[287] }),
  .A3({ S14952 }),
  .ZN({ S14953 })
);
NAND3_X1 #() 
NAND3_X1_2079_ (
  .A1({ S14953 }),
  .A2({ S12112 }),
  .A3({ S14903 }),
  .ZN({ S14954 })
);
INV_X1 #() 
INV_X1_577_ (
  .A({ S14954 }),
  .ZN({ S14955 })
);
AOI21_X1 #() 
AOI21_X1_1078_ (
  .A({ S12112 }),
  .B1({ S14953 }),
  .B2({ S14903 }),
  .ZN({ S14957 })
);
NOR2_X1 #() 
NOR2_X1_424_ (
  .A1({ S14955 }),
  .A2({ S14957 }),
  .ZN({ S25957[199] })
);
AND2_X1 #() 
AND2_X1_107_ (
  .A1({ S25957[199] }),
  .A2({ S25957[295] }),
  .ZN({ S14958 })
);
NOR2_X1 #() 
NOR2_X1_425_ (
  .A1({ S25957[199] }),
  .A2({ S25957[295] }),
  .ZN({ S14959 })
);
NOR2_X1 #() 
NOR2_X1_426_ (
  .A1({ S14958 }),
  .A2({ S14959 }),
  .ZN({ S25957[167] })
);
INV_X1 #() 
INV_X1_578_ (
  .A({ S25957[167] }),
  .ZN({ S14960 })
);
NAND2_X1 #() 
NAND2_X1_1791_ (
  .A1({ S14960 }),
  .A2({ S12121 }),
  .ZN({ S14961 })
);
NAND2_X1 #() 
NAND2_X1_1792_ (
  .A1({ S25957[167] }),
  .A2({ S25957[263] }),
  .ZN({ S14962 })
);
AND2_X1 #() 
AND2_X1_108_ (
  .A1({ S14961 }),
  .A2({ S14962 }),
  .ZN({ S25957[135] })
);
NAND2_X1 #() 
NAND2_X1_1793_ (
  .A1({ S14866 }),
  .A2({ S14830 }),
  .ZN({ S14963 })
);
OAI21_X1 #() 
OAI21_X1_984_ (
  .A({ S14852 }),
  .B1({ S14963 }),
  .B2({ S14914 }),
  .ZN({ S14965 })
);
INV_X1 #() 
INV_X1_579_ (
  .A({ S14965 }),
  .ZN({ S14966 })
);
NAND3_X1 #() 
NAND3_X1_2080_ (
  .A1({ S14932 }),
  .A2({ S14845 }),
  .A3({ S14842 }),
  .ZN({ S14967 })
);
NAND2_X1 #() 
NAND2_X1_1794_ (
  .A1({ S49 }),
  .A2({ S14854 }),
  .ZN({ S14968 })
);
INV_X1 #() 
INV_X1_580_ (
  .A({ S14968 }),
  .ZN({ S14969 })
);
AOI21_X1 #() 
AOI21_X1_1079_ (
  .A({ S14852 }),
  .B1({ S14969 }),
  .B2({ S25957[283] }),
  .ZN({ S14970 })
);
AOI21_X1 #() 
AOI21_X1_1080_ (
  .A({ S14966 }),
  .B1({ S14967 }),
  .B2({ S14970 }),
  .ZN({ S14971 })
);
NAND3_X1 #() 
NAND3_X1_2081_ (
  .A1({ S14830 }),
  .A2({ S14854 }),
  .A3({ S14842 }),
  .ZN({ S14972 })
);
NAND2_X1 #() 
NAND2_X1_1795_ (
  .A1({ S14972 }),
  .A2({ S25957[283] }),
  .ZN({ S14973 })
);
AND2_X1 #() 
AND2_X1_109_ (
  .A1({ S14885 }),
  .A2({ S14973 }),
  .ZN({ S14974 })
);
NAND2_X1 #() 
NAND2_X1_1796_ (
  .A1({ S14911 }),
  .A2({ S14836 }),
  .ZN({ S14976 })
);
AOI21_X1 #() 
AOI21_X1_1081_ (
  .A({ S14852 }),
  .B1({ S14976 }),
  .B2({ S41 }),
  .ZN({ S14977 })
);
INV_X1 #() 
INV_X1_581_ (
  .A({ S14977 }),
  .ZN({ S14978 })
);
OAI22_X1 #() 
OAI22_X1_48_ (
  .A1({ S14974 }),
  .A2({ S25957[284] }),
  .B1({ S14898 }),
  .B2({ S14978 }),
  .ZN({ S14979 })
);
NAND2_X1 #() 
NAND2_X1_1797_ (
  .A1({ S14979 }),
  .A2({ S14919 }),
  .ZN({ S14980 })
);
OAI21_X1 #() 
OAI21_X1_985_ (
  .A({ S14980 }),
  .B1({ S14919 }),
  .B2({ S14971 }),
  .ZN({ S14981 })
);
NAND2_X1 #() 
NAND2_X1_1798_ (
  .A1({ S14853 }),
  .A2({ S25957[283] }),
  .ZN({ S14982 })
);
NAND2_X1 #() 
NAND2_X1_1799_ (
  .A1({ S14939 }),
  .A2({ S25957[280] }),
  .ZN({ S14983 })
);
NAND2_X1 #() 
NAND2_X1_1800_ (
  .A1({ S14983 }),
  .A2({ S14896 }),
  .ZN({ S14984 })
);
OAI21_X1 #() 
OAI21_X1_986_ (
  .A({ S14984 }),
  .B1({ S14847 }),
  .B2({ S14982 }),
  .ZN({ S14985 })
);
NAND2_X1 #() 
NAND2_X1_1801_ (
  .A1({ S14904 }),
  .A2({ S14841 }),
  .ZN({ S14987 })
);
NAND2_X1 #() 
NAND2_X1_1802_ (
  .A1({ S14987 }),
  .A2({ S14935 }),
  .ZN({ S14988 })
);
NOR2_X1 #() 
NOR2_X1_427_ (
  .A1({ S14988 }),
  .A2({ S41 }),
  .ZN({ S14989 })
);
NAND2_X1 #() 
NAND2_X1_1803_ (
  .A1({ S14854 }),
  .A2({ S41 }),
  .ZN({ S14990 })
);
NAND2_X1 #() 
NAND2_X1_1804_ (
  .A1({ S14990 }),
  .A2({ S25957[284] }),
  .ZN({ S14991 })
);
OAI221_X1 #() 
OAI221_X1_39_ (
  .A({ S25957[285] }),
  .B1({ S14989 }),
  .B2({ S14991 }),
  .C1({ S25957[284] }),
  .C2({ S14985 }),
  .ZN({ S14992 })
);
OAI211_X1 #() 
OAI211_X1_657_ (
  .A({ S14836 }),
  .B({ S14854 }),
  .C1({ S14841 }),
  .C2({ S14842 }),
  .ZN({ S14993 })
);
NAND2_X1 #() 
NAND2_X1_1805_ (
  .A1({ S14993 }),
  .A2({ S25957[283] }),
  .ZN({ S14994 })
);
INV_X1 #() 
INV_X1_582_ (
  .A({ S14994 }),
  .ZN({ S14995 })
);
NAND2_X1 #() 
NAND2_X1_1806_ (
  .A1({ S14990 }),
  .A2({ S14944 }),
  .ZN({ S14996 })
);
NOR2_X1 #() 
NOR2_X1_428_ (
  .A1({ S14996 }),
  .A2({ S14852 }),
  .ZN({ S14998 })
);
AOI22_X1 #() 
AOI22_X1_245_ (
  .A1({ S14995 }),
  .A2({ S14852 }),
  .B1({ S14998 }),
  .B2({ S14856 }),
  .ZN({ S14999 })
);
OAI211_X1 #() 
OAI211_X1_658_ (
  .A({ S14992 }),
  .B({ S14823 }),
  .C1({ S25957[285] }),
  .C2({ S14999 }),
  .ZN({ S15000 })
);
OAI211_X1 #() 
OAI211_X1_659_ (
  .A({ S15000 }),
  .B({ S14822 }),
  .C1({ S14981 }),
  .C2({ S14823 }),
  .ZN({ S15001 })
);
INV_X1 #() 
INV_X1_583_ (
  .A({ S14874 }),
  .ZN({ S15002 })
);
NAND2_X1 #() 
NAND2_X1_1807_ (
  .A1({ S14864 }),
  .A2({ S14937 }),
  .ZN({ S15003 })
);
NAND3_X1 #() 
NAND3_X1_2082_ (
  .A1({ S15003 }),
  .A2({ S25957[284] }),
  .A3({ S14973 }),
  .ZN({ S15004 })
);
NAND2_X1 #() 
NAND2_X1_1808_ (
  .A1({ S14837 }),
  .A2({ S25957[281] }),
  .ZN({ S15005 })
);
AOI21_X1 #() 
AOI21_X1_1082_ (
  .A({ S41 }),
  .B1({ S15005 }),
  .B2({ S14827 }),
  .ZN({ S15006 })
);
OAI211_X1 #() 
OAI211_X1_660_ (
  .A({ S15004 }),
  .B({ S14919 }),
  .C1({ S15002 }),
  .C2({ S15006 }),
  .ZN({ S15007 })
);
NOR2_X1 #() 
NOR2_X1_429_ (
  .A1({ S14884 }),
  .A2({ S25957[283] }),
  .ZN({ S15009 })
);
OAI21_X1 #() 
OAI21_X1_987_ (
  .A({ S14852 }),
  .B1({ S14922 }),
  .B2({ S14910 }),
  .ZN({ S15010 })
);
NAND2_X1 #() 
NAND2_X1_1809_ (
  .A1({ S14842 }),
  .A2({ S25957[283] }),
  .ZN({ S15011 })
);
OAI21_X1 #() 
OAI21_X1_988_ (
  .A({ S25957[284] }),
  .B1({ S14855 }),
  .B2({ S15011 }),
  .ZN({ S15012 })
);
OAI21_X1 #() 
OAI21_X1_989_ (
  .A({ S15010 }),
  .B1({ S15009 }),
  .B2({ S15012 }),
  .ZN({ S15013 })
);
NAND2_X1 #() 
NAND2_X1_1810_ (
  .A1({ S15013 }),
  .A2({ S25957[285] }),
  .ZN({ S15014 })
);
AOI21_X1 #() 
AOI21_X1_1083_ (
  .A({ S14823 }),
  .B1({ S15007 }),
  .B2({ S15014 }),
  .ZN({ S15015 })
);
AND3_X1 #() 
AND3_X1_83_ (
  .A1({ S14834 }),
  .A2({ S13209 }),
  .A3({ S13239 }),
  .ZN({ S15016 })
);
NAND3_X1 #() 
NAND3_X1_2083_ (
  .A1({ S14845 }),
  .A2({ S14827 }),
  .A3({ S25957[283] }),
  .ZN({ S15017 })
);
OAI21_X1 #() 
OAI21_X1_990_ (
  .A({ S15003 }),
  .B1({ S15016 }),
  .B2({ S15017 }),
  .ZN({ S15018 })
);
OAI21_X1 #() 
OAI21_X1_991_ (
  .A({ S14946 }),
  .B1({ S25957[283] }),
  .B2({ S14908 }),
  .ZN({ S15020 })
);
NAND2_X1 #() 
NAND2_X1_1811_ (
  .A1({ S15020 }),
  .A2({ S25957[284] }),
  .ZN({ S15021 })
);
OAI211_X1 #() 
OAI211_X1_661_ (
  .A({ S15021 }),
  .B({ S14919 }),
  .C1({ S15018 }),
  .C2({ S25957[284] }),
  .ZN({ S15022 })
);
NAND2_X1 #() 
NAND2_X1_1812_ (
  .A1({ S15016 }),
  .A2({ S14910 }),
  .ZN({ S15023 })
);
AOI21_X1 #() 
AOI21_X1_1084_ (
  .A({ S14852 }),
  .B1({ S25957[283] }),
  .B2({ S14895 }),
  .ZN({ S15024 })
);
NAND3_X1 #() 
NAND3_X1_2084_ (
  .A1({ S14880 }),
  .A2({ S15023 }),
  .A3({ S15024 }),
  .ZN({ S15025 })
);
NOR2_X1 #() 
NOR2_X1_430_ (
  .A1({ S14841 }),
  .A2({ S14837 }),
  .ZN({ S15026 })
);
NOR2_X1 #() 
NOR2_X1_431_ (
  .A1({ S15026 }),
  .A2({ S14847 }),
  .ZN({ S15027 })
);
NAND3_X1 #() 
NAND3_X1_2085_ (
  .A1({ S25957[281] }),
  .A2({ S25957[280] }),
  .A3({ S25957[282] }),
  .ZN({ S15028 })
);
NAND3_X1 #() 
NAND3_X1_2086_ (
  .A1({ S15028 }),
  .A2({ S41 }),
  .A3({ S49 }),
  .ZN({ S15029 })
);
OAI211_X1 #() 
OAI211_X1_662_ (
  .A({ S14852 }),
  .B({ S15029 }),
  .C1({ S15027 }),
  .C2({ S41 }),
  .ZN({ S15031 })
);
NAND3_X1 #() 
NAND3_X1_2087_ (
  .A1({ S15025 }),
  .A2({ S15031 }),
  .A3({ S25957[285] }),
  .ZN({ S15032 })
);
AOI21_X1 #() 
AOI21_X1_1085_ (
  .A({ S25957[286] }),
  .B1({ S15022 }),
  .B2({ S15032 }),
  .ZN({ S15033 })
);
OAI21_X1 #() 
OAI21_X1_992_ (
  .A({ S25957[287] }),
  .B1({ S15033 }),
  .B2({ S15015 }),
  .ZN({ S15034 })
);
AOI21_X1 #() 
AOI21_X1_1086_ (
  .A({ S25957[454] }),
  .B1({ S15001 }),
  .B2({ S15034 }),
  .ZN({ S15035 })
);
NAND2_X1 #() 
NAND2_X1_1813_ (
  .A1({ S15001 }),
  .A2({ S15034 }),
  .ZN({ S15036 })
);
NOR2_X1 #() 
NOR2_X1_432_ (
  .A1({ S15036 }),
  .A2({ S12195 }),
  .ZN({ S15037 })
);
OAI21_X1 #() 
OAI21_X1_993_ (
  .A({ S11418 }),
  .B1({ S15037 }),
  .B2({ S15035 }),
  .ZN({ S15038 })
);
NOR2_X1 #() 
NOR2_X1_433_ (
  .A1({ S15037 }),
  .A2({ S15035 }),
  .ZN({ S25957[198] })
);
NAND2_X1 #() 
NAND2_X1_1814_ (
  .A1({ S25957[198] }),
  .A2({ S25957[390] }),
  .ZN({ S15039 })
);
NAND2_X1 #() 
NAND2_X1_1815_ (
  .A1({ S15039 }),
  .A2({ S15038 }),
  .ZN({ S15041 })
);
INV_X1 #() 
INV_X1_584_ (
  .A({ S15041 }),
  .ZN({ S25957[134] })
);
XNOR2_X1 #() 
XNOR2_X1_61_ (
  .A({ S12200 }),
  .B({ S25957[549] }),
  .ZN({ S25957[421] })
);
INV_X1 #() 
INV_X1_585_ (
  .A({ S25957[421] }),
  .ZN({ S15042 })
);
NOR2_X1 #() 
NOR2_X1_434_ (
  .A1({ S25957[280] }),
  .A2({ S41 }),
  .ZN({ S15043 })
);
AOI21_X1 #() 
AOI21_X1_1087_ (
  .A({ S15043 }),
  .B1({ S14932 }),
  .B2({ S14866 }),
  .ZN({ S15044 })
);
OAI21_X1 #() 
OAI21_X1_994_ (
  .A({ S25957[283] }),
  .B1({ S14841 }),
  .B2({ S14837 }),
  .ZN({ S15045 })
);
NAND4_X1 #() 
NAND4_X1_259_ (
  .A1({ S14853 }),
  .A2({ S14845 }),
  .A3({ S14837 }),
  .A4({ S41 }),
  .ZN({ S15046 })
);
OAI211_X1 #() 
OAI211_X1_663_ (
  .A({ S25957[284] }),
  .B({ S15046 }),
  .C1({ S14878 }),
  .C2({ S15045 }),
  .ZN({ S15047 })
);
OAI21_X1 #() 
OAI21_X1_995_ (
  .A({ S15047 }),
  .B1({ S25957[284] }),
  .B2({ S15044 }),
  .ZN({ S15048 })
);
NAND2_X1 #() 
NAND2_X1_1816_ (
  .A1({ S15048 }),
  .A2({ S25957[285] }),
  .ZN({ S15050 })
);
AOI21_X1 #() 
AOI21_X1_1088_ (
  .A({ S25957[283] }),
  .B1({ S14861 }),
  .B2({ S14882 }),
  .ZN({ S15051 })
);
NOR2_X1 #() 
NOR2_X1_435_ (
  .A1({ S15051 }),
  .A2({ S14909 }),
  .ZN({ S15052 })
);
AOI21_X1 #() 
AOI21_X1_1089_ (
  .A({ S41 }),
  .B1({ S25957[280] }),
  .B2({ S14834 }),
  .ZN({ S15053 })
);
NAND3_X1 #() 
NAND3_X1_2088_ (
  .A1({ S15053 }),
  .A2({ S14845 }),
  .A3({ S14842 }),
  .ZN({ S15054 })
);
OAI21_X1 #() 
OAI21_X1_996_ (
  .A({ S41 }),
  .B1({ S14841 }),
  .B2({ S14837 }),
  .ZN({ S15055 })
);
AOI21_X1 #() 
AOI21_X1_1090_ (
  .A({ S25957[284] }),
  .B1({ S15054 }),
  .B2({ S15055 }),
  .ZN({ S15056 })
);
INV_X1 #() 
INV_X1_586_ (
  .A({ S15056 }),
  .ZN({ S15057 })
);
AOI21_X1 #() 
AOI21_X1_1091_ (
  .A({ S15057 }),
  .B1({ S15054 }),
  .B2({ S14943 }),
  .ZN({ S15058 })
);
OAI21_X1 #() 
OAI21_X1_997_ (
  .A({ S14919 }),
  .B1({ S15058 }),
  .B2({ S15052 }),
  .ZN({ S15059 })
);
NAND3_X1 #() 
NAND3_X1_2089_ (
  .A1({ S15059 }),
  .A2({ S25957[286] }),
  .A3({ S15050 }),
  .ZN({ S15061 })
);
OAI211_X1 #() 
OAI211_X1_664_ (
  .A({ S15023 }),
  .B({ S25957[284] }),
  .C1({ S41 }),
  .C2({ S14838 }),
  .ZN({ S15062 })
);
NOR2_X1 #() 
NOR2_X1_436_ (
  .A1({ S14937 }),
  .A2({ S14914 }),
  .ZN({ S15063 })
);
OAI21_X1 #() 
OAI21_X1_998_ (
  .A({ S15062 }),
  .B1({ S14965 }),
  .B2({ S15063 }),
  .ZN({ S15064 })
);
NAND2_X1 #() 
NAND2_X1_1817_ (
  .A1({ S15064 }),
  .A2({ S25957[285] }),
  .ZN({ S15065 })
);
OAI21_X1 #() 
OAI21_X1_999_ (
  .A({ S14927 }),
  .B1({ S25957[283] }),
  .B2({ S15028 }),
  .ZN({ S15066 })
);
NOR2_X1 #() 
NOR2_X1_437_ (
  .A1({ S14988 }),
  .A2({ S15053 }),
  .ZN({ S15067 })
);
NAND4_X1 #() 
NAND4_X1_260_ (
  .A1({ S14866 }),
  .A2({ S14862 }),
  .A3({ S25957[283] }),
  .A4({ S25957[282] }),
  .ZN({ S15068 })
);
NAND2_X1 #() 
NAND2_X1_1818_ (
  .A1({ S15068 }),
  .A2({ S25957[284] }),
  .ZN({ S15069 })
);
OAI211_X1 #() 
OAI211_X1_665_ (
  .A({ S15066 }),
  .B({ S14919 }),
  .C1({ S15067 }),
  .C2({ S15069 }),
  .ZN({ S15070 })
);
NAND3_X1 #() 
NAND3_X1_2090_ (
  .A1({ S15070 }),
  .A2({ S15065 }),
  .A3({ S14823 }),
  .ZN({ S15072 })
);
NAND3_X1 #() 
NAND3_X1_2091_ (
  .A1({ S15061 }),
  .A2({ S14822 }),
  .A3({ S15072 }),
  .ZN({ S15073 })
);
NAND2_X1 #() 
NAND2_X1_1819_ (
  .A1({ S14921 }),
  .A2({ S14908 }),
  .ZN({ S15074 })
);
OAI21_X1 #() 
OAI21_X1_1000_ (
  .A({ S15074 }),
  .B1({ S41 }),
  .B2({ S14976 }),
  .ZN({ S15075 })
);
NAND2_X1 #() 
NAND2_X1_1820_ (
  .A1({ S15075 }),
  .A2({ S25957[284] }),
  .ZN({ S15076 })
);
NAND2_X1 #() 
NAND2_X1_1821_ (
  .A1({ S15005 }),
  .A2({ S25957[283] }),
  .ZN({ S15077 })
);
NAND4_X1 #() 
NAND4_X1_261_ (
  .A1({ S15077 }),
  .A2({ S14944 }),
  .A3({ S14827 }),
  .A4({ S14852 }),
  .ZN({ S15078 })
);
NAND3_X1 #() 
NAND3_X1_2092_ (
  .A1({ S15076 }),
  .A2({ S25957[285] }),
  .A3({ S15078 }),
  .ZN({ S15079 })
);
AOI21_X1 #() 
AOI21_X1_1092_ (
  .A({ S14881 }),
  .B1({ S25957[283] }),
  .B2({ S14972 }),
  .ZN({ S15080 })
);
NAND2_X1 #() 
NAND2_X1_1822_ (
  .A1({ S14845 }),
  .A2({ S14827 }),
  .ZN({ S15081 })
);
NAND2_X1 #() 
NAND2_X1_1823_ (
  .A1({ S15081 }),
  .A2({ S41 }),
  .ZN({ S15083 })
);
NAND2_X1 #() 
NAND2_X1_1824_ (
  .A1({ S15053 }),
  .A2({ S14836 }),
  .ZN({ S15084 })
);
NAND2_X1 #() 
NAND2_X1_1825_ (
  .A1({ S15083 }),
  .A2({ S15084 }),
  .ZN({ S15085 })
);
INV_X1 #() 
INV_X1_587_ (
  .A({ S15085 }),
  .ZN({ S15086 })
);
AOI21_X1 #() 
AOI21_X1_1093_ (
  .A({ S15080 }),
  .B1({ S25957[284] }),
  .B2({ S15086 }),
  .ZN({ S15087 })
);
NAND2_X1 #() 
NAND2_X1_1826_ (
  .A1({ S15087 }),
  .A2({ S14919 }),
  .ZN({ S15088 })
);
NAND3_X1 #() 
NAND3_X1_2093_ (
  .A1({ S15088 }),
  .A2({ S25957[286] }),
  .A3({ S15079 }),
  .ZN({ S15089 })
);
NAND3_X1 #() 
NAND3_X1_2094_ (
  .A1({ S14866 }),
  .A2({ S41 }),
  .A3({ S14836 }),
  .ZN({ S15090 })
);
NOR2_X1 #() 
NOR2_X1_438_ (
  .A1({ S14926 }),
  .A2({ S25957[284] }),
  .ZN({ S15091 })
);
NOR2_X1 #() 
NOR2_X1_439_ (
  .A1({ S14891 }),
  .A2({ S14841 }),
  .ZN({ S15092 })
);
INV_X1 #() 
INV_X1_588_ (
  .A({ S15092 }),
  .ZN({ S15094 })
);
NAND2_X1 #() 
NAND2_X1_1827_ (
  .A1({ S14837 }),
  .A2({ S41 }),
  .ZN({ S15095 })
);
OAI21_X1 #() 
OAI21_X1_1001_ (
  .A({ S15095 }),
  .B1({ S14873 }),
  .B2({ S41 }),
  .ZN({ S15096 })
);
AOI21_X1 #() 
AOI21_X1_1094_ (
  .A({ S14852 }),
  .B1({ S15096 }),
  .B2({ S15094 }),
  .ZN({ S15097 })
);
AOI21_X1 #() 
AOI21_X1_1095_ (
  .A({ S15097 }),
  .B1({ S15091 }),
  .B2({ S15090 }),
  .ZN({ S15098 })
);
AOI21_X1 #() 
AOI21_X1_1096_ (
  .A({ S25957[282] }),
  .B1({ S14866 }),
  .B2({ S14862 }),
  .ZN({ S15099 })
);
NAND2_X1 #() 
NAND2_X1_1828_ (
  .A1({ S15099 }),
  .A2({ S25957[283] }),
  .ZN({ S15100 })
);
AOI21_X1 #() 
AOI21_X1_1097_ (
  .A({ S14852 }),
  .B1({ S14932 }),
  .B2({ S14841 }),
  .ZN({ S15101 })
);
NAND2_X1 #() 
NAND2_X1_1829_ (
  .A1({ S15100 }),
  .A2({ S15101 }),
  .ZN({ S15102 })
);
NOR2_X1 #() 
NOR2_X1_440_ (
  .A1({ S14884 }),
  .A2({ S48 }),
  .ZN({ S15103 })
);
OAI21_X1 #() 
OAI21_X1_1002_ (
  .A({ S25957[283] }),
  .B1({ S14837 }),
  .B2({ S25957[281] }),
  .ZN({ S15105 })
);
OAI221_X1 #() 
OAI221_X1_40_ (
  .A({ S14852 }),
  .B1({ S14853 }),
  .B2({ S14891 }),
  .C1({ S15103 }),
  .C2({ S15105 }),
  .ZN({ S15106 })
);
AOI21_X1 #() 
AOI21_X1_1098_ (
  .A({ S25957[285] }),
  .B1({ S15106 }),
  .B2({ S15102 }),
  .ZN({ S15107 })
);
AOI21_X1 #() 
AOI21_X1_1099_ (
  .A({ S15107 }),
  .B1({ S15098 }),
  .B2({ S25957[285] }),
  .ZN({ S15108 })
);
NAND2_X1 #() 
NAND2_X1_1830_ (
  .A1({ S15108 }),
  .A2({ S14823 }),
  .ZN({ S15109 })
);
NAND3_X1 #() 
NAND3_X1_2095_ (
  .A1({ S15089 }),
  .A2({ S15109 }),
  .A3({ S25957[287] }),
  .ZN({ S15110 })
);
NAND3_X1 #() 
NAND3_X1_2096_ (
  .A1({ S15110 }),
  .A2({ S25957[357] }),
  .A3({ S15073 }),
  .ZN({ S15111 })
);
INV_X1 #() 
INV_X1_589_ (
  .A({ S25957[357] }),
  .ZN({ S15112 })
);
NAND2_X1 #() 
NAND2_X1_1831_ (
  .A1({ S15076 }),
  .A2({ S15078 }),
  .ZN({ S15113 })
);
NAND2_X1 #() 
NAND2_X1_1832_ (
  .A1({ S15113 }),
  .A2({ S25957[285] }),
  .ZN({ S15114 })
);
OAI211_X1 #() 
OAI211_X1_666_ (
  .A({ S15114 }),
  .B({ S25957[286] }),
  .C1({ S15087 }),
  .C2({ S25957[285] }),
  .ZN({ S15116 })
);
OAI211_X1 #() 
OAI211_X1_667_ (
  .A({ S15116 }),
  .B({ S25957[287] }),
  .C1({ S25957[286] }),
  .C2({ S15108 }),
  .ZN({ S15117 })
);
NAND2_X1 #() 
NAND2_X1_1833_ (
  .A1({ S15061 }),
  .A2({ S15072 }),
  .ZN({ S15118 })
);
NAND2_X1 #() 
NAND2_X1_1834_ (
  .A1({ S15118 }),
  .A2({ S14822 }),
  .ZN({ S15119 })
);
NAND3_X1 #() 
NAND3_X1_2097_ (
  .A1({ S15117 }),
  .A2({ S15119 }),
  .A3({ S15112 }),
  .ZN({ S15120 })
);
NAND3_X1 #() 
NAND3_X1_2098_ (
  .A1({ S15120 }),
  .A2({ S15111 }),
  .A3({ S15042 }),
  .ZN({ S15121 })
);
NAND3_X1 #() 
NAND3_X1_2099_ (
  .A1({ S15110 }),
  .A2({ S15112 }),
  .A3({ S15073 }),
  .ZN({ S15122 })
);
NAND3_X1 #() 
NAND3_X1_2100_ (
  .A1({ S15117 }),
  .A2({ S15119 }),
  .A3({ S25957[357] }),
  .ZN({ S15123 })
);
NAND3_X1 #() 
NAND3_X1_2101_ (
  .A1({ S15123 }),
  .A2({ S15122 }),
  .A3({ S25957[421] }),
  .ZN({ S15124 })
);
NAND3_X1 #() 
NAND3_X1_2102_ (
  .A1({ S15121 }),
  .A2({ S15124 }),
  .A3({ S14186 }),
  .ZN({ S15125 })
);
NAND2_X1 #() 
NAND2_X1_1835_ (
  .A1({ S12273 }),
  .A2({ S12277 }),
  .ZN({ S25957[325] })
);
XNOR2_X1 #() 
XNOR2_X1_62_ (
  .A({ S25957[325] }),
  .B({ S15042 }),
  .ZN({ S25957[293] })
);
NAND3_X1 #() 
NAND3_X1_2103_ (
  .A1({ S15110 }),
  .A2({ S25957[453] }),
  .A3({ S15073 }),
  .ZN({ S15127 })
);
NAND3_X1 #() 
NAND3_X1_2104_ (
  .A1({ S15117 }),
  .A2({ S15119 }),
  .A3({ S12200 }),
  .ZN({ S15128 })
);
NAND3_X1 #() 
NAND3_X1_2105_ (
  .A1({ S15128 }),
  .A2({ S15127 }),
  .A3({ S25957[293] }),
  .ZN({ S15129 })
);
INV_X1 #() 
INV_X1_590_ (
  .A({ S25957[293] }),
  .ZN({ S15130 })
);
AOI21_X1 #() 
AOI21_X1_1100_ (
  .A({ S12200 }),
  .B1({ S15117 }),
  .B2({ S15119 }),
  .ZN({ S15131 })
);
AOI21_X1 #() 
AOI21_X1_1101_ (
  .A({ S25957[453] }),
  .B1({ S15110 }),
  .B2({ S15073 }),
  .ZN({ S15132 })
);
OAI21_X1 #() 
OAI21_X1_1003_ (
  .A({ S15130 }),
  .B1({ S15131 }),
  .B2({ S15132 }),
  .ZN({ S15133 })
);
NAND3_X1 #() 
NAND3_X1_2106_ (
  .A1({ S15133 }),
  .A2({ S15129 }),
  .A3({ S25957[261] }),
  .ZN({ S15134 })
);
AND2_X1 #() 
AND2_X1_110_ (
  .A1({ S15134 }),
  .A2({ S15125 }),
  .ZN({ S25957[133] })
);
NOR2_X1 #() 
NOR2_X1_441_ (
  .A1({ S12352 }),
  .A2({ S12355 }),
  .ZN({ S25957[292] })
);
XOR2_X1 #() 
XOR2_X1_28_ (
  .A({ S25957[356] }),
  .B({ S25957[452] }),
  .Z({ S25957[324] })
);
INV_X1 #() 
INV_X1_591_ (
  .A({ S25957[356] }),
  .ZN({ S15136 })
);
NAND3_X1 #() 
NAND3_X1_2107_ (
  .A1({ S14884 }),
  .A2({ S41 }),
  .A3({ S14836 }),
  .ZN({ S15137 })
);
NAND3_X1 #() 
NAND3_X1_2108_ (
  .A1({ S14946 }),
  .A2({ S15137 }),
  .A3({ S25957[284] }),
  .ZN({ S15138 })
);
NAND3_X1 #() 
NAND3_X1_2109_ (
  .A1({ S14827 }),
  .A2({ S14836 }),
  .A3({ S14837 }),
  .ZN({ S15139 })
);
NAND2_X1 #() 
NAND2_X1_1836_ (
  .A1({ S15139 }),
  .A2({ S41 }),
  .ZN({ S15140 })
);
NAND3_X1 #() 
NAND3_X1_2110_ (
  .A1({ S15140 }),
  .A2({ S14852 }),
  .A3({ S14913 }),
  .ZN({ S15141 })
);
NAND3_X1 #() 
NAND3_X1_2111_ (
  .A1({ S15138 }),
  .A2({ S15141 }),
  .A3({ S14919 }),
  .ZN({ S15142 })
);
INV_X1 #() 
INV_X1_592_ (
  .A({ S150 }),
  .ZN({ S15144 })
);
OAI21_X1 #() 
OAI21_X1_1004_ (
  .A({ S25957[284] }),
  .B1({ S15144 }),
  .B2({ S25957[282] }),
  .ZN({ S15145 })
);
NAND3_X1 #() 
NAND3_X1_2112_ (
  .A1({ S14838 }),
  .A2({ S41 }),
  .A3({ S49 }),
  .ZN({ S15146 })
);
NAND2_X1 #() 
NAND2_X1_1837_ (
  .A1({ S15083 }),
  .A2({ S15146 }),
  .ZN({ S15147 })
);
NAND2_X1 #() 
NAND2_X1_1838_ (
  .A1({ S15054 }),
  .A2({ S14852 }),
  .ZN({ S15148 })
);
OAI211_X1 #() 
OAI211_X1_668_ (
  .A({ S15145 }),
  .B({ S25957[285] }),
  .C1({ S15147 }),
  .C2({ S15148 }),
  .ZN({ S15149 })
);
AOI21_X1 #() 
AOI21_X1_1102_ (
  .A({ S14823 }),
  .B1({ S15142 }),
  .B2({ S15149 }),
  .ZN({ S15150 })
);
AOI21_X1 #() 
AOI21_X1_1103_ (
  .A({ S25957[284] }),
  .B1({ S15100 }),
  .B2({ S15094 }),
  .ZN({ S15151 })
);
NAND3_X1 #() 
NAND3_X1_2113_ (
  .A1({ S14856 }),
  .A2({ S15083 }),
  .A3({ S25957[284] }),
  .ZN({ S15152 })
);
INV_X1 #() 
INV_X1_593_ (
  .A({ S15152 }),
  .ZN({ S15153 })
);
OAI21_X1 #() 
OAI21_X1_1005_ (
  .A({ S25957[285] }),
  .B1({ S15151 }),
  .B2({ S15153 }),
  .ZN({ S15155 })
);
NAND2_X1 #() 
NAND2_X1_1839_ (
  .A1({ S14871 }),
  .A2({ S49 }),
  .ZN({ S15156 })
);
NAND2_X1 #() 
NAND2_X1_1840_ (
  .A1({ S49 }),
  .A2({ S14834 }),
  .ZN({ S15157 })
);
NAND3_X1 #() 
NAND3_X1_2114_ (
  .A1({ S14987 }),
  .A2({ S15157 }),
  .A3({ S41 }),
  .ZN({ S15158 })
);
AOI21_X1 #() 
AOI21_X1_1104_ (
  .A({ S25957[284] }),
  .B1({ S15158 }),
  .B2({ S15156 }),
  .ZN({ S15159 })
);
NAND2_X1 #() 
NAND2_X1_1841_ (
  .A1({ S14908 }),
  .A2({ S14871 }),
  .ZN({ S15160 })
);
NAND3_X1 #() 
NAND3_X1_2115_ (
  .A1({ S15160 }),
  .A2({ S25957[284] }),
  .A3({ S15090 }),
  .ZN({ S15161 })
);
INV_X1 #() 
INV_X1_594_ (
  .A({ S15161 }),
  .ZN({ S15162 })
);
OAI21_X1 #() 
OAI21_X1_1006_ (
  .A({ S14919 }),
  .B1({ S15162 }),
  .B2({ S15159 }),
  .ZN({ S15163 })
);
AOI21_X1 #() 
AOI21_X1_1105_ (
  .A({ S25957[286] }),
  .B1({ S15155 }),
  .B2({ S15163 }),
  .ZN({ S15164 })
);
OAI21_X1 #() 
OAI21_X1_1007_ (
  .A({ S14822 }),
  .B1({ S15164 }),
  .B2({ S15150 }),
  .ZN({ S15166 })
);
OAI211_X1 #() 
OAI211_X1_669_ (
  .A({ S15090 }),
  .B({ S25957[284] }),
  .C1({ S41 }),
  .C2({ S14855 }),
  .ZN({ S15167 })
);
INV_X1 #() 
INV_X1_595_ (
  .A({ S14862 }),
  .ZN({ S15168 })
);
NAND2_X1 #() 
NAND2_X1_1842_ (
  .A1({ S14937 }),
  .A2({ S14836 }),
  .ZN({ S15169 })
);
OAI211_X1 #() 
OAI211_X1_670_ (
  .A({ S15169 }),
  .B({ S14852 }),
  .C1({ S15168 }),
  .C2({ S14982 }),
  .ZN({ S15170 })
);
NAND3_X1 #() 
NAND3_X1_2116_ (
  .A1({ S15170 }),
  .A2({ S14919 }),
  .A3({ S15167 }),
  .ZN({ S15171 })
);
NAND2_X1 #() 
NAND2_X1_1843_ (
  .A1({ S14848 }),
  .A2({ S14944 }),
  .ZN({ S15172 })
);
NAND3_X1 #() 
NAND3_X1_2117_ (
  .A1({ S14853 }),
  .A2({ S14911 }),
  .A3({ S41 }),
  .ZN({ S15173 })
);
NAND3_X1 #() 
NAND3_X1_2118_ (
  .A1({ S14892 }),
  .A2({ S14852 }),
  .A3({ S15173 }),
  .ZN({ S15174 })
);
OAI211_X1 #() 
OAI211_X1_671_ (
  .A({ S15174 }),
  .B({ S25957[285] }),
  .C1({ S14909 }),
  .C2({ S15172 }),
  .ZN({ S15175 })
);
NAND3_X1 #() 
NAND3_X1_2119_ (
  .A1({ S15171 }),
  .A2({ S25957[286] }),
  .A3({ S15175 }),
  .ZN({ S15177 })
);
AOI22_X1 #() 
AOI22_X1_246_ (
  .A1({ S14836 }),
  .A2({ S14854 }),
  .B1({ S14841 }),
  .B2({ S25957[280] }),
  .ZN({ S15178 })
);
OAI21_X1 #() 
OAI21_X1_1008_ (
  .A({ S41 }),
  .B1({ S15178 }),
  .B2({ S14860 }),
  .ZN({ S15179 })
);
NAND4_X1 #() 
NAND4_X1_262_ (
  .A1({ S14862 }),
  .A2({ S14845 }),
  .A3({ S14827 }),
  .A4({ S25957[283] }),
  .ZN({ S15180 })
);
NAND3_X1 #() 
NAND3_X1_2120_ (
  .A1({ S15179 }),
  .A2({ S14852 }),
  .A3({ S15180 }),
  .ZN({ S15181 })
);
AOI21_X1 #() 
AOI21_X1_1106_ (
  .A({ S14852 }),
  .B1({ S14972 }),
  .B2({ S41 }),
  .ZN({ S15182 })
);
NAND2_X1 #() 
NAND2_X1_1844_ (
  .A1({ S14939 }),
  .A2({ S41 }),
  .ZN({ S15183 })
);
OAI211_X1 #() 
OAI211_X1_672_ (
  .A({ S15182 }),
  .B({ S15183 }),
  .C1({ S15045 }),
  .C2({ S15168 }),
  .ZN({ S15184 })
);
NAND3_X1 #() 
NAND3_X1_2121_ (
  .A1({ S15181 }),
  .A2({ S15184 }),
  .A3({ S25957[285] }),
  .ZN({ S15185 })
);
OAI21_X1 #() 
OAI21_X1_1009_ (
  .A({ S41 }),
  .B1({ S15005 }),
  .B2({ S14943 }),
  .ZN({ S15186 })
);
OAI21_X1 #() 
OAI21_X1_1010_ (
  .A({ S25957[283] }),
  .B1({ S14887 }),
  .B2({ S14939 }),
  .ZN({ S15188 })
);
NAND3_X1 #() 
NAND3_X1_2122_ (
  .A1({ S15188 }),
  .A2({ S25957[284] }),
  .A3({ S15186 }),
  .ZN({ S15189 })
);
NAND2_X1 #() 
NAND2_X1_1845_ (
  .A1({ S14993 }),
  .A2({ S41 }),
  .ZN({ S15190 })
);
NAND2_X1 #() 
NAND2_X1_1846_ (
  .A1({ S14871 }),
  .A2({ S14841 }),
  .ZN({ S15191 })
);
NAND3_X1 #() 
NAND3_X1_2123_ (
  .A1({ S15190 }),
  .A2({ S14852 }),
  .A3({ S15191 }),
  .ZN({ S15192 })
);
NAND3_X1 #() 
NAND3_X1_2124_ (
  .A1({ S15192 }),
  .A2({ S15189 }),
  .A3({ S14919 }),
  .ZN({ S15193 })
);
NAND3_X1 #() 
NAND3_X1_2125_ (
  .A1({ S15185 }),
  .A2({ S15193 }),
  .A3({ S14823 }),
  .ZN({ S15194 })
);
NAND3_X1 #() 
NAND3_X1_2126_ (
  .A1({ S15194 }),
  .A2({ S15177 }),
  .A3({ S25957[287] }),
  .ZN({ S15195 })
);
NAND3_X1 #() 
NAND3_X1_2127_ (
  .A1({ S15166 }),
  .A2({ S15136 }),
  .A3({ S15195 }),
  .ZN({ S15196 })
);
NAND2_X1 #() 
NAND2_X1_1847_ (
  .A1({ S15142 }),
  .A2({ S15149 }),
  .ZN({ S15197 })
);
NAND2_X1 #() 
NAND2_X1_1848_ (
  .A1({ S15197 }),
  .A2({ S25957[286] }),
  .ZN({ S15199 })
);
AND2_X1 #() 
AND2_X1_111_ (
  .A1({ S15158 }),
  .A2({ S15156 }),
  .ZN({ S15200 })
);
OAI211_X1 #() 
OAI211_X1_673_ (
  .A({ S14919 }),
  .B({ S15161 }),
  .C1({ S15200 }),
  .C2({ S25957[284] }),
  .ZN({ S15201 })
);
NOR2_X1 #() 
NOR2_X1_442_ (
  .A1({ S14936 }),
  .A2({ S41 }),
  .ZN({ S15202 })
);
OAI21_X1 #() 
OAI21_X1_1011_ (
  .A({ S14852 }),
  .B1({ S15202 }),
  .B2({ S15092 }),
  .ZN({ S15203 })
);
NAND3_X1 #() 
NAND3_X1_2128_ (
  .A1({ S15203 }),
  .A2({ S25957[285] }),
  .A3({ S15152 }),
  .ZN({ S15204 })
);
NAND3_X1 #() 
NAND3_X1_2129_ (
  .A1({ S15201 }),
  .A2({ S15204 }),
  .A3({ S14823 }),
  .ZN({ S15205 })
);
AOI21_X1 #() 
AOI21_X1_1107_ (
  .A({ S25957[287] }),
  .B1({ S15205 }),
  .B2({ S15199 }),
  .ZN({ S15206 })
);
AND3_X1 #() 
AND3_X1_84_ (
  .A1({ S15194 }),
  .A2({ S15177 }),
  .A3({ S25957[287] }),
  .ZN({ S15207 })
);
OAI21_X1 #() 
OAI21_X1_1012_ (
  .A({ S25957[356] }),
  .B1({ S15207 }),
  .B2({ S15206 }),
  .ZN({ S15208 })
);
NAND3_X1 #() 
NAND3_X1_2130_ (
  .A1({ S15208 }),
  .A2({ S15196 }),
  .A3({ S25957[324] }),
  .ZN({ S15210 })
);
INV_X1 #() 
INV_X1_596_ (
  .A({ S25957[324] }),
  .ZN({ S15211 })
);
NAND3_X1 #() 
NAND3_X1_2131_ (
  .A1({ S15166 }),
  .A2({ S25957[356] }),
  .A3({ S15195 }),
  .ZN({ S15212 })
);
OAI21_X1 #() 
OAI21_X1_1013_ (
  .A({ S15136 }),
  .B1({ S15207 }),
  .B2({ S15206 }),
  .ZN({ S15213 })
);
NAND3_X1 #() 
NAND3_X1_2132_ (
  .A1({ S15213 }),
  .A2({ S15212 }),
  .A3({ S15211 }),
  .ZN({ S15214 })
);
NAND3_X1 #() 
NAND3_X1_2133_ (
  .A1({ S15210 }),
  .A2({ S15214 }),
  .A3({ S11332 }),
  .ZN({ S15215 })
);
NAND3_X1 #() 
NAND3_X1_2134_ (
  .A1({ S15213 }),
  .A2({ S15212 }),
  .A3({ S25957[324] }),
  .ZN({ S15216 })
);
NAND3_X1 #() 
NAND3_X1_2135_ (
  .A1({ S15208 }),
  .A2({ S15196 }),
  .A3({ S15211 }),
  .ZN({ S15217 })
);
NAND3_X1 #() 
NAND3_X1_2136_ (
  .A1({ S15216 }),
  .A2({ S15217 }),
  .A3({ S25957[388] }),
  .ZN({ S15218 })
);
AND2_X1 #() 
AND2_X1_112_ (
  .A1({ S15218 }),
  .A2({ S15215 }),
  .ZN({ S25957[132] })
);
NOR2_X1 #() 
NOR2_X1_443_ (
  .A1({ S12438 }),
  .A2({ S12437 }),
  .ZN({ S25957[291] })
);
NAND2_X1 #() 
NAND2_X1_1849_ (
  .A1({ S9512 }),
  .A2({ S9513 }),
  .ZN({ S25957[451] })
);
INV_X1 #() 
INV_X1_597_ (
  .A({ S25957[451] }),
  .ZN({ S15220 })
);
NAND3_X1 #() 
NAND3_X1_2137_ (
  .A1({ S14867 }),
  .A2({ S41 }),
  .A3({ S14983 }),
  .ZN({ S15221 })
);
NAND2_X1 #() 
NAND2_X1_1850_ (
  .A1({ S15221 }),
  .A2({ S15077 }),
  .ZN({ S15222 })
);
AND3_X1 #() 
AND3_X1_85_ (
  .A1({ S14969 }),
  .A2({ S14913 }),
  .A3({ S14852 }),
  .ZN({ S15223 })
);
AOI21_X1 #() 
AOI21_X1_1108_ (
  .A({ S15223 }),
  .B1({ S15222 }),
  .B2({ S25957[284] }),
  .ZN({ S15224 })
);
INV_X1 #() 
INV_X1_598_ (
  .A({ S49 }),
  .ZN({ S15225 })
);
OAI21_X1 #() 
OAI21_X1_1014_ (
  .A({ S25957[283] }),
  .B1({ S15225 }),
  .B2({ S14943 }),
  .ZN({ S15226 })
);
OAI21_X1 #() 
OAI21_X1_1015_ (
  .A({ S41 }),
  .B1({ S14887 }),
  .B2({ S15168 }),
  .ZN({ S15227 })
);
NAND3_X1 #() 
NAND3_X1_2138_ (
  .A1({ S15227 }),
  .A2({ S25957[284] }),
  .A3({ S15226 }),
  .ZN({ S15229 })
);
NAND2_X1 #() 
NAND2_X1_1851_ (
  .A1({ S14836 }),
  .A2({ S25957[283] }),
  .ZN({ S15230 })
);
NAND3_X1 #() 
NAND3_X1_2139_ (
  .A1({ S14976 }),
  .A2({ S41 }),
  .A3({ S14862 }),
  .ZN({ S15231 })
);
OAI211_X1 #() 
OAI211_X1_674_ (
  .A({ S15231 }),
  .B({ S14852 }),
  .C1({ S15230 }),
  .C2({ S14972 }),
  .ZN({ S15232 })
);
NAND3_X1 #() 
NAND3_X1_2140_ (
  .A1({ S15229 }),
  .A2({ S15232 }),
  .A3({ S25957[285] }),
  .ZN({ S15233 })
);
OAI211_X1 #() 
OAI211_X1_675_ (
  .A({ S25957[286] }),
  .B({ S15233 }),
  .C1({ S15224 }),
  .C2({ S25957[285] }),
  .ZN({ S15234 })
);
NAND3_X1 #() 
NAND3_X1_2141_ (
  .A1({ S14936 }),
  .A2({ S14987 }),
  .A3({ S25957[283] }),
  .ZN({ S15235 })
);
NAND2_X1 #() 
NAND2_X1_1852_ (
  .A1({ S14860 }),
  .A2({ S49 }),
  .ZN({ S15236 })
);
NAND3_X1 #() 
NAND3_X1_2142_ (
  .A1({ S15236 }),
  .A2({ S41 }),
  .A3({ S14836 }),
  .ZN({ S15237 })
);
NAND4_X1 #() 
NAND4_X1_263_ (
  .A1({ S14854 }),
  .A2({ S14842 }),
  .A3({ S25957[281] }),
  .A4({ S25957[283] }),
  .ZN({ S15238 })
);
AND2_X1 #() 
AND2_X1_113_ (
  .A1({ S15238 }),
  .A2({ S14852 }),
  .ZN({ S15240 })
);
AOI22_X1 #() 
AOI22_X1_247_ (
  .A1({ S15240 }),
  .A2({ S15237 }),
  .B1({ S15235 }),
  .B2({ S15182 }),
  .ZN({ S15241 })
);
NAND3_X1 #() 
NAND3_X1_2143_ (
  .A1({ S14853 }),
  .A2({ S14827 }),
  .A3({ S41 }),
  .ZN({ S15242 })
);
OAI211_X1 #() 
OAI211_X1_676_ (
  .A({ S25957[284] }),
  .B({ S15242 }),
  .C1({ S14864 }),
  .C2({ S41 }),
  .ZN({ S15243 })
);
AOI21_X1 #() 
AOI21_X1_1109_ (
  .A({ S25957[284] }),
  .B1({ S14932 }),
  .B2({ S49 }),
  .ZN({ S15244 })
);
OAI21_X1 #() 
OAI21_X1_1016_ (
  .A({ S15244 }),
  .B1({ S15103 }),
  .B2({ S14982 }),
  .ZN({ S15245 })
);
NAND3_X1 #() 
NAND3_X1_2144_ (
  .A1({ S15245 }),
  .A2({ S15243 }),
  .A3({ S14919 }),
  .ZN({ S15246 })
);
OAI211_X1 #() 
OAI211_X1_677_ (
  .A({ S14823 }),
  .B({ S15246 }),
  .C1({ S15241 }),
  .C2({ S14919 }),
  .ZN({ S15247 })
);
NAND3_X1 #() 
NAND3_X1_2145_ (
  .A1({ S15234 }),
  .A2({ S25957[287] }),
  .A3({ S15247 }),
  .ZN({ S15248 })
);
NAND2_X1 #() 
NAND2_X1_1853_ (
  .A1({ S15043 }),
  .A2({ S14830 }),
  .ZN({ S15249 })
);
AOI21_X1 #() 
AOI21_X1_1110_ (
  .A({ S25957[283] }),
  .B1({ S25957[281] }),
  .B2({ S14834 }),
  .ZN({ S15251 })
);
NAND2_X1 #() 
NAND2_X1_1854_ (
  .A1({ S15251 }),
  .A2({ S14862 }),
  .ZN({ S15252 })
);
AOI21_X1 #() 
AOI21_X1_1111_ (
  .A({ S25957[284] }),
  .B1({ S15252 }),
  .B2({ S15249 }),
  .ZN({ S15253 })
);
OAI21_X1 #() 
OAI21_X1_1017_ (
  .A({ S25957[284] }),
  .B1({ S14891 }),
  .B2({ S14853 }),
  .ZN({ S15254 })
);
AOI21_X1 #() 
AOI21_X1_1112_ (
  .A({ S15254 }),
  .B1({ S14885 }),
  .B2({ S14973 }),
  .ZN({ S15255 })
);
OAI21_X1 #() 
OAI21_X1_1018_ (
  .A({ S25957[285] }),
  .B1({ S15255 }),
  .B2({ S15253 }),
  .ZN({ S15256 })
);
NAND2_X1 #() 
NAND2_X1_1855_ (
  .A1({ S14836 }),
  .A2({ S25957[280] }),
  .ZN({ S15257 })
);
NAND2_X1 #() 
NAND2_X1_1856_ (
  .A1({ S15257 }),
  .A2({ S41 }),
  .ZN({ S15258 })
);
NOR2_X1 #() 
NOR2_X1_444_ (
  .A1({ S15258 }),
  .A2({ S14852 }),
  .ZN({ S15259 })
);
NAND3_X1 #() 
NAND3_X1_2146_ (
  .A1({ S14853 }),
  .A2({ S14827 }),
  .A3({ S14837 }),
  .ZN({ S15260 })
);
NAND2_X1 #() 
NAND2_X1_1857_ (
  .A1({ S15260 }),
  .A2({ S25957[283] }),
  .ZN({ S15262 })
);
NAND4_X1 #() 
NAND4_X1_264_ (
  .A1({ S14853 }),
  .A2({ S14845 }),
  .A3({ S25957[280] }),
  .A4({ S41 }),
  .ZN({ S15263 })
);
AOI21_X1 #() 
AOI21_X1_1113_ (
  .A({ S25957[284] }),
  .B1({ S15262 }),
  .B2({ S15263 }),
  .ZN({ S15264 })
);
OAI21_X1 #() 
OAI21_X1_1019_ (
  .A({ S14919 }),
  .B1({ S15264 }),
  .B2({ S15259 }),
  .ZN({ S15265 })
);
AOI21_X1 #() 
AOI21_X1_1114_ (
  .A({ S14823 }),
  .B1({ S15256 }),
  .B2({ S15265 }),
  .ZN({ S15266 })
);
OAI21_X1 #() 
OAI21_X1_1020_ (
  .A({ S25957[283] }),
  .B1({ S14842 }),
  .B2({ S25957[281] }),
  .ZN({ S15267 })
);
OAI211_X1 #() 
OAI211_X1_678_ (
  .A({ S25957[284] }),
  .B({ S15267 }),
  .C1({ S14878 }),
  .C2({ S25957[283] }),
  .ZN({ S15268 })
);
OAI211_X1 #() 
OAI211_X1_679_ (
  .A({ S14852 }),
  .B({ S25957[280] }),
  .C1({ S15251 }),
  .C2({ S14847 }),
  .ZN({ S15269 })
);
NAND3_X1 #() 
NAND3_X1_2147_ (
  .A1({ S15268 }),
  .A2({ S25957[285] }),
  .A3({ S15269 }),
  .ZN({ S15270 })
);
AOI21_X1 #() 
AOI21_X1_1115_ (
  .A({ S15016 }),
  .B1({ S15081 }),
  .B2({ S14862 }),
  .ZN({ S15271 })
);
NAND2_X1 #() 
NAND2_X1_1858_ (
  .A1({ S15139 }),
  .A2({ S25957[283] }),
  .ZN({ S15273 })
);
OAI211_X1 #() 
OAI211_X1_680_ (
  .A({ S14852 }),
  .B({ S15273 }),
  .C1({ S15271 }),
  .C2({ S25957[283] }),
  .ZN({ S15274 })
);
OAI21_X1 #() 
OAI21_X1_1021_ (
  .A({ S49 }),
  .B1({ S14935 }),
  .B2({ S25957[282] }),
  .ZN({ S15275 })
);
OAI211_X1 #() 
OAI211_X1_681_ (
  .A({ S25957[284] }),
  .B({ S15046 }),
  .C1({ S15275 }),
  .C2({ S41 }),
  .ZN({ S15276 })
);
NAND3_X1 #() 
NAND3_X1_2148_ (
  .A1({ S15274 }),
  .A2({ S14919 }),
  .A3({ S15276 }),
  .ZN({ S15277 })
);
AOI21_X1 #() 
AOI21_X1_1116_ (
  .A({ S25957[286] }),
  .B1({ S15277 }),
  .B2({ S15270 }),
  .ZN({ S15278 })
);
OAI21_X1 #() 
OAI21_X1_1022_ (
  .A({ S14822 }),
  .B1({ S15278 }),
  .B2({ S15266 }),
  .ZN({ S15279 })
);
AOI21_X1 #() 
AOI21_X1_1117_ (
  .A({ S15220 }),
  .B1({ S15279 }),
  .B2({ S15248 }),
  .ZN({ S15280 })
);
AND3_X1 #() 
AND3_X1_86_ (
  .A1({ S15279 }),
  .A2({ S15248 }),
  .A3({ S15220 }),
  .ZN({ S15281 })
);
OAI21_X1 #() 
OAI21_X1_1023_ (
  .A({ S25957[291] }),
  .B1({ S15281 }),
  .B2({ S15280 }),
  .ZN({ S15282 })
);
INV_X1 #() 
INV_X1_599_ (
  .A({ S25957[291] }),
  .ZN({ S15284 })
);
AND3_X1 #() 
AND3_X1_87_ (
  .A1({ S15234 }),
  .A2({ S25957[287] }),
  .A3({ S15247 }),
  .ZN({ S15285 })
);
NAND2_X1 #() 
NAND2_X1_1859_ (
  .A1({ S15252 }),
  .A2({ S15249 }),
  .ZN({ S15286 })
);
NAND2_X1 #() 
NAND2_X1_1860_ (
  .A1({ S15286 }),
  .A2({ S14852 }),
  .ZN({ S15287 })
);
OAI211_X1 #() 
OAI211_X1_682_ (
  .A({ S15287 }),
  .B({ S25957[285] }),
  .C1({ S14974 }),
  .C2({ S15254 }),
  .ZN({ S15288 })
);
INV_X1 #() 
INV_X1_600_ (
  .A({ S15259 }),
  .ZN({ S15289 })
);
NAND2_X1 #() 
NAND2_X1_1861_ (
  .A1({ S14874 }),
  .A2({ S15160 }),
  .ZN({ S15290 })
);
NAND3_X1 #() 
NAND3_X1_2149_ (
  .A1({ S15290 }),
  .A2({ S14919 }),
  .A3({ S15289 }),
  .ZN({ S15291 })
);
NAND3_X1 #() 
NAND3_X1_2150_ (
  .A1({ S15288 }),
  .A2({ S25957[286] }),
  .A3({ S15291 }),
  .ZN({ S15292 })
);
AND2_X1 #() 
AND2_X1_114_ (
  .A1({ S15139 }),
  .A2({ S25957[283] }),
  .ZN({ S15293 })
);
NOR3_X1 #() 
NOR3_X1_61_ (
  .A1({ S14869 }),
  .A2({ S15293 }),
  .A3({ S25957[284] }),
  .ZN({ S15294 })
);
NAND2_X1 #() 
NAND2_X1_1862_ (
  .A1({ S15276 }),
  .A2({ S14919 }),
  .ZN({ S15295 })
);
OAI21_X1 #() 
OAI21_X1_1024_ (
  .A({ S15270 }),
  .B1({ S15294 }),
  .B2({ S15295 }),
  .ZN({ S15296 })
);
NAND2_X1 #() 
NAND2_X1_1863_ (
  .A1({ S15296 }),
  .A2({ S14823 }),
  .ZN({ S15297 })
);
AOI21_X1 #() 
AOI21_X1_1118_ (
  .A({ S25957[287] }),
  .B1({ S15297 }),
  .B2({ S15292 }),
  .ZN({ S15298 })
);
OAI21_X1 #() 
OAI21_X1_1025_ (
  .A({ S25957[451] }),
  .B1({ S15285 }),
  .B2({ S15298 }),
  .ZN({ S15299 })
);
NAND3_X1 #() 
NAND3_X1_2151_ (
  .A1({ S15279 }),
  .A2({ S15220 }),
  .A3({ S15248 }),
  .ZN({ S15300 })
);
NAND3_X1 #() 
NAND3_X1_2152_ (
  .A1({ S15299 }),
  .A2({ S15284 }),
  .A3({ S15300 }),
  .ZN({ S15301 })
);
NAND3_X1 #() 
NAND3_X1_2153_ (
  .A1({ S15282 }),
  .A2({ S25957[259] }),
  .A3({ S15301 }),
  .ZN({ S15302 })
);
OAI21_X1 #() 
OAI21_X1_1026_ (
  .A({ S15284 }),
  .B1({ S15281 }),
  .B2({ S15280 }),
  .ZN({ S15303 })
);
NAND3_X1 #() 
NAND3_X1_2154_ (
  .A1({ S15299 }),
  .A2({ S25957[291] }),
  .A3({ S15300 }),
  .ZN({ S15305 })
);
NAND3_X1 #() 
NAND3_X1_2155_ (
  .A1({ S15303 }),
  .A2({ S38 }),
  .A3({ S15305 }),
  .ZN({ S15306 })
);
NAND2_X1 #() 
NAND2_X1_1864_ (
  .A1({ S15302 }),
  .A2({ S15306 }),
  .ZN({ S51 })
);
AND2_X1 #() 
AND2_X1_115_ (
  .A1({ S15306 }),
  .A2({ S15302 }),
  .ZN({ S25957[131] })
);
NAND2_X1 #() 
NAND2_X1_1865_ (
  .A1({ S15160 }),
  .A2({ S14852 }),
  .ZN({ S15307 })
);
AOI21_X1 #() 
AOI21_X1_1119_ (
  .A({ S25957[283] }),
  .B1({ S14936 }),
  .B2({ S14830 }),
  .ZN({ S15308 })
);
NAND3_X1 #() 
NAND3_X1_2156_ (
  .A1({ S14866 }),
  .A2({ S25957[283] }),
  .A3({ S25957[282] }),
  .ZN({ S15309 })
);
OAI211_X1 #() 
OAI211_X1_683_ (
  .A({ S25957[284] }),
  .B({ S15309 }),
  .C1({ S14925 }),
  .C2({ S25957[283] }),
  .ZN({ S15310 })
);
OAI211_X1 #() 
OAI211_X1_684_ (
  .A({ S15310 }),
  .B({ S25957[285] }),
  .C1({ S15307 }),
  .C2({ S15308 }),
  .ZN({ S15311 })
);
NAND2_X1 #() 
NAND2_X1_1866_ (
  .A1({ S14972 }),
  .A2({ S41 }),
  .ZN({ S15312 })
);
NAND3_X1 #() 
NAND3_X1_2157_ (
  .A1({ S15312 }),
  .A2({ S15068 }),
  .A3({ S15183 }),
  .ZN({ S15314 })
);
AOI21_X1 #() 
AOI21_X1_1120_ (
  .A({ S15056 }),
  .B1({ S15314 }),
  .B2({ S25957[284] }),
  .ZN({ S15315 })
);
OAI211_X1 #() 
OAI211_X1_685_ (
  .A({ S15311 }),
  .B({ S25957[286] }),
  .C1({ S15315 }),
  .C2({ S25957[285] }),
  .ZN({ S15316 })
);
NOR2_X1 #() 
NOR2_X1_445_ (
  .A1({ S14842 }),
  .A2({ S25957[281] }),
  .ZN({ S15317 })
);
AOI21_X1 #() 
AOI21_X1_1121_ (
  .A({ S15317 }),
  .B1({ S14996 }),
  .B2({ S14842 }),
  .ZN({ S15318 })
);
NAND4_X1 #() 
NAND4_X1_265_ (
  .A1({ S15180 }),
  .A2({ S14848 }),
  .A3({ S14944 }),
  .A4({ S14852 }),
  .ZN({ S15319 })
);
OAI211_X1 #() 
OAI211_X1_686_ (
  .A({ S25957[285] }),
  .B({ S15319 }),
  .C1({ S15318 }),
  .C2({ S14852 }),
  .ZN({ S15320 })
);
OAI21_X1 #() 
OAI21_X1_1027_ (
  .A({ S15249 }),
  .B1({ S15081 }),
  .B2({ S15095 }),
  .ZN({ S15321 })
);
NAND2_X1 #() 
NAND2_X1_1867_ (
  .A1({ S14830 }),
  .A2({ S25957[283] }),
  .ZN({ S15322 })
);
OAI211_X1 #() 
OAI211_X1_687_ (
  .A({ S25957[284] }),
  .B({ S15322 }),
  .C1({ S15099 }),
  .C2({ S25957[283] }),
  .ZN({ S15323 })
);
OAI211_X1 #() 
OAI211_X1_688_ (
  .A({ S15323 }),
  .B({ S14919 }),
  .C1({ S25957[284] }),
  .C2({ S15321 }),
  .ZN({ S15325 })
);
NAND3_X1 #() 
NAND3_X1_2158_ (
  .A1({ S15325 }),
  .A2({ S15320 }),
  .A3({ S14823 }),
  .ZN({ S15326 })
);
NAND3_X1 #() 
NAND3_X1_2159_ (
  .A1({ S15316 }),
  .A2({ S25957[287] }),
  .A3({ S15326 }),
  .ZN({ S15327 })
);
AOI21_X1 #() 
AOI21_X1_1122_ (
  .A({ S25957[283] }),
  .B1({ S14987 }),
  .B2({ S14935 }),
  .ZN({ S15328 })
);
NAND2_X1 #() 
NAND2_X1_1868_ (
  .A1({ S14932 }),
  .A2({ S14866 }),
  .ZN({ S15329 })
);
NAND3_X1 #() 
NAND3_X1_2160_ (
  .A1({ S15156 }),
  .A2({ S15329 }),
  .A3({ S25957[284] }),
  .ZN({ S15330 })
);
OAI21_X1 #() 
OAI21_X1_1028_ (
  .A({ S14852 }),
  .B1({ S14855 }),
  .B2({ S15011 }),
  .ZN({ S15331 })
);
OAI211_X1 #() 
OAI211_X1_689_ (
  .A({ S15330 }),
  .B({ S25957[285] }),
  .C1({ S15328 }),
  .C2({ S15331 }),
  .ZN({ S15332 })
);
OAI211_X1 #() 
OAI211_X1_690_ (
  .A({ S41 }),
  .B({ S14853 }),
  .C1({ S14884 }),
  .C2({ S48 }),
  .ZN({ S15333 })
);
OAI211_X1 #() 
OAI211_X1_691_ (
  .A({ S15333 }),
  .B({ S25957[284] }),
  .C1({ S41 }),
  .C2({ S15178 }),
  .ZN({ S15334 })
);
NAND2_X1 #() 
NAND2_X1_1869_ (
  .A1({ S15028 }),
  .A2({ S49 }),
  .ZN({ S15336 })
);
NAND2_X1 #() 
NAND2_X1_1870_ (
  .A1({ S15336 }),
  .A2({ S25957[283] }),
  .ZN({ S15337 })
);
NOR2_X1 #() 
NOR2_X1_446_ (
  .A1({ S14911 }),
  .A2({ S14836 }),
  .ZN({ S15338 })
);
OAI21_X1 #() 
OAI21_X1_1029_ (
  .A({ S41 }),
  .B1({ S15338 }),
  .B2({ S15317 }),
  .ZN({ S15339 })
);
NAND3_X1 #() 
NAND3_X1_2161_ (
  .A1({ S15337 }),
  .A2({ S15339 }),
  .A3({ S14852 }),
  .ZN({ S15340 })
);
NAND3_X1 #() 
NAND3_X1_2162_ (
  .A1({ S15334 }),
  .A2({ S15340 }),
  .A3({ S14919 }),
  .ZN({ S15341 })
);
NAND3_X1 #() 
NAND3_X1_2163_ (
  .A1({ S15341 }),
  .A2({ S14823 }),
  .A3({ S15332 }),
  .ZN({ S15342 })
);
AOI21_X1 #() 
AOI21_X1_1123_ (
  .A({ S25957[284] }),
  .B1({ S14993 }),
  .B2({ S25957[283] }),
  .ZN({ S15343 })
);
OAI21_X1 #() 
OAI21_X1_1030_ (
  .A({ S25957[283] }),
  .B1({ S15103 }),
  .B2({ S14883 }),
  .ZN({ S15344 })
);
AOI22_X1 #() 
AOI22_X1_248_ (
  .A1({ S15344 }),
  .A2({ S14977 }),
  .B1({ S15343 }),
  .B2({ S15095 }),
  .ZN({ S15345 })
);
NAND2_X1 #() 
NAND2_X1_1871_ (
  .A1({ S14827 }),
  .A2({ S14841 }),
  .ZN({ S15347 })
);
NAND2_X1 #() 
NAND2_X1_1872_ (
  .A1({ S15347 }),
  .A2({ S41 }),
  .ZN({ S15348 })
);
INV_X1 #() 
INV_X1_601_ (
  .A({ S15348 }),
  .ZN({ S15349 })
);
NAND2_X1 #() 
NAND2_X1_1873_ (
  .A1({ S14911 }),
  .A2({ S25957[283] }),
  .ZN({ S15350 })
);
NAND2_X1 #() 
NAND2_X1_1874_ (
  .A1({ S15016 }),
  .A2({ S25957[281] }),
  .ZN({ S15351 })
);
NAND3_X1 #() 
NAND3_X1_2164_ (
  .A1({ S15351 }),
  .A2({ S15350 }),
  .A3({ S14845 }),
  .ZN({ S15352 })
);
OAI221_X1 #() 
OAI221_X1_41_ (
  .A({ S14919 }),
  .B1({ S15352 }),
  .B2({ S14852 }),
  .C1({ S15148 }),
  .C2({ S15349 }),
  .ZN({ S15353 })
);
OAI211_X1 #() 
OAI211_X1_692_ (
  .A({ S25957[286] }),
  .B({ S15353 }),
  .C1({ S15345 }),
  .C2({ S14919 }),
  .ZN({ S15354 })
);
NAND3_X1 #() 
NAND3_X1_2165_ (
  .A1({ S15354 }),
  .A2({ S15342 }),
  .A3({ S14822 }),
  .ZN({ S15355 })
);
NAND3_X1 #() 
NAND3_X1_2166_ (
  .A1({ S15355 }),
  .A2({ S15327 }),
  .A3({ S25957[640] }),
  .ZN({ S15356 })
);
OAI21_X1 #() 
OAI21_X1_1031_ (
  .A({ S15310 }),
  .B1({ S15307 }),
  .B2({ S15308 }),
  .ZN({ S15358 })
);
NAND2_X1 #() 
NAND2_X1_1875_ (
  .A1({ S15358 }),
  .A2({ S25957[285] }),
  .ZN({ S15359 })
);
NAND2_X1 #() 
NAND2_X1_1876_ (
  .A1({ S15314 }),
  .A2({ S25957[284] }),
  .ZN({ S15360 })
);
NOR2_X1 #() 
NOR2_X1_447_ (
  .A1({ S15056 }),
  .A2({ S25957[285] }),
  .ZN({ S15361 })
);
NAND2_X1 #() 
NAND2_X1_1877_ (
  .A1({ S15361 }),
  .A2({ S15360 }),
  .ZN({ S15362 })
);
NAND3_X1 #() 
NAND3_X1_2167_ (
  .A1({ S15359 }),
  .A2({ S15362 }),
  .A3({ S25957[286] }),
  .ZN({ S15363 })
);
NAND2_X1 #() 
NAND2_X1_1878_ (
  .A1({ S15318 }),
  .A2({ S25957[284] }),
  .ZN({ S15364 })
);
INV_X1 #() 
INV_X1_602_ (
  .A({ S15180 }),
  .ZN({ S15365 })
);
OAI21_X1 #() 
OAI21_X1_1032_ (
  .A({ S14852 }),
  .B1({ S15365 }),
  .B2({ S15172 }),
  .ZN({ S15366 })
);
NAND3_X1 #() 
NAND3_X1_2168_ (
  .A1({ S15364 }),
  .A2({ S25957[285] }),
  .A3({ S15366 }),
  .ZN({ S15367 })
);
NAND2_X1 #() 
NAND2_X1_1879_ (
  .A1({ S15024 }),
  .A2({ S15146 }),
  .ZN({ S15369 })
);
NAND2_X1 #() 
NAND2_X1_1880_ (
  .A1({ S15321 }),
  .A2({ S14852 }),
  .ZN({ S15370 })
);
NAND3_X1 #() 
NAND3_X1_2169_ (
  .A1({ S15370 }),
  .A2({ S14919 }),
  .A3({ S15369 }),
  .ZN({ S15371 })
);
NAND3_X1 #() 
NAND3_X1_2170_ (
  .A1({ S15367 }),
  .A2({ S15371 }),
  .A3({ S14823 }),
  .ZN({ S15372 })
);
NAND3_X1 #() 
NAND3_X1_2171_ (
  .A1({ S15363 }),
  .A2({ S15372 }),
  .A3({ S25957[287] }),
  .ZN({ S15373 })
);
NAND2_X1 #() 
NAND2_X1_1881_ (
  .A1({ S15352 }),
  .A2({ S25957[284] }),
  .ZN({ S15374 })
);
AOI22_X1 #() 
AOI22_X1_249_ (
  .A1({ S14861 }),
  .A2({ S15053 }),
  .B1({ S15347 }),
  .B2({ S41 }),
  .ZN({ S15375 })
);
OAI211_X1 #() 
OAI211_X1_693_ (
  .A({ S15374 }),
  .B({ S14919 }),
  .C1({ S15375 }),
  .C2({ S25957[284] }),
  .ZN({ S15376 })
);
AND2_X1 #() 
AND2_X1_116_ (
  .A1({ S15343 }),
  .A2({ S15095 }),
  .ZN({ S15377 })
);
AOI21_X1 #() 
AOI21_X1_1124_ (
  .A({ S41 }),
  .B1({ S15236 }),
  .B2({ S14882 }),
  .ZN({ S15378 })
);
OAI21_X1 #() 
OAI21_X1_1033_ (
  .A({ S25957[285] }),
  .B1({ S15378 }),
  .B2({ S14978 }),
  .ZN({ S15380 })
);
OAI211_X1 #() 
OAI211_X1_694_ (
  .A({ S15376 }),
  .B({ S25957[286] }),
  .C1({ S15380 }),
  .C2({ S15377 }),
  .ZN({ S15381 })
);
AOI21_X1 #() 
AOI21_X1_1125_ (
  .A({ S41 }),
  .B1({ S14863 }),
  .B2({ S14862 }),
  .ZN({ S15382 })
);
AOI21_X1 #() 
AOI21_X1_1126_ (
  .A({ S25957[283] }),
  .B1({ S15347 }),
  .B2({ S15028 }),
  .ZN({ S15383 })
);
OAI21_X1 #() 
OAI21_X1_1034_ (
  .A({ S25957[284] }),
  .B1({ S15383 }),
  .B2({ S15382 }),
  .ZN({ S15384 })
);
NAND2_X1 #() 
NAND2_X1_1882_ (
  .A1({ S14996 }),
  .A2({ S14987 }),
  .ZN({ S15385 })
);
OAI211_X1 #() 
OAI211_X1_695_ (
  .A({ S15385 }),
  .B({ S14852 }),
  .C1({ S41 }),
  .C2({ S15336 }),
  .ZN({ S15386 })
);
NAND3_X1 #() 
NAND3_X1_2172_ (
  .A1({ S15386 }),
  .A2({ S15384 }),
  .A3({ S14919 }),
  .ZN({ S15387 })
);
OAI21_X1 #() 
OAI21_X1_1035_ (
  .A({ S15330 }),
  .B1({ S15328 }),
  .B2({ S15331 }),
  .ZN({ S15388 })
);
AOI21_X1 #() 
AOI21_X1_1127_ (
  .A({ S25957[286] }),
  .B1({ S15388 }),
  .B2({ S25957[285] }),
  .ZN({ S15389 })
);
NAND2_X1 #() 
NAND2_X1_1883_ (
  .A1({ S15389 }),
  .A2({ S15387 }),
  .ZN({ S15391 })
);
NAND3_X1 #() 
NAND3_X1_2173_ (
  .A1({ S15391 }),
  .A2({ S15381 }),
  .A3({ S14822 }),
  .ZN({ S15392 })
);
NAND3_X1 #() 
NAND3_X1_2174_ (
  .A1({ S15373 }),
  .A2({ S15392 }),
  .A3({ S5479 }),
  .ZN({ S15393 })
);
AND2_X1 #() 
AND2_X1_117_ (
  .A1({ S15393 }),
  .A2({ S15356 }),
  .ZN({ S25957[128] })
);
NAND2_X1 #() 
NAND2_X1_1884_ (
  .A1({ S6821 }),
  .A2({ S6825 }),
  .ZN({ S25957[545] })
);
XNOR2_X1 #() 
XNOR2_X1_63_ (
  .A({ S12518 }),
  .B({ S25957[545] }),
  .ZN({ S25957[417] })
);
NAND2_X1 #() 
NAND2_X1_1885_ (
  .A1({ S12570 }),
  .A2({ S12573 }),
  .ZN({ S15394 })
);
NAND2_X1 #() 
NAND2_X1_1886_ (
  .A1({ S15394 }),
  .A2({ S25957[417] }),
  .ZN({ S15395 })
);
OR2_X1 #() 
OR2_X1_27_ (
  .A1({ S15394 }),
  .A2({ S25957[417] }),
  .ZN({ S15396 })
);
NAND2_X1 #() 
NAND2_X1_1887_ (
  .A1({ S15396 }),
  .A2({ S15395 }),
  .ZN({ S25957[289] })
);
AOI21_X1 #() 
AOI21_X1_1128_ (
  .A({ S41 }),
  .B1({ S14867 }),
  .B2({ S14837 }),
  .ZN({ S15398 })
);
NAND3_X1 #() 
NAND3_X1_2175_ (
  .A1({ S15252 }),
  .A2({ S14852 }),
  .A3({ S15084 }),
  .ZN({ S15399 })
);
OAI211_X1 #() 
OAI211_X1_696_ (
  .A({ S15399 }),
  .B({ S25957[285] }),
  .C1({ S15398 }),
  .C2({ S14844 }),
  .ZN({ S15400 })
);
NAND2_X1 #() 
NAND2_X1_1888_ (
  .A1({ S14897 }),
  .A2({ S25957[283] }),
  .ZN({ S15401 })
);
NAND3_X1 #() 
NAND3_X1_2176_ (
  .A1({ S15351 }),
  .A2({ S41 }),
  .A3({ S14845 }),
  .ZN({ S15402 })
);
NAND3_X1 #() 
NAND3_X1_2177_ (
  .A1({ S15402 }),
  .A2({ S25957[284] }),
  .A3({ S15401 }),
  .ZN({ S15403 })
);
NAND2_X1 #() 
NAND2_X1_1889_ (
  .A1({ S15190 }),
  .A2({ S14852 }),
  .ZN({ S15404 })
);
OAI211_X1 #() 
OAI211_X1_697_ (
  .A({ S14919 }),
  .B({ S15403 }),
  .C1({ S15404 }),
  .C2({ S14865 }),
  .ZN({ S15405 })
);
NAND3_X1 #() 
NAND3_X1_2178_ (
  .A1({ S15405 }),
  .A2({ S14823 }),
  .A3({ S15400 }),
  .ZN({ S15406 })
);
NAND3_X1 #() 
NAND3_X1_2179_ (
  .A1({ S14830 }),
  .A2({ S14911 }),
  .A3({ S41 }),
  .ZN({ S15407 })
);
OAI211_X1 #() 
OAI211_X1_698_ (
  .A({ S25957[284] }),
  .B({ S15407 }),
  .C1({ S14878 }),
  .C2({ S15045 }),
  .ZN({ S15409 })
);
INV_X1 #() 
INV_X1_603_ (
  .A({ S15257 }),
  .ZN({ S15410 })
);
NAND3_X1 #() 
NAND3_X1_2180_ (
  .A1({ S14935 }),
  .A2({ S25957[283] }),
  .A3({ S14842 }),
  .ZN({ S15411 })
);
OAI211_X1 #() 
OAI211_X1_699_ (
  .A({ S15411 }),
  .B({ S14852 }),
  .C1({ S15410 }),
  .C2({ S14948 }),
  .ZN({ S15412 })
);
NAND3_X1 #() 
NAND3_X1_2181_ (
  .A1({ S15409 }),
  .A2({ S15412 }),
  .A3({ S14919 }),
  .ZN({ S15413 })
);
OAI21_X1 #() 
OAI21_X1_1036_ (
  .A({ S14852 }),
  .B1({ S14887 }),
  .B2({ S25957[283] }),
  .ZN({ S15414 })
);
OAI211_X1 #() 
OAI211_X1_700_ (
  .A({ S15077 }),
  .B({ S25957[284] }),
  .C1({ S14847 }),
  .C2({ S14848 }),
  .ZN({ S15415 })
);
OAI211_X1 #() 
OAI211_X1_701_ (
  .A({ S25957[285] }),
  .B({ S15415 }),
  .C1({ S15378 }),
  .C2({ S15414 }),
  .ZN({ S15416 })
);
NAND3_X1 #() 
NAND3_X1_2182_ (
  .A1({ S15416 }),
  .A2({ S25957[286] }),
  .A3({ S15413 }),
  .ZN({ S15417 })
);
NAND3_X1 #() 
NAND3_X1_2183_ (
  .A1({ S15406 }),
  .A2({ S25957[287] }),
  .A3({ S15417 }),
  .ZN({ S15418 })
);
NAND2_X1 #() 
NAND2_X1_1890_ (
  .A1({ S15275 }),
  .A2({ S25957[283] }),
  .ZN({ S15420 })
);
NAND2_X1 #() 
NAND2_X1_1891_ (
  .A1({ S15172 }),
  .A2({ S14854 }),
  .ZN({ S15421 })
);
NAND3_X1 #() 
NAND3_X1_2184_ (
  .A1({ S15420 }),
  .A2({ S15421 }),
  .A3({ S25957[284] }),
  .ZN({ S15422 })
);
NAND2_X1 #() 
NAND2_X1_1892_ (
  .A1({ S14976 }),
  .A2({ S14854 }),
  .ZN({ S15423 })
);
AOI21_X1 #() 
AOI21_X1_1129_ (
  .A({ S14919 }),
  .B1({ S15423 }),
  .B2({ S15091 }),
  .ZN({ S15424 })
);
NAND2_X1 #() 
NAND2_X1_1893_ (
  .A1({ S15422 }),
  .A2({ S15424 }),
  .ZN({ S15425 })
);
INV_X1 #() 
INV_X1_604_ (
  .A({ S15028 }),
  .ZN({ S15426 })
);
OAI21_X1 #() 
OAI21_X1_1037_ (
  .A({ S25957[284] }),
  .B1({ S15426 }),
  .B2({ S14948 }),
  .ZN({ S15427 })
);
NAND3_X1 #() 
NAND3_X1_2185_ (
  .A1({ S14967 }),
  .A2({ S15068 }),
  .A3({ S14852 }),
  .ZN({ S15428 })
);
OAI211_X1 #() 
OAI211_X1_702_ (
  .A({ S14919 }),
  .B({ S15428 }),
  .C1({ S15378 }),
  .C2({ S15427 }),
  .ZN({ S15429 })
);
NAND3_X1 #() 
NAND3_X1_2186_ (
  .A1({ S15429 }),
  .A2({ S15425 }),
  .A3({ S25957[286] }),
  .ZN({ S15431 })
);
NAND3_X1 #() 
NAND3_X1_2187_ (
  .A1({ S15263 }),
  .A2({ S14852 }),
  .A3({ S14940 }),
  .ZN({ S15432 })
);
NAND3_X1 #() 
NAND3_X1_2188_ (
  .A1({ S15169 }),
  .A2({ S14946 }),
  .A3({ S25957[284] }),
  .ZN({ S15433 })
);
NAND3_X1 #() 
NAND3_X1_2189_ (
  .A1({ S15433 }),
  .A2({ S14919 }),
  .A3({ S15432 }),
  .ZN({ S15434 })
);
AOI21_X1 #() 
AOI21_X1_1130_ (
  .A({ S14852 }),
  .B1({ S15238 }),
  .B2({ S15173 }),
  .ZN({ S15435 })
);
OAI21_X1 #() 
OAI21_X1_1038_ (
  .A({ S25957[285] }),
  .B1({ S14874 }),
  .B2({ S15435 }),
  .ZN({ S15436 })
);
NAND3_X1 #() 
NAND3_X1_2190_ (
  .A1({ S15434 }),
  .A2({ S15436 }),
  .A3({ S14823 }),
  .ZN({ S15437 })
);
NAND3_X1 #() 
NAND3_X1_2191_ (
  .A1({ S15431 }),
  .A2({ S15437 }),
  .A3({ S14822 }),
  .ZN({ S15438 })
);
NAND3_X1 #() 
NAND3_X1_2192_ (
  .A1({ S15418 }),
  .A2({ S15438 }),
  .A3({ S25957[449] }),
  .ZN({ S15439 })
);
NAND2_X1 #() 
NAND2_X1_1894_ (
  .A1({ S15418 }),
  .A2({ S15438 }),
  .ZN({ S15440 })
);
NAND2_X1 #() 
NAND2_X1_1895_ (
  .A1({ S15440 }),
  .A2({ S12518 }),
  .ZN({ S15442 })
);
AOI21_X1 #() 
AOI21_X1_1131_ (
  .A({ S25957[289] }),
  .B1({ S15442 }),
  .B2({ S15439 }),
  .ZN({ S15443 })
);
INV_X1 #() 
INV_X1_605_ (
  .A({ S25957[289] }),
  .ZN({ S15444 })
);
INV_X1 #() 
INV_X1_606_ (
  .A({ S15439 }),
  .ZN({ S15445 })
);
AOI21_X1 #() 
AOI21_X1_1132_ (
  .A({ S25957[449] }),
  .B1({ S15418 }),
  .B2({ S15438 }),
  .ZN({ S15446 })
);
NOR3_X1 #() 
NOR3_X1_62_ (
  .A1({ S15445 }),
  .A2({ S15446 }),
  .A3({ S15444 }),
  .ZN({ S15447 })
);
OAI21_X1 #() 
OAI21_X1_1039_ (
  .A({ S25957[257] }),
  .B1({ S15447 }),
  .B2({ S15443 }),
  .ZN({ S15448 })
);
OAI21_X1 #() 
OAI21_X1_1040_ (
  .A({ S15444 }),
  .B1({ S15445 }),
  .B2({ S15446 }),
  .ZN({ S15449 })
);
NAND3_X1 #() 
NAND3_X1_2193_ (
  .A1({ S15442 }),
  .A2({ S25957[289] }),
  .A3({ S15439 }),
  .ZN({ S15450 })
);
NAND3_X1 #() 
NAND3_X1_2194_ (
  .A1({ S15449 }),
  .A2({ S15450 }),
  .A3({ S14141 }),
  .ZN({ S15451 })
);
NAND2_X1 #() 
NAND2_X1_1896_ (
  .A1({ S15448 }),
  .A2({ S15451 }),
  .ZN({ S25957[129] })
);
AOI22_X1 #() 
AOI22_X1_250_ (
  .A1({ S14830 }),
  .A2({ S41 }),
  .B1({ S14851 }),
  .B2({ S14850 }),
  .ZN({ S15453 })
);
OAI21_X1 #() 
OAI21_X1_1041_ (
  .A({ S15453 }),
  .B1({ S15099 }),
  .B2({ S15017 }),
  .ZN({ S15454 })
);
NAND2_X1 #() 
NAND2_X1_1897_ (
  .A1({ S14872 }),
  .A2({ S25957[284] }),
  .ZN({ S15455 })
);
OAI211_X1 #() 
OAI211_X1_703_ (
  .A({ S15454 }),
  .B({ S25957[285] }),
  .C1({ S15308 }),
  .C2({ S15455 }),
  .ZN({ S15456 })
);
NAND2_X1 #() 
NAND2_X1_1898_ (
  .A1({ S14862 }),
  .A2({ S25957[282] }),
  .ZN({ S15457 })
);
NAND3_X1 #() 
NAND3_X1_2195_ (
  .A1({ S14936 }),
  .A2({ S25957[283] }),
  .A3({ S15457 }),
  .ZN({ S15458 })
);
NAND2_X1 #() 
NAND2_X1_1899_ (
  .A1({ S15458 }),
  .A2({ S15101 }),
  .ZN({ S15459 })
);
OAI211_X1 #() 
OAI211_X1_704_ (
  .A({ S15183 }),
  .B({ S14852 }),
  .C1({ S14982 }),
  .C2({ S15168 }),
  .ZN({ S15460 })
);
NAND3_X1 #() 
NAND3_X1_2196_ (
  .A1({ S15459 }),
  .A2({ S15460 }),
  .A3({ S14919 }),
  .ZN({ S15461 })
);
NAND3_X1 #() 
NAND3_X1_2197_ (
  .A1({ S15461 }),
  .A2({ S15456 }),
  .A3({ S25957[286] }),
  .ZN({ S15463 })
);
OAI211_X1 #() 
OAI211_X1_705_ (
  .A({ S14866 }),
  .B({ S25957[283] }),
  .C1({ S14862 }),
  .C2({ S14834 }),
  .ZN({ S15464 })
);
OAI211_X1 #() 
OAI211_X1_706_ (
  .A({ S15464 }),
  .B({ S14852 }),
  .C1({ S25957[283] }),
  .C2({ S14831 }),
  .ZN({ S15465 })
);
OAI211_X1 #() 
OAI211_X1_707_ (
  .A({ S15263 }),
  .B({ S25957[284] }),
  .C1({ S41 }),
  .C2({ S15257 }),
  .ZN({ S15466 })
);
NAND3_X1 #() 
NAND3_X1_2198_ (
  .A1({ S15465 }),
  .A2({ S15466 }),
  .A3({ S25957[285] }),
  .ZN({ S15467 })
);
INV_X1 #() 
INV_X1_607_ (
  .A({ S15053 }),
  .ZN({ S15468 })
);
NOR2_X1 #() 
NOR2_X1_448_ (
  .A1({ S15468 }),
  .A2({ S14841 }),
  .ZN({ S15469 })
);
OAI21_X1 #() 
OAI21_X1_1042_ (
  .A({ S25957[284] }),
  .B1({ S14897 }),
  .B2({ S25957[283] }),
  .ZN({ S15470 })
);
OAI211_X1 #() 
OAI211_X1_708_ (
  .A({ S15023 }),
  .B({ S14852 }),
  .C1({ S14841 }),
  .C2({ S14913 }),
  .ZN({ S15471 })
);
OAI211_X1 #() 
OAI211_X1_709_ (
  .A({ S15471 }),
  .B({ S14919 }),
  .C1({ S15469 }),
  .C2({ S15470 }),
  .ZN({ S15472 })
);
NAND3_X1 #() 
NAND3_X1_2199_ (
  .A1({ S15467 }),
  .A2({ S15472 }),
  .A3({ S14823 }),
  .ZN({ S15474 })
);
NAND3_X1 #() 
NAND3_X1_2200_ (
  .A1({ S15463 }),
  .A2({ S25957[287] }),
  .A3({ S15474 }),
  .ZN({ S15475 })
);
OAI21_X1 #() 
OAI21_X1_1043_ (
  .A({ S14852 }),
  .B1({ S14897 }),
  .B2({ S14891 }),
  .ZN({ S15476 })
);
AOI21_X1 #() 
AOI21_X1_1133_ (
  .A({ S15476 }),
  .B1({ S14931 }),
  .B2({ S14867 }),
  .ZN({ S15477 })
);
NAND3_X1 #() 
NAND3_X1_2201_ (
  .A1({ S14862 }),
  .A2({ S25957[283] }),
  .A3({ S14836 }),
  .ZN({ S15478 })
);
AOI21_X1 #() 
AOI21_X1_1134_ (
  .A({ S14852 }),
  .B1({ S15258 }),
  .B2({ S15478 }),
  .ZN({ S15479 })
);
OAI21_X1 #() 
OAI21_X1_1044_ (
  .A({ S25957[285] }),
  .B1({ S15477 }),
  .B2({ S15479 }),
  .ZN({ S15480 })
);
NAND3_X1 #() 
NAND3_X1_2202_ (
  .A1({ S14866 }),
  .A2({ S25957[283] }),
  .A3({ S14830 }),
  .ZN({ S15481 })
);
NAND4_X1 #() 
NAND4_X1_266_ (
  .A1({ S15312 }),
  .A2({ S14852 }),
  .A3({ S15183 }),
  .A4({ S15481 }),
  .ZN({ S15482 })
);
OAI21_X1 #() 
OAI21_X1_1045_ (
  .A({ S41 }),
  .B1({ S15257 }),
  .B2({ S14895 }),
  .ZN({ S15483 })
);
NAND2_X1 #() 
NAND2_X1_1900_ (
  .A1({ S15351 }),
  .A2({ S14871 }),
  .ZN({ S15485 })
);
NAND3_X1 #() 
NAND3_X1_2203_ (
  .A1({ S15483 }),
  .A2({ S15485 }),
  .A3({ S25957[284] }),
  .ZN({ S15486 })
);
NAND3_X1 #() 
NAND3_X1_2204_ (
  .A1({ S15482 }),
  .A2({ S14919 }),
  .A3({ S15486 }),
  .ZN({ S15487 })
);
NAND3_X1 #() 
NAND3_X1_2205_ (
  .A1({ S15480 }),
  .A2({ S15487 }),
  .A3({ S25957[286] }),
  .ZN({ S15488 })
);
NAND3_X1 #() 
NAND3_X1_2206_ (
  .A1({ S14936 }),
  .A2({ S41 }),
  .A3({ S14830 }),
  .ZN({ S15489 })
);
NAND2_X1 #() 
NAND2_X1_1901_ (
  .A1({ S15343 }),
  .A2({ S15489 }),
  .ZN({ S15490 })
);
AOI21_X1 #() 
AOI21_X1_1135_ (
  .A({ S14852 }),
  .B1({ S15053 }),
  .B2({ S25957[281] }),
  .ZN({ S15491 })
);
AOI21_X1 #() 
AOI21_X1_1136_ (
  .A({ S25957[285] }),
  .B1({ S15491 }),
  .B2({ S15186 }),
  .ZN({ S15492 })
);
NAND2_X1 #() 
NAND2_X1_1902_ (
  .A1({ S15490 }),
  .A2({ S15492 }),
  .ZN({ S15493 })
);
AOI211_X1 #() 
AOI211_X1_26_ (
  .A({ S25957[283] }),
  .B({ S14939 }),
  .C1({ S14860 }),
  .C2({ S49 }),
  .ZN({ S15494 })
);
AOI22_X1 #() 
AOI22_X1_251_ (
  .A1({ S15016 }),
  .A2({ S14910 }),
  .B1({ S14851 }),
  .B2({ S14850 }),
  .ZN({ S15496 })
);
NAND4_X1 #() 
NAND4_X1_267_ (
  .A1({ S15028 }),
  .A2({ S14837 }),
  .A3({ S14836 }),
  .A4({ S25957[283] }),
  .ZN({ S15497 })
);
NAND2_X1 #() 
NAND2_X1_1903_ (
  .A1({ S15497 }),
  .A2({ S15496 }),
  .ZN({ S15498 })
);
OAI21_X1 #() 
OAI21_X1_1046_ (
  .A({ S25957[284] }),
  .B1({ S15105 }),
  .B2({ S14943 }),
  .ZN({ S15499 })
);
OAI211_X1 #() 
OAI211_X1_710_ (
  .A({ S25957[285] }),
  .B({ S15498 }),
  .C1({ S15494 }),
  .C2({ S15499 }),
  .ZN({ S15500 })
);
NAND3_X1 #() 
NAND3_X1_2207_ (
  .A1({ S15493 }),
  .A2({ S15500 }),
  .A3({ S14823 }),
  .ZN({ S15501 })
);
NAND3_X1 #() 
NAND3_X1_2208_ (
  .A1({ S15488 }),
  .A2({ S15501 }),
  .A3({ S14822 }),
  .ZN({ S15502 })
);
AND3_X1 #() 
AND3_X1_88_ (
  .A1({ S15502 }),
  .A2({ S15475 }),
  .A3({ S12662 }),
  .ZN({ S15503 })
);
AOI21_X1 #() 
AOI21_X1_1137_ (
  .A({ S12662 }),
  .B1({ S15502 }),
  .B2({ S15475 }),
  .ZN({ S15504 })
);
OAI21_X1 #() 
OAI21_X1_1047_ (
  .A({ S25957[386] }),
  .B1({ S15503 }),
  .B2({ S15504 }),
  .ZN({ S15505 })
);
NAND3_X1 #() 
NAND3_X1_2209_ (
  .A1({ S15502 }),
  .A2({ S15475 }),
  .A3({ S12662 }),
  .ZN({ S15507 })
);
NAND2_X1 #() 
NAND2_X1_1904_ (
  .A1({ S15502 }),
  .A2({ S15475 }),
  .ZN({ S15508 })
);
NAND2_X1 #() 
NAND2_X1_1905_ (
  .A1({ S15508 }),
  .A2({ S25957[450] }),
  .ZN({ S15509 })
);
NAND3_X1 #() 
NAND3_X1_2210_ (
  .A1({ S15509 }),
  .A2({ S11298 }),
  .A3({ S15507 }),
  .ZN({ S15510 })
);
AND2_X1 #() 
AND2_X1_118_ (
  .A1({ S15505 }),
  .A2({ S15510 }),
  .ZN({ S25957[130] })
);
NAND3_X1 #() 
NAND3_X1_2211_ (
  .A1({ S11082 }),
  .A2({ S25957[400] }),
  .A3({ S11084 }),
  .ZN({ S15511 })
);
NAND3_X1 #() 
NAND3_X1_2212_ (
  .A1({ S11074 }),
  .A2({ S11081 }),
  .A3({ S11077 }),
  .ZN({ S15512 })
);
OAI21_X1 #() 
OAI21_X1_1048_ (
  .A({ S11179 }),
  .B1({ S11175 }),
  .B2({ S11174 }),
  .ZN({ S15513 })
);
NAND3_X1 #() 
NAND3_X1_2213_ (
  .A1({ S11183 }),
  .A2({ S25957[401] }),
  .A3({ S11184 }),
  .ZN({ S15514 })
);
NAND4_X1 #() 
NAND4_X1_268_ (
  .A1({ S15513 }),
  .A2({ S15511 }),
  .A3({ S15512 }),
  .A4({ S15514 }),
  .ZN({ S15515 })
);
INV_X1 #() 
INV_X1_608_ (
  .A({ S15515 }),
  .ZN({ S52 })
);
NAND4_X1 #() 
NAND4_X1_269_ (
  .A1({ S11176 }),
  .A2({ S11078 }),
  .A3({ S11085 }),
  .A4({ S11185 }),
  .ZN({ S53 })
);
NAND2_X1 #() 
NAND2_X1_1906_ (
  .A1({ S10652 }),
  .A2({ S10654 }),
  .ZN({ S15517 })
);
NAND4_X1 #() 
NAND4_X1_270_ (
  .A1({ S11176 }),
  .A2({ S15511 }),
  .A3({ S15512 }),
  .A4({ S11185 }),
  .ZN({ S15518 })
);
NAND2_X1 #() 
NAND2_X1_1907_ (
  .A1({ S15511 }),
  .A2({ S15512 }),
  .ZN({ S15519 })
);
NAND3_X1 #() 
NAND3_X1_2214_ (
  .A1({ S25957[274] }),
  .A2({ S25957[273] }),
  .A3({ S15519 }),
  .ZN({ S15520 })
);
NAND3_X1 #() 
NAND3_X1_2215_ (
  .A1({ S15520 }),
  .A2({ S25957[275] }),
  .A3({ S15518 }),
  .ZN({ S15521 })
);
OAI21_X1 #() 
OAI21_X1_1049_ (
  .A({ S11281 }),
  .B1({ S11273 }),
  .B2({ S11277 }),
  .ZN({ S15522 })
);
NAND3_X1 #() 
NAND3_X1_2216_ (
  .A1({ S11282 }),
  .A2({ S11283 }),
  .A3({ S25957[402] }),
  .ZN({ S15523 })
);
AOI22_X1 #() 
AOI22_X1_252_ (
  .A1({ S15522 }),
  .A2({ S15523 }),
  .B1({ S11085 }),
  .B2({ S11078 }),
  .ZN({ S15524 })
);
NAND2_X1 #() 
NAND2_X1_1908_ (
  .A1({ S15524 }),
  .A2({ S25957[273] }),
  .ZN({ S15526 })
);
NAND2_X1 #() 
NAND2_X1_1909_ (
  .A1({ S15513 }),
  .A2({ S15514 }),
  .ZN({ S15527 })
);
NAND3_X1 #() 
NAND3_X1_2217_ (
  .A1({ S25957[274] }),
  .A2({ S15527 }),
  .A3({ S15519 }),
  .ZN({ S15528 })
);
NAND2_X1 #() 
NAND2_X1_1910_ (
  .A1({ S15526 }),
  .A2({ S15528 }),
  .ZN({ S15529 })
);
OAI21_X1 #() 
OAI21_X1_1050_ (
  .A({ S15521 }),
  .B1({ S25957[275] }),
  .B2({ S15529 }),
  .ZN({ S15530 })
);
NAND4_X1 #() 
NAND4_X1_271_ (
  .A1({ S15522 }),
  .A2({ S15523 }),
  .A3({ S11078 }),
  .A4({ S11085 }),
  .ZN({ S15531 })
);
OAI211_X1 #() 
OAI211_X1_711_ (
  .A({ S15531 }),
  .B({ S25957[275] }),
  .C1({ S15518 }),
  .C2({ S25957[274] }),
  .ZN({ S15532 })
);
NAND4_X1 #() 
NAND4_X1_272_ (
  .A1({ S11278 }),
  .A2({ S11284 }),
  .A3({ S11078 }),
  .A4({ S11085 }),
  .ZN({ S15533 })
);
NAND2_X1 #() 
NAND2_X1_1911_ (
  .A1({ S15533 }),
  .A2({ S25957[273] }),
  .ZN({ S15534 })
);
OAI21_X1 #() 
OAI21_X1_1051_ (
  .A({ S15532 }),
  .B1({ S25957[275] }),
  .B2({ S15534 }),
  .ZN({ S15535 })
);
OAI21_X1 #() 
OAI21_X1_1052_ (
  .A({ S25957[277] }),
  .B1({ S15535 }),
  .B2({ S13772 }),
  .ZN({ S15537 })
);
AOI21_X1 #() 
AOI21_X1_1138_ (
  .A({ S15537 }),
  .B1({ S15530 }),
  .B2({ S13772 }),
  .ZN({ S15538 })
);
NAND4_X1 #() 
NAND4_X1_273_ (
  .A1({ S15513 }),
  .A2({ S11078 }),
  .A3({ S11085 }),
  .A4({ S15514 }),
  .ZN({ S15539 })
);
INV_X1 #() 
INV_X1_609_ (
  .A({ S15539 }),
  .ZN({ S15540 })
);
NAND4_X1 #() 
NAND4_X1_274_ (
  .A1({ S15522 }),
  .A2({ S11176 }),
  .A3({ S11185 }),
  .A4({ S15523 }),
  .ZN({ S15541 })
);
NAND4_X1 #() 
NAND4_X1_275_ (
  .A1({ S10985 }),
  .A2({ S10988 }),
  .A3({ S11176 }),
  .A4({ S11185 }),
  .ZN({ S15542 })
);
NAND2_X1 #() 
NAND2_X1_1912_ (
  .A1({ S25957[275] }),
  .A2({ S15519 }),
  .ZN({ S15543 })
);
NAND2_X1 #() 
NAND2_X1_1913_ (
  .A1({ S15543 }),
  .A2({ S15542 }),
  .ZN({ S15544 })
);
NAND2_X1 #() 
NAND2_X1_1914_ (
  .A1({ S15544 }),
  .A2({ S15541 }),
  .ZN({ S15545 })
);
OAI21_X1 #() 
OAI21_X1_1053_ (
  .A({ S15545 }),
  .B1({ S25957[275] }),
  .B2({ S15540 }),
  .ZN({ S15546 })
);
NAND2_X1 #() 
NAND2_X1_1915_ (
  .A1({ S15546 }),
  .A2({ S25957[276] }),
  .ZN({ S15548 })
);
NAND4_X1 #() 
NAND4_X1_276_ (
  .A1({ S15522 }),
  .A2({ S15523 }),
  .A3({ S15511 }),
  .A4({ S15512 }),
  .ZN({ S15549 })
);
INV_X1 #() 
INV_X1_610_ (
  .A({ S15549 }),
  .ZN({ S15550 })
);
NAND2_X1 #() 
NAND2_X1_1916_ (
  .A1({ S25957[274] }),
  .A2({ S25957[273] }),
  .ZN({ S15551 })
);
INV_X1 #() 
INV_X1_611_ (
  .A({ S15551 }),
  .ZN({ S15552 })
);
NAND2_X1 #() 
NAND2_X1_1917_ (
  .A1({ S15522 }),
  .A2({ S15523 }),
  .ZN({ S15553 })
);
NAND3_X1 #() 
NAND3_X1_2218_ (
  .A1({ S15553 }),
  .A2({ S15527 }),
  .A3({ S15519 }),
  .ZN({ S15554 })
);
NAND2_X1 #() 
NAND2_X1_1918_ (
  .A1({ S15554 }),
  .A2({ S13772 }),
  .ZN({ S15555 })
);
NOR3_X1 #() 
NOR3_X1_63_ (
  .A1({ S15555 }),
  .A2({ S15552 }),
  .A3({ S15550 }),
  .ZN({ S15556 })
);
OAI21_X1 #() 
OAI21_X1_1054_ (
  .A({ S15556 }),
  .B1({ S32 }),
  .B2({ S15518 }),
  .ZN({ S15557 })
);
AOI21_X1 #() 
AOI21_X1_1139_ (
  .A({ S25957[277] }),
  .B1({ S15548 }),
  .B2({ S15557 }),
  .ZN({ S15559 })
);
OAI21_X1 #() 
OAI21_X1_1055_ (
  .A({ S25957[278] }),
  .B1({ S15538 }),
  .B2({ S15559 }),
  .ZN({ S15560 })
);
AOI22_X1 #() 
AOI22_X1_253_ (
  .A1({ S10985 }),
  .A2({ S10988 }),
  .B1({ S11176 }),
  .B2({ S11185 }),
  .ZN({ S15561 })
);
INV_X1 #() 
INV_X1_612_ (
  .A({ S15561 }),
  .ZN({ S15562 })
);
OAI21_X1 #() 
OAI21_X1_1056_ (
  .A({ S25957[275] }),
  .B1({ S15550 }),
  .B2({ S15527 }),
  .ZN({ S15563 })
);
OAI21_X1 #() 
OAI21_X1_1057_ (
  .A({ S15563 }),
  .B1({ S15550 }),
  .B2({ S15562 }),
  .ZN({ S15564 })
);
NAND2_X1 #() 
NAND2_X1_1919_ (
  .A1({ S15564 }),
  .A2({ S25957[276] }),
  .ZN({ S15565 })
);
OAI21_X1 #() 
OAI21_X1_1058_ (
  .A({ S15565 }),
  .B1({ S15544 }),
  .B2({ S15555 }),
  .ZN({ S15566 })
);
NAND4_X1 #() 
NAND4_X1_277_ (
  .A1({ S11278 }),
  .A2({ S11176 }),
  .A3({ S11185 }),
  .A4({ S11284 }),
  .ZN({ S15567 })
);
INV_X1 #() 
INV_X1_613_ (
  .A({ S15567 }),
  .ZN({ S15568 })
);
AOI21_X1 #() 
AOI21_X1_1140_ (
  .A({ S25957[274] }),
  .B1({ S15518 }),
  .B2({ S15539 }),
  .ZN({ S15570 })
);
NAND2_X1 #() 
NAND2_X1_1920_ (
  .A1({ S15518 }),
  .A2({ S25957[274] }),
  .ZN({ S15571 })
);
INV_X1 #() 
INV_X1_614_ (
  .A({ S15571 }),
  .ZN({ S15572 })
);
OAI21_X1 #() 
OAI21_X1_1059_ (
  .A({ S32 }),
  .B1({ S15572 }),
  .B2({ S15570 }),
  .ZN({ S15573 })
);
OAI21_X1 #() 
OAI21_X1_1060_ (
  .A({ S15573 }),
  .B1({ S32 }),
  .B2({ S15568 }),
  .ZN({ S15574 })
);
NOR2_X1 #() 
NOR2_X1_449_ (
  .A1({ S15574 }),
  .A2({ S25957[276] }),
  .ZN({ S15575 })
);
NAND3_X1 #() 
NAND3_X1_2219_ (
  .A1({ S15515 }),
  .A2({ S53 }),
  .A3({ S15553 }),
  .ZN({ S15576 })
);
NAND3_X1 #() 
NAND3_X1_2220_ (
  .A1({ S15518 }),
  .A2({ S15539 }),
  .A3({ S25957[274] }),
  .ZN({ S15577 })
);
NAND3_X1 #() 
NAND3_X1_2221_ (
  .A1({ S15576 }),
  .A2({ S15577 }),
  .A3({ S25957[275] }),
  .ZN({ S15578 })
);
AOI22_X1 #() 
AOI22_X1_254_ (
  .A1({ S15553 }),
  .A2({ S25957[272] }),
  .B1({ S10988 }),
  .B2({ S10985 }),
  .ZN({ S15579 })
);
AOI21_X1 #() 
AOI21_X1_1141_ (
  .A({ S13772 }),
  .B1({ S15579 }),
  .B2({ S15551 }),
  .ZN({ S15581 })
);
AOI211_X1 #() 
AOI211_X1_27_ (
  .A({ S25957[277] }),
  .B({ S15575 }),
  .C1({ S15578 }),
  .C2({ S15581 }),
  .ZN({ S15582 })
);
AOI21_X1 #() 
AOI21_X1_1142_ (
  .A({ S15582 }),
  .B1({ S15566 }),
  .B2({ S25957[277] }),
  .ZN({ S15583 })
);
OAI21_X1 #() 
OAI21_X1_1061_ (
  .A({ S15560 }),
  .B1({ S15583 }),
  .B2({ S25957[278] }),
  .ZN({ S15584 })
);
INV_X1 #() 
INV_X1_615_ (
  .A({ S25957[278] }),
  .ZN({ S15585 })
);
AOI21_X1 #() 
AOI21_X1_1143_ (
  .A({ S25957[275] }),
  .B1({ S15515 }),
  .B2({ S25957[274] }),
  .ZN({ S15586 })
);
NAND2_X1 #() 
NAND2_X1_1921_ (
  .A1({ S15518 }),
  .A2({ S15553 }),
  .ZN({ S15587 })
);
NAND2_X1 #() 
NAND2_X1_1922_ (
  .A1({ S15587 }),
  .A2({ S15541 }),
  .ZN({ S15588 })
);
OAI21_X1 #() 
OAI21_X1_1062_ (
  .A({ S13772 }),
  .B1({ S15588 }),
  .B2({ S32 }),
  .ZN({ S15589 })
);
NOR2_X1 #() 
NOR2_X1_450_ (
  .A1({ S15529 }),
  .A2({ S32 }),
  .ZN({ S15590 })
);
AOI21_X1 #() 
AOI21_X1_1144_ (
  .A({ S25957[272] }),
  .B1({ S25957[274] }),
  .B2({ S15527 }),
  .ZN({ S15592 })
);
OAI21_X1 #() 
OAI21_X1_1063_ (
  .A({ S25957[276] }),
  .B1({ S15592 }),
  .B2({ S25957[275] }),
  .ZN({ S15593 })
);
OAI22_X1 #() 
OAI22_X1_49_ (
  .A1({ S15589 }),
  .A2({ S15586 }),
  .B1({ S15590 }),
  .B2({ S15593 }),
  .ZN({ S15594 })
);
AOI21_X1 #() 
AOI21_X1_1145_ (
  .A({ S25957[275] }),
  .B1({ S15577 }),
  .B2({ S15533 }),
  .ZN({ S15595 })
);
NAND2_X1 #() 
NAND2_X1_1923_ (
  .A1({ S15515 }),
  .A2({ S25957[274] }),
  .ZN({ S15596 })
);
NAND3_X1 #() 
NAND3_X1_2222_ (
  .A1({ S15518 }),
  .A2({ S15539 }),
  .A3({ S15553 }),
  .ZN({ S15597 })
);
AOI21_X1 #() 
AOI21_X1_1146_ (
  .A({ S32 }),
  .B1({ S15597 }),
  .B2({ S15596 }),
  .ZN({ S15598 })
);
OR3_X1 #() 
OR3_X1_8_ (
  .A1({ S15598 }),
  .A2({ S15595 }),
  .A3({ S13772 }),
  .ZN({ S15599 })
);
NAND4_X1 #() 
NAND4_X1_278_ (
  .A1({ S11278 }),
  .A2({ S15513 }),
  .A3({ S15514 }),
  .A4({ S11284 }),
  .ZN({ S15600 })
);
AOI22_X1 #() 
AOI22_X1_255_ (
  .A1({ S25957[274] }),
  .A2({ S25957[272] }),
  .B1({ S10991 }),
  .B2({ S10989 }),
  .ZN({ S15601 })
);
NAND2_X1 #() 
NAND2_X1_1924_ (
  .A1({ S15601 }),
  .A2({ S15600 }),
  .ZN({ S15603 })
);
NAND3_X1 #() 
NAND3_X1_2223_ (
  .A1({ S15600 }),
  .A2({ S15541 }),
  .A3({ S25957[272] }),
  .ZN({ S15604 })
);
AOI21_X1 #() 
AOI21_X1_1147_ (
  .A({ S25957[276] }),
  .B1({ S15604 }),
  .B2({ S32 }),
  .ZN({ S15605 })
);
AOI21_X1 #() 
AOI21_X1_1148_ (
  .A({ S25957[277] }),
  .B1({ S15605 }),
  .B2({ S15603 }),
  .ZN({ S15606 })
);
AOI22_X1 #() 
AOI22_X1_256_ (
  .A1({ S15594 }),
  .A2({ S25957[277] }),
  .B1({ S15599 }),
  .B2({ S15606 }),
  .ZN({ S15607 })
);
NAND2_X1 #() 
NAND2_X1_1925_ (
  .A1({ S32 }),
  .A2({ S25957[272] }),
  .ZN({ S15608 })
);
NAND2_X1 #() 
NAND2_X1_1926_ (
  .A1({ S15601 }),
  .A2({ S15567 }),
  .ZN({ S15609 })
);
NAND3_X1 #() 
NAND3_X1_2224_ (
  .A1({ S15609 }),
  .A2({ S25957[276] }),
  .A3({ S15608 }),
  .ZN({ S15610 })
);
NAND2_X1 #() 
NAND2_X1_1927_ (
  .A1({ S15515 }),
  .A2({ S15553 }),
  .ZN({ S15611 })
);
NAND2_X1 #() 
NAND2_X1_1928_ (
  .A1({ S15551 }),
  .A2({ S32 }),
  .ZN({ S15612 })
);
INV_X1 #() 
INV_X1_616_ (
  .A({ S15612 }),
  .ZN({ S15614 })
);
NAND3_X1 #() 
NAND3_X1_2225_ (
  .A1({ S15600 }),
  .A2({ S15518 }),
  .A3({ S25957[275] }),
  .ZN({ S15615 })
);
INV_X1 #() 
INV_X1_617_ (
  .A({ S15615 }),
  .ZN({ S15616 })
);
AOI21_X1 #() 
AOI21_X1_1149_ (
  .A({ S15616 }),
  .B1({ S15614 }),
  .B2({ S15611 }),
  .ZN({ S15617 })
);
OAI211_X1 #() 
OAI211_X1_712_ (
  .A({ S25957[277] }),
  .B({ S15610 }),
  .C1({ S15617 }),
  .C2({ S25957[276] }),
  .ZN({ S15618 })
);
NAND3_X1 #() 
NAND3_X1_2226_ (
  .A1({ S10804 }),
  .A2({ S10805 }),
  .A3({ S10807 }),
  .ZN({ S15619 })
);
NAND3_X1 #() 
NAND3_X1_2227_ (
  .A1({ S10808 }),
  .A2({ S10809 }),
  .A3({ S25957[405] }),
  .ZN({ S15620 })
);
NAND2_X1 #() 
NAND2_X1_1929_ (
  .A1({ S15619 }),
  .A2({ S15620 }),
  .ZN({ S15621 })
);
AOI21_X1 #() 
AOI21_X1_1150_ (
  .A({ S15553 }),
  .B1({ S15518 }),
  .B2({ S15539 }),
  .ZN({ S15622 })
);
NAND2_X1 #() 
NAND2_X1_1930_ (
  .A1({ S15526 }),
  .A2({ S32 }),
  .ZN({ S15623 })
);
NOR2_X1 #() 
NOR2_X1_451_ (
  .A1({ S15623 }),
  .A2({ S15622 }),
  .ZN({ S15625 })
);
NOR2_X1 #() 
NOR2_X1_452_ (
  .A1({ S15539 }),
  .A2({ S15553 }),
  .ZN({ S15626 })
);
OAI21_X1 #() 
OAI21_X1_1064_ (
  .A({ S25957[276] }),
  .B1({ S15626 }),
  .B2({ S32 }),
  .ZN({ S15627 })
);
NOR2_X1 #() 
NOR2_X1_453_ (
  .A1({ S15577 }),
  .A2({ S25957[275] }),
  .ZN({ S15628 })
);
OAI21_X1 #() 
OAI21_X1_1065_ (
  .A({ S13772 }),
  .B1({ S15596 }),
  .B2({ S32 }),
  .ZN({ S15629 })
);
OAI221_X1 #() 
OAI221_X1_42_ (
  .A({ S15621 }),
  .B1({ S15628 }),
  .B2({ S15629 }),
  .C1({ S15625 }),
  .C2({ S15627 }),
  .ZN({ S15630 })
);
NAND3_X1 #() 
NAND3_X1_2228_ (
  .A1({ S15630 }),
  .A2({ S15585 }),
  .A3({ S15618 }),
  .ZN({ S15631 })
);
OAI211_X1 #() 
OAI211_X1_713_ (
  .A({ S15517 }),
  .B({ S15631 }),
  .C1({ S15607 }),
  .C2({ S15585 }),
  .ZN({ S15632 })
);
OAI21_X1 #() 
OAI21_X1_1066_ (
  .A({ S15632 }),
  .B1({ S15584 }),
  .B2({ S15517 }),
  .ZN({ S15633 })
);
NOR2_X1 #() 
NOR2_X1_454_ (
  .A1({ S15633 }),
  .A2({ S9904 }),
  .ZN({ S15634 })
);
INV_X1 #() 
INV_X1_618_ (
  .A({ S15634 }),
  .ZN({ S15636 })
);
NAND2_X1 #() 
NAND2_X1_1931_ (
  .A1({ S15633 }),
  .A2({ S9904 }),
  .ZN({ S15637 })
);
NAND3_X1 #() 
NAND3_X1_2229_ (
  .A1({ S15636 }),
  .A2({ S9910 }),
  .A3({ S15637 }),
  .ZN({ S15638 })
);
NAND2_X1 #() 
NAND2_X1_1932_ (
  .A1({ S15636 }),
  .A2({ S15637 }),
  .ZN({ S25957[223] })
);
NAND2_X1 #() 
NAND2_X1_1933_ (
  .A1({ S25957[223] }),
  .A2({ S25957[415] }),
  .ZN({ S15639 })
);
NAND2_X1 #() 
NAND2_X1_1934_ (
  .A1({ S15639 }),
  .A2({ S15638 }),
  .ZN({ S15640 })
);
INV_X1 #() 
INV_X1_619_ (
  .A({ S15640 }),
  .ZN({ S25957[159] })
);
NAND2_X1 #() 
NAND2_X1_1935_ (
  .A1({ S9997 }),
  .A2({ S10003 }),
  .ZN({ S15641 })
);
INV_X1 #() 
INV_X1_620_ (
  .A({ S15641 }),
  .ZN({ S25957[446] })
);
NAND3_X1 #() 
NAND3_X1_2230_ (
  .A1({ S15567 }),
  .A2({ S32 }),
  .A3({ S15519 }),
  .ZN({ S15642 })
);
INV_X1 #() 
INV_X1_621_ (
  .A({ S15600 }),
  .ZN({ S15644 })
);
NAND2_X1 #() 
NAND2_X1_1936_ (
  .A1({ S15644 }),
  .A2({ S25957[275] }),
  .ZN({ S15645 })
);
NAND3_X1 #() 
NAND3_X1_2231_ (
  .A1({ S15645 }),
  .A2({ S25957[276] }),
  .A3({ S15642 }),
  .ZN({ S15646 })
);
NAND3_X1 #() 
NAND3_X1_2232_ (
  .A1({ S15515 }),
  .A2({ S53 }),
  .A3({ S25957[274] }),
  .ZN({ S15647 })
);
NAND2_X1 #() 
NAND2_X1_1937_ (
  .A1({ S15647 }),
  .A2({ S32 }),
  .ZN({ S15648 })
);
NAND3_X1 #() 
NAND3_X1_2233_ (
  .A1({ S25957[274] }),
  .A2({ S15527 }),
  .A3({ S25957[272] }),
  .ZN({ S15649 })
);
NAND3_X1 #() 
NAND3_X1_2234_ (
  .A1({ S15649 }),
  .A2({ S25957[275] }),
  .A3({ S15533 }),
  .ZN({ S15650 })
);
NAND3_X1 #() 
NAND3_X1_2235_ (
  .A1({ S15648 }),
  .A2({ S13772 }),
  .A3({ S15650 }),
  .ZN({ S15651 })
);
NAND2_X1 #() 
NAND2_X1_1938_ (
  .A1({ S15651 }),
  .A2({ S15646 }),
  .ZN({ S15652 })
);
NAND4_X1 #() 
NAND4_X1_279_ (
  .A1({ S11278 }),
  .A2({ S11284 }),
  .A3({ S15511 }),
  .A4({ S15512 }),
  .ZN({ S15653 })
);
NAND2_X1 #() 
NAND2_X1_1939_ (
  .A1({ S15653 }),
  .A2({ S53 }),
  .ZN({ S15655 })
);
OAI21_X1 #() 
OAI21_X1_1067_ (
  .A({ S25957[276] }),
  .B1({ S15655 }),
  .B2({ S32 }),
  .ZN({ S15656 })
);
AOI21_X1 #() 
AOI21_X1_1151_ (
  .A({ S15656 }),
  .B1({ S15579 }),
  .B2({ S15596 }),
  .ZN({ S15657 })
);
NAND2_X1 #() 
NAND2_X1_1940_ (
  .A1({ S15653 }),
  .A2({ S25957[273] }),
  .ZN({ S15658 })
);
OAI21_X1 #() 
OAI21_X1_1068_ (
  .A({ S15658 }),
  .B1({ S32 }),
  .B2({ S15549 }),
  .ZN({ S15659 })
);
AOI21_X1 #() 
AOI21_X1_1152_ (
  .A({ S15657 }),
  .B1({ S13772 }),
  .B2({ S15659 }),
  .ZN({ S15660 })
);
MUX2_X1 #() 
MUX2_X1_6_ (
  .A({ S15652 }),
  .B({ S15660 }),
  .S({ S25957[277] }),
  .Z({ S15661 })
);
AOI22_X1 #() 
AOI22_X1_257_ (
  .A1({ S25957[273] }),
  .A2({ S15519 }),
  .B1({ S15522 }),
  .B2({ S15523 }),
  .ZN({ S15662 })
);
OAI21_X1 #() 
OAI21_X1_1069_ (
  .A({ S25957[275] }),
  .B1({ S15626 }),
  .B2({ S15662 }),
  .ZN({ S15663 })
);
NAND2_X1 #() 
NAND2_X1_1941_ (
  .A1({ S15663 }),
  .A2({ S13772 }),
  .ZN({ S15664 })
);
NAND2_X1 #() 
NAND2_X1_1942_ (
  .A1({ S15568 }),
  .A2({ S32 }),
  .ZN({ S15666 })
);
NAND2_X1 #() 
NAND2_X1_1943_ (
  .A1({ S15588 }),
  .A2({ S25957[275] }),
  .ZN({ S15667 })
);
OAI21_X1 #() 
OAI21_X1_1070_ (
  .A({ S15667 }),
  .B1({ S15519 }),
  .B2({ S15666 }),
  .ZN({ S15668 })
);
OAI21_X1 #() 
OAI21_X1_1071_ (
  .A({ S15664 }),
  .B1({ S15668 }),
  .B2({ S13772 }),
  .ZN({ S15669 })
);
NOR2_X1 #() 
NOR2_X1_455_ (
  .A1({ S15518 }),
  .A2({ S25957[274] }),
  .ZN({ S15670 })
);
NAND2_X1 #() 
NAND2_X1_1944_ (
  .A1({ S15541 }),
  .A2({ S25957[275] }),
  .ZN({ S15671 })
);
OAI221_X1 #() 
OAI221_X1_43_ (
  .A({ S13772 }),
  .B1({ S15671 }),
  .B2({ S15644 }),
  .C1({ S15612 }),
  .C2({ S15670 }),
  .ZN({ S15672 })
);
NAND2_X1 #() 
NAND2_X1_1945_ (
  .A1({ S15653 }),
  .A2({ S32 }),
  .ZN({ S15673 })
);
OAI21_X1 #() 
OAI21_X1_1072_ (
  .A({ S15515 }),
  .B1({ S53 }),
  .B2({ S15553 }),
  .ZN({ S15674 })
);
OAI211_X1 #() 
OAI211_X1_714_ (
  .A({ S25957[276] }),
  .B({ S15673 }),
  .C1({ S15674 }),
  .C2({ S32 }),
  .ZN({ S15675 })
);
NAND3_X1 #() 
NAND3_X1_2236_ (
  .A1({ S15672 }),
  .A2({ S25957[277] }),
  .A3({ S15675 }),
  .ZN({ S15677 })
);
OAI21_X1 #() 
OAI21_X1_1073_ (
  .A({ S15677 }),
  .B1({ S15669 }),
  .B2({ S25957[277] }),
  .ZN({ S15678 })
);
NAND2_X1 #() 
NAND2_X1_1946_ (
  .A1({ S15678 }),
  .A2({ S15585 }),
  .ZN({ S15679 })
);
OAI21_X1 #() 
OAI21_X1_1074_ (
  .A({ S15679 }),
  .B1({ S15661 }),
  .B2({ S15585 }),
  .ZN({ S15680 })
);
NOR2_X1 #() 
NOR2_X1_456_ (
  .A1({ S15542 }),
  .A2({ S15524 }),
  .ZN({ S15681 })
);
NAND2_X1 #() 
NAND2_X1_1947_ (
  .A1({ S15681 }),
  .A2({ S15531 }),
  .ZN({ S15682 })
);
NAND3_X1 #() 
NAND3_X1_2237_ (
  .A1({ S53 }),
  .A2({ S32 }),
  .A3({ S25957[274] }),
  .ZN({ S15683 })
);
AND2_X1 #() 
AND2_X1_119_ (
  .A1({ S15682 }),
  .A2({ S15683 }),
  .ZN({ S15684 })
);
NAND2_X1 #() 
NAND2_X1_1948_ (
  .A1({ S15684 }),
  .A2({ S25957[276] }),
  .ZN({ S15685 })
);
INV_X1 #() 
INV_X1_622_ (
  .A({ S15545 }),
  .ZN({ S15686 })
);
OAI21_X1 #() 
OAI21_X1_1075_ (
  .A({ S13772 }),
  .B1({ S15686 }),
  .B2({ S15561 }),
  .ZN({ S15688 })
);
AOI21_X1 #() 
AOI21_X1_1153_ (
  .A({ S15621 }),
  .B1({ S15685 }),
  .B2({ S15688 }),
  .ZN({ S15689 })
);
INV_X1 #() 
INV_X1_623_ (
  .A({ S15650 }),
  .ZN({ S15690 })
);
AOI21_X1 #() 
AOI21_X1_1154_ (
  .A({ S25957[275] }),
  .B1({ S15576 }),
  .B2({ S15549 }),
  .ZN({ S15691 })
);
OAI21_X1 #() 
OAI21_X1_1076_ (
  .A({ S25957[276] }),
  .B1({ S15690 }),
  .B2({ S15691 }),
  .ZN({ S15692 })
);
NAND4_X1 #() 
NAND4_X1_280_ (
  .A1({ S15600 }),
  .A2({ S15541 }),
  .A3({ S32 }),
  .A4({ S25957[272] }),
  .ZN({ S15693 })
);
AOI21_X1 #() 
AOI21_X1_1155_ (
  .A({ S32 }),
  .B1({ S15533 }),
  .B2({ S25957[273] }),
  .ZN({ S15694 })
);
INV_X1 #() 
INV_X1_624_ (
  .A({ S15694 }),
  .ZN({ S15695 })
);
OAI211_X1 #() 
OAI211_X1_715_ (
  .A({ S13772 }),
  .B({ S15693 }),
  .C1({ S15695 }),
  .C2({ S15550 }),
  .ZN({ S15696 })
);
AOI21_X1 #() 
AOI21_X1_1156_ (
  .A({ S25957[277] }),
  .B1({ S15692 }),
  .B2({ S15696 }),
  .ZN({ S15697 })
);
OAI21_X1 #() 
OAI21_X1_1077_ (
  .A({ S25957[278] }),
  .B1({ S15689 }),
  .B2({ S15697 }),
  .ZN({ S15699 })
);
NAND3_X1 #() 
NAND3_X1_2238_ (
  .A1({ S25957[275] }),
  .A2({ S25957[273] }),
  .A3({ S25957[274] }),
  .ZN({ S15700 })
);
OAI21_X1 #() 
OAI21_X1_1078_ (
  .A({ S15700 }),
  .B1({ S15562 }),
  .B2({ S15533 }),
  .ZN({ S15701 })
);
OAI21_X1 #() 
OAI21_X1_1079_ (
  .A({ S25957[276] }),
  .B1({ S15701 }),
  .B2({ S15628 }),
  .ZN({ S15702 })
);
AOI22_X1 #() 
AOI22_X1_258_ (
  .A1({ S15522 }),
  .A2({ S15523 }),
  .B1({ S15512 }),
  .B2({ S15511 }),
  .ZN({ S15703 })
);
NAND2_X1 #() 
NAND2_X1_1949_ (
  .A1({ S15703 }),
  .A2({ S25957[273] }),
  .ZN({ S15704 })
);
INV_X1 #() 
INV_X1_625_ (
  .A({ S15704 }),
  .ZN({ S15705 })
);
NAND3_X1 #() 
NAND3_X1_2239_ (
  .A1({ S25957[274] }),
  .A2({ S25957[273] }),
  .A3({ S25957[272] }),
  .ZN({ S15706 })
);
NAND2_X1 #() 
NAND2_X1_1950_ (
  .A1({ S15706 }),
  .A2({ S53 }),
  .ZN({ S15707 })
);
AOI21_X1 #() 
AOI21_X1_1157_ (
  .A({ S25957[276] }),
  .B1({ S15707 }),
  .B2({ S32 }),
  .ZN({ S15708 })
);
OAI21_X1 #() 
OAI21_X1_1080_ (
  .A({ S15708 }),
  .B1({ S15671 }),
  .B2({ S15705 }),
  .ZN({ S15710 })
);
NAND3_X1 #() 
NAND3_X1_2240_ (
  .A1({ S15710 }),
  .A2({ S25957[277] }),
  .A3({ S15702 }),
  .ZN({ S15711 })
);
OAI21_X1 #() 
OAI21_X1_1081_ (
  .A({ S15653 }),
  .B1({ S15539 }),
  .B2({ S15553 }),
  .ZN({ S15712 })
);
AOI21_X1 #() 
AOI21_X1_1158_ (
  .A({ S15691 }),
  .B1({ S25957[275] }),
  .B2({ S15712 }),
  .ZN({ S15713 })
);
NOR2_X1 #() 
NOR2_X1_457_ (
  .A1({ S15587 }),
  .A2({ S25957[275] }),
  .ZN({ S15714 })
);
NAND2_X1 #() 
NAND2_X1_1951_ (
  .A1({ S15563 }),
  .A2({ S25957[276] }),
  .ZN({ S15715 })
);
OAI22_X1 #() 
OAI22_X1_50_ (
  .A1({ S15713 }),
  .A2({ S25957[276] }),
  .B1({ S15714 }),
  .B2({ S15715 }),
  .ZN({ S15716 })
);
OAI211_X1 #() 
OAI211_X1_716_ (
  .A({ S15585 }),
  .B({ S15711 }),
  .C1({ S15716 }),
  .C2({ S25957[277] }),
  .ZN({ S15717 })
);
NAND3_X1 #() 
NAND3_X1_2241_ (
  .A1({ S15717 }),
  .A2({ S25957[279] }),
  .A3({ S15699 }),
  .ZN({ S15718 })
);
OAI21_X1 #() 
OAI21_X1_1082_ (
  .A({ S15718 }),
  .B1({ S15680 }),
  .B2({ S25957[279] }),
  .ZN({ S15719 })
);
NAND2_X1 #() 
NAND2_X1_1952_ (
  .A1({ S15719 }),
  .A2({ S12880 }),
  .ZN({ S15721 })
);
OR2_X1 #() 
OR2_X1_28_ (
  .A1({ S15719 }),
  .A2({ S12880 }),
  .ZN({ S15722 })
);
NAND2_X1 #() 
NAND2_X1_1953_ (
  .A1({ S15722 }),
  .A2({ S15721 }),
  .ZN({ S25957[254] })
);
NAND2_X1 #() 
NAND2_X1_1954_ (
  .A1({ S25957[254] }),
  .A2({ S25957[446] }),
  .ZN({ S15723 })
);
INV_X1 #() 
INV_X1_626_ (
  .A({ S15723 }),
  .ZN({ S15724 })
);
NOR2_X1 #() 
NOR2_X1_458_ (
  .A1({ S25957[254] }),
  .A2({ S25957[446] }),
  .ZN({ S15725 })
);
OAI21_X1 #() 
OAI21_X1_1083_ (
  .A({ S14823 }),
  .B1({ S15724 }),
  .B2({ S15725 }),
  .ZN({ S15726 })
);
INV_X1 #() 
INV_X1_627_ (
  .A({ S15725 }),
  .ZN({ S15727 })
);
NAND3_X1 #() 
NAND3_X1_2242_ (
  .A1({ S15727 }),
  .A2({ S25957[286] }),
  .A3({ S15723 }),
  .ZN({ S15728 })
);
NAND2_X1 #() 
NAND2_X1_1955_ (
  .A1({ S15726 }),
  .A2({ S15728 }),
  .ZN({ S15729 })
);
INV_X1 #() 
INV_X1_628_ (
  .A({ S15729 }),
  .ZN({ S25957[158] })
);
NAND2_X1 #() 
NAND2_X1_1956_ (
  .A1({ S10086 }),
  .A2({ S10085 }),
  .ZN({ S25957[477] })
);
NAND2_X1 #() 
NAND2_X1_1957_ (
  .A1({ S12963 }),
  .A2({ S12958 }),
  .ZN({ S15731 })
);
XNOR2_X1 #() 
XNOR2_X1_64_ (
  .A({ S15731 }),
  .B({ S25957[477] }),
  .ZN({ S25957[349] })
);
INV_X1 #() 
INV_X1_629_ (
  .A({ S15731 }),
  .ZN({ S25957[381] })
);
AOI22_X1 #() 
AOI22_X1_259_ (
  .A1({ S11278 }),
  .A2({ S11284 }),
  .B1({ S15512 }),
  .B2({ S15511 }),
  .ZN({ S15732 })
);
NAND2_X1 #() 
NAND2_X1_1958_ (
  .A1({ S15561 }),
  .A2({ S15732 }),
  .ZN({ S15733 })
);
NAND2_X1 #() 
NAND2_X1_1959_ (
  .A1({ S15567 }),
  .A2({ S15519 }),
  .ZN({ S15734 })
);
AOI21_X1 #() 
AOI21_X1_1159_ (
  .A({ S15714 }),
  .B1({ S15734 }),
  .B2({ S25957[275] }),
  .ZN({ S15735 })
);
AOI21_X1 #() 
AOI21_X1_1160_ (
  .A({ S13772 }),
  .B1({ S15735 }),
  .B2({ S15733 }),
  .ZN({ S15736 })
);
AND2_X1 #() 
AND2_X1_120_ (
  .A1({ S53 }),
  .A2({ S32 }),
  .ZN({ S15738 })
);
NAND2_X1 #() 
NAND2_X1_1960_ (
  .A1({ S15738 }),
  .A2({ S15567 }),
  .ZN({ S15739 })
);
NAND2_X1 #() 
NAND2_X1_1961_ (
  .A1({ S15539 }),
  .A2({ S25957[274] }),
  .ZN({ S15740 })
);
NAND2_X1 #() 
NAND2_X1_1962_ (
  .A1({ S15611 }),
  .A2({ S15740 }),
  .ZN({ S15741 })
);
NAND2_X1 #() 
NAND2_X1_1963_ (
  .A1({ S15741 }),
  .A2({ S25957[275] }),
  .ZN({ S15742 })
);
AOI21_X1 #() 
AOI21_X1_1161_ (
  .A({ S25957[276] }),
  .B1({ S15742 }),
  .B2({ S15739 }),
  .ZN({ S15743 })
);
OAI21_X1 #() 
OAI21_X1_1084_ (
  .A({ S25957[277] }),
  .B1({ S15736 }),
  .B2({ S15743 }),
  .ZN({ S15744 })
);
INV_X1 #() 
INV_X1_630_ (
  .A({ S15628 }),
  .ZN({ S15745 })
);
AOI21_X1 #() 
AOI21_X1_1162_ (
  .A({ S25957[276] }),
  .B1({ S15745 }),
  .B2({ S15650 }),
  .ZN({ S15746 })
);
NAND3_X1 #() 
NAND3_X1_2243_ (
  .A1({ S15567 }),
  .A2({ S15653 }),
  .A3({ S25957[275] }),
  .ZN({ S15747 })
);
INV_X1 #() 
INV_X1_631_ (
  .A({ S15740 }),
  .ZN({ S15749 })
);
NAND2_X1 #() 
NAND2_X1_1964_ (
  .A1({ S15749 }),
  .A2({ S32 }),
  .ZN({ S15750 })
);
AOI21_X1 #() 
AOI21_X1_1163_ (
  .A({ S13772 }),
  .B1({ S15750 }),
  .B2({ S15747 }),
  .ZN({ S15751 })
);
OAI21_X1 #() 
OAI21_X1_1085_ (
  .A({ S15621 }),
  .B1({ S15746 }),
  .B2({ S15751 }),
  .ZN({ S15752 })
);
AOI21_X1 #() 
AOI21_X1_1164_ (
  .A({ S15585 }),
  .B1({ S15744 }),
  .B2({ S15752 }),
  .ZN({ S15753 })
);
NAND2_X1 #() 
NAND2_X1_1965_ (
  .A1({ S15541 }),
  .A2({ S15515 }),
  .ZN({ S15754 })
);
INV_X1 #() 
INV_X1_632_ (
  .A({ S15542 }),
  .ZN({ S15755 })
);
AOI21_X1 #() 
AOI21_X1_1165_ (
  .A({ S15755 }),
  .B1({ S15754 }),
  .B2({ S32 }),
  .ZN({ S15756 })
);
NAND3_X1 #() 
NAND3_X1_2244_ (
  .A1({ S15533 }),
  .A2({ S15515 }),
  .A3({ S32 }),
  .ZN({ S15757 })
);
OAI21_X1 #() 
OAI21_X1_1086_ (
  .A({ S15757 }),
  .B1({ S15604 }),
  .B2({ S32 }),
  .ZN({ S15758 })
);
NAND2_X1 #() 
NAND2_X1_1966_ (
  .A1({ S15758 }),
  .A2({ S25957[276] }),
  .ZN({ S15760 })
);
OAI21_X1 #() 
OAI21_X1_1087_ (
  .A({ S15760 }),
  .B1({ S25957[276] }),
  .B2({ S15756 }),
  .ZN({ S15761 })
);
NOR2_X1 #() 
NOR2_X1_459_ (
  .A1({ S53 }),
  .A2({ S25957[274] }),
  .ZN({ S15762 })
);
OAI21_X1 #() 
OAI21_X1_1088_ (
  .A({ S25957[275] }),
  .B1({ S15622 }),
  .B2({ S15762 }),
  .ZN({ S15763 })
);
NAND3_X1 #() 
NAND3_X1_2245_ (
  .A1({ S15763 }),
  .A2({ S13772 }),
  .A3({ S15623 }),
  .ZN({ S15764 })
);
NAND2_X1 #() 
NAND2_X1_1967_ (
  .A1({ S15570 }),
  .A2({ S25957[275] }),
  .ZN({ S15765 })
);
NAND2_X1 #() 
NAND2_X1_1968_ (
  .A1({ S15579 }),
  .A2({ S15527 }),
  .ZN({ S15766 })
);
NAND2_X1 #() 
NAND2_X1_1969_ (
  .A1({ S15765 }),
  .A2({ S15766 }),
  .ZN({ S15767 })
);
AOI21_X1 #() 
AOI21_X1_1166_ (
  .A({ S25957[277] }),
  .B1({ S15767 }),
  .B2({ S25957[276] }),
  .ZN({ S15768 })
);
AOI22_X1 #() 
AOI22_X1_260_ (
  .A1({ S15764 }),
  .A2({ S15768 }),
  .B1({ S15761 }),
  .B2({ S25957[277] }),
  .ZN({ S15769 })
);
NOR2_X1 #() 
NOR2_X1_460_ (
  .A1({ S15769 }),
  .A2({ S25957[278] }),
  .ZN({ S15771 })
);
OAI21_X1 #() 
OAI21_X1_1089_ (
  .A({ S25957[279] }),
  .B1({ S15771 }),
  .B2({ S15753 }),
  .ZN({ S15772 })
);
NAND3_X1 #() 
NAND3_X1_2246_ (
  .A1({ S15611 }),
  .A2({ S15706 }),
  .A3({ S32 }),
  .ZN({ S15773 })
);
NAND3_X1 #() 
NAND3_X1_2247_ (
  .A1({ S15518 }),
  .A2({ S25957[275] }),
  .A3({ S15553 }),
  .ZN({ S15774 })
);
NAND3_X1 #() 
NAND3_X1_2248_ (
  .A1({ S15773 }),
  .A2({ S25957[276] }),
  .A3({ S15774 }),
  .ZN({ S15775 })
);
NAND4_X1 #() 
NAND4_X1_281_ (
  .A1({ S15541 }),
  .A2({ S15653 }),
  .A3({ S15531 }),
  .A4({ S25957[275] }),
  .ZN({ S15776 })
);
INV_X1 #() 
INV_X1_633_ (
  .A({ S15776 }),
  .ZN({ S15777 })
);
NAND2_X1 #() 
NAND2_X1_1970_ (
  .A1({ S15539 }),
  .A2({ S15553 }),
  .ZN({ S15778 })
);
AOI21_X1 #() 
AOI21_X1_1167_ (
  .A({ S25957[275] }),
  .B1({ S15778 }),
  .B2({ S15531 }),
  .ZN({ S15779 })
);
OAI21_X1 #() 
OAI21_X1_1090_ (
  .A({ S13772 }),
  .B1({ S15779 }),
  .B2({ S15777 }),
  .ZN({ S15780 })
);
AND3_X1 #() 
AND3_X1_89_ (
  .A1({ S15780 }),
  .A2({ S15775 }),
  .A3({ S25957[278] }),
  .ZN({ S15782 })
);
NAND2_X1 #() 
NAND2_X1_1971_ (
  .A1({ S15520 }),
  .A2({ S15567 }),
  .ZN({ S15783 })
);
NAND3_X1 #() 
NAND3_X1_2249_ (
  .A1({ S15553 }),
  .A2({ S15527 }),
  .A3({ S25957[272] }),
  .ZN({ S15784 })
);
NAND3_X1 #() 
NAND3_X1_2250_ (
  .A1({ S15577 }),
  .A2({ S25957[275] }),
  .A3({ S15784 }),
  .ZN({ S15785 })
);
NAND3_X1 #() 
NAND3_X1_2251_ (
  .A1({ S15649 }),
  .A2({ S32 }),
  .A3({ S15533 }),
  .ZN({ S15786 })
);
OAI211_X1 #() 
OAI211_X1_717_ (
  .A({ S15785 }),
  .B({ S25957[276] }),
  .C1({ S15783 }),
  .C2({ S15786 }),
  .ZN({ S15787 })
);
AOI21_X1 #() 
AOI21_X1_1168_ (
  .A({ S25957[276] }),
  .B1({ S15551 }),
  .B2({ S32 }),
  .ZN({ S15788 })
);
OAI211_X1 #() 
OAI211_X1_718_ (
  .A({ S15788 }),
  .B({ S25957[272] }),
  .C1({ S15527 }),
  .C2({ S32 }),
  .ZN({ S15789 })
);
AND3_X1 #() 
AND3_X1_90_ (
  .A1({ S15787 }),
  .A2({ S15585 }),
  .A3({ S15789 }),
  .ZN({ S15790 })
);
OAI21_X1 #() 
OAI21_X1_1091_ (
  .A({ S15621 }),
  .B1({ S15782 }),
  .B2({ S15790 }),
  .ZN({ S15791 })
);
AOI22_X1 #() 
AOI22_X1_261_ (
  .A1({ S15541 }),
  .A2({ S15549 }),
  .B1({ S15527 }),
  .B2({ S25957[272] }),
  .ZN({ S15793 })
);
NAND3_X1 #() 
NAND3_X1_2252_ (
  .A1({ S15587 }),
  .A2({ S32 }),
  .A3({ S15541 }),
  .ZN({ S15794 })
);
OAI21_X1 #() 
OAI21_X1_1092_ (
  .A({ S25957[275] }),
  .B1({ S15539 }),
  .B2({ S25957[274] }),
  .ZN({ S15795 })
);
OAI211_X1 #() 
OAI211_X1_719_ (
  .A({ S15794 }),
  .B({ S25957[276] }),
  .C1({ S15793 }),
  .C2({ S15795 }),
  .ZN({ S15796 })
);
NOR2_X1 #() 
NOR2_X1_461_ (
  .A1({ S32 }),
  .A2({ S25957[272] }),
  .ZN({ S15797 })
);
AOI21_X1 #() 
AOI21_X1_1169_ (
  .A({ S25957[275] }),
  .B1({ S15549 }),
  .B2({ S53 }),
  .ZN({ S15798 })
);
OAI21_X1 #() 
OAI21_X1_1093_ (
  .A({ S13772 }),
  .B1({ S15798 }),
  .B2({ S15797 }),
  .ZN({ S15799 })
);
NAND3_X1 #() 
NAND3_X1_2253_ (
  .A1({ S15796 }),
  .A2({ S25957[278] }),
  .A3({ S15799 }),
  .ZN({ S15800 })
);
AOI21_X1 #() 
AOI21_X1_1170_ (
  .A({ S25957[275] }),
  .B1({ S15596 }),
  .B2({ S15778 }),
  .ZN({ S15801 })
);
OAI21_X1 #() 
OAI21_X1_1094_ (
  .A({ S32 }),
  .B1({ S15539 }),
  .B2({ S25957[274] }),
  .ZN({ S15802 })
);
OAI21_X1 #() 
OAI21_X1_1095_ (
  .A({ S15802 }),
  .B1({ S32 }),
  .B2({ S15611 }),
  .ZN({ S15804 })
);
NAND2_X1 #() 
NAND2_X1_1972_ (
  .A1({ S15804 }),
  .A2({ S25957[276] }),
  .ZN({ S15805 })
);
OAI21_X1 #() 
OAI21_X1_1096_ (
  .A({ S13772 }),
  .B1({ S15550 }),
  .B2({ S32 }),
  .ZN({ S15806 })
);
OAI21_X1 #() 
OAI21_X1_1097_ (
  .A({ S15805 }),
  .B1({ S15801 }),
  .B2({ S15806 }),
  .ZN({ S15807 })
);
OAI21_X1 #() 
OAI21_X1_1098_ (
  .A({ S15800 }),
  .B1({ S15807 }),
  .B2({ S25957[278] }),
  .ZN({ S15808 })
);
NAND2_X1 #() 
NAND2_X1_1973_ (
  .A1({ S15808 }),
  .A2({ S25957[277] }),
  .ZN({ S15809 })
);
NAND3_X1 #() 
NAND3_X1_2254_ (
  .A1({ S15791 }),
  .A2({ S15809 }),
  .A3({ S15517 }),
  .ZN({ S15810 })
);
NAND3_X1 #() 
NAND3_X1_2255_ (
  .A1({ S15772 }),
  .A2({ S15810 }),
  .A3({ S25957[381] }),
  .ZN({ S15811 })
);
NAND2_X1 #() 
NAND2_X1_1974_ (
  .A1({ S15791 }),
  .A2({ S15809 }),
  .ZN({ S15812 })
);
NAND2_X1 #() 
NAND2_X1_1975_ (
  .A1({ S15812 }),
  .A2({ S15517 }),
  .ZN({ S15813 })
);
OR3_X1 #() 
OR3_X1_9_ (
  .A1({ S15771 }),
  .A2({ S15753 }),
  .A3({ S15517 }),
  .ZN({ S15815 })
);
NAND3_X1 #() 
NAND3_X1_2256_ (
  .A1({ S15815 }),
  .A2({ S15813 }),
  .A3({ S15731 }),
  .ZN({ S15816 })
);
NAND3_X1 #() 
NAND3_X1_2257_ (
  .A1({ S15816 }),
  .A2({ S15811 }),
  .A3({ S25957[349] }),
  .ZN({ S15817 })
);
INV_X1 #() 
INV_X1_634_ (
  .A({ S25957[349] }),
  .ZN({ S15818 })
);
NAND3_X1 #() 
NAND3_X1_2258_ (
  .A1({ S15815 }),
  .A2({ S15813 }),
  .A3({ S25957[381] }),
  .ZN({ S15819 })
);
NAND3_X1 #() 
NAND3_X1_2259_ (
  .A1({ S15772 }),
  .A2({ S15810 }),
  .A3({ S15731 }),
  .ZN({ S15820 })
);
NAND3_X1 #() 
NAND3_X1_2260_ (
  .A1({ S15819 }),
  .A2({ S15820 }),
  .A3({ S15818 }),
  .ZN({ S15821 })
);
NAND3_X1 #() 
NAND3_X1_2261_ (
  .A1({ S15817 }),
  .A2({ S15821 }),
  .A3({ S12034 }),
  .ZN({ S15822 })
);
NAND3_X1 #() 
NAND3_X1_2262_ (
  .A1({ S15816 }),
  .A2({ S15811 }),
  .A3({ S15818 }),
  .ZN({ S15823 })
);
NAND3_X1 #() 
NAND3_X1_2263_ (
  .A1({ S15819 }),
  .A2({ S15820 }),
  .A3({ S25957[349] }),
  .ZN({ S15824 })
);
NAND3_X1 #() 
NAND3_X1_2264_ (
  .A1({ S15823 }),
  .A2({ S15824 }),
  .A3({ S25957[413] }),
  .ZN({ S15826 })
);
NAND2_X1 #() 
NAND2_X1_1976_ (
  .A1({ S15822 }),
  .A2({ S15826 }),
  .ZN({ S25957[157] })
);
NAND2_X1 #() 
NAND2_X1_1977_ (
  .A1({ S13074 }),
  .A2({ S13078 }),
  .ZN({ S25957[316] })
);
NAND2_X1 #() 
NAND2_X1_1978_ (
  .A1({ S13031 }),
  .A2({ S13073 }),
  .ZN({ S25957[380] })
);
AOI21_X1 #() 
AOI21_X1_1171_ (
  .A({ S25957[276] }),
  .B1({ S25957[275] }),
  .B2({ S25957[274] }),
  .ZN({ S15827 })
);
OAI21_X1 #() 
OAI21_X1_1099_ (
  .A({ S15827 }),
  .B1({ S15623 }),
  .B2({ S15732 }),
  .ZN({ S15828 })
);
NAND3_X1 #() 
NAND3_X1_2265_ (
  .A1({ S15551 }),
  .A2({ S32 }),
  .A3({ S15549 }),
  .ZN({ S15829 })
);
OAI211_X1 #() 
OAI211_X1_720_ (
  .A({ S15563 }),
  .B({ S25957[276] }),
  .C1({ S15568 }),
  .C2({ S15829 }),
  .ZN({ S15830 })
);
NAND2_X1 #() 
NAND2_X1_1979_ (
  .A1({ S15830 }),
  .A2({ S15828 }),
  .ZN({ S15831 })
);
AOI21_X1 #() 
AOI21_X1_1172_ (
  .A({ S13772 }),
  .B1({ S151 }),
  .B2({ S15553 }),
  .ZN({ S15832 })
);
OAI21_X1 #() 
OAI21_X1_1100_ (
  .A({ S32 }),
  .B1({ S15749 }),
  .B2({ S15570 }),
  .ZN({ S15834 })
);
NAND2_X1 #() 
NAND2_X1_1980_ (
  .A1({ S15706 }),
  .A2({ S15533 }),
  .ZN({ S15835 })
);
AOI21_X1 #() 
AOI21_X1_1173_ (
  .A({ S25957[276] }),
  .B1({ S15835 }),
  .B2({ S25957[275] }),
  .ZN({ S15836 })
);
AOI21_X1 #() 
AOI21_X1_1174_ (
  .A({ S15832 }),
  .B1({ S15836 }),
  .B2({ S15834 }),
  .ZN({ S15837 })
);
NAND2_X1 #() 
NAND2_X1_1981_ (
  .A1({ S15837 }),
  .A2({ S25957[277] }),
  .ZN({ S15838 })
);
OAI211_X1 #() 
OAI211_X1_721_ (
  .A({ S15838 }),
  .B({ S25957[278] }),
  .C1({ S25957[277] }),
  .C2({ S15831 }),
  .ZN({ S15839 })
);
AOI21_X1 #() 
AOI21_X1_1175_ (
  .A({ S32 }),
  .B1({ S15653 }),
  .B2({ S15539 }),
  .ZN({ S15840 })
);
NAND4_X1 #() 
NAND4_X1_282_ (
  .A1({ S32 }),
  .A2({ S15553 }),
  .A3({ S15519 }),
  .A4({ S15527 }),
  .ZN({ S15841 })
);
NAND2_X1 #() 
NAND2_X1_1982_ (
  .A1({ S15841 }),
  .A2({ S15683 }),
  .ZN({ S15842 })
);
OAI21_X1 #() 
OAI21_X1_1101_ (
  .A({ S13772 }),
  .B1({ S15842 }),
  .B2({ S15840 }),
  .ZN({ S15843 })
);
AOI21_X1 #() 
AOI21_X1_1176_ (
  .A({ S13772 }),
  .B1({ S15754 }),
  .B2({ S32 }),
  .ZN({ S15845 })
);
NAND3_X1 #() 
NAND3_X1_2266_ (
  .A1({ S15587 }),
  .A2({ S25957[275] }),
  .A3({ S15549 }),
  .ZN({ S15846 })
);
NAND2_X1 #() 
NAND2_X1_1983_ (
  .A1({ S15845 }),
  .A2({ S15846 }),
  .ZN({ S15847 })
);
AND2_X1 #() 
AND2_X1_121_ (
  .A1({ S15843 }),
  .A2({ S15847 }),
  .ZN({ S15848 })
);
NAND2_X1 #() 
NAND2_X1_1984_ (
  .A1({ S15740 }),
  .A2({ S32 }),
  .ZN({ S15849 })
);
NAND3_X1 #() 
NAND3_X1_2267_ (
  .A1({ S15667 }),
  .A2({ S25957[276] }),
  .A3({ S15849 }),
  .ZN({ S15850 })
);
OAI211_X1 #() 
OAI211_X1_722_ (
  .A({ S15765 }),
  .B({ S13772 }),
  .C1({ S25957[275] }),
  .C2({ S15515 }),
  .ZN({ S15851 })
);
NAND3_X1 #() 
NAND3_X1_2268_ (
  .A1({ S15851 }),
  .A2({ S15850 }),
  .A3({ S25957[277] }),
  .ZN({ S15852 })
);
OAI211_X1 #() 
OAI211_X1_723_ (
  .A({ S15852 }),
  .B({ S15585 }),
  .C1({ S15848 }),
  .C2({ S25957[277] }),
  .ZN({ S15853 })
);
NAND3_X1 #() 
NAND3_X1_2269_ (
  .A1({ S15839 }),
  .A2({ S15517 }),
  .A3({ S15853 }),
  .ZN({ S15854 })
);
AOI21_X1 #() 
AOI21_X1_1177_ (
  .A({ S25957[275] }),
  .B1({ S15611 }),
  .B2({ S15740 }),
  .ZN({ S15856 })
);
AOI21_X1 #() 
AOI21_X1_1178_ (
  .A({ S15856 }),
  .B1({ S15783 }),
  .B2({ S25957[275] }),
  .ZN({ S15857 })
);
NAND2_X1 #() 
NAND2_X1_1985_ (
  .A1({ S15857 }),
  .A2({ S25957[276] }),
  .ZN({ S15858 })
);
INV_X1 #() 
INV_X1_635_ (
  .A({ S15518 }),
  .ZN({ S15859 })
);
AOI22_X1 #() 
AOI22_X1_262_ (
  .A1({ S15600 }),
  .A2({ S15549 }),
  .B1({ S25957[273] }),
  .B2({ S25957[272] }),
  .ZN({ S15860 })
);
OAI221_X1 #() 
OAI221_X1_44_ (
  .A({ S25957[276] }),
  .B1({ S15795 }),
  .B2({ S15859 }),
  .C1({ S15860 }),
  .C2({ S25957[275] }),
  .ZN({ S15861 })
);
NAND2_X1 #() 
NAND2_X1_1986_ (
  .A1({ S15597 }),
  .A2({ S15596 }),
  .ZN({ S15862 })
);
NAND2_X1 #() 
NAND2_X1_1987_ (
  .A1({ S15862 }),
  .A2({ S32 }),
  .ZN({ S15863 })
);
NAND4_X1 #() 
NAND4_X1_283_ (
  .A1({ S25957[275] }),
  .A2({ S25957[274] }),
  .A3({ S15519 }),
  .A4({ S25957[273] }),
  .ZN({ S15864 })
);
AND3_X1 #() 
AND3_X1_91_ (
  .A1({ S15864 }),
  .A2({ S15774 }),
  .A3({ S13772 }),
  .ZN({ S15865 })
);
AOI21_X1 #() 
AOI21_X1_1179_ (
  .A({ S15621 }),
  .B1({ S15863 }),
  .B2({ S15865 }),
  .ZN({ S15867 })
);
OAI21_X1 #() 
OAI21_X1_1102_ (
  .A({ S32 }),
  .B1({ S15626 }),
  .B2({ S15662 }),
  .ZN({ S15868 })
);
AOI21_X1 #() 
AOI21_X1_1180_ (
  .A({ S25957[276] }),
  .B1({ S15601 }),
  .B2({ S15527 }),
  .ZN({ S15869 })
);
AOI21_X1 #() 
AOI21_X1_1181_ (
  .A({ S25957[277] }),
  .B1({ S15868 }),
  .B2({ S15869 }),
  .ZN({ S15870 })
);
AOI22_X1 #() 
AOI22_X1_263_ (
  .A1({ S15858 }),
  .A2({ S15870 }),
  .B1({ S15867 }),
  .B2({ S15861 }),
  .ZN({ S15871 })
);
OAI21_X1 #() 
OAI21_X1_1103_ (
  .A({ S32 }),
  .B1({ S53 }),
  .B2({ S15553 }),
  .ZN({ S15872 })
);
NAND3_X1 #() 
NAND3_X1_2270_ (
  .A1({ S15872 }),
  .A2({ S15774 }),
  .A3({ S25957[276] }),
  .ZN({ S15873 })
);
NAND3_X1 #() 
NAND3_X1_2271_ (
  .A1({ S15600 }),
  .A2({ S32 }),
  .A3({ S15519 }),
  .ZN({ S15874 })
);
NAND3_X1 #() 
NAND3_X1_2272_ (
  .A1({ S15609 }),
  .A2({ S13772 }),
  .A3({ S15874 }),
  .ZN({ S15875 })
);
NAND3_X1 #() 
NAND3_X1_2273_ (
  .A1({ S15875 }),
  .A2({ S25957[277] }),
  .A3({ S15873 }),
  .ZN({ S15876 })
);
INV_X1 #() 
INV_X1_636_ (
  .A({ S15845 }),
  .ZN({ S15878 })
);
NAND3_X1 #() 
NAND3_X1_2274_ (
  .A1({ S15567 }),
  .A2({ S15531 }),
  .A3({ S32 }),
  .ZN({ S15879 })
);
NAND3_X1 #() 
NAND3_X1_2275_ (
  .A1({ S15879 }),
  .A2({ S15615 }),
  .A3({ S13772 }),
  .ZN({ S15880 })
);
OAI211_X1 #() 
OAI211_X1_724_ (
  .A({ S15621 }),
  .B({ S15880 }),
  .C1({ S15878 }),
  .C2({ S15681 }),
  .ZN({ S15881 })
);
NAND2_X1 #() 
NAND2_X1_1988_ (
  .A1({ S15881 }),
  .A2({ S15876 }),
  .ZN({ S15882 })
);
NAND2_X1 #() 
NAND2_X1_1989_ (
  .A1({ S15882 }),
  .A2({ S25957[278] }),
  .ZN({ S15883 })
);
OAI21_X1 #() 
OAI21_X1_1104_ (
  .A({ S15883 }),
  .B1({ S15871 }),
  .B2({ S25957[278] }),
  .ZN({ S15884 })
);
NAND2_X1 #() 
NAND2_X1_1990_ (
  .A1({ S15884 }),
  .A2({ S25957[279] }),
  .ZN({ S15885 })
);
NAND3_X1 #() 
NAND3_X1_2276_ (
  .A1({ S15885 }),
  .A2({ S25957[380] }),
  .A3({ S15854 }),
  .ZN({ S15886 })
);
INV_X1 #() 
INV_X1_637_ (
  .A({ S25957[380] }),
  .ZN({ S15887 })
);
OAI211_X1 #() 
OAI211_X1_725_ (
  .A({ S15883 }),
  .B({ S25957[279] }),
  .C1({ S15871 }),
  .C2({ S25957[278] }),
  .ZN({ S15889 })
);
AOI211_X1 #() 
AOI211_X1_28_ (
  .A({ S15832 }),
  .B({ S15621 }),
  .C1({ S15836 }),
  .C2({ S15834 }),
  .ZN({ S15890 })
);
NOR2_X1 #() 
NOR2_X1_462_ (
  .A1({ S15831 }),
  .A2({ S25957[277] }),
  .ZN({ S15891 })
);
OAI21_X1 #() 
OAI21_X1_1105_ (
  .A({ S25957[278] }),
  .B1({ S15891 }),
  .B2({ S15890 }),
  .ZN({ S15892 })
);
AOI21_X1 #() 
AOI21_X1_1182_ (
  .A({ S25957[277] }),
  .B1({ S15843 }),
  .B2({ S15847 }),
  .ZN({ S15893 })
);
INV_X1 #() 
INV_X1_638_ (
  .A({ S15852 }),
  .ZN({ S15894 })
);
OAI21_X1 #() 
OAI21_X1_1106_ (
  .A({ S15585 }),
  .B1({ S15894 }),
  .B2({ S15893 }),
  .ZN({ S15895 })
);
NAND3_X1 #() 
NAND3_X1_2277_ (
  .A1({ S15895 }),
  .A2({ S15892 }),
  .A3({ S15517 }),
  .ZN({ S15896 })
);
NAND3_X1 #() 
NAND3_X1_2278_ (
  .A1({ S15896 }),
  .A2({ S15887 }),
  .A3({ S15889 }),
  .ZN({ S15897 })
);
AOI21_X1 #() 
AOI21_X1_1183_ (
  .A({ S25957[444] }),
  .B1({ S15886 }),
  .B2({ S15897 }),
  .ZN({ S15898 })
);
INV_X1 #() 
INV_X1_639_ (
  .A({ S25957[444] }),
  .ZN({ S15900 })
);
NAND3_X1 #() 
NAND3_X1_2279_ (
  .A1({ S15885 }),
  .A2({ S15887 }),
  .A3({ S15854 }),
  .ZN({ S15901 })
);
NAND3_X1 #() 
NAND3_X1_2280_ (
  .A1({ S15896 }),
  .A2({ S25957[380] }),
  .A3({ S15889 }),
  .ZN({ S15902 })
);
AOI21_X1 #() 
AOI21_X1_1184_ (
  .A({ S15900 }),
  .B1({ S15901 }),
  .B2({ S15902 }),
  .ZN({ S15903 })
);
OAI21_X1 #() 
OAI21_X1_1107_ (
  .A({ S14852 }),
  .B1({ S15898 }),
  .B2({ S15903 }),
  .ZN({ S15904 })
);
NAND3_X1 #() 
NAND3_X1_2281_ (
  .A1({ S15901 }),
  .A2({ S15902 }),
  .A3({ S15900 }),
  .ZN({ S15905 })
);
NAND3_X1 #() 
NAND3_X1_2282_ (
  .A1({ S15886 }),
  .A2({ S15897 }),
  .A3({ S25957[444] }),
  .ZN({ S15906 })
);
NAND3_X1 #() 
NAND3_X1_2283_ (
  .A1({ S15905 }),
  .A2({ S15906 }),
  .A3({ S25957[284] }),
  .ZN({ S15907 })
);
NAND2_X1 #() 
NAND2_X1_1991_ (
  .A1({ S15904 }),
  .A2({ S15907 }),
  .ZN({ S25957[156] })
);
NAND2_X1 #() 
NAND2_X1_1992_ (
  .A1({ S2001 }),
  .A2({ S2002 }),
  .ZN({ S25957[859] })
);
XOR2_X1 #() 
XOR2_X1_29_ (
  .A({ S10161 }),
  .B({ S25957[859] }),
  .Z({ S25957[603] })
);
NAND2_X1 #() 
NAND2_X1_1993_ (
  .A1({ S13148 }),
  .A2({ S13157 }),
  .ZN({ S15909 })
);
XOR2_X1 #() 
XOR2_X1_30_ (
  .A({ S15909 }),
  .B({ S25957[603] }),
  .Z({ S15910 })
);
INV_X1 #() 
INV_X1_640_ (
  .A({ S15910 }),
  .ZN({ S25957[347] })
);
NAND2_X1 #() 
NAND2_X1_1994_ (
  .A1({ S10239 }),
  .A2({ S10214 }),
  .ZN({ S25957[507] })
);
XNOR2_X1 #() 
XNOR2_X1_65_ (
  .A({ S15909 }),
  .B({ S25957[507] }),
  .ZN({ S25957[379] })
);
INV_X1 #() 
INV_X1_641_ (
  .A({ S25957[379] }),
  .ZN({ S15911 })
);
OAI211_X1 #() 
OAI211_X1_726_ (
  .A({ S15650 }),
  .B({ S25957[276] }),
  .C1({ S15623 }),
  .C2({ S15622 }),
  .ZN({ S15912 })
);
NAND3_X1 #() 
NAND3_X1_2284_ (
  .A1({ S15600 }),
  .A2({ S15518 }),
  .A3({ S32 }),
  .ZN({ S15913 })
);
AOI21_X1 #() 
AOI21_X1_1185_ (
  .A({ S25957[272] }),
  .B1({ S25957[274] }),
  .B2({ S25957[273] }),
  .ZN({ S15914 })
);
AOI21_X1 #() 
AOI21_X1_1186_ (
  .A({ S25957[276] }),
  .B1({ S15914 }),
  .B2({ S25957[275] }),
  .ZN({ S15916 })
);
AOI21_X1 #() 
AOI21_X1_1187_ (
  .A({ S15621 }),
  .B1({ S15916 }),
  .B2({ S15913 }),
  .ZN({ S15917 })
);
NAND2_X1 #() 
NAND2_X1_1995_ (
  .A1({ S15912 }),
  .A2({ S15917 }),
  .ZN({ S15918 })
);
NAND4_X1 #() 
NAND4_X1_284_ (
  .A1({ S25957[276] }),
  .A2({ S15549 }),
  .A3({ S15515 }),
  .A4({ S32 }),
  .ZN({ S15919 })
);
INV_X1 #() 
INV_X1_642_ (
  .A({ S15919 }),
  .ZN({ S15920 })
);
AOI21_X1 #() 
AOI21_X1_1188_ (
  .A({ S25957[276] }),
  .B1({ S15693 }),
  .B2({ S15532 }),
  .ZN({ S15921 })
);
OAI21_X1 #() 
OAI21_X1_1108_ (
  .A({ S15621 }),
  .B1({ S15921 }),
  .B2({ S15920 }),
  .ZN({ S15922 })
);
AOI21_X1 #() 
AOI21_X1_1189_ (
  .A({ S15585 }),
  .B1({ S15918 }),
  .B2({ S15922 }),
  .ZN({ S15923 })
);
INV_X1 #() 
INV_X1_643_ (
  .A({ S15923 }),
  .ZN({ S15924 })
);
OAI21_X1 #() 
OAI21_X1_1109_ (
  .A({ S25957[275] }),
  .B1({ S15515 }),
  .B2({ S25957[274] }),
  .ZN({ S15925 })
);
OAI21_X1 #() 
OAI21_X1_1110_ (
  .A({ S13772 }),
  .B1({ S15925 }),
  .B2({ S15732 }),
  .ZN({ S15927 })
);
OAI211_X1 #() 
OAI211_X1_727_ (
  .A({ S25957[275] }),
  .B({ S53 }),
  .C1({ S15515 }),
  .C2({ S25957[274] }),
  .ZN({ S15928 })
);
NAND3_X1 #() 
NAND3_X1_2285_ (
  .A1({ S15794 }),
  .A2({ S15928 }),
  .A3({ S25957[276] }),
  .ZN({ S15929 })
);
OAI21_X1 #() 
OAI21_X1_1111_ (
  .A({ S15929 }),
  .B1({ S15927 }),
  .B2({ S15595 }),
  .ZN({ S15930 })
);
NAND2_X1 #() 
NAND2_X1_1996_ (
  .A1({ S15930 }),
  .A2({ S15621 }),
  .ZN({ S15931 })
);
NAND2_X1 #() 
NAND2_X1_1997_ (
  .A1({ S15649 }),
  .A2({ S25957[275] }),
  .ZN({ S15932 })
);
INV_X1 #() 
INV_X1_644_ (
  .A({ S15932 }),
  .ZN({ S15933 })
);
AOI21_X1 #() 
AOI21_X1_1190_ (
  .A({ S25957[275] }),
  .B1({ S15600 }),
  .B2({ S25957[272] }),
  .ZN({ S15934 })
);
OAI21_X1 #() 
OAI21_X1_1112_ (
  .A({ S13772 }),
  .B1({ S15933 }),
  .B2({ S15934 }),
  .ZN({ S15935 })
);
NAND2_X1 #() 
NAND2_X1_1998_ (
  .A1({ S15528 }),
  .A2({ S25957[275] }),
  .ZN({ S15936 })
);
OAI21_X1 #() 
OAI21_X1_1113_ (
  .A({ S15936 }),
  .B1({ S15793 }),
  .B2({ S25957[275] }),
  .ZN({ S15938 })
);
NAND2_X1 #() 
NAND2_X1_1999_ (
  .A1({ S15938 }),
  .A2({ S25957[276] }),
  .ZN({ S15939 })
);
NAND3_X1 #() 
NAND3_X1_2286_ (
  .A1({ S15939 }),
  .A2({ S15935 }),
  .A3({ S25957[277] }),
  .ZN({ S15940 })
);
NAND3_X1 #() 
NAND3_X1_2287_ (
  .A1({ S15931 }),
  .A2({ S15940 }),
  .A3({ S15585 }),
  .ZN({ S15941 })
);
NAND3_X1 #() 
NAND3_X1_2288_ (
  .A1({ S15924 }),
  .A2({ S15941 }),
  .A3({ S15517 }),
  .ZN({ S15942 })
);
NAND3_X1 #() 
NAND3_X1_2289_ (
  .A1({ S15571 }),
  .A2({ S15778 }),
  .A3({ S25957[275] }),
  .ZN({ S15943 })
);
NAND3_X1 #() 
NAND3_X1_2290_ (
  .A1({ S15734 }),
  .A2({ S32 }),
  .A3({ S15518 }),
  .ZN({ S15944 })
);
AND2_X1 #() 
AND2_X1_122_ (
  .A1({ S15944 }),
  .A2({ S15943 }),
  .ZN({ S15945 })
);
NAND2_X1 #() 
NAND2_X1_2000_ (
  .A1({ S15601 }),
  .A2({ S53 }),
  .ZN({ S15946 })
);
NAND3_X1 #() 
NAND3_X1_2291_ (
  .A1({ S15520 }),
  .A2({ S32 }),
  .A3({ S15518 }),
  .ZN({ S15947 })
);
NAND3_X1 #() 
NAND3_X1_2292_ (
  .A1({ S15946 }),
  .A2({ S15947 }),
  .A3({ S25957[276] }),
  .ZN({ S15949 })
);
OAI211_X1 #() 
OAI211_X1_728_ (
  .A({ S25957[277] }),
  .B({ S15949 }),
  .C1({ S15945 }),
  .C2({ S25957[276] }),
  .ZN({ S15950 })
);
NAND3_X1 #() 
NAND3_X1_2293_ (
  .A1({ S15577 }),
  .A2({ S32 }),
  .A3({ S15784 }),
  .ZN({ S15951 })
);
NAND2_X1 #() 
NAND2_X1_2001_ (
  .A1({ S15951 }),
  .A2({ S15695 }),
  .ZN({ S15952 })
);
NAND2_X1 #() 
NAND2_X1_2002_ (
  .A1({ S15952 }),
  .A2({ S25957[276] }),
  .ZN({ S15953 })
);
OAI21_X1 #() 
OAI21_X1_1114_ (
  .A({ S13772 }),
  .B1({ S32 }),
  .B2({ S15553 }),
  .ZN({ S15954 })
);
NOR2_X1 #() 
NOR2_X1_463_ (
  .A1({ S15954 }),
  .A2({ S15655 }),
  .ZN({ S15955 })
);
INV_X1 #() 
INV_X1_645_ (
  .A({ S15955 }),
  .ZN({ S15956 })
);
NAND3_X1 #() 
NAND3_X1_2294_ (
  .A1({ S15953 }),
  .A2({ S15621 }),
  .A3({ S15956 }),
  .ZN({ S15957 })
);
NAND3_X1 #() 
NAND3_X1_2295_ (
  .A1({ S15957 }),
  .A2({ S15950 }),
  .A3({ S25957[278] }),
  .ZN({ S15958 })
);
OAI211_X1 #() 
OAI211_X1_729_ (
  .A({ S25957[276] }),
  .B({ S15879 }),
  .C1({ S15925 }),
  .C2({ S15762 }),
  .ZN({ S15960 })
);
AOI21_X1 #() 
AOI21_X1_1191_ (
  .A({ S32 }),
  .B1({ S25957[273] }),
  .B2({ S15553 }),
  .ZN({ S15961 })
);
AOI22_X1 #() 
AOI22_X1_264_ (
  .A1({ S15961 }),
  .A2({ S15647 }),
  .B1({ S15579 }),
  .B2({ S53 }),
  .ZN({ S15962 })
);
OAI211_X1 #() 
OAI211_X1_730_ (
  .A({ S15621 }),
  .B({ S15960 }),
  .C1({ S15962 }),
  .C2({ S25957[276] }),
  .ZN({ S15963 })
);
OAI211_X1 #() 
OAI211_X1_731_ (
  .A({ S15786 }),
  .B({ S25957[276] }),
  .C1({ S15936 }),
  .C2({ S15570 }),
  .ZN({ S15964 })
);
NAND3_X1 #() 
NAND3_X1_2296_ (
  .A1({ S15647 }),
  .A2({ S32 }),
  .A3({ S15567 }),
  .ZN({ S15965 })
);
NAND4_X1 #() 
NAND4_X1_285_ (
  .A1({ S15531 }),
  .A2({ S15653 }),
  .A3({ S25957[275] }),
  .A4({ S25957[273] }),
  .ZN({ S15966 })
);
NAND3_X1 #() 
NAND3_X1_2297_ (
  .A1({ S15965 }),
  .A2({ S13772 }),
  .A3({ S15966 }),
  .ZN({ S15967 })
);
NAND3_X1 #() 
NAND3_X1_2298_ (
  .A1({ S15967 }),
  .A2({ S15964 }),
  .A3({ S25957[277] }),
  .ZN({ S15968 })
);
NAND3_X1 #() 
NAND3_X1_2299_ (
  .A1({ S15968 }),
  .A2({ S15963 }),
  .A3({ S15585 }),
  .ZN({ S15969 })
);
NAND3_X1 #() 
NAND3_X1_2300_ (
  .A1({ S15958 }),
  .A2({ S25957[279] }),
  .A3({ S15969 }),
  .ZN({ S15971 })
);
NAND3_X1 #() 
NAND3_X1_2301_ (
  .A1({ S15942 }),
  .A2({ S15971 }),
  .A3({ S15911 }),
  .ZN({ S15972 })
);
NAND3_X1 #() 
NAND3_X1_2302_ (
  .A1({ S15600 }),
  .A2({ S13772 }),
  .A3({ S25957[272] }),
  .ZN({ S15973 })
);
OAI221_X1 #() 
OAI221_X1_45_ (
  .A({ S25957[277] }),
  .B1({ S15933 }),
  .B2({ S15973 }),
  .C1({ S15938 }),
  .C2({ S13772 }),
  .ZN({ S15974 })
);
OAI211_X1 #() 
OAI211_X1_732_ (
  .A({ S15929 }),
  .B({ S15621 }),
  .C1({ S15595 }),
  .C2({ S15927 }),
  .ZN({ S15975 })
);
AOI21_X1 #() 
AOI21_X1_1192_ (
  .A({ S25957[278] }),
  .B1({ S15974 }),
  .B2({ S15975 }),
  .ZN({ S15976 })
);
OAI21_X1 #() 
OAI21_X1_1115_ (
  .A({ S15517 }),
  .B1({ S15976 }),
  .B2({ S15923 }),
  .ZN({ S15977 })
);
AOI21_X1 #() 
AOI21_X1_1193_ (
  .A({ S25957[276] }),
  .B1({ S15944 }),
  .B2({ S15943 }),
  .ZN({ S15978 })
);
AND3_X1 #() 
AND3_X1_92_ (
  .A1({ S15946 }),
  .A2({ S15947 }),
  .A3({ S25957[276] }),
  .ZN({ S15979 })
);
OAI21_X1 #() 
OAI21_X1_1116_ (
  .A({ S25957[277] }),
  .B1({ S15979 }),
  .B2({ S15978 }),
  .ZN({ S15980 })
);
AOI21_X1 #() 
AOI21_X1_1194_ (
  .A({ S13772 }),
  .B1({ S15951 }),
  .B2({ S15695 }),
  .ZN({ S15982 })
);
OAI21_X1 #() 
OAI21_X1_1117_ (
  .A({ S15621 }),
  .B1({ S15982 }),
  .B2({ S15955 }),
  .ZN({ S15983 })
);
AOI21_X1 #() 
AOI21_X1_1195_ (
  .A({ S15585 }),
  .B1({ S15980 }),
  .B2({ S15983 }),
  .ZN({ S15984 })
);
INV_X1 #() 
INV_X1_646_ (
  .A({ S15969 }),
  .ZN({ S15985 })
);
OAI21_X1 #() 
OAI21_X1_1118_ (
  .A({ S25957[279] }),
  .B1({ S15984 }),
  .B2({ S15985 }),
  .ZN({ S15986 })
);
NAND3_X1 #() 
NAND3_X1_2303_ (
  .A1({ S15986 }),
  .A2({ S15977 }),
  .A3({ S25957[379] }),
  .ZN({ S15987 })
);
NAND3_X1 #() 
NAND3_X1_2304_ (
  .A1({ S15987 }),
  .A2({ S25957[347] }),
  .A3({ S15972 }),
  .ZN({ S15988 })
);
NAND3_X1 #() 
NAND3_X1_2305_ (
  .A1({ S15942 }),
  .A2({ S15971 }),
  .A3({ S25957[379] }),
  .ZN({ S15989 })
);
NAND3_X1 #() 
NAND3_X1_2306_ (
  .A1({ S15986 }),
  .A2({ S15977 }),
  .A3({ S15911 }),
  .ZN({ S15990 })
);
NAND3_X1 #() 
NAND3_X1_2307_ (
  .A1({ S15990 }),
  .A2({ S15910 }),
  .A3({ S15989 }),
  .ZN({ S15991 })
);
NAND3_X1 #() 
NAND3_X1_2308_ (
  .A1({ S15988 }),
  .A2({ S15991 }),
  .A3({ S28 }),
  .ZN({ S15993 })
);
NAND3_X1 #() 
NAND3_X1_2309_ (
  .A1({ S15990 }),
  .A2({ S25957[347] }),
  .A3({ S15989 }),
  .ZN({ S15994 })
);
NAND3_X1 #() 
NAND3_X1_2310_ (
  .A1({ S15987 }),
  .A2({ S15910 }),
  .A3({ S15972 }),
  .ZN({ S15995 })
);
NAND3_X1 #() 
NAND3_X1_2311_ (
  .A1({ S15994 }),
  .A2({ S15995 }),
  .A3({ S25957[411] }),
  .ZN({ S15996 })
);
NAND2_X1 #() 
NAND2_X1_2003_ (
  .A1({ S15993 }),
  .A2({ S15996 }),
  .ZN({ S54 })
);
NAND3_X1 #() 
NAND3_X1_2312_ (
  .A1({ S15994 }),
  .A2({ S15995 }),
  .A3({ S28 }),
  .ZN({ S15997 })
);
NAND3_X1 #() 
NAND3_X1_2313_ (
  .A1({ S15988 }),
  .A2({ S15991 }),
  .A3({ S25957[411] }),
  .ZN({ S15998 })
);
NAND2_X1 #() 
NAND2_X1_2004_ (
  .A1({ S15997 }),
  .A2({ S15998 }),
  .ZN({ S25957[155] })
);
NOR2_X1 #() 
NOR2_X1_464_ (
  .A1({ S13207 }),
  .A2({ S13208 }),
  .ZN({ S25957[344] })
);
NAND2_X1 #() 
NAND2_X1_2005_ (
  .A1({ S10304 }),
  .A2({ S10281 }),
  .ZN({ S15999 })
);
XNOR2_X1 #() 
XNOR2_X1_66_ (
  .A({ S15999 }),
  .B({ S25957[632] }),
  .ZN({ S25957[504] })
);
NAND2_X1 #() 
NAND2_X1_2006_ (
  .A1({ S13185 }),
  .A2({ S13206 }),
  .ZN({ S16001 })
);
XNOR2_X1 #() 
XNOR2_X1_67_ (
  .A({ S16001 }),
  .B({ S25957[504] }),
  .ZN({ S25957[376] })
);
INV_X1 #() 
INV_X1_647_ (
  .A({ S25957[376] }),
  .ZN({ S16002 })
);
OAI211_X1 #() 
OAI211_X1_733_ (
  .A({ S15946 }),
  .B({ S25957[276] }),
  .C1({ S15540 }),
  .C2({ S15673 }),
  .ZN({ S16003 })
);
AOI22_X1 #() 
AOI22_X1_265_ (
  .A1({ S15681 }),
  .A2({ S15531 }),
  .B1({ S15674 }),
  .B2({ S32 }),
  .ZN({ S16004 })
);
NAND2_X1 #() 
NAND2_X1_2007_ (
  .A1({ S16004 }),
  .A2({ S13772 }),
  .ZN({ S16005 })
);
NAND3_X1 #() 
NAND3_X1_2314_ (
  .A1({ S16005 }),
  .A2({ S25957[277] }),
  .A3({ S16003 }),
  .ZN({ S16006 })
);
NAND2_X1 #() 
NAND2_X1_2008_ (
  .A1({ S15707 }),
  .A2({ S25957[275] }),
  .ZN({ S16007 })
);
NOR2_X1 #() 
NOR2_X1_465_ (
  .A1({ S53 }),
  .A2({ S15553 }),
  .ZN({ S16008 })
);
OAI21_X1 #() 
OAI21_X1_1119_ (
  .A({ S32 }),
  .B1({ S15670 }),
  .B2({ S16008 }),
  .ZN({ S16010 })
);
NAND3_X1 #() 
NAND3_X1_2315_ (
  .A1({ S16010 }),
  .A2({ S16007 }),
  .A3({ S13772 }),
  .ZN({ S16011 })
);
NAND2_X1 #() 
NAND2_X1_2009_ (
  .A1({ S15597 }),
  .A2({ S25957[275] }),
  .ZN({ S16012 })
);
OAI211_X1 #() 
OAI211_X1_734_ (
  .A({ S25957[276] }),
  .B({ S16012 }),
  .C1({ S15648 }),
  .C2({ S15644 }),
  .ZN({ S16013 })
);
NAND3_X1 #() 
NAND3_X1_2316_ (
  .A1({ S16011 }),
  .A2({ S16013 }),
  .A3({ S15621 }),
  .ZN({ S16014 })
);
NAND3_X1 #() 
NAND3_X1_2317_ (
  .A1({ S16006 }),
  .A2({ S16014 }),
  .A3({ S15585 }),
  .ZN({ S16015 })
);
AOI21_X1 #() 
AOI21_X1_1196_ (
  .A({ S25957[276] }),
  .B1({ S32 }),
  .B2({ S15533 }),
  .ZN({ S16016 })
);
OAI21_X1 #() 
OAI21_X1_1120_ (
  .A({ S15642 }),
  .B1({ S15622 }),
  .B2({ S15925 }),
  .ZN({ S16017 })
);
AOI22_X1 #() 
AOI22_X1_266_ (
  .A1({ S16017 }),
  .A2({ S25957[276] }),
  .B1({ S15663 }),
  .B2({ S16016 }),
  .ZN({ S16018 })
);
NAND3_X1 #() 
NAND3_X1_2318_ (
  .A1({ S15739 }),
  .A2({ S13772 }),
  .A3({ S15776 }),
  .ZN({ S16019 })
);
NAND3_X1 #() 
NAND3_X1_2319_ (
  .A1({ S15704 }),
  .A2({ S15541 }),
  .A3({ S15543 }),
  .ZN({ S16021 })
);
OAI211_X1 #() 
OAI211_X1_735_ (
  .A({ S16019 }),
  .B({ S15621 }),
  .C1({ S13772 }),
  .C2({ S16021 }),
  .ZN({ S16022 })
);
OAI211_X1 #() 
OAI211_X1_736_ (
  .A({ S16022 }),
  .B({ S25957[278] }),
  .C1({ S15621 }),
  .C2({ S16018 }),
  .ZN({ S16023 })
);
NAND3_X1 #() 
NAND3_X1_2320_ (
  .A1({ S16023 }),
  .A2({ S16015 }),
  .A3({ S15517 }),
  .ZN({ S16024 })
);
NAND3_X1 #() 
NAND3_X1_2321_ (
  .A1({ S15549 }),
  .A2({ S15515 }),
  .A3({ S32 }),
  .ZN({ S16025 })
);
AOI22_X1 #() 
AOI22_X1_267_ (
  .A1({ S15936 }),
  .A2({ S16025 }),
  .B1({ S15914 }),
  .B2({ S32 }),
  .ZN({ S16026 })
);
NAND4_X1 #() 
NAND4_X1_286_ (
  .A1({ S15872 }),
  .A2({ S15864 }),
  .A3({ S15774 }),
  .A4({ S13772 }),
  .ZN({ S16027 })
);
OAI211_X1 #() 
OAI211_X1_737_ (
  .A({ S25957[277] }),
  .B({ S16027 }),
  .C1({ S16026 }),
  .C2({ S13772 }),
  .ZN({ S16028 })
);
OAI211_X1 #() 
OAI211_X1_738_ (
  .A({ S25957[276] }),
  .B({ S15700 }),
  .C1({ S15576 }),
  .C2({ S25957[275] }),
  .ZN({ S16029 })
);
INV_X1 #() 
INV_X1_648_ (
  .A({ S16029 }),
  .ZN({ S16030 })
);
NAND2_X1 #() 
NAND2_X1_2010_ (
  .A1({ S15914 }),
  .A2({ S25957[275] }),
  .ZN({ S16032 })
);
NAND4_X1 #() 
NAND4_X1_287_ (
  .A1({ S15549 }),
  .A2({ S15533 }),
  .A3({ S53 }),
  .A4({ S32 }),
  .ZN({ S16033 })
);
AOI21_X1 #() 
AOI21_X1_1197_ (
  .A({ S25957[276] }),
  .B1({ S16032 }),
  .B2({ S16033 }),
  .ZN({ S16034 })
);
OAI21_X1 #() 
OAI21_X1_1121_ (
  .A({ S15621 }),
  .B1({ S16030 }),
  .B2({ S16034 }),
  .ZN({ S16035 })
);
NAND3_X1 #() 
NAND3_X1_2322_ (
  .A1({ S16035 }),
  .A2({ S16028 }),
  .A3({ S15585 }),
  .ZN({ S16036 })
);
NAND2_X1 #() 
NAND2_X1_2011_ (
  .A1({ S15835 }),
  .A2({ S15562 }),
  .ZN({ S16037 })
);
NAND2_X1 #() 
NAND2_X1_2012_ (
  .A1({ S16037 }),
  .A2({ S16016 }),
  .ZN({ S16038 })
);
NAND4_X1 #() 
NAND4_X1_288_ (
  .A1({ S15518 }),
  .A2({ S15539 }),
  .A3({ S25957[275] }),
  .A4({ S25957[274] }),
  .ZN({ S16039 })
);
OAI211_X1 #() 
OAI211_X1_739_ (
  .A({ S25957[276] }),
  .B({ S16039 }),
  .C1({ S15860 }),
  .C2({ S25957[275] }),
  .ZN({ S16040 })
);
NAND3_X1 #() 
NAND3_X1_2323_ (
  .A1({ S16038 }),
  .A2({ S15621 }),
  .A3({ S16040 }),
  .ZN({ S16041 })
);
NAND3_X1 #() 
NAND3_X1_2324_ (
  .A1({ S15658 }),
  .A2({ S15784 }),
  .A3({ S32 }),
  .ZN({ S16043 })
);
AND2_X1 #() 
AND2_X1_123_ (
  .A1({ S15532 }),
  .A2({ S13772 }),
  .ZN({ S16044 })
);
NAND3_X1 #() 
NAND3_X1_2325_ (
  .A1({ S15539 }),
  .A2({ S25957[275] }),
  .A3({ S25957[274] }),
  .ZN({ S16045 })
);
NAND3_X1 #() 
NAND3_X1_2326_ (
  .A1({ S15841 }),
  .A2({ S15683 }),
  .A3({ S16045 }),
  .ZN({ S16046 })
);
AOI22_X1 #() 
AOI22_X1_268_ (
  .A1({ S16044 }),
  .A2({ S16043 }),
  .B1({ S16046 }),
  .B2({ S25957[276] }),
  .ZN({ S16047 })
);
OAI211_X1 #() 
OAI211_X1_740_ (
  .A({ S16041 }),
  .B({ S25957[278] }),
  .C1({ S16047 }),
  .C2({ S15621 }),
  .ZN({ S16048 })
);
NAND3_X1 #() 
NAND3_X1_2327_ (
  .A1({ S16048 }),
  .A2({ S16036 }),
  .A3({ S25957[279] }),
  .ZN({ S16049 })
);
NAND3_X1 #() 
NAND3_X1_2328_ (
  .A1({ S16024 }),
  .A2({ S16049 }),
  .A3({ S16002 }),
  .ZN({ S16050 })
);
AOI22_X1 #() 
AOI22_X1_269_ (
  .A1({ S15712 }),
  .A2({ S32 }),
  .B1({ S15797 }),
  .B2({ S15551 }),
  .ZN({ S16051 })
);
OAI211_X1 #() 
OAI211_X1_741_ (
  .A({ S15585 }),
  .B({ S16029 }),
  .C1({ S16051 }),
  .C2({ S25957[276] }),
  .ZN({ S16052 })
);
AOI21_X1 #() 
AOI21_X1_1198_ (
  .A({ S25957[275] }),
  .B1({ S15571 }),
  .B2({ S15778 }),
  .ZN({ S16054 })
);
AND4_X1 #() 
AND4_X1_5_ (
  .A1({ S25957[275] }),
  .A2({ S15518 }),
  .A3({ S15539 }),
  .A4({ S25957[274] }),
  .ZN({ S16055 })
);
OAI21_X1 #() 
OAI21_X1_1122_ (
  .A({ S25957[276] }),
  .B1({ S16054 }),
  .B2({ S16055 }),
  .ZN({ S16056 })
);
NAND2_X1 #() 
NAND2_X1_2013_ (
  .A1({ S15776 }),
  .A2({ S15802 }),
  .ZN({ S16057 })
);
NAND2_X1 #() 
NAND2_X1_2014_ (
  .A1({ S16057 }),
  .A2({ S13772 }),
  .ZN({ S16058 })
);
NAND3_X1 #() 
NAND3_X1_2329_ (
  .A1({ S16056 }),
  .A2({ S25957[278] }),
  .A3({ S16058 }),
  .ZN({ S16059 })
);
AOI21_X1 #() 
AOI21_X1_1199_ (
  .A({ S15517 }),
  .B1({ S16059 }),
  .B2({ S16052 }),
  .ZN({ S16060 })
);
NAND2_X1 #() 
NAND2_X1_2015_ (
  .A1({ S16021 }),
  .A2({ S25957[276] }),
  .ZN({ S16061 })
);
AOI22_X1 #() 
AOI22_X1_270_ (
  .A1({ S15835 }),
  .A2({ S25957[275] }),
  .B1({ S15738 }),
  .B2({ S15567 }),
  .ZN({ S16062 })
);
OAI211_X1 #() 
OAI211_X1_742_ (
  .A({ S16061 }),
  .B({ S25957[278] }),
  .C1({ S16062 }),
  .C2({ S25957[276] }),
  .ZN({ S16063 })
);
AOI21_X1 #() 
AOI21_X1_1200_ (
  .A({ S32 }),
  .B1({ S15662 }),
  .B2({ S15518 }),
  .ZN({ S16065 })
);
AOI21_X1 #() 
AOI21_X1_1201_ (
  .A({ S25957[275] }),
  .B1({ S15577 }),
  .B2({ S15567 }),
  .ZN({ S16066 })
);
OAI21_X1 #() 
OAI21_X1_1123_ (
  .A({ S25957[276] }),
  .B1({ S16066 }),
  .B2({ S16065 }),
  .ZN({ S16067 })
);
NAND3_X1 #() 
NAND3_X1_2330_ (
  .A1({ S15706 }),
  .A2({ S25957[275] }),
  .A3({ S53 }),
  .ZN({ S16068 })
);
OAI211_X1 #() 
OAI211_X1_743_ (
  .A({ S16068 }),
  .B({ S13772 }),
  .C1({ S15670 }),
  .C2({ S15872 }),
  .ZN({ S16069 })
);
NAND3_X1 #() 
NAND3_X1_2331_ (
  .A1({ S16067 }),
  .A2({ S15585 }),
  .A3({ S16069 }),
  .ZN({ S16070 })
);
AOI21_X1 #() 
AOI21_X1_1202_ (
  .A({ S25957[279] }),
  .B1({ S16070 }),
  .B2({ S16063 }),
  .ZN({ S16071 })
);
OAI21_X1 #() 
OAI21_X1_1124_ (
  .A({ S15621 }),
  .B1({ S16071 }),
  .B2({ S16060 }),
  .ZN({ S16072 })
);
NAND2_X1 #() 
NAND2_X1_2016_ (
  .A1({ S15663 }),
  .A2({ S16016 }),
  .ZN({ S16073 })
);
NAND2_X1 #() 
NAND2_X1_2017_ (
  .A1({ S16017 }),
  .A2({ S25957[276] }),
  .ZN({ S16074 })
);
NAND3_X1 #() 
NAND3_X1_2332_ (
  .A1({ S16074 }),
  .A2({ S25957[278] }),
  .A3({ S16073 }),
  .ZN({ S16076 })
);
OAI21_X1 #() 
OAI21_X1_1125_ (
  .A({ S25957[276] }),
  .B1({ S15798 }),
  .B2({ S15840 }),
  .ZN({ S16077 })
);
OAI211_X1 #() 
OAI211_X1_744_ (
  .A({ S15585 }),
  .B({ S16077 }),
  .C1({ S16004 }),
  .C2({ S25957[276] }),
  .ZN({ S16078 })
);
AOI21_X1 #() 
AOI21_X1_1203_ (
  .A({ S25957[279] }),
  .B1({ S16076 }),
  .B2({ S16078 }),
  .ZN({ S16079 })
);
AOI21_X1 #() 
AOI21_X1_1204_ (
  .A({ S25957[275] }),
  .B1({ S15567 }),
  .B2({ S25957[272] }),
  .ZN({ S16080 })
);
AOI21_X1 #() 
AOI21_X1_1205_ (
  .A({ S32 }),
  .B1({ S15732 }),
  .B2({ S15527 }),
  .ZN({ S16081 })
);
NAND3_X1 #() 
NAND3_X1_2333_ (
  .A1({ S15551 }),
  .A2({ S32 }),
  .A3({ S15519 }),
  .ZN({ S16082 })
);
OAI211_X1 #() 
OAI211_X1_745_ (
  .A({ S25957[276] }),
  .B({ S16082 }),
  .C1({ S16081 }),
  .C2({ S16080 }),
  .ZN({ S16083 })
);
NAND3_X1 #() 
NAND3_X1_2334_ (
  .A1({ S15872 }),
  .A2({ S15864 }),
  .A3({ S15774 }),
  .ZN({ S16084 })
);
NAND2_X1 #() 
NAND2_X1_2018_ (
  .A1({ S16084 }),
  .A2({ S13772 }),
  .ZN({ S16085 })
);
NAND3_X1 #() 
NAND3_X1_2335_ (
  .A1({ S16085 }),
  .A2({ S16083 }),
  .A3({ S15585 }),
  .ZN({ S16087 })
);
NAND3_X1 #() 
NAND3_X1_2336_ (
  .A1({ S16043 }),
  .A2({ S13772 }),
  .A3({ S15532 }),
  .ZN({ S16088 })
);
NAND2_X1 #() 
NAND2_X1_2019_ (
  .A1({ S16046 }),
  .A2({ S25957[276] }),
  .ZN({ S16089 })
);
NAND3_X1 #() 
NAND3_X1_2337_ (
  .A1({ S16089 }),
  .A2({ S16088 }),
  .A3({ S25957[278] }),
  .ZN({ S16090 })
);
AOI21_X1 #() 
AOI21_X1_1206_ (
  .A({ S15517 }),
  .B1({ S16087 }),
  .B2({ S16090 }),
  .ZN({ S16091 })
);
OAI21_X1 #() 
OAI21_X1_1126_ (
  .A({ S25957[277] }),
  .B1({ S16079 }),
  .B2({ S16091 }),
  .ZN({ S16092 })
);
NAND3_X1 #() 
NAND3_X1_2338_ (
  .A1({ S16072 }),
  .A2({ S16092 }),
  .A3({ S25957[376] }),
  .ZN({ S16093 })
);
AOI21_X1 #() 
AOI21_X1_1207_ (
  .A({ S25957[344] }),
  .B1({ S16093 }),
  .B2({ S16050 }),
  .ZN({ S16094 })
);
INV_X1 #() 
INV_X1_649_ (
  .A({ S25957[344] }),
  .ZN({ S16095 })
);
NAND3_X1 #() 
NAND3_X1_2339_ (
  .A1({ S16024 }),
  .A2({ S16049 }),
  .A3({ S25957[376] }),
  .ZN({ S16096 })
);
NAND3_X1 #() 
NAND3_X1_2340_ (
  .A1({ S16072 }),
  .A2({ S16092 }),
  .A3({ S16002 }),
  .ZN({ S16097 })
);
AOI21_X1 #() 
AOI21_X1_1208_ (
  .A({ S16095 }),
  .B1({ S16097 }),
  .B2({ S16096 }),
  .ZN({ S16098 })
);
OAI21_X1 #() 
OAI21_X1_1127_ (
  .A({ S25957[408] }),
  .B1({ S16094 }),
  .B2({ S16098 }),
  .ZN({ S16099 })
);
NAND3_X1 #() 
NAND3_X1_2341_ (
  .A1({ S16097 }),
  .A2({ S16096 }),
  .A3({ S16095 }),
  .ZN({ S16100 })
);
NAND3_X1 #() 
NAND3_X1_2342_ (
  .A1({ S16093 }),
  .A2({ S16050 }),
  .A3({ S25957[344] }),
  .ZN({ S16101 })
);
NAND3_X1 #() 
NAND3_X1_2343_ (
  .A1({ S16100 }),
  .A2({ S16101 }),
  .A3({ S12012 }),
  .ZN({ S16102 })
);
NAND2_X1 #() 
NAND2_X1_2020_ (
  .A1({ S16099 }),
  .A2({ S16102 }),
  .ZN({ S25957[152] })
);
NAND2_X1 #() 
NAND2_X1_2021_ (
  .A1({ S10405 }),
  .A2({ S10404 }),
  .ZN({ S16103 })
);
NAND2_X1 #() 
NAND2_X1_2022_ (
  .A1({ S7462 }),
  .A2({ S7461 }),
  .ZN({ S25957[633] })
);
XNOR2_X1 #() 
XNOR2_X1_68_ (
  .A({ S10399 }),
  .B({ S25957[633] }),
  .ZN({ S25957[505] })
);
NAND2_X1 #() 
NAND2_X1_2023_ (
  .A1({ S13266 }),
  .A2({ S13293 }),
  .ZN({ S16105 })
);
XOR2_X1 #() 
XOR2_X1_31_ (
  .A({ S16105 }),
  .B({ S25957[505] }),
  .Z({ S25957[377] })
);
OAI21_X1 #() 
OAI21_X1_1128_ (
  .A({ S25957[276] }),
  .B1({ S15586 }),
  .B2({ S15694 }),
  .ZN({ S16106 })
);
OAI211_X1 #() 
OAI211_X1_746_ (
  .A({ S13772 }),
  .B({ S15733 }),
  .C1({ S15622 }),
  .C2({ S15925 }),
  .ZN({ S16107 })
);
AOI21_X1 #() 
AOI21_X1_1209_ (
  .A({ S15621 }),
  .B1({ S16107 }),
  .B2({ S16106 }),
  .ZN({ S16108 })
);
OAI211_X1 #() 
OAI211_X1_747_ (
  .A({ S25957[276] }),
  .B({ S16082 }),
  .C1({ S15793 }),
  .C2({ S15795 }),
  .ZN({ S16109 })
);
NAND3_X1 #() 
NAND3_X1_2344_ (
  .A1({ S15531 }),
  .A2({ S15515 }),
  .A3({ S25957[275] }),
  .ZN({ S16110 })
);
OAI211_X1 #() 
OAI211_X1_748_ (
  .A({ S13772 }),
  .B({ S16110 }),
  .C1({ S16025 }),
  .C2({ S15762 }),
  .ZN({ S16111 })
);
NAND3_X1 #() 
NAND3_X1_2345_ (
  .A1({ S16109 }),
  .A2({ S16111 }),
  .A3({ S15621 }),
  .ZN({ S16112 })
);
NAND2_X1 #() 
NAND2_X1_2024_ (
  .A1({ S16112 }),
  .A2({ S25957[278] }),
  .ZN({ S16113 })
);
AOI21_X1 #() 
AOI21_X1_1210_ (
  .A({ S25957[275] }),
  .B1({ S15778 }),
  .B2({ S15520 }),
  .ZN({ S16115 })
);
NOR3_X1 #() 
NOR3_X1_64_ (
  .A1({ S15598 }),
  .A2({ S16115 }),
  .A3({ S25957[276] }),
  .ZN({ S16116 })
);
AOI21_X1 #() 
AOI21_X1_1211_ (
  .A({ S32 }),
  .B1({ S15577 }),
  .B2({ S15533 }),
  .ZN({ S16117 })
);
NAND3_X1 #() 
NAND3_X1_2346_ (
  .A1({ S15747 }),
  .A2({ S15913 }),
  .A3({ S13772 }),
  .ZN({ S16118 })
);
OAI211_X1 #() 
OAI211_X1_749_ (
  .A({ S16118 }),
  .B({ S25957[277] }),
  .C1({ S16117 }),
  .C2({ S15593 }),
  .ZN({ S16119 })
);
OAI211_X1 #() 
OAI211_X1_750_ (
  .A({ S15541 }),
  .B({ S32 }),
  .C1({ S15533 }),
  .C2({ S15527 }),
  .ZN({ S16120 })
);
NAND2_X1 #() 
NAND2_X1_2025_ (
  .A1({ S15645 }),
  .A2({ S16120 }),
  .ZN({ S16121 })
);
OAI21_X1 #() 
OAI21_X1_1129_ (
  .A({ S15621 }),
  .B1({ S16121 }),
  .B2({ S13772 }),
  .ZN({ S16122 })
);
OAI211_X1 #() 
OAI211_X1_751_ (
  .A({ S16119 }),
  .B({ S15585 }),
  .C1({ S16116 }),
  .C2({ S16122 }),
  .ZN({ S16123 })
);
OAI211_X1 #() 
OAI211_X1_752_ (
  .A({ S16123 }),
  .B({ S25957[279] }),
  .C1({ S16108 }),
  .C2({ S16113 }),
  .ZN({ S16124 })
);
NAND3_X1 #() 
NAND3_X1_2347_ (
  .A1({ S15647 }),
  .A2({ S25957[275] }),
  .A3({ S15526 }),
  .ZN({ S16125 })
);
NAND3_X1 #() 
NAND3_X1_2348_ (
  .A1({ S15579 }),
  .A2({ S15600 }),
  .A3({ S15596 }),
  .ZN({ S16126 })
);
AOI21_X1 #() 
AOI21_X1_1212_ (
  .A({ S13772 }),
  .B1({ S16125 }),
  .B2({ S16126 }),
  .ZN({ S16127 })
);
NAND4_X1 #() 
NAND4_X1_289_ (
  .A1({ S15541 }),
  .A2({ S15653 }),
  .A3({ S15531 }),
  .A4({ S32 }),
  .ZN({ S16128 })
);
NAND2_X1 #() 
NAND2_X1_2026_ (
  .A1({ S16128 }),
  .A2({ S16039 }),
  .ZN({ S16129 })
);
OAI21_X1 #() 
OAI21_X1_1130_ (
  .A({ S15621 }),
  .B1({ S16129 }),
  .B2({ S25957[276] }),
  .ZN({ S16130 })
);
OAI21_X1 #() 
OAI21_X1_1131_ (
  .A({ S53 }),
  .B1({ S15515 }),
  .B2({ S25957[274] }),
  .ZN({ S16131 })
);
AND2_X1 #() 
AND2_X1_124_ (
  .A1({ S16131 }),
  .A2({ S25957[275] }),
  .ZN({ S16132 })
);
NAND4_X1 #() 
NAND4_X1_290_ (
  .A1({ S15554 }),
  .A2({ S15542 }),
  .A3({ S15549 }),
  .A4({ S13772 }),
  .ZN({ S16133 })
);
OAI21_X1 #() 
OAI21_X1_1132_ (
  .A({ S25957[276] }),
  .B1({ S16008 }),
  .B2({ S15673 }),
  .ZN({ S16134 })
);
OAI211_X1 #() 
OAI211_X1_753_ (
  .A({ S25957[277] }),
  .B({ S16133 }),
  .C1({ S16132 }),
  .C2({ S16134 }),
  .ZN({ S16136 })
);
OAI211_X1 #() 
OAI211_X1_754_ (
  .A({ S16136 }),
  .B({ S25957[278] }),
  .C1({ S16127 }),
  .C2({ S16130 }),
  .ZN({ S16137 })
);
AOI21_X1 #() 
AOI21_X1_1213_ (
  .A({ S13772 }),
  .B1({ S15966 }),
  .B2({ S15874 }),
  .ZN({ S16138 })
);
OAI21_X1 #() 
OAI21_X1_1133_ (
  .A({ S25957[277] }),
  .B1({ S16138 }),
  .B2({ S15605 }),
  .ZN({ S16139 })
);
INV_X1 #() 
INV_X1_650_ (
  .A({ S15879 }),
  .ZN({ S16140 })
);
NAND2_X1 #() 
NAND2_X1_2027_ (
  .A1({ S15568 }),
  .A2({ S25957[275] }),
  .ZN({ S16141 })
);
NAND3_X1 #() 
NAND3_X1_2349_ (
  .A1({ S16141 }),
  .A2({ S15693 }),
  .A3({ S13772 }),
  .ZN({ S16142 })
);
OAI211_X1 #() 
OAI211_X1_755_ (
  .A({ S15621 }),
  .B({ S16142 }),
  .C1({ S15715 }),
  .C2({ S16140 }),
  .ZN({ S16143 })
);
NAND3_X1 #() 
NAND3_X1_2350_ (
  .A1({ S16143 }),
  .A2({ S16139 }),
  .A3({ S15585 }),
  .ZN({ S16144 })
);
NAND3_X1 #() 
NAND3_X1_2351_ (
  .A1({ S16137 }),
  .A2({ S16144 }),
  .A3({ S15517 }),
  .ZN({ S16145 })
);
NAND3_X1 #() 
NAND3_X1_2352_ (
  .A1({ S16124 }),
  .A2({ S16145 }),
  .A3({ S25957[377] }),
  .ZN({ S16147 })
);
INV_X1 #() 
INV_X1_651_ (
  .A({ S25957[377] }),
  .ZN({ S16148 })
);
AND3_X1 #() 
AND3_X1_93_ (
  .A1({ S16109 }),
  .A2({ S16111 }),
  .A3({ S15621 }),
  .ZN({ S16149 })
);
OAI21_X1 #() 
OAI21_X1_1134_ (
  .A({ S25957[278] }),
  .B1({ S16149 }),
  .B2({ S16108 }),
  .ZN({ S16150 })
);
NAND2_X1 #() 
NAND2_X1_2028_ (
  .A1({ S16121 }),
  .A2({ S25957[276] }),
  .ZN({ S16151 })
);
OAI21_X1 #() 
OAI21_X1_1135_ (
  .A({ S13772 }),
  .B1({ S15598 }),
  .B2({ S16115 }),
  .ZN({ S16152 })
);
NAND3_X1 #() 
NAND3_X1_2353_ (
  .A1({ S16152 }),
  .A2({ S15621 }),
  .A3({ S16151 }),
  .ZN({ S16153 })
);
OAI21_X1 #() 
OAI21_X1_1136_ (
  .A({ S16118 }),
  .B1({ S16117 }),
  .B2({ S15593 }),
  .ZN({ S16154 })
);
NAND2_X1 #() 
NAND2_X1_2029_ (
  .A1({ S16154 }),
  .A2({ S25957[277] }),
  .ZN({ S16155 })
);
NAND3_X1 #() 
NAND3_X1_2354_ (
  .A1({ S16153 }),
  .A2({ S16155 }),
  .A3({ S15585 }),
  .ZN({ S16156 })
);
NAND3_X1 #() 
NAND3_X1_2355_ (
  .A1({ S16150 }),
  .A2({ S16156 }),
  .A3({ S25957[279] }),
  .ZN({ S16158 })
);
AOI22_X1 #() 
AOI22_X1_271_ (
  .A1({ S16131 }),
  .A2({ S25957[275] }),
  .B1({ S15579 }),
  .B2({ S15528 }),
  .ZN({ S16159 })
);
NAND3_X1 #() 
NAND3_X1_2356_ (
  .A1({ S15554 }),
  .A2({ S15549 }),
  .A3({ S15542 }),
  .ZN({ S16160 })
);
NAND2_X1 #() 
NAND2_X1_2030_ (
  .A1({ S16160 }),
  .A2({ S13772 }),
  .ZN({ S16161 })
);
OAI211_X1 #() 
OAI211_X1_756_ (
  .A({ S16161 }),
  .B({ S25957[277] }),
  .C1({ S16159 }),
  .C2({ S13772 }),
  .ZN({ S16162 })
);
NAND2_X1 #() 
NAND2_X1_2031_ (
  .A1({ S16129 }),
  .A2({ S13772 }),
  .ZN({ S16163 })
);
NAND3_X1 #() 
NAND3_X1_2357_ (
  .A1({ S16125 }),
  .A2({ S25957[276] }),
  .A3({ S16126 }),
  .ZN({ S16164 })
);
NAND3_X1 #() 
NAND3_X1_2358_ (
  .A1({ S16164 }),
  .A2({ S16163 }),
  .A3({ S15621 }),
  .ZN({ S16165 })
);
NAND3_X1 #() 
NAND3_X1_2359_ (
  .A1({ S16165 }),
  .A2({ S16162 }),
  .A3({ S25957[278] }),
  .ZN({ S16166 })
);
AND2_X1 #() 
AND2_X1_125_ (
  .A1({ S16141 }),
  .A2({ S15693 }),
  .ZN({ S16167 })
);
OAI211_X1 #() 
OAI211_X1_757_ (
  .A({ S15542 }),
  .B({ S15549 }),
  .C1({ S15600 }),
  .C2({ S25957[275] }),
  .ZN({ S16169 })
);
NAND2_X1 #() 
NAND2_X1_2032_ (
  .A1({ S16169 }),
  .A2({ S25957[276] }),
  .ZN({ S16170 })
);
OAI211_X1 #() 
OAI211_X1_758_ (
  .A({ S15621 }),
  .B({ S16170 }),
  .C1({ S16167 }),
  .C2({ S25957[276] }),
  .ZN({ S16171 })
);
OR3_X1 #() 
OR3_X1_10_ (
  .A1({ S16138 }),
  .A2({ S15605 }),
  .A3({ S15621 }),
  .ZN({ S16172 })
);
NAND3_X1 #() 
NAND3_X1_2360_ (
  .A1({ S16172 }),
  .A2({ S15585 }),
  .A3({ S16171 }),
  .ZN({ S16173 })
);
NAND3_X1 #() 
NAND3_X1_2361_ (
  .A1({ S16173 }),
  .A2({ S16166 }),
  .A3({ S15517 }),
  .ZN({ S16174 })
);
NAND3_X1 #() 
NAND3_X1_2362_ (
  .A1({ S16158 }),
  .A2({ S16174 }),
  .A3({ S16148 }),
  .ZN({ S16175 })
);
AOI21_X1 #() 
AOI21_X1_1214_ (
  .A({ S16103 }),
  .B1({ S16175 }),
  .B2({ S16147 }),
  .ZN({ S16176 })
);
INV_X1 #() 
INV_X1_652_ (
  .A({ S16103 }),
  .ZN({ S25957[441] })
);
NAND3_X1 #() 
NAND3_X1_2363_ (
  .A1({ S16124 }),
  .A2({ S16145 }),
  .A3({ S16148 }),
  .ZN({ S16177 })
);
NAND3_X1 #() 
NAND3_X1_2364_ (
  .A1({ S16158 }),
  .A2({ S16174 }),
  .A3({ S25957[377] }),
  .ZN({ S16179 })
);
AOI21_X1 #() 
AOI21_X1_1215_ (
  .A({ S25957[441] }),
  .B1({ S16179 }),
  .B2({ S16177 }),
  .ZN({ S16180 })
);
OAI21_X1 #() 
OAI21_X1_1137_ (
  .A({ S25957[281] }),
  .B1({ S16176 }),
  .B2({ S16180 }),
  .ZN({ S16181 })
);
NAND3_X1 #() 
NAND3_X1_2365_ (
  .A1({ S16179 }),
  .A2({ S16177 }),
  .A3({ S25957[441] }),
  .ZN({ S16182 })
);
NAND3_X1 #() 
NAND3_X1_2366_ (
  .A1({ S16175 }),
  .A2({ S16147 }),
  .A3({ S16103 }),
  .ZN({ S16183 })
);
NAND3_X1 #() 
NAND3_X1_2367_ (
  .A1({ S16182 }),
  .A2({ S16183 }),
  .A3({ S14841 }),
  .ZN({ S16184 })
);
NAND2_X1 #() 
NAND2_X1_2033_ (
  .A1({ S16181 }),
  .A2({ S16184 }),
  .ZN({ S25957[153] })
);
NAND2_X1 #() 
NAND2_X1_2034_ (
  .A1({ S10498 }),
  .A2({ S10502 }),
  .ZN({ S25957[442] })
);
NAND2_X1 #() 
NAND2_X1_2035_ (
  .A1({ S13369 }),
  .A2({ S13344 }),
  .ZN({ S16185 })
);
XNOR2_X1 #() 
XNOR2_X1_69_ (
  .A({ S16185 }),
  .B({ S25957[602] }),
  .ZN({ S25957[346] })
);
XOR2_X1 #() 
XOR2_X1_32_ (
  .A({ S25957[346] }),
  .B({ S25957[442] }),
  .Z({ S25957[314] })
);
INV_X1 #() 
INV_X1_653_ (
  .A({ S25957[314] }),
  .ZN({ S16187 })
);
NAND2_X1 #() 
NAND2_X1_2036_ (
  .A1({ S7549 }),
  .A2({ S7527 }),
  .ZN({ S25957[634] })
);
NAND2_X1 #() 
NAND2_X1_2037_ (
  .A1({ S10480 }),
  .A2({ S10496 }),
  .ZN({ S16188 })
);
XNOR2_X1 #() 
XNOR2_X1_70_ (
  .A({ S16188 }),
  .B({ S25957[634] }),
  .ZN({ S25957[506] })
);
XNOR2_X1 #() 
XNOR2_X1_71_ (
  .A({ S16185 }),
  .B({ S25957[506] }),
  .ZN({ S25957[378] })
);
NAND3_X1 #() 
NAND3_X1_2368_ (
  .A1({ S15554 }),
  .A2({ S25957[275] }),
  .A3({ S15549 }),
  .ZN({ S16189 })
);
NAND3_X1 #() 
NAND3_X1_2369_ (
  .A1({ S15965 }),
  .A2({ S25957[276] }),
  .A3({ S16189 }),
  .ZN({ S16190 })
);
NAND3_X1 #() 
NAND3_X1_2370_ (
  .A1({ S15611 }),
  .A2({ S15706 }),
  .A3({ S25957[275] }),
  .ZN({ S16191 })
);
AOI21_X1 #() 
AOI21_X1_1216_ (
  .A({ S25957[276] }),
  .B1({ S15561 }),
  .B2({ S15703 }),
  .ZN({ S16192 })
);
AOI21_X1 #() 
AOI21_X1_1217_ (
  .A({ S15621 }),
  .B1({ S16191 }),
  .B2({ S16192 }),
  .ZN({ S16194 })
);
NAND2_X1 #() 
NAND2_X1_2038_ (
  .A1({ S16190 }),
  .A2({ S16194 }),
  .ZN({ S16195 })
);
AND3_X1 #() 
AND3_X1_94_ (
  .A1({ S15663 }),
  .A2({ S13772 }),
  .A3({ S16043 }),
  .ZN({ S16196 })
);
NAND3_X1 #() 
NAND3_X1_2371_ (
  .A1({ S15653 }),
  .A2({ S25957[275] }),
  .A3({ S25957[273] }),
  .ZN({ S16197 })
);
NAND2_X1 #() 
NAND2_X1_2039_ (
  .A1({ S16197 }),
  .A2({ S25957[276] }),
  .ZN({ S16198 })
);
OAI21_X1 #() 
OAI21_X1_1138_ (
  .A({ S15621 }),
  .B1({ S15856 }),
  .B2({ S16198 }),
  .ZN({ S16199 })
);
OAI21_X1 #() 
OAI21_X1_1139_ (
  .A({ S16195 }),
  .B1({ S16196 }),
  .B2({ S16199 }),
  .ZN({ S16200 })
);
AOI21_X1 #() 
AOI21_X1_1218_ (
  .A({ S15608 }),
  .B1({ S15541 }),
  .B2({ S15600 }),
  .ZN({ S16201 })
);
NAND3_X1 #() 
NAND3_X1_2372_ (
  .A1({ S15778 }),
  .A2({ S25957[275] }),
  .A3({ S15531 }),
  .ZN({ S16202 })
);
NAND2_X1 #() 
NAND2_X1_2040_ (
  .A1({ S16202 }),
  .A2({ S25957[276] }),
  .ZN({ S16203 })
);
OAI211_X1 #() 
OAI211_X1_759_ (
  .A({ S13772 }),
  .B({ S16197 }),
  .C1({ S15879 }),
  .C2({ S52 }),
  .ZN({ S16205 })
);
OAI211_X1 #() 
OAI211_X1_760_ (
  .A({ S15621 }),
  .B({ S16205 }),
  .C1({ S16203 }),
  .C2({ S16201 }),
  .ZN({ S16206 })
);
OAI211_X1 #() 
OAI211_X1_761_ (
  .A({ S15578 }),
  .B({ S13772 }),
  .C1({ S15644 }),
  .C2({ S15608 }),
  .ZN({ S16207 })
);
NAND2_X1 #() 
NAND2_X1_2041_ (
  .A1({ S25957[276] }),
  .A2({ S15567 }),
  .ZN({ S16208 })
);
OAI211_X1 #() 
OAI211_X1_762_ (
  .A({ S25957[277] }),
  .B({ S15919 }),
  .C1({ S15932 }),
  .C2({ S16208 }),
  .ZN({ S16209 })
);
INV_X1 #() 
INV_X1_654_ (
  .A({ S16209 }),
  .ZN({ S16210 })
);
AOI21_X1 #() 
AOI21_X1_1219_ (
  .A({ S15585 }),
  .B1({ S16207 }),
  .B2({ S16210 }),
  .ZN({ S16211 })
);
AOI22_X1 #() 
AOI22_X1_272_ (
  .A1({ S16200 }),
  .A2({ S15585 }),
  .B1({ S16211 }),
  .B2({ S16206 }),
  .ZN({ S16212 })
);
OAI21_X1 #() 
OAI21_X1_1140_ (
  .A({ S32 }),
  .B1({ S15570 }),
  .B2({ S15552 }),
  .ZN({ S16213 })
);
NAND3_X1 #() 
NAND3_X1_2373_ (
  .A1({ S16213 }),
  .A2({ S25957[276] }),
  .A3({ S15603 }),
  .ZN({ S16214 })
);
NAND3_X1 #() 
NAND3_X1_2374_ (
  .A1({ S15576 }),
  .A2({ S25957[275] }),
  .A3({ S15740 }),
  .ZN({ S16216 })
);
AOI21_X1 #() 
AOI21_X1_1220_ (
  .A({ S15621 }),
  .B1({ S16216 }),
  .B2({ S15788 }),
  .ZN({ S16217 })
);
NAND2_X1 #() 
NAND2_X1_2042_ (
  .A1({ S16214 }),
  .A2({ S16217 }),
  .ZN({ S16218 })
);
NAND2_X1 #() 
NAND2_X1_2043_ (
  .A1({ S15766 }),
  .A2({ S25957[276] }),
  .ZN({ S16219 })
);
NOR3_X1 #() 
NOR3_X1_65_ (
  .A1({ S15572 }),
  .A2({ S15570 }),
  .A3({ S32 }),
  .ZN({ S16220 })
);
NAND3_X1 #() 
NAND3_X1_2375_ (
  .A1({ S15666 }),
  .A2({ S13772 }),
  .A3({ S15615 }),
  .ZN({ S16221 })
);
OAI211_X1 #() 
OAI211_X1_763_ (
  .A({ S15621 }),
  .B({ S16221 }),
  .C1({ S16220 }),
  .C2({ S16219 }),
  .ZN({ S16222 })
);
NAND3_X1 #() 
NAND3_X1_2376_ (
  .A1({ S16222 }),
  .A2({ S16218 }),
  .A3({ S25957[278] }),
  .ZN({ S16223 })
);
NAND3_X1 #() 
NAND3_X1_2377_ (
  .A1({ S15649 }),
  .A2({ S25957[275] }),
  .A3({ S15539 }),
  .ZN({ S16224 })
);
AOI21_X1 #() 
AOI21_X1_1221_ (
  .A({ S25957[276] }),
  .B1({ S16224 }),
  .B2({ S15829 }),
  .ZN({ S16225 })
);
NAND3_X1 #() 
NAND3_X1_2378_ (
  .A1({ S15567 }),
  .A2({ S25957[275] }),
  .A3({ S25957[272] }),
  .ZN({ S16227 })
);
AOI21_X1 #() 
AOI21_X1_1222_ (
  .A({ S13772 }),
  .B1({ S15693 }),
  .B2({ S16227 }),
  .ZN({ S16228 })
);
OAI21_X1 #() 
OAI21_X1_1141_ (
  .A({ S25957[277] }),
  .B1({ S16225 }),
  .B2({ S16228 }),
  .ZN({ S16229 })
);
OAI211_X1 #() 
OAI211_X1_764_ (
  .A({ S16197 }),
  .B({ S25957[276] }),
  .C1({ S15644 }),
  .C2({ S25957[275] }),
  .ZN({ S16230 })
);
AOI21_X1 #() 
AOI21_X1_1223_ (
  .A({ S25957[277] }),
  .B1({ S16192 }),
  .B2({ S15700 }),
  .ZN({ S16231 })
);
AOI21_X1 #() 
AOI21_X1_1224_ (
  .A({ S25957[278] }),
  .B1({ S16231 }),
  .B2({ S16230 }),
  .ZN({ S16232 })
);
AOI21_X1 #() 
AOI21_X1_1225_ (
  .A({ S15517 }),
  .B1({ S16229 }),
  .B2({ S16232 }),
  .ZN({ S16233 })
);
NAND2_X1 #() 
NAND2_X1_2044_ (
  .A1({ S16233 }),
  .A2({ S16223 }),
  .ZN({ S16234 })
);
OAI211_X1 #() 
OAI211_X1_765_ (
  .A({ S16234 }),
  .B({ S25957[378] }),
  .C1({ S16212 }),
  .C2({ S25957[279] }),
  .ZN({ S16235 })
);
INV_X1 #() 
INV_X1_655_ (
  .A({ S25957[378] }),
  .ZN({ S16236 })
);
NAND2_X1 #() 
NAND2_X1_2045_ (
  .A1({ S16200 }),
  .A2({ S15585 }),
  .ZN({ S16238 })
);
NAND2_X1 #() 
NAND2_X1_2046_ (
  .A1({ S16211 }),
  .A2({ S16206 }),
  .ZN({ S16239 })
);
AOI21_X1 #() 
AOI21_X1_1226_ (
  .A({ S25957[279] }),
  .B1({ S16238 }),
  .B2({ S16239 }),
  .ZN({ S16240 })
);
AND2_X1 #() 
AND2_X1_126_ (
  .A1({ S16233 }),
  .A2({ S16223 }),
  .ZN({ S16241 })
);
OAI21_X1 #() 
OAI21_X1_1142_ (
  .A({ S16236 }),
  .B1({ S16240 }),
  .B2({ S16241 }),
  .ZN({ S16242 })
);
NAND3_X1 #() 
NAND3_X1_2379_ (
  .A1({ S16242 }),
  .A2({ S25957[346] }),
  .A3({ S16235 }),
  .ZN({ S16243 })
);
INV_X1 #() 
INV_X1_656_ (
  .A({ S25957[346] }),
  .ZN({ S16244 })
);
OAI211_X1 #() 
OAI211_X1_766_ (
  .A({ S16234 }),
  .B({ S16236 }),
  .C1({ S16212 }),
  .C2({ S25957[279] }),
  .ZN({ S16245 })
);
OAI21_X1 #() 
OAI21_X1_1143_ (
  .A({ S25957[378] }),
  .B1({ S16240 }),
  .B2({ S16241 }),
  .ZN({ S16246 })
);
NAND3_X1 #() 
NAND3_X1_2380_ (
  .A1({ S16246 }),
  .A2({ S16244 }),
  .A3({ S16245 }),
  .ZN({ S16247 })
);
NAND3_X1 #() 
NAND3_X1_2381_ (
  .A1({ S16243 }),
  .A2({ S16247 }),
  .A3({ S16187 }),
  .ZN({ S16249 })
);
NAND3_X1 #() 
NAND3_X1_2382_ (
  .A1({ S16242 }),
  .A2({ S16244 }),
  .A3({ S16235 }),
  .ZN({ S16250 })
);
NAND3_X1 #() 
NAND3_X1_2383_ (
  .A1({ S16246 }),
  .A2({ S25957[346] }),
  .A3({ S16245 }),
  .ZN({ S16251 })
);
NAND3_X1 #() 
NAND3_X1_2384_ (
  .A1({ S16250 }),
  .A2({ S16251 }),
  .A3({ S25957[314] }),
  .ZN({ S16252 })
);
NAND3_X1 #() 
NAND3_X1_2385_ (
  .A1({ S16249 }),
  .A2({ S16252 }),
  .A3({ S25957[282] }),
  .ZN({ S16253 })
);
NAND3_X1 #() 
NAND3_X1_2386_ (
  .A1({ S16243 }),
  .A2({ S16247 }),
  .A3({ S25957[314] }),
  .ZN({ S16254 })
);
NAND3_X1 #() 
NAND3_X1_2387_ (
  .A1({ S16250 }),
  .A2({ S16251 }),
  .A3({ S16187 }),
  .ZN({ S16255 })
);
NAND3_X1 #() 
NAND3_X1_2388_ (
  .A1({ S16254 }),
  .A2({ S16255 }),
  .A3({ S14834 }),
  .ZN({ S16256 })
);
NAND2_X1 #() 
NAND2_X1_2047_ (
  .A1({ S16253 }),
  .A2({ S16256 }),
  .ZN({ S25957[154] })
);
NAND2_X1 #() 
NAND2_X1_2048_ (
  .A1({ S17944 }),
  .A2({ S17976 }),
  .ZN({ S25957[1194] })
);
NAND2_X1 #() 
NAND2_X1_2049_ (
  .A1({ S11432 }),
  .A2({ S11465 }),
  .ZN({ S25957[1202] })
);
NOR2_X1 #() 
NOR2_X1_466_ (
  .A1({ S20066 }),
  .A2({ S20067 }),
  .ZN({ S25957[1209] })
);
NAND2_X1 #() 
NAND2_X1_2050_ (
  .A1({ S22638 }),
  .A2({ S22639 }),
  .ZN({ S25957[1098] })
);
NAND2_X1 #() 
NAND2_X1_2051_ (
  .A1({ S21178 }),
  .A2({ S21179 }),
  .ZN({ S25957[1099] })
);
XNOR2_X1 #() 
XNOR2_X1_72_ (
  .A({ S25957[1138] }),
  .B({ S23272 }),
  .ZN({ S25957[1106] })
);
NOR2_X1 #() 
NOR2_X1_467_ (
  .A1({ S20469 }),
  .A2({ S20470 }),
  .ZN({ S25957[1108] })
);
INV_X1 #() 
INV_X1_657_ (
  .A({ S22837 }),
  .ZN({ S25957[1109] })
);
NAND2_X1 #() 
NAND2_X1_2052_ (
  .A1({ S24018 }),
  .A2({ S24019 }),
  .ZN({ S25957[1113] })
);
NOR2_X1 #() 
NOR2_X1_468_ (
  .A1({ S22620 }),
  .A2({ S22619 }),
  .ZN({ S25957[1082] })
);
NOR2_X1 #() 
NOR2_X1_469_ (
  .A1({ S24542 }),
  .A2({ S24543 }),
  .ZN({ S25957[960] })
);
NAND2_X1 #() 
NAND2_X1_2053_ (
  .A1({ S24281 }),
  .A2({ S24289 }),
  .ZN({ S25957[965] })
);
INV_X1 #() 
INV_X1_658_ (
  .A({ S23623 }),
  .ZN({ S25957[973] })
);
NAND2_X1 #() 
NAND2_X1_2054_ (
  .A1({ S23202 }),
  .A2({ S23201 }),
  .ZN({ S25957[976] })
);
NOR2_X1 #() 
NOR2_X1_470_ (
  .A1({ S23239 }),
  .A2({ S23240 }),
  .ZN({ S25957[977] })
);
NOR2_X1 #() 
NOR2_X1_471_ (
  .A1({ S22752 }),
  .A2({ S22750 }),
  .ZN({ S25957[983] })
);
NAND2_X1 #() 
NAND2_X1_2055_ (
  .A1({ S25261 }),
  .A2({ S25260 }),
  .ZN({ S25957[984] })
);
NOR2_X1 #() 
NOR2_X1_472_ (
  .A1({ S25173 }),
  .A2({ S25174 }),
  .ZN({ S25957[987] })
);
NOR2_X1 #() 
NOR2_X1_473_ (
  .A1({ S25060 }),
  .A2({ S25061 }),
  .ZN({ S25957[988] })
);
XNOR2_X1 #() 
XNOR2_X1_73_ (
  .A({ S25957[962] }),
  .B({ S1614 }),
  .ZN({ S25957[930] })
);
XNOR2_X1 #() 
XNOR2_X1_74_ (
  .A({ S25957[966] }),
  .B({ S1215 }),
  .ZN({ S25957[934] })
);
NAND2_X1 #() 
NAND2_X1_2056_ (
  .A1({ S24009 }),
  .A2({ S24006 }),
  .ZN({ S25957[938] })
);
NAND2_X1 #() 
NAND2_X1_2057_ (
  .A1({ S23789 }),
  .A2({ S23793 }),
  .ZN({ S25957[939] })
);
XNOR2_X1 #() 
XNOR2_X1_75_ (
  .A({ S25957[978] }),
  .B({ S268 }),
  .ZN({ S25957[946] })
);
INV_X1 #() 
INV_X1_659_ (
  .A({ S2445 }),
  .ZN({ S25957[949] })
);
NOR2_X1 #() 
NOR2_X1_474_ (
  .A1({ S1549 }),
  .A2({ S1550 }),
  .ZN({ S25957[833] })
);
INV_X1 #() 
INV_X1_660_ (
  .A({ S25957[972] }),
  .ZN({ S16260 })
);
XNOR2_X1 #() 
XNOR2_X1_76_ (
  .A({ S25957[876] }),
  .B({ S16260 }),
  .ZN({ S25957[844] })
);
NAND2_X1 #() 
NAND2_X1_2058_ (
  .A1({ S548 }),
  .A2({ S551 }),
  .ZN({ S25957[846] })
);
XNOR2_X1 #() 
XNOR2_X1_77_ (
  .A({ S25957[882] }),
  .B({ S2866 }),
  .ZN({ S25957[850] })
);
NAND2_X1 #() 
NAND2_X1_2059_ (
  .A1({ S2224 }),
  .A2({ S2225 }),
  .ZN({ S25957[858] })
);
NOR2_X1 #() 
NOR2_X1_475_ (
  .A1({ S25667 }),
  .A2({ S25668 }),
  .ZN({ S25957[821] })
);
XNOR2_X1 #() 
XNOR2_X1_78_ (
  .A({ S25957[859] }),
  .B({ S4503 }),
  .ZN({ S25957[827] })
);
XNOR2_X1 #() 
XNOR2_X1_79_ (
  .A({ S1804 }),
  .B({ S25957[958] }),
  .ZN({ S25957[830] })
);
INV_X1 #() 
INV_X1_661_ (
  .A({ S9041 }),
  .ZN({ S25957[711] })
);
NOR2_X1 #() 
NOR2_X1_476_ (
  .A1({ S3472 }),
  .A2({ S3460 }),
  .ZN({ S16262 })
);
INV_X1 #() 
INV_X1_662_ (
  .A({ S16262 }),
  .ZN({ S25957[714] })
);
NOR2_X1 #() 
NOR2_X1_477_ (
  .A1({ S2659 }),
  .A2({ S2660 }),
  .ZN({ S25957[723] })
);
XNOR2_X1 #() 
XNOR2_X1_80_ (
  .A({ S25957[757] }),
  .B({ S4996 }),
  .ZN({ S25957[725] })
);
XOR2_X1 #() 
XOR2_X1_33_ (
  .A({ S25957[763] }),
  .B({ S25957[859] }),
  .Z({ S25957[731] })
);
INV_X1 #() 
INV_X1_663_ (
  .A({ S10093 }),
  .ZN({ S25957[732] })
);
XNOR2_X1 #() 
XNOR2_X1_81_ (
  .A({ S25957[766] }),
  .B({ S1804 }),
  .ZN({ S25957[734] })
);
NAND2_X1 #() 
NAND2_X1_2060_ (
  .A1({ S3352 }),
  .A2({ S3353 }),
  .ZN({ S25957[680] })
);
NAND2_X1 #() 
NAND2_X1_2061_ (
  .A1({ S3406 }),
  .A2({ S3403 }),
  .ZN({ S25957[681] })
);
NAND2_X1 #() 
NAND2_X1_2062_ (
  .A1({ S2742 }),
  .A2({ S2745 }),
  .ZN({ S25957[688] })
);
XNOR2_X1 #() 
XNOR2_X1_82_ (
  .A({ S8203 }),
  .B({ S25957[818] }),
  .ZN({ S25957[690] })
);
NOR2_X1 #() 
NOR2_X1_478_ (
  .A1({ S4672 }),
  .A2({ S4675 }),
  .ZN({ S25957[696] })
);
NAND2_X1 #() 
NAND2_X1_2063_ (
  .A1({ S4729 }),
  .A2({ S4733 }),
  .ZN({ S25957[697] })
);
NAND2_X1 #() 
NAND2_X1_2064_ (
  .A1({ S6710 }),
  .A2({ S6747 }),
  .ZN({ S25957[576] })
);
NAND2_X1 #() 
NAND2_X1_2065_ (
  .A1({ S6823 }),
  .A2({ S6824 }),
  .ZN({ S25957[577] })
);
NOR2_X1 #() 
NOR2_X1_479_ (
  .A1({ S6886 }),
  .A2({ S6885 }),
  .ZN({ S25957[578] })
);
NAND2_X1 #() 
NAND2_X1_2066_ (
  .A1({ S6495 }),
  .A2({ S6498 }),
  .ZN({ S25957[581] })
);
XNOR2_X1 #() 
XNOR2_X1_83_ (
  .A({ S25957[616] }),
  .B({ S8811 }),
  .ZN({ S25957[584] })
);
XOR2_X1 #() 
XOR2_X1_34_ (
  .A({ S25957[623] }),
  .B({ S25957[719] }),
  .Z({ S25957[591] })
);
NAND2_X1 #() 
NAND2_X1_2067_ (
  .A1({ S8275 }),
  .A2({ S8276 }),
  .ZN({ S25957[594] })
);
NAND2_X1 #() 
NAND2_X1_2068_ (
  .A1({ S7264 }),
  .A2({ S7262 }),
  .ZN({ S25957[604] })
);
XNOR2_X1 #() 
XNOR2_X1_84_ (
  .A({ S25957[582] }),
  .B({ S9185 }),
  .ZN({ S25957[550] })
);
NAND2_X1 #() 
NAND2_X1_2069_ (
  .A1({ S6097 }),
  .A2({ S6098 }),
  .ZN({ S25957[553] })
);
XNOR2_X1 #() 
XNOR2_X1_85_ (
  .A({ S25957[587] }),
  .B({ S8685 }),
  .ZN({ S25957[555] })
);
NAND2_X1 #() 
NAND2_X1_2070_ (
  .A1({ S5742 }),
  .A2({ S5743 }),
  .ZN({ S25957[557] })
);
NAND2_X1 #() 
NAND2_X1_2071_ (
  .A1({ S5350 }),
  .A2({ S5353 }),
  .ZN({ S25957[561] })
);
XNOR2_X1 #() 
XNOR2_X1_86_ (
  .A({ S25957[603] }),
  .B({ S10241 }),
  .ZN({ S25957[571] })
);
NAND2_X1 #() 
NAND2_X1_2072_ (
  .A1({ S9521 }),
  .A2({ S9522 }),
  .ZN({ S25957[483] })
);
XNOR2_X1 #() 
XNOR2_X1_87_ (
  .A({ S8126 }),
  .B({ S25957[624] }),
  .ZN({ S25957[496] })
);
NAND2_X1 #() 
NAND2_X1_2073_ (
  .A1({ S8939 }),
  .A2({ S8940 }),
  .ZN({ S25957[457] })
);
NOR2_X1 #() 
NOR2_X1_480_ (
  .A1({ S8677 }),
  .A2({ S8678 }),
  .ZN({ S25957[460] })
);
XNOR2_X1 #() 
XNOR2_X1_88_ (
  .A({ S25957[493] }),
  .B({ S11576 }),
  .ZN({ S25957[461] })
);
XOR2_X1 #() 
XOR2_X1_35_ (
  .A({ S8417 }),
  .B({ S25957[719] }),
  .Z({ S25957[463] })
);
NOR2_X1 #() 
NOR2_X1_481_ (
  .A1({ S7699 }),
  .A2({ S7700 }),
  .ZN({ S25957[471] })
);
NOR2_X1 #() 
NOR2_X1_482_ (
  .A1({ S10339 }),
  .A2({ S10340 }),
  .ZN({ S16266 })
);
INV_X1 #() 
INV_X1_664_ (
  .A({ S16266 }),
  .ZN({ S25957[472] })
);
NOR2_X1 #() 
NOR2_X1_483_ (
  .A1({ S10396 }),
  .A2({ S10395 }),
  .ZN({ S25957[473] })
);
NOR2_X1 #() 
NOR2_X1_484_ (
  .A1({ S10459 }),
  .A2({ S10497 }),
  .ZN({ S25957[474] })
);
XOR2_X1 #() 
XOR2_X1_36_ (
  .A({ S25957[507] }),
  .B({ S25957[603] }),
  .Z({ S25957[475] })
);
NAND2_X1 #() 
NAND2_X1_2074_ (
  .A1({ S10152 }),
  .A2({ S10149 }),
  .ZN({ S25957[476] })
);
NAND2_X1 #() 
NAND2_X1_2075_ (
  .A1({ S10001 }),
  .A2({ S10002 }),
  .ZN({ S25957[478] })
);
NAND2_X1 #() 
NAND2_X1_2076_ (
  .A1({ S9267 }),
  .A2({ S9268 }),
  .ZN({ S25957[422] })
);
XOR2_X1 #() 
XOR2_X1_37_ (
  .A({ S25957[457] }),
  .B({ S25957[553] }),
  .Z({ S25957[425] })
);
NOR2_X1 #() 
NOR2_X1_485_ (
  .A1({ S8273 }),
  .A2({ S8272 }),
  .ZN({ S25957[434] })
);
NOR2_X1 #() 
NOR2_X1_486_ (
  .A1({ S8059 }),
  .A2({ S8063 }),
  .ZN({ S25957[435] })
);
XNOR2_X1 #() 
XNOR2_X1_89_ (
  .A({ S13616 }),
  .B({ S25957[565] }),
  .ZN({ S25957[437] })
);
NOR2_X1 #() 
NOR2_X1_487_ (
  .A1({ S10341 }),
  .A2({ S10337 }),
  .ZN({ S25957[440] })
);
NAND2_X1 #() 
NAND2_X1_2077_ (
  .A1({ S10247 }),
  .A2({ S10248 }),
  .ZN({ S25957[443] })
);
XNOR2_X1 #() 
XNOR2_X1_90_ (
  .A({ S25957[477] }),
  .B({ S12888 }),
  .ZN({ S25957[445] })
);
NAND2_X1 #() 
NAND2_X1_2078_ (
  .A1({ S9907 }),
  .A2({ S9908 }),
  .ZN({ S25957[447] })
);
NAND2_X1 #() 
NAND2_X1_2079_ (
  .A1({ S12505 }),
  .A2({ S12506 }),
  .ZN({ S25957[352] })
);
NAND2_X1 #() 
NAND2_X1_2080_ (
  .A1({ S12571 }),
  .A2({ S12572 }),
  .ZN({ S25957[353] })
);
NAND2_X1 #() 
NAND2_X1_2081_ (
  .A1({ S12664 }),
  .A2({ S12663 }),
  .ZN({ S25957[354] })
);
NAND2_X1 #() 
NAND2_X1_2082_ (
  .A1({ S12392 }),
  .A2({ S12416 }),
  .ZN({ S16269 })
);
XNOR2_X1 #() 
XNOR2_X1_91_ (
  .A({ S16269 }),
  .B({ S25957[483] }),
  .ZN({ S25957[355] })
);
XOR2_X1 #() 
XOR2_X1_38_ (
  .A({ S11726 }),
  .B({ S25957[491] }),
  .Z({ S25957[363] })
);
NAND2_X1 #() 
NAND2_X1_2083_ (
  .A1({ S11492 }),
  .A2({ S11493 }),
  .ZN({ S25957[366] })
);
NAND2_X1 #() 
NAND2_X1_2084_ (
  .A1({ S11071 }),
  .A2({ S11054 }),
  .ZN({ S16271 })
);
XNOR2_X1 #() 
XNOR2_X1_92_ (
  .A({ S16271 }),
  .B({ S25957[496] }),
  .ZN({ S25957[368] })
);
NAND2_X1 #() 
NAND2_X1_2085_ (
  .A1({ S11127 }),
  .A2({ S11108 }),
  .ZN({ S16272 })
);
XNOR2_X1 #() 
XNOR2_X1_93_ (
  .A({ S16272 }),
  .B({ S25957[497] }),
  .ZN({ S25957[369] })
);
NAND2_X1 #() 
NAND2_X1_2086_ (
  .A1({ S11272 }),
  .A2({ S11236 }),
  .ZN({ S25957[370] })
);
NAND2_X1 #() 
NAND2_X1_2087_ (
  .A1({ S12510 }),
  .A2({ S12511 }),
  .ZN({ S25957[320] })
);
INV_X1 #() 
INV_X1_665_ (
  .A({ S15394 }),
  .ZN({ S25957[321] })
);
NAND2_X1 #() 
NAND2_X1_2088_ (
  .A1({ S12669 }),
  .A2({ S12670 }),
  .ZN({ S25957[322] })
);
NAND2_X1 #() 
NAND2_X1_2089_ (
  .A1({ S12417 }),
  .A2({ S12436 }),
  .ZN({ S25957[323] })
);
INV_X1 #() 
INV_X1_666_ (
  .A({ S12198 }),
  .ZN({ S25957[326] })
);
NAND2_X1 #() 
NAND2_X1_2090_ (
  .A1({ S12111 }),
  .A2({ S12113 }),
  .ZN({ S16274 })
);
INV_X1 #() 
INV_X1_667_ (
  .A({ S16274 }),
  .ZN({ S25957[327] })
);
XNOR2_X1 #() 
XNOR2_X1_94_ (
  .A({ S14744 }),
  .B({ S25957[458] }),
  .ZN({ S25957[330] })
);
NOR2_X1 #() 
NOR2_X1_488_ (
  .A1({ S11721 }),
  .A2({ S11722 }),
  .ZN({ S25957[331] })
);
NAND2_X1 #() 
NAND2_X1_2091_ (
  .A1({ S11497 }),
  .A2({ S11499 }),
  .ZN({ S25957[334] })
);
XOR2_X1 #() 
XOR2_X1_39_ (
  .A({ S11409 }),
  .B({ S25957[591] }),
  .Z({ S25957[335] })
);
NOR2_X1 #() 
NOR2_X1_489_ (
  .A1({ S11041 }),
  .A2({ S11073 }),
  .ZN({ S16275 })
);
INV_X1 #() 
INV_X1_668_ (
  .A({ S16275 }),
  .ZN({ S25957[336] })
);
NAND2_X1 #() 
NAND2_X1_2092_ (
  .A1({ S11173 }),
  .A2({ S11128 }),
  .ZN({ S25957[337] })
);
XNOR2_X1 #() 
XNOR2_X1_95_ (
  .A({ S25957[370] }),
  .B({ S14119 }),
  .ZN({ S25957[338] })
);
XNOR2_X1 #() 
XNOR2_X1_96_ (
  .A({ S25957[373] }),
  .B({ S13616 }),
  .ZN({ S25957[341] })
);
INV_X1 #() 
INV_X1_669_ (
  .A({ S10726 }),
  .ZN({ S25957[342] })
);
NOR2_X1 #() 
NOR2_X1_490_ (
  .A1({ S13294 }),
  .A2({ S13317 }),
  .ZN({ S25957[345] })
);
XOR2_X1 #() 
XOR2_X1_40_ (
  .A({ S25957[380] }),
  .B({ S25957[476] }),
  .Z({ S25957[348] })
);
XNOR2_X1 #() 
XNOR2_X1_97_ (
  .A({ S12877 }),
  .B({ S9995 }),
  .ZN({ S25957[350] })
);
XNOR2_X1 #() 
XNOR2_X1_98_ (
  .A({ S25957[383] }),
  .B({ S9904 }),
  .ZN({ S25957[351] })
);
NAND2_X1 #() 
NAND2_X1_2093_ (
  .A1({ S12515 }),
  .A2({ S12516 }),
  .ZN({ S25957[288] })
);
NAND2_X1 #() 
NAND2_X1_2094_ (
  .A1({ S12673 }),
  .A2({ S12674 }),
  .ZN({ S25957[290] })
);
XNOR2_X1 #() 
XNOR2_X1_99_ (
  .A({ S12198 }),
  .B({ S25957[422] }),
  .ZN({ S25957[294] })
);
XOR2_X1 #() 
XOR2_X1_41_ (
  .A({ S25957[329] }),
  .B({ S25957[425] }),
  .Z({ S25957[297] })
);
NOR2_X1 #() 
NOR2_X1_491_ (
  .A1({ S11966 }),
  .A2({ S11969 }),
  .ZN({ S25957[298] })
);
NAND2_X1 #() 
NAND2_X1_2095_ (
  .A1({ S11732 }),
  .A2({ S11731 }),
  .ZN({ S16278 })
);
INV_X1 #() 
INV_X1_670_ (
  .A({ S16278 }),
  .ZN({ S25957[299] })
);
NOR2_X1 #() 
NOR2_X1_492_ (
  .A1({ S11584 }),
  .A2({ S11582 }),
  .ZN({ S25957[301] })
);
NAND2_X1 #() 
NAND2_X1_2096_ (
  .A1({ S11502 }),
  .A2({ S11503 }),
  .ZN({ S25957[302] })
);
NAND2_X1 #() 
NAND2_X1_2097_ (
  .A1({ S11082 }),
  .A2({ S11084 }),
  .ZN({ S16279 })
);
INV_X1 #() 
INV_X1_671_ (
  .A({ S16279 }),
  .ZN({ S25957[304] })
);
NOR2_X1 #() 
NOR2_X1_493_ (
  .A1({ S11175 }),
  .A2({ S11174 }),
  .ZN({ S25957[305] })
);
NOR2_X1 #() 
NOR2_X1_494_ (
  .A1({ S11273 }),
  .A2({ S11277 }),
  .ZN({ S25957[306] })
);
NAND2_X1 #() 
NAND2_X1_2098_ (
  .A1({ S10804 }),
  .A2({ S10805 }),
  .ZN({ S25957[309] })
);
XNOR2_X1 #() 
XNOR2_X1_100_ (
  .A({ S10726 }),
  .B({ S25957[438] }),
  .ZN({ S25957[310] })
);
INV_X1 #() 
INV_X1_672_ (
  .A({ S10651 }),
  .ZN({ S25957[311] })
);
XOR2_X1 #() 
XOR2_X1_42_ (
  .A({ S25957[344] }),
  .B({ S25957[440] }),
  .Z({ S25957[312] })
);
XNOR2_X1 #() 
XNOR2_X1_101_ (
  .A({ S25957[345] }),
  .B({ S16103 }),
  .ZN({ S25957[313] })
);
XNOR2_X1 #() 
XNOR2_X1_102_ (
  .A({ S15910 }),
  .B({ S25957[443] }),
  .ZN({ S25957[315] })
);
NOR2_X1 #() 
NOR2_X1_495_ (
  .A1({ S12881 }),
  .A2({ S12882 }),
  .ZN({ S25957[318] })
);
NAND4_X1 #() 
NAND4_X1_291_ (
  .A1({ S15355 }),
  .A2({ S15327 }),
  .A3({ S12506 }),
  .A4({ S12505 }),
  .ZN({ S16281 })
);
NAND3_X1 #() 
NAND3_X1_2389_ (
  .A1({ S15373 }),
  .A2({ S15392 }),
  .A3({ S25957[352] }),
  .ZN({ S16282 })
);
NAND2_X1 #() 
NAND2_X1_2099_ (
  .A1({ S16281 }),
  .A2({ S16282 }),
  .ZN({ S25957[224] })
);
XNOR2_X1 #() 
XNOR2_X1_103_ (
  .A({ S15440 }),
  .B({ S25957[353] }),
  .ZN({ S25957[225] })
);
XNOR2_X1 #() 
XNOR2_X1_104_ (
  .A({ S15508 }),
  .B({ S25957[354] }),
  .ZN({ S25957[226] })
);
NAND2_X1 #() 
NAND2_X1_2100_ (
  .A1({ S15279 }),
  .A2({ S15248 }),
  .ZN({ S16284 })
);
XNOR2_X1 #() 
XNOR2_X1_105_ (
  .A({ S16284 }),
  .B({ S25957[355] }),
  .ZN({ S25957[227] })
);
NAND2_X1 #() 
NAND2_X1_2101_ (
  .A1({ S15208 }),
  .A2({ S15196 }),
  .ZN({ S25957[228] })
);
NAND2_X1 #() 
NAND2_X1_2102_ (
  .A1({ S15120 }),
  .A2({ S15111 }),
  .ZN({ S16285 })
);
INV_X1 #() 
INV_X1_673_ (
  .A({ S16285 }),
  .ZN({ S25957[229] })
);
XNOR2_X1 #() 
XNOR2_X1_106_ (
  .A({ S15036 }),
  .B({ S25957[358] }),
  .ZN({ S25957[230] })
);
NAND2_X1 #() 
NAND2_X1_2103_ (
  .A1({ S14953 }),
  .A2({ S14903 }),
  .ZN({ S16286 })
);
NAND2_X1 #() 
NAND2_X1_2104_ (
  .A1({ S16286 }),
  .A2({ S25957[359] }),
  .ZN({ S16287 })
);
OR2_X1 #() 
OR2_X1_29_ (
  .A1({ S16286 }),
  .A2({ S25957[359] }),
  .ZN({ S16289 })
);
NAND2_X1 #() 
NAND2_X1_2105_ (
  .A1({ S16289 }),
  .A2({ S16287 }),
  .ZN({ S16290 })
);
INV_X1 #() 
INV_X1_674_ (
  .A({ S16290 }),
  .ZN({ S25957[231] })
);
NAND2_X1 #() 
NAND2_X1_2106_ (
  .A1({ S14659 }),
  .A2({ S14646 }),
  .ZN({ S25957[232] })
);
NAND2_X1 #() 
NAND2_X1_2107_ (
  .A1({ S14736 }),
  .A2({ S14735 }),
  .ZN({ S25957[233] })
);
NAND2_X1 #() 
NAND2_X1_2108_ (
  .A1({ S14815 }),
  .A2({ S14814 }),
  .ZN({ S25957[234] })
);
NAND2_X1 #() 
NAND2_X1_2109_ (
  .A1({ S14561 }),
  .A2({ S14585 }),
  .ZN({ S16291 })
);
XNOR2_X1 #() 
XNOR2_X1_107_ (
  .A({ S16291 }),
  .B({ S25957[363] }),
  .ZN({ S25957[235] })
);
NAND2_X1 #() 
NAND2_X1_2110_ (
  .A1({ S14519 }),
  .A2({ S14516 }),
  .ZN({ S25957[236] })
);
XNOR2_X1 #() 
XNOR2_X1_108_ (
  .A({ S14354 }),
  .B({ S25957[366] }),
  .ZN({ S25957[238] })
);
NAND2_X1 #() 
NAND2_X1_2111_ (
  .A1({ S13980 }),
  .A2({ S13958 }),
  .ZN({ S16293 })
);
XOR2_X1 #() 
XOR2_X1_43_ (
  .A({ S16293 }),
  .B({ S25957[368] }),
  .Z({ S25957[240] })
);
NAND2_X1 #() 
NAND2_X1_2112_ (
  .A1({ S14047 }),
  .A2({ S14068 }),
  .ZN({ S16294 })
);
XOR2_X1 #() 
XOR2_X1_44_ (
  .A({ S16294 }),
  .B({ S25957[369] }),
  .Z({ S25957[241] })
);
NAND2_X1 #() 
NAND2_X1_2113_ (
  .A1({ S14133 }),
  .A2({ S14130 }),
  .ZN({ S16295 })
);
XNOR2_X1 #() 
XNOR2_X1_109_ (
  .A({ S16295 }),
  .B({ S25957[370] }),
  .ZN({ S25957[242] })
);
NAND2_X1 #() 
NAND2_X1_2114_ (
  .A1({ S13887 }),
  .A2({ S13888 }),
  .ZN({ S25957[243] })
);
NAND2_X1 #() 
NAND2_X1_2115_ (
  .A1({ S13765 }),
  .A2({ S13750 }),
  .ZN({ S25957[244] })
);
XOR2_X1 #() 
XOR2_X1_45_ (
  .A({ S13683 }),
  .B({ S25957[373] }),
  .Z({ S16296 })
);
INV_X1 #() 
INV_X1_675_ (
  .A({ S16296 }),
  .ZN({ S25957[245] })
);
NAND2_X1 #() 
NAND2_X1_2116_ (
  .A1({ S13607 }),
  .A2({ S13608 }),
  .ZN({ S25957[246] })
);
NAND2_X1 #() 
NAND2_X1_2117_ (
  .A1({ S16097 }),
  .A2({ S16096 }),
  .ZN({ S25957[248] })
);
NAND2_X1 #() 
NAND2_X1_2118_ (
  .A1({ S16175 }),
  .A2({ S16147 }),
  .ZN({ S25957[249] })
);
NAND2_X1 #() 
NAND2_X1_2119_ (
  .A1({ S16246 }),
  .A2({ S16245 }),
  .ZN({ S25957[250] })
);
NAND2_X1 #() 
NAND2_X1_2120_ (
  .A1({ S15987 }),
  .A2({ S15972 }),
  .ZN({ S25957[251] })
);
NAND2_X1 #() 
NAND2_X1_2121_ (
  .A1({ S15886 }),
  .A2({ S15897 }),
  .ZN({ S25957[252] })
);
NAND2_X1 #() 
NAND2_X1_2122_ (
  .A1({ S15819 }),
  .A2({ S15820 }),
  .ZN({ S25957[253] })
);
XOR2_X1 #() 
XOR2_X1_46_ (
  .A({ S15633 }),
  .B({ S25957[383] }),
  .Z({ S25957[255] })
);
XOR2_X1 #() 
XOR2_X1_47_ (
  .A({ S25957[224] }),
  .B({ S25957[320] }),
  .Z({ S25957[192] })
);
NOR2_X1 #() 
NOR2_X1_496_ (
  .A1({ S15445 }),
  .A2({ S15446 }),
  .ZN({ S25957[193] })
);
NOR2_X1 #() 
NOR2_X1_497_ (
  .A1({ S15503 }),
  .A2({ S15504 }),
  .ZN({ S16299 })
);
INV_X1 #() 
INV_X1_676_ (
  .A({ S16299 }),
  .ZN({ S25957[194] })
);
NOR2_X1 #() 
NOR2_X1_498_ (
  .A1({ S15281 }),
  .A2({ S15280 }),
  .ZN({ S16300 })
);
INV_X1 #() 
INV_X1_677_ (
  .A({ S16300 }),
  .ZN({ S25957[195] })
);
NAND2_X1 #() 
NAND2_X1_2123_ (
  .A1({ S15210 }),
  .A2({ S15214 }),
  .ZN({ S25957[196] })
);
NOR2_X1 #() 
NOR2_X1_499_ (
  .A1({ S15131 }),
  .A2({ S15132 }),
  .ZN({ S25957[197] })
);
NOR2_X1 #() 
NOR2_X1_500_ (
  .A1({ S14660 }),
  .A2({ S14664 }),
  .ZN({ S25957[200] })
);
NAND2_X1 #() 
NAND2_X1_2124_ (
  .A1({ S14732 }),
  .A2({ S14737 }),
  .ZN({ S16301 })
);
INV_X1 #() 
INV_X1_678_ (
  .A({ S16301 }),
  .ZN({ S25957[201] })
);
INV_X1 #() 
INV_X1_679_ (
  .A({ S25957[330] }),
  .ZN({ S16302 })
);
XNOR2_X1 #() 
XNOR2_X1_110_ (
  .A({ S25957[234] }),
  .B({ S16302 }),
  .ZN({ S25957[202] })
);
NAND2_X1 #() 
NAND2_X1_2125_ (
  .A1({ S14586 }),
  .A2({ S14588 }),
  .ZN({ S25957[203] })
);
NAND2_X1 #() 
NAND2_X1_2126_ (
  .A1({ S14525 }),
  .A2({ S14527 }),
  .ZN({ S16304 })
);
INV_X1 #() 
INV_X1_680_ (
  .A({ S16304 }),
  .ZN({ S25957[204] })
);
INV_X1 #() 
INV_X1_681_ (
  .A({ S25957[335] }),
  .ZN({ S16305 })
);
XNOR2_X1 #() 
XNOR2_X1_111_ (
  .A({ S25957[239] }),
  .B({ S16305 }),
  .ZN({ S25957[207] })
);
AOI21_X1 #() 
AOI21_X1_1227_ (
  .A({ S25957[464] }),
  .B1({ S13980 }),
  .B2({ S13958 }),
  .ZN({ S16306 })
);
AOI21_X1 #() 
AOI21_X1_1228_ (
  .A({ S10993 }),
  .B1({ S13948 }),
  .B2({ S13926 }),
  .ZN({ S16307 })
);
NOR2_X1 #() 
NOR2_X1_501_ (
  .A1({ S16306 }),
  .A2({ S16307 }),
  .ZN({ S16308 })
);
INV_X1 #() 
INV_X1_682_ (
  .A({ S16308 }),
  .ZN({ S25957[208] })
);
NOR2_X1 #() 
NOR2_X1_502_ (
  .A1({ S14025 }),
  .A2({ S14026 }),
  .ZN({ S16310 })
);
INV_X1 #() 
INV_X1_683_ (
  .A({ S16310 }),
  .ZN({ S25957[209] })
);
NAND2_X1 #() 
NAND2_X1_2127_ (
  .A1({ S14134 }),
  .A2({ S14118 }),
  .ZN({ S25957[210] })
);
NAND2_X1 #() 
NAND2_X1_2128_ (
  .A1({ S13886 }),
  .A2({ S13889 }),
  .ZN({ S25957[211] })
);
INV_X1 #() 
INV_X1_684_ (
  .A({ S25957[340] }),
  .ZN({ S16311 })
);
XNOR2_X1 #() 
XNOR2_X1_112_ (
  .A({ S25957[244] }),
  .B({ S16311 }),
  .ZN({ S25957[212] })
);
AND2_X1 #() 
AND2_X1_127_ (
  .A1({ S13685 }),
  .A2({ S13682 }),
  .ZN({ S25957[213] })
);
NOR2_X1 #() 
NOR2_X1_503_ (
  .A1({ S13614 }),
  .A2({ S13609 }),
  .ZN({ S25957[214] })
);
NOR2_X1 #() 
NOR2_X1_504_ (
  .A1({ S16094 }),
  .A2({ S16098 }),
  .ZN({ S25957[216] })
);
INV_X1 #() 
INV_X1_685_ (
  .A({ S25957[345] }),
  .ZN({ S16312 })
);
XNOR2_X1 #() 
XNOR2_X1_113_ (
  .A({ S25957[249] }),
  .B({ S16312 }),
  .ZN({ S25957[217] })
);
NAND2_X1 #() 
NAND2_X1_2129_ (
  .A1({ S16250 }),
  .A2({ S16251 }),
  .ZN({ S25957[218] })
);
NAND2_X1 #() 
NAND2_X1_2130_ (
  .A1({ S15988 }),
  .A2({ S15991 }),
  .ZN({ S25957[219] })
);
INV_X1 #() 
INV_X1_686_ (
  .A({ S25957[348] }),
  .ZN({ S16314 })
);
XNOR2_X1 #() 
XNOR2_X1_114_ (
  .A({ S25957[252] }),
  .B({ S16314 }),
  .ZN({ S25957[220] })
);
NAND2_X1 #() 
NAND2_X1_2131_ (
  .A1({ S15823 }),
  .A2({ S15824 }),
  .ZN({ S25957[221] })
);
XOR2_X1 #() 
XOR2_X1_48_ (
  .A({ S25957[254] }),
  .B({ S25957[350] }),
  .Z({ S25957[222] })
);
XOR2_X1 #() 
XOR2_X1_49_ (
  .A({ S25957[192] }),
  .B({ S25957[288] }),
  .Z({ S25957[160] })
);
NOR2_X1 #() 
NOR2_X1_505_ (
  .A1({ S15447 }),
  .A2({ S15443 }),
  .ZN({ S25957[161] })
);
XNOR2_X1 #() 
XNOR2_X1_115_ (
  .A({ S16299 }),
  .B({ S25957[290] }),
  .ZN({ S25957[162] })
);
NAND2_X1 #() 
NAND2_X1_2132_ (
  .A1({ S15282 }),
  .A2({ S15301 }),
  .ZN({ S16316 })
);
INV_X1 #() 
INV_X1_687_ (
  .A({ S16316 }),
  .ZN({ S25957[163] })
);
XOR2_X1 #() 
XOR2_X1_50_ (
  .A({ S25957[196] }),
  .B({ S25957[292] }),
  .Z({ S25957[164] })
);
NAND2_X1 #() 
NAND2_X1_2133_ (
  .A1({ S15133 }),
  .A2({ S15129 }),
  .ZN({ S16317 })
);
INV_X1 #() 
INV_X1_688_ (
  .A({ S16317 }),
  .ZN({ S25957[165] })
);
XOR2_X1 #() 
XOR2_X1_51_ (
  .A({ S25957[198] }),
  .B({ S25957[294] }),
  .Z({ S25957[166] })
);
NAND2_X1 #() 
NAND2_X1_2134_ (
  .A1({ S14665 }),
  .A2({ S14669 }),
  .ZN({ S25957[168] })
);
XNOR2_X1 #() 
XNOR2_X1_116_ (
  .A({ S16301 }),
  .B({ S25957[297] }),
  .ZN({ S25957[169] })
);
NOR2_X1 #() 
NOR2_X1_506_ (
  .A1({ S14813 }),
  .A2({ S14816 }),
  .ZN({ S16318 })
);
INV_X1 #() 
INV_X1_689_ (
  .A({ S16318 }),
  .ZN({ S25957[170] })
);
XNOR2_X1 #() 
XNOR2_X1_117_ (
  .A({ S25957[203] }),
  .B({ S16278 }),
  .ZN({ S25957[171] })
);
XNOR2_X1 #() 
XNOR2_X1_118_ (
  .A({ S16304 }),
  .B({ S25957[300] }),
  .ZN({ S25957[172] })
);
INV_X1 #() 
INV_X1_690_ (
  .A({ S25957[301] }),
  .ZN({ S16320 })
);
XNOR2_X1 #() 
XNOR2_X1_119_ (
  .A({ S25957[205] }),
  .B({ S16320 }),
  .ZN({ S25957[173] })
);
XOR2_X1 #() 
XOR2_X1_52_ (
  .A({ S25957[206] }),
  .B({ S25957[302] }),
  .Z({ S25957[174] })
);
NAND2_X1 #() 
NAND2_X1_2135_ (
  .A1({ S25957[208] }),
  .A2({ S16279 }),
  .ZN({ S16321 })
);
NAND2_X1 #() 
NAND2_X1_2136_ (
  .A1({ S16308 }),
  .A2({ S25957[304] }),
  .ZN({ S16322 })
);
NAND2_X1 #() 
NAND2_X1_2137_ (
  .A1({ S16321 }),
  .A2({ S16322 }),
  .ZN({ S25957[176] })
);
XNOR2_X1 #() 
XNOR2_X1_120_ (
  .A({ S16310 }),
  .B({ S25957[305] }),
  .ZN({ S25957[177] })
);
XNOR2_X1 #() 
XNOR2_X1_121_ (
  .A({ S25957[210] }),
  .B({ S25957[306] }),
  .ZN({ S16323 })
);
INV_X1 #() 
INV_X1_691_ (
  .A({ S16323 }),
  .ZN({ S25957[178] })
);
NOR2_X1 #() 
NOR2_X1_507_ (
  .A1({ S13890 }),
  .A2({ S13894 }),
  .ZN({ S25957[179] })
);
NOR2_X1 #() 
NOR2_X1_508_ (
  .A1({ S13767 }),
  .A2({ S13770 }),
  .ZN({ S25957[180] })
);
XNOR2_X1 #() 
XNOR2_X1_122_ (
  .A({ S25957[213] }),
  .B({ S25957[309] }),
  .ZN({ S16325 })
);
INV_X1 #() 
INV_X1_692_ (
  .A({ S16325 }),
  .ZN({ S25957[181] })
);
INV_X1 #() 
INV_X1_693_ (
  .A({ S25957[310] }),
  .ZN({ S16326 })
);
XNOR2_X1 #() 
XNOR2_X1_123_ (
  .A({ S25957[214] }),
  .B({ S16326 }),
  .ZN({ S25957[182] })
);
XNOR2_X1 #() 
XNOR2_X1_124_ (
  .A({ S25957[215] }),
  .B({ S10651 }),
  .ZN({ S25957[183] })
);
XOR2_X1 #() 
XOR2_X1_53_ (
  .A({ S25957[216] }),
  .B({ S25957[312] }),
  .Z({ S25957[184] })
);
NOR2_X1 #() 
NOR2_X1_509_ (
  .A1({ S16176 }),
  .A2({ S16180 }),
  .ZN({ S25957[185] })
);
NAND2_X1 #() 
NAND2_X1_2138_ (
  .A1({ S16254 }),
  .A2({ S16255 }),
  .ZN({ S16328 })
);
INV_X1 #() 
INV_X1_694_ (
  .A({ S16328 }),
  .ZN({ S25957[186] })
);
XOR2_X1 #() 
XOR2_X1_54_ (
  .A({ S25957[251] }),
  .B({ S25957[443] }),
  .Z({ S25957[187] })
);
NOR2_X1 #() 
NOR2_X1_510_ (
  .A1({ S15898 }),
  .A2({ S15903 }),
  .ZN({ S16329 })
);
INV_X1 #() 
INV_X1_695_ (
  .A({ S16329 }),
  .ZN({ S25957[188] })
);
XOR2_X1 #() 
XOR2_X1_55_ (
  .A({ S25957[221] }),
  .B({ S25957[317] }),
  .Z({ S25957[189] })
);
NOR2_X1 #() 
NOR2_X1_511_ (
  .A1({ S15724 }),
  .A2({ S15725 }),
  .ZN({ S25957[190] })
);
XOR2_X1 #() 
XOR2_X1_56_ (
  .A({ S25957[223] }),
  .B({ S25957[319] }),
  .Z({ S25957[191] })
);
NAND3_X1 #() 
NAND3_X1_2390_ (
  .A1({ S16100 }),
  .A2({ S16101 }),
  .A3({ S25957[408] }),
  .ZN({ S16330 })
);
OAI21_X1 #() 
OAI21_X1_1144_ (
  .A({ S12012 }),
  .B1({ S16094 }),
  .B2({ S16098 }),
  .ZN({ S16331 })
);
OAI21_X1 #() 
OAI21_X1_1145_ (
  .A({ S14841 }),
  .B1({ S16176 }),
  .B2({ S16180 }),
  .ZN({ S16333 })
);
NAND3_X1 #() 
NAND3_X1_2391_ (
  .A1({ S16182 }),
  .A2({ S16183 }),
  .A3({ S25957[281] }),
  .ZN({ S16334 })
);
NAND4_X1 #() 
NAND4_X1_292_ (
  .A1({ S16331 }),
  .A2({ S16330 }),
  .A3({ S16333 }),
  .A4({ S16334 }),
  .ZN({ S16335 })
);
INV_X1 #() 
INV_X1_696_ (
  .A({ S16335 }),
  .ZN({ S55 })
);
NAND4_X1 #() 
NAND4_X1_293_ (
  .A1({ S16099 }),
  .A2({ S16102 }),
  .A3({ S16181 }),
  .A4({ S16184 }),
  .ZN({ S57 })
);
INV_X1 #() 
INV_X1_697_ (
  .A({ S25957[224] }),
  .ZN({ S16336 })
);
NAND2_X1 #() 
NAND2_X1_2139_ (
  .A1({ S16331 }),
  .A2({ S16330 }),
  .ZN({ S16337 })
);
NAND2_X1 #() 
NAND2_X1_2140_ (
  .A1({ S16333 }),
  .A2({ S16334 }),
  .ZN({ S16338 })
);
NAND3_X1 #() 
NAND3_X1_2392_ (
  .A1({ S16254 }),
  .A2({ S16255 }),
  .A3({ S25957[282] }),
  .ZN({ S16339 })
);
NAND3_X1 #() 
NAND3_X1_2393_ (
  .A1({ S16249 }),
  .A2({ S16252 }),
  .A3({ S14834 }),
  .ZN({ S16340 })
);
NAND4_X1 #() 
NAND4_X1_294_ (
  .A1({ S16339 }),
  .A2({ S16340 }),
  .A3({ S16337 }),
  .A4({ S16338 }),
  .ZN({ S16342 })
);
AOI21_X1 #() 
AOI21_X1_1229_ (
  .A({ S25957[155] }),
  .B1({ S25957[152] }),
  .B2({ S25957[153] }),
  .ZN({ S16343 })
);
NAND4_X1 #() 
NAND4_X1_295_ (
  .A1({ S16253 }),
  .A2({ S16256 }),
  .A3({ S16337 }),
  .A4({ S16338 }),
  .ZN({ S16344 })
);
NAND4_X1 #() 
NAND4_X1_296_ (
  .A1({ S16331 }),
  .A2({ S16330 }),
  .A3({ S16181 }),
  .A4({ S16184 }),
  .ZN({ S16345 })
);
INV_X1 #() 
INV_X1_698_ (
  .A({ S16345 }),
  .ZN({ S16346 })
);
AOI21_X1 #() 
AOI21_X1_1230_ (
  .A({ S54 }),
  .B1({ S25957[154] }),
  .B2({ S16346 }),
  .ZN({ S16347 })
);
AOI22_X1 #() 
AOI22_X1_273_ (
  .A1({ S16347 }),
  .A2({ S16344 }),
  .B1({ S16343 }),
  .B2({ S16342 }),
  .ZN({ S16348 })
);
NAND3_X1 #() 
NAND3_X1_2394_ (
  .A1({ S16253 }),
  .A2({ S16256 }),
  .A3({ S25957[152] }),
  .ZN({ S16349 })
);
AOI21_X1 #() 
AOI21_X1_1231_ (
  .A({ S25957[155] }),
  .B1({ S16337 }),
  .B2({ S25957[153] }),
  .ZN({ S16350 })
);
NAND2_X1 #() 
NAND2_X1_2141_ (
  .A1({ S16350 }),
  .A2({ S16349 }),
  .ZN({ S16351 })
);
NAND3_X1 #() 
NAND3_X1_2395_ (
  .A1({ S16339 }),
  .A2({ S16340 }),
  .A3({ S25957[152] }),
  .ZN({ S16353 })
);
NAND3_X1 #() 
NAND3_X1_2396_ (
  .A1({ S16353 }),
  .A2({ S25957[155] }),
  .A3({ S57 }),
  .ZN({ S16354 })
);
NAND3_X1 #() 
NAND3_X1_2397_ (
  .A1({ S16354 }),
  .A2({ S16351 }),
  .A3({ S25957[156] }),
  .ZN({ S16355 })
);
OAI211_X1 #() 
OAI211_X1_767_ (
  .A({ S16355 }),
  .B({ S25957[157] }),
  .C1({ S16348 }),
  .C2({ S25957[156] }),
  .ZN({ S16356 })
);
OAI21_X1 #() 
OAI21_X1_1146_ (
  .A({ S25957[284] }),
  .B1({ S15898 }),
  .B2({ S15903 }),
  .ZN({ S16357 })
);
NAND3_X1 #() 
NAND3_X1_2398_ (
  .A1({ S15905 }),
  .A2({ S15906 }),
  .A3({ S14852 }),
  .ZN({ S16358 })
);
NAND2_X1 #() 
NAND2_X1_2142_ (
  .A1({ S16357 }),
  .A2({ S16358 }),
  .ZN({ S16359 })
);
NAND4_X1 #() 
NAND4_X1_297_ (
  .A1({ S16099 }),
  .A2({ S16102 }),
  .A3({ S16333 }),
  .A4({ S16334 }),
  .ZN({ S16360 })
);
NAND2_X1 #() 
NAND2_X1_2143_ (
  .A1({ S16360 }),
  .A2({ S16345 }),
  .ZN({ S16361 })
);
NOR2_X1 #() 
NOR2_X1_512_ (
  .A1({ S16361 }),
  .A2({ S25957[154] }),
  .ZN({ S16362 })
);
AOI21_X1 #() 
AOI21_X1_1232_ (
  .A({ S16359 }),
  .B1({ S16362 }),
  .B2({ S25957[155] }),
  .ZN({ S16364 })
);
NAND4_X1 #() 
NAND4_X1_298_ (
  .A1({ S16360 }),
  .A2({ S16345 }),
  .A3({ S16339 }),
  .A4({ S16340 }),
  .ZN({ S16365 })
);
NAND3_X1 #() 
NAND3_X1_2399_ (
  .A1({ S16253 }),
  .A2({ S16256 }),
  .A3({ S16338 }),
  .ZN({ S16366 })
);
NAND3_X1 #() 
NAND3_X1_2400_ (
  .A1({ S16365 }),
  .A2({ S54 }),
  .A3({ S16366 }),
  .ZN({ S16367 })
);
NAND4_X1 #() 
NAND4_X1_299_ (
  .A1({ S16253 }),
  .A2({ S16256 }),
  .A3({ S25957[152] }),
  .A4({ S16338 }),
  .ZN({ S16368 })
);
NAND3_X1 #() 
NAND3_X1_2401_ (
  .A1({ S16342 }),
  .A2({ S16368 }),
  .A3({ S54 }),
  .ZN({ S16369 })
);
NAND4_X1 #() 
NAND4_X1_300_ (
  .A1({ S16339 }),
  .A2({ S16340 }),
  .A3({ S25957[152] }),
  .A4({ S25957[153] }),
  .ZN({ S16370 })
);
AOI21_X1 #() 
AOI21_X1_1233_ (
  .A({ S54 }),
  .B1({ S16337 }),
  .B2({ S16338 }),
  .ZN({ S16371 })
);
AOI21_X1 #() 
AOI21_X1_1234_ (
  .A({ S25957[156] }),
  .B1({ S16370 }),
  .B2({ S16371 }),
  .ZN({ S16372 })
);
AOI22_X1 #() 
AOI22_X1_274_ (
  .A1({ S16364 }),
  .A2({ S16367 }),
  .B1({ S16372 }),
  .B2({ S16369 }),
  .ZN({ S16373 })
);
OAI211_X1 #() 
OAI211_X1_768_ (
  .A({ S16356 }),
  .B({ S15729 }),
  .C1({ S16373 }),
  .C2({ S25957[157] }),
  .ZN({ S16375 })
);
INV_X1 #() 
INV_X1_699_ (
  .A({ S25957[157] }),
  .ZN({ S16376 })
);
NAND3_X1 #() 
NAND3_X1_2402_ (
  .A1({ S16253 }),
  .A2({ S16256 }),
  .A3({ S16337 }),
  .ZN({ S16377 })
);
NAND2_X1 #() 
NAND2_X1_2144_ (
  .A1({ S16377 }),
  .A2({ S54 }),
  .ZN({ S16378 })
);
NAND3_X1 #() 
NAND3_X1_2403_ (
  .A1({ S16339 }),
  .A2({ S16340 }),
  .A3({ S16338 }),
  .ZN({ S16379 })
);
NAND4_X1 #() 
NAND4_X1_301_ (
  .A1({ S16253 }),
  .A2({ S16256 }),
  .A3({ S16337 }),
  .A4({ S25957[153] }),
  .ZN({ S16380 })
);
NAND4_X1 #() 
NAND4_X1_302_ (
  .A1({ S16380 }),
  .A2({ S16353 }),
  .A3({ S16379 }),
  .A4({ S25957[155] }),
  .ZN({ S16381 })
);
NAND3_X1 #() 
NAND3_X1_2404_ (
  .A1({ S16381 }),
  .A2({ S16359 }),
  .A3({ S16378 }),
  .ZN({ S16382 })
);
NAND3_X1 #() 
NAND3_X1_2405_ (
  .A1({ S16339 }),
  .A2({ S16340 }),
  .A3({ S16337 }),
  .ZN({ S16383 })
);
NAND2_X1 #() 
NAND2_X1_2145_ (
  .A1({ S16350 }),
  .A2({ S16383 }),
  .ZN({ S16384 })
);
NAND2_X1 #() 
NAND2_X1_2146_ (
  .A1({ S16339 }),
  .A2({ S16340 }),
  .ZN({ S16386 })
);
NAND2_X1 #() 
NAND2_X1_2147_ (
  .A1({ S16386 }),
  .A2({ S16335 }),
  .ZN({ S16387 })
);
NAND3_X1 #() 
NAND3_X1_2406_ (
  .A1({ S16387 }),
  .A2({ S16365 }),
  .A3({ S25957[155] }),
  .ZN({ S16388 })
);
NAND3_X1 #() 
NAND3_X1_2407_ (
  .A1({ S16388 }),
  .A2({ S25957[156] }),
  .A3({ S16384 }),
  .ZN({ S16389 })
);
AND2_X1 #() 
AND2_X1_128_ (
  .A1({ S16389 }),
  .A2({ S16382 }),
  .ZN({ S16390 })
);
NAND3_X1 #() 
NAND3_X1_2408_ (
  .A1({ S16380 }),
  .A2({ S54 }),
  .A3({ S16379 }),
  .ZN({ S16391 })
);
NAND3_X1 #() 
NAND3_X1_2409_ (
  .A1({ S16335 }),
  .A2({ S16339 }),
  .A3({ S16340 }),
  .ZN({ S16392 })
);
NAND3_X1 #() 
NAND3_X1_2410_ (
  .A1({ S16392 }),
  .A2({ S16377 }),
  .A3({ S25957[155] }),
  .ZN({ S16393 })
);
AND2_X1 #() 
AND2_X1_129_ (
  .A1({ S16391 }),
  .A2({ S16393 }),
  .ZN({ S16394 })
);
NAND3_X1 #() 
NAND3_X1_2411_ (
  .A1({ S16392 }),
  .A2({ S16349 }),
  .A3({ S25957[155] }),
  .ZN({ S16395 })
);
NAND2_X1 #() 
NAND2_X1_2148_ (
  .A1({ S25957[152] }),
  .A2({ S54 }),
  .ZN({ S16397 })
);
NAND2_X1 #() 
NAND2_X1_2149_ (
  .A1({ S54 }),
  .A2({ S25957[153] }),
  .ZN({ S16398 })
);
OAI211_X1 #() 
OAI211_X1_769_ (
  .A({ S16359 }),
  .B({ S16398 }),
  .C1({ S16386 }),
  .C2({ S16397 }),
  .ZN({ S16399 })
);
INV_X1 #() 
INV_X1_700_ (
  .A({ S16399 }),
  .ZN({ S16400 })
);
NAND2_X1 #() 
NAND2_X1_2150_ (
  .A1({ S16400 }),
  .A2({ S16395 }),
  .ZN({ S16401 })
);
OAI211_X1 #() 
OAI211_X1_770_ (
  .A({ S16401 }),
  .B({ S16376 }),
  .C1({ S16394 }),
  .C2({ S16359 }),
  .ZN({ S16402 })
);
OAI211_X1 #() 
OAI211_X1_771_ (
  .A({ S16402 }),
  .B({ S25957[158] }),
  .C1({ S16390 }),
  .C2({ S16376 }),
  .ZN({ S16403 })
);
NAND3_X1 #() 
NAND3_X1_2412_ (
  .A1({ S16403 }),
  .A2({ S16375 }),
  .A3({ S15640 }),
  .ZN({ S16404 })
);
NAND2_X1 #() 
NAND2_X1_2151_ (
  .A1({ S16342 }),
  .A2({ S54 }),
  .ZN({ S16405 })
);
INV_X1 #() 
INV_X1_701_ (
  .A({ S16360 }),
  .ZN({ S16406 })
);
AOI21_X1 #() 
AOI21_X1_1235_ (
  .A({ S16406 }),
  .B1({ S16386 }),
  .B2({ S16345 }),
  .ZN({ S16408 })
);
OAI211_X1 #() 
OAI211_X1_772_ (
  .A({ S16359 }),
  .B({ S16405 }),
  .C1({ S16408 }),
  .C2({ S54 }),
  .ZN({ S16409 })
);
NAND3_X1 #() 
NAND3_X1_2413_ (
  .A1({ S16386 }),
  .A2({ S16346 }),
  .A3({ S54 }),
  .ZN({ S16410 })
);
NAND2_X1 #() 
NAND2_X1_2152_ (
  .A1({ S16342 }),
  .A2({ S25957[155] }),
  .ZN({ S16411 })
);
AOI21_X1 #() 
AOI21_X1_1236_ (
  .A({ S25957[152] }),
  .B1({ S16253 }),
  .B2({ S16256 }),
  .ZN({ S16412 })
);
AOI22_X1 #() 
AOI22_X1_275_ (
  .A1({ S15996 }),
  .A2({ S15993 }),
  .B1({ S16181 }),
  .B2({ S16184 }),
  .ZN({ S16413 })
);
NAND2_X1 #() 
NAND2_X1_2153_ (
  .A1({ S16412 }),
  .A2({ S16413 }),
  .ZN({ S16414 })
);
NAND3_X1 #() 
NAND3_X1_2414_ (
  .A1({ S16411 }),
  .A2({ S16414 }),
  .A3({ S16410 }),
  .ZN({ S16415 })
);
OAI211_X1 #() 
OAI211_X1_773_ (
  .A({ S16409 }),
  .B({ S25957[157] }),
  .C1({ S16359 }),
  .C2({ S16415 }),
  .ZN({ S16416 })
);
NAND4_X1 #() 
NAND4_X1_303_ (
  .A1({ S16339 }),
  .A2({ S16340 }),
  .A3({ S16337 }),
  .A4({ S25957[153] }),
  .ZN({ S16417 })
);
NAND2_X1 #() 
NAND2_X1_2154_ (
  .A1({ S16417 }),
  .A2({ S16349 }),
  .ZN({ S16419 })
);
NAND2_X1 #() 
NAND2_X1_2155_ (
  .A1({ S16419 }),
  .A2({ S54 }),
  .ZN({ S16420 })
);
NAND2_X1 #() 
NAND2_X1_2156_ (
  .A1({ S16337 }),
  .A2({ S25957[155] }),
  .ZN({ S16421 })
);
NAND2_X1 #() 
NAND2_X1_2157_ (
  .A1({ S16421 }),
  .A2({ S16359 }),
  .ZN({ S16422 })
);
NAND3_X1 #() 
NAND3_X1_2415_ (
  .A1({ S25957[154] }),
  .A2({ S16359 }),
  .A3({ S25957[153] }),
  .ZN({ S16423 })
);
NAND2_X1 #() 
NAND2_X1_2158_ (
  .A1({ S16423 }),
  .A2({ S16422 }),
  .ZN({ S16424 })
);
NAND2_X1 #() 
NAND2_X1_2159_ (
  .A1({ S16420 }),
  .A2({ S16424 }),
  .ZN({ S16425 })
);
NAND2_X1 #() 
NAND2_X1_2160_ (
  .A1({ S16335 }),
  .A2({ S57 }),
  .ZN({ S16426 })
);
NOR2_X1 #() 
NOR2_X1_513_ (
  .A1({ S16426 }),
  .A2({ S25957[154] }),
  .ZN({ S16427 })
);
NAND3_X1 #() 
NAND3_X1_2416_ (
  .A1({ S16339 }),
  .A2({ S16340 }),
  .A3({ S25957[153] }),
  .ZN({ S16428 })
);
NAND2_X1 #() 
NAND2_X1_2161_ (
  .A1({ S16428 }),
  .A2({ S25957[155] }),
  .ZN({ S16430 })
);
OAI211_X1 #() 
OAI211_X1_774_ (
  .A({ S16430 }),
  .B({ S25957[156] }),
  .C1({ S16427 }),
  .C2({ S25957[155] }),
  .ZN({ S16431 })
);
NAND3_X1 #() 
NAND3_X1_2417_ (
  .A1({ S16425 }),
  .A2({ S16376 }),
  .A3({ S16431 }),
  .ZN({ S16432 })
);
NAND3_X1 #() 
NAND3_X1_2418_ (
  .A1({ S16416 }),
  .A2({ S16432 }),
  .A3({ S15729 }),
  .ZN({ S16433 })
);
AOI21_X1 #() 
AOI21_X1_1237_ (
  .A({ S25957[155] }),
  .B1({ S16344 }),
  .B2({ S16353 }),
  .ZN({ S16434 })
);
NAND3_X1 #() 
NAND3_X1_2419_ (
  .A1({ S16339 }),
  .A2({ S16340 }),
  .A3({ S25957[155] }),
  .ZN({ S16435 })
);
OAI22_X1 #() 
OAI22_X1_51_ (
  .A1({ S16435 }),
  .A2({ S16406 }),
  .B1({ S16386 }),
  .B2({ S16398 }),
  .ZN({ S16436 })
);
OAI21_X1 #() 
OAI21_X1_1147_ (
  .A({ S25957[156] }),
  .B1({ S16434 }),
  .B2({ S16436 }),
  .ZN({ S16437 })
);
NAND3_X1 #() 
NAND3_X1_2420_ (
  .A1({ S16368 }),
  .A2({ S25957[155] }),
  .A3({ S16383 }),
  .ZN({ S16438 })
);
NAND2_X1 #() 
NAND2_X1_2162_ (
  .A1({ S16361 }),
  .A2({ S16386 }),
  .ZN({ S16439 })
);
NAND3_X1 #() 
NAND3_X1_2421_ (
  .A1({ S16439 }),
  .A2({ S54 }),
  .A3({ S16428 }),
  .ZN({ S16441 })
);
NAND3_X1 #() 
NAND3_X1_2422_ (
  .A1({ S16441 }),
  .A2({ S16359 }),
  .A3({ S16438 }),
  .ZN({ S16442 })
);
AOI21_X1 #() 
AOI21_X1_1238_ (
  .A({ S16376 }),
  .B1({ S16442 }),
  .B2({ S16437 }),
  .ZN({ S16443 })
);
NOR2_X1 #() 
NOR2_X1_514_ (
  .A1({ S16435 }),
  .A2({ S16361 }),
  .ZN({ S16444 })
);
NAND3_X1 #() 
NAND3_X1_2423_ (
  .A1({ S16360 }),
  .A2({ S16253 }),
  .A3({ S16256 }),
  .ZN({ S16445 })
);
NAND3_X1 #() 
NAND3_X1_2424_ (
  .A1({ S16345 }),
  .A2({ S16339 }),
  .A3({ S16340 }),
  .ZN({ S16446 })
);
AOI21_X1 #() 
AOI21_X1_1239_ (
  .A({ S25957[155] }),
  .B1({ S16446 }),
  .B2({ S16445 }),
  .ZN({ S16447 })
);
NOR3_X1 #() 
NOR3_X1_66_ (
  .A1({ S16447 }),
  .A2({ S16444 }),
  .A3({ S16359 }),
  .ZN({ S16448 })
);
AOI21_X1 #() 
AOI21_X1_1240_ (
  .A({ S16360 }),
  .B1({ S16340 }),
  .B2({ S16339 }),
  .ZN({ S16449 })
);
NOR2_X1 #() 
NOR2_X1_515_ (
  .A1({ S16449 }),
  .A2({ S25957[155] }),
  .ZN({ S16450 })
);
NAND2_X1 #() 
NAND2_X1_2163_ (
  .A1({ S16395 }),
  .A2({ S16359 }),
  .ZN({ S16452 })
);
OAI21_X1 #() 
OAI21_X1_1148_ (
  .A({ S16376 }),
  .B1({ S16452 }),
  .B2({ S16450 }),
  .ZN({ S16453 })
);
OAI21_X1 #() 
OAI21_X1_1149_ (
  .A({ S25957[158] }),
  .B1({ S16453 }),
  .B2({ S16448 }),
  .ZN({ S16454 })
);
OAI211_X1 #() 
OAI211_X1_775_ (
  .A({ S16433 }),
  .B({ S25957[159] }),
  .C1({ S16443 }),
  .C2({ S16454 }),
  .ZN({ S16455 })
);
NAND3_X1 #() 
NAND3_X1_2425_ (
  .A1({ S16404 }),
  .A2({ S16455 }),
  .A3({ S16336 }),
  .ZN({ S16456 })
);
NAND3_X1 #() 
NAND3_X1_2426_ (
  .A1({ S16389 }),
  .A2({ S16382 }),
  .A3({ S25957[157] }),
  .ZN({ S16457 })
);
AOI21_X1 #() 
AOI21_X1_1241_ (
  .A({ S16359 }),
  .B1({ S16391 }),
  .B2({ S16393 }),
  .ZN({ S16458 })
);
AOI21_X1 #() 
AOI21_X1_1242_ (
  .A({ S54 }),
  .B1({ S16370 }),
  .B2({ S16377 }),
  .ZN({ S16459 })
);
NOR2_X1 #() 
NOR2_X1_516_ (
  .A1({ S16459 }),
  .A2({ S16399 }),
  .ZN({ S16460 })
);
OAI21_X1 #() 
OAI21_X1_1150_ (
  .A({ S16376 }),
  .B1({ S16458 }),
  .B2({ S16460 }),
  .ZN({ S16461 })
);
NAND3_X1 #() 
NAND3_X1_2427_ (
  .A1({ S16461 }),
  .A2({ S16457 }),
  .A3({ S25957[158] }),
  .ZN({ S16463 })
);
NAND2_X1 #() 
NAND2_X1_2164_ (
  .A1({ S16354 }),
  .A2({ S16351 }),
  .ZN({ S16464 })
);
NAND2_X1 #() 
NAND2_X1_2165_ (
  .A1({ S16464 }),
  .A2({ S25957[156] }),
  .ZN({ S16465 })
);
NAND2_X1 #() 
NAND2_X1_2166_ (
  .A1({ S16342 }),
  .A2({ S16343 }),
  .ZN({ S16466 })
);
INV_X1 #() 
INV_X1_702_ (
  .A({ S16344 }),
  .ZN({ S16467 })
);
NAND2_X1 #() 
NAND2_X1_2167_ (
  .A1({ S25957[154] }),
  .A2({ S16346 }),
  .ZN({ S16468 })
);
NAND2_X1 #() 
NAND2_X1_2168_ (
  .A1({ S16468 }),
  .A2({ S25957[155] }),
  .ZN({ S16469 })
);
OAI211_X1 #() 
OAI211_X1_776_ (
  .A({ S16359 }),
  .B({ S16466 }),
  .C1({ S16469 }),
  .C2({ S16467 }),
  .ZN({ S16470 })
);
NAND3_X1 #() 
NAND3_X1_2428_ (
  .A1({ S16470 }),
  .A2({ S16465 }),
  .A3({ S25957[157] }),
  .ZN({ S16471 })
);
NAND2_X1 #() 
NAND2_X1_2169_ (
  .A1({ S16364 }),
  .A2({ S16367 }),
  .ZN({ S16472 })
);
AOI21_X1 #() 
AOI21_X1_1243_ (
  .A({ S25957[157] }),
  .B1({ S16372 }),
  .B2({ S16369 }),
  .ZN({ S16474 })
);
NAND2_X1 #() 
NAND2_X1_2170_ (
  .A1({ S16472 }),
  .A2({ S16474 }),
  .ZN({ S16475 })
);
NAND3_X1 #() 
NAND3_X1_2429_ (
  .A1({ S16471 }),
  .A2({ S16475 }),
  .A3({ S15729 }),
  .ZN({ S16476 })
);
NAND3_X1 #() 
NAND3_X1_2430_ (
  .A1({ S16476 }),
  .A2({ S16463 }),
  .A3({ S15640 }),
  .ZN({ S16477 })
);
NOR2_X1 #() 
NOR2_X1_517_ (
  .A1({ S16452 }),
  .A2({ S16450 }),
  .ZN({ S16478 })
);
OAI21_X1 #() 
OAI21_X1_1151_ (
  .A({ S16376 }),
  .B1({ S16478 }),
  .B2({ S16448 }),
  .ZN({ S16479 })
);
NAND3_X1 #() 
NAND3_X1_2431_ (
  .A1({ S16442 }),
  .A2({ S16437 }),
  .A3({ S25957[157] }),
  .ZN({ S16480 })
);
NAND3_X1 #() 
NAND3_X1_2432_ (
  .A1({ S16479 }),
  .A2({ S25957[158] }),
  .A3({ S16480 }),
  .ZN({ S16481 })
);
AOI22_X1 #() 
AOI22_X1_276_ (
  .A1({ S16419 }),
  .A2({ S54 }),
  .B1({ S16423 }),
  .B2({ S16422 }),
  .ZN({ S16482 })
);
NAND3_X1 #() 
NAND3_X1_2433_ (
  .A1({ S25957[154] }),
  .A2({ S25957[155] }),
  .A3({ S25957[153] }),
  .ZN({ S16483 })
);
NAND3_X1 #() 
NAND3_X1_2434_ (
  .A1({ S16361 }),
  .A2({ S54 }),
  .A3({ S16386 }),
  .ZN({ S16485 })
);
AOI21_X1 #() 
AOI21_X1_1244_ (
  .A({ S16359 }),
  .B1({ S16485 }),
  .B2({ S16483 }),
  .ZN({ S16486 })
);
OAI21_X1 #() 
OAI21_X1_1152_ (
  .A({ S16376 }),
  .B1({ S16482 }),
  .B2({ S16486 }),
  .ZN({ S16487 })
);
NAND2_X1 #() 
NAND2_X1_2171_ (
  .A1({ S16415 }),
  .A2({ S25957[156] }),
  .ZN({ S16488 })
);
INV_X1 #() 
INV_X1_703_ (
  .A({ S57 }),
  .ZN({ S16489 })
);
AOI21_X1 #() 
AOI21_X1_1245_ (
  .A({ S25957[155] }),
  .B1({ S25957[154] }),
  .B2({ S16489 }),
  .ZN({ S16490 })
);
NAND3_X1 #() 
NAND3_X1_2435_ (
  .A1({ S16345 }),
  .A2({ S16253 }),
  .A3({ S16256 }),
  .ZN({ S16491 })
);
AOI21_X1 #() 
AOI21_X1_1246_ (
  .A({ S54 }),
  .B1({ S16491 }),
  .B2({ S16360 }),
  .ZN({ S16492 })
);
OAI21_X1 #() 
OAI21_X1_1153_ (
  .A({ S16359 }),
  .B1({ S16492 }),
  .B2({ S16490 }),
  .ZN({ S16493 })
);
NAND3_X1 #() 
NAND3_X1_2436_ (
  .A1({ S16488 }),
  .A2({ S16493 }),
  .A3({ S25957[157] }),
  .ZN({ S16494 })
);
NAND3_X1 #() 
NAND3_X1_2437_ (
  .A1({ S16494 }),
  .A2({ S15729 }),
  .A3({ S16487 }),
  .ZN({ S16496 })
);
NAND3_X1 #() 
NAND3_X1_2438_ (
  .A1({ S16481 }),
  .A2({ S25957[159] }),
  .A3({ S16496 }),
  .ZN({ S16497 })
);
NAND3_X1 #() 
NAND3_X1_2439_ (
  .A1({ S16497 }),
  .A2({ S25957[224] }),
  .A3({ S16477 }),
  .ZN({ S16498 })
);
NAND2_X1 #() 
NAND2_X1_2172_ (
  .A1({ S16456 }),
  .A2({ S16498 }),
  .ZN({ S25957[96] })
);
INV_X1 #() 
INV_X1_704_ (
  .A({ S25957[225] }),
  .ZN({ S16499 })
);
NAND3_X1 #() 
NAND3_X1_2440_ (
  .A1({ S16365 }),
  .A2({ S25957[155] }),
  .A3({ S16377 }),
  .ZN({ S16500 })
);
AOI21_X1 #() 
AOI21_X1_1247_ (
  .A({ S16337 }),
  .B1({ S16339 }),
  .B2({ S16340 }),
  .ZN({ S16501 })
);
NOR2_X1 #() 
NOR2_X1_518_ (
  .A1({ S16501 }),
  .A2({ S25957[155] }),
  .ZN({ S16502 })
);
NAND2_X1 #() 
NAND2_X1_2173_ (
  .A1({ S25957[154] }),
  .A2({ S16360 }),
  .ZN({ S16503 })
);
NAND2_X1 #() 
NAND2_X1_2174_ (
  .A1({ S16502 }),
  .A2({ S16503 }),
  .ZN({ S16504 })
);
NAND3_X1 #() 
NAND3_X1_2441_ (
  .A1({ S16504 }),
  .A2({ S25957[156] }),
  .A3({ S16500 }),
  .ZN({ S16506 })
);
NAND2_X1 #() 
NAND2_X1_2175_ (
  .A1({ S16386 }),
  .A2({ S25957[153] }),
  .ZN({ S16507 })
);
AOI21_X1 #() 
AOI21_X1_1248_ (
  .A({ S25957[155] }),
  .B1({ S25957[152] }),
  .B2({ S16338 }),
  .ZN({ S16508 })
);
AOI22_X1 #() 
AOI22_X1_277_ (
  .A1({ S16507 }),
  .A2({ S16508 }),
  .B1({ S25957[155] }),
  .B2({ S16445 }),
  .ZN({ S16509 })
);
OAI211_X1 #() 
OAI211_X1_777_ (
  .A({ S16506 }),
  .B({ S25957[157] }),
  .C1({ S25957[156] }),
  .C2({ S16509 }),
  .ZN({ S16510 })
);
NOR2_X1 #() 
NOR2_X1_519_ (
  .A1({ S25957[154] }),
  .A2({ S16338 }),
  .ZN({ S16511 })
);
AOI21_X1 #() 
AOI21_X1_1249_ (
  .A({ S16359 }),
  .B1({ S16511 }),
  .B2({ S25957[155] }),
  .ZN({ S16512 })
);
NAND2_X1 #() 
NAND2_X1_2176_ (
  .A1({ S16426 }),
  .A2({ S16386 }),
  .ZN({ S16513 })
);
AOI21_X1 #() 
AOI21_X1_1250_ (
  .A({ S54 }),
  .B1({ S16513 }),
  .B2({ S16392 }),
  .ZN({ S16514 })
);
INV_X1 #() 
INV_X1_705_ (
  .A({ S16514 }),
  .ZN({ S16515 })
);
AOI22_X1 #() 
AOI22_X1_278_ (
  .A1({ S16256 }),
  .A2({ S16253 }),
  .B1({ S16337 }),
  .B2({ S25957[153] }),
  .ZN({ S16517 })
);
NOR2_X1 #() 
NOR2_X1_520_ (
  .A1({ S16517 }),
  .A2({ S25957[155] }),
  .ZN({ S16518 })
);
AOI21_X1 #() 
AOI21_X1_1251_ (
  .A({ S25957[156] }),
  .B1({ S16518 }),
  .B2({ S16380 }),
  .ZN({ S16519 })
);
AOI22_X1 #() 
AOI22_X1_279_ (
  .A1({ S16515 }),
  .A2({ S16519 }),
  .B1({ S16512 }),
  .B2({ S16391 }),
  .ZN({ S16520 })
);
OAI21_X1 #() 
OAI21_X1_1154_ (
  .A({ S16510 }),
  .B1({ S25957[157] }),
  .B2({ S16520 }),
  .ZN({ S16521 })
);
NOR2_X1 #() 
NOR2_X1_521_ (
  .A1({ S16521 }),
  .A2({ S25957[158] }),
  .ZN({ S16522 })
);
NAND3_X1 #() 
NAND3_X1_2442_ (
  .A1({ S16383 }),
  .A2({ S25957[155] }),
  .A3({ S16335 }),
  .ZN({ S16523 })
);
OAI21_X1 #() 
OAI21_X1_1155_ (
  .A({ S54 }),
  .B1({ S16427 }),
  .B2({ S16412 }),
  .ZN({ S16524 })
);
AOI21_X1 #() 
AOI21_X1_1252_ (
  .A({ S25957[156] }),
  .B1({ S16524 }),
  .B2({ S16523 }),
  .ZN({ S16525 })
);
OAI211_X1 #() 
OAI211_X1_778_ (
  .A({ S16445 }),
  .B({ S25957[155] }),
  .C1({ S16426 }),
  .C2({ S16386 }),
  .ZN({ S16526 })
);
AND2_X1 #() 
AND2_X1_130_ (
  .A1({ S16397 }),
  .A2({ S25957[156] }),
  .ZN({ S16528 })
);
NAND2_X1 #() 
NAND2_X1_2177_ (
  .A1({ S16526 }),
  .A2({ S16528 }),
  .ZN({ S16529 })
);
AOI21_X1 #() 
AOI21_X1_1253_ (
  .A({ S16529 }),
  .B1({ S16413 }),
  .B2({ S25957[154] }),
  .ZN({ S16530 })
);
NOR3_X1 #() 
NOR3_X1_67_ (
  .A1({ S16530 }),
  .A2({ S16525 }),
  .A3({ S25957[157] }),
  .ZN({ S16531 })
);
NAND2_X1 #() 
NAND2_X1_2178_ (
  .A1({ S16417 }),
  .A2({ S54 }),
  .ZN({ S16532 })
);
AND2_X1 #() 
AND2_X1_131_ (
  .A1({ S16388 }),
  .A2({ S16532 }),
  .ZN({ S16533 })
);
NOR2_X1 #() 
NOR2_X1_522_ (
  .A1({ S16533 }),
  .A2({ S25957[156] }),
  .ZN({ S16534 })
);
AND4_X1 #() 
AND4_X1_6_ (
  .A1({ S54 }),
  .A2({ S16335 }),
  .A3({ S16339 }),
  .A4({ S16340 }),
  .ZN({ S16535 })
);
NAND3_X1 #() 
NAND3_X1_2443_ (
  .A1({ S16377 }),
  .A2({ S25957[155] }),
  .A3({ S25957[153] }),
  .ZN({ S16536 })
);
NAND2_X1 #() 
NAND2_X1_2179_ (
  .A1({ S16536 }),
  .A2({ S25957[156] }),
  .ZN({ S16537 })
);
OAI21_X1 #() 
OAI21_X1_1156_ (
  .A({ S25957[157] }),
  .B1({ S16537 }),
  .B2({ S16535 }),
  .ZN({ S16539 })
);
OAI21_X1 #() 
OAI21_X1_1157_ (
  .A({ S25957[158] }),
  .B1({ S16534 }),
  .B2({ S16539 }),
  .ZN({ S16540 })
);
NOR2_X1 #() 
NOR2_X1_523_ (
  .A1({ S16540 }),
  .A2({ S16531 }),
  .ZN({ S16541 })
);
OAI21_X1 #() 
OAI21_X1_1158_ (
  .A({ S25957[159] }),
  .B1({ S16522 }),
  .B2({ S16541 }),
  .ZN({ S16542 })
);
NAND2_X1 #() 
NAND2_X1_2180_ (
  .A1({ S16428 }),
  .A2({ S16360 }),
  .ZN({ S16543 })
);
NAND3_X1 #() 
NAND3_X1_2444_ (
  .A1({ S16543 }),
  .A2({ S25957[155] }),
  .A3({ S16383 }),
  .ZN({ S16544 })
);
NAND3_X1 #() 
NAND3_X1_2445_ (
  .A1({ S16507 }),
  .A2({ S54 }),
  .A3({ S16337 }),
  .ZN({ S16545 })
);
AND3_X1 #() 
AND3_X1_95_ (
  .A1({ S16544 }),
  .A2({ S25957[157] }),
  .A3({ S16545 }),
  .ZN({ S16546 })
);
NAND3_X1 #() 
NAND3_X1_2446_ (
  .A1({ S16383 }),
  .A2({ S16366 }),
  .A3({ S54 }),
  .ZN({ S16547 })
);
AOI21_X1 #() 
AOI21_X1_1254_ (
  .A({ S25957[153] }),
  .B1({ S16339 }),
  .B2({ S16340 }),
  .ZN({ S16548 })
);
OAI21_X1 #() 
OAI21_X1_1159_ (
  .A({ S25957[155] }),
  .B1({ S16517 }),
  .B2({ S16548 }),
  .ZN({ S16550 })
);
NAND3_X1 #() 
NAND3_X1_2447_ (
  .A1({ S16550 }),
  .A2({ S16376 }),
  .A3({ S16547 }),
  .ZN({ S16551 })
);
NAND2_X1 #() 
NAND2_X1_2181_ (
  .A1({ S16551 }),
  .A2({ S25957[156] }),
  .ZN({ S16552 })
);
NAND3_X1 #() 
NAND3_X1_2448_ (
  .A1({ S16370 }),
  .A2({ S16368 }),
  .A3({ S54 }),
  .ZN({ S16553 })
);
NAND2_X1 #() 
NAND2_X1_2182_ (
  .A1({ S16366 }),
  .A2({ S25957[155] }),
  .ZN({ S16554 })
);
OAI211_X1 #() 
OAI211_X1_779_ (
  .A({ S16553 }),
  .B({ S16359 }),
  .C1({ S25957[157] }),
  .C2({ S16554 }),
  .ZN({ S16555 })
);
OAI211_X1 #() 
OAI211_X1_780_ (
  .A({ S15729 }),
  .B({ S16555 }),
  .C1({ S16552 }),
  .C2({ S16546 }),
  .ZN({ S16556 })
);
AOI21_X1 #() 
AOI21_X1_1255_ (
  .A({ S54 }),
  .B1({ S25957[154] }),
  .B2({ S16489 }),
  .ZN({ S16557 })
);
NAND2_X1 #() 
NAND2_X1_2183_ (
  .A1({ S16557 }),
  .A2({ S16513 }),
  .ZN({ S16558 })
);
INV_X1 #() 
INV_X1_706_ (
  .A({ S16377 }),
  .ZN({ S16559 })
);
NOR2_X1 #() 
NOR2_X1_524_ (
  .A1({ S16559 }),
  .A2({ S25957[155] }),
  .ZN({ S16561 })
);
NAND2_X1 #() 
NAND2_X1_2184_ (
  .A1({ S25957[154] }),
  .A2({ S57 }),
  .ZN({ S16562 })
);
AOI21_X1 #() 
AOI21_X1_1256_ (
  .A({ S16359 }),
  .B1({ S16561 }),
  .B2({ S16562 }),
  .ZN({ S16563 })
);
NAND2_X1 #() 
NAND2_X1_2185_ (
  .A1({ S16344 }),
  .A2({ S16353 }),
  .ZN({ S16564 })
);
NAND2_X1 #() 
NAND2_X1_2186_ (
  .A1({ S16564 }),
  .A2({ S54 }),
  .ZN({ S16565 })
);
AOI21_X1 #() 
AOI21_X1_1257_ (
  .A({ S25957[156] }),
  .B1({ S16565 }),
  .B2({ S16550 }),
  .ZN({ S16566 })
);
AOI21_X1 #() 
AOI21_X1_1258_ (
  .A({ S16566 }),
  .B1({ S16563 }),
  .B2({ S16558 }),
  .ZN({ S16567 })
);
NAND3_X1 #() 
NAND3_X1_2449_ (
  .A1({ S16370 }),
  .A2({ S16344 }),
  .A3({ S54 }),
  .ZN({ S16568 })
);
AOI21_X1 #() 
AOI21_X1_1259_ (
  .A({ S16359 }),
  .B1({ S16388 }),
  .B2({ S16568 }),
  .ZN({ S16569 })
);
INV_X1 #() 
INV_X1_707_ (
  .A({ S16444 }),
  .ZN({ S16570 })
);
NAND2_X1 #() 
NAND2_X1_2187_ (
  .A1({ S16502 }),
  .A2({ S16392 }),
  .ZN({ S16572 })
);
AOI21_X1 #() 
AOI21_X1_1260_ (
  .A({ S25957[156] }),
  .B1({ S16572 }),
  .B2({ S16570 }),
  .ZN({ S16573 })
);
OAI21_X1 #() 
OAI21_X1_1160_ (
  .A({ S16376 }),
  .B1({ S16573 }),
  .B2({ S16569 }),
  .ZN({ S16574 })
);
OAI211_X1 #() 
OAI211_X1_781_ (
  .A({ S16574 }),
  .B({ S25957[158] }),
  .C1({ S16567 }),
  .C2({ S16376 }),
  .ZN({ S16575 })
);
NAND3_X1 #() 
NAND3_X1_2450_ (
  .A1({ S16575 }),
  .A2({ S15640 }),
  .A3({ S16556 }),
  .ZN({ S16576 })
);
NAND3_X1 #() 
NAND3_X1_2451_ (
  .A1({ S16542 }),
  .A2({ S16499 }),
  .A3({ S16576 }),
  .ZN({ S16577 })
);
NAND2_X1 #() 
NAND2_X1_2188_ (
  .A1({ S16575 }),
  .A2({ S16556 }),
  .ZN({ S16578 })
);
NAND2_X1 #() 
NAND2_X1_2189_ (
  .A1({ S16578 }),
  .A2({ S15640 }),
  .ZN({ S16579 })
);
OAI221_X1 #() 
OAI221_X1_46_ (
  .A({ S25957[159] }),
  .B1({ S16540 }),
  .B2({ S16531 }),
  .C1({ S16521 }),
  .C2({ S25957[158] }),
  .ZN({ S16580 })
);
NAND3_X1 #() 
NAND3_X1_2452_ (
  .A1({ S16580 }),
  .A2({ S16579 }),
  .A3({ S25957[225] }),
  .ZN({ S16581 })
);
NAND2_X1 #() 
NAND2_X1_2190_ (
  .A1({ S16577 }),
  .A2({ S16581 }),
  .ZN({ S25957[97] })
);
AOI21_X1 #() 
AOI21_X1_1261_ (
  .A({ S54 }),
  .B1({ S16428 }),
  .B2({ S16360 }),
  .ZN({ S16583 })
);
NOR2_X1 #() 
NOR2_X1_525_ (
  .A1({ S16583 }),
  .A2({ S16359 }),
  .ZN({ S16584 })
);
OAI21_X1 #() 
OAI21_X1_1161_ (
  .A({ S16584 }),
  .B1({ S25957[155] }),
  .B2({ S16511 }),
  .ZN({ S16585 })
);
AOI21_X1 #() 
AOI21_X1_1262_ (
  .A({ S25957[156] }),
  .B1({ S16449 }),
  .B2({ S54 }),
  .ZN({ S16586 })
);
AOI21_X1 #() 
AOI21_X1_1263_ (
  .A({ S25957[157] }),
  .B1({ S16586 }),
  .B2({ S16483 }),
  .ZN({ S16587 })
);
NAND2_X1 #() 
NAND2_X1_2191_ (
  .A1({ S16585 }),
  .A2({ S16587 }),
  .ZN({ S16588 })
);
NAND2_X1 #() 
NAND2_X1_2192_ (
  .A1({ S16562 }),
  .A2({ S54 }),
  .ZN({ S16589 })
);
OAI211_X1 #() 
OAI211_X1_782_ (
  .A({ S16359 }),
  .B({ S16589 }),
  .C1({ S16469 }),
  .C2({ S16406 }),
  .ZN({ S16590 })
);
NAND4_X1 #() 
NAND4_X1_304_ (
  .A1({ S16413 }),
  .A2({ S16340 }),
  .A3({ S16339 }),
  .A4({ S25957[152] }),
  .ZN({ S16591 })
);
OAI211_X1 #() 
OAI211_X1_783_ (
  .A({ S16591 }),
  .B({ S16410 }),
  .C1({ S16554 }),
  .C2({ S16337 }),
  .ZN({ S16593 })
);
OAI211_X1 #() 
OAI211_X1_784_ (
  .A({ S16590 }),
  .B({ S25957[157] }),
  .C1({ S16359 }),
  .C2({ S16593 }),
  .ZN({ S16594 })
);
AND2_X1 #() 
AND2_X1_132_ (
  .A1({ S16594 }),
  .A2({ S16588 }),
  .ZN({ S16595 })
);
INV_X1 #() 
INV_X1_708_ (
  .A({ S16435 }),
  .ZN({ S16596 })
);
NOR2_X1 #() 
NOR2_X1_526_ (
  .A1({ S54 }),
  .A2({ S25957[153] }),
  .ZN({ S16597 })
);
AOI21_X1 #() 
AOI21_X1_1264_ (
  .A({ S25957[156] }),
  .B1({ S16597 }),
  .B2({ S25957[152] }),
  .ZN({ S16598 })
);
OAI21_X1 #() 
OAI21_X1_1162_ (
  .A({ S16598 }),
  .B1({ S16596 }),
  .B2({ S16548 }),
  .ZN({ S16599 })
);
NOR2_X1 #() 
NOR2_X1_527_ (
  .A1({ S16469 }),
  .A2({ S16362 }),
  .ZN({ S16600 })
);
AOI21_X1 #() 
AOI21_X1_1265_ (
  .A({ S25957[155] }),
  .B1({ S16349 }),
  .B2({ S16338 }),
  .ZN({ S16601 })
);
OR2_X1 #() 
OR2_X1_30_ (
  .A1({ S16601 }),
  .A2({ S16359 }),
  .ZN({ S16602 })
);
OAI211_X1 #() 
OAI211_X1_785_ (
  .A({ S16376 }),
  .B({ S16599 }),
  .C1({ S16602 }),
  .C2({ S16600 }),
  .ZN({ S16604 })
);
NAND2_X1 #() 
NAND2_X1_2193_ (
  .A1({ S16417 }),
  .A2({ S25957[155] }),
  .ZN({ S16605 })
);
NOR2_X1 #() 
NOR2_X1_528_ (
  .A1({ S16605 }),
  .A2({ S16362 }),
  .ZN({ S16606 })
);
OAI21_X1 #() 
OAI21_X1_1163_ (
  .A({ S16359 }),
  .B1({ S16386 }),
  .B2({ S16398 }),
  .ZN({ S16607 })
);
NAND3_X1 #() 
NAND3_X1_2453_ (
  .A1({ S25957[154] }),
  .A2({ S25957[155] }),
  .A3({ S25957[152] }),
  .ZN({ S16608 })
);
NAND3_X1 #() 
NAND3_X1_2454_ (
  .A1({ S16512 }),
  .A2({ S16441 }),
  .A3({ S16608 }),
  .ZN({ S16609 })
);
OAI211_X1 #() 
OAI211_X1_786_ (
  .A({ S16609 }),
  .B({ S25957[157] }),
  .C1({ S16606 }),
  .C2({ S16607 }),
  .ZN({ S16610 })
);
NAND3_X1 #() 
NAND3_X1_2455_ (
  .A1({ S16610 }),
  .A2({ S16604 }),
  .A3({ S25957[158] }),
  .ZN({ S16611 })
);
OAI211_X1 #() 
OAI211_X1_787_ (
  .A({ S25957[159] }),
  .B({ S16611 }),
  .C1({ S16595 }),
  .C2({ S25957[158] }),
  .ZN({ S16612 })
);
INV_X1 #() 
INV_X1_709_ (
  .A({ S16365 }),
  .ZN({ S16613 })
);
OAI21_X1 #() 
OAI21_X1_1164_ (
  .A({ S54 }),
  .B1({ S16613 }),
  .B2({ S16511 }),
  .ZN({ S16614 })
);
OAI21_X1 #() 
OAI21_X1_1165_ (
  .A({ S16614 }),
  .B1({ S54 }),
  .B2({ S16564 }),
  .ZN({ S16615 })
);
NAND3_X1 #() 
NAND3_X1_2456_ (
  .A1({ S16387 }),
  .A2({ S25957[155] }),
  .A3({ S16370 }),
  .ZN({ S16616 })
);
AOI21_X1 #() 
AOI21_X1_1266_ (
  .A({ S16376 }),
  .B1({ S16586 }),
  .B2({ S16616 }),
  .ZN({ S16617 })
);
OAI21_X1 #() 
OAI21_X1_1166_ (
  .A({ S16617 }),
  .B1({ S16615 }),
  .B2({ S16359 }),
  .ZN({ S16618 })
);
NAND3_X1 #() 
NAND3_X1_2457_ (
  .A1({ S16441 }),
  .A2({ S16381 }),
  .A3({ S16359 }),
  .ZN({ S16619 })
);
AOI22_X1 #() 
AOI22_X1_280_ (
  .A1({ S16340 }),
  .A2({ S16339 }),
  .B1({ S25957[152] }),
  .B2({ S25957[153] }),
  .ZN({ S16620 })
);
OAI21_X1 #() 
OAI21_X1_1167_ (
  .A({ S54 }),
  .B1({ S16620 }),
  .B2({ S16517 }),
  .ZN({ S16621 })
);
NAND2_X1 #() 
NAND2_X1_2194_ (
  .A1({ S16584 }),
  .A2({ S16621 }),
  .ZN({ S16622 })
);
NAND3_X1 #() 
NAND3_X1_2458_ (
  .A1({ S16622 }),
  .A2({ S16376 }),
  .A3({ S16619 }),
  .ZN({ S16623 })
);
AND2_X1 #() 
AND2_X1_133_ (
  .A1({ S16618 }),
  .A2({ S16623 }),
  .ZN({ S16625 })
);
NAND2_X1 #() 
NAND2_X1_2195_ (
  .A1({ S16428 }),
  .A2({ S54 }),
  .ZN({ S16626 })
);
NAND3_X1 #() 
NAND3_X1_2459_ (
  .A1({ S16445 }),
  .A2({ S16383 }),
  .A3({ S25957[155] }),
  .ZN({ S16627 })
);
NAND3_X1 #() 
NAND3_X1_2460_ (
  .A1({ S16627 }),
  .A2({ S25957[156] }),
  .A3({ S16626 }),
  .ZN({ S16628 })
);
INV_X1 #() 
INV_X1_710_ (
  .A({ S16583 }),
  .ZN({ S16629 })
);
NAND3_X1 #() 
NAND3_X1_2461_ (
  .A1({ S16445 }),
  .A2({ S16446 }),
  .A3({ S54 }),
  .ZN({ S16630 })
);
NAND3_X1 #() 
NAND3_X1_2462_ (
  .A1({ S16629 }),
  .A2({ S16359 }),
  .A3({ S16630 }),
  .ZN({ S16631 })
);
NAND3_X1 #() 
NAND3_X1_2463_ (
  .A1({ S16343 }),
  .A2({ S16353 }),
  .A3({ S25957[156] }),
  .ZN({ S16632 })
);
NAND4_X1 #() 
NAND4_X1_305_ (
  .A1({ S16631 }),
  .A2({ S16632 }),
  .A3({ S16376 }),
  .A4({ S16628 }),
  .ZN({ S16633 })
);
NAND2_X1 #() 
NAND2_X1_2196_ (
  .A1({ S16427 }),
  .A2({ S25957[155] }),
  .ZN({ S16634 })
);
NAND2_X1 #() 
NAND2_X1_2197_ (
  .A1({ S16508 }),
  .A2({ S16353 }),
  .ZN({ S16636 })
);
NAND3_X1 #() 
NAND3_X1_2464_ (
  .A1({ S16634 }),
  .A2({ S16570 }),
  .A3({ S16636 }),
  .ZN({ S16637 })
);
NAND2_X1 #() 
NAND2_X1_2198_ (
  .A1({ S16637 }),
  .A2({ S16359 }),
  .ZN({ S16638 })
);
NOR3_X1 #() 
NOR3_X1_68_ (
  .A1({ S16548 }),
  .A2({ S16346 }),
  .A3({ S54 }),
  .ZN({ S16639 })
);
NAND2_X1 #() 
NAND2_X1_2199_ (
  .A1({ S16639 }),
  .A2({ S25957[156] }),
  .ZN({ S16640 })
);
NAND4_X1 #() 
NAND4_X1_306_ (
  .A1({ S16638 }),
  .A2({ S16640 }),
  .A3({ S25957[157] }),
  .A4({ S16632 }),
  .ZN({ S16641 })
);
NAND3_X1 #() 
NAND3_X1_2465_ (
  .A1({ S16641 }),
  .A2({ S25957[158] }),
  .A3({ S16633 }),
  .ZN({ S16642 })
);
OAI211_X1 #() 
OAI211_X1_788_ (
  .A({ S16642 }),
  .B({ S15640 }),
  .C1({ S16625 }),
  .C2({ S25957[158] }),
  .ZN({ S16643 })
);
NAND3_X1 #() 
NAND3_X1_2466_ (
  .A1({ S16643 }),
  .A2({ S25957[226] }),
  .A3({ S16612 }),
  .ZN({ S16644 })
);
INV_X1 #() 
INV_X1_711_ (
  .A({ S25957[226] }),
  .ZN({ S16645 })
);
AOI21_X1 #() 
AOI21_X1_1267_ (
  .A({ S25957[158] }),
  .B1({ S16618 }),
  .B2({ S16623 }),
  .ZN({ S16647 })
);
NAND3_X1 #() 
NAND3_X1_2467_ (
  .A1({ S16631 }),
  .A2({ S16628 }),
  .A3({ S16632 }),
  .ZN({ S16648 })
);
NAND2_X1 #() 
NAND2_X1_2200_ (
  .A1({ S16648 }),
  .A2({ S16376 }),
  .ZN({ S16649 })
);
INV_X1 #() 
INV_X1_712_ (
  .A({ S16343 }),
  .ZN({ S16650 })
);
INV_X1 #() 
INV_X1_713_ (
  .A({ S16353 }),
  .ZN({ S16651 })
);
OAI21_X1 #() 
OAI21_X1_1168_ (
  .A({ S25957[156] }),
  .B1({ S16650 }),
  .B2({ S16651 }),
  .ZN({ S16652 })
);
NAND4_X1 #() 
NAND4_X1_307_ (
  .A1({ S16634 }),
  .A2({ S16570 }),
  .A3({ S16359 }),
  .A4({ S16636 }),
  .ZN({ S16653 })
);
OAI211_X1 #() 
OAI211_X1_789_ (
  .A({ S16653 }),
  .B({ S25957[157] }),
  .C1({ S16652 }),
  .C2({ S16639 }),
  .ZN({ S16654 })
);
AOI21_X1 #() 
AOI21_X1_1268_ (
  .A({ S15729 }),
  .B1({ S16649 }),
  .B2({ S16654 }),
  .ZN({ S16655 })
);
OAI21_X1 #() 
OAI21_X1_1169_ (
  .A({ S15640 }),
  .B1({ S16655 }),
  .B2({ S16647 }),
  .ZN({ S16656 })
);
AOI21_X1 #() 
AOI21_X1_1269_ (
  .A({ S25957[158] }),
  .B1({ S16594 }),
  .B2({ S16588 }),
  .ZN({ S16658 })
);
AND3_X1 #() 
AND3_X1_96_ (
  .A1({ S16610 }),
  .A2({ S16604 }),
  .A3({ S25957[158] }),
  .ZN({ S16659 })
);
OAI21_X1 #() 
OAI21_X1_1170_ (
  .A({ S25957[159] }),
  .B1({ S16659 }),
  .B2({ S16658 }),
  .ZN({ S16660 })
);
NAND3_X1 #() 
NAND3_X1_2468_ (
  .A1({ S16656 }),
  .A2({ S16660 }),
  .A3({ S16645 }),
  .ZN({ S16661 })
);
NAND2_X1 #() 
NAND2_X1_2201_ (
  .A1({ S16644 }),
  .A2({ S16661 }),
  .ZN({ S25957[98] })
);
INV_X1 #() 
INV_X1_714_ (
  .A({ S25957[227] }),
  .ZN({ S16662 })
);
OAI211_X1 #() 
OAI211_X1_790_ (
  .A({ S25957[156] }),
  .B({ S16354 }),
  .C1({ S16532 }),
  .C2({ S16346 }),
  .ZN({ S16663 })
);
NAND3_X1 #() 
NAND3_X1_2469_ (
  .A1({ S16468 }),
  .A2({ S25957[155] }),
  .A3({ S16380 }),
  .ZN({ S16664 })
);
OAI211_X1 #() 
OAI211_X1_791_ (
  .A({ S16664 }),
  .B({ S16359 }),
  .C1({ S16650 }),
  .C2({ S16467 }),
  .ZN({ S16665 })
);
NAND3_X1 #() 
NAND3_X1_2470_ (
  .A1({ S16665 }),
  .A2({ S25957[157] }),
  .A3({ S16663 }),
  .ZN({ S16666 })
);
AOI21_X1 #() 
AOI21_X1_1270_ (
  .A({ S25957[155] }),
  .B1({ S16365 }),
  .B2({ S16368 }),
  .ZN({ S16668 })
);
NAND2_X1 #() 
NAND2_X1_2202_ (
  .A1({ S16353 }),
  .A2({ S16360 }),
  .ZN({ S16669 })
);
NOR2_X1 #() 
NOR2_X1_529_ (
  .A1({ S16596 }),
  .A2({ S25957[156] }),
  .ZN({ S16670 })
);
NAND2_X1 #() 
NAND2_X1_2203_ (
  .A1({ S16670 }),
  .A2({ S16669 }),
  .ZN({ S16671 })
);
OAI211_X1 #() 
OAI211_X1_792_ (
  .A({ S16671 }),
  .B({ S16376 }),
  .C1({ S16537 }),
  .C2({ S16668 }),
  .ZN({ S16672 })
);
AND3_X1 #() 
AND3_X1_97_ (
  .A1({ S16666 }),
  .A2({ S16672 }),
  .A3({ S25957[158] }),
  .ZN({ S16673 })
);
NAND2_X1 #() 
NAND2_X1_2204_ (
  .A1({ S16365 }),
  .A2({ S54 }),
  .ZN({ S16674 })
);
INV_X1 #() 
INV_X1_715_ (
  .A({ S16674 }),
  .ZN({ S16675 })
);
AOI21_X1 #() 
AOI21_X1_1271_ (
  .A({ S54 }),
  .B1({ S16543 }),
  .B2({ S16383 }),
  .ZN({ S16676 })
);
AOI21_X1 #() 
AOI21_X1_1272_ (
  .A({ S16676 }),
  .B1({ S16675 }),
  .B2({ S16507 }),
  .ZN({ S16677 })
);
NAND2_X1 #() 
NAND2_X1_2205_ (
  .A1({ S16677 }),
  .A2({ S16359 }),
  .ZN({ S16679 })
);
NOR2_X1 #() 
NOR2_X1_530_ (
  .A1({ S16411 }),
  .A2({ S16427 }),
  .ZN({ S16680 })
);
NAND2_X1 #() 
NAND2_X1_2206_ (
  .A1({ S16468 }),
  .A2({ S16377 }),
  .ZN({ S16681 })
);
NOR2_X1 #() 
NOR2_X1_531_ (
  .A1({ S16681 }),
  .A2({ S25957[155] }),
  .ZN({ S16682 })
);
OAI21_X1 #() 
OAI21_X1_1171_ (
  .A({ S25957[156] }),
  .B1({ S16682 }),
  .B2({ S16680 }),
  .ZN({ S16683 })
);
NAND3_X1 #() 
NAND3_X1_2471_ (
  .A1({ S16679 }),
  .A2({ S25957[157] }),
  .A3({ S16683 }),
  .ZN({ S16684 })
);
NAND2_X1 #() 
NAND2_X1_2207_ (
  .A1({ S16669 }),
  .A2({ S54 }),
  .ZN({ S16685 })
);
OAI21_X1 #() 
OAI21_X1_1172_ (
  .A({ S25957[155] }),
  .B1({ S16613 }),
  .B2({ S16548 }),
  .ZN({ S16686 })
);
AOI21_X1 #() 
AOI21_X1_1273_ (
  .A({ S25957[156] }),
  .B1({ S16686 }),
  .B2({ S16685 }),
  .ZN({ S16687 })
);
AOI21_X1 #() 
AOI21_X1_1274_ (
  .A({ S16359 }),
  .B1({ S16513 }),
  .B2({ S25957[155] }),
  .ZN({ S16688 })
);
NAND2_X1 #() 
NAND2_X1_2208_ (
  .A1({ S16688 }),
  .A2({ S16547 }),
  .ZN({ S16690 })
);
INV_X1 #() 
INV_X1_716_ (
  .A({ S16690 }),
  .ZN({ S16691 })
);
OAI21_X1 #() 
OAI21_X1_1173_ (
  .A({ S16376 }),
  .B1({ S16687 }),
  .B2({ S16691 }),
  .ZN({ S16692 })
);
AOI21_X1 #() 
AOI21_X1_1275_ (
  .A({ S25957[158] }),
  .B1({ S16684 }),
  .B2({ S16692 }),
  .ZN({ S16693 })
);
OAI21_X1 #() 
OAI21_X1_1174_ (
  .A({ S25957[159] }),
  .B1({ S16693 }),
  .B2({ S16673 }),
  .ZN({ S16694 })
);
AOI21_X1 #() 
AOI21_X1_1276_ (
  .A({ S25957[155] }),
  .B1({ S16387 }),
  .B2({ S16365 }),
  .ZN({ S16695 })
);
NAND2_X1 #() 
NAND2_X1_2209_ (
  .A1({ S16347 }),
  .A2({ S16377 }),
  .ZN({ S16696 })
);
NAND2_X1 #() 
NAND2_X1_2210_ (
  .A1({ S16696 }),
  .A2({ S25957[156] }),
  .ZN({ S16697 })
);
NAND2_X1 #() 
NAND2_X1_2211_ (
  .A1({ S16507 }),
  .A2({ S16508 }),
  .ZN({ S16698 })
);
NAND2_X1 #() 
NAND2_X1_2212_ (
  .A1({ S16424 }),
  .A2({ S16698 }),
  .ZN({ S16699 })
);
OAI21_X1 #() 
OAI21_X1_1175_ (
  .A({ S16699 }),
  .B1({ S16697 }),
  .B2({ S16695 }),
  .ZN({ S16701 })
);
INV_X1 #() 
INV_X1_717_ (
  .A({ S16438 }),
  .ZN({ S16702 })
);
NAND3_X1 #() 
NAND3_X1_2472_ (
  .A1({ S16410 }),
  .A2({ S16359 }),
  .A3({ S16591 }),
  .ZN({ S16703 })
);
OAI21_X1 #() 
OAI21_X1_1176_ (
  .A({ S16652 }),
  .B1({ S16702 }),
  .B2({ S16703 }),
  .ZN({ S16704 })
);
OR2_X1 #() 
OR2_X1_31_ (
  .A1({ S16704 }),
  .A2({ S25957[157] }),
  .ZN({ S16705 })
);
OAI211_X1 #() 
OAI211_X1_793_ (
  .A({ S16705 }),
  .B({ S25957[158] }),
  .C1({ S16376 }),
  .C2({ S16701 }),
  .ZN({ S16706 })
);
NAND2_X1 #() 
NAND2_X1_2213_ (
  .A1({ S16469 }),
  .A2({ S16636 }),
  .ZN({ S16707 })
);
NAND2_X1 #() 
NAND2_X1_2214_ (
  .A1({ S16707 }),
  .A2({ S16359 }),
  .ZN({ S16708 })
);
NAND3_X1 #() 
NAND3_X1_2473_ (
  .A1({ S16591 }),
  .A2({ S25957[156] }),
  .A3({ S16342 }),
  .ZN({ S16709 })
);
AND2_X1 #() 
AND2_X1_134_ (
  .A1({ S16708 }),
  .A2({ S16709 }),
  .ZN({ S16710 })
);
NAND3_X1 #() 
NAND3_X1_2474_ (
  .A1({ S16491 }),
  .A2({ S16379 }),
  .A3({ S54 }),
  .ZN({ S16712 })
);
AND2_X1 #() 
AND2_X1_135_ (
  .A1({ S16558 }),
  .A2({ S16712 }),
  .ZN({ S16713 })
);
AOI21_X1 #() 
AOI21_X1_1277_ (
  .A({ S25957[155] }),
  .B1({ S16365 }),
  .B2({ S16377 }),
  .ZN({ S16714 })
);
AOI21_X1 #() 
AOI21_X1_1278_ (
  .A({ S54 }),
  .B1({ S16387 }),
  .B2({ S16353 }),
  .ZN({ S16715 })
);
OAI21_X1 #() 
OAI21_X1_1177_ (
  .A({ S16359 }),
  .B1({ S16715 }),
  .B2({ S16714 }),
  .ZN({ S16716 })
);
OAI21_X1 #() 
OAI21_X1_1178_ (
  .A({ S16716 }),
  .B1({ S16713 }),
  .B2({ S16359 }),
  .ZN({ S16717 })
);
NAND2_X1 #() 
NAND2_X1_2215_ (
  .A1({ S16717 }),
  .A2({ S16376 }),
  .ZN({ S16718 })
);
OAI211_X1 #() 
OAI211_X1_794_ (
  .A({ S16718 }),
  .B({ S15729 }),
  .C1({ S16376 }),
  .C2({ S16710 }),
  .ZN({ S16719 })
);
NAND3_X1 #() 
NAND3_X1_2475_ (
  .A1({ S16719 }),
  .A2({ S16706 }),
  .A3({ S15640 }),
  .ZN({ S16720 })
);
NAND3_X1 #() 
NAND3_X1_2476_ (
  .A1({ S16694 }),
  .A2({ S16720 }),
  .A3({ S16662 }),
  .ZN({ S16721 })
);
OAI211_X1 #() 
OAI211_X1_795_ (
  .A({ S25957[158] }),
  .B({ S16671 }),
  .C1({ S16668 }),
  .C2({ S16537 }),
  .ZN({ S16723 })
);
NAND2_X1 #() 
NAND2_X1_2216_ (
  .A1({ S16690 }),
  .A2({ S15729 }),
  .ZN({ S16724 })
);
OR2_X1 #() 
OR2_X1_32_ (
  .A1({ S16724 }),
  .A2({ S16687 }),
  .ZN({ S16725 })
);
AOI21_X1 #() 
AOI21_X1_1279_ (
  .A({ S15640 }),
  .B1({ S16725 }),
  .B2({ S16723 }),
  .ZN({ S16726 })
);
OAI211_X1 #() 
OAI211_X1_796_ (
  .A({ S15729 }),
  .B({ S16716 }),
  .C1({ S16713 }),
  .C2({ S16359 }),
  .ZN({ S16727 })
);
NAND2_X1 #() 
NAND2_X1_2217_ (
  .A1({ S16704 }),
  .A2({ S25957[158] }),
  .ZN({ S16728 })
);
AOI21_X1 #() 
AOI21_X1_1280_ (
  .A({ S25957[159] }),
  .B1({ S16727 }),
  .B2({ S16728 }),
  .ZN({ S16729 })
);
OAI21_X1 #() 
OAI21_X1_1179_ (
  .A({ S16376 }),
  .B1({ S16726 }),
  .B2({ S16729 }),
  .ZN({ S16730 })
);
NAND2_X1 #() 
NAND2_X1_2218_ (
  .A1({ S16701 }),
  .A2({ S25957[158] }),
  .ZN({ S16731 })
);
NAND3_X1 #() 
NAND3_X1_2477_ (
  .A1({ S16708 }),
  .A2({ S15729 }),
  .A3({ S16709 }),
  .ZN({ S16732 })
);
AOI21_X1 #() 
AOI21_X1_1281_ (
  .A({ S25957[159] }),
  .B1({ S16731 }),
  .B2({ S16732 }),
  .ZN({ S16734 })
);
NAND3_X1 #() 
NAND3_X1_2478_ (
  .A1({ S16665 }),
  .A2({ S25957[158] }),
  .A3({ S16663 }),
  .ZN({ S16735 })
);
OAI221_X1 #() 
OAI221_X1_47_ (
  .A({ S25957[156] }),
  .B1({ S16411 }),
  .B2({ S16427 }),
  .C1({ S16681 }),
  .C2({ S25957[155] }),
  .ZN({ S16736 })
);
OAI211_X1 #() 
OAI211_X1_797_ (
  .A({ S16736 }),
  .B({ S15729 }),
  .C1({ S16677 }),
  .C2({ S25957[156] }),
  .ZN({ S16737 })
);
AOI21_X1 #() 
AOI21_X1_1282_ (
  .A({ S15640 }),
  .B1({ S16737 }),
  .B2({ S16735 }),
  .ZN({ S16738 })
);
OAI21_X1 #() 
OAI21_X1_1180_ (
  .A({ S25957[157] }),
  .B1({ S16738 }),
  .B2({ S16734 }),
  .ZN({ S16739 })
);
NAND3_X1 #() 
NAND3_X1_2479_ (
  .A1({ S16730 }),
  .A2({ S16739 }),
  .A3({ S25957[227] }),
  .ZN({ S16740 })
);
NAND2_X1 #() 
NAND2_X1_2219_ (
  .A1({ S16721 }),
  .A2({ S16740 }),
  .ZN({ S25957[99] })
);
NOR2_X1 #() 
NOR2_X1_532_ (
  .A1({ S16532 }),
  .A2({ S16362 }),
  .ZN({ S16741 })
);
AND2_X1 #() 
AND2_X1_136_ (
  .A1({ S16386 }),
  .A2({ S152 }),
  .ZN({ S16742 })
);
OAI22_X1 #() 
OAI22_X1_52_ (
  .A1({ S16741 }),
  .A2({ S16452 }),
  .B1({ S16359 }),
  .B2({ S16742 }),
  .ZN({ S16744 })
);
AOI21_X1 #() 
AOI21_X1_1283_ (
  .A({ S25957[155] }),
  .B1({ S16507 }),
  .B2({ S16342 }),
  .ZN({ S16745 })
);
NAND2_X1 #() 
NAND2_X1_2220_ (
  .A1({ S16550 }),
  .A2({ S25957[156] }),
  .ZN({ S16746 })
);
NAND2_X1 #() 
NAND2_X1_2221_ (
  .A1({ S16386 }),
  .A2({ S55 }),
  .ZN({ S16747 })
);
NAND3_X1 #() 
NAND3_X1_2480_ (
  .A1({ S16747 }),
  .A2({ S54 }),
  .A3({ S16383 }),
  .ZN({ S16748 })
);
AOI21_X1 #() 
AOI21_X1_1284_ (
  .A({ S25957[157] }),
  .B1({ S16670 }),
  .B2({ S16748 }),
  .ZN({ S16749 })
);
OAI21_X1 #() 
OAI21_X1_1181_ (
  .A({ S16749 }),
  .B1({ S16746 }),
  .B2({ S16745 }),
  .ZN({ S16750 })
);
OAI21_X1 #() 
OAI21_X1_1182_ (
  .A({ S16750 }),
  .B1({ S16376 }),
  .B2({ S16744 }),
  .ZN({ S16751 })
);
NOR2_X1 #() 
NOR2_X1_533_ (
  .A1({ S16434 }),
  .A2({ S16607 }),
  .ZN({ S16752 })
);
NAND2_X1 #() 
NAND2_X1_2222_ (
  .A1({ S16752 }),
  .A2({ S16354 }),
  .ZN({ S16753 })
);
INV_X1 #() 
INV_X1_718_ (
  .A({ S16379 }),
  .ZN({ S16755 })
);
OAI211_X1 #() 
OAI211_X1_798_ (
  .A({ S16438 }),
  .B({ S25957[156] }),
  .C1({ S16755 }),
  .C2({ S16650 }),
  .ZN({ S16756 })
);
NAND2_X1 #() 
NAND2_X1_2223_ (
  .A1({ S16753 }),
  .A2({ S16756 }),
  .ZN({ S16757 })
);
AOI21_X1 #() 
AOI21_X1_1285_ (
  .A({ S54 }),
  .B1({ S16491 }),
  .B2({ S16379 }),
  .ZN({ S16758 })
);
OAI21_X1 #() 
OAI21_X1_1183_ (
  .A({ S25957[156] }),
  .B1({ S16758 }),
  .B2({ S16518 }),
  .ZN({ S16759 })
);
AOI21_X1 #() 
AOI21_X1_1286_ (
  .A({ S54 }),
  .B1({ S16361 }),
  .B2({ S16386 }),
  .ZN({ S16760 })
);
NAND2_X1 #() 
NAND2_X1_2224_ (
  .A1({ S16650 }),
  .A2({ S16359 }),
  .ZN({ S16761 })
);
OAI21_X1 #() 
OAI21_X1_1184_ (
  .A({ S16759 }),
  .B1({ S16760 }),
  .B2({ S16761 }),
  .ZN({ S16762 })
);
NAND2_X1 #() 
NAND2_X1_2225_ (
  .A1({ S16762 }),
  .A2({ S25957[157] }),
  .ZN({ S16763 })
);
OAI211_X1 #() 
OAI211_X1_799_ (
  .A({ S16763 }),
  .B({ S15729 }),
  .C1({ S25957[157] }),
  .C2({ S16757 }),
  .ZN({ S16764 })
);
OAI211_X1 #() 
OAI211_X1_800_ (
  .A({ S16764 }),
  .B({ S15640 }),
  .C1({ S15729 }),
  .C2({ S16751 }),
  .ZN({ S16766 })
);
NAND3_X1 #() 
NAND3_X1_2481_ (
  .A1({ S16405 }),
  .A2({ S25957[156] }),
  .A3({ S16491 }),
  .ZN({ S16767 })
);
NOR2_X1 #() 
NOR2_X1_534_ (
  .A1({ S16548 }),
  .A2({ S54 }),
  .ZN({ S16768 })
);
NAND2_X1 #() 
NAND2_X1_2226_ (
  .A1({ S16768 }),
  .A2({ S16353 }),
  .ZN({ S16769 })
);
NAND3_X1 #() 
NAND3_X1_2482_ (
  .A1({ S16769 }),
  .A2({ S16359 }),
  .A3({ S16545 }),
  .ZN({ S16770 })
);
NAND3_X1 #() 
NAND3_X1_2483_ (
  .A1({ S16770 }),
  .A2({ S25957[157] }),
  .A3({ S16767 }),
  .ZN({ S16771 })
);
NAND2_X1 #() 
NAND2_X1_2227_ (
  .A1({ S16360 }),
  .A2({ S54 }),
  .ZN({ S16772 })
);
NAND2_X1 #() 
NAND2_X1_2228_ (
  .A1({ S25957[155] }),
  .A2({ S16338 }),
  .ZN({ S16773 })
);
OAI221_X1 #() 
OAI221_X1_48_ (
  .A({ S25957[156] }),
  .B1({ S16501 }),
  .B2({ S16773 }),
  .C1({ S16548 }),
  .C2({ S16772 }),
  .ZN({ S16774 })
);
AOI21_X1 #() 
AOI21_X1_1287_ (
  .A({ S54 }),
  .B1({ S16428 }),
  .B2({ S57 }),
  .ZN({ S16775 })
);
NOR2_X1 #() 
NOR2_X1_535_ (
  .A1({ S16775 }),
  .A2({ S25957[156] }),
  .ZN({ S16777 })
);
NAND2_X1 #() 
NAND2_X1_2229_ (
  .A1({ S16777 }),
  .A2({ S16547 }),
  .ZN({ S16778 })
);
NAND3_X1 #() 
NAND3_X1_2484_ (
  .A1({ S16778 }),
  .A2({ S16376 }),
  .A3({ S16774 }),
  .ZN({ S16779 })
);
NAND2_X1 #() 
NAND2_X1_2230_ (
  .A1({ S16771 }),
  .A2({ S16779 }),
  .ZN({ S16780 })
);
NAND2_X1 #() 
NAND2_X1_2231_ (
  .A1({ S16780 }),
  .A2({ S25957[158] }),
  .ZN({ S16781 })
);
NOR2_X1 #() 
NOR2_X1_536_ (
  .A1({ S16492 }),
  .A2({ S25957[156] }),
  .ZN({ S16782 })
);
AOI21_X1 #() 
AOI21_X1_1288_ (
  .A({ S16447 }),
  .B1({ S16439 }),
  .B2({ S16347 }),
  .ZN({ S16783 })
);
NAND2_X1 #() 
NAND2_X1_2232_ (
  .A1({ S16513 }),
  .A2({ S16392 }),
  .ZN({ S16784 })
);
NAND2_X1 #() 
NAND2_X1_2233_ (
  .A1({ S16784 }),
  .A2({ S54 }),
  .ZN({ S16785 })
);
AOI22_X1 #() 
AOI22_X1_281_ (
  .A1({ S16783 }),
  .A2({ S25957[156] }),
  .B1({ S16785 }),
  .B2({ S16782 }),
  .ZN({ S16786 })
);
NAND2_X1 #() 
NAND2_X1_2234_ (
  .A1({ S16391 }),
  .A2({ S16773 }),
  .ZN({ S16788 })
);
NAND3_X1 #() 
NAND3_X1_2485_ (
  .A1({ S16788 }),
  .A2({ S16359 }),
  .A3({ S16353 }),
  .ZN({ S16789 })
);
NAND3_X1 #() 
NAND3_X1_2486_ (
  .A1({ S16387 }),
  .A2({ S16503 }),
  .A3({ S54 }),
  .ZN({ S16790 })
);
OAI211_X1 #() 
OAI211_X1_801_ (
  .A({ S16790 }),
  .B({ S25957[156] }),
  .C1({ S16548 }),
  .C2({ S16605 }),
  .ZN({ S16791 })
);
AOI21_X1 #() 
AOI21_X1_1289_ (
  .A({ S25957[157] }),
  .B1({ S16791 }),
  .B2({ S16789 }),
  .ZN({ S16792 })
);
AOI21_X1 #() 
AOI21_X1_1290_ (
  .A({ S16792 }),
  .B1({ S16786 }),
  .B2({ S25957[157] }),
  .ZN({ S16793 })
);
OAI21_X1 #() 
OAI21_X1_1185_ (
  .A({ S16781 }),
  .B1({ S16793 }),
  .B2({ S25957[158] }),
  .ZN({ S16794 })
);
NAND2_X1 #() 
NAND2_X1_2235_ (
  .A1({ S16794 }),
  .A2({ S25957[159] }),
  .ZN({ S16795 })
);
NAND2_X1 #() 
NAND2_X1_2236_ (
  .A1({ S16795 }),
  .A2({ S16766 }),
  .ZN({ S16796 })
);
XNOR2_X1 #() 
XNOR2_X1_125_ (
  .A({ S16796 }),
  .B({ S25957[228] }),
  .ZN({ S25957[100] })
);
AOI21_X1 #() 
AOI21_X1_1291_ (
  .A({ S25957[155] }),
  .B1({ S16383 }),
  .B2({ S16345 }),
  .ZN({ S16798 })
);
AOI21_X1 #() 
AOI21_X1_1292_ (
  .A({ S54 }),
  .B1({ S16370 }),
  .B2({ S16368 }),
  .ZN({ S16799 })
);
OAI21_X1 #() 
OAI21_X1_1186_ (
  .A({ S25957[156] }),
  .B1({ S16799 }),
  .B2({ S16798 }),
  .ZN({ S16800 })
);
OAI21_X1 #() 
OAI21_X1_1187_ (
  .A({ S16773 }),
  .B1({ S16548 }),
  .B2({ S16772 }),
  .ZN({ S16801 })
);
NAND2_X1 #() 
NAND2_X1_2237_ (
  .A1({ S16801 }),
  .A2({ S16359 }),
  .ZN({ S16802 })
);
NAND3_X1 #() 
NAND3_X1_2487_ (
  .A1({ S16800 }),
  .A2({ S25957[157] }),
  .A3({ S16802 }),
  .ZN({ S16803 })
);
OAI21_X1 #() 
OAI21_X1_1188_ (
  .A({ S25957[156] }),
  .B1({ S16601 }),
  .B2({ S16760 }),
  .ZN({ S16804 })
);
OAI211_X1 #() 
OAI211_X1_802_ (
  .A({ S16344 }),
  .B({ S25957[155] }),
  .C1({ S16426 }),
  .C2({ S16386 }),
  .ZN({ S16805 })
);
AOI21_X1 #() 
AOI21_X1_1293_ (
  .A({ S25957[156] }),
  .B1({ S16501 }),
  .B2({ S16413 }),
  .ZN({ S16806 })
);
NAND2_X1 #() 
NAND2_X1_2238_ (
  .A1({ S16805 }),
  .A2({ S16806 }),
  .ZN({ S16807 })
);
NAND3_X1 #() 
NAND3_X1_2488_ (
  .A1({ S16804 }),
  .A2({ S16376 }),
  .A3({ S16807 }),
  .ZN({ S16809 })
);
AOI21_X1 #() 
AOI21_X1_1294_ (
  .A({ S25957[158] }),
  .B1({ S16803 }),
  .B2({ S16809 }),
  .ZN({ S16810 })
);
AOI21_X1 #() 
AOI21_X1_1295_ (
  .A({ S16359 }),
  .B1({ S16412 }),
  .B2({ S16413 }),
  .ZN({ S16811 })
);
AOI21_X1 #() 
AOI21_X1_1296_ (
  .A({ S54 }),
  .B1({ S16337 }),
  .B2({ S25957[153] }),
  .ZN({ S16812 })
);
AOI22_X1 #() 
AOI22_X1_282_ (
  .A1({ S16812 }),
  .A2({ S16383 }),
  .B1({ S16508 }),
  .B2({ S16386 }),
  .ZN({ S16813 })
);
NAND2_X1 #() 
NAND2_X1_2239_ (
  .A1({ S16813 }),
  .A2({ S16811 }),
  .ZN({ S16814 })
);
OAI21_X1 #() 
OAI21_X1_1189_ (
  .A({ S25957[155] }),
  .B1({ S16620 }),
  .B2({ S16517 }),
  .ZN({ S16815 })
);
AOI21_X1 #() 
AOI21_X1_1297_ (
  .A({ S16376 }),
  .B1({ S16400 }),
  .B2({ S16815 }),
  .ZN({ S16816 })
);
AND2_X1 #() 
AND2_X1_137_ (
  .A1({ S16816 }),
  .A2({ S16814 }),
  .ZN({ S16817 })
);
NAND4_X1 #() 
NAND4_X1_308_ (
  .A1({ S16383 }),
  .A2({ S16349 }),
  .A3({ S25957[155] }),
  .A4({ S16335 }),
  .ZN({ S16818 })
);
AOI21_X1 #() 
AOI21_X1_1298_ (
  .A({ S25957[156] }),
  .B1({ S16365 }),
  .B2({ S54 }),
  .ZN({ S16820 })
);
NAND2_X1 #() 
NAND2_X1_2240_ (
  .A1({ S16406 }),
  .A2({ S54 }),
  .ZN({ S16821 })
);
AOI21_X1 #() 
AOI21_X1_1299_ (
  .A({ S16359 }),
  .B1({ S16386 }),
  .B2({ S16360 }),
  .ZN({ S16822 })
);
AOI22_X1 #() 
AOI22_X1_283_ (
  .A1({ S16820 }),
  .A2({ S16818 }),
  .B1({ S16821 }),
  .B2({ S16822 }),
  .ZN({ S16823 })
);
OAI21_X1 #() 
OAI21_X1_1190_ (
  .A({ S25957[158] }),
  .B1({ S16823 }),
  .B2({ S25957[157] }),
  .ZN({ S16824 })
);
OAI21_X1 #() 
OAI21_X1_1191_ (
  .A({ S25957[159] }),
  .B1({ S16817 }),
  .B2({ S16824 }),
  .ZN({ S16825 })
);
NAND3_X1 #() 
NAND3_X1_2489_ (
  .A1({ S16368 }),
  .A2({ S54 }),
  .A3({ S16428 }),
  .ZN({ S16826 })
);
NAND3_X1 #() 
NAND3_X1_2490_ (
  .A1({ S16526 }),
  .A2({ S25957[156] }),
  .A3({ S16826 }),
  .ZN({ S16827 })
);
INV_X1 #() 
INV_X1_719_ (
  .A({ S16422 }),
  .ZN({ S16828 })
);
AOI21_X1 #() 
AOI21_X1_1300_ (
  .A({ S16376 }),
  .B1({ S16828 }),
  .B2({ S16351 }),
  .ZN({ S16829 })
);
NAND2_X1 #() 
NAND2_X1_2241_ (
  .A1({ S16827 }),
  .A2({ S16829 }),
  .ZN({ S16831 })
);
AOI21_X1 #() 
AOI21_X1_1301_ (
  .A({ S25957[155] }),
  .B1({ S16445 }),
  .B2({ S16383 }),
  .ZN({ S16832 })
);
AOI22_X1 #() 
AOI22_X1_284_ (
  .A1({ S16335 }),
  .A2({ S54 }),
  .B1({ S16339 }),
  .B2({ S16340 }),
  .ZN({ S16833 })
);
AOI21_X1 #() 
AOI21_X1_1302_ (
  .A({ S16359 }),
  .B1({ S16597 }),
  .B2({ S25957[152] }),
  .ZN({ S16834 })
);
OAI21_X1 #() 
OAI21_X1_1192_ (
  .A({ S16834 }),
  .B1({ S16535 }),
  .B2({ S16833 }),
  .ZN({ S16835 })
);
OAI211_X1 #() 
OAI211_X1_803_ (
  .A({ S16835 }),
  .B({ S16376 }),
  .C1({ S16452 }),
  .C2({ S16832 }),
  .ZN({ S16836 })
);
NAND3_X1 #() 
NAND3_X1_2491_ (
  .A1({ S16836 }),
  .A2({ S16831 }),
  .A3({ S25957[158] }),
  .ZN({ S16837 })
);
AOI21_X1 #() 
AOI21_X1_1303_ (
  .A({ S54 }),
  .B1({ S16365 }),
  .B2({ S16368 }),
  .ZN({ S16838 })
);
NAND2_X1 #() 
NAND2_X1_2242_ (
  .A1({ S16466 }),
  .A2({ S25957[156] }),
  .ZN({ S16839 })
);
AOI21_X1 #() 
AOI21_X1_1304_ (
  .A({ S25957[157] }),
  .B1({ S16598 }),
  .B2({ S16591 }),
  .ZN({ S16840 })
);
OAI21_X1 #() 
OAI21_X1_1193_ (
  .A({ S16840 }),
  .B1({ S16839 }),
  .B2({ S16838 }),
  .ZN({ S16842 })
);
NAND2_X1 #() 
NAND2_X1_2243_ (
  .A1({ S16608 }),
  .A2({ S16359 }),
  .ZN({ S16843 })
);
AOI21_X1 #() 
AOI21_X1_1305_ (
  .A({ S16398 }),
  .B1({ S16353 }),
  .B2({ S16377 }),
  .ZN({ S16844 })
);
NAND4_X1 #() 
NAND4_X1_309_ (
  .A1({ S16335 }),
  .A2({ S16256 }),
  .A3({ S16253 }),
  .A4({ S25957[155] }),
  .ZN({ S16845 })
);
OAI211_X1 #() 
OAI211_X1_804_ (
  .A({ S25957[156] }),
  .B({ S16845 }),
  .C1({ S16449 }),
  .C2({ S25957[155] }),
  .ZN({ S16846 })
);
OAI211_X1 #() 
OAI211_X1_805_ (
  .A({ S16846 }),
  .B({ S25957[157] }),
  .C1({ S16843 }),
  .C2({ S16844 }),
  .ZN({ S16847 })
);
NAND3_X1 #() 
NAND3_X1_2492_ (
  .A1({ S16847 }),
  .A2({ S16842 }),
  .A3({ S15729 }),
  .ZN({ S16848 })
);
NAND3_X1 #() 
NAND3_X1_2493_ (
  .A1({ S16837 }),
  .A2({ S16848 }),
  .A3({ S15640 }),
  .ZN({ S16849 })
);
OAI211_X1 #() 
OAI211_X1_806_ (
  .A({ S16849 }),
  .B({ S16285 }),
  .C1({ S16825 }),
  .C2({ S16810 }),
  .ZN({ S16850 })
);
NAND2_X1 #() 
NAND2_X1_2244_ (
  .A1({ S16820 }),
  .A2({ S16818 }),
  .ZN({ S16851 })
);
AOI21_X1 #() 
AOI21_X1_1306_ (
  .A({ S25957[157] }),
  .B1({ S16822 }),
  .B2({ S16821 }),
  .ZN({ S16853 })
);
NAND2_X1 #() 
NAND2_X1_2245_ (
  .A1({ S16851 }),
  .A2({ S16853 }),
  .ZN({ S16854 })
);
AOI22_X1 #() 
AOI22_X1_285_ (
  .A1({ S16400 }),
  .A2({ S16815 }),
  .B1({ S16813 }),
  .B2({ S16811 }),
  .ZN({ S16855 })
);
OAI211_X1 #() 
OAI211_X1_807_ (
  .A({ S25957[158] }),
  .B({ S16854 }),
  .C1({ S16855 }),
  .C2({ S16376 }),
  .ZN({ S16856 })
);
NAND3_X1 #() 
NAND3_X1_2494_ (
  .A1({ S16803 }),
  .A2({ S15729 }),
  .A3({ S16809 }),
  .ZN({ S16857 })
);
AOI21_X1 #() 
AOI21_X1_1307_ (
  .A({ S15640 }),
  .B1({ S16857 }),
  .B2({ S16856 }),
  .ZN({ S16858 })
);
AND3_X1 #() 
AND3_X1_98_ (
  .A1({ S16837 }),
  .A2({ S15640 }),
  .A3({ S16848 }),
  .ZN({ S16859 })
);
OAI21_X1 #() 
OAI21_X1_1194_ (
  .A({ S25957[229] }),
  .B1({ S16858 }),
  .B2({ S16859 }),
  .ZN({ S16860 })
);
NAND2_X1 #() 
NAND2_X1_2246_ (
  .A1({ S16860 }),
  .A2({ S16850 }),
  .ZN({ S25957[101] })
);
AND2_X1 #() 
AND2_X1_138_ (
  .A1({ S16366 }),
  .A2({ S16428 }),
  .ZN({ S16861 })
);
OAI211_X1 #() 
OAI211_X1_808_ (
  .A({ S16359 }),
  .B({ S16826 }),
  .C1({ S16861 }),
  .C2({ S54 }),
  .ZN({ S16863 })
);
NAND2_X1 #() 
NAND2_X1_2247_ (
  .A1({ S16421 }),
  .A2({ S16773 }),
  .ZN({ S16864 })
);
AND2_X1 #() 
AND2_X1_139_ (
  .A1({ S16864 }),
  .A2({ S16342 }),
  .ZN({ S16865 })
);
OAI21_X1 #() 
OAI21_X1_1195_ (
  .A({ S25957[156] }),
  .B1({ S16501 }),
  .B2({ S25957[155] }),
  .ZN({ S16866 })
);
OAI211_X1 #() 
OAI211_X1_809_ (
  .A({ S16863 }),
  .B({ S25957[157] }),
  .C1({ S16865 }),
  .C2({ S16866 }),
  .ZN({ S16867 })
);
NAND2_X1 #() 
NAND2_X1_2248_ (
  .A1({ S16381 }),
  .A2({ S16359 }),
  .ZN({ S16868 })
);
NAND2_X1 #() 
NAND2_X1_2249_ (
  .A1({ S16410 }),
  .A2({ S25957[156] }),
  .ZN({ S16869 })
);
OAI211_X1 #() 
OAI211_X1_810_ (
  .A({ S16868 }),
  .B({ S16376 }),
  .C1({ S16869 }),
  .C2({ S16758 }),
  .ZN({ S16870 })
);
AOI21_X1 #() 
AOI21_X1_1308_ (
  .A({ S25957[158] }),
  .B1({ S16867 }),
  .B2({ S16870 }),
  .ZN({ S16871 })
);
NAND3_X1 #() 
NAND3_X1_2495_ (
  .A1({ S16370 }),
  .A2({ S54 }),
  .A3({ S16377 }),
  .ZN({ S16872 })
);
OAI211_X1 #() 
OAI211_X1_811_ (
  .A({ S16872 }),
  .B({ S25957[156] }),
  .C1({ S54 }),
  .C2({ S16669 }),
  .ZN({ S16874 })
);
OAI211_X1 #() 
OAI211_X1_812_ (
  .A({ S16874 }),
  .B({ S25957[157] }),
  .C1({ S16543 }),
  .C2({ S16843 }),
  .ZN({ S16875 })
);
AND3_X1 #() 
AND3_X1_99_ (
  .A1({ S16528 }),
  .A2({ S16366 }),
  .A3({ S16435 }),
  .ZN({ S16876 })
);
OAI21_X1 #() 
OAI21_X1_1196_ (
  .A({ S54 }),
  .B1({ S16426 }),
  .B2({ S16386 }),
  .ZN({ S16877 })
);
AOI21_X1 #() 
AOI21_X1_1309_ (
  .A({ S25957[156] }),
  .B1({ S16696 }),
  .B2({ S16877 }),
  .ZN({ S16878 })
);
OAI21_X1 #() 
OAI21_X1_1197_ (
  .A({ S16376 }),
  .B1({ S16878 }),
  .B2({ S16876 }),
  .ZN({ S16879 })
);
AOI21_X1 #() 
AOI21_X1_1310_ (
  .A({ S15729 }),
  .B1({ S16879 }),
  .B2({ S16875 }),
  .ZN({ S16880 })
);
OAI21_X1 #() 
OAI21_X1_1198_ (
  .A({ S15640 }),
  .B1({ S16880 }),
  .B2({ S16871 }),
  .ZN({ S16881 })
);
NAND2_X1 #() 
NAND2_X1_2250_ (
  .A1({ S16508 }),
  .A2({ S16386 }),
  .ZN({ S16882 })
);
NAND2_X1 #() 
NAND2_X1_2251_ (
  .A1({ S16550 }),
  .A2({ S16882 }),
  .ZN({ S16883 })
);
NAND2_X1 #() 
NAND2_X1_2252_ (
  .A1({ S16883 }),
  .A2({ S25957[156] }),
  .ZN({ S16885 })
);
NAND2_X1 #() 
NAND2_X1_2253_ (
  .A1({ S16651 }),
  .A2({ S54 }),
  .ZN({ S16886 })
);
NAND2_X1 #() 
NAND2_X1_2254_ (
  .A1({ S16419 }),
  .A2({ S25957[155] }),
  .ZN({ S16887 })
);
NAND3_X1 #() 
NAND3_X1_2496_ (
  .A1({ S16887 }),
  .A2({ S16886 }),
  .A3({ S16485 }),
  .ZN({ S16888 })
);
OAI211_X1 #() 
OAI211_X1_813_ (
  .A({ S16885 }),
  .B({ S16376 }),
  .C1({ S25957[156] }),
  .C2({ S16888 }),
  .ZN({ S16889 })
);
INV_X1 #() 
INV_X1_720_ (
  .A({ S16445 }),
  .ZN({ S16890 })
);
OAI211_X1 #() 
OAI211_X1_814_ (
  .A({ S25957[156] }),
  .B({ S16483 }),
  .C1({ S16877 }),
  .C2({ S16890 }),
  .ZN({ S16891 })
);
OAI21_X1 #() 
OAI21_X1_1199_ (
  .A({ S25957[155] }),
  .B1({ S16755 }),
  .B2({ S16449 }),
  .ZN({ S16892 })
);
NAND3_X1 #() 
NAND3_X1_2497_ (
  .A1({ S16370 }),
  .A2({ S54 }),
  .A3({ S57 }),
  .ZN({ S16893 })
);
NAND3_X1 #() 
NAND3_X1_2498_ (
  .A1({ S16892 }),
  .A2({ S16359 }),
  .A3({ S16893 }),
  .ZN({ S16894 })
);
NAND3_X1 #() 
NAND3_X1_2499_ (
  .A1({ S16894 }),
  .A2({ S16891 }),
  .A3({ S25957[157] }),
  .ZN({ S16896 })
);
NAND3_X1 #() 
NAND3_X1_2500_ (
  .A1({ S16889 }),
  .A2({ S15729 }),
  .A3({ S16896 }),
  .ZN({ S16897 })
);
NAND2_X1 #() 
NAND2_X1_2255_ (
  .A1({ S16886 }),
  .A2({ S16485 }),
  .ZN({ S16898 })
);
AOI21_X1 #() 
AOI21_X1_1311_ (
  .A({ S25957[157] }),
  .B1({ S16553 }),
  .B2({ S16359 }),
  .ZN({ S16899 })
);
NOR4_X1 #() 
NOR4_X1_1_ (
  .A1({ S16554 }),
  .A2({ S16559 }),
  .A3({ S16489 }),
  .A4({ S25957[157] }),
  .ZN({ S16900 })
);
OAI22_X1 #() 
OAI22_X1_53_ (
  .A1({ S16900 }),
  .A2({ S16899 }),
  .B1({ S16697 }),
  .B2({ S16898 }),
  .ZN({ S16901 })
);
OAI21_X1 #() 
OAI21_X1_1200_ (
  .A({ S16589 }),
  .B1({ S16469 }),
  .B2({ S16467 }),
  .ZN({ S16902 })
);
NAND2_X1 #() 
NAND2_X1_2256_ (
  .A1({ S16864 }),
  .A2({ S16379 }),
  .ZN({ S16903 })
);
AOI21_X1 #() 
AOI21_X1_1312_ (
  .A({ S25957[156] }),
  .B1({ S16903 }),
  .B2({ S16398 }),
  .ZN({ S16904 })
);
AOI21_X1 #() 
AOI21_X1_1313_ (
  .A({ S16904 }),
  .B1({ S16902 }),
  .B2({ S25957[156] }),
  .ZN({ S16905 })
);
OAI211_X1 #() 
OAI211_X1_815_ (
  .A({ S16901 }),
  .B({ S25957[158] }),
  .C1({ S16376 }),
  .C2({ S16905 }),
  .ZN({ S16907 })
);
NAND3_X1 #() 
NAND3_X1_2501_ (
  .A1({ S16897 }),
  .A2({ S16907 }),
  .A3({ S25957[159] }),
  .ZN({ S16908 })
);
NAND2_X1 #() 
NAND2_X1_2257_ (
  .A1({ S16881 }),
  .A2({ S16908 }),
  .ZN({ S16909 })
);
XNOR2_X1 #() 
XNOR2_X1_126_ (
  .A({ S16909 }),
  .B({ S25957[230] }),
  .ZN({ S25957[102] })
);
OAI21_X1 #() 
OAI21_X1_1201_ (
  .A({ S16438 }),
  .B1({ S16338 }),
  .B2({ S16378 }),
  .ZN({ S16910 })
);
NAND2_X1 #() 
NAND2_X1_2258_ (
  .A1({ S16910 }),
  .A2({ S25957[156] }),
  .ZN({ S16911 })
);
NAND2_X1 #() 
NAND2_X1_2259_ (
  .A1({ S16747 }),
  .A2({ S16342 }),
  .ZN({ S16912 })
);
OAI221_X1 #() 
OAI221_X1_49_ (
  .A({ S16359 }),
  .B1({ S16605 }),
  .B2({ S16346 }),
  .C1({ S16912 }),
  .C2({ S25957[155] }),
  .ZN({ S16913 })
);
NAND2_X1 #() 
NAND2_X1_2260_ (
  .A1({ S16913 }),
  .A2({ S16911 }),
  .ZN({ S16914 })
);
NOR2_X1 #() 
NOR2_X1_537_ (
  .A1({ S16914 }),
  .A2({ S16376 }),
  .ZN({ S16915 })
);
NOR2_X1 #() 
NOR2_X1_538_ (
  .A1({ S16411 }),
  .A2({ S16511 }),
  .ZN({ S16917 })
);
NOR3_X1 #() 
NOR3_X1_69_ (
  .A1({ S16917 }),
  .A2({ S16607 }),
  .A3({ S16434 }),
  .ZN({ S16918 })
);
NOR2_X1 #() 
NOR2_X1_539_ (
  .A1({ S25957[157] }),
  .A2({ S16350 }),
  .ZN({ S16919 })
);
AOI22_X1 #() 
AOI22_X1_286_ (
  .A1({ S16919 }),
  .A2({ S16903 }),
  .B1({ S16376 }),
  .B2({ S16359 }),
  .ZN({ S16920 })
);
NOR2_X1 #() 
NOR2_X1_540_ (
  .A1({ S16918 }),
  .A2({ S16920 }),
  .ZN({ S16921 })
);
OAI21_X1 #() 
OAI21_X1_1202_ (
  .A({ S25957[158] }),
  .B1({ S16915 }),
  .B2({ S16921 }),
  .ZN({ S16922 })
);
OAI211_X1 #() 
OAI211_X1_816_ (
  .A({ S16634 }),
  .B({ S16570 }),
  .C1({ S16378 }),
  .C2({ S16755 }),
  .ZN({ S16923 })
);
NOR2_X1 #() 
NOR2_X1_541_ (
  .A1({ S25957[157] }),
  .A2({ S16359 }),
  .ZN({ S16924 })
);
NAND2_X1 #() 
NAND2_X1_2261_ (
  .A1({ S16923 }),
  .A2({ S16924 }),
  .ZN({ S16925 })
);
NAND3_X1 #() 
NAND3_X1_2502_ (
  .A1({ S16513 }),
  .A2({ S54 }),
  .A3({ S16468 }),
  .ZN({ S16926 })
);
NAND4_X1 #() 
NAND4_X1_310_ (
  .A1({ S16926 }),
  .A2({ S16554 }),
  .A3({ S16359 }),
  .A4({ S16376 }),
  .ZN({ S16928 })
);
NAND2_X1 #() 
NAND2_X1_2262_ (
  .A1({ S16353 }),
  .A2({ S16413 }),
  .ZN({ S16929 })
);
AOI21_X1 #() 
AOI21_X1_1314_ (
  .A({ S16359 }),
  .B1({ S16550 }),
  .B2({ S16929 }),
  .ZN({ S16930 })
);
NAND2_X1 #() 
NAND2_X1_2263_ (
  .A1({ S16344 }),
  .A2({ S16359 }),
  .ZN({ S16931 })
);
OAI21_X1 #() 
OAI21_X1_1203_ (
  .A({ S25957[157] }),
  .B1({ S16931 }),
  .B2({ S16864 }),
  .ZN({ S16932 })
);
OAI211_X1 #() 
OAI211_X1_817_ (
  .A({ S16925 }),
  .B({ S16928 }),
  .C1({ S16932 }),
  .C2({ S16930 }),
  .ZN({ S16933 })
);
NAND2_X1 #() 
NAND2_X1_2264_ (
  .A1({ S16933 }),
  .A2({ S15729 }),
  .ZN({ S16934 })
);
NAND3_X1 #() 
NAND3_X1_2503_ (
  .A1({ S16922 }),
  .A2({ S16934 }),
  .A3({ S25957[159] }),
  .ZN({ S16935 })
);
NOR2_X1 #() 
NOR2_X1_542_ (
  .A1({ S16626 }),
  .A2({ S16620 }),
  .ZN({ S16936 })
);
OAI21_X1 #() 
OAI21_X1_1204_ (
  .A({ S16359 }),
  .B1({ S16936 }),
  .B2({ S16775 }),
  .ZN({ S16937 })
);
NAND2_X1 #() 
NAND2_X1_2265_ (
  .A1({ S16769 }),
  .A2({ S16528 }),
  .ZN({ S16939 })
);
NAND2_X1 #() 
NAND2_X1_2266_ (
  .A1({ S16937 }),
  .A2({ S16939 }),
  .ZN({ S16940 })
);
INV_X1 #() 
INV_X1_721_ (
  .A({ S16940 }),
  .ZN({ S16941 })
);
INV_X1 #() 
INV_X1_722_ (
  .A({ S16605 }),
  .ZN({ S16942 })
);
NOR3_X1 #() 
NOR3_X1_70_ (
  .A1({ S16695 }),
  .A2({ S16942 }),
  .A3({ S16359 }),
  .ZN({ S16943 })
);
NAND2_X1 #() 
NAND2_X1_2267_ (
  .A1({ S16392 }),
  .A2({ S25957[155] }),
  .ZN({ S16944 })
);
AOI21_X1 #() 
AOI21_X1_1315_ (
  .A({ S25957[156] }),
  .B1({ S16674 }),
  .B2({ S16944 }),
  .ZN({ S16945 })
);
OAI21_X1 #() 
OAI21_X1_1205_ (
  .A({ S16376 }),
  .B1({ S16943 }),
  .B2({ S16945 }),
  .ZN({ S16946 })
);
OAI211_X1 #() 
OAI211_X1_818_ (
  .A({ S16946 }),
  .B({ S15729 }),
  .C1({ S16941 }),
  .C2({ S16376 }),
  .ZN({ S16947 })
);
NOR3_X1 #() 
NOR3_X1_71_ (
  .A1({ S16514 }),
  .A2({ S16714 }),
  .A3({ S16359 }),
  .ZN({ S16948 })
);
NAND2_X1 #() 
NAND2_X1_2268_ (
  .A1({ S16912 }),
  .A2({ S25957[155] }),
  .ZN({ S16950 })
);
NAND3_X1 #() 
NAND3_X1_2504_ (
  .A1({ S16950 }),
  .A2({ S25957[156] }),
  .A3({ S16504 }),
  .ZN({ S16951 })
);
OR3_X1 #() 
OR3_X1_11_ (
  .A1({ S16758 }),
  .A2({ S16535 }),
  .A3({ S25957[156] }),
  .ZN({ S16952 })
);
NAND2_X1 #() 
NAND2_X1_2269_ (
  .A1({ S16951 }),
  .A2({ S16952 }),
  .ZN({ S16953 })
);
NAND2_X1 #() 
NAND2_X1_2270_ (
  .A1({ S16553 }),
  .A2({ S16359 }),
  .ZN({ S16954 })
);
AOI21_X1 #() 
AOI21_X1_1316_ (
  .A({ S54 }),
  .B1({ S16383 }),
  .B2({ S16366 }),
  .ZN({ S16955 })
);
OAI21_X1 #() 
OAI21_X1_1206_ (
  .A({ S16376 }),
  .B1({ S16954 }),
  .B2({ S16955 }),
  .ZN({ S16956 })
);
OAI221_X1 #() 
OAI221_X1_50_ (
  .A({ S25957[158] }),
  .B1({ S16956 }),
  .B2({ S16948 }),
  .C1({ S16953 }),
  .C2({ S16376 }),
  .ZN({ S16957 })
);
NAND3_X1 #() 
NAND3_X1_2505_ (
  .A1({ S16957 }),
  .A2({ S16947 }),
  .A3({ S15640 }),
  .ZN({ S16958 })
);
NAND2_X1 #() 
NAND2_X1_2271_ (
  .A1({ S16935 }),
  .A2({ S16958 }),
  .ZN({ S16959 })
);
XNOR2_X1 #() 
XNOR2_X1_127_ (
  .A({ S16959 }),
  .B({ S25957[231] }),
  .ZN({ S25957[103] })
);
OAI21_X1 #() 
OAI21_X1_1207_ (
  .A({ S14141 }),
  .B1({ S15447 }),
  .B2({ S15443 }),
  .ZN({ S16961 })
);
NAND3_X1 #() 
NAND3_X1_2506_ (
  .A1({ S15449 }),
  .A2({ S15450 }),
  .A3({ S25957[257] }),
  .ZN({ S16962 })
);
NAND3_X1 #() 
NAND3_X1_2507_ (
  .A1({ S16961 }),
  .A2({ S25957[128] }),
  .A3({ S16962 }),
  .ZN({ S16963 })
);
INV_X1 #() 
INV_X1_723_ (
  .A({ S16963 }),
  .ZN({ S59 })
);
NAND2_X1 #() 
NAND2_X1_2272_ (
  .A1({ S15393 }),
  .A2({ S15356 }),
  .ZN({ S16964 })
);
NAND3_X1 #() 
NAND3_X1_2508_ (
  .A1({ S15448 }),
  .A2({ S16964 }),
  .A3({ S15451 }),
  .ZN({ S60 })
);
INV_X1 #() 
INV_X1_724_ (
  .A({ S25957[232] }),
  .ZN({ S16965 })
);
NAND2_X1 #() 
NAND2_X1_2273_ (
  .A1({ S14961 }),
  .A2({ S14962 }),
  .ZN({ S16966 })
);
NAND2_X1 #() 
NAND2_X1_2274_ (
  .A1({ S15134 }),
  .A2({ S15125 }),
  .ZN({ S16967 })
);
AOI21_X1 #() 
AOI21_X1_1317_ (
  .A({ S16964 }),
  .B1({ S15505 }),
  .B2({ S15510 }),
  .ZN({ S16969 })
);
NAND2_X1 #() 
NAND2_X1_2275_ (
  .A1({ S16963 }),
  .A2({ S25957[130] }),
  .ZN({ S16970 })
);
NAND2_X1 #() 
NAND2_X1_2276_ (
  .A1({ S16970 }),
  .A2({ S25957[131] }),
  .ZN({ S16971 })
);
AND3_X1 #() 
AND3_X1_100_ (
  .A1({ S25957[128] }),
  .A2({ S15505 }),
  .A3({ S15510 }),
  .ZN({ S16972 })
);
OAI21_X1 #() 
OAI21_X1_1208_ (
  .A({ S51 }),
  .B1({ S25957[129] }),
  .B2({ S16972 }),
  .ZN({ S16973 })
);
OAI21_X1 #() 
OAI21_X1_1209_ (
  .A({ S16973 }),
  .B1({ S16971 }),
  .B2({ S16969 }),
  .ZN({ S16974 })
);
AOI21_X1 #() 
AOI21_X1_1318_ (
  .A({ S25957[128] }),
  .B1({ S15505 }),
  .B2({ S15510 }),
  .ZN({ S16975 })
);
NAND2_X1 #() 
NAND2_X1_2277_ (
  .A1({ S25957[129] }),
  .A2({ S16975 }),
  .ZN({ S16976 })
);
NAND2_X1 #() 
NAND2_X1_2278_ (
  .A1({ S16961 }),
  .A2({ S16962 }),
  .ZN({ S16977 })
);
NAND2_X1 #() 
NAND2_X1_2279_ (
  .A1({ S16977 }),
  .A2({ S25957[130] }),
  .ZN({ S16978 })
);
NAND3_X1 #() 
NAND3_X1_2509_ (
  .A1({ S15302 }),
  .A2({ S15306 }),
  .A3({ S16964 }),
  .ZN({ S16980 })
);
NAND4_X1 #() 
NAND4_X1_311_ (
  .A1({ S16976 }),
  .A2({ S16978 }),
  .A3({ S25957[132] }),
  .A4({ S16980 }),
  .ZN({ S16981 })
);
OAI21_X1 #() 
OAI21_X1_1210_ (
  .A({ S16981 }),
  .B1({ S16974 }),
  .B2({ S25957[132] }),
  .ZN({ S16982 })
);
NAND2_X1 #() 
NAND2_X1_2280_ (
  .A1({ S16982 }),
  .A2({ S16967 }),
  .ZN({ S16983 })
);
NAND3_X1 #() 
NAND3_X1_2510_ (
  .A1({ S16961 }),
  .A2({ S16964 }),
  .A3({ S16962 }),
  .ZN({ S16984 })
);
NAND3_X1 #() 
NAND3_X1_2511_ (
  .A1({ S15505 }),
  .A2({ S15510 }),
  .A3({ S16964 }),
  .ZN({ S16985 })
);
NAND2_X1 #() 
NAND2_X1_2281_ (
  .A1({ S16984 }),
  .A2({ S16985 }),
  .ZN({ S16986 })
);
NAND3_X1 #() 
NAND3_X1_2512_ (
  .A1({ S15448 }),
  .A2({ S25957[128] }),
  .A3({ S15451 }),
  .ZN({ S16987 })
);
NAND3_X1 #() 
NAND3_X1_2513_ (
  .A1({ S16987 }),
  .A2({ S16984 }),
  .A3({ S25957[130] }),
  .ZN({ S16988 })
);
NAND2_X1 #() 
NAND2_X1_2282_ (
  .A1({ S15505 }),
  .A2({ S15510 }),
  .ZN({ S16989 })
);
NAND2_X1 #() 
NAND2_X1_2283_ (
  .A1({ S16977 }),
  .A2({ S16989 }),
  .ZN({ S16991 })
);
NAND2_X1 #() 
NAND2_X1_2284_ (
  .A1({ S16989 }),
  .A2({ S16964 }),
  .ZN({ S16992 })
);
NAND3_X1 #() 
NAND3_X1_2514_ (
  .A1({ S15302 }),
  .A2({ S15306 }),
  .A3({ S16992 }),
  .ZN({ S16993 })
);
INV_X1 #() 
INV_X1_725_ (
  .A({ S16993 }),
  .ZN({ S16994 })
);
NAND3_X1 #() 
NAND3_X1_2515_ (
  .A1({ S16988 }),
  .A2({ S16994 }),
  .A3({ S16991 }),
  .ZN({ S16995 })
);
OAI211_X1 #() 
OAI211_X1_819_ (
  .A({ S16995 }),
  .B({ S25957[132] }),
  .C1({ S25957[131] }),
  .C2({ S16986 }),
  .ZN({ S16996 })
);
AOI21_X1 #() 
AOI21_X1_1319_ (
  .A({ S16975 }),
  .B1({ S15306 }),
  .B2({ S15302 }),
  .ZN({ S16997 })
);
INV_X1 #() 
INV_X1_726_ (
  .A({ S16997 }),
  .ZN({ S16998 })
);
INV_X1 #() 
INV_X1_727_ (
  .A({ S16972 }),
  .ZN({ S16999 })
);
OAI21_X1 #() 
OAI21_X1_1211_ (
  .A({ S16999 }),
  .B1({ S16977 }),
  .B2({ S16992 }),
  .ZN({ S17000 })
);
INV_X1 #() 
INV_X1_728_ (
  .A({ S17000 }),
  .ZN({ S17002 })
);
NOR2_X1 #() 
NOR2_X1_543_ (
  .A1({ S25957[129] }),
  .A2({ S16989 }),
  .ZN({ S17003 })
);
NOR2_X1 #() 
NOR2_X1_544_ (
  .A1({ S17003 }),
  .A2({ S51 }),
  .ZN({ S17004 })
);
AOI21_X1 #() 
AOI21_X1_1320_ (
  .A({ S25957[132] }),
  .B1({ S17004 }),
  .B2({ S17002 }),
  .ZN({ S17005 })
);
NAND2_X1 #() 
NAND2_X1_2285_ (
  .A1({ S17005 }),
  .A2({ S16998 }),
  .ZN({ S17006 })
);
NAND3_X1 #() 
NAND3_X1_2516_ (
  .A1({ S17006 }),
  .A2({ S16996 }),
  .A3({ S25957[133] }),
  .ZN({ S17007 })
);
AND2_X1 #() 
AND2_X1_140_ (
  .A1({ S16983 }),
  .A2({ S17007 }),
  .ZN({ S17008 })
);
NAND2_X1 #() 
NAND2_X1_2286_ (
  .A1({ S16963 }),
  .A2({ S60 }),
  .ZN({ S17009 })
);
NAND2_X1 #() 
NAND2_X1_2287_ (
  .A1({ S17009 }),
  .A2({ S16992 }),
  .ZN({ S17010 })
);
NAND2_X1 #() 
NAND2_X1_2288_ (
  .A1({ S17010 }),
  .A2({ S51 }),
  .ZN({ S17011 })
);
NAND2_X1 #() 
NAND2_X1_2289_ (
  .A1({ S16977 }),
  .A2({ S16975 }),
  .ZN({ S17013 })
);
NAND3_X1 #() 
NAND3_X1_2517_ (
  .A1({ S15448 }),
  .A2({ S16972 }),
  .A3({ S15451 }),
  .ZN({ S17014 })
);
NAND3_X1 #() 
NAND3_X1_2518_ (
  .A1({ S17014 }),
  .A2({ S15302 }),
  .A3({ S15306 }),
  .ZN({ S17015 })
);
INV_X1 #() 
INV_X1_729_ (
  .A({ S17015 }),
  .ZN({ S17016 })
);
NAND2_X1 #() 
NAND2_X1_2290_ (
  .A1({ S17016 }),
  .A2({ S17013 }),
  .ZN({ S17017 })
);
NAND2_X1 #() 
NAND2_X1_2291_ (
  .A1({ S17011 }),
  .A2({ S17017 }),
  .ZN({ S17018 })
);
NAND2_X1 #() 
NAND2_X1_2292_ (
  .A1({ S16989 }),
  .A2({ S25957[128] }),
  .ZN({ S17019 })
);
NAND2_X1 #() 
NAND2_X1_2293_ (
  .A1({ S16984 }),
  .A2({ S17019 }),
  .ZN({ S17020 })
);
NOR2_X1 #() 
NOR2_X1_545_ (
  .A1({ S17020 }),
  .A2({ S25957[131] }),
  .ZN({ S17021 })
);
NAND3_X1 #() 
NAND3_X1_2519_ (
  .A1({ S25957[131] }),
  .A2({ S60 }),
  .A3({ S16999 }),
  .ZN({ S17022 })
);
INV_X1 #() 
INV_X1_730_ (
  .A({ S17022 }),
  .ZN({ S17024 })
);
OAI21_X1 #() 
OAI21_X1_1212_ (
  .A({ S25957[132] }),
  .B1({ S17024 }),
  .B2({ S17021 }),
  .ZN({ S17025 })
);
OAI21_X1 #() 
OAI21_X1_1213_ (
  .A({ S17025 }),
  .B1({ S17018 }),
  .B2({ S25957[132] }),
  .ZN({ S17026 })
);
NAND2_X1 #() 
NAND2_X1_2294_ (
  .A1({ S17026 }),
  .A2({ S25957[133] }),
  .ZN({ S17027 })
);
NAND2_X1 #() 
NAND2_X1_2295_ (
  .A1({ S15215 }),
  .A2({ S15218 }),
  .ZN({ S17028 })
);
NAND4_X1 #() 
NAND4_X1_312_ (
  .A1({ S16961 }),
  .A2({ S25957[128] }),
  .A3({ S16962 }),
  .A4({ S25957[130] }),
  .ZN({ S17029 })
);
NAND3_X1 #() 
NAND3_X1_2520_ (
  .A1({ S15448 }),
  .A2({ S15451 }),
  .A3({ S16969 }),
  .ZN({ S17030 })
);
AND4_X1 #() 
AND4_X1_7_ (
  .A1({ S51 }),
  .A2({ S17029 }),
  .A3({ S17030 }),
  .A4({ S60 }),
  .ZN({ S17031 })
);
AOI21_X1 #() 
AOI21_X1_1321_ (
  .A({ S25957[130] }),
  .B1({ S16963 }),
  .B2({ S60 }),
  .ZN({ S17032 })
);
AOI21_X1 #() 
AOI21_X1_1322_ (
  .A({ S17031 }),
  .B1({ S25957[131] }),
  .B2({ S17032 }),
  .ZN({ S17033 })
);
NAND2_X1 #() 
NAND2_X1_2296_ (
  .A1({ S16988 }),
  .A2({ S17013 }),
  .ZN({ S17035 })
);
INV_X1 #() 
INV_X1_731_ (
  .A({ S16985 }),
  .ZN({ S17036 })
);
NAND3_X1 #() 
NAND3_X1_2521_ (
  .A1({ S17036 }),
  .A2({ S15448 }),
  .A3({ S15451 }),
  .ZN({ S17037 })
);
NAND3_X1 #() 
NAND3_X1_2522_ (
  .A1({ S17037 }),
  .A2({ S51 }),
  .A3({ S17030 }),
  .ZN({ S17038 })
);
OAI21_X1 #() 
OAI21_X1_1214_ (
  .A({ S17038 }),
  .B1({ S17035 }),
  .B2({ S51 }),
  .ZN({ S17039 })
);
NAND2_X1 #() 
NAND2_X1_2297_ (
  .A1({ S17039 }),
  .A2({ S17028 }),
  .ZN({ S17040 })
);
OAI211_X1 #() 
OAI211_X1_820_ (
  .A({ S17040 }),
  .B({ S16967 }),
  .C1({ S17028 }),
  .C2({ S17033 }),
  .ZN({ S17041 })
);
NAND3_X1 #() 
NAND3_X1_2523_ (
  .A1({ S17027 }),
  .A2({ S17041 }),
  .A3({ S15041 }),
  .ZN({ S17042 })
);
OAI211_X1 #() 
OAI211_X1_821_ (
  .A({ S17042 }),
  .B({ S16966 }),
  .C1({ S15041 }),
  .C2({ S17008 }),
  .ZN({ S17043 })
);
AOI21_X1 #() 
AOI21_X1_1323_ (
  .A({ S16989 }),
  .B1({ S15448 }),
  .B2({ S15451 }),
  .ZN({ S17044 })
);
NAND2_X1 #() 
NAND2_X1_2298_ (
  .A1({ S17044 }),
  .A2({ S51 }),
  .ZN({ S17046 })
);
NOR2_X1 #() 
NOR2_X1_546_ (
  .A1({ S25957[129] }),
  .A2({ S16992 }),
  .ZN({ S17047 })
);
OAI21_X1 #() 
OAI21_X1_1215_ (
  .A({ S51 }),
  .B1({ S17047 }),
  .B2({ S16972 }),
  .ZN({ S17048 })
);
NAND2_X1 #() 
NAND2_X1_2299_ (
  .A1({ S17048 }),
  .A2({ S17046 }),
  .ZN({ S17049 })
);
NAND2_X1 #() 
NAND2_X1_2300_ (
  .A1({ S16984 }),
  .A2({ S25957[130] }),
  .ZN({ S17050 })
);
NOR2_X1 #() 
NOR2_X1_547_ (
  .A1({ S17050 }),
  .A2({ S51 }),
  .ZN({ S17051 })
);
OAI21_X1 #() 
OAI21_X1_1216_ (
  .A({ S25957[132] }),
  .B1({ S17049 }),
  .B2({ S17051 }),
  .ZN({ S17052 })
);
NAND3_X1 #() 
NAND3_X1_2524_ (
  .A1({ S16963 }),
  .A2({ S60 }),
  .A3({ S16989 }),
  .ZN({ S17053 })
);
NOR2_X1 #() 
NOR2_X1_548_ (
  .A1({ S25957[131] }),
  .A2({ S17044 }),
  .ZN({ S17054 })
);
NAND2_X1 #() 
NAND2_X1_2301_ (
  .A1({ S17054 }),
  .A2({ S17053 }),
  .ZN({ S17055 })
);
NAND3_X1 #() 
NAND3_X1_2525_ (
  .A1({ S25957[131] }),
  .A2({ S16985 }),
  .A3({ S17030 }),
  .ZN({ S17057 })
);
NAND3_X1 #() 
NAND3_X1_2526_ (
  .A1({ S17055 }),
  .A2({ S17028 }),
  .A3({ S17057 }),
  .ZN({ S17058 })
);
AOI21_X1 #() 
AOI21_X1_1324_ (
  .A({ S16967 }),
  .B1({ S17052 }),
  .B2({ S17058 }),
  .ZN({ S17059 })
);
NOR2_X1 #() 
NOR2_X1_549_ (
  .A1({ S16988 }),
  .A2({ S51 }),
  .ZN({ S17060 })
);
AOI21_X1 #() 
AOI21_X1_1325_ (
  .A({ S17044 }),
  .B1({ S16976 }),
  .B2({ S16999 }),
  .ZN({ S17061 })
);
OAI21_X1 #() 
OAI21_X1_1217_ (
  .A({ S25957[132] }),
  .B1({ S17061 }),
  .B2({ S25957[131] }),
  .ZN({ S17062 })
);
NAND2_X1 #() 
NAND2_X1_2302_ (
  .A1({ S16976 }),
  .A2({ S51 }),
  .ZN({ S17063 })
);
AOI21_X1 #() 
AOI21_X1_1326_ (
  .A({ S51 }),
  .B1({ S17029 }),
  .B2({ S16992 }),
  .ZN({ S17064 })
);
NOR2_X1 #() 
NOR2_X1_550_ (
  .A1({ S17064 }),
  .A2({ S25957[132] }),
  .ZN({ S17065 })
);
NAND2_X1 #() 
NAND2_X1_2303_ (
  .A1({ S17065 }),
  .A2({ S17063 }),
  .ZN({ S17066 })
);
OAI21_X1 #() 
OAI21_X1_1218_ (
  .A({ S17066 }),
  .B1({ S17062 }),
  .B2({ S17060 }),
  .ZN({ S17068 })
);
OAI21_X1 #() 
OAI21_X1_1219_ (
  .A({ S25957[134] }),
  .B1({ S17068 }),
  .B2({ S25957[133] }),
  .ZN({ S17069 })
);
AOI21_X1 #() 
AOI21_X1_1327_ (
  .A({ S16985 }),
  .B1({ S16961 }),
  .B2({ S16962 }),
  .ZN({ S17070 })
);
AOI21_X1 #() 
AOI21_X1_1328_ (
  .A({ S17036 }),
  .B1({ S15306 }),
  .B2({ S15302 }),
  .ZN({ S17071 })
);
NOR2_X1 #() 
NOR2_X1_551_ (
  .A1({ S25957[129] }),
  .A2({ S25957[130] }),
  .ZN({ S17072 })
);
AOI21_X1 #() 
AOI21_X1_1329_ (
  .A({ S16964 }),
  .B1({ S15306 }),
  .B2({ S15302 }),
  .ZN({ S17073 })
);
AOI21_X1 #() 
AOI21_X1_1330_ (
  .A({ S17028 }),
  .B1({ S17072 }),
  .B2({ S17073 }),
  .ZN({ S17074 })
);
OAI21_X1 #() 
OAI21_X1_1220_ (
  .A({ S17074 }),
  .B1({ S17070 }),
  .B2({ S17071 }),
  .ZN({ S17075 })
);
NAND3_X1 #() 
NAND3_X1_2527_ (
  .A1({ S17036 }),
  .A2({ S16961 }),
  .A3({ S16962 }),
  .ZN({ S17076 })
);
INV_X1 #() 
INV_X1_732_ (
  .A({ S17076 }),
  .ZN({ S17077 })
);
NAND3_X1 #() 
NAND3_X1_2528_ (
  .A1({ S16961 }),
  .A2({ S16962 }),
  .A3({ S16989 }),
  .ZN({ S17079 })
);
NAND2_X1 #() 
NAND2_X1_2304_ (
  .A1({ S17079 }),
  .A2({ S16992 }),
  .ZN({ S17080 })
);
NOR2_X1 #() 
NOR2_X1_552_ (
  .A1({ S17080 }),
  .A2({ S17077 }),
  .ZN({ S17081 })
);
NOR2_X1 #() 
NOR2_X1_553_ (
  .A1({ S17081 }),
  .A2({ S51 }),
  .ZN({ S17082 })
);
OAI21_X1 #() 
OAI21_X1_1221_ (
  .A({ S17028 }),
  .B1({ S25957[131] }),
  .B2({ S17070 }),
  .ZN({ S17083 })
);
OAI211_X1 #() 
OAI211_X1_822_ (
  .A({ S17075 }),
  .B({ S25957[133] }),
  .C1({ S17082 }),
  .C2({ S17083 }),
  .ZN({ S17084 })
);
NAND2_X1 #() 
NAND2_X1_2305_ (
  .A1({ S17020 }),
  .A2({ S16992 }),
  .ZN({ S17085 })
);
NOR2_X1 #() 
NOR2_X1_554_ (
  .A1({ S17085 }),
  .A2({ S25957[131] }),
  .ZN({ S17086 })
);
OAI21_X1 #() 
OAI21_X1_1222_ (
  .A({ S17028 }),
  .B1({ S16980 }),
  .B2({ S17044 }),
  .ZN({ S17087 })
);
NAND2_X1 #() 
NAND2_X1_2306_ (
  .A1({ S25957[131] }),
  .A2({ S17044 }),
  .ZN({ S17088 })
);
OAI21_X1 #() 
OAI21_X1_1223_ (
  .A({ S17088 }),
  .B1({ S17053 }),
  .B2({ S25957[131] }),
  .ZN({ S17090 })
);
AOI21_X1 #() 
AOI21_X1_1331_ (
  .A({ S25957[133] }),
  .B1({ S17090 }),
  .B2({ S25957[132] }),
  .ZN({ S17091 })
);
OAI21_X1 #() 
OAI21_X1_1224_ (
  .A({ S17091 }),
  .B1({ S17086 }),
  .B2({ S17087 }),
  .ZN({ S17092 })
);
NAND2_X1 #() 
NAND2_X1_2307_ (
  .A1({ S17092 }),
  .A2({ S17084 }),
  .ZN({ S17093 })
);
OAI221_X1 #() 
OAI221_X1_51_ (
  .A({ S25957[135] }),
  .B1({ S17093 }),
  .B2({ S25957[134] }),
  .C1({ S17069 }),
  .C2({ S17059 }),
  .ZN({ S17094 })
);
NAND3_X1 #() 
NAND3_X1_2529_ (
  .A1({ S17043 }),
  .A2({ S17094 }),
  .A3({ S16965 }),
  .ZN({ S17095 })
);
NOR2_X1 #() 
NOR2_X1_555_ (
  .A1({ S17068 }),
  .A2({ S25957[133] }),
  .ZN({ S17096 })
);
OAI21_X1 #() 
OAI21_X1_1225_ (
  .A({ S25957[134] }),
  .B1({ S17096 }),
  .B2({ S17059 }),
  .ZN({ S17097 })
);
NAND2_X1 #() 
NAND2_X1_2308_ (
  .A1({ S17093 }),
  .A2({ S15041 }),
  .ZN({ S17098 })
);
NAND3_X1 #() 
NAND3_X1_2530_ (
  .A1({ S17097 }),
  .A2({ S25957[135] }),
  .A3({ S17098 }),
  .ZN({ S17099 })
);
NAND3_X1 #() 
NAND3_X1_2531_ (
  .A1({ S16983 }),
  .A2({ S17007 }),
  .A3({ S25957[134] }),
  .ZN({ S17101 })
);
NAND2_X1 #() 
NAND2_X1_2309_ (
  .A1({ S17033 }),
  .A2({ S25957[132] }),
  .ZN({ S17102 })
);
OAI211_X1 #() 
OAI211_X1_823_ (
  .A({ S17102 }),
  .B({ S16967 }),
  .C1({ S25957[132] }),
  .C2({ S17039 }),
  .ZN({ S17103 })
);
OAI211_X1 #() 
OAI211_X1_824_ (
  .A({ S25957[133] }),
  .B({ S17025 }),
  .C1({ S17018 }),
  .C2({ S25957[132] }),
  .ZN({ S17104 })
);
NAND3_X1 #() 
NAND3_X1_2532_ (
  .A1({ S17103 }),
  .A2({ S17104 }),
  .A3({ S15041 }),
  .ZN({ S17105 })
);
NAND3_X1 #() 
NAND3_X1_2533_ (
  .A1({ S17105 }),
  .A2({ S16966 }),
  .A3({ S17101 }),
  .ZN({ S17106 })
);
NAND3_X1 #() 
NAND3_X1_2534_ (
  .A1({ S17099 }),
  .A2({ S17106 }),
  .A3({ S25957[232] }),
  .ZN({ S17107 })
);
NAND2_X1 #() 
NAND2_X1_2310_ (
  .A1({ S17095 }),
  .A2({ S17107 }),
  .ZN({ S25957[104] })
);
INV_X1 #() 
INV_X1_733_ (
  .A({ S25957[233] }),
  .ZN({ S17108 })
);
NAND2_X1 #() 
NAND2_X1_2311_ (
  .A1({ S17076 }),
  .A2({ S51 }),
  .ZN({ S17109 })
);
NAND3_X1 #() 
NAND3_X1_2535_ (
  .A1({ S16995 }),
  .A2({ S17028 }),
  .A3({ S17109 }),
  .ZN({ S17111 })
);
NAND2_X1 #() 
NAND2_X1_2312_ (
  .A1({ S16978 }),
  .A2({ S16985 }),
  .ZN({ S17112 })
);
NAND2_X1 #() 
NAND2_X1_2313_ (
  .A1({ S25957[129] }),
  .A2({ S16992 }),
  .ZN({ S17113 })
);
NAND2_X1 #() 
NAND2_X1_2314_ (
  .A1({ S17113 }),
  .A2({ S25957[131] }),
  .ZN({ S17114 })
);
OAI211_X1 #() 
OAI211_X1_825_ (
  .A({ S25957[132] }),
  .B({ S17114 }),
  .C1({ S17112 }),
  .C2({ S25957[131] }),
  .ZN({ S17115 })
);
NAND3_X1 #() 
NAND3_X1_2536_ (
  .A1({ S17111 }),
  .A2({ S25957[133] }),
  .A3({ S17115 }),
  .ZN({ S17116 })
);
NAND3_X1 #() 
NAND3_X1_2537_ (
  .A1({ S16963 }),
  .A2({ S60 }),
  .A3({ S25957[130] }),
  .ZN({ S17117 })
);
NAND2_X1 #() 
NAND2_X1_2315_ (
  .A1({ S16991 }),
  .A2({ S25957[131] }),
  .ZN({ S17118 })
);
NOR2_X1 #() 
NOR2_X1_556_ (
  .A1({ S17118 }),
  .A2({ S16969 }),
  .ZN({ S17119 })
);
NAND2_X1 #() 
NAND2_X1_2316_ (
  .A1({ S17119 }),
  .A2({ S17117 }),
  .ZN({ S17120 })
);
INV_X1 #() 
INV_X1_734_ (
  .A({ S17046 }),
  .ZN({ S17122 })
);
NOR3_X1 #() 
NOR3_X1_72_ (
  .A1({ S17122 }),
  .A2({ S17073 }),
  .A3({ S17028 }),
  .ZN({ S17123 })
);
NAND2_X1 #() 
NAND2_X1_2317_ (
  .A1({ S17072 }),
  .A2({ S17073 }),
  .ZN({ S17124 })
);
NAND2_X1 #() 
NAND2_X1_2318_ (
  .A1({ S16986 }),
  .A2({ S51 }),
  .ZN({ S17125 })
);
NAND2_X1 #() 
NAND2_X1_2319_ (
  .A1({ S25957[131] }),
  .A2({ S16963 }),
  .ZN({ S17126 })
);
OAI211_X1 #() 
OAI211_X1_826_ (
  .A({ S17125 }),
  .B({ S17124 }),
  .C1({ S17036 }),
  .C2({ S17126 }),
  .ZN({ S17127 })
);
AOI22_X1 #() 
AOI22_X1_287_ (
  .A1({ S17120 }),
  .A2({ S17123 }),
  .B1({ S17127 }),
  .B2({ S17028 }),
  .ZN({ S17128 })
);
OAI211_X1 #() 
OAI211_X1_827_ (
  .A({ S25957[134] }),
  .B({ S17116 }),
  .C1({ S17128 }),
  .C2({ S25957[133] }),
  .ZN({ S17129 })
);
NAND3_X1 #() 
NAND3_X1_2538_ (
  .A1({ S17050 }),
  .A2({ S51 }),
  .A3({ S17019 }),
  .ZN({ S17130 })
);
INV_X1 #() 
INV_X1_735_ (
  .A({ S17130 }),
  .ZN({ S17131 })
);
AOI21_X1 #() 
AOI21_X1_1332_ (
  .A({ S51 }),
  .B1({ S17117 }),
  .B2({ S17019 }),
  .ZN({ S17133 })
);
OAI21_X1 #() 
OAI21_X1_1226_ (
  .A({ S25957[132] }),
  .B1({ S17131 }),
  .B2({ S17133 }),
  .ZN({ S17134 })
);
INV_X1 #() 
INV_X1_736_ (
  .A({ S16987 }),
  .ZN({ S17135 })
);
NAND2_X1 #() 
NAND2_X1_2320_ (
  .A1({ S51 }),
  .A2({ S17079 }),
  .ZN({ S17136 })
);
OAI221_X1 #() 
OAI221_X1_52_ (
  .A({ S17028 }),
  .B1({ S17136 }),
  .B2({ S17135 }),
  .C1({ S17118 }),
  .C2({ S16969 }),
  .ZN({ S17137 })
);
NAND3_X1 #() 
NAND3_X1_2539_ (
  .A1({ S17134 }),
  .A2({ S17137 }),
  .A3({ S25957[133] }),
  .ZN({ S17138 })
);
NAND2_X1 #() 
NAND2_X1_2321_ (
  .A1({ S17009 }),
  .A2({ S16989 }),
  .ZN({ S17139 })
);
AOI21_X1 #() 
AOI21_X1_1333_ (
  .A({ S51 }),
  .B1({ S17139 }),
  .B2({ S16970 }),
  .ZN({ S17140 })
);
NAND3_X1 #() 
NAND3_X1_2540_ (
  .A1({ S17050 }),
  .A2({ S51 }),
  .A3({ S16976 }),
  .ZN({ S17141 })
);
NAND2_X1 #() 
NAND2_X1_2322_ (
  .A1({ S17141 }),
  .A2({ S17028 }),
  .ZN({ S17142 })
);
NAND3_X1 #() 
NAND3_X1_2541_ (
  .A1({ S25957[131] }),
  .A2({ S25957[129] }),
  .A3({ S16989 }),
  .ZN({ S17144 })
);
OAI21_X1 #() 
OAI21_X1_1227_ (
  .A({ S17144 }),
  .B1({ S17063 }),
  .B2({ S17003 }),
  .ZN({ S17145 })
);
OAI221_X1 #() 
OAI221_X1_53_ (
  .A({ S16967 }),
  .B1({ S17145 }),
  .B2({ S17028 }),
  .C1({ S17140 }),
  .C2({ S17142 }),
  .ZN({ S17146 })
);
NAND3_X1 #() 
NAND3_X1_2542_ (
  .A1({ S17146 }),
  .A2({ S17138 }),
  .A3({ S15041 }),
  .ZN({ S17147 })
);
NAND3_X1 #() 
NAND3_X1_2543_ (
  .A1({ S17129 }),
  .A2({ S17147 }),
  .A3({ S25957[135] }),
  .ZN({ S17148 })
);
OAI21_X1 #() 
OAI21_X1_1228_ (
  .A({ S25957[131] }),
  .B1({ S16977 }),
  .B2({ S16972 }),
  .ZN({ S17149 })
);
NAND3_X1 #() 
NAND3_X1_2544_ (
  .A1({ S25957[133] }),
  .A2({ S17048 }),
  .A3({ S17149 }),
  .ZN({ S17150 })
);
NAND2_X1 #() 
NAND2_X1_2323_ (
  .A1({ S51 }),
  .A2({ S17019 }),
  .ZN({ S17151 })
);
NOR2_X1 #() 
NOR2_X1_557_ (
  .A1({ S17112 }),
  .A2({ S17151 }),
  .ZN({ S17152 })
);
OAI21_X1 #() 
OAI21_X1_1229_ (
  .A({ S16967 }),
  .B1({ S16988 }),
  .B2({ S51 }),
  .ZN({ S17153 })
);
OAI211_X1 #() 
OAI211_X1_828_ (
  .A({ S17150 }),
  .B({ S17028 }),
  .C1({ S17152 }),
  .C2({ S17153 }),
  .ZN({ S17155 })
);
OAI21_X1 #() 
OAI21_X1_1230_ (
  .A({ S60 }),
  .B1({ S16963 }),
  .B2({ S25957[130] }),
  .ZN({ S17156 })
);
NOR2_X1 #() 
NOR2_X1_558_ (
  .A1({ S17156 }),
  .A2({ S51 }),
  .ZN({ S17157 })
);
NAND2_X1 #() 
NAND2_X1_2324_ (
  .A1({ S60 }),
  .A2({ S25957[130] }),
  .ZN({ S17158 })
);
AND2_X1 #() 
AND2_X1_141_ (
  .A1({ S17158 }),
  .A2({ S16997 }),
  .ZN({ S17159 })
);
OAI21_X1 #() 
OAI21_X1_1231_ (
  .A({ S25957[133] }),
  .B1({ S17157 }),
  .B2({ S17159 }),
  .ZN({ S17160 })
);
NAND2_X1 #() 
NAND2_X1_2325_ (
  .A1({ S17079 }),
  .A2({ S16985 }),
  .ZN({ S17161 })
);
OAI21_X1 #() 
OAI21_X1_1232_ (
  .A({ S51 }),
  .B1({ S17161 }),
  .B2({ S17135 }),
  .ZN({ S17162 })
);
NAND3_X1 #() 
NAND3_X1_2545_ (
  .A1({ S16995 }),
  .A2({ S17162 }),
  .A3({ S16967 }),
  .ZN({ S17163 })
);
NAND3_X1 #() 
NAND3_X1_2546_ (
  .A1({ S17160 }),
  .A2({ S25957[132] }),
  .A3({ S17163 }),
  .ZN({ S17164 })
);
AOI21_X1 #() 
AOI21_X1_1334_ (
  .A({ S15041 }),
  .B1({ S17164 }),
  .B2({ S17155 }),
  .ZN({ S17166 })
);
NAND3_X1 #() 
NAND3_X1_2547_ (
  .A1({ S17029 }),
  .A2({ S51 }),
  .A3({ S17030 }),
  .ZN({ S17167 })
);
INV_X1 #() 
INV_X1_737_ (
  .A({ S17118 }),
  .ZN({ S17168 })
);
NAND2_X1 #() 
NAND2_X1_2326_ (
  .A1({ S17168 }),
  .A2({ S16967 }),
  .ZN({ S17169 })
);
AOI21_X1 #() 
AOI21_X1_1335_ (
  .A({ S25957[132] }),
  .B1({ S17169 }),
  .B2({ S17167 }),
  .ZN({ S17170 })
);
AOI22_X1 #() 
AOI22_X1_288_ (
  .A1({ S25957[129] }),
  .A2({ S16989 }),
  .B1({ S15306 }),
  .B2({ S15302 }),
  .ZN({ S17171 })
);
NAND2_X1 #() 
NAND2_X1_2327_ (
  .A1({ S17171 }),
  .A2({ S16964 }),
  .ZN({ S17172 })
);
NAND3_X1 #() 
NAND3_X1_2548_ (
  .A1({ S25957[129] }),
  .A2({ S16985 }),
  .A3({ S17019 }),
  .ZN({ S17173 })
);
OAI211_X1 #() 
OAI211_X1_829_ (
  .A({ S25957[133] }),
  .B({ S17172 }),
  .C1({ S51 }),
  .C2({ S17173 }),
  .ZN({ S17174 })
);
INV_X1 #() 
INV_X1_738_ (
  .A({ S17071 }),
  .ZN({ S17175 })
);
OAI211_X1 #() 
OAI211_X1_830_ (
  .A({ S16967 }),
  .B({ S17149 }),
  .C1({ S17072 }),
  .C2({ S17175 }),
  .ZN({ S17177 })
);
AOI21_X1 #() 
AOI21_X1_1336_ (
  .A({ S17028 }),
  .B1({ S17174 }),
  .B2({ S17177 }),
  .ZN({ S17178 })
);
NOR3_X1 #() 
NOR3_X1_73_ (
  .A1({ S17178 }),
  .A2({ S17170 }),
  .A3({ S25957[134] }),
  .ZN({ S17179 })
);
OAI21_X1 #() 
OAI21_X1_1233_ (
  .A({ S16966 }),
  .B1({ S17179 }),
  .B2({ S17166 }),
  .ZN({ S17180 })
);
NAND3_X1 #() 
NAND3_X1_2549_ (
  .A1({ S17180 }),
  .A2({ S17148 }),
  .A3({ S17108 }),
  .ZN({ S17181 })
);
NAND2_X1 #() 
NAND2_X1_2328_ (
  .A1({ S17180 }),
  .A2({ S17148 }),
  .ZN({ S17182 })
);
NAND2_X1 #() 
NAND2_X1_2329_ (
  .A1({ S17182 }),
  .A2({ S25957[233] }),
  .ZN({ S17183 })
);
NAND2_X1 #() 
NAND2_X1_2330_ (
  .A1({ S17183 }),
  .A2({ S17181 }),
  .ZN({ S25957[105] })
);
INV_X1 #() 
INV_X1_739_ (
  .A({ S16984 }),
  .ZN({ S17184 })
);
NAND2_X1 #() 
NAND2_X1_2331_ (
  .A1({ S17158 }),
  .A2({ S51 }),
  .ZN({ S17185 })
);
OAI211_X1 #() 
OAI211_X1_831_ (
  .A({ S17185 }),
  .B({ S17028 }),
  .C1({ S17184 }),
  .C2({ S17015 }),
  .ZN({ S17187 })
);
AOI22_X1 #() 
AOI22_X1_289_ (
  .A1({ S17029 }),
  .A2({ S17030 }),
  .B1({ S15306 }),
  .B2({ S15302 }),
  .ZN({ S17188 })
);
INV_X1 #() 
INV_X1_740_ (
  .A({ S17188 }),
  .ZN({ S17189 })
);
NAND2_X1 #() 
NAND2_X1_2332_ (
  .A1({ S17168 }),
  .A2({ S25957[128] }),
  .ZN({ S17190 })
);
NAND3_X1 #() 
NAND3_X1_2550_ (
  .A1({ S17190 }),
  .A2({ S25957[132] }),
  .A3({ S17189 }),
  .ZN({ S17191 })
);
NAND3_X1 #() 
NAND3_X1_2551_ (
  .A1({ S17191 }),
  .A2({ S25957[133] }),
  .A3({ S17187 }),
  .ZN({ S17192 })
);
NAND2_X1 #() 
NAND2_X1_2333_ (
  .A1({ S25957[129] }),
  .A2({ S17019 }),
  .ZN({ S17193 })
);
NOR2_X1 #() 
NOR2_X1_559_ (
  .A1({ S17193 }),
  .A2({ S51 }),
  .ZN({ S17194 })
);
NOR2_X1 #() 
NOR2_X1_560_ (
  .A1({ S17194 }),
  .A2({ S17028 }),
  .ZN({ S17195 })
);
INV_X1 #() 
INV_X1_741_ (
  .A({ S16976 }),
  .ZN({ S17196 })
);
NAND2_X1 #() 
NAND2_X1_2334_ (
  .A1({ S17196 }),
  .A2({ S51 }),
  .ZN({ S17198 })
);
NAND3_X1 #() 
NAND3_X1_2552_ (
  .A1({ S16961 }),
  .A2({ S16962 }),
  .A3({ S25957[130] }),
  .ZN({ S17199 })
);
NOR2_X1 #() 
NOR2_X1_561_ (
  .A1({ S51 }),
  .A2({ S17199 }),
  .ZN({ S17200 })
);
NOR2_X1 #() 
NOR2_X1_562_ (
  .A1({ S17200 }),
  .A2({ S25957[132] }),
  .ZN({ S17201 })
);
AOI22_X1 #() 
AOI22_X1_290_ (
  .A1({ S17195 }),
  .A2({ S17136 }),
  .B1({ S17201 }),
  .B2({ S17198 }),
  .ZN({ S17202 })
);
NAND2_X1 #() 
NAND2_X1_2335_ (
  .A1({ S17202 }),
  .A2({ S16967 }),
  .ZN({ S17203 })
);
AOI21_X1 #() 
AOI21_X1_1337_ (
  .A({ S25957[134] }),
  .B1({ S17192 }),
  .B2({ S17203 }),
  .ZN({ S17204 })
);
NAND3_X1 #() 
NAND3_X1_2553_ (
  .A1({ S17019 }),
  .A2({ S15448 }),
  .A3({ S15451 }),
  .ZN({ S17205 })
);
INV_X1 #() 
INV_X1_742_ (
  .A({ S17205 }),
  .ZN({ S17206 })
);
OAI221_X1 #() 
OAI221_X1_54_ (
  .A({ S25957[132] }),
  .B1({ S17206 }),
  .B2({ S25957[131] }),
  .C1({ S17032 }),
  .C2({ S17015 }),
  .ZN({ S17207 })
);
NOR2_X1 #() 
NOR2_X1_563_ (
  .A1({ S51 }),
  .A2({ S16989 }),
  .ZN({ S17209 })
);
NAND2_X1 #() 
NAND2_X1_2336_ (
  .A1({ S17135 }),
  .A2({ S25957[131] }),
  .ZN({ S17210 })
);
OAI211_X1 #() 
OAI211_X1_832_ (
  .A({ S17210 }),
  .B({ S17028 }),
  .C1({ S17209 }),
  .C2({ S17072 }),
  .ZN({ S17211 })
);
NAND3_X1 #() 
NAND3_X1_2554_ (
  .A1({ S17207 }),
  .A2({ S16967 }),
  .A3({ S17211 }),
  .ZN({ S17212 })
);
NAND2_X1 #() 
NAND2_X1_2337_ (
  .A1({ S25957[131] }),
  .A2({ S17076 }),
  .ZN({ S17213 })
);
OAI211_X1 #() 
OAI211_X1_833_ (
  .A({ S17046 }),
  .B({ S17028 }),
  .C1({ S17032 }),
  .C2({ S17213 }),
  .ZN({ S17214 })
);
OAI211_X1 #() 
OAI211_X1_834_ (
  .A({ S17055 }),
  .B({ S25957[132] }),
  .C1({ S17036 }),
  .C2({ S17118 }),
  .ZN({ S17215 })
);
NAND3_X1 #() 
NAND3_X1_2555_ (
  .A1({ S17215 }),
  .A2({ S17214 }),
  .A3({ S25957[133] }),
  .ZN({ S17216 })
);
AND3_X1 #() 
AND3_X1_101_ (
  .A1({ S17216 }),
  .A2({ S17212 }),
  .A3({ S25957[134] }),
  .ZN({ S17217 })
);
OAI21_X1 #() 
OAI21_X1_1234_ (
  .A({ S25957[135] }),
  .B1({ S17204 }),
  .B2({ S17217 }),
  .ZN({ S17218 })
);
OAI21_X1 #() 
OAI21_X1_1235_ (
  .A({ S25957[132] }),
  .B1({ S16986 }),
  .B2({ S51 }),
  .ZN({ S17220 })
);
NAND2_X1 #() 
NAND2_X1_2338_ (
  .A1({ S25957[132] }),
  .A2({ S16969 }),
  .ZN({ S17221 })
);
AOI22_X1 #() 
AOI22_X1_291_ (
  .A1({ S17220 }),
  .A2({ S17221 }),
  .B1({ S17171 }),
  .B2({ S16988 }),
  .ZN({ S17222 })
);
NAND3_X1 #() 
NAND3_X1_2556_ (
  .A1({ S16961 }),
  .A2({ S16962 }),
  .A3({ S16969 }),
  .ZN({ S17223 })
);
INV_X1 #() 
INV_X1_743_ (
  .A({ S17223 }),
  .ZN({ S17224 })
);
OAI21_X1 #() 
OAI21_X1_1236_ (
  .A({ S25957[131] }),
  .B1({ S17112 }),
  .B2({ S17224 }),
  .ZN({ S17225 })
);
AOI21_X1 #() 
AOI21_X1_1338_ (
  .A({ S25957[132] }),
  .B1({ S17225 }),
  .B2({ S17198 }),
  .ZN({ S17226 })
);
OAI21_X1 #() 
OAI21_X1_1237_ (
  .A({ S25957[133] }),
  .B1({ S17226 }),
  .B2({ S17222 }),
  .ZN({ S17227 })
);
OAI21_X1 #() 
OAI21_X1_1238_ (
  .A({ S25957[129] }),
  .B1({ S17036 }),
  .B2({ S16969 }),
  .ZN({ S17228 })
);
NAND2_X1 #() 
NAND2_X1_2339_ (
  .A1({ S17228 }),
  .A2({ S51 }),
  .ZN({ S17229 })
);
AOI22_X1 #() 
AOI22_X1_292_ (
  .A1({ S17005 }),
  .A2({ S17055 }),
  .B1({ S17195 }),
  .B2({ S17229 }),
  .ZN({ S17231 })
);
NAND2_X1 #() 
NAND2_X1_2340_ (
  .A1({ S17231 }),
  .A2({ S16967 }),
  .ZN({ S17232 })
);
NAND3_X1 #() 
NAND3_X1_2557_ (
  .A1({ S17232 }),
  .A2({ S17227 }),
  .A3({ S15041 }),
  .ZN({ S17233 })
);
NAND2_X1 #() 
NAND2_X1_2341_ (
  .A1({ S17053 }),
  .A2({ S25957[131] }),
  .ZN({ S17234 })
);
INV_X1 #() 
INV_X1_744_ (
  .A({ S17234 }),
  .ZN({ S17235 })
);
NAND2_X1 #() 
NAND2_X1_2342_ (
  .A1({ S17235 }),
  .A2({ S16988 }),
  .ZN({ S17236 })
);
AOI21_X1 #() 
AOI21_X1_1339_ (
  .A({ S25957[132] }),
  .B1({ S17073 }),
  .B2({ S17079 }),
  .ZN({ S17237 })
);
NAND3_X1 #() 
NAND3_X1_2558_ (
  .A1({ S51 }),
  .A2({ S16963 }),
  .A3({ S16999 }),
  .ZN({ S17238 })
);
OAI21_X1 #() 
OAI21_X1_1239_ (
  .A({ S17238 }),
  .B1({ S17118 }),
  .B2({ S17135 }),
  .ZN({ S17239 })
);
AOI22_X1 #() 
AOI22_X1_293_ (
  .A1({ S17236 }),
  .A2({ S17237 }),
  .B1({ S25957[132] }),
  .B2({ S17239 }),
  .ZN({ S17240 })
);
NOR2_X1 #() 
NOR2_X1_564_ (
  .A1({ S17194 }),
  .A2({ S17054 }),
  .ZN({ S17242 })
);
NAND2_X1 #() 
NAND2_X1_2343_ (
  .A1({ S17002 }),
  .A2({ S51 }),
  .ZN({ S17243 })
);
NAND2_X1 #() 
NAND2_X1_2344_ (
  .A1({ S17243 }),
  .A2({ S17028 }),
  .ZN({ S17244 })
);
NAND2_X1 #() 
NAND2_X1_2345_ (
  .A1({ S17238 }),
  .A2({ S25957[132] }),
  .ZN({ S17245 })
);
OAI21_X1 #() 
OAI21_X1_1240_ (
  .A({ S17046 }),
  .B1({ S17000 }),
  .B2({ S51 }),
  .ZN({ S17246 })
);
OAI221_X1 #() 
OAI221_X1_55_ (
  .A({ S16967 }),
  .B1({ S17245 }),
  .B2({ S17246 }),
  .C1({ S17244 }),
  .C2({ S17242 }),
  .ZN({ S17247 })
);
OAI21_X1 #() 
OAI21_X1_1241_ (
  .A({ S17247 }),
  .B1({ S17240 }),
  .B2({ S16967 }),
  .ZN({ S17248 })
);
OAI211_X1 #() 
OAI211_X1_835_ (
  .A({ S16966 }),
  .B({ S17233 }),
  .C1({ S17248 }),
  .C2({ S15041 }),
  .ZN({ S17249 })
);
NAND2_X1 #() 
NAND2_X1_2346_ (
  .A1({ S17249 }),
  .A2({ S17218 }),
  .ZN({ S17250 })
);
XNOR2_X1 #() 
XNOR2_X1_128_ (
  .A({ S17250 }),
  .B({ S25957[234] }),
  .ZN({ S25957[106] })
);
INV_X1 #() 
INV_X1_745_ (
  .A({ S25957[235] }),
  .ZN({ S17252 })
);
NAND3_X1 #() 
NAND3_X1_2559_ (
  .A1({ S17029 }),
  .A2({ S60 }),
  .A3({ S17030 }),
  .ZN({ S17253 })
);
NAND3_X1 #() 
NAND3_X1_2560_ (
  .A1({ S51 }),
  .A2({ S16984 }),
  .A3({ S16999 }),
  .ZN({ S17254 })
);
OAI211_X1 #() 
OAI211_X1_836_ (
  .A({ S17028 }),
  .B({ S17254 }),
  .C1({ S17253 }),
  .C2({ S51 }),
  .ZN({ S17255 })
);
AOI21_X1 #() 
AOI21_X1_1340_ (
  .A({ S17028 }),
  .B1({ S16991 }),
  .B2({ S17071 }),
  .ZN({ S17256 })
);
OAI21_X1 #() 
OAI21_X1_1242_ (
  .A({ S17256 }),
  .B1({ S51 }),
  .B2({ S17032 }),
  .ZN({ S17257 })
);
NAND3_X1 #() 
NAND3_X1_2561_ (
  .A1({ S17257 }),
  .A2({ S16967 }),
  .A3({ S17255 }),
  .ZN({ S17258 })
);
AOI21_X1 #() 
AOI21_X1_1341_ (
  .A({ S16989 }),
  .B1({ S16963 }),
  .B2({ S60 }),
  .ZN({ S17259 })
);
NAND2_X1 #() 
NAND2_X1_2347_ (
  .A1({ S17173 }),
  .A2({ S25957[131] }),
  .ZN({ S17260 })
);
OAI21_X1 #() 
OAI21_X1_1243_ (
  .A({ S17260 }),
  .B1({ S17259 }),
  .B2({ S17136 }),
  .ZN({ S17261 })
);
NAND2_X1 #() 
NAND2_X1_2348_ (
  .A1({ S17261 }),
  .A2({ S17028 }),
  .ZN({ S17263 })
);
NOR2_X1 #() 
NOR2_X1_565_ (
  .A1({ S17070 }),
  .A2({ S51 }),
  .ZN({ S17264 })
);
NAND2_X1 #() 
NAND2_X1_2349_ (
  .A1({ S17264 }),
  .A2({ S17053 }),
  .ZN({ S17265 })
);
AOI21_X1 #() 
AOI21_X1_1342_ (
  .A({ S17028 }),
  .B1({ S16997 }),
  .B2({ S17014 }),
  .ZN({ S17266 })
);
AOI21_X1 #() 
AOI21_X1_1343_ (
  .A({ S16967 }),
  .B1({ S17265 }),
  .B2({ S17266 }),
  .ZN({ S17267 })
);
AOI21_X1 #() 
AOI21_X1_1344_ (
  .A({ S25957[134] }),
  .B1({ S17263 }),
  .B2({ S17267 }),
  .ZN({ S17268 })
);
OAI21_X1 #() 
OAI21_X1_1244_ (
  .A({ S16992 }),
  .B1({ S51 }),
  .B2({ S25957[129] }),
  .ZN({ S17269 })
);
OAI21_X1 #() 
OAI21_X1_1245_ (
  .A({ S25957[132] }),
  .B1({ S17031 }),
  .B2({ S17269 }),
  .ZN({ S17270 })
);
NAND2_X1 #() 
NAND2_X1_2350_ (
  .A1({ S16984 }),
  .A2({ S16999 }),
  .ZN({ S17271 })
);
NOR2_X1 #() 
NOR2_X1_566_ (
  .A1({ S17209 }),
  .A2({ S25957[132] }),
  .ZN({ S17272 })
);
NAND2_X1 #() 
NAND2_X1_2351_ (
  .A1({ S17272 }),
  .A2({ S17271 }),
  .ZN({ S17274 })
);
NAND3_X1 #() 
NAND3_X1_2562_ (
  .A1({ S17270 }),
  .A2({ S16967 }),
  .A3({ S17274 }),
  .ZN({ S17275 })
);
OAI211_X1 #() 
OAI211_X1_837_ (
  .A({ S51 }),
  .B({ S16963 }),
  .C1({ S60 }),
  .C2({ S25957[130] }),
  .ZN({ S17276 })
);
OAI211_X1 #() 
OAI211_X1_838_ (
  .A({ S17028 }),
  .B({ S17276 }),
  .C1({ S17061 }),
  .C2({ S51 }),
  .ZN({ S17277 })
);
NAND3_X1 #() 
NAND3_X1_2563_ (
  .A1({ S17076 }),
  .A2({ S51 }),
  .A3({ S16987 }),
  .ZN({ S17278 })
);
AOI21_X1 #() 
AOI21_X1_1345_ (
  .A({ S17028 }),
  .B1({ S17020 }),
  .B2({ S25957[131] }),
  .ZN({ S17279 })
);
AOI21_X1 #() 
AOI21_X1_1346_ (
  .A({ S16967 }),
  .B1({ S17279 }),
  .B2({ S17278 }),
  .ZN({ S17280 })
);
AOI21_X1 #() 
AOI21_X1_1347_ (
  .A({ S15041 }),
  .B1({ S17280 }),
  .B2({ S17277 }),
  .ZN({ S17281 })
);
AOI22_X1 #() 
AOI22_X1_294_ (
  .A1({ S17258 }),
  .A2({ S17268 }),
  .B1({ S17281 }),
  .B2({ S17275 }),
  .ZN({ S17282 })
);
NAND4_X1 #() 
NAND4_X1_313_ (
  .A1({ S17029 }),
  .A2({ S17030 }),
  .A3({ S60 }),
  .A4({ S16992 }),
  .ZN({ S17283 })
);
INV_X1 #() 
INV_X1_746_ (
  .A({ S17014 }),
  .ZN({ S17285 })
);
OAI21_X1 #() 
OAI21_X1_1246_ (
  .A({ S25957[132] }),
  .B1({ S17285 }),
  .B2({ S16993 }),
  .ZN({ S17286 })
);
AOI21_X1 #() 
AOI21_X1_1348_ (
  .A({ S17286 }),
  .B1({ S17283 }),
  .B2({ S51 }),
  .ZN({ S17287 })
);
AOI22_X1 #() 
AOI22_X1_295_ (
  .A1({ S60 }),
  .A2({ S17199 }),
  .B1({ S15306 }),
  .B2({ S15302 }),
  .ZN({ S17288 })
);
OAI21_X1 #() 
OAI21_X1_1247_ (
  .A({ S25957[133] }),
  .B1({ S17087 }),
  .B2({ S17288 }),
  .ZN({ S17289 })
);
NAND2_X1 #() 
NAND2_X1_2352_ (
  .A1({ S17057 }),
  .A2({ S17028 }),
  .ZN({ S17290 })
);
OAI211_X1 #() 
OAI211_X1_839_ (
  .A({ S16967 }),
  .B({ S17245 }),
  .C1({ S17290 }),
  .C2({ S17188 }),
  .ZN({ S17291 })
);
OAI211_X1 #() 
OAI211_X1_840_ (
  .A({ S17291 }),
  .B({ S25957[134] }),
  .C1({ S17287 }),
  .C2({ S17289 }),
  .ZN({ S17292 })
);
NAND2_X1 #() 
NAND2_X1_2353_ (
  .A1({ S25957[131] }),
  .A2({ S17037 }),
  .ZN({ S17293 })
);
OAI21_X1 #() 
OAI21_X1_1248_ (
  .A({ S17293 }),
  .B1({ S17259 }),
  .B2({ S25957[131] }),
  .ZN({ S17294 })
);
NAND3_X1 #() 
NAND3_X1_2564_ (
  .A1({ S51 }),
  .A2({ S16987 }),
  .A3({ S16999 }),
  .ZN({ S17296 })
);
AOI21_X1 #() 
AOI21_X1_1349_ (
  .A({ S25957[132] }),
  .B1({ S17296 }),
  .B2({ S17015 }),
  .ZN({ S17297 })
);
AOI21_X1 #() 
AOI21_X1_1350_ (
  .A({ S17297 }),
  .B1({ S17294 }),
  .B2({ S25957[132] }),
  .ZN({ S17298 })
);
AOI21_X1 #() 
AOI21_X1_1351_ (
  .A({ S16989 }),
  .B1({ S16987 }),
  .B2({ S16984 }),
  .ZN({ S17299 })
);
NAND4_X1 #() 
NAND4_X1_314_ (
  .A1({ S17223 }),
  .A2({ S16985 }),
  .A3({ S15306 }),
  .A4({ S15302 }),
  .ZN({ S17300 })
);
OAI211_X1 #() 
OAI211_X1_841_ (
  .A({ S17028 }),
  .B({ S17300 }),
  .C1({ S17299 }),
  .C2({ S17151 }),
  .ZN({ S17301 })
);
NAND3_X1 #() 
NAND3_X1_2565_ (
  .A1({ S17205 }),
  .A2({ S51 }),
  .A3({ S17079 }),
  .ZN({ S17302 })
);
OAI211_X1 #() 
OAI211_X1_842_ (
  .A({ S25957[132] }),
  .B({ S17302 }),
  .C1({ S17156 }),
  .C2({ S51 }),
  .ZN({ S17303 })
);
NAND3_X1 #() 
NAND3_X1_2566_ (
  .A1({ S17301 }),
  .A2({ S17303 }),
  .A3({ S16967 }),
  .ZN({ S17304 })
);
OAI211_X1 #() 
OAI211_X1_843_ (
  .A({ S15041 }),
  .B({ S17304 }),
  .C1({ S17298 }),
  .C2({ S16967 }),
  .ZN({ S17305 })
);
NAND3_X1 #() 
NAND3_X1_2567_ (
  .A1({ S17305 }),
  .A2({ S16966 }),
  .A3({ S17292 }),
  .ZN({ S17307 })
);
OAI211_X1 #() 
OAI211_X1_844_ (
  .A({ S17307 }),
  .B({ S17252 }),
  .C1({ S17282 }),
  .C2({ S16966 }),
  .ZN({ S17308 })
);
NAND3_X1 #() 
NAND3_X1_2568_ (
  .A1({ S17257 }),
  .A2({ S15041 }),
  .A3({ S17255 }),
  .ZN({ S17309 })
);
AOI21_X1 #() 
AOI21_X1_1352_ (
  .A({ S15041 }),
  .B1({ S17272 }),
  .B2({ S17271 }),
  .ZN({ S17310 })
);
NAND2_X1 #() 
NAND2_X1_2354_ (
  .A1({ S17310 }),
  .A2({ S17270 }),
  .ZN({ S17311 })
);
AOI21_X1 #() 
AOI21_X1_1353_ (
  .A({ S16966 }),
  .B1({ S17311 }),
  .B2({ S17309 }),
  .ZN({ S17312 })
);
NAND2_X1 #() 
NAND2_X1_2355_ (
  .A1({ S51 }),
  .A2({ S16963 }),
  .ZN({ S17313 })
);
INV_X1 #() 
INV_X1_747_ (
  .A({ S17313 }),
  .ZN({ S17314 })
);
NAND3_X1 #() 
NAND3_X1_2569_ (
  .A1({ S17314 }),
  .A2({ S25957[132] }),
  .A3({ S16999 }),
  .ZN({ S17315 })
);
AND3_X1 #() 
AND3_X1_102_ (
  .A1({ S25957[131] }),
  .A2({ S16985 }),
  .A3({ S17030 }),
  .ZN({ S17316 })
);
OAI21_X1 #() 
OAI21_X1_1249_ (
  .A({ S17028 }),
  .B1({ S17316 }),
  .B2({ S17188 }),
  .ZN({ S17318 })
);
NAND3_X1 #() 
NAND3_X1_2570_ (
  .A1({ S17318 }),
  .A2({ S25957[134] }),
  .A3({ S17315 }),
  .ZN({ S17319 })
);
NAND2_X1 #() 
NAND2_X1_2356_ (
  .A1({ S17301 }),
  .A2({ S17303 }),
  .ZN({ S17320 })
);
NAND2_X1 #() 
NAND2_X1_2357_ (
  .A1({ S17320 }),
  .A2({ S15041 }),
  .ZN({ S17321 })
);
AOI21_X1 #() 
AOI21_X1_1354_ (
  .A({ S25957[135] }),
  .B1({ S17321 }),
  .B2({ S17319 }),
  .ZN({ S17322 })
);
OAI21_X1 #() 
OAI21_X1_1250_ (
  .A({ S16967 }),
  .B1({ S17322 }),
  .B2({ S17312 }),
  .ZN({ S17323 })
);
AOI22_X1 #() 
AOI22_X1_296_ (
  .A1({ S17283 }),
  .A2({ S51 }),
  .B1({ S16994 }),
  .B2({ S17014 }),
  .ZN({ S17324 })
);
NOR2_X1 #() 
NOR2_X1_567_ (
  .A1({ S16980 }),
  .A2({ S17044 }),
  .ZN({ S17325 })
);
OAI21_X1 #() 
OAI21_X1_1251_ (
  .A({ S17028 }),
  .B1({ S17288 }),
  .B2({ S17325 }),
  .ZN({ S17326 })
);
OAI211_X1 #() 
OAI211_X1_845_ (
  .A({ S17326 }),
  .B({ S25957[134] }),
  .C1({ S17324 }),
  .C2({ S17028 }),
  .ZN({ S17327 })
);
AOI21_X1 #() 
AOI21_X1_1355_ (
  .A({ S17264 }),
  .B1({ S16988 }),
  .B2({ S51 }),
  .ZN({ S17329 })
);
NAND2_X1 #() 
NAND2_X1_2358_ (
  .A1({ S17285 }),
  .A2({ S25957[131] }),
  .ZN({ S17330 })
);
AOI21_X1 #() 
AOI21_X1_1356_ (
  .A({ S25957[134] }),
  .B1({ S17237 }),
  .B2({ S17330 }),
  .ZN({ S17331 })
);
OAI21_X1 #() 
OAI21_X1_1252_ (
  .A({ S17331 }),
  .B1({ S17028 }),
  .B2({ S17329 }),
  .ZN({ S17332 })
);
AOI21_X1 #() 
AOI21_X1_1357_ (
  .A({ S25957[135] }),
  .B1({ S17327 }),
  .B2({ S17332 }),
  .ZN({ S17333 })
);
AOI22_X1 #() 
AOI22_X1_297_ (
  .A1({ S16988 }),
  .A2({ S17171 }),
  .B1({ S17173 }),
  .B2({ S25957[131] }),
  .ZN({ S17334 })
);
AOI21_X1 #() 
AOI21_X1_1358_ (
  .A({ S25957[130] }),
  .B1({ S16987 }),
  .B2({ S16984 }),
  .ZN({ S17335 })
);
OAI21_X1 #() 
OAI21_X1_1253_ (
  .A({ S17266 }),
  .B1({ S17335 }),
  .B2({ S17293 }),
  .ZN({ S17336 })
);
OAI211_X1 #() 
OAI211_X1_846_ (
  .A({ S17336 }),
  .B({ S15041 }),
  .C1({ S17334 }),
  .C2({ S25957[132] }),
  .ZN({ S17337 })
);
NAND3_X1 #() 
NAND3_X1_2571_ (
  .A1({ S17022 }),
  .A2({ S25957[132] }),
  .A3({ S17278 }),
  .ZN({ S17338 })
);
AOI21_X1 #() 
AOI21_X1_1359_ (
  .A({ S51 }),
  .B1({ S17000 }),
  .B2({ S17199 }),
  .ZN({ S17339 })
);
OAI21_X1 #() 
OAI21_X1_1254_ (
  .A({ S17028 }),
  .B1({ S17313 }),
  .B2({ S17047 }),
  .ZN({ S17340 })
);
OAI211_X1 #() 
OAI211_X1_847_ (
  .A({ S17338 }),
  .B({ S25957[134] }),
  .C1({ S17339 }),
  .C2({ S17340 }),
  .ZN({ S17341 })
);
AOI21_X1 #() 
AOI21_X1_1360_ (
  .A({ S16966 }),
  .B1({ S17337 }),
  .B2({ S17341 }),
  .ZN({ S17342 })
);
OAI21_X1 #() 
OAI21_X1_1255_ (
  .A({ S25957[133] }),
  .B1({ S17333 }),
  .B2({ S17342 }),
  .ZN({ S17343 })
);
NAND3_X1 #() 
NAND3_X1_2572_ (
  .A1({ S17323 }),
  .A2({ S17343 }),
  .A3({ S25957[235] }),
  .ZN({ S17344 })
);
NAND2_X1 #() 
NAND2_X1_2359_ (
  .A1({ S17344 }),
  .A2({ S17308 }),
  .ZN({ S25957[107] })
);
INV_X1 #() 
INV_X1_748_ (
  .A({ S25957[236] }),
  .ZN({ S17345 })
);
NOR3_X1 #() 
NOR3_X1_74_ (
  .A1({ S17196 }),
  .A2({ S17135 }),
  .A3({ S51 }),
  .ZN({ S17346 })
);
OR2_X1 #() 
OR2_X1_33_ (
  .A1({ S17062 }),
  .A2({ S17346 }),
  .ZN({ S17347 })
);
NOR2_X1 #() 
NOR2_X1_568_ (
  .A1({ S17082 }),
  .A2({ S25957[132] }),
  .ZN({ S17349 })
);
OAI21_X1 #() 
OAI21_X1_1256_ (
  .A({ S51 }),
  .B1({ S17112 }),
  .B2({ S17032 }),
  .ZN({ S17350 })
);
AOI21_X1 #() 
AOI21_X1_1361_ (
  .A({ S16967 }),
  .B1({ S17349 }),
  .B2({ S17350 }),
  .ZN({ S17351 })
);
NAND3_X1 #() 
NAND3_X1_2573_ (
  .A1({ S16978 }),
  .A2({ S25957[131] }),
  .A3({ S17079 }),
  .ZN({ S17352 })
);
OAI211_X1 #() 
OAI211_X1_848_ (
  .A({ S17229 }),
  .B({ S25957[132] }),
  .C1({ S17352 }),
  .C2({ S16972 }),
  .ZN({ S17353 })
);
NOR2_X1 #() 
NOR2_X1_569_ (
  .A1({ S51 }),
  .A2({ S25957[129] }),
  .ZN({ S17354 })
);
AOI21_X1 #() 
AOI21_X1_1362_ (
  .A({ S25957[132] }),
  .B1({ S17354 }),
  .B2({ S16999 }),
  .ZN({ S17355 })
);
AOI21_X1 #() 
AOI21_X1_1363_ (
  .A({ S25957[133] }),
  .B1({ S17355 }),
  .B2({ S17141 }),
  .ZN({ S17356 })
);
AOI22_X1 #() 
AOI22_X1_298_ (
  .A1({ S17351 }),
  .A2({ S17347 }),
  .B1({ S17353 }),
  .B2({ S17356 }),
  .ZN({ S17357 })
);
NAND2_X1 #() 
NAND2_X1_2360_ (
  .A1({ S17357 }),
  .A2({ S15041 }),
  .ZN({ S17358 })
);
OAI221_X1 #() 
OAI221_X1_56_ (
  .A({ S25957[132] }),
  .B1({ S25957[131] }),
  .B2({ S17070 }),
  .C1({ S25957[130] }),
  .C2({ S17135 }),
  .ZN({ S17360 })
);
NAND2_X1 #() 
NAND2_X1_2361_ (
  .A1({ S17161 }),
  .A2({ S25957[131] }),
  .ZN({ S17361 })
);
NAND3_X1 #() 
NAND3_X1_2574_ (
  .A1({ S17172 }),
  .A2({ S17028 }),
  .A3({ S17361 }),
  .ZN({ S17362 })
);
NAND3_X1 #() 
NAND3_X1_2575_ (
  .A1({ S17362 }),
  .A2({ S25957[133] }),
  .A3({ S17360 }),
  .ZN({ S17363 })
);
NAND3_X1 #() 
NAND3_X1_2576_ (
  .A1({ S25957[131] }),
  .A2({ S16987 }),
  .A3({ S17079 }),
  .ZN({ S17364 })
);
OAI21_X1 #() 
OAI21_X1_1257_ (
  .A({ S17364 }),
  .B1({ S17072 }),
  .B2({ S17175 }),
  .ZN({ S17365 })
);
NAND2_X1 #() 
NAND2_X1_2362_ (
  .A1({ S25957[131] }),
  .A2({ S16977 }),
  .ZN({ S17366 })
);
AND2_X1 #() 
AND2_X1_142_ (
  .A1({ S51 }),
  .A2({ S16984 }),
  .ZN({ S17367 })
);
NAND2_X1 #() 
NAND2_X1_2363_ (
  .A1({ S17367 }),
  .A2({ S16991 }),
  .ZN({ S17368 })
);
OAI211_X1 #() 
OAI211_X1_849_ (
  .A({ S17368 }),
  .B({ S25957[132] }),
  .C1({ S16969 }),
  .C2({ S17366 }),
  .ZN({ S17369 })
);
OAI211_X1 #() 
OAI211_X1_850_ (
  .A({ S17369 }),
  .B({ S16967 }),
  .C1({ S17365 }),
  .C2({ S25957[132] }),
  .ZN({ S17371 })
);
NAND3_X1 #() 
NAND3_X1_2577_ (
  .A1({ S17371 }),
  .A2({ S25957[134] }),
  .A3({ S17363 }),
  .ZN({ S17372 })
);
AND2_X1 #() 
AND2_X1_143_ (
  .A1({ S17372 }),
  .A2({ S25957[135] }),
  .ZN({ S17373 })
);
NAND2_X1 #() 
NAND2_X1_2364_ (
  .A1({ S17358 }),
  .A2({ S17373 }),
  .ZN({ S17374 })
);
NAND2_X1 #() 
NAND2_X1_2365_ (
  .A1({ S17050 }),
  .A2({ S51 }),
  .ZN({ S17375 })
);
NAND2_X1 #() 
NAND2_X1_2366_ (
  .A1({ S17205 }),
  .A2({ S17079 }),
  .ZN({ S17376 })
);
NAND2_X1 #() 
NAND2_X1_2367_ (
  .A1({ S17376 }),
  .A2({ S25957[131] }),
  .ZN({ S17377 })
);
AOI21_X1 #() 
AOI21_X1_1364_ (
  .A({ S17028 }),
  .B1({ S17377 }),
  .B2({ S17375 }),
  .ZN({ S17378 })
);
NOR3_X1 #() 
NOR3_X1_75_ (
  .A1({ S17235 }),
  .A2({ S17314 }),
  .A3({ S25957[132] }),
  .ZN({ S17379 })
);
OAI21_X1 #() 
OAI21_X1_1258_ (
  .A({ S25957[133] }),
  .B1({ S17379 }),
  .B2({ S17378 }),
  .ZN({ S17380 })
);
OAI211_X1 #() 
OAI211_X1_851_ (
  .A({ S17057 }),
  .B({ S25957[132] }),
  .C1({ S17003 }),
  .C2({ S17313 }),
  .ZN({ S17382 })
);
NAND2_X1 #() 
NAND2_X1_2368_ (
  .A1({ S17022 }),
  .A2({ S17028 }),
  .ZN({ S17383 })
);
OAI211_X1 #() 
OAI211_X1_852_ (
  .A({ S17382 }),
  .B({ S16967 }),
  .C1({ S17049 }),
  .C2({ S17383 }),
  .ZN({ S17384 })
);
NAND3_X1 #() 
NAND3_X1_2578_ (
  .A1({ S17380 }),
  .A2({ S15041 }),
  .A3({ S17384 }),
  .ZN({ S17385 })
);
NAND2_X1 #() 
NAND2_X1_2369_ (
  .A1({ S51 }),
  .A2({ S17223 }),
  .ZN({ S17386 })
);
OAI21_X1 #() 
OAI21_X1_1259_ (
  .A({ S17272 }),
  .B1({ S17036 }),
  .B2({ S17386 }),
  .ZN({ S17387 })
);
INV_X1 #() 
INV_X1_749_ (
  .A({ S17054 }),
  .ZN({ S17388 })
);
INV_X1 #() 
INV_X1_750_ (
  .A({ S17161 }),
  .ZN({ S17389 })
);
OAI21_X1 #() 
OAI21_X1_1260_ (
  .A({ S17149 }),
  .B1({ S17388 }),
  .B2({ S17389 }),
  .ZN({ S17390 })
);
OAI21_X1 #() 
OAI21_X1_1261_ (
  .A({ S17387 }),
  .B1({ S17028 }),
  .B2({ S17390 }),
  .ZN({ S17391 })
);
INV_X1 #() 
INV_X1_751_ (
  .A({ S153 }),
  .ZN({ S17393 })
);
OAI21_X1 #() 
OAI21_X1_1262_ (
  .A({ S25957[132] }),
  .B1({ S17393 }),
  .B2({ S25957[130] }),
  .ZN({ S17394 })
);
OAI21_X1 #() 
OAI21_X1_1263_ (
  .A({ S17065 }),
  .B1({ S17032 }),
  .B2({ S17109 }),
  .ZN({ S17395 })
);
NAND3_X1 #() 
NAND3_X1_2579_ (
  .A1({ S17395 }),
  .A2({ S25957[133] }),
  .A3({ S17394 }),
  .ZN({ S17396 })
);
OAI211_X1 #() 
OAI211_X1_853_ (
  .A({ S25957[134] }),
  .B({ S17396 }),
  .C1({ S17391 }),
  .C2({ S25957[133] }),
  .ZN({ S17397 })
);
NAND3_X1 #() 
NAND3_X1_2580_ (
  .A1({ S17385 }),
  .A2({ S17397 }),
  .A3({ S16966 }),
  .ZN({ S17398 })
);
NAND3_X1 #() 
NAND3_X1_2581_ (
  .A1({ S17374 }),
  .A2({ S17398 }),
  .A3({ S17345 }),
  .ZN({ S17399 })
);
NAND2_X1 #() 
NAND2_X1_2370_ (
  .A1({ S17385 }),
  .A2({ S17397 }),
  .ZN({ S17400 })
);
NAND2_X1 #() 
NAND2_X1_2371_ (
  .A1({ S17400 }),
  .A2({ S16966 }),
  .ZN({ S17401 })
);
NAND2_X1 #() 
NAND2_X1_2372_ (
  .A1({ S17371 }),
  .A2({ S17363 }),
  .ZN({ S17402 })
);
NAND2_X1 #() 
NAND2_X1_2373_ (
  .A1({ S17402 }),
  .A2({ S25957[134] }),
  .ZN({ S17404 })
);
OAI211_X1 #() 
OAI211_X1_854_ (
  .A({ S25957[135] }),
  .B({ S17404 }),
  .C1({ S17357 }),
  .C2({ S25957[134] }),
  .ZN({ S17405 })
);
NAND3_X1 #() 
NAND3_X1_2582_ (
  .A1({ S17405 }),
  .A2({ S17401 }),
  .A3({ S25957[236] }),
  .ZN({ S17406 })
);
NAND2_X1 #() 
NAND2_X1_2374_ (
  .A1({ S17399 }),
  .A2({ S17406 }),
  .ZN({ S25957[108] })
);
NAND2_X1 #() 
NAND2_X1_2375_ (
  .A1({ S17228 }),
  .A2({ S25957[131] }),
  .ZN({ S17407 })
);
NAND3_X1 #() 
NAND3_X1_2583_ (
  .A1({ S17407 }),
  .A2({ S16973 }),
  .A3({ S17028 }),
  .ZN({ S17408 })
);
NOR2_X1 #() 
NOR2_X1_570_ (
  .A1({ S17081 }),
  .A2({ S25957[131] }),
  .ZN({ S17409 })
);
OAI21_X1 #() 
OAI21_X1_1264_ (
  .A({ S17408 }),
  .B1({ S17409 }),
  .B2({ S17220 }),
  .ZN({ S17410 })
);
NOR2_X1 #() 
NOR2_X1_571_ (
  .A1({ S16988 }),
  .A2({ S25957[131] }),
  .ZN({ S17411 })
);
OAI21_X1 #() 
OAI21_X1_1265_ (
  .A({ S17028 }),
  .B1({ S17285 }),
  .B2({ S16993 }),
  .ZN({ S17412 })
);
OAI211_X1 #() 
OAI211_X1_855_ (
  .A({ S17050 }),
  .B({ S25957[132] }),
  .C1({ S51 }),
  .C2({ S16984 }),
  .ZN({ S17414 })
);
OAI211_X1 #() 
OAI211_X1_856_ (
  .A({ S16967 }),
  .B({ S17414 }),
  .C1({ S17411 }),
  .C2({ S17412 }),
  .ZN({ S17415 })
);
OAI211_X1 #() 
OAI211_X1_857_ (
  .A({ S25957[134] }),
  .B({ S17415 }),
  .C1({ S17410 }),
  .C2({ S16967 }),
  .ZN({ S17416 })
);
OAI21_X1 #() 
OAI21_X1_1266_ (
  .A({ S17234 }),
  .B1({ S17206 }),
  .B2({ S25957[131] }),
  .ZN({ S17417 })
);
OAI21_X1 #() 
OAI21_X1_1267_ (
  .A({ S25957[131] }),
  .B1({ S17299 }),
  .B2({ S17047 }),
  .ZN({ S17418 })
);
NAND3_X1 #() 
NAND3_X1_2584_ (
  .A1({ S17418 }),
  .A2({ S17028 }),
  .A3({ S17386 }),
  .ZN({ S17419 })
);
OAI21_X1 #() 
OAI21_X1_1268_ (
  .A({ S17419 }),
  .B1({ S17028 }),
  .B2({ S17417 }),
  .ZN({ S17420 })
);
NAND3_X1 #() 
NAND3_X1_2585_ (
  .A1({ S17368 }),
  .A2({ S17028 }),
  .A3({ S17366 }),
  .ZN({ S17421 })
);
OAI221_X1 #() 
OAI221_X1_57_ (
  .A({ S25957[132] }),
  .B1({ S16998 }),
  .B2({ S59 }),
  .C1({ S17352 }),
  .C2({ S16964 }),
  .ZN({ S17422 })
);
NAND3_X1 #() 
NAND3_X1_2586_ (
  .A1({ S17422 }),
  .A2({ S25957[133] }),
  .A3({ S17421 }),
  .ZN({ S17423 })
);
OAI211_X1 #() 
OAI211_X1_858_ (
  .A({ S17423 }),
  .B({ S15041 }),
  .C1({ S17420 }),
  .C2({ S25957[133] }),
  .ZN({ S17425 })
);
NAND3_X1 #() 
NAND3_X1_2587_ (
  .A1({ S17425 }),
  .A2({ S25957[135] }),
  .A3({ S17416 }),
  .ZN({ S17426 })
);
AOI22_X1 #() 
AOI22_X1_299_ (
  .A1({ S17119 }),
  .A2({ S17117 }),
  .B1({ S17376 }),
  .B2({ S51 }),
  .ZN({ S17427 })
);
AND2_X1 #() 
AND2_X1_144_ (
  .A1({ S17427 }),
  .A2({ S25957[132] }),
  .ZN({ S17428 })
);
OAI21_X1 #() 
OAI21_X1_1269_ (
  .A({ S16980 }),
  .B1({ S17020 }),
  .B2({ S25957[131] }),
  .ZN({ S17429 })
);
OAI21_X1 #() 
OAI21_X1_1270_ (
  .A({ S25957[133] }),
  .B1({ S17429 }),
  .B2({ S25957[132] }),
  .ZN({ S17430 })
);
NAND3_X1 #() 
NAND3_X1_2588_ (
  .A1({ S16970 }),
  .A2({ S51 }),
  .A3({ S17223 }),
  .ZN({ S17431 })
);
NOR2_X1 #() 
NOR2_X1_572_ (
  .A1({ S17209 }),
  .A2({ S17028 }),
  .ZN({ S17432 })
);
NAND3_X1 #() 
NAND3_X1_2589_ (
  .A1({ S17432 }),
  .A2({ S17431 }),
  .A3({ S17210 }),
  .ZN({ S17433 })
);
OAI211_X1 #() 
OAI211_X1_859_ (
  .A({ S16967 }),
  .B({ S17433 }),
  .C1({ S17244 }),
  .C2({ S17064 }),
  .ZN({ S17434 })
);
OAI211_X1 #() 
OAI211_X1_860_ (
  .A({ S25957[134] }),
  .B({ S17434 }),
  .C1({ S17428 }),
  .C2({ S17430 }),
  .ZN({ S17436 })
);
AOI21_X1 #() 
AOI21_X1_1365_ (
  .A({ S16994 }),
  .B1({ S17010 }),
  .B2({ S51 }),
  .ZN({ S17437 })
);
OAI21_X1 #() 
OAI21_X1_1271_ (
  .A({ S25957[132] }),
  .B1({ S17253 }),
  .B2({ S51 }),
  .ZN({ S17438 })
);
OAI211_X1 #() 
OAI211_X1_861_ (
  .A({ S25957[128] }),
  .B({ S17028 }),
  .C1({ S17122 }),
  .C2({ S17354 }),
  .ZN({ S17439 })
);
OAI211_X1 #() 
OAI211_X1_862_ (
  .A({ S17439 }),
  .B({ S16967 }),
  .C1({ S17437 }),
  .C2({ S17438 }),
  .ZN({ S17440 })
);
INV_X1 #() 
INV_X1_752_ (
  .A({ S17126 }),
  .ZN({ S17441 })
);
AOI22_X1 #() 
AOI22_X1_300_ (
  .A1({ S17441 }),
  .A2({ S16989 }),
  .B1({ S51 }),
  .B2({ S16976 }),
  .ZN({ S17442 })
);
NAND2_X1 #() 
NAND2_X1_2376_ (
  .A1({ S25957[131] }),
  .A2({ S16972 }),
  .ZN({ S17443 })
);
OAI21_X1 #() 
OAI21_X1_1272_ (
  .A({ S17443 }),
  .B1({ S25957[131] }),
  .B2({ S17173 }),
  .ZN({ S17444 })
);
NAND2_X1 #() 
NAND2_X1_2377_ (
  .A1({ S17444 }),
  .A2({ S17028 }),
  .ZN({ S17445 })
);
OAI21_X1 #() 
OAI21_X1_1273_ (
  .A({ S17445 }),
  .B1({ S17442 }),
  .B2({ S17028 }),
  .ZN({ S17447 })
);
OAI21_X1 #() 
OAI21_X1_1274_ (
  .A({ S17440 }),
  .B1({ S17447 }),
  .B2({ S16967 }),
  .ZN({ S17448 })
);
NAND2_X1 #() 
NAND2_X1_2378_ (
  .A1({ S17448 }),
  .A2({ S15041 }),
  .ZN({ S17449 })
);
NAND3_X1 #() 
NAND3_X1_2590_ (
  .A1({ S17436 }),
  .A2({ S16966 }),
  .A3({ S17449 }),
  .ZN({ S17450 })
);
NAND3_X1 #() 
NAND3_X1_2591_ (
  .A1({ S17450 }),
  .A2({ S17426 }),
  .A3({ S14448 }),
  .ZN({ S17451 })
);
NAND2_X1 #() 
NAND2_X1_2379_ (
  .A1({ S17425 }),
  .A2({ S17416 }),
  .ZN({ S17452 })
);
NAND2_X1 #() 
NAND2_X1_2380_ (
  .A1({ S17452 }),
  .A2({ S25957[135] }),
  .ZN({ S17453 })
);
OAI21_X1 #() 
OAI21_X1_1275_ (
  .A({ S17433 }),
  .B1({ S17244 }),
  .B2({ S17064 }),
  .ZN({ S17454 })
);
NAND2_X1 #() 
NAND2_X1_2381_ (
  .A1({ S17454 }),
  .A2({ S16967 }),
  .ZN({ S17455 })
);
NAND2_X1 #() 
NAND2_X1_2382_ (
  .A1({ S17429 }),
  .A2({ S17028 }),
  .ZN({ S17456 })
);
OAI211_X1 #() 
OAI211_X1_863_ (
  .A({ S25957[133] }),
  .B({ S17456 }),
  .C1({ S17427 }),
  .C2({ S17028 }),
  .ZN({ S17458 })
);
NAND3_X1 #() 
NAND3_X1_2592_ (
  .A1({ S17455 }),
  .A2({ S17458 }),
  .A3({ S25957[134] }),
  .ZN({ S17459 })
);
OAI211_X1 #() 
OAI211_X1_864_ (
  .A({ S17459 }),
  .B({ S16966 }),
  .C1({ S25957[134] }),
  .C2({ S17448 }),
  .ZN({ S17460 })
);
NAND3_X1 #() 
NAND3_X1_2593_ (
  .A1({ S17453 }),
  .A2({ S17460 }),
  .A3({ S25957[237] }),
  .ZN({ S17461 })
);
NAND2_X1 #() 
NAND2_X1_2383_ (
  .A1({ S17461 }),
  .A2({ S17451 }),
  .ZN({ S25957[109] })
);
INV_X1 #() 
INV_X1_753_ (
  .A({ S25957[238] }),
  .ZN({ S17462 })
);
OAI221_X1 #() 
OAI221_X1_58_ (
  .A({ S17028 }),
  .B1({ S16977 }),
  .B2({ S25957[131] }),
  .C1({ S17126 }),
  .C2({ S17003 }),
  .ZN({ S17463 })
);
NAND3_X1 #() 
NAND3_X1_2594_ (
  .A1({ S17017 }),
  .A2({ S25957[132] }),
  .A3({ S17185 }),
  .ZN({ S17464 })
);
NAND3_X1 #() 
NAND3_X1_2595_ (
  .A1({ S17464 }),
  .A2({ S25957[133] }),
  .A3({ S17463 }),
  .ZN({ S17465 })
);
NOR2_X1 #() 
NOR2_X1_573_ (
  .A1({ S17032 }),
  .A2({ S17175 }),
  .ZN({ S17466 })
);
NOR2_X1 #() 
NOR2_X1_574_ (
  .A1({ S17466 }),
  .A2({ S17286 }),
  .ZN({ S17468 })
);
AND2_X1 #() 
AND2_X1_145_ (
  .A1({ S17190 }),
  .A2({ S17167 }),
  .ZN({ S17469 })
);
AOI21_X1 #() 
AOI21_X1_1366_ (
  .A({ S17468 }),
  .B1({ S17469 }),
  .B2({ S17201 }),
  .ZN({ S17470 })
);
NAND2_X1 #() 
NAND2_X1_2384_ (
  .A1({ S17470 }),
  .A2({ S16967 }),
  .ZN({ S17471 })
);
NAND3_X1 #() 
NAND3_X1_2596_ (
  .A1({ S17471 }),
  .A2({ S25957[134] }),
  .A3({ S17465 }),
  .ZN({ S17472 })
);
NAND3_X1 #() 
NAND3_X1_2597_ (
  .A1({ S16991 }),
  .A2({ S17113 }),
  .A3({ S25957[131] }),
  .ZN({ S17473 })
);
OAI211_X1 #() 
OAI211_X1_865_ (
  .A({ S17028 }),
  .B({ S17473 }),
  .C1({ S17035 }),
  .C2({ S25957[131] }),
  .ZN({ S17474 })
);
NAND2_X1 #() 
NAND2_X1_2385_ (
  .A1({ S16984 }),
  .A2({ S16989 }),
  .ZN({ S17475 })
);
NOR2_X1 #() 
NOR2_X1_575_ (
  .A1({ S17299 }),
  .A2({ S25957[131] }),
  .ZN({ S17476 })
);
NAND2_X1 #() 
NAND2_X1_2386_ (
  .A1({ S17476 }),
  .A2({ S17475 }),
  .ZN({ S17477 })
);
NAND3_X1 #() 
NAND3_X1_2598_ (
  .A1({ S17477 }),
  .A2({ S25957[132] }),
  .A3({ S17088 }),
  .ZN({ S17479 })
);
NAND3_X1 #() 
NAND3_X1_2599_ (
  .A1({ S17479 }),
  .A2({ S17474 }),
  .A3({ S25957[133] }),
  .ZN({ S17480 })
);
INV_X1 #() 
INV_X1_754_ (
  .A({ S17149 }),
  .ZN({ S17481 })
);
AOI21_X1 #() 
AOI21_X1_1367_ (
  .A({ S17481 }),
  .B1({ S17080 }),
  .B2({ S51 }),
  .ZN({ S17482 })
);
NOR2_X1 #() 
NOR2_X1_576_ (
  .A1({ S17085 }),
  .A2({ S51 }),
  .ZN({ S17483 })
);
NOR2_X1 #() 
NOR2_X1_577_ (
  .A1({ S17483 }),
  .A2({ S17466 }),
  .ZN({ S17484 })
);
NAND2_X1 #() 
NAND2_X1_2387_ (
  .A1({ S17484 }),
  .A2({ S17028 }),
  .ZN({ S17485 })
);
OAI211_X1 #() 
OAI211_X1_866_ (
  .A({ S17485 }),
  .B({ S16967 }),
  .C1({ S17028 }),
  .C2({ S17482 }),
  .ZN({ S17486 })
);
NAND3_X1 #() 
NAND3_X1_2600_ (
  .A1({ S17486 }),
  .A2({ S15041 }),
  .A3({ S17480 }),
  .ZN({ S17487 })
);
NAND3_X1 #() 
NAND3_X1_2601_ (
  .A1({ S17472 }),
  .A2({ S25957[135] }),
  .A3({ S17487 }),
  .ZN({ S17488 })
);
NAND3_X1 #() 
NAND3_X1_2602_ (
  .A1({ S17125 }),
  .A2({ S17144 }),
  .A3({ S25957[132] }),
  .ZN({ S17490 })
);
OAI21_X1 #() 
OAI21_X1_1276_ (
  .A({ S17490 }),
  .B1({ S17476 }),
  .B2({ S17412 }),
  .ZN({ S17491 })
);
AOI21_X1 #() 
AOI21_X1_1368_ (
  .A({ S51 }),
  .B1({ S16984 }),
  .B2({ S16999 }),
  .ZN({ S17492 })
);
NOR3_X1 #() 
NOR3_X1_76_ (
  .A1({ S17152 }),
  .A2({ S17492 }),
  .A3({ S17028 }),
  .ZN({ S17493 })
);
AOI21_X1 #() 
AOI21_X1_1369_ (
  .A({ S25957[132] }),
  .B1({ S17443 }),
  .B2({ S17193 }),
  .ZN({ S17494 })
);
OAI21_X1 #() 
OAI21_X1_1277_ (
  .A({ S25957[133] }),
  .B1({ S17493 }),
  .B2({ S17494 }),
  .ZN({ S17495 })
);
OAI21_X1 #() 
OAI21_X1_1278_ (
  .A({ S17495 }),
  .B1({ S25957[133] }),
  .B2({ S17491 }),
  .ZN({ S17496 })
);
OAI21_X1 #() 
OAI21_X1_1279_ (
  .A({ S17151 }),
  .B1({ S17293 }),
  .B2({ S59 }),
  .ZN({ S17497 })
);
NAND2_X1 #() 
NAND2_X1_2388_ (
  .A1({ S17497 }),
  .A2({ S25957[132] }),
  .ZN({ S17498 })
);
NAND2_X1 #() 
NAND2_X1_2389_ (
  .A1({ S17376 }),
  .A2({ S51 }),
  .ZN({ S17499 })
);
AND2_X1 #() 
AND2_X1_146_ (
  .A1({ S17499 }),
  .A2({ S17352 }),
  .ZN({ S17501 })
);
OAI211_X1 #() 
OAI211_X1_867_ (
  .A({ S17498 }),
  .B({ S25957[133] }),
  .C1({ S17501 }),
  .C2({ S25957[132] }),
  .ZN({ S17502 })
);
AND2_X1 #() 
AND2_X1_147_ (
  .A1({ S17074 }),
  .A2({ S17377 }),
  .ZN({ S17503 })
);
OAI21_X1 #() 
OAI21_X1_1280_ (
  .A({ S16967 }),
  .B1({ S17503 }),
  .B2({ S17005 }),
  .ZN({ S17504 })
);
NAND2_X1 #() 
NAND2_X1_2390_ (
  .A1({ S17502 }),
  .A2({ S17504 }),
  .ZN({ S17505 })
);
NAND2_X1 #() 
NAND2_X1_2391_ (
  .A1({ S17505 }),
  .A2({ S15041 }),
  .ZN({ S17506 })
);
OAI211_X1 #() 
OAI211_X1_868_ (
  .A({ S17506 }),
  .B({ S16966 }),
  .C1({ S17496 }),
  .C2({ S15041 }),
  .ZN({ S17507 })
);
NAND3_X1 #() 
NAND3_X1_2603_ (
  .A1({ S17488 }),
  .A2({ S17507 }),
  .A3({ S17462 }),
  .ZN({ S17508 })
);
NAND2_X1 #() 
NAND2_X1_2392_ (
  .A1({ S17496 }),
  .A2({ S25957[134] }),
  .ZN({ S17509 })
);
NAND3_X1 #() 
NAND3_X1_2604_ (
  .A1({ S17502 }),
  .A2({ S17504 }),
  .A3({ S15041 }),
  .ZN({ S17510 })
);
NAND3_X1 #() 
NAND3_X1_2605_ (
  .A1({ S17509 }),
  .A2({ S16966 }),
  .A3({ S17510 }),
  .ZN({ S17512 })
);
NAND2_X1 #() 
NAND2_X1_2393_ (
  .A1({ S17464 }),
  .A2({ S17463 }),
  .ZN({ S17513 })
);
NAND2_X1 #() 
NAND2_X1_2394_ (
  .A1({ S17513 }),
  .A2({ S25957[133] }),
  .ZN({ S17514 })
);
OAI211_X1 #() 
OAI211_X1_869_ (
  .A({ S17514 }),
  .B({ S25957[134] }),
  .C1({ S17470 }),
  .C2({ S25957[133] }),
  .ZN({ S17515 })
);
NAND2_X1 #() 
NAND2_X1_2395_ (
  .A1({ S17482 }),
  .A2({ S25957[132] }),
  .ZN({ S17516 })
);
OAI211_X1 #() 
OAI211_X1_870_ (
  .A({ S17516 }),
  .B({ S16967 }),
  .C1({ S17484 }),
  .C2({ S25957[132] }),
  .ZN({ S17517 })
);
AND2_X1 #() 
AND2_X1_148_ (
  .A1({ S17479 }),
  .A2({ S17474 }),
  .ZN({ S17518 })
);
OAI211_X1 #() 
OAI211_X1_871_ (
  .A({ S17517 }),
  .B({ S15041 }),
  .C1({ S17518 }),
  .C2({ S16967 }),
  .ZN({ S17519 })
);
NAND3_X1 #() 
NAND3_X1_2606_ (
  .A1({ S17519 }),
  .A2({ S17515 }),
  .A3({ S25957[135] }),
  .ZN({ S17520 })
);
NAND3_X1 #() 
NAND3_X1_2607_ (
  .A1({ S17520 }),
  .A2({ S17512 }),
  .A3({ S25957[238] }),
  .ZN({ S17521 })
);
NAND2_X1 #() 
NAND2_X1_2396_ (
  .A1({ S17508 }),
  .A2({ S17521 }),
  .ZN({ S25957[110] })
);
AOI21_X1 #() 
AOI21_X1_1370_ (
  .A({ S17028 }),
  .B1({ S16997 }),
  .B2({ S25957[129] }),
  .ZN({ S17523 })
);
NAND3_X1 #() 
NAND3_X1_2608_ (
  .A1({ S25957[131] }),
  .A2({ S16987 }),
  .A3({ S17076 }),
  .ZN({ S17524 })
);
NAND3_X1 #() 
NAND3_X1_2609_ (
  .A1({ S17037 }),
  .A2({ S51 }),
  .A3({ S17223 }),
  .ZN({ S17525 })
);
AOI21_X1 #() 
AOI21_X1_1371_ (
  .A({ S25957[132] }),
  .B1({ S17524 }),
  .B2({ S17525 }),
  .ZN({ S17526 })
);
AOI211_X1 #() 
AOI211_X1_29_ (
  .A({ S16967 }),
  .B({ S17526 }),
  .C1({ S17057 }),
  .C2({ S17523 }),
  .ZN({ S17527 })
);
NAND2_X1 #() 
NAND2_X1_2397_ (
  .A1({ S17389 }),
  .A2({ S25957[131] }),
  .ZN({ S17528 })
);
NAND4_X1 #() 
NAND4_X1_315_ (
  .A1({ S17528 }),
  .A2({ S17201 }),
  .A3({ S17048 }),
  .A4({ S17046 }),
  .ZN({ S17529 })
);
NOR2_X1 #() 
NOR2_X1_578_ (
  .A1({ S17126 }),
  .A2({ S17003 }),
  .ZN({ S17530 })
);
OAI21_X1 #() 
OAI21_X1_1281_ (
  .A({ S25957[132] }),
  .B1({ S17530 }),
  .B2({ S17367 }),
  .ZN({ S17531 })
);
AOI21_X1 #() 
AOI21_X1_1372_ (
  .A({ S25957[133] }),
  .B1({ S17529 }),
  .B2({ S17531 }),
  .ZN({ S17533 })
);
OR3_X1 #() 
OR3_X1_12_ (
  .A1({ S17527 }),
  .A2({ S17533 }),
  .A3({ S15041 }),
  .ZN({ S17534 })
);
AOI21_X1 #() 
AOI21_X1_1373_ (
  .A({ S17028 }),
  .B1({ S17054 }),
  .B2({ S17019 }),
  .ZN({ S17535 })
);
AND2_X1 #() 
AND2_X1_149_ (
  .A1({ S17236 }),
  .A2({ S17535 }),
  .ZN({ S17536 })
);
NAND3_X1 #() 
NAND3_X1_2610_ (
  .A1({ S51 }),
  .A2({ S25957[129] }),
  .A3({ S16999 }),
  .ZN({ S17537 })
);
AOI21_X1 #() 
AOI21_X1_1374_ (
  .A({ S17028 }),
  .B1({ S17149 }),
  .B2({ S17537 }),
  .ZN({ S17538 })
);
NOR3_X1 #() 
NOR3_X1_77_ (
  .A1({ S17441 }),
  .A2({ S17047 }),
  .A3({ S25957[132] }),
  .ZN({ S17539 })
);
OAI21_X1 #() 
OAI21_X1_1282_ (
  .A({ S25957[133] }),
  .B1({ S17539 }),
  .B2({ S17538 }),
  .ZN({ S17540 })
);
NOR2_X1 #() 
NOR2_X1_579_ (
  .A1({ S17072 }),
  .A2({ S17073 }),
  .ZN({ S17541 })
);
NAND3_X1 #() 
NAND3_X1_2611_ (
  .A1({ S17124 }),
  .A2({ S17028 }),
  .A3({ S17199 }),
  .ZN({ S17542 })
);
OAI21_X1 #() 
OAI21_X1_1283_ (
  .A({ S16967 }),
  .B1({ S17542 }),
  .B2({ S17541 }),
  .ZN({ S17544 })
);
OAI211_X1 #() 
OAI211_X1_872_ (
  .A({ S17540 }),
  .B({ S15041 }),
  .C1({ S17536 }),
  .C2({ S17544 }),
  .ZN({ S17545 })
);
NAND3_X1 #() 
NAND3_X1_2612_ (
  .A1({ S17534 }),
  .A2({ S25957[135] }),
  .A3({ S17545 }),
  .ZN({ S17546 })
);
NAND2_X1 #() 
NAND2_X1_2398_ (
  .A1({ S17283 }),
  .A2({ S51 }),
  .ZN({ S17547 })
);
NAND3_X1 #() 
NAND3_X1_2613_ (
  .A1({ S17547 }),
  .A2({ S25957[132] }),
  .A3({ S17213 }),
  .ZN({ S17548 })
);
OAI21_X1 #() 
OAI21_X1_1284_ (
  .A({ S16971 }),
  .B1({ S17259 }),
  .B2({ S25957[131] }),
  .ZN({ S17549 })
);
AOI21_X1 #() 
AOI21_X1_1375_ (
  .A({ S25957[134] }),
  .B1({ S17549 }),
  .B2({ S17028 }),
  .ZN({ S17550 })
);
NOR2_X1 #() 
NOR2_X1_580_ (
  .A1({ S17299 }),
  .A2({ S17151 }),
  .ZN({ S17551 })
);
OAI21_X1 #() 
OAI21_X1_1285_ (
  .A({ S25957[132] }),
  .B1({ S17140 }),
  .B2({ S17551 }),
  .ZN({ S17552 })
);
AOI21_X1 #() 
AOI21_X1_1376_ (
  .A({ S25957[132] }),
  .B1({ S17168 }),
  .B2({ S16985 }),
  .ZN({ S17553 })
);
AOI21_X1 #() 
AOI21_X1_1377_ (
  .A({ S15041 }),
  .B1({ S17553 }),
  .B2({ S17189 }),
  .ZN({ S17555 })
);
AOI22_X1 #() 
AOI22_X1_301_ (
  .A1({ S17555 }),
  .A2({ S17552 }),
  .B1({ S17550 }),
  .B2({ S17548 }),
  .ZN({ S17556 })
);
NAND3_X1 #() 
NAND3_X1_2614_ (
  .A1({ S16991 }),
  .A2({ S16997 }),
  .A3({ S17199 }),
  .ZN({ S17557 })
);
NAND2_X1 #() 
NAND2_X1_2399_ (
  .A1({ S17557 }),
  .A2({ S17364 }),
  .ZN({ S17558 })
);
NAND2_X1 #() 
NAND2_X1_2400_ (
  .A1({ S17558 }),
  .A2({ S17028 }),
  .ZN({ S17559 })
);
OAI211_X1 #() 
OAI211_X1_873_ (
  .A({ S17361 }),
  .B({ S25957[132] }),
  .C1({ S25957[131] }),
  .C2({ S16964 }),
  .ZN({ S17560 })
);
AND3_X1 #() 
AND3_X1_103_ (
  .A1({ S17559 }),
  .A2({ S15041 }),
  .A3({ S17560 }),
  .ZN({ S17561 })
);
NAND2_X1 #() 
NAND2_X1_2401_ (
  .A1({ S17112 }),
  .A2({ S51 }),
  .ZN({ S17562 })
);
AOI21_X1 #() 
AOI21_X1_1378_ (
  .A({ S25957[132] }),
  .B1({ S17562 }),
  .B2({ S17377 }),
  .ZN({ S17563 })
);
OAI21_X1 #() 
OAI21_X1_1286_ (
  .A({ S25957[131] }),
  .B1({ S17224 }),
  .B2({ S17070 }),
  .ZN({ S17564 })
);
AOI21_X1 #() 
AOI21_X1_1379_ (
  .A({ S17028 }),
  .B1({ S17130 }),
  .B2({ S17564 }),
  .ZN({ S17566 })
);
NOR3_X1 #() 
NOR3_X1_78_ (
  .A1({ S17563 }),
  .A2({ S17566 }),
  .A3({ S15041 }),
  .ZN({ S17567 })
);
OAI21_X1 #() 
OAI21_X1_1287_ (
  .A({ S25957[133] }),
  .B1({ S17567 }),
  .B2({ S17561 }),
  .ZN({ S17568 })
);
OAI211_X1 #() 
OAI211_X1_874_ (
  .A({ S17568 }),
  .B({ S16966 }),
  .C1({ S25957[133] }),
  .C2({ S17556 }),
  .ZN({ S17569 })
);
NAND2_X1 #() 
NAND2_X1_2402_ (
  .A1({ S17546 }),
  .A2({ S17569 }),
  .ZN({ S17570 })
);
XNOR2_X1 #() 
XNOR2_X1_129_ (
  .A({ S17570 }),
  .B({ S25957[239] }),
  .ZN({ S25957[111] })
);
NAND3_X1 #() 
NAND3_X1_2615_ (
  .A1({ S14673 }),
  .A2({ S25957[264] }),
  .A3({ S14672 }),
  .ZN({ S17571 })
);
NAND3_X1 #() 
NAND3_X1_2616_ (
  .A1({ S14665 }),
  .A2({ S13424 }),
  .A3({ S14669 }),
  .ZN({ S17572 })
);
NAND3_X1 #() 
NAND3_X1_2617_ (
  .A1({ S17571 }),
  .A2({ S17572 }),
  .A3({ S25957[137] }),
  .ZN({ S17573 })
);
INV_X1 #() 
INV_X1_755_ (
  .A({ S17573 }),
  .ZN({ S61 })
);
AND2_X1 #() 
AND2_X1_150_ (
  .A1({ S14741 }),
  .A2({ S14738 }),
  .ZN({ S17575 })
);
NAND3_X1 #() 
NAND3_X1_2618_ (
  .A1({ S14670 }),
  .A2({ S14674 }),
  .A3({ S17575 }),
  .ZN({ S62 })
);
INV_X1 #() 
INV_X1_756_ (
  .A({ S25957[240] }),
  .ZN({ S17576 })
);
NAND2_X1 #() 
NAND2_X1_2403_ (
  .A1({ S14451 }),
  .A2({ S14452 }),
  .ZN({ S17577 })
);
AND2_X1 #() 
AND2_X1_151_ (
  .A1({ S14528 }),
  .A2({ S14524 }),
  .ZN({ S17578 })
);
OAI21_X1 #() 
OAI21_X1_1288_ (
  .A({ S25957[266] }),
  .B1({ S14813 }),
  .B2({ S14816 }),
  .ZN({ S17579 })
);
NAND3_X1 #() 
NAND3_X1_2619_ (
  .A1({ S14819 }),
  .A2({ S14820 }),
  .A3({ S13416 }),
  .ZN({ S17580 })
);
NAND2_X1 #() 
NAND2_X1_2404_ (
  .A1({ S17579 }),
  .A2({ S17580 }),
  .ZN({ S17581 })
);
NAND3_X1 #() 
NAND3_X1_2620_ (
  .A1({ S14670 }),
  .A2({ S14674 }),
  .A3({ S17581 }),
  .ZN({ S17582 })
);
NAND2_X1 #() 
NAND2_X1_2405_ (
  .A1({ S17582 }),
  .A2({ S47 }),
  .ZN({ S17583 })
);
NAND2_X1 #() 
NAND2_X1_2406_ (
  .A1({ S17575 }),
  .A2({ S25957[138] }),
  .ZN({ S17585 })
);
NAND4_X1 #() 
NAND4_X1_316_ (
  .A1({ S14670 }),
  .A2({ S14674 }),
  .A3({ S25957[137] }),
  .A4({ S17581 }),
  .ZN({ S17586 })
);
NAND3_X1 #() 
NAND3_X1_2621_ (
  .A1({ S17571 }),
  .A2({ S17572 }),
  .A3({ S25957[138] }),
  .ZN({ S17587 })
);
NAND4_X1 #() 
NAND4_X1_317_ (
  .A1({ S17586 }),
  .A2({ S17587 }),
  .A3({ S17585 }),
  .A4({ S25957[139] }),
  .ZN({ S17588 })
);
NAND3_X1 #() 
NAND3_X1_2622_ (
  .A1({ S17588 }),
  .A2({ S17578 }),
  .A3({ S17583 }),
  .ZN({ S17589 })
);
NAND3_X1 #() 
NAND3_X1_2623_ (
  .A1({ S14670 }),
  .A2({ S14674 }),
  .A3({ S25957[137] }),
  .ZN({ S17590 })
);
NAND3_X1 #() 
NAND3_X1_2624_ (
  .A1({ S17571 }),
  .A2({ S17572 }),
  .A3({ S17575 }),
  .ZN({ S17591 })
);
NAND3_X1 #() 
NAND3_X1_2625_ (
  .A1({ S17591 }),
  .A2({ S17590 }),
  .A3({ S25957[138] }),
  .ZN({ S17592 })
);
NAND2_X1 #() 
NAND2_X1_2407_ (
  .A1({ S17573 }),
  .A2({ S17581 }),
  .ZN({ S17593 })
);
NAND3_X1 #() 
NAND3_X1_2626_ (
  .A1({ S17592 }),
  .A2({ S17593 }),
  .A3({ S25957[139] }),
  .ZN({ S17594 })
);
NAND4_X1 #() 
NAND4_X1_318_ (
  .A1({ S14818 }),
  .A2({ S14738 }),
  .A3({ S14741 }),
  .A4({ S14821 }),
  .ZN({ S17596 })
);
NAND3_X1 #() 
NAND3_X1_2627_ (
  .A1({ S17596 }),
  .A2({ S14670 }),
  .A3({ S14674 }),
  .ZN({ S17597 })
);
AOI21_X1 #() 
AOI21_X1_1380_ (
  .A({ S17578 }),
  .B1({ S47 }),
  .B2({ S17597 }),
  .ZN({ S17598 })
);
NAND2_X1 #() 
NAND2_X1_2408_ (
  .A1({ S17594 }),
  .A2({ S17598 }),
  .ZN({ S17599 })
);
AND2_X1 #() 
AND2_X1_152_ (
  .A1({ S17599 }),
  .A2({ S17589 }),
  .ZN({ S17600 })
);
INV_X1 #() 
INV_X1_757_ (
  .A({ S62 }),
  .ZN({ S17601 })
);
NAND3_X1 #() 
NAND3_X1_2628_ (
  .A1({ S14670 }),
  .A2({ S14674 }),
  .A3({ S25957[138] }),
  .ZN({ S17602 })
);
NAND3_X1 #() 
NAND3_X1_2629_ (
  .A1({ S17571 }),
  .A2({ S17572 }),
  .A3({ S17581 }),
  .ZN({ S17603 })
);
NAND4_X1 #() 
NAND4_X1_319_ (
  .A1({ S17603 }),
  .A2({ S17602 }),
  .A3({ S17585 }),
  .A4({ S25957[139] }),
  .ZN({ S17604 })
);
NAND2_X1 #() 
NAND2_X1_2409_ (
  .A1({ S17596 }),
  .A2({ S47 }),
  .ZN({ S17605 })
);
OAI211_X1 #() 
OAI211_X1_875_ (
  .A({ S17604 }),
  .B({ S17578 }),
  .C1({ S17601 }),
  .C2({ S17605 }),
  .ZN({ S17607 })
);
NAND2_X1 #() 
NAND2_X1_2410_ (
  .A1({ S17581 }),
  .A2({ S25957[137] }),
  .ZN({ S17608 })
);
AOI21_X1 #() 
AOI21_X1_1381_ (
  .A({ S25957[136] }),
  .B1({ S47 }),
  .B2({ S17608 }),
  .ZN({ S17609 })
);
NAND2_X1 #() 
NAND2_X1_2411_ (
  .A1({ S25957[140] }),
  .A2({ S17585 }),
  .ZN({ S17610 })
);
NOR2_X1 #() 
NOR2_X1_581_ (
  .A1({ S17609 }),
  .A2({ S17610 }),
  .ZN({ S17611 })
);
NOR2_X1 #() 
NOR2_X1_582_ (
  .A1({ S17611 }),
  .A2({ S25957[141] }),
  .ZN({ S17612 })
);
AOI21_X1 #() 
AOI21_X1_1382_ (
  .A({ S14361 }),
  .B1({ S17612 }),
  .B2({ S17607 }),
  .ZN({ S17613 })
);
OAI21_X1 #() 
OAI21_X1_1289_ (
  .A({ S17613 }),
  .B1({ S17600 }),
  .B2({ S17577 }),
  .ZN({ S17614 })
);
AOI21_X1 #() 
AOI21_X1_1383_ (
  .A({ S25957[138] }),
  .B1({ S62 }),
  .B2({ S17573 }),
  .ZN({ S17615 })
);
AOI21_X1 #() 
AOI21_X1_1384_ (
  .A({ S17578 }),
  .B1({ S17615 }),
  .B2({ S25957[139] }),
  .ZN({ S17616 })
);
NAND3_X1 #() 
NAND3_X1_2630_ (
  .A1({ S62 }),
  .A2({ S17573 }),
  .A3({ S25957[138] }),
  .ZN({ S17618 })
);
NAND2_X1 #() 
NAND2_X1_2412_ (
  .A1({ S17618 }),
  .A2({ S17608 }),
  .ZN({ S17619 })
);
NAND2_X1 #() 
NAND2_X1_2413_ (
  .A1({ S17619 }),
  .A2({ S47 }),
  .ZN({ S17620 })
);
NAND2_X1 #() 
NAND2_X1_2414_ (
  .A1({ S17571 }),
  .A2({ S17572 }),
  .ZN({ S17621 })
);
NAND2_X1 #() 
NAND2_X1_2415_ (
  .A1({ S25957[138] }),
  .A2({ S25957[137] }),
  .ZN({ S17622 })
);
OAI211_X1 #() 
OAI211_X1_876_ (
  .A({ S62 }),
  .B({ S25957[139] }),
  .C1({ S17621 }),
  .C2({ S17622 }),
  .ZN({ S17623 })
);
NOR2_X1 #() 
NOR2_X1_583_ (
  .A1({ S17581 }),
  .A2({ S25957[137] }),
  .ZN({ S17624 })
);
AOI21_X1 #() 
AOI21_X1_1385_ (
  .A({ S25957[139] }),
  .B1({ S17621 }),
  .B2({ S17624 }),
  .ZN({ S17625 })
);
NAND4_X1 #() 
NAND4_X1_320_ (
  .A1({ S17571 }),
  .A2({ S17572 }),
  .A3({ S17575 }),
  .A4({ S17581 }),
  .ZN({ S17626 })
);
AOI21_X1 #() 
AOI21_X1_1386_ (
  .A({ S25957[140] }),
  .B1({ S17625 }),
  .B2({ S17626 }),
  .ZN({ S17627 })
);
AOI22_X1 #() 
AOI22_X1_302_ (
  .A1({ S17620 }),
  .A2({ S17616 }),
  .B1({ S17623 }),
  .B2({ S17627 }),
  .ZN({ S17629 })
);
INV_X1 #() 
INV_X1_758_ (
  .A({ S17596 }),
  .ZN({ S17630 })
);
NAND2_X1 #() 
NAND2_X1_2416_ (
  .A1({ S17621 }),
  .A2({ S17630 }),
  .ZN({ S17631 })
);
NAND4_X1 #() 
NAND4_X1_321_ (
  .A1({ S17571 }),
  .A2({ S17572 }),
  .A3({ S17575 }),
  .A4({ S25957[138] }),
  .ZN({ S17632 })
);
NAND3_X1 #() 
NAND3_X1_2631_ (
  .A1({ S17631 }),
  .A2({ S25957[139] }),
  .A3({ S17632 }),
  .ZN({ S17633 })
);
OAI211_X1 #() 
OAI211_X1_877_ (
  .A({ S17573 }),
  .B({ S47 }),
  .C1({ S25957[136] }),
  .C2({ S17585 }),
  .ZN({ S17634 })
);
NAND2_X1 #() 
NAND2_X1_2417_ (
  .A1({ S17633 }),
  .A2({ S17634 }),
  .ZN({ S17635 })
);
NAND2_X1 #() 
NAND2_X1_2418_ (
  .A1({ S17635 }),
  .A2({ S17578 }),
  .ZN({ S17636 })
);
INV_X1 #() 
INV_X1_759_ (
  .A({ S17590 }),
  .ZN({ S17637 })
);
NAND2_X1 #() 
NAND2_X1_2419_ (
  .A1({ S17603 }),
  .A2({ S47 }),
  .ZN({ S17638 })
);
NAND3_X1 #() 
NAND3_X1_2632_ (
  .A1({ S62 }),
  .A2({ S17587 }),
  .A3({ S25957[139] }),
  .ZN({ S17640 })
);
OAI211_X1 #() 
OAI211_X1_878_ (
  .A({ S17640 }),
  .B({ S25957[140] }),
  .C1({ S17637 }),
  .C2({ S17638 }),
  .ZN({ S17641 })
);
NAND3_X1 #() 
NAND3_X1_2633_ (
  .A1({ S17636 }),
  .A2({ S17641 }),
  .A3({ S25957[141] }),
  .ZN({ S17642 })
);
OAI211_X1 #() 
OAI211_X1_879_ (
  .A({ S17642 }),
  .B({ S14361 }),
  .C1({ S17629 }),
  .C2({ S25957[141] }),
  .ZN({ S17643 })
);
NAND3_X1 #() 
NAND3_X1_2634_ (
  .A1({ S17643 }),
  .A2({ S17614 }),
  .A3({ S14271 }),
  .ZN({ S17644 })
);
NAND2_X1 #() 
NAND2_X1_2420_ (
  .A1({ S17621 }),
  .A2({ S17622 }),
  .ZN({ S17645 })
);
NOR2_X1 #() 
NOR2_X1_584_ (
  .A1({ S17645 }),
  .A2({ S47 }),
  .ZN({ S17646 })
);
NAND4_X1 #() 
NAND4_X1_322_ (
  .A1({ S14670 }),
  .A2({ S14674 }),
  .A3({ S25957[137] }),
  .A4({ S25957[138] }),
  .ZN({ S17647 })
);
AOI21_X1 #() 
AOI21_X1_1387_ (
  .A({ S25957[139] }),
  .B1({ S17647 }),
  .B2({ S17603 }),
  .ZN({ S17648 })
);
OAI21_X1 #() 
OAI21_X1_1290_ (
  .A({ S17578 }),
  .B1({ S17646 }),
  .B2({ S17648 }),
  .ZN({ S17649 })
);
NOR2_X1 #() 
NOR2_X1_585_ (
  .A1({ S17581 }),
  .A2({ S47 }),
  .ZN({ S17651 })
);
NAND2_X1 #() 
NAND2_X1_2421_ (
  .A1({ S17651 }),
  .A2({ S25957[137] }),
  .ZN({ S17652 })
);
NAND2_X1 #() 
NAND2_X1_2422_ (
  .A1({ S17652 }),
  .A2({ S25957[140] }),
  .ZN({ S17653 })
);
INV_X1 #() 
INV_X1_760_ (
  .A({ S17653 }),
  .ZN({ S17654 })
);
NAND2_X1 #() 
NAND2_X1_2423_ (
  .A1({ S25957[136] }),
  .A2({ S17596 }),
  .ZN({ S17655 })
);
NAND2_X1 #() 
NAND2_X1_2424_ (
  .A1({ S17621 }),
  .A2({ S17608 }),
  .ZN({ S17656 })
);
NAND3_X1 #() 
NAND3_X1_2635_ (
  .A1({ S17655 }),
  .A2({ S17656 }),
  .A3({ S47 }),
  .ZN({ S17657 })
);
NAND2_X1 #() 
NAND2_X1_2425_ (
  .A1({ S17654 }),
  .A2({ S17657 }),
  .ZN({ S17658 })
);
NAND3_X1 #() 
NAND3_X1_2636_ (
  .A1({ S17658 }),
  .A2({ S17649 }),
  .A3({ S17577 }),
  .ZN({ S17659 })
);
AOI21_X1 #() 
AOI21_X1_1388_ (
  .A({ S47 }),
  .B1({ S17621 }),
  .B2({ S17624 }),
  .ZN({ S17660 })
);
AOI21_X1 #() 
AOI21_X1_1389_ (
  .A({ S25957[139] }),
  .B1({ S17626 }),
  .B2({ S17647 }),
  .ZN({ S17662 })
);
OAI21_X1 #() 
OAI21_X1_1291_ (
  .A({ S25957[140] }),
  .B1({ S17662 }),
  .B2({ S17660 }),
  .ZN({ S17663 })
);
NAND3_X1 #() 
NAND3_X1_2637_ (
  .A1({ S17590 }),
  .A2({ S17582 }),
  .A3({ S17608 }),
  .ZN({ S17664 })
);
AOI21_X1 #() 
AOI21_X1_1390_ (
  .A({ S17625 }),
  .B1({ S17664 }),
  .B2({ S25957[139] }),
  .ZN({ S17665 })
);
OAI211_X1 #() 
OAI211_X1_880_ (
  .A({ S17663 }),
  .B({ S25957[141] }),
  .C1({ S25957[140] }),
  .C2({ S17665 }),
  .ZN({ S17666 })
);
AND2_X1 #() 
AND2_X1_153_ (
  .A1({ S17666 }),
  .A2({ S17659 }),
  .ZN({ S17667 })
);
AOI22_X1 #() 
AOI22_X1_303_ (
  .A1({ S14674 }),
  .A2({ S14670 }),
  .B1({ S17575 }),
  .B2({ S17581 }),
  .ZN({ S17668 })
);
AOI22_X1 #() 
AOI22_X1_304_ (
  .A1({ S17571 }),
  .A2({ S17572 }),
  .B1({ S17581 }),
  .B2({ S25957[137] }),
  .ZN({ S17669 })
);
AOI21_X1 #() 
AOI21_X1_1391_ (
  .A({ S25957[139] }),
  .B1({ S25957[137] }),
  .B2({ S25957[138] }),
  .ZN({ S17670 })
);
OAI21_X1 #() 
OAI21_X1_1292_ (
  .A({ S17670 }),
  .B1({ S17668 }),
  .B2({ S17669 }),
  .ZN({ S17671 })
);
NAND3_X1 #() 
NAND3_X1_2638_ (
  .A1({ S17597 }),
  .A2({ S17603 }),
  .A3({ S47 }),
  .ZN({ S17673 })
);
NAND2_X1 #() 
NAND2_X1_2426_ (
  .A1({ S17590 }),
  .A2({ S17651 }),
  .ZN({ S17674 })
);
NAND3_X1 #() 
NAND3_X1_2639_ (
  .A1({ S25957[138] }),
  .A2({ S47 }),
  .A3({ S25957[137] }),
  .ZN({ S17675 })
);
NAND3_X1 #() 
NAND3_X1_2640_ (
  .A1({ S17673 }),
  .A2({ S17674 }),
  .A3({ S17675 }),
  .ZN({ S17676 })
);
NAND3_X1 #() 
NAND3_X1_2641_ (
  .A1({ S17626 }),
  .A2({ S25957[139] }),
  .A3({ S17602 }),
  .ZN({ S17677 })
);
AND2_X1 #() 
AND2_X1_154_ (
  .A1({ S17677 }),
  .A2({ S17578 }),
  .ZN({ S17678 })
);
AOI22_X1 #() 
AOI22_X1_305_ (
  .A1({ S17678 }),
  .A2({ S17671 }),
  .B1({ S17676 }),
  .B2({ S25957[140] }),
  .ZN({ S17679 })
);
INV_X1 #() 
INV_X1_761_ (
  .A({ S17586 }),
  .ZN({ S17680 })
);
NAND3_X1 #() 
NAND3_X1_2642_ (
  .A1({ S17591 }),
  .A2({ S17590 }),
  .A3({ S17651 }),
  .ZN({ S17681 })
);
NAND2_X1 #() 
NAND2_X1_2427_ (
  .A1({ S17632 }),
  .A2({ S47 }),
  .ZN({ S17682 })
);
OAI211_X1 #() 
OAI211_X1_881_ (
  .A({ S17681 }),
  .B({ S25957[140] }),
  .C1({ S17682 }),
  .C2({ S17680 }),
  .ZN({ S17684 })
);
NAND2_X1 #() 
NAND2_X1_2428_ (
  .A1({ S17586 }),
  .A2({ S47 }),
  .ZN({ S17685 })
);
NAND3_X1 #() 
NAND3_X1_2643_ (
  .A1({ S17604 }),
  .A2({ S17578 }),
  .A3({ S17685 }),
  .ZN({ S17686 })
);
NAND3_X1 #() 
NAND3_X1_2644_ (
  .A1({ S17684 }),
  .A2({ S17686 }),
  .A3({ S17577 }),
  .ZN({ S17687 })
);
OAI211_X1 #() 
OAI211_X1_882_ (
  .A({ S25957[142] }),
  .B({ S17687 }),
  .C1({ S17679 }),
  .C2({ S17577 }),
  .ZN({ S17688 })
);
OAI211_X1 #() 
OAI211_X1_883_ (
  .A({ S25957[143] }),
  .B({ S17688 }),
  .C1({ S17667 }),
  .C2({ S25957[142] }),
  .ZN({ S17689 })
);
NAND3_X1 #() 
NAND3_X1_2645_ (
  .A1({ S17689 }),
  .A2({ S17644 }),
  .A3({ S17576 }),
  .ZN({ S17690 })
);
AOI21_X1 #() 
AOI21_X1_1392_ (
  .A({ S17577 }),
  .B1({ S17599 }),
  .B2({ S17589 }),
  .ZN({ S17691 })
);
OR2_X1 #() 
OR2_X1_34_ (
  .A1({ S17609 }),
  .A2({ S17610 }),
  .ZN({ S17692 })
);
AND3_X1 #() 
AND3_X1_104_ (
  .A1({ S17607 }),
  .A2({ S17692 }),
  .A3({ S17577 }),
  .ZN({ S17693 })
);
OAI21_X1 #() 
OAI21_X1_1293_ (
  .A({ S25957[142] }),
  .B1({ S17691 }),
  .B2({ S17693 }),
  .ZN({ S17695 })
);
NAND2_X1 #() 
NAND2_X1_2429_ (
  .A1({ S17603 }),
  .A2({ S17596 }),
  .ZN({ S17696 })
);
NAND2_X1 #() 
NAND2_X1_2430_ (
  .A1({ S17696 }),
  .A2({ S17591 }),
  .ZN({ S17697 })
);
OAI21_X1 #() 
OAI21_X1_1294_ (
  .A({ S25957[140] }),
  .B1({ S17697 }),
  .B2({ S47 }),
  .ZN({ S17698 })
);
AOI21_X1 #() 
AOI21_X1_1393_ (
  .A({ S25957[139] }),
  .B1({ S17618 }),
  .B2({ S17608 }),
  .ZN({ S17699 })
);
NAND2_X1 #() 
NAND2_X1_2431_ (
  .A1({ S17625 }),
  .A2({ S17626 }),
  .ZN({ S17700 })
);
NAND3_X1 #() 
NAND3_X1_2646_ (
  .A1({ S17700 }),
  .A2({ S17578 }),
  .A3({ S17623 }),
  .ZN({ S17701 })
);
OAI211_X1 #() 
OAI211_X1_884_ (
  .A({ S17701 }),
  .B({ S17577 }),
  .C1({ S17698 }),
  .C2({ S17699 }),
  .ZN({ S17702 })
);
OAI21_X1 #() 
OAI21_X1_1295_ (
  .A({ S17640 }),
  .B1({ S17637 }),
  .B2({ S17638 }),
  .ZN({ S17703 })
);
NAND2_X1 #() 
NAND2_X1_2432_ (
  .A1({ S17703 }),
  .A2({ S25957[140] }),
  .ZN({ S17704 })
);
OAI211_X1 #() 
OAI211_X1_885_ (
  .A({ S17704 }),
  .B({ S25957[141] }),
  .C1({ S25957[140] }),
  .C2({ S17635 }),
  .ZN({ S17706 })
);
NAND3_X1 #() 
NAND3_X1_2647_ (
  .A1({ S17706 }),
  .A2({ S17702 }),
  .A3({ S14361 }),
  .ZN({ S17707 })
);
AOI21_X1 #() 
AOI21_X1_1394_ (
  .A({ S25957[143] }),
  .B1({ S17695 }),
  .B2({ S17707 }),
  .ZN({ S17708 })
);
NAND2_X1 #() 
NAND2_X1_2433_ (
  .A1({ S17676 }),
  .A2({ S25957[140] }),
  .ZN({ S17709 })
);
NAND3_X1 #() 
NAND3_X1_2648_ (
  .A1({ S17671 }),
  .A2({ S17578 }),
  .A3({ S17677 }),
  .ZN({ S17710 })
);
AOI21_X1 #() 
AOI21_X1_1395_ (
  .A({ S17577 }),
  .B1({ S17709 }),
  .B2({ S17710 }),
  .ZN({ S17711 })
);
AND3_X1 #() 
AND3_X1_105_ (
  .A1({ S17684 }),
  .A2({ S17686 }),
  .A3({ S17577 }),
  .ZN({ S17712 })
);
OAI21_X1 #() 
OAI21_X1_1296_ (
  .A({ S25957[142] }),
  .B1({ S17711 }),
  .B2({ S17712 }),
  .ZN({ S17713 })
);
NAND3_X1 #() 
NAND3_X1_2649_ (
  .A1({ S17666 }),
  .A2({ S17659 }),
  .A3({ S14361 }),
  .ZN({ S17714 })
);
AOI21_X1 #() 
AOI21_X1_1396_ (
  .A({ S14271 }),
  .B1({ S17713 }),
  .B2({ S17714 }),
  .ZN({ S17715 })
);
OAI21_X1 #() 
OAI21_X1_1297_ (
  .A({ S25957[240] }),
  .B1({ S17708 }),
  .B2({ S17715 }),
  .ZN({ S17717 })
);
NAND2_X1 #() 
NAND2_X1_2434_ (
  .A1({ S17717 }),
  .A2({ S17690 }),
  .ZN({ S25957[112] })
);
INV_X1 #() 
INV_X1_762_ (
  .A({ S25957[241] }),
  .ZN({ S17718 })
);
NOR2_X1 #() 
NOR2_X1_586_ (
  .A1({ S25957[136] }),
  .A2({ S25957[139] }),
  .ZN({ S17719 })
);
AOI21_X1 #() 
AOI21_X1_1397_ (
  .A({ S17578 }),
  .B1({ S17719 }),
  .B2({ S17585 }),
  .ZN({ S17720 })
);
XNOR2_X1 #() 
XNOR2_X1_130_ (
  .A({ S25957[136] }),
  .B({ S17622 }),
  .ZN({ S17721 })
);
NAND2_X1 #() 
NAND2_X1_2435_ (
  .A1({ S17721 }),
  .A2({ S25957[139] }),
  .ZN({ S17722 })
);
AND2_X1 #() 
AND2_X1_155_ (
  .A1({ S17722 }),
  .A2({ S17720 }),
  .ZN({ S17723 })
);
NOR2_X1 #() 
NOR2_X1_587_ (
  .A1({ S17630 }),
  .A2({ S47 }),
  .ZN({ S17724 })
);
NAND2_X1 #() 
NAND2_X1_2436_ (
  .A1({ S17724 }),
  .A2({ S17603 }),
  .ZN({ S17725 })
);
NAND2_X1 #() 
NAND2_X1_2437_ (
  .A1({ S17608 }),
  .A2({ S47 }),
  .ZN({ S17727 })
);
INV_X1 #() 
INV_X1_763_ (
  .A({ S17727 }),
  .ZN({ S17728 })
);
NAND2_X1 #() 
NAND2_X1_2438_ (
  .A1({ S17728 }),
  .A2({ S17591 }),
  .ZN({ S17729 })
);
AOI21_X1 #() 
AOI21_X1_1398_ (
  .A({ S25957[140] }),
  .B1({ S17729 }),
  .B2({ S17725 }),
  .ZN({ S17730 })
);
NOR3_X1 #() 
NOR3_X1_79_ (
  .A1({ S17723 }),
  .A2({ S17730 }),
  .A3({ S25957[142] }),
  .ZN({ S17731 })
);
NAND2_X1 #() 
NAND2_X1_2439_ (
  .A1({ S17647 }),
  .A2({ S47 }),
  .ZN({ S17732 })
);
AOI21_X1 #() 
AOI21_X1_1399_ (
  .A({ S25957[140] }),
  .B1({ S17594 }),
  .B2({ S17732 }),
  .ZN({ S17733 })
);
NAND2_X1 #() 
NAND2_X1_2440_ (
  .A1({ S17573 }),
  .A2({ S25957[138] }),
  .ZN({ S17734 })
);
INV_X1 #() 
INV_X1_764_ (
  .A({ S17734 }),
  .ZN({ S17735 })
);
NAND2_X1 #() 
NAND2_X1_2441_ (
  .A1({ S17735 }),
  .A2({ S47 }),
  .ZN({ S17736 })
);
NOR2_X1 #() 
NOR2_X1_588_ (
  .A1({ S17573 }),
  .A2({ S47 }),
  .ZN({ S17738 })
);
NOR2_X1 #() 
NOR2_X1_589_ (
  .A1({ S17653 }),
  .A2({ S17738 }),
  .ZN({ S17739 })
);
AND2_X1 #() 
AND2_X1_156_ (
  .A1({ S17739 }),
  .A2({ S17736 }),
  .ZN({ S17740 })
);
NOR3_X1 #() 
NOR3_X1_80_ (
  .A1({ S17740 }),
  .A2({ S17733 }),
  .A3({ S14361 }),
  .ZN({ S17741 })
);
OAI21_X1 #() 
OAI21_X1_1298_ (
  .A({ S25957[141] }),
  .B1({ S17731 }),
  .B2({ S17741 }),
  .ZN({ S17742 })
);
AOI21_X1 #() 
AOI21_X1_1400_ (
  .A({ S47 }),
  .B1({ S17697 }),
  .B2({ S17734 }),
  .ZN({ S17743 })
);
NAND2_X1 #() 
NAND2_X1_2442_ (
  .A1({ S17586 }),
  .A2({ S17585 }),
  .ZN({ S17744 })
);
NAND2_X1 #() 
NAND2_X1_2443_ (
  .A1({ S17587 }),
  .A2({ S47 }),
  .ZN({ S17745 })
);
OAI21_X1 #() 
OAI21_X1_1299_ (
  .A({ S17578 }),
  .B1({ S17744 }),
  .B2({ S17745 }),
  .ZN({ S17746 })
);
OAI221_X1 #() 
OAI221_X1_59_ (
  .A({ S25957[140] }),
  .B1({ S17608 }),
  .B2({ S47 }),
  .C1({ S17685 }),
  .C2({ S17624 }),
  .ZN({ S17747 })
);
OAI21_X1 #() 
OAI21_X1_1300_ (
  .A({ S17747 }),
  .B1({ S17743 }),
  .B2({ S17746 }),
  .ZN({ S17749 })
);
INV_X1 #() 
INV_X1_765_ (
  .A({ S17618 }),
  .ZN({ S17750 })
);
NAND2_X1 #() 
NAND2_X1_2444_ (
  .A1({ S25957[136] }),
  .A2({ S47 }),
  .ZN({ S17751 })
);
NAND2_X1 #() 
NAND2_X1_2445_ (
  .A1({ S17751 }),
  .A2({ S25957[140] }),
  .ZN({ S17752 })
);
INV_X1 #() 
INV_X1_766_ (
  .A({ S17752 }),
  .ZN({ S17753 })
);
OAI211_X1 #() 
OAI211_X1_886_ (
  .A({ S17753 }),
  .B({ S17675 }),
  .C1({ S17750 }),
  .C2({ S17725 }),
  .ZN({ S17754 })
);
NAND2_X1 #() 
NAND2_X1_2446_ (
  .A1({ S17655 }),
  .A2({ S47 }),
  .ZN({ S17755 })
);
AOI211_X1 #() 
AOI211_X1_30_ (
  .A({ S25957[140] }),
  .B({ S17755 }),
  .C1({ S17621 }),
  .C2({ S17630 }),
  .ZN({ S17756 })
);
NAND2_X1 #() 
NAND2_X1_2447_ (
  .A1({ S17602 }),
  .A2({ S25957[139] }),
  .ZN({ S17757 })
);
NOR3_X1 #() 
NOR3_X1_81_ (
  .A1({ S17757 }),
  .A2({ S61 }),
  .A3({ S25957[140] }),
  .ZN({ S17758 })
);
NOR3_X1 #() 
NOR3_X1_82_ (
  .A1({ S17756 }),
  .A2({ S17758 }),
  .A3({ S14361 }),
  .ZN({ S17760 })
);
AOI22_X1 #() 
AOI22_X1_306_ (
  .A1({ S17760 }),
  .A2({ S17754 }),
  .B1({ S17749 }),
  .B2({ S14361 }),
  .ZN({ S17761 })
);
OAI211_X1 #() 
OAI211_X1_887_ (
  .A({ S17742 }),
  .B({ S25957[143] }),
  .C1({ S17761 }),
  .C2({ S25957[141] }),
  .ZN({ S17762 })
);
NAND2_X1 #() 
NAND2_X1_2448_ (
  .A1({ S17590 }),
  .A2({ S17622 }),
  .ZN({ S17763 })
);
NAND2_X1 #() 
NAND2_X1_2449_ (
  .A1({ S17763 }),
  .A2({ S17602 }),
  .ZN({ S17764 })
);
OAI221_X1 #() 
OAI221_X1_60_ (
  .A({ S25957[141] }),
  .B1({ S25957[136] }),
  .B2({ S17727 }),
  .C1({ S17764 }),
  .C2({ S47 }),
  .ZN({ S17765 })
);
NOR2_X1 #() 
NOR2_X1_590_ (
  .A1({ S47 }),
  .A2({ S25957[137] }),
  .ZN({ S17766 })
);
NOR2_X1 #() 
NOR2_X1_591_ (
  .A1({ S17587 }),
  .A2({ S47 }),
  .ZN({ S17767 })
);
NOR2_X1 #() 
NOR2_X1_592_ (
  .A1({ S17767 }),
  .A2({ S17766 }),
  .ZN({ S17768 })
);
NAND2_X1 #() 
NAND2_X1_2450_ (
  .A1({ S17587 }),
  .A2({ S17608 }),
  .ZN({ S17769 })
);
NAND2_X1 #() 
NAND2_X1_2451_ (
  .A1({ S17769 }),
  .A2({ S47 }),
  .ZN({ S17771 })
);
NAND3_X1 #() 
NAND3_X1_2650_ (
  .A1({ S17768 }),
  .A2({ S17577 }),
  .A3({ S17771 }),
  .ZN({ S17772 })
);
AND2_X1 #() 
AND2_X1_157_ (
  .A1({ S17765 }),
  .A2({ S17772 }),
  .ZN({ S17773 })
);
NAND2_X1 #() 
NAND2_X1_2452_ (
  .A1({ S17773 }),
  .A2({ S25957[140] }),
  .ZN({ S17774 })
);
NAND2_X1 #() 
NAND2_X1_2453_ (
  .A1({ S17622 }),
  .A2({ S17596 }),
  .ZN({ S17775 })
);
AOI21_X1 #() 
AOI21_X1_1401_ (
  .A({ S25957[139] }),
  .B1({ S17775 }),
  .B2({ S25957[136] }),
  .ZN({ S17776 })
);
NOR2_X1 #() 
NOR2_X1_593_ (
  .A1({ S17776 }),
  .A2({ S25957[140] }),
  .ZN({ S17777 })
);
INV_X1 #() 
INV_X1_767_ (
  .A({ S17724 }),
  .ZN({ S17778 })
);
NOR2_X1 #() 
NOR2_X1_594_ (
  .A1({ S25957[141] }),
  .A2({ S17778 }),
  .ZN({ S17779 })
);
INV_X1 #() 
INV_X1_768_ (
  .A({ S17779 }),
  .ZN({ S17780 })
);
AOI21_X1 #() 
AOI21_X1_1402_ (
  .A({ S25957[142] }),
  .B1({ S17780 }),
  .B2({ S17777 }),
  .ZN({ S17782 })
);
NAND2_X1 #() 
NAND2_X1_2454_ (
  .A1({ S17774 }),
  .A2({ S17782 }),
  .ZN({ S17783 })
);
NAND2_X1 #() 
NAND2_X1_2455_ (
  .A1({ S17591 }),
  .A2({ S25957[139] }),
  .ZN({ S17784 })
);
INV_X1 #() 
INV_X1_769_ (
  .A({ S17784 }),
  .ZN({ S17785 })
);
NAND2_X1 #() 
NAND2_X1_2456_ (
  .A1({ S62 }),
  .A2({ S17603 }),
  .ZN({ S17786 })
);
NAND2_X1 #() 
NAND2_X1_2457_ (
  .A1({ S17785 }),
  .A2({ S17786 }),
  .ZN({ S17787 })
);
OAI211_X1 #() 
OAI211_X1_888_ (
  .A({ S17603 }),
  .B({ S47 }),
  .C1({ S25957[136] }),
  .C2({ S17585 }),
  .ZN({ S17788 })
);
AOI21_X1 #() 
AOI21_X1_1403_ (
  .A({ S17578 }),
  .B1({ S17787 }),
  .B2({ S17788 }),
  .ZN({ S17789 })
);
AOI21_X1 #() 
AOI21_X1_1404_ (
  .A({ S25957[140] }),
  .B1({ S17768 }),
  .B2({ S17673 }),
  .ZN({ S17790 })
);
OAI21_X1 #() 
OAI21_X1_1301_ (
  .A({ S25957[141] }),
  .B1({ S17789 }),
  .B2({ S17790 }),
  .ZN({ S17791 })
);
NAND3_X1 #() 
NAND3_X1_2651_ (
  .A1({ S17734 }),
  .A2({ S47 }),
  .A3({ S17603 }),
  .ZN({ S17793 })
);
NAND3_X1 #() 
NAND3_X1_2652_ (
  .A1({ S17793 }),
  .A2({ S17578 }),
  .A3({ S17681 }),
  .ZN({ S17794 })
);
NOR2_X1 #() 
NOR2_X1_595_ (
  .A1({ S17621 }),
  .A2({ S17622 }),
  .ZN({ S17795 })
);
NAND2_X1 #() 
NAND2_X1_2458_ (
  .A1({ S17631 }),
  .A2({ S47 }),
  .ZN({ S17796 })
);
OAI211_X1 #() 
OAI211_X1_889_ (
  .A({ S17594 }),
  .B({ S25957[140] }),
  .C1({ S17795 }),
  .C2({ S17796 }),
  .ZN({ S17797 })
);
NAND3_X1 #() 
NAND3_X1_2653_ (
  .A1({ S17797 }),
  .A2({ S17577 }),
  .A3({ S17794 }),
  .ZN({ S17798 })
);
NAND3_X1 #() 
NAND3_X1_2654_ (
  .A1({ S17791 }),
  .A2({ S17798 }),
  .A3({ S25957[142] }),
  .ZN({ S17799 })
);
NAND3_X1 #() 
NAND3_X1_2655_ (
  .A1({ S17783 }),
  .A2({ S14271 }),
  .A3({ S17799 }),
  .ZN({ S17800 })
);
NAND3_X1 #() 
NAND3_X1_2656_ (
  .A1({ S17762 }),
  .A2({ S17800 }),
  .A3({ S17718 }),
  .ZN({ S17801 })
);
OAI21_X1 #() 
OAI21_X1_1302_ (
  .A({ S25957[141] }),
  .B1({ S17723 }),
  .B2({ S17730 }),
  .ZN({ S17802 })
);
OAI211_X1 #() 
OAI211_X1_890_ (
  .A({ S17747 }),
  .B({ S17577 }),
  .C1({ S17743 }),
  .C2({ S17746 }),
  .ZN({ S17804 })
);
AND2_X1 #() 
AND2_X1_158_ (
  .A1({ S17802 }),
  .A2({ S17804 }),
  .ZN({ S17805 })
);
NOR2_X1 #() 
NOR2_X1_596_ (
  .A1({ S17757 }),
  .A2({ S61 }),
  .ZN({ S17806 })
);
AOI21_X1 #() 
AOI21_X1_1405_ (
  .A({ S25957[139] }),
  .B1({ S17626 }),
  .B2({ S17597 }),
  .ZN({ S17807 })
);
OAI21_X1 #() 
OAI21_X1_1303_ (
  .A({ S17578 }),
  .B1({ S17806 }),
  .B2({ S17807 }),
  .ZN({ S17808 })
);
NAND3_X1 #() 
NAND3_X1_2657_ (
  .A1({ S17754 }),
  .A2({ S17577 }),
  .A3({ S17808 }),
  .ZN({ S17809 })
);
OR3_X1 #() 
OR3_X1_13_ (
  .A1({ S17740 }),
  .A2({ S17733 }),
  .A3({ S17577 }),
  .ZN({ S17810 })
);
NAND3_X1 #() 
NAND3_X1_2658_ (
  .A1({ S17810 }),
  .A2({ S25957[142] }),
  .A3({ S17809 }),
  .ZN({ S17811 })
);
OAI211_X1 #() 
OAI211_X1_891_ (
  .A({ S17811 }),
  .B({ S25957[143] }),
  .C1({ S17805 }),
  .C2({ S25957[142] }),
  .ZN({ S17812 })
);
AND2_X1 #() 
AND2_X1_159_ (
  .A1({ S17791 }),
  .A2({ S17798 }),
  .ZN({ S17813 })
);
OAI21_X1 #() 
OAI21_X1_1304_ (
  .A({ S17578 }),
  .B1({ S17779 }),
  .B2({ S17776 }),
  .ZN({ S17815 })
);
OAI211_X1 #() 
OAI211_X1_892_ (
  .A({ S14361 }),
  .B({ S17815 }),
  .C1({ S17773 }),
  .C2({ S17578 }),
  .ZN({ S17816 })
);
OAI211_X1 #() 
OAI211_X1_893_ (
  .A({ S17816 }),
  .B({ S14271 }),
  .C1({ S14361 }),
  .C2({ S17813 }),
  .ZN({ S17817 })
);
NAND3_X1 #() 
NAND3_X1_2659_ (
  .A1({ S17817 }),
  .A2({ S17812 }),
  .A3({ S25957[241] }),
  .ZN({ S17818 })
);
NAND2_X1 #() 
NAND2_X1_2459_ (
  .A1({ S17818 }),
  .A2({ S17801 }),
  .ZN({ S25957[113] })
);
NAND3_X1 #() 
NAND3_X1_2660_ (
  .A1({ S17632 }),
  .A2({ S25957[139] }),
  .A3({ S17590 }),
  .ZN({ S17819 })
);
NAND2_X1 #() 
NAND2_X1_2460_ (
  .A1({ S17670 }),
  .A2({ S17587 }),
  .ZN({ S17820 })
);
AOI21_X1 #() 
AOI21_X1_1406_ (
  .A({ S25957[140] }),
  .B1({ S17819 }),
  .B2({ S17820 }),
  .ZN({ S17821 })
);
NAND2_X1 #() 
NAND2_X1_2461_ (
  .A1({ S17585 }),
  .A2({ S17608 }),
  .ZN({ S17822 })
);
NOR2_X1 #() 
NOR2_X1_597_ (
  .A1({ S17751 }),
  .A2({ S17822 }),
  .ZN({ S17823 })
);
AOI21_X1 #() 
AOI21_X1_1407_ (
  .A({ S17823 }),
  .B1({ S17724 }),
  .B2({ S25957[136] }),
  .ZN({ S17825 })
);
OAI21_X1 #() 
OAI21_X1_1305_ (
  .A({ S25957[141] }),
  .B1({ S17825 }),
  .B2({ S17578 }),
  .ZN({ S17826 })
);
AOI21_X1 #() 
AOI21_X1_1408_ (
  .A({ S17578 }),
  .B1({ S17763 }),
  .B2({ S25957[139] }),
  .ZN({ S17827 })
);
NAND2_X1 #() 
NAND2_X1_2462_ (
  .A1({ S17827 }),
  .A2({ S17727 }),
  .ZN({ S17828 })
);
NAND2_X1 #() 
NAND2_X1_2463_ (
  .A1({ S17680 }),
  .A2({ S47 }),
  .ZN({ S17829 })
);
NAND3_X1 #() 
NAND3_X1_2661_ (
  .A1({ S17829 }),
  .A2({ S17578 }),
  .A3({ S17652 }),
  .ZN({ S17830 })
);
AND2_X1 #() 
AND2_X1_160_ (
  .A1({ S17828 }),
  .A2({ S17830 }),
  .ZN({ S17831 })
);
OAI22_X1 #() 
OAI22_X1_54_ (
  .A1({ S17826 }),
  .A2({ S17821 }),
  .B1({ S17831 }),
  .B2({ S25957[141] }),
  .ZN({ S17832 })
);
NAND2_X1 #() 
NAND2_X1_2464_ (
  .A1({ S17832 }),
  .A2({ S14361 }),
  .ZN({ S17833 })
);
NAND2_X1 #() 
NAND2_X1_2465_ (
  .A1({ S17632 }),
  .A2({ S25957[139] }),
  .ZN({ S17834 })
);
NOR2_X1 #() 
NOR2_X1_598_ (
  .A1({ S17624 }),
  .A2({ S25957[139] }),
  .ZN({ S17836 })
);
AOI21_X1 #() 
AOI21_X1_1409_ (
  .A({ S17578 }),
  .B1({ S17836 }),
  .B2({ S62 }),
  .ZN({ S17837 })
);
OAI21_X1 #() 
OAI21_X1_1306_ (
  .A({ S17837 }),
  .B1({ S17615 }),
  .B2({ S17834 }),
  .ZN({ S17838 })
);
AOI22_X1 #() 
AOI22_X1_307_ (
  .A1({ S17785 }),
  .A2({ S17608 }),
  .B1({ S17630 }),
  .B2({ S47 }),
  .ZN({ S17839 })
);
OAI211_X1 #() 
OAI211_X1_894_ (
  .A({ S17838 }),
  .B({ S17577 }),
  .C1({ S25957[140] }),
  .C2({ S17839 }),
  .ZN({ S17840 })
);
NAND2_X1 #() 
NAND2_X1_2466_ (
  .A1({ S17724 }),
  .A2({ S17602 }),
  .ZN({ S17841 })
);
NAND3_X1 #() 
NAND3_X1_2662_ (
  .A1({ S17671 }),
  .A2({ S25957[140] }),
  .A3({ S17841 }),
  .ZN({ S17842 })
);
NAND2_X1 #() 
NAND2_X1_2467_ (
  .A1({ S17647 }),
  .A2({ S25957[139] }),
  .ZN({ S17843 })
);
AND2_X1 #() 
AND2_X1_161_ (
  .A1({ S17578 }),
  .A2({ S17675 }),
  .ZN({ S17844 })
);
OAI21_X1 #() 
OAI21_X1_1307_ (
  .A({ S17844 }),
  .B1({ S17615 }),
  .B2({ S17843 }),
  .ZN({ S17845 })
);
NAND3_X1 #() 
NAND3_X1_2663_ (
  .A1({ S17845 }),
  .A2({ S17842 }),
  .A3({ S25957[141] }),
  .ZN({ S17847 })
);
NAND2_X1 #() 
NAND2_X1_2468_ (
  .A1({ S17840 }),
  .A2({ S17847 }),
  .ZN({ S17848 })
);
NAND2_X1 #() 
NAND2_X1_2469_ (
  .A1({ S17848 }),
  .A2({ S25957[142] }),
  .ZN({ S17849 })
);
NAND3_X1 #() 
NAND3_X1_2664_ (
  .A1({ S17833 }),
  .A2({ S25957[143] }),
  .A3({ S17849 }),
  .ZN({ S17850 })
);
INV_X1 #() 
INV_X1_770_ (
  .A({ S17597 }),
  .ZN({ S17851 })
);
OAI21_X1 #() 
OAI21_X1_1308_ (
  .A({ S25957[140] }),
  .B1({ S17851 }),
  .B2({ S47 }),
  .ZN({ S17852 })
);
INV_X1 #() 
INV_X1_771_ (
  .A({ S17603 }),
  .ZN({ S17853 })
);
NAND2_X1 #() 
NAND2_X1_2470_ (
  .A1({ S17853 }),
  .A2({ S25957[140] }),
  .ZN({ S17854 })
);
AOI22_X1 #() 
AOI22_X1_308_ (
  .A1({ S17852 }),
  .A2({ S17854 }),
  .B1({ S17728 }),
  .B2({ S17592 }),
  .ZN({ S17855 })
);
NOR2_X1 #() 
NOR2_X1_599_ (
  .A1({ S17621 }),
  .A2({ S17608 }),
  .ZN({ S17856 })
);
OAI21_X1 #() 
OAI21_X1_1309_ (
  .A({ S25957[139] }),
  .B1({ S17735 }),
  .B2({ S17856 }),
  .ZN({ S17858 })
);
AOI21_X1 #() 
AOI21_X1_1410_ (
  .A({ S25957[140] }),
  .B1({ S17858 }),
  .B2({ S17829 }),
  .ZN({ S17859 })
);
OAI21_X1 #() 
OAI21_X1_1310_ (
  .A({ S25957[141] }),
  .B1({ S17859 }),
  .B2({ S17855 }),
  .ZN({ S17860 })
);
NAND2_X1 #() 
NAND2_X1_2471_ (
  .A1({ S17588 }),
  .A2({ S17578 }),
  .ZN({ S17861 })
);
INV_X1 #() 
INV_X1_772_ (
  .A({ S17671 }),
  .ZN({ S17862 })
);
NAND2_X1 #() 
NAND2_X1_2472_ (
  .A1({ S17590 }),
  .A2({ S25957[138] }),
  .ZN({ S17863 })
);
INV_X1 #() 
INV_X1_773_ (
  .A({ S17863 }),
  .ZN({ S17864 })
);
INV_X1 #() 
INV_X1_774_ (
  .A({ S17593 }),
  .ZN({ S17865 })
);
OAI21_X1 #() 
OAI21_X1_1311_ (
  .A({ S47 }),
  .B1({ S17865 }),
  .B2({ S17864 }),
  .ZN({ S17866 })
);
NAND2_X1 #() 
NAND2_X1_2473_ (
  .A1({ S17866 }),
  .A2({ S17827 }),
  .ZN({ S17867 })
);
OAI211_X1 #() 
OAI211_X1_895_ (
  .A({ S17867 }),
  .B({ S17577 }),
  .C1({ S17861 }),
  .C2({ S17862 }),
  .ZN({ S17869 })
);
NAND3_X1 #() 
NAND3_X1_2665_ (
  .A1({ S17860 }),
  .A2({ S17869 }),
  .A3({ S14361 }),
  .ZN({ S17870 })
);
NAND3_X1 #() 
NAND3_X1_2666_ (
  .A1({ S17586 }),
  .A2({ S25957[139] }),
  .A3({ S17587 }),
  .ZN({ S17871 })
);
INV_X1 #() 
INV_X1_775_ (
  .A({ S17856 }),
  .ZN({ S17872 })
);
NAND3_X1 #() 
NAND3_X1_2667_ (
  .A1({ S17872 }),
  .A2({ S47 }),
  .A3({ S17632 }),
  .ZN({ S17873 })
);
AOI21_X1 #() 
AOI21_X1_1411_ (
  .A({ S17578 }),
  .B1({ S17873 }),
  .B2({ S17871 }),
  .ZN({ S17874 })
);
OAI22_X1 #() 
OAI22_X1_55_ (
  .A1({ S17682 }),
  .A2({ S17680 }),
  .B1({ S17763 }),
  .B2({ S47 }),
  .ZN({ S17875 })
);
AOI21_X1 #() 
AOI21_X1_1412_ (
  .A({ S17874 }),
  .B1({ S17578 }),
  .B2({ S17875 }),
  .ZN({ S17876 })
);
NOR2_X1 #() 
NOR2_X1_600_ (
  .A1({ S17668 }),
  .A2({ S17669 }),
  .ZN({ S17877 })
);
NOR2_X1 #() 
NOR2_X1_601_ (
  .A1({ S17877 }),
  .A2({ S47 }),
  .ZN({ S17878 })
);
OAI21_X1 #() 
OAI21_X1_1312_ (
  .A({ S17578 }),
  .B1({ S17727 }),
  .B2({ S17621 }),
  .ZN({ S17880 })
);
AOI21_X1 #() 
AOI21_X1_1413_ (
  .A({ S17880 }),
  .B1({ S17878 }),
  .B2({ S17592 }),
  .ZN({ S17881 })
);
NAND2_X1 #() 
NAND2_X1_2474_ (
  .A1({ S17724 }),
  .A2({ S17591 }),
  .ZN({ S17882 })
);
AOI21_X1 #() 
AOI21_X1_1414_ (
  .A({ S17578 }),
  .B1({ S17882 }),
  .B2({ S17755 }),
  .ZN({ S17883 })
);
OAI21_X1 #() 
OAI21_X1_1313_ (
  .A({ S25957[141] }),
  .B1({ S17881 }),
  .B2({ S17883 }),
  .ZN({ S17884 })
);
OAI211_X1 #() 
OAI211_X1_896_ (
  .A({ S17884 }),
  .B({ S25957[142] }),
  .C1({ S17876 }),
  .C2({ S25957[141] }),
  .ZN({ S17885 })
);
NAND3_X1 #() 
NAND3_X1_2668_ (
  .A1({ S17885 }),
  .A2({ S14271 }),
  .A3({ S17870 }),
  .ZN({ S17886 })
);
NAND2_X1 #() 
NAND2_X1_2475_ (
  .A1({ S17850 }),
  .A2({ S17886 }),
  .ZN({ S17887 })
);
XNOR2_X1 #() 
XNOR2_X1_131_ (
  .A({ S17887 }),
  .B({ S25957[242] }),
  .ZN({ S25957[114] })
);
INV_X1 #() 
INV_X1_776_ (
  .A({ S17632 }),
  .ZN({ S17888 })
);
OAI21_X1 #() 
OAI21_X1_1314_ (
  .A({ S25957[139] }),
  .B1({ S25957[136] }),
  .B2({ S17585 }),
  .ZN({ S17890 })
);
OAI22_X1 #() 
OAI22_X1_56_ (
  .A1({ S17877 }),
  .A2({ S17890 }),
  .B1({ S17888 }),
  .B2({ S17583 }),
  .ZN({ S17891 })
);
AOI22_X1 #() 
AOI22_X1_309_ (
  .A1({ S17764 }),
  .A2({ S25957[139] }),
  .B1({ S17592 }),
  .B2({ S17728 }),
  .ZN({ S17892 })
);
MUX2_X1 #() 
MUX2_X1_7_ (
  .A({ S17891 }),
  .B({ S17892 }),
  .S({ S17578 }),
  .Z({ S17893 })
);
NAND2_X1 #() 
NAND2_X1_2476_ (
  .A1({ S17893 }),
  .A2({ S25957[141] }),
  .ZN({ S17894 })
);
NAND2_X1 #() 
NAND2_X1_2477_ (
  .A1({ S17619 }),
  .A2({ S25957[139] }),
  .ZN({ S17895 })
);
INV_X1 #() 
INV_X1_777_ (
  .A({ S17587 }),
  .ZN({ S17896 })
);
OAI22_X1 #() 
OAI22_X1_57_ (
  .A1({ S17697 }),
  .A2({ S47 }),
  .B1({ S17896 }),
  .B2({ S17727 }),
  .ZN({ S17897 })
);
AOI21_X1 #() 
AOI21_X1_1415_ (
  .A({ S25957[140] }),
  .B1({ S17786 }),
  .B2({ S47 }),
  .ZN({ S17898 })
);
AOI22_X1 #() 
AOI22_X1_310_ (
  .A1({ S17897 }),
  .A2({ S25957[140] }),
  .B1({ S17898 }),
  .B2({ S17895 }),
  .ZN({ S17899 })
);
NAND2_X1 #() 
NAND2_X1_2478_ (
  .A1({ S17899 }),
  .A2({ S17577 }),
  .ZN({ S17901 })
);
NAND2_X1 #() 
NAND2_X1_2479_ (
  .A1({ S17894 }),
  .A2({ S17901 }),
  .ZN({ S17902 })
);
NAND2_X1 #() 
NAND2_X1_2480_ (
  .A1({ S17902 }),
  .A2({ S14361 }),
  .ZN({ S17903 })
);
INV_X1 #() 
INV_X1_778_ (
  .A({ S17591 }),
  .ZN({ S17904 })
);
OAI211_X1 #() 
OAI211_X1_897_ (
  .A({ S17640 }),
  .B({ S25957[140] }),
  .C1({ S17732 }),
  .C2({ S17904 }),
  .ZN({ S17905 })
);
NOR2_X1 #() 
NOR2_X1_602_ (
  .A1({ S61 }),
  .A2({ S25957[140] }),
  .ZN({ S17906 })
);
NAND3_X1 #() 
NAND3_X1_2669_ (
  .A1({ S17906 }),
  .A2({ S25957[139] }),
  .A3({ S17769 }),
  .ZN({ S17907 })
);
NOR2_X1 #() 
NOR2_X1_603_ (
  .A1({ S17851 }),
  .A2({ S25957[139] }),
  .ZN({ S17908 })
);
NOR2_X1 #() 
NOR2_X1_604_ (
  .A1({ S17904 }),
  .A2({ S25957[140] }),
  .ZN({ S17909 })
);
AOI21_X1 #() 
AOI21_X1_1416_ (
  .A({ S17577 }),
  .B1({ S17908 }),
  .B2({ S17909 }),
  .ZN({ S17910 })
);
AND3_X1 #() 
AND3_X1_106_ (
  .A1({ S17905 }),
  .A2({ S17910 }),
  .A3({ S17907 }),
  .ZN({ S17912 })
);
NAND4_X1 #() 
NAND4_X1_323_ (
  .A1({ S17618 }),
  .A2({ S17608 }),
  .A3({ S17582 }),
  .A4({ S47 }),
  .ZN({ S17913 })
);
INV_X1 #() 
INV_X1_779_ (
  .A({ S17651 }),
  .ZN({ S17914 })
);
NAND2_X1 #() 
NAND2_X1_2481_ (
  .A1({ S17578 }),
  .A2({ S17914 }),
  .ZN({ S17915 })
);
OAI21_X1 #() 
OAI21_X1_1315_ (
  .A({ S17577 }),
  .B1({ S17915 }),
  .B2({ S17786 }),
  .ZN({ S17916 })
);
AOI21_X1 #() 
AOI21_X1_1417_ (
  .A({ S17916 }),
  .B1({ S17913 }),
  .B2({ S17739 }),
  .ZN({ S17917 })
);
OAI21_X1 #() 
OAI21_X1_1316_ (
  .A({ S25957[142] }),
  .B1({ S17912 }),
  .B2({ S17917 }),
  .ZN({ S17918 })
);
NAND3_X1 #() 
NAND3_X1_2670_ (
  .A1({ S17903 }),
  .A2({ S17918 }),
  .A3({ S25957[143] }),
  .ZN({ S17919 })
);
NOR2_X1 #() 
NOR2_X1_605_ (
  .A1({ S17856 }),
  .A2({ S25957[139] }),
  .ZN({ S17920 })
);
NAND2_X1 #() 
NAND2_X1_2482_ (
  .A1({ S17920 }),
  .A2({ S17618 }),
  .ZN({ S17921 })
);
NAND3_X1 #() 
NAND3_X1_2671_ (
  .A1({ S17632 }),
  .A2({ S25957[139] }),
  .A3({ S17582 }),
  .ZN({ S17923 })
);
NAND2_X1 #() 
NAND2_X1_2483_ (
  .A1({ S17923 }),
  .A2({ S25957[140] }),
  .ZN({ S17924 })
);
INV_X1 #() 
INV_X1_780_ (
  .A({ S17924 }),
  .ZN({ S17925 })
);
AOI21_X1 #() 
AOI21_X1_1418_ (
  .A({ S17646 }),
  .B1({ S17728 }),
  .B2({ S17591 }),
  .ZN({ S17926 })
);
AOI22_X1 #() 
AOI22_X1_311_ (
  .A1({ S17926 }),
  .A2({ S17578 }),
  .B1({ S17925 }),
  .B2({ S17921 }),
  .ZN({ S17927 })
);
NAND2_X1 #() 
NAND2_X1_2484_ (
  .A1({ S17927 }),
  .A2({ S25957[141] }),
  .ZN({ S17928 })
);
INV_X1 #() 
INV_X1_781_ (
  .A({ S17677 }),
  .ZN({ S17929 })
);
NAND2_X1 #() 
NAND2_X1_2485_ (
  .A1({ S17755 }),
  .A2({ S25957[140] }),
  .ZN({ S17930 })
);
OAI21_X1 #() 
OAI21_X1_1317_ (
  .A({ S17578 }),
  .B1({ S17751 }),
  .B2({ S17822 }),
  .ZN({ S17931 })
);
OAI211_X1 #() 
OAI211_X1_898_ (
  .A({ S17930 }),
  .B({ S17577 }),
  .C1({ S17929 }),
  .C2({ S17931 }),
  .ZN({ S17932 })
);
NAND3_X1 #() 
NAND3_X1_2672_ (
  .A1({ S17928 }),
  .A2({ S25957[142] }),
  .A3({ S17932 }),
  .ZN({ S17934 })
);
NOR2_X1 #() 
NOR2_X1_606_ (
  .A1({ S17757 }),
  .A2({ S17856 }),
  .ZN({ S17935 })
);
NOR2_X1 #() 
NOR2_X1_607_ (
  .A1({ S17721 }),
  .A2({ S25957[139] }),
  .ZN({ S17936 })
);
OAI21_X1 #() 
OAI21_X1_1318_ (
  .A({ S17578 }),
  .B1({ S17936 }),
  .B2({ S17935 }),
  .ZN({ S17937 })
);
INV_X1 #() 
INV_X1_782_ (
  .A({ S17626 }),
  .ZN({ S17938 })
);
NAND2_X1 #() 
NAND2_X1_2486_ (
  .A1({ S17622 }),
  .A2({ S47 }),
  .ZN({ S17939 })
);
NOR2_X1 #() 
NOR2_X1_608_ (
  .A1({ S17938 }),
  .A2({ S17939 }),
  .ZN({ S17940 })
);
AOI21_X1 #() 
AOI21_X1_1419_ (
  .A({ S17940 }),
  .B1({ S17785 }),
  .B2({ S17786 }),
  .ZN({ S17941 })
);
AOI21_X1 #() 
AOI21_X1_1420_ (
  .A({ S25957[141] }),
  .B1({ S17941 }),
  .B2({ S25957[140] }),
  .ZN({ S17942 })
);
INV_X1 #() 
INV_X1_783_ (
  .A({ S17592 }),
  .ZN({ S17943 })
);
OAI21_X1 #() 
OAI21_X1_1319_ (
  .A({ S17890 }),
  .B1({ S17943 }),
  .B2({ S25957[139] }),
  .ZN({ S17945 })
);
OAI21_X1 #() 
OAI21_X1_1320_ (
  .A({ S25957[141] }),
  .B1({ S17880 }),
  .B2({ S17888 }),
  .ZN({ S17946 })
);
AOI21_X1 #() 
AOI21_X1_1421_ (
  .A({ S17946 }),
  .B1({ S17945 }),
  .B2({ S25957[140] }),
  .ZN({ S17947 })
);
AOI21_X1 #() 
AOI21_X1_1422_ (
  .A({ S17947 }),
  .B1({ S17942 }),
  .B2({ S17937 }),
  .ZN({ S17948 })
);
OAI211_X1 #() 
OAI211_X1_899_ (
  .A({ S17934 }),
  .B({ S14271 }),
  .C1({ S17948 }),
  .C2({ S25957[142] }),
  .ZN({ S17949 })
);
NAND2_X1 #() 
NAND2_X1_2487_ (
  .A1({ S17919 }),
  .A2({ S17949 }),
  .ZN({ S17950 })
);
XNOR2_X1 #() 
XNOR2_X1_132_ (
  .A({ S17950 }),
  .B({ S25957[243] }),
  .ZN({ S25957[115] })
);
AOI21_X1 #() 
AOI21_X1_1423_ (
  .A({ S25957[139] }),
  .B1({ S17697 }),
  .B2({ S17734 }),
  .ZN({ S17951 })
);
AOI211_X1 #() 
AOI211_X1_31_ (
  .A({ S25957[140] }),
  .B({ S17951 }),
  .C1({ S25957[139] }),
  .C2({ S17664 }),
  .ZN({ S17952 })
);
AOI21_X1 #() 
AOI21_X1_1424_ (
  .A({ S17680 }),
  .B1({ S17682 }),
  .B2({ S17784 }),
  .ZN({ S17953 })
);
OAI21_X1 #() 
OAI21_X1_1321_ (
  .A({ S25957[141] }),
  .B1({ S17953 }),
  .B2({ S17578 }),
  .ZN({ S17955 })
);
INV_X1 #() 
INV_X1_784_ (
  .A({ S17766 }),
  .ZN({ S17956 })
);
NOR2_X1 #() 
NOR2_X1_609_ (
  .A1({ S17896 }),
  .A2({ S17956 }),
  .ZN({ S17957 })
);
NOR2_X1 #() 
NOR2_X1_610_ (
  .A1({ S17822 }),
  .A2({ S47 }),
  .ZN({ S17958 })
);
AOI21_X1 #() 
AOI21_X1_1425_ (
  .A({ S17578 }),
  .B1({ S17958 }),
  .B2({ S17655 }),
  .ZN({ S17959 })
);
AOI21_X1 #() 
AOI21_X1_1426_ (
  .A({ S25957[141] }),
  .B1({ S17866 }),
  .B2({ S17959 }),
  .ZN({ S17960 })
);
OAI21_X1 #() 
OAI21_X1_1322_ (
  .A({ S17960 }),
  .B1({ S17746 }),
  .B2({ S17957 }),
  .ZN({ S17961 })
);
OAI211_X1 #() 
OAI211_X1_900_ (
  .A({ S14361 }),
  .B({ S17961 }),
  .C1({ S17952 }),
  .C2({ S17955 }),
  .ZN({ S17962 })
);
NAND2_X1 #() 
NAND2_X1_2488_ (
  .A1({ S17785 }),
  .A2({ S17608 }),
  .ZN({ S17963 })
);
NAND2_X1 #() 
NAND2_X1_2489_ (
  .A1({ S17963 }),
  .A2({ S17771 }),
  .ZN({ S17964 })
);
NAND2_X1 #() 
NAND2_X1_2490_ (
  .A1({ S17590 }),
  .A2({ S47 }),
  .ZN({ S17966 })
);
INV_X1 #() 
INV_X1_785_ (
  .A({ S17966 }),
  .ZN({ S17967 })
);
AOI22_X1 #() 
AOI22_X1_312_ (
  .A1({ S17967 }),
  .A2({ S17596 }),
  .B1({ S17603 }),
  .B2({ S17766 }),
  .ZN({ S17968 })
);
NAND2_X1 #() 
NAND2_X1_2491_ (
  .A1({ S17968 }),
  .A2({ S25957[140] }),
  .ZN({ S17969 })
);
OAI211_X1 #() 
OAI211_X1_901_ (
  .A({ S17969 }),
  .B({ S17577 }),
  .C1({ S25957[140] }),
  .C2({ S17964 }),
  .ZN({ S17970 })
);
NAND2_X1 #() 
NAND2_X1_2492_ (
  .A1({ S17582 }),
  .A2({ S17608 }),
  .ZN({ S17971 })
);
OAI21_X1 #() 
OAI21_X1_1323_ (
  .A({ S25957[140] }),
  .B1({ S17625 }),
  .B2({ S17971 }),
  .ZN({ S17972 })
);
NOR2_X1 #() 
NOR2_X1_611_ (
  .A1({ S17727 }),
  .A2({ S25957[136] }),
  .ZN({ S17973 })
);
NOR2_X1 #() 
NOR2_X1_612_ (
  .A1({ S17778 }),
  .A2({ S17896 }),
  .ZN({ S17974 })
);
OAI21_X1 #() 
OAI21_X1_1324_ (
  .A({ S17578 }),
  .B1({ S17974 }),
  .B2({ S17973 }),
  .ZN({ S17975 })
);
AND2_X1 #() 
AND2_X1_162_ (
  .A1({ S17975 }),
  .A2({ S17972 }),
  .ZN({ S17977 })
);
OAI211_X1 #() 
OAI211_X1_902_ (
  .A({ S17970 }),
  .B({ S25957[142] }),
  .C1({ S17577 }),
  .C2({ S17977 }),
  .ZN({ S17978 })
);
NAND3_X1 #() 
NAND3_X1_2673_ (
  .A1({ S17962 }),
  .A2({ S25957[143] }),
  .A3({ S17978 }),
  .ZN({ S17979 })
);
NAND2_X1 #() 
NAND2_X1_2493_ (
  .A1({ S17590 }),
  .A2({ S17608 }),
  .ZN({ S17980 })
);
AOI22_X1 #() 
AOI22_X1_313_ (
  .A1({ S17625 }),
  .A2({ S17608 }),
  .B1({ S17980 }),
  .B2({ S25957[139] }),
  .ZN({ S17981 })
);
NOR2_X1 #() 
NOR2_X1_613_ (
  .A1({ S17981 }),
  .A2({ S17578 }),
  .ZN({ S17982 })
);
AOI21_X1 #() 
AOI21_X1_1427_ (
  .A({ S17915 }),
  .B1({ S17920 }),
  .B2({ S17602 }),
  .ZN({ S17983 })
);
OAI21_X1 #() 
OAI21_X1_1325_ (
  .A({ S17577 }),
  .B1({ S17982 }),
  .B2({ S17983 }),
  .ZN({ S17984 })
);
NAND3_X1 #() 
NAND3_X1_2674_ (
  .A1({ S25957[140] }),
  .A2({ S154 }),
  .A3({ S17581 }),
  .ZN({ S17985 })
);
OAI21_X1 #() 
OAI21_X1_1326_ (
  .A({ S17604 }),
  .B1({ S17615 }),
  .B2({ S17732 }),
  .ZN({ S17986 })
);
NAND2_X1 #() 
NAND2_X1_2494_ (
  .A1({ S17986 }),
  .A2({ S17578 }),
  .ZN({ S17988 })
);
NAND2_X1 #() 
NAND2_X1_2495_ (
  .A1({ S17988 }),
  .A2({ S17985 }),
  .ZN({ S17989 })
);
OAI21_X1 #() 
OAI21_X1_1327_ (
  .A({ S17984 }),
  .B1({ S17577 }),
  .B2({ S17989 }),
  .ZN({ S17990 })
);
NAND3_X1 #() 
NAND3_X1_2675_ (
  .A1({ S17844 }),
  .A2({ S17640 }),
  .A3({ S17673 }),
  .ZN({ S17991 })
);
NAND2_X1 #() 
NAND2_X1_2496_ (
  .A1({ S17573 }),
  .A2({ S47 }),
  .ZN({ S17992 })
);
OAI211_X1 #() 
OAI211_X1_903_ (
  .A({ S17677 }),
  .B({ S25957[140] }),
  .C1({ S17624 }),
  .C2({ S17992 }),
  .ZN({ S17993 })
);
AND2_X1 #() 
AND2_X1_163_ (
  .A1({ S17991 }),
  .A2({ S17993 }),
  .ZN({ S17994 })
);
NAND2_X1 #() 
NAND2_X1_2497_ (
  .A1({ S17863 }),
  .A2({ S47 }),
  .ZN({ S17995 })
);
NAND2_X1 #() 
NAND2_X1_2498_ (
  .A1({ S17784 }),
  .A2({ S17914 }),
  .ZN({ S17996 })
);
NAND2_X1 #() 
NAND2_X1_2499_ (
  .A1({ S17996 }),
  .A2({ S17622 }),
  .ZN({ S17997 })
);
AND2_X1 #() 
AND2_X1_164_ (
  .A1({ S17997 }),
  .A2({ S17995 }),
  .ZN({ S17999 })
);
NAND2_X1 #() 
NAND2_X1_2500_ (
  .A1({ S17996 }),
  .A2({ S17586 }),
  .ZN({ S18000 })
);
NAND3_X1 #() 
NAND3_X1_2676_ (
  .A1({ S18000 }),
  .A2({ S17578 }),
  .A3({ S17992 }),
  .ZN({ S18001 })
);
OAI211_X1 #() 
OAI211_X1_904_ (
  .A({ S25957[141] }),
  .B({ S18001 }),
  .C1({ S17999 }),
  .C2({ S17578 }),
  .ZN({ S18002 })
);
OAI211_X1 #() 
OAI211_X1_905_ (
  .A({ S18002 }),
  .B({ S14361 }),
  .C1({ S25957[141] }),
  .C2({ S17994 }),
  .ZN({ S18003 })
);
OAI21_X1 #() 
OAI21_X1_1328_ (
  .A({ S18003 }),
  .B1({ S14361 }),
  .B2({ S17990 }),
  .ZN({ S18004 })
);
NAND2_X1 #() 
NAND2_X1_2501_ (
  .A1({ S18004 }),
  .A2({ S14271 }),
  .ZN({ S18005 })
);
NAND2_X1 #() 
NAND2_X1_2502_ (
  .A1({ S18005 }),
  .A2({ S17979 }),
  .ZN({ S18006 })
);
XNOR2_X1 #() 
XNOR2_X1_133_ (
  .A({ S18006 }),
  .B({ S25957[244] }),
  .ZN({ S25957[116] })
);
AOI21_X1 #() 
AOI21_X1_1428_ (
  .A({ S17852 }),
  .B1({ S17664 }),
  .B2({ S47 }),
  .ZN({ S18007 })
);
OAI21_X1 #() 
OAI21_X1_1329_ (
  .A({ S17578 }),
  .B1({ S17601 }),
  .B2({ S17605 }),
  .ZN({ S18009 })
);
NAND2_X1 #() 
NAND2_X1_2503_ (
  .A1({ S17980 }),
  .A2({ S17582 }),
  .ZN({ S18010 })
);
AOI21_X1 #() 
AOI21_X1_1429_ (
  .A({ S18009 }),
  .B1({ S25957[139] }),
  .B2({ S18010 }),
  .ZN({ S18011 })
);
NOR2_X1 #() 
NOR2_X1_614_ (
  .A1({ S18007 }),
  .A2({ S18011 }),
  .ZN({ S18012 })
);
NAND2_X1 #() 
NAND2_X1_2504_ (
  .A1({ S18012 }),
  .A2({ S25957[141] }),
  .ZN({ S18013 })
);
NAND2_X1 #() 
NAND2_X1_2505_ (
  .A1({ S17943 }),
  .A2({ S47 }),
  .ZN({ S18014 })
);
AOI21_X1 #() 
AOI21_X1_1430_ (
  .A({ S25957[140] }),
  .B1({ S18014 }),
  .B2({ S17923 }),
  .ZN({ S18015 })
);
AOI211_X1 #() 
AOI211_X1_32_ (
  .A({ S17578 }),
  .B({ S17696 }),
  .C1({ S47 }),
  .C2({ S17637 }),
  .ZN({ S18016 })
);
OAI21_X1 #() 
OAI21_X1_1330_ (
  .A({ S17577 }),
  .B1({ S18015 }),
  .B2({ S18016 }),
  .ZN({ S18017 })
);
NAND3_X1 #() 
NAND3_X1_2677_ (
  .A1({ S18013 }),
  .A2({ S25957[142] }),
  .A3({ S18017 }),
  .ZN({ S18018 })
);
OAI21_X1 #() 
OAI21_X1_1331_ (
  .A({ S17956 }),
  .B1({ S17966 }),
  .B2({ S17630 }),
  .ZN({ S18020 })
);
NOR2_X1 #() 
NOR2_X1_615_ (
  .A1({ S17583 }),
  .A2({ S61 }),
  .ZN({ S18021 })
);
NAND2_X1 #() 
NAND2_X1_2506_ (
  .A1({ S17958 }),
  .A2({ S25957[136] }),
  .ZN({ S18022 })
);
NAND2_X1 #() 
NAND2_X1_2507_ (
  .A1({ S18022 }),
  .A2({ S25957[140] }),
  .ZN({ S18023 })
);
OAI22_X1 #() 
OAI22_X1_58_ (
  .A1({ S18023 }),
  .A2({ S18021 }),
  .B1({ S18020 }),
  .B2({ S25957[140] }),
  .ZN({ S18024 })
);
NAND2_X1 #() 
NAND2_X1_2508_ (
  .A1({ S18024 }),
  .A2({ S25957[141] }),
  .ZN({ S18025 })
);
OAI21_X1 #() 
OAI21_X1_1332_ (
  .A({ S17660 }),
  .B1({ S17735 }),
  .B2({ S17601 }),
  .ZN({ S18026 })
);
NOR2_X1 #() 
NOR2_X1_616_ (
  .A1({ S17920 }),
  .A2({ S25957[140] }),
  .ZN({ S18027 })
);
AOI22_X1 #() 
AOI22_X1_314_ (
  .A1({ S18027 }),
  .A2({ S18026 }),
  .B1({ S18000 }),
  .B2({ S17837 }),
  .ZN({ S18028 })
);
OAI21_X1 #() 
OAI21_X1_1333_ (
  .A({ S18025 }),
  .B1({ S18028 }),
  .B2({ S25957[141] }),
  .ZN({ S18029 })
);
NAND2_X1 #() 
NAND2_X1_2509_ (
  .A1({ S18029 }),
  .A2({ S14361 }),
  .ZN({ S18030 })
);
NAND3_X1 #() 
NAND3_X1_2678_ (
  .A1({ S18030 }),
  .A2({ S25957[143] }),
  .A3({ S18018 }),
  .ZN({ S18031 })
);
OAI21_X1 #() 
OAI21_X1_1334_ (
  .A({ S17685 }),
  .B1({ S17593 }),
  .B2({ S47 }),
  .ZN({ S18032 })
);
OAI221_X1 #() 
OAI221_X1_61_ (
  .A({ S17578 }),
  .B1({ S17621 }),
  .B2({ S17914 }),
  .C1({ S17764 }),
  .C2({ S25957[139] }),
  .ZN({ S18033 })
);
OAI21_X1 #() 
OAI21_X1_1335_ (
  .A({ S18033 }),
  .B1({ S17578 }),
  .B2({ S18032 }),
  .ZN({ S18034 })
);
NOR3_X1 #() 
NOR3_X1_83_ (
  .A1({ S17750 }),
  .A2({ S17971 }),
  .A3({ S47 }),
  .ZN({ S18035 })
);
NAND2_X1 #() 
NAND2_X1_2510_ (
  .A1({ S17634 }),
  .A2({ S25957[140] }),
  .ZN({ S18036 })
);
AOI21_X1 #() 
AOI21_X1_1431_ (
  .A({ S17621 }),
  .B1({ S17956 }),
  .B2({ S17675 }),
  .ZN({ S18037 })
);
OAI221_X1 #() 
OAI221_X1_62_ (
  .A({ S17577 }),
  .B1({ S25957[140] }),
  .B2({ S18037 }),
  .C1({ S18035 }),
  .C2({ S18036 }),
  .ZN({ S18038 })
);
OAI211_X1 #() 
OAI211_X1_906_ (
  .A({ S18038 }),
  .B({ S14361 }),
  .C1({ S17577 }),
  .C2({ S18034 }),
  .ZN({ S18039 })
);
OAI211_X1 #() 
OAI211_X1_907_ (
  .A({ S17604 }),
  .B({ S17578 }),
  .C1({ S17680 }),
  .C2({ S17745 }),
  .ZN({ S18041 })
);
AOI22_X1 #() 
AOI22_X1_315_ (
  .A1({ S17735 }),
  .A2({ S47 }),
  .B1({ S17992 }),
  .B2({ S17971 }),
  .ZN({ S18042 })
);
OAI21_X1 #() 
OAI21_X1_1336_ (
  .A({ S18041 }),
  .B1({ S18042 }),
  .B2({ S17578 }),
  .ZN({ S18043 })
);
NOR2_X1 #() 
NOR2_X1_617_ (
  .A1({ S17750 }),
  .A2({ S17725 }),
  .ZN({ S18044 })
);
OAI21_X1 #() 
OAI21_X1_1337_ (
  .A({ S25957[140] }),
  .B1({ S17938 }),
  .B2({ S17939 }),
  .ZN({ S18045 })
);
OAI22_X1 #() 
OAI22_X1_59_ (
  .A1({ S17966 }),
  .A2({ S17853 }),
  .B1({ S25957[136] }),
  .B2({ S47 }),
  .ZN({ S18046 })
);
OAI221_X1 #() 
OAI221_X1_63_ (
  .A({ S25957[141] }),
  .B1({ S25957[140] }),
  .B2({ S18046 }),
  .C1({ S18044 }),
  .C2({ S18045 }),
  .ZN({ S18047 })
);
OAI211_X1 #() 
OAI211_X1_908_ (
  .A({ S18047 }),
  .B({ S25957[142] }),
  .C1({ S25957[141] }),
  .C2({ S18043 }),
  .ZN({ S18048 })
);
NAND3_X1 #() 
NAND3_X1_2679_ (
  .A1({ S18039 }),
  .A2({ S14271 }),
  .A3({ S18048 }),
  .ZN({ S18049 })
);
NAND2_X1 #() 
NAND2_X1_2511_ (
  .A1({ S18031 }),
  .A2({ S18049 }),
  .ZN({ S18050 })
);
XNOR2_X1 #() 
XNOR2_X1_134_ (
  .A({ S18050 }),
  .B({ S25957[245] }),
  .ZN({ S25957[117] })
);
INV_X1 #() 
INV_X1_786_ (
  .A({ S25957[246] }),
  .ZN({ S18051 })
);
NAND3_X1 #() 
NAND3_X1_2680_ (
  .A1({ S17573 }),
  .A2({ S25957[139] }),
  .A3({ S17585 }),
  .ZN({ S18052 })
);
OAI211_X1 #() 
OAI211_X1_909_ (
  .A({ S18052 }),
  .B({ S17578 }),
  .C1({ S25957[139] }),
  .C2({ S17575 }),
  .ZN({ S18053 })
);
NAND3_X1 #() 
NAND3_X1_2681_ (
  .A1({ S17633 }),
  .A2({ S17820 }),
  .A3({ S25957[140] }),
  .ZN({ S18054 })
);
NAND3_X1 #() 
NAND3_X1_2682_ (
  .A1({ S18054 }),
  .A2({ S25957[141] }),
  .A3({ S18053 }),
  .ZN({ S18055 })
);
NAND2_X1 #() 
NAND2_X1_2512_ (
  .A1({ S17920 }),
  .A2({ S17656 }),
  .ZN({ S18056 })
);
NAND2_X1 #() 
NAND2_X1_2513_ (
  .A1({ S17925 }),
  .A2({ S18056 }),
  .ZN({ S18057 })
);
OAI21_X1 #() 
OAI21_X1_1338_ (
  .A({ S17777 }),
  .B1({ S17865 }),
  .B2({ S17890 }),
  .ZN({ S18058 })
);
NAND3_X1 #() 
NAND3_X1_2683_ (
  .A1({ S18058 }),
  .A2({ S18057 }),
  .A3({ S17577 }),
  .ZN({ S18059 })
);
AOI21_X1 #() 
AOI21_X1_1432_ (
  .A({ S14361 }),
  .B1({ S18059 }),
  .B2({ S18055 }),
  .ZN({ S18061 })
);
NAND2_X1 #() 
NAND2_X1_2514_ (
  .A1({ S17591 }),
  .A2({ S17590 }),
  .ZN({ S18062 })
);
OAI22_X1 #() 
OAI22_X1_60_ (
  .A1({ S17744 }),
  .A2({ S47 }),
  .B1({ S18062 }),
  .B2({ S17727 }),
  .ZN({ S18063 })
);
NAND2_X1 #() 
NAND2_X1_2515_ (
  .A1({ S18063 }),
  .A2({ S17578 }),
  .ZN({ S18064 })
);
NAND2_X1 #() 
NAND2_X1_2516_ (
  .A1({ S17618 }),
  .A2({ S47 }),
  .ZN({ S18065 })
);
OAI21_X1 #() 
OAI21_X1_1339_ (
  .A({ S17654 }),
  .B1({ S18065 }),
  .B2({ S17696 }),
  .ZN({ S18066 })
);
NAND3_X1 #() 
NAND3_X1_2684_ (
  .A1({ S18064 }),
  .A2({ S18066 }),
  .A3({ S25957[141] }),
  .ZN({ S18067 })
);
AOI21_X1 #() 
AOI21_X1_1433_ (
  .A({ S17578 }),
  .B1({ S17980 }),
  .B2({ S25957[139] }),
  .ZN({ S18068 })
);
OAI21_X1 #() 
OAI21_X1_1340_ (
  .A({ S18068 }),
  .B1({ S25957[139] }),
  .B2({ S17971 }),
  .ZN({ S18069 })
);
NAND3_X1 #() 
NAND3_X1_2685_ (
  .A1({ S17645 }),
  .A2({ S25957[139] }),
  .A3({ S17587 }),
  .ZN({ S18070 })
);
NAND3_X1 #() 
NAND3_X1_2686_ (
  .A1({ S18056 }),
  .A2({ S17578 }),
  .A3({ S18070 }),
  .ZN({ S18071 })
);
NAND3_X1 #() 
NAND3_X1_2687_ (
  .A1({ S18071 }),
  .A2({ S17577 }),
  .A3({ S18069 }),
  .ZN({ S18072 })
);
AOI21_X1 #() 
AOI21_X1_1434_ (
  .A({ S25957[142] }),
  .B1({ S18072 }),
  .B2({ S18067 }),
  .ZN({ S18073 })
);
OAI21_X1 #() 
OAI21_X1_1341_ (
  .A({ S25957[143] }),
  .B1({ S18061 }),
  .B2({ S18073 }),
  .ZN({ S18074 })
);
OAI21_X1 #() 
OAI21_X1_1342_ (
  .A({ S17793 }),
  .B1({ S17786 }),
  .B2({ S47 }),
  .ZN({ S18075 })
);
OAI21_X1 #() 
OAI21_X1_1343_ (
  .A({ S17578 }),
  .B1({ S17767 }),
  .B2({ S17763 }),
  .ZN({ S18076 })
);
OAI211_X1 #() 
OAI211_X1_910_ (
  .A({ S25957[141] }),
  .B({ S18076 }),
  .C1({ S18075 }),
  .C2({ S17578 }),
  .ZN({ S18077 })
);
NAND2_X1 #() 
NAND2_X1_2517_ (
  .A1({ S17914 }),
  .A2({ S17596 }),
  .ZN({ S18078 })
);
NAND2_X1 #() 
NAND2_X1_2518_ (
  .A1({ S18065 }),
  .A2({ S17923 }),
  .ZN({ S18079 })
);
NAND2_X1 #() 
NAND2_X1_2519_ (
  .A1({ S18079 }),
  .A2({ S17578 }),
  .ZN({ S18080 })
);
OAI211_X1 #() 
OAI211_X1_911_ (
  .A({ S18080 }),
  .B({ S17577 }),
  .C1({ S17752 }),
  .C2({ S18078 }),
  .ZN({ S18082 })
);
NAND2_X1 #() 
NAND2_X1_2520_ (
  .A1({ S18082 }),
  .A2({ S18077 }),
  .ZN({ S18083 })
);
NAND2_X1 #() 
NAND2_X1_2521_ (
  .A1({ S18083 }),
  .A2({ S25957[142] }),
  .ZN({ S18084 })
);
OAI21_X1 #() 
OAI21_X1_1344_ (
  .A({ S17752 }),
  .B1({ S17578 }),
  .B2({ S17630 }),
  .ZN({ S18085 })
);
NAND2_X1 #() 
NAND2_X1_2522_ (
  .A1({ S18085 }),
  .A2({ S17997 }),
  .ZN({ S18086 })
);
NAND3_X1 #() 
NAND3_X1_2688_ (
  .A1({ S18086 }),
  .A2({ S17577 }),
  .A3({ S17861 }),
  .ZN({ S18087 })
);
OR3_X1 #() 
OR3_X1_14_ (
  .A1({ S17940 }),
  .A2({ S17958 }),
  .A3({ S25957[140] }),
  .ZN({ S18088 })
);
NAND3_X1 #() 
NAND3_X1_2689_ (
  .A1({ S17872 }),
  .A2({ S25957[139] }),
  .A3({ S17592 }),
  .ZN({ S18089 })
);
NAND3_X1 #() 
NAND3_X1_2690_ (
  .A1({ S18089 }),
  .A2({ S25957[140] }),
  .A3({ S17638 }),
  .ZN({ S18090 })
);
NAND3_X1 #() 
NAND3_X1_2691_ (
  .A1({ S18088 }),
  .A2({ S25957[141] }),
  .A3({ S18090 }),
  .ZN({ S18091 })
);
NAND3_X1 #() 
NAND3_X1_2692_ (
  .A1({ S18091 }),
  .A2({ S18087 }),
  .A3({ S14361 }),
  .ZN({ S18093 })
);
NAND3_X1 #() 
NAND3_X1_2693_ (
  .A1({ S18084 }),
  .A2({ S14271 }),
  .A3({ S18093 }),
  .ZN({ S18094 })
);
NAND3_X1 #() 
NAND3_X1_2694_ (
  .A1({ S18094 }),
  .A2({ S18074 }),
  .A3({ S18051 }),
  .ZN({ S18095 })
);
AOI21_X1 #() 
AOI21_X1_1435_ (
  .A({ S25957[143] }),
  .B1({ S18082 }),
  .B2({ S18077 }),
  .ZN({ S18096 })
);
AND3_X1 #() 
AND3_X1_107_ (
  .A1({ S18059 }),
  .A2({ S18055 }),
  .A3({ S25957[143] }),
  .ZN({ S18097 })
);
OAI21_X1 #() 
OAI21_X1_1345_ (
  .A({ S25957[142] }),
  .B1({ S18096 }),
  .B2({ S18097 }),
  .ZN({ S18098 })
);
NAND3_X1 #() 
NAND3_X1_2695_ (
  .A1({ S18091 }),
  .A2({ S18087 }),
  .A3({ S14271 }),
  .ZN({ S18099 })
);
NAND3_X1 #() 
NAND3_X1_2696_ (
  .A1({ S18072 }),
  .A2({ S18067 }),
  .A3({ S25957[143] }),
  .ZN({ S18100 })
);
NAND2_X1 #() 
NAND2_X1_2523_ (
  .A1({ S18099 }),
  .A2({ S18100 }),
  .ZN({ S18101 })
);
NAND2_X1 #() 
NAND2_X1_2524_ (
  .A1({ S18101 }),
  .A2({ S14361 }),
  .ZN({ S18102 })
);
NAND3_X1 #() 
NAND3_X1_2697_ (
  .A1({ S18098 }),
  .A2({ S18102 }),
  .A3({ S25957[246] }),
  .ZN({ S18104 })
);
NAND2_X1 #() 
NAND2_X1_2525_ (
  .A1({ S18095 }),
  .A2({ S18104 }),
  .ZN({ S25957[118] })
);
NAND3_X1 #() 
NAND3_X1_2698_ (
  .A1({ S17582 }),
  .A2({ S47 }),
  .A3({ S25957[137] }),
  .ZN({ S18105 })
);
AOI21_X1 #() 
AOI21_X1_1436_ (
  .A({ S17578 }),
  .B1({ S17677 }),
  .B2({ S18105 }),
  .ZN({ S18106 })
);
NOR2_X1 #() 
NOR2_X1_618_ (
  .A1({ S17843 }),
  .A2({ S17904 }),
  .ZN({ S18107 })
);
AOI21_X1 #() 
AOI21_X1_1437_ (
  .A({ S25957[139] }),
  .B1({ S17786 }),
  .B2({ S17596 }),
  .ZN({ S18108 })
);
NOR3_X1 #() 
NOR3_X1_84_ (
  .A1({ S18108 }),
  .A2({ S18107 }),
  .A3({ S25957[140] }),
  .ZN({ S18109 })
);
OAI21_X1 #() 
OAI21_X1_1346_ (
  .A({ S25957[141] }),
  .B1({ S18109 }),
  .B2({ S18106 }),
  .ZN({ S18110 })
);
AOI21_X1 #() 
AOI21_X1_1438_ (
  .A({ S17578 }),
  .B1({ S18052 }),
  .B2({ S17966 }),
  .ZN({ S18111 })
);
NAND2_X1 #() 
NAND2_X1_2526_ (
  .A1({ S17660 }),
  .A2({ S17608 }),
  .ZN({ S18112 })
);
AND3_X1 #() 
AND3_X1_108_ (
  .A1({ S17844 }),
  .A2({ S18112 }),
  .A3({ S17673 }),
  .ZN({ S18114 })
);
OAI21_X1 #() 
OAI21_X1_1347_ (
  .A({ S17577 }),
  .B1({ S18114 }),
  .B2({ S18111 }),
  .ZN({ S18115 })
);
NAND2_X1 #() 
NAND2_X1_2527_ (
  .A1({ S18110 }),
  .A2({ S18115 }),
  .ZN({ S18116 })
);
NAND2_X1 #() 
NAND2_X1_2528_ (
  .A1({ S18116 }),
  .A2({ S25957[142] }),
  .ZN({ S18117 })
);
NAND2_X1 #() 
NAND2_X1_2529_ (
  .A1({ S17980 }),
  .A2({ S47 }),
  .ZN({ S18118 })
);
NAND3_X1 #() 
NAND3_X1_2699_ (
  .A1({ S17768 }),
  .A2({ S25957[140] }),
  .A3({ S18118 }),
  .ZN({ S18119 })
);
NAND2_X1 #() 
NAND2_X1_2530_ (
  .A1({ S17906 }),
  .A2({ S17796 }),
  .ZN({ S18120 })
);
NAND3_X1 #() 
NAND3_X1_2700_ (
  .A1({ S18119 }),
  .A2({ S25957[141] }),
  .A3({ S18120 }),
  .ZN({ S18121 })
);
NAND2_X1 #() 
NAND2_X1_2531_ (
  .A1({ S17670 }),
  .A2({ S17603 }),
  .ZN({ S18122 })
);
OAI211_X1 #() 
OAI211_X1_912_ (
  .A({ S25957[140] }),
  .B({ S18122 }),
  .C1({ S18000 }),
  .C2({ S17943 }),
  .ZN({ S18123 })
);
OAI211_X1 #() 
OAI211_X1_913_ (
  .A({ S17578 }),
  .B({ S17778 }),
  .C1({ S17615 }),
  .C2({ S17682 }),
  .ZN({ S18125 })
);
NAND3_X1 #() 
NAND3_X1_2701_ (
  .A1({ S18123 }),
  .A2({ S18125 }),
  .A3({ S17577 }),
  .ZN({ S18126 })
);
AND2_X1 #() 
AND2_X1_165_ (
  .A1({ S18126 }),
  .A2({ S18121 }),
  .ZN({ S18127 })
);
OAI211_X1 #() 
OAI211_X1_914_ (
  .A({ S18117 }),
  .B({ S25957[143] }),
  .C1({ S25957[142] }),
  .C2({ S18127 }),
  .ZN({ S18128 })
);
INV_X1 #() 
INV_X1_787_ (
  .A({ S17841 }),
  .ZN({ S18129 })
);
OAI21_X1 #() 
OAI21_X1_1348_ (
  .A({ S25957[140] }),
  .B1({ S17936 }),
  .B2({ S17743 }),
  .ZN({ S18130 })
);
OAI211_X1 #() 
OAI211_X1_915_ (
  .A({ S18130 }),
  .B({ S17577 }),
  .C1({ S18129 }),
  .C2({ S17931 }),
  .ZN({ S18131 })
);
NAND3_X1 #() 
NAND3_X1_2702_ (
  .A1({ S17997 }),
  .A2({ S17578 }),
  .A3({ S17736 }),
  .ZN({ S18132 })
);
NAND3_X1 #() 
NAND3_X1_2703_ (
  .A1({ S17786 }),
  .A2({ S25957[139] }),
  .A3({ S17596 }),
  .ZN({ S18133 })
);
NAND2_X1 #() 
NAND2_X1_2532_ (
  .A1({ S17720 }),
  .A2({ S18133 }),
  .ZN({ S18134 })
);
NAND2_X1 #() 
NAND2_X1_2533_ (
  .A1({ S18132 }),
  .A2({ S18134 }),
  .ZN({ S18136 })
);
AOI21_X1 #() 
AOI21_X1_1439_ (
  .A({ S14361 }),
  .B1({ S18136 }),
  .B2({ S25957[141] }),
  .ZN({ S18137 })
);
NAND2_X1 #() 
NAND2_X1_2534_ (
  .A1({ S18131 }),
  .A2({ S18137 }),
  .ZN({ S18138 })
);
NAND3_X1 #() 
NAND3_X1_2704_ (
  .A1({ S17921 }),
  .A2({ S25957[140] }),
  .A3({ S17843 }),
  .ZN({ S18139 })
);
OAI211_X1 #() 
OAI211_X1_916_ (
  .A({ S18014 }),
  .B({ S17578 }),
  .C1({ S47 }),
  .C2({ S17734 }),
  .ZN({ S18140 })
);
NAND3_X1 #() 
NAND3_X1_2705_ (
  .A1({ S18140 }),
  .A2({ S18139 }),
  .A3({ S17577 }),
  .ZN({ S18141 })
);
NAND2_X1 #() 
NAND2_X1_2535_ (
  .A1({ S17967 }),
  .A2({ S17822 }),
  .ZN({ S18142 })
);
AOI21_X1 #() 
AOI21_X1_1440_ (
  .A({ S25957[140] }),
  .B1({ S17963 }),
  .B2({ S18142 }),
  .ZN({ S18143 })
);
NOR2_X1 #() 
NOR2_X1_619_ (
  .A1({ S17974 }),
  .A2({ S17752 }),
  .ZN({ S18144 })
);
OR3_X1 #() 
OR3_X1_15_ (
  .A1({ S18143 }),
  .A2({ S18144 }),
  .A3({ S17577 }),
  .ZN({ S18145 })
);
NAND3_X1 #() 
NAND3_X1_2706_ (
  .A1({ S18145 }),
  .A2({ S14361 }),
  .A3({ S18141 }),
  .ZN({ S18147 })
);
NAND3_X1 #() 
NAND3_X1_2707_ (
  .A1({ S18138 }),
  .A2({ S18147 }),
  .A3({ S14271 }),
  .ZN({ S18148 })
);
NAND3_X1 #() 
NAND3_X1_2708_ (
  .A1({ S18128 }),
  .A2({ S18148 }),
  .A3({ S25957[247] }),
  .ZN({ S18149 })
);
AND2_X1 #() 
AND2_X1_166_ (
  .A1({ S18138 }),
  .A2({ S18147 }),
  .ZN({ S18150 })
);
AOI21_X1 #() 
AOI21_X1_1441_ (
  .A({ S14361 }),
  .B1({ S18110 }),
  .B2({ S18115 }),
  .ZN({ S18151 })
);
AOI21_X1 #() 
AOI21_X1_1442_ (
  .A({ S25957[142] }),
  .B1({ S18126 }),
  .B2({ S18121 }),
  .ZN({ S18152 })
);
OAI21_X1 #() 
OAI21_X1_1349_ (
  .A({ S25957[143] }),
  .B1({ S18152 }),
  .B2({ S18151 }),
  .ZN({ S18153 })
);
OAI211_X1 #() 
OAI211_X1_917_ (
  .A({ S18153 }),
  .B({ S13519 }),
  .C1({ S18150 }),
  .C2({ S25957[143] }),
  .ZN({ S18154 })
);
NAND2_X1 #() 
NAND2_X1_2536_ (
  .A1({ S18154 }),
  .A2({ S18149 }),
  .ZN({ S25957[119] })
);
OAI21_X1 #() 
OAI21_X1_1350_ (
  .A({ S25957[400] }),
  .B1({ S16306 }),
  .B2({ S16307 }),
  .ZN({ S18155 })
);
NAND3_X1 #() 
NAND3_X1_2709_ (
  .A1({ S13981 }),
  .A2({ S13949 }),
  .A3({ S11081 }),
  .ZN({ S18157 })
);
AOI21_X1 #() 
AOI21_X1_1443_ (
  .A({ S25957[401] }),
  .B1({ S14069 }),
  .B2({ S14028 }),
  .ZN({ S18158 })
);
AND3_X1 #() 
AND3_X1_109_ (
  .A1({ S14069 }),
  .A2({ S14028 }),
  .A3({ S25957[401] }),
  .ZN({ S18159 })
);
OAI211_X1 #() 
OAI211_X1_918_ (
  .A({ S18155 }),
  .B({ S18157 }),
  .C1({ S18159 }),
  .C2({ S18158 }),
  .ZN({ S18160 })
);
INV_X1 #() 
INV_X1_788_ (
  .A({ S18160 }),
  .ZN({ S63 })
);
OAI211_X1 #() 
OAI211_X1_919_ (
  .A({ S14027 }),
  .B({ S14070 }),
  .C1({ S13983 }),
  .C2({ S13982 }),
  .ZN({ S64 })
);
NOR2_X1 #() 
NOR2_X1_620_ (
  .A1({ S18159 }),
  .A2({ S18158 }),
  .ZN({ S18161 })
);
AOI21_X1 #() 
AOI21_X1_1444_ (
  .A({ S14119 }),
  .B1({ S14133 }),
  .B2({ S14130 }),
  .ZN({ S18162 })
);
AOI21_X1 #() 
AOI21_X1_1445_ (
  .A({ S25957[466] }),
  .B1({ S14093 }),
  .B2({ S14116 }),
  .ZN({ S18163 })
);
OAI21_X1 #() 
OAI21_X1_1351_ (
  .A({ S25957[402] }),
  .B1({ S18162 }),
  .B2({ S18163 }),
  .ZN({ S18164 })
);
NAND3_X1 #() 
NAND3_X1_2710_ (
  .A1({ S14134 }),
  .A2({ S14118 }),
  .A3({ S11281 }),
  .ZN({ S18166 })
);
NAND2_X1 #() 
NAND2_X1_2537_ (
  .A1({ S18164 }),
  .A2({ S18166 }),
  .ZN({ S18167 })
);
AOI21_X1 #() 
AOI21_X1_1446_ (
  .A({ S25957[144] }),
  .B1({ S18161 }),
  .B2({ S18167 }),
  .ZN({ S18168 })
);
NOR2_X1 #() 
NOR2_X1_621_ (
  .A1({ S25957[147] }),
  .A2({ S18168 }),
  .ZN({ S18169 })
);
NAND2_X1 #() 
NAND2_X1_2538_ (
  .A1({ S18155 }),
  .A2({ S18157 }),
  .ZN({ S18170 })
);
NAND2_X1 #() 
NAND2_X1_2539_ (
  .A1({ S18167 }),
  .A2({ S18170 }),
  .ZN({ S18171 })
);
NAND3_X1 #() 
NAND3_X1_2711_ (
  .A1({ S25957[146] }),
  .A2({ S25957[144] }),
  .A3({ S25957[145] }),
  .ZN({ S18172 })
);
NAND4_X1 #() 
NAND4_X1_324_ (
  .A1({ S18164 }),
  .A2({ S18155 }),
  .A3({ S18157 }),
  .A4({ S18166 }),
  .ZN({ S18173 })
);
NAND2_X1 #() 
NAND2_X1_2540_ (
  .A1({ S18173 }),
  .A2({ S18161 }),
  .ZN({ S18174 })
);
NAND4_X1 #() 
NAND4_X1_325_ (
  .A1({ S25957[147] }),
  .A2({ S18171 }),
  .A3({ S18172 }),
  .A4({ S18174 }),
  .ZN({ S18175 })
);
NAND2_X1 #() 
NAND2_X1_2541_ (
  .A1({ S18175 }),
  .A2({ S25957[148] }),
  .ZN({ S18177 })
);
INV_X1 #() 
INV_X1_789_ (
  .A({ S25957[148] }),
  .ZN({ S18178 })
);
NAND4_X1 #() 
NAND4_X1_326_ (
  .A1({ S18164 }),
  .A2({ S18166 }),
  .A3({ S14027 }),
  .A4({ S14070 }),
  .ZN({ S18179 })
);
OAI22_X1 #() 
OAI22_X1_61_ (
  .A1({ S14136 }),
  .A2({ S14135 }),
  .B1({ S18159 }),
  .B2({ S18158 }),
  .ZN({ S18180 })
);
OAI211_X1 #() 
OAI211_X1_920_ (
  .A({ S18173 }),
  .B({ S18179 }),
  .C1({ S18180 }),
  .C2({ S25957[144] }),
  .ZN({ S18181 })
);
NAND2_X1 #() 
NAND2_X1_2542_ (
  .A1({ S44 }),
  .A2({ S18171 }),
  .ZN({ S18182 })
);
OAI211_X1 #() 
OAI211_X1_921_ (
  .A({ S18182 }),
  .B({ S18178 }),
  .C1({ S44 }),
  .C2({ S18181 }),
  .ZN({ S18183 })
);
OAI211_X1 #() 
OAI211_X1_922_ (
  .A({ S18183 }),
  .B({ S25957[149] }),
  .C1({ S18177 }),
  .C2({ S18169 }),
  .ZN({ S18184 })
);
OR2_X1 #() 
OR2_X1_35_ (
  .A1({ S13613 }),
  .A2({ S13615 }),
  .ZN({ S18185 })
);
INV_X1 #() 
INV_X1_790_ (
  .A({ S18179 }),
  .ZN({ S18186 })
);
OAI22_X1 #() 
OAI22_X1_62_ (
  .A1({ S13983 }),
  .A2({ S13982 }),
  .B1({ S18159 }),
  .B2({ S18158 }),
  .ZN({ S18188 })
);
INV_X1 #() 
INV_X1_791_ (
  .A({ S18188 }),
  .ZN({ S18189 })
);
AOI21_X1 #() 
AOI21_X1_1447_ (
  .A({ S18186 }),
  .B1({ S18167 }),
  .B2({ S18189 }),
  .ZN({ S18190 })
);
NAND2_X1 #() 
NAND2_X1_2543_ (
  .A1({ S25957[147] }),
  .A2({ S18170 }),
  .ZN({ S18191 })
);
NAND3_X1 #() 
NAND3_X1_2712_ (
  .A1({ S18191 }),
  .A2({ S25957[148] }),
  .A3({ S18190 }),
  .ZN({ S18192 })
);
NAND2_X1 #() 
NAND2_X1_2544_ (
  .A1({ S18172 }),
  .A2({ S18171 }),
  .ZN({ S18193 })
);
NAND2_X1 #() 
NAND2_X1_2545_ (
  .A1({ S18193 }),
  .A2({ S25957[147] }),
  .ZN({ S18194 })
);
AOI21_X1 #() 
AOI21_X1_1448_ (
  .A({ S25957[148] }),
  .B1({ S44 }),
  .B2({ S18174 }),
  .ZN({ S18195 })
);
NAND2_X1 #() 
NAND2_X1_2546_ (
  .A1({ S18195 }),
  .A2({ S18194 }),
  .ZN({ S18196 })
);
NAND2_X1 #() 
NAND2_X1_2547_ (
  .A1({ S18196 }),
  .A2({ S18192 }),
  .ZN({ S18197 })
);
AOI21_X1 #() 
AOI21_X1_1449_ (
  .A({ S18185 }),
  .B1({ S18197 }),
  .B2({ S13688 }),
  .ZN({ S18199 })
);
NAND2_X1 #() 
NAND2_X1_2548_ (
  .A1({ S18199 }),
  .A2({ S18184 }),
  .ZN({ S18200 })
);
NAND2_X1 #() 
NAND2_X1_2549_ (
  .A1({ S64 }),
  .A2({ S18173 }),
  .ZN({ S18201 })
);
NAND2_X1 #() 
NAND2_X1_2550_ (
  .A1({ S44 }),
  .A2({ S18201 }),
  .ZN({ S18202 })
);
NAND3_X1 #() 
NAND3_X1_2713_ (
  .A1({ S25957[147] }),
  .A2({ S64 }),
  .A3({ S18173 }),
  .ZN({ S18203 })
);
AND3_X1 #() 
AND3_X1_110_ (
  .A1({ S18203 }),
  .A2({ S18202 }),
  .A3({ S25957[148] }),
  .ZN({ S18204 })
);
NAND3_X1 #() 
NAND3_X1_2714_ (
  .A1({ S18167 }),
  .A2({ S18161 }),
  .A3({ S18170 }),
  .ZN({ S18205 })
);
NAND3_X1 #() 
NAND3_X1_2715_ (
  .A1({ S25957[146] }),
  .A2({ S25957[144] }),
  .A3({ S18161 }),
  .ZN({ S18206 })
);
NAND4_X1 #() 
NAND4_X1_327_ (
  .A1({ S18206 }),
  .A2({ S13895 }),
  .A3({ S18205 }),
  .A4({ S13898 }),
  .ZN({ S18207 })
);
NAND4_X1 #() 
NAND4_X1_328_ (
  .A1({ S18155 }),
  .A2({ S14027 }),
  .A3({ S18157 }),
  .A4({ S14070 }),
  .ZN({ S18208 })
);
NAND3_X1 #() 
NAND3_X1_2716_ (
  .A1({ S18188 }),
  .A2({ S25957[146] }),
  .A3({ S18208 }),
  .ZN({ S18210 })
);
NAND3_X1 #() 
NAND3_X1_2717_ (
  .A1({ S25957[144] }),
  .A2({ S18167 }),
  .A3({ S25957[145] }),
  .ZN({ S18211 })
);
NAND3_X1 #() 
NAND3_X1_2718_ (
  .A1({ S44 }),
  .A2({ S18210 }),
  .A3({ S18211 }),
  .ZN({ S18212 })
);
AOI21_X1 #() 
AOI21_X1_1450_ (
  .A({ S25957[148] }),
  .B1({ S18212 }),
  .B2({ S18207 }),
  .ZN({ S18213 })
);
OAI21_X1 #() 
OAI21_X1_1352_ (
  .A({ S25957[149] }),
  .B1({ S18204 }),
  .B2({ S18213 }),
  .ZN({ S18214 })
);
AOI21_X1 #() 
AOI21_X1_1451_ (
  .A({ S25957[146] }),
  .B1({ S64 }),
  .B2({ S18160 }),
  .ZN({ S18215 })
);
NAND2_X1 #() 
NAND2_X1_2551_ (
  .A1({ S25957[147] }),
  .A2({ S18215 }),
  .ZN({ S18216 })
);
NAND3_X1 #() 
NAND3_X1_2719_ (
  .A1({ S44 }),
  .A2({ S18172 }),
  .A3({ S18174 }),
  .ZN({ S18217 })
);
NAND3_X1 #() 
NAND3_X1_2720_ (
  .A1({ S18217 }),
  .A2({ S25957[148] }),
  .A3({ S18216 }),
  .ZN({ S18218 })
);
NAND3_X1 #() 
NAND3_X1_2721_ (
  .A1({ S25957[146] }),
  .A2({ S18170 }),
  .A3({ S18161 }),
  .ZN({ S18219 })
);
NAND2_X1 #() 
NAND2_X1_2552_ (
  .A1({ S44 }),
  .A2({ S18219 }),
  .ZN({ S18221 })
);
NAND3_X1 #() 
NAND3_X1_2722_ (
  .A1({ S25957[144] }),
  .A2({ S18167 }),
  .A3({ S18161 }),
  .ZN({ S18222 })
);
INV_X1 #() 
INV_X1_792_ (
  .A({ S18222 }),
  .ZN({ S18223 })
);
NAND3_X1 #() 
NAND3_X1_2723_ (
  .A1({ S25957[147] }),
  .A2({ S18205 }),
  .A3({ S18210 }),
  .ZN({ S18224 })
);
OAI211_X1 #() 
OAI211_X1_923_ (
  .A({ S18224 }),
  .B({ S18178 }),
  .C1({ S18221 }),
  .C2({ S18223 }),
  .ZN({ S18225 })
);
NAND3_X1 #() 
NAND3_X1_2724_ (
  .A1({ S18225 }),
  .A2({ S18218 }),
  .A3({ S13688 }),
  .ZN({ S18226 })
);
NAND3_X1 #() 
NAND3_X1_2725_ (
  .A1({ S18214 }),
  .A2({ S18226 }),
  .A3({ S18185 }),
  .ZN({ S18227 })
);
AOI21_X1 #() 
AOI21_X1_1452_ (
  .A({ S25957[151] }),
  .B1({ S18200 }),
  .B2({ S18227 }),
  .ZN({ S18228 })
);
NAND2_X1 #() 
NAND2_X1_2553_ (
  .A1({ S18208 }),
  .A2({ S18167 }),
  .ZN({ S18229 })
);
NAND2_X1 #() 
NAND2_X1_2554_ (
  .A1({ S18229 }),
  .A2({ S18173 }),
  .ZN({ S18230 })
);
NAND2_X1 #() 
NAND2_X1_2555_ (
  .A1({ S25957[147] }),
  .A2({ S18230 }),
  .ZN({ S18232 })
);
NAND3_X1 #() 
NAND3_X1_2726_ (
  .A1({ S25957[145] }),
  .A2({ S18164 }),
  .A3({ S18166 }),
  .ZN({ S18233 })
);
NAND3_X1 #() 
NAND3_X1_2727_ (
  .A1({ S64 }),
  .A2({ S18160 }),
  .A3({ S18167 }),
  .ZN({ S18234 })
);
NAND3_X1 #() 
NAND3_X1_2728_ (
  .A1({ S44 }),
  .A2({ S18233 }),
  .A3({ S18234 }),
  .ZN({ S18235 })
);
AND2_X1 #() 
AND2_X1_167_ (
  .A1({ S18235 }),
  .A2({ S18232 }),
  .ZN({ S18236 })
);
NAND2_X1 #() 
NAND2_X1_2556_ (
  .A1({ S64 }),
  .A2({ S18167 }),
  .ZN({ S18237 })
);
NAND3_X1 #() 
NAND3_X1_2729_ (
  .A1({ S44 }),
  .A2({ S18219 }),
  .A3({ S18237 }),
  .ZN({ S18238 })
);
NAND2_X1 #() 
NAND2_X1_2557_ (
  .A1({ S18179 }),
  .A2({ S18173 }),
  .ZN({ S18239 })
);
NAND2_X1 #() 
NAND2_X1_2558_ (
  .A1({ S25957[147] }),
  .A2({ S18239 }),
  .ZN({ S18240 })
);
NAND3_X1 #() 
NAND3_X1_2730_ (
  .A1({ S18238 }),
  .A2({ S25957[148] }),
  .A3({ S18240 }),
  .ZN({ S18241 })
);
OAI211_X1 #() 
OAI211_X1_924_ (
  .A({ S25957[149] }),
  .B({ S18241 }),
  .C1({ S18236 }),
  .C2({ S25957[148] }),
  .ZN({ S18243 })
);
INV_X1 #() 
INV_X1_793_ (
  .A({ S18210 }),
  .ZN({ S18244 })
);
NAND2_X1 #() 
NAND2_X1_2559_ (
  .A1({ S18244 }),
  .A2({ S25957[147] }),
  .ZN({ S18245 })
);
NAND2_X1 #() 
NAND2_X1_2560_ (
  .A1({ S18189 }),
  .A2({ S18167 }),
  .ZN({ S18246 })
);
NAND3_X1 #() 
NAND3_X1_2731_ (
  .A1({ S44 }),
  .A2({ S18246 }),
  .A3({ S18206 }),
  .ZN({ S18247 })
);
NAND3_X1 #() 
NAND3_X1_2732_ (
  .A1({ S18247 }),
  .A2({ S18245 }),
  .A3({ S25957[148] }),
  .ZN({ S18248 })
);
NAND2_X1 #() 
NAND2_X1_2561_ (
  .A1({ S44 }),
  .A2({ S18246 }),
  .ZN({ S18249 })
);
NAND3_X1 #() 
NAND3_X1_2733_ (
  .A1({ S18194 }),
  .A2({ S18249 }),
  .A3({ S18178 }),
  .ZN({ S18250 })
);
NAND3_X1 #() 
NAND3_X1_2734_ (
  .A1({ S18248 }),
  .A2({ S18250 }),
  .A3({ S13688 }),
  .ZN({ S18251 })
);
NAND3_X1 #() 
NAND3_X1_2735_ (
  .A1({ S18243 }),
  .A2({ S18251 }),
  .A3({ S25957[150] }),
  .ZN({ S18252 })
);
INV_X1 #() 
INV_X1_794_ (
  .A({ S18221 }),
  .ZN({ S18254 })
);
INV_X1 #() 
INV_X1_795_ (
  .A({ S18171 }),
  .ZN({ S18255 })
);
NAND2_X1 #() 
NAND2_X1_2562_ (
  .A1({ S18180 }),
  .A2({ S18188 }),
  .ZN({ S18256 })
);
NOR2_X1 #() 
NOR2_X1_622_ (
  .A1({ S18255 }),
  .A2({ S18256 }),
  .ZN({ S18257 })
);
OAI21_X1 #() 
OAI21_X1_1353_ (
  .A({ S18178 }),
  .B1({ S18257 }),
  .B2({ S44 }),
  .ZN({ S18258 })
);
OAI211_X1 #() 
OAI211_X1_925_ (
  .A({ S14027 }),
  .B({ S14070 }),
  .C1({ S14136 }),
  .C2({ S14135 }),
  .ZN({ S18259 })
);
NAND2_X1 #() 
NAND2_X1_2563_ (
  .A1({ S18259 }),
  .A2({ S18188 }),
  .ZN({ S18260 })
);
NAND2_X1 #() 
NAND2_X1_2564_ (
  .A1({ S44 }),
  .A2({ S18260 }),
  .ZN({ S18261 })
);
NAND3_X1 #() 
NAND3_X1_2736_ (
  .A1({ S18219 }),
  .A2({ S13895 }),
  .A3({ S13898 }),
  .ZN({ S18262 })
);
OAI211_X1 #() 
OAI211_X1_926_ (
  .A({ S25957[148] }),
  .B({ S18262 }),
  .C1({ S18261 }),
  .C2({ S18255 }),
  .ZN({ S18263 })
);
OAI211_X1 #() 
OAI211_X1_927_ (
  .A({ S18263 }),
  .B({ S25957[149] }),
  .C1({ S18254 }),
  .C2({ S18258 }),
  .ZN({ S18265 })
);
NOR2_X1 #() 
NOR2_X1_623_ (
  .A1({ S18182 }),
  .A2({ S18201 }),
  .ZN({ S18266 })
);
NAND2_X1 #() 
NAND2_X1_2565_ (
  .A1({ S18233 }),
  .A2({ S18170 }),
  .ZN({ S18267 })
);
INV_X1 #() 
INV_X1_796_ (
  .A({ S18267 }),
  .ZN({ S18268 })
);
NAND2_X1 #() 
NAND2_X1_2566_ (
  .A1({ S18268 }),
  .A2({ S25957[147] }),
  .ZN({ S18269 })
);
NAND2_X1 #() 
NAND2_X1_2567_ (
  .A1({ S18269 }),
  .A2({ S18178 }),
  .ZN({ S18270 })
);
NOR2_X1 #() 
NOR2_X1_624_ (
  .A1({ S18167 }),
  .A2({ S18161 }),
  .ZN({ S18271 })
);
NAND2_X1 #() 
NAND2_X1_2568_ (
  .A1({ S44 }),
  .A2({ S18234 }),
  .ZN({ S18272 })
);
OAI211_X1 #() 
OAI211_X1_928_ (
  .A({ S18272 }),
  .B({ S25957[148] }),
  .C1({ S44 }),
  .C2({ S18271 }),
  .ZN({ S18273 })
);
OAI211_X1 #() 
OAI211_X1_929_ (
  .A({ S18273 }),
  .B({ S13688 }),
  .C1({ S18266 }),
  .C2({ S18270 }),
  .ZN({ S18274 })
);
NAND3_X1 #() 
NAND3_X1_2737_ (
  .A1({ S18265 }),
  .A2({ S18274 }),
  .A3({ S18185 }),
  .ZN({ S18276 })
);
AND3_X1 #() 
AND3_X1_111_ (
  .A1({ S18252 }),
  .A2({ S18276 }),
  .A3({ S25957[151] }),
  .ZN({ S18277 })
);
NOR2_X1 #() 
NOR2_X1_625_ (
  .A1({ S18277 }),
  .A2({ S18228 }),
  .ZN({ S18278 })
);
XOR2_X1 #() 
XOR2_X1_57_ (
  .A({ S18278 }),
  .B({ S25957[248] }),
  .Z({ S25957[120] })
);
NAND2_X1 #() 
NAND2_X1_2569_ (
  .A1({ S18178 }),
  .A2({ S18173 }),
  .ZN({ S18279 })
);
NAND3_X1 #() 
NAND3_X1_2738_ (
  .A1({ S64 }),
  .A2({ S18160 }),
  .A3({ S25957[146] }),
  .ZN({ S18280 })
);
INV_X1 #() 
INV_X1_797_ (
  .A({ S18280 }),
  .ZN({ S18281 })
);
NAND2_X1 #() 
NAND2_X1_2570_ (
  .A1({ S18188 }),
  .A2({ S18167 }),
  .ZN({ S18282 })
);
NAND2_X1 #() 
NAND2_X1_2571_ (
  .A1({ S25957[147] }),
  .A2({ S18282 }),
  .ZN({ S18283 })
);
OAI221_X1 #() 
OAI221_X1_64_ (
  .A({ S25957[148] }),
  .B1({ S18268 }),
  .B2({ S25957[147] }),
  .C1({ S18283 }),
  .C2({ S18281 }),
  .ZN({ S18284 })
);
NAND2_X1 #() 
NAND2_X1_2572_ (
  .A1({ S25957[146] }),
  .A2({ S18170 }),
  .ZN({ S18286 })
);
INV_X1 #() 
INV_X1_798_ (
  .A({ S18286 }),
  .ZN({ S18287 })
);
NOR2_X1 #() 
NOR2_X1_626_ (
  .A1({ S44 }),
  .A2({ S18287 }),
  .ZN({ S18288 })
);
NOR2_X1 #() 
NOR2_X1_627_ (
  .A1({ S25957[148] }),
  .A2({ S63 }),
  .ZN({ S18289 })
);
NAND2_X1 #() 
NAND2_X1_2573_ (
  .A1({ S18288 }),
  .A2({ S18289 }),
  .ZN({ S18290 })
);
NAND3_X1 #() 
NAND3_X1_2739_ (
  .A1({ S18188 }),
  .A2({ S18167 }),
  .A3({ S18208 }),
  .ZN({ S18291 })
);
NAND2_X1 #() 
NAND2_X1_2574_ (
  .A1({ S44 }),
  .A2({ S18291 }),
  .ZN({ S18292 })
);
OAI211_X1 #() 
OAI211_X1_930_ (
  .A({ S18284 }),
  .B({ S18290 }),
  .C1({ S18292 }),
  .C2({ S18279 }),
  .ZN({ S18293 })
);
NAND2_X1 #() 
NAND2_X1_2575_ (
  .A1({ S18160 }),
  .A2({ S25957[146] }),
  .ZN({ S18294 })
);
INV_X1 #() 
INV_X1_799_ (
  .A({ S18294 }),
  .ZN({ S18295 })
);
NAND2_X1 #() 
NAND2_X1_2576_ (
  .A1({ S44 }),
  .A2({ S18295 }),
  .ZN({ S18297 })
);
INV_X1 #() 
INV_X1_800_ (
  .A({ S18297 }),
  .ZN({ S18298 })
);
NAND3_X1 #() 
NAND3_X1_2740_ (
  .A1({ S13895 }),
  .A2({ S18271 }),
  .A3({ S13898 }),
  .ZN({ S18299 })
);
NAND3_X1 #() 
NAND3_X1_2741_ (
  .A1({ S25957[148] }),
  .A2({ S13899 }),
  .A3({ S13900 }),
  .ZN({ S18300 })
);
NAND2_X1 #() 
NAND2_X1_2577_ (
  .A1({ S25957[148] }),
  .A2({ S18160 }),
  .ZN({ S18301 })
);
NAND2_X1 #() 
NAND2_X1_2578_ (
  .A1({ S18300 }),
  .A2({ S18301 }),
  .ZN({ S18302 })
);
NAND2_X1 #() 
NAND2_X1_2579_ (
  .A1({ S18302 }),
  .A2({ S18299 }),
  .ZN({ S18303 })
);
NAND2_X1 #() 
NAND2_X1_2580_ (
  .A1({ S18271 }),
  .A2({ S18170 }),
  .ZN({ S18304 })
);
INV_X1 #() 
INV_X1_801_ (
  .A({ S18304 }),
  .ZN({ S18305 })
);
OAI21_X1 #() 
OAI21_X1_1354_ (
  .A({ S18175 }),
  .B1({ S25957[147] }),
  .B2({ S18305 }),
  .ZN({ S18306 })
);
NAND2_X1 #() 
NAND2_X1_2581_ (
  .A1({ S18306 }),
  .A2({ S18178 }),
  .ZN({ S18308 })
);
OAI211_X1 #() 
OAI211_X1_931_ (
  .A({ S18308 }),
  .B({ S25957[149] }),
  .C1({ S18298 }),
  .C2({ S18303 }),
  .ZN({ S18309 })
);
OAI211_X1 #() 
OAI211_X1_932_ (
  .A({ S18309 }),
  .B({ S25957[150] }),
  .C1({ S25957[149] }),
  .C2({ S18293 }),
  .ZN({ S18310 })
);
NAND3_X1 #() 
NAND3_X1_2742_ (
  .A1({ S44 }),
  .A2({ S18180 }),
  .A3({ S18208 }),
  .ZN({ S18311 })
);
NAND2_X1 #() 
NAND2_X1_2582_ (
  .A1({ S18311 }),
  .A2({ S18283 }),
  .ZN({ S18312 })
);
NAND2_X1 #() 
NAND2_X1_2583_ (
  .A1({ S18312 }),
  .A2({ S18178 }),
  .ZN({ S18313 })
);
NOR3_X1 #() 
NOR3_X1_85_ (
  .A1({ S18244 }),
  .A2({ S44 }),
  .A3({ S18255 }),
  .ZN({ S18314 })
);
NAND2_X1 #() 
NAND2_X1_2584_ (
  .A1({ S44 }),
  .A2({ S18170 }),
  .ZN({ S18315 })
);
OAI21_X1 #() 
OAI21_X1_1355_ (
  .A({ S25957[148] }),
  .B1({ S18315 }),
  .B2({ S18186 }),
  .ZN({ S18316 })
);
OR2_X1 #() 
OR2_X1_36_ (
  .A1({ S18316 }),
  .A2({ S18314 }),
  .ZN({ S18317 })
);
AOI21_X1 #() 
AOI21_X1_1453_ (
  .A({ S13688 }),
  .B1({ S18317 }),
  .B2({ S18313 }),
  .ZN({ S18319 })
);
INV_X1 #() 
INV_X1_802_ (
  .A({ S18239 }),
  .ZN({ S18320 })
);
NAND3_X1 #() 
NAND3_X1_2743_ (
  .A1({ S18320 }),
  .A2({ S44 }),
  .A3({ S18246 }),
  .ZN({ S18321 })
);
NOR2_X1 #() 
NOR2_X1_628_ (
  .A1({ S18295 }),
  .A2({ S18215 }),
  .ZN({ S18322 })
);
OAI211_X1 #() 
OAI211_X1_933_ (
  .A({ S18321 }),
  .B({ S18178 }),
  .C1({ S18322 }),
  .C2({ S44 }),
  .ZN({ S18323 })
);
NAND2_X1 #() 
NAND2_X1_2585_ (
  .A1({ S18190 }),
  .A2({ S44 }),
  .ZN({ S18324 })
);
INV_X1 #() 
INV_X1_803_ (
  .A({ S18180 }),
  .ZN({ S18325 })
);
NAND3_X1 #() 
NAND3_X1_2744_ (
  .A1({ S13895 }),
  .A2({ S18325 }),
  .A3({ S13898 }),
  .ZN({ S18326 })
);
NAND3_X1 #() 
NAND3_X1_2745_ (
  .A1({ S18324 }),
  .A2({ S25957[148] }),
  .A3({ S18326 }),
  .ZN({ S18327 })
);
AND3_X1 #() 
AND3_X1_112_ (
  .A1({ S18323 }),
  .A2({ S18327 }),
  .A3({ S13688 }),
  .ZN({ S18328 })
);
OAI21_X1 #() 
OAI21_X1_1356_ (
  .A({ S18185 }),
  .B1({ S18319 }),
  .B2({ S18328 }),
  .ZN({ S18330 })
);
NAND3_X1 #() 
NAND3_X1_2746_ (
  .A1({ S18330 }),
  .A2({ S18310 }),
  .A3({ S25957[151] }),
  .ZN({ S18331 })
);
INV_X1 #() 
INV_X1_804_ (
  .A({ S18172 }),
  .ZN({ S18332 })
);
NAND2_X1 #() 
NAND2_X1_2586_ (
  .A1({ S44 }),
  .A2({ S18205 }),
  .ZN({ S18333 })
);
NOR2_X1 #() 
NOR2_X1_629_ (
  .A1({ S18333 }),
  .A2({ S18332 }),
  .ZN({ S18334 })
);
NAND2_X1 #() 
NAND2_X1_2587_ (
  .A1({ S18193 }),
  .A2({ S44 }),
  .ZN({ S18335 })
);
NAND3_X1 #() 
NAND3_X1_2747_ (
  .A1({ S18245 }),
  .A2({ S18335 }),
  .A3({ S18178 }),
  .ZN({ S18336 })
);
OAI211_X1 #() 
OAI211_X1_934_ (
  .A({ S18336 }),
  .B({ S13688 }),
  .C1({ S18177 }),
  .C2({ S18334 }),
  .ZN({ S18337 })
);
INV_X1 #() 
INV_X1_805_ (
  .A({ S18208 }),
  .ZN({ S18338 })
);
NAND2_X1 #() 
NAND2_X1_2588_ (
  .A1({ S18188 }),
  .A2({ S18173 }),
  .ZN({ S18339 })
);
NOR3_X1 #() 
NOR3_X1_86_ (
  .A1({ S44 }),
  .A2({ S18338 }),
  .A3({ S18339 }),
  .ZN({ S18341 })
);
NOR2_X1 #() 
NOR2_X1_630_ (
  .A1({ S18179 }),
  .A2({ S25957[144] }),
  .ZN({ S18342 })
);
OAI211_X1 #() 
OAI211_X1_935_ (
  .A({ S13899 }),
  .B({ S13900 }),
  .C1({ S25957[146] }),
  .C2({ S18170 }),
  .ZN({ S18343 })
);
OAI21_X1 #() 
OAI21_X1_1357_ (
  .A({ S25957[148] }),
  .B1({ S18343 }),
  .B2({ S18342 }),
  .ZN({ S18344 })
);
INV_X1 #() 
INV_X1_806_ (
  .A({ S18173 }),
  .ZN({ S18345 })
);
AOI21_X1 #() 
AOI21_X1_1454_ (
  .A({ S18345 }),
  .B1({ S18182 }),
  .B2({ S18161 }),
  .ZN({ S18346 })
);
AOI21_X1 #() 
AOI21_X1_1455_ (
  .A({ S13688 }),
  .B1({ S18346 }),
  .B2({ S18178 }),
  .ZN({ S18347 })
);
OAI21_X1 #() 
OAI21_X1_1358_ (
  .A({ S18347 }),
  .B1({ S18341 }),
  .B2({ S18344 }),
  .ZN({ S18348 })
);
AND2_X1 #() 
AND2_X1_168_ (
  .A1({ S18348 }),
  .A2({ S18337 }),
  .ZN({ S18349 })
);
NAND2_X1 #() 
NAND2_X1_2589_ (
  .A1({ S25957[147] }),
  .A2({ S18259 }),
  .ZN({ S18350 })
);
NAND4_X1 #() 
NAND4_X1_329_ (
  .A1({ S18172 }),
  .A2({ S18222 }),
  .A3({ S13899 }),
  .A4({ S13900 }),
  .ZN({ S18352 })
);
OAI21_X1 #() 
OAI21_X1_1359_ (
  .A({ S18352 }),
  .B1({ S25957[149] }),
  .B2({ S18350 }),
  .ZN({ S18353 })
);
NAND2_X1 #() 
NAND2_X1_2590_ (
  .A1({ S18353 }),
  .A2({ S18178 }),
  .ZN({ S18354 })
);
INV_X1 #() 
INV_X1_807_ (
  .A({ S18256 }),
  .ZN({ S18355 })
);
NAND2_X1 #() 
NAND2_X1_2591_ (
  .A1({ S18355 }),
  .A2({ S25957[147] }),
  .ZN({ S18356 })
);
NAND3_X1 #() 
NAND3_X1_2748_ (
  .A1({ S44 }),
  .A2({ S18259 }),
  .A3({ S18286 }),
  .ZN({ S18357 })
);
NAND3_X1 #() 
NAND3_X1_2749_ (
  .A1({ S18357 }),
  .A2({ S18356 }),
  .A3({ S13688 }),
  .ZN({ S18358 })
);
NAND3_X1 #() 
NAND3_X1_2750_ (
  .A1({ S44 }),
  .A2({ S18170 }),
  .A3({ S18180 }),
  .ZN({ S18359 })
);
NAND2_X1 #() 
NAND2_X1_2592_ (
  .A1({ S18233 }),
  .A2({ S18188 }),
  .ZN({ S18360 })
);
NAND2_X1 #() 
NAND2_X1_2593_ (
  .A1({ S18360 }),
  .A2({ S18286 }),
  .ZN({ S18361 })
);
OAI211_X1 #() 
OAI211_X1_936_ (
  .A({ S25957[149] }),
  .B({ S18359 }),
  .C1({ S44 }),
  .C2({ S18361 }),
  .ZN({ S18363 })
);
AND2_X1 #() 
AND2_X1_169_ (
  .A1({ S18363 }),
  .A2({ S18358 }),
  .ZN({ S18364 })
);
OAI211_X1 #() 
OAI211_X1_937_ (
  .A({ S18185 }),
  .B({ S18354 }),
  .C1({ S18364 }),
  .C2({ S18178 }),
  .ZN({ S18365 })
);
OAI211_X1 #() 
OAI211_X1_938_ (
  .A({ S13526 }),
  .B({ S18365 }),
  .C1({ S18349 }),
  .C2({ S18185 }),
  .ZN({ S18366 })
);
NAND2_X1 #() 
NAND2_X1_2594_ (
  .A1({ S18366 }),
  .A2({ S18331 }),
  .ZN({ S18367 })
);
XNOR2_X1 #() 
XNOR2_X1_135_ (
  .A({ S18367 }),
  .B({ S25957[249] }),
  .ZN({ S25957[121] })
);
NAND2_X1 #() 
NAND2_X1_2595_ (
  .A1({ S25957[147] }),
  .A2({ S25957[146] }),
  .ZN({ S18368 })
);
NAND2_X1 #() 
NAND2_X1_2596_ (
  .A1({ S18368 }),
  .A2({ S18259 }),
  .ZN({ S18369 })
);
AOI21_X1 #() 
AOI21_X1_1456_ (
  .A({ S25957[148] }),
  .B1({ S25957[147] }),
  .B2({ S18338 }),
  .ZN({ S18370 })
);
NAND2_X1 #() 
NAND2_X1_2597_ (
  .A1({ S18369 }),
  .A2({ S18370 }),
  .ZN({ S18371 })
);
NOR2_X1 #() 
NOR2_X1_631_ (
  .A1({ S18160 }),
  .A2({ S25957[146] }),
  .ZN({ S18373 })
);
NOR2_X1 #() 
NOR2_X1_632_ (
  .A1({ S18207 }),
  .A2({ S18373 }),
  .ZN({ S18374 })
);
OAI21_X1 #() 
OAI21_X1_1360_ (
  .A({ S18161 }),
  .B1({ S25957[146] }),
  .B2({ S18170 }),
  .ZN({ S18375 })
);
NAND2_X1 #() 
NAND2_X1_2598_ (
  .A1({ S44 }),
  .A2({ S18375 }),
  .ZN({ S18376 })
);
NAND2_X1 #() 
NAND2_X1_2599_ (
  .A1({ S18376 }),
  .A2({ S25957[148] }),
  .ZN({ S18377 })
);
OAI211_X1 #() 
OAI211_X1_939_ (
  .A({ S18371 }),
  .B({ S13688 }),
  .C1({ S18374 }),
  .C2({ S18377 }),
  .ZN({ S18378 })
);
NAND2_X1 #() 
NAND2_X1_2600_ (
  .A1({ S25957[147] }),
  .A2({ S18291 }),
  .ZN({ S18379 })
);
NAND3_X1 #() 
NAND3_X1_2751_ (
  .A1({ S13899 }),
  .A2({ S13900 }),
  .A3({ S25957[145] }),
  .ZN({ S18380 })
);
OAI221_X1 #() 
OAI221_X1_65_ (
  .A({ S18178 }),
  .B1({ S18380 }),
  .B2({ S18167 }),
  .C1({ S18379 }),
  .C2({ S18305 }),
  .ZN({ S18381 })
);
NAND3_X1 #() 
NAND3_X1_2752_ (
  .A1({ S25957[147] }),
  .A2({ S18259 }),
  .A3({ S18286 }),
  .ZN({ S18382 })
);
NAND3_X1 #() 
NAND3_X1_2753_ (
  .A1({ S18235 }),
  .A2({ S18382 }),
  .A3({ S25957[148] }),
  .ZN({ S18384 })
);
NAND3_X1 #() 
NAND3_X1_2754_ (
  .A1({ S18381 }),
  .A2({ S25957[149] }),
  .A3({ S18384 }),
  .ZN({ S18385 })
);
NAND3_X1 #() 
NAND3_X1_2755_ (
  .A1({ S18378 }),
  .A2({ S18385 }),
  .A3({ S25957[150] }),
  .ZN({ S18386 })
);
NAND2_X1 #() 
NAND2_X1_2601_ (
  .A1({ S25957[147] }),
  .A2({ S18206 }),
  .ZN({ S18387 })
);
NAND2_X1 #() 
NAND2_X1_2602_ (
  .A1({ S64 }),
  .A2({ S25957[146] }),
  .ZN({ S18388 })
);
NAND3_X1 #() 
NAND3_X1_2756_ (
  .A1({ S18388 }),
  .A2({ S13899 }),
  .A3({ S13900 }),
  .ZN({ S18389 })
);
OAI211_X1 #() 
OAI211_X1_940_ (
  .A({ S18178 }),
  .B({ S18389 }),
  .C1({ S18387 }),
  .C2({ S18189 }),
  .ZN({ S18390 })
);
NAND2_X1 #() 
NAND2_X1_2603_ (
  .A1({ S18233 }),
  .A2({ S18259 }),
  .ZN({ S18391 })
);
NAND3_X1 #() 
NAND3_X1_2757_ (
  .A1({ S44 }),
  .A2({ S25957[144] }),
  .A3({ S18391 }),
  .ZN({ S18392 })
);
OAI211_X1 #() 
OAI211_X1_941_ (
  .A({ S18302 }),
  .B({ S18392 }),
  .C1({ S18368 }),
  .C2({ S18170 }),
  .ZN({ S18393 })
);
NAND3_X1 #() 
NAND3_X1_2758_ (
  .A1({ S18393 }),
  .A2({ S18390 }),
  .A3({ S25957[149] }),
  .ZN({ S18395 })
);
OAI211_X1 #() 
OAI211_X1_942_ (
  .A({ S18299 }),
  .B({ S18178 }),
  .C1({ S25957[147] }),
  .C2({ S18246 }),
  .ZN({ S18396 })
);
NAND2_X1 #() 
NAND2_X1_2604_ (
  .A1({ S44 }),
  .A2({ S18180 }),
  .ZN({ S18397 })
);
NAND2_X1 #() 
NAND2_X1_2605_ (
  .A1({ S25957[147] }),
  .A2({ S18360 }),
  .ZN({ S18398 })
);
NAND3_X1 #() 
NAND3_X1_2759_ (
  .A1({ S18397 }),
  .A2({ S18398 }),
  .A3({ S25957[148] }),
  .ZN({ S18399 })
);
NAND3_X1 #() 
NAND3_X1_2760_ (
  .A1({ S18399 }),
  .A2({ S13688 }),
  .A3({ S18396 }),
  .ZN({ S18400 })
);
AND2_X1 #() 
AND2_X1_170_ (
  .A1({ S18395 }),
  .A2({ S18400 }),
  .ZN({ S18401 })
);
OAI211_X1 #() 
OAI211_X1_943_ (
  .A({ S18386 }),
  .B({ S25957[151] }),
  .C1({ S18401 }),
  .C2({ S25957[150] }),
  .ZN({ S18402 })
);
NAND2_X1 #() 
NAND2_X1_2606_ (
  .A1({ S18246 }),
  .A2({ S18173 }),
  .ZN({ S18403 })
);
NOR2_X1 #() 
NOR2_X1_633_ (
  .A1({ S18403 }),
  .A2({ S44 }),
  .ZN({ S18404 })
);
NAND2_X1 #() 
NAND2_X1_2607_ (
  .A1({ S18180 }),
  .A2({ S18179 }),
  .ZN({ S18406 })
);
AOI21_X1 #() 
AOI21_X1_1457_ (
  .A({ S25957[147] }),
  .B1({ S25957[144] }),
  .B2({ S18406 }),
  .ZN({ S18407 })
);
OAI21_X1 #() 
OAI21_X1_1361_ (
  .A({ S25957[148] }),
  .B1({ S18404 }),
  .B2({ S18407 }),
  .ZN({ S18408 })
);
NAND2_X1 #() 
NAND2_X1_2608_ (
  .A1({ S18246 }),
  .A2({ S18206 }),
  .ZN({ S18409 })
);
NAND2_X1 #() 
NAND2_X1_2609_ (
  .A1({ S18409 }),
  .A2({ S44 }),
  .ZN({ S18410 })
);
NAND3_X1 #() 
NAND3_X1_2761_ (
  .A1({ S18410 }),
  .A2({ S18178 }),
  .A3({ S18398 }),
  .ZN({ S18411 })
);
NAND3_X1 #() 
NAND3_X1_2762_ (
  .A1({ S18408 }),
  .A2({ S13688 }),
  .A3({ S18411 }),
  .ZN({ S18412 })
);
NAND3_X1 #() 
NAND3_X1_2763_ (
  .A1({ S25957[147] }),
  .A2({ S18234 }),
  .A3({ S18210 }),
  .ZN({ S18413 })
);
OAI211_X1 #() 
OAI211_X1_944_ (
  .A({ S18413 }),
  .B({ S18178 }),
  .C1({ S18397 }),
  .C2({ S18170 }),
  .ZN({ S18414 })
);
NOR3_X1 #() 
NOR3_X1_87_ (
  .A1({ S18300 }),
  .A2({ S18373 }),
  .A3({ S18345 }),
  .ZN({ S18415 })
);
INV_X1 #() 
INV_X1_808_ (
  .A({ S18259 }),
  .ZN({ S18417 })
);
NOR3_X1 #() 
NOR3_X1_88_ (
  .A1({ S18387 }),
  .A2({ S18417 }),
  .A3({ S18178 }),
  .ZN({ S18418 })
);
NOR3_X1 #() 
NOR3_X1_89_ (
  .A1({ S18418 }),
  .A2({ S18415 }),
  .A3({ S13688 }),
  .ZN({ S18419 })
);
NAND2_X1 #() 
NAND2_X1_2610_ (
  .A1({ S18419 }),
  .A2({ S18414 }),
  .ZN({ S18420 })
);
NAND3_X1 #() 
NAND3_X1_2764_ (
  .A1({ S18420 }),
  .A2({ S25957[150] }),
  .A3({ S18412 }),
  .ZN({ S18421 })
);
NAND2_X1 #() 
NAND2_X1_2611_ (
  .A1({ S44 }),
  .A2({ S18210 }),
  .ZN({ S18422 })
);
AOI21_X1 #() 
AOI21_X1_1458_ (
  .A({ S18178 }),
  .B1({ S18288 }),
  .B2({ S18237 }),
  .ZN({ S18423 })
);
OAI21_X1 #() 
OAI21_X1_1362_ (
  .A({ S18423 }),
  .B1({ S18325 }),
  .B2({ S18422 }),
  .ZN({ S18424 })
);
NAND3_X1 #() 
NAND3_X1_2765_ (
  .A1({ S18380 }),
  .A2({ S18211 }),
  .A3({ S18294 }),
  .ZN({ S18425 })
);
NAND3_X1 #() 
NAND3_X1_2766_ (
  .A1({ S18425 }),
  .A2({ S18178 }),
  .A3({ S18182 }),
  .ZN({ S18426 })
);
NAND3_X1 #() 
NAND3_X1_2767_ (
  .A1({ S18424 }),
  .A2({ S25957[149] }),
  .A3({ S18426 }),
  .ZN({ S18428 })
);
NAND2_X1 #() 
NAND2_X1_2612_ (
  .A1({ S18171 }),
  .A2({ S18259 }),
  .ZN({ S18429 })
);
OAI21_X1 #() 
OAI21_X1_1363_ (
  .A({ S44 }),
  .B1({ S18429 }),
  .B2({ S18239 }),
  .ZN({ S18430 })
);
AOI21_X1 #() 
AOI21_X1_1459_ (
  .A({ S18178 }),
  .B1({ S25957[147] }),
  .B2({ S18360 }),
  .ZN({ S18431 })
);
AOI22_X1 #() 
AOI22_X1_316_ (
  .A1({ S18431 }),
  .A2({ S18430 }),
  .B1({ S18235 }),
  .B2({ S18178 }),
  .ZN({ S18432 })
);
NAND4_X1 #() 
NAND4_X1_330_ (
  .A1({ S25957[147] }),
  .A2({ S18320 }),
  .A3({ S18246 }),
  .A4({ S18178 }),
  .ZN({ S18433 })
);
NAND2_X1 #() 
NAND2_X1_2613_ (
  .A1({ S18433 }),
  .A2({ S13688 }),
  .ZN({ S18434 })
);
OAI211_X1 #() 
OAI211_X1_945_ (
  .A({ S18428 }),
  .B({ S18185 }),
  .C1({ S18432 }),
  .C2({ S18434 }),
  .ZN({ S18435 })
);
NAND3_X1 #() 
NAND3_X1_2768_ (
  .A1({ S18435 }),
  .A2({ S13526 }),
  .A3({ S18421 }),
  .ZN({ S18436 })
);
NAND2_X1 #() 
NAND2_X1_2614_ (
  .A1({ S18436 }),
  .A2({ S18402 }),
  .ZN({ S18437 })
);
XNOR2_X1 #() 
XNOR2_X1_136_ (
  .A({ S18437 }),
  .B({ S25957[250] }),
  .ZN({ S25957[122] })
);
OAI21_X1 #() 
OAI21_X1_1364_ (
  .A({ S44 }),
  .B1({ S18332 }),
  .B2({ S18215 }),
  .ZN({ S18439 })
);
NAND2_X1 #() 
NAND2_X1_2615_ (
  .A1({ S18409 }),
  .A2({ S25957[147] }),
  .ZN({ S18440 })
);
NAND3_X1 #() 
NAND3_X1_2769_ (
  .A1({ S18440 }),
  .A2({ S18178 }),
  .A3({ S18439 }),
  .ZN({ S18441 })
);
NOR2_X1 #() 
NOR2_X1_634_ (
  .A1({ S44 }),
  .A2({ S18201 }),
  .ZN({ S18442 })
);
NAND2_X1 #() 
NAND2_X1_2616_ (
  .A1({ S18280 }),
  .A2({ S18222 }),
  .ZN({ S18443 })
);
NOR2_X1 #() 
NOR2_X1_635_ (
  .A1({ S18443 }),
  .A2({ S25957[147] }),
  .ZN({ S18444 })
);
OAI21_X1 #() 
OAI21_X1_1365_ (
  .A({ S25957[148] }),
  .B1({ S18444 }),
  .B2({ S18442 }),
  .ZN({ S18445 })
);
AOI21_X1 #() 
AOI21_X1_1460_ (
  .A({ S18185 }),
  .B1({ S18445 }),
  .B2({ S18441 }),
  .ZN({ S18446 })
);
AOI21_X1 #() 
AOI21_X1_1461_ (
  .A({ S25957[148] }),
  .B1({ S18361 }),
  .B2({ S25957[147] }),
  .ZN({ S18447 })
);
OAI21_X1 #() 
OAI21_X1_1366_ (
  .A({ S18447 }),
  .B1({ S18244 }),
  .B2({ S18397 }),
  .ZN({ S18449 })
);
INV_X1 #() 
INV_X1_809_ (
  .A({ S18234 }),
  .ZN({ S18450 })
);
INV_X1 #() 
INV_X1_810_ (
  .A({ S18206 }),
  .ZN({ S18451 })
);
OAI22_X1 #() 
OAI22_X1_63_ (
  .A1({ S18182 }),
  .A2({ S18451 }),
  .B1({ S18450 }),
  .B2({ S18262 }),
  .ZN({ S18452 })
);
NAND2_X1 #() 
NAND2_X1_2617_ (
  .A1({ S18452 }),
  .A2({ S25957[148] }),
  .ZN({ S18453 })
);
AOI21_X1 #() 
AOI21_X1_1462_ (
  .A({ S25957[150] }),
  .B1({ S18453 }),
  .B2({ S18449 }),
  .ZN({ S18454 })
);
OAI21_X1 #() 
OAI21_X1_1367_ (
  .A({ S25957[149] }),
  .B1({ S18454 }),
  .B2({ S18446 }),
  .ZN({ S18455 })
);
NAND3_X1 #() 
NAND3_X1_2770_ (
  .A1({ S25957[147] }),
  .A2({ S18172 }),
  .A3({ S18174 }),
  .ZN({ S18456 })
);
OAI211_X1 #() 
OAI211_X1_946_ (
  .A({ S18456 }),
  .B({ S18178 }),
  .C1({ S25957[147] }),
  .C2({ S18339 }),
  .ZN({ S18457 })
);
NAND3_X1 #() 
NAND3_X1_2771_ (
  .A1({ S18357 }),
  .A2({ S25957[148] }),
  .A3({ S18379 }),
  .ZN({ S18458 })
);
NAND3_X1 #() 
NAND3_X1_2772_ (
  .A1({ S18185 }),
  .A2({ S18457 }),
  .A3({ S18458 }),
  .ZN({ S18460 })
);
INV_X1 #() 
INV_X1_811_ (
  .A({ S18229 }),
  .ZN({ S18461 })
);
NOR3_X1 #() 
NOR3_X1_90_ (
  .A1({ S18281 }),
  .A2({ S25957[147] }),
  .A3({ S18461 }),
  .ZN({ S18462 })
);
AOI21_X1 #() 
AOI21_X1_1463_ (
  .A({ S25957[148] }),
  .B1({ S25957[147] }),
  .B2({ S25957[146] }),
  .ZN({ S18463 })
);
NAND2_X1 #() 
NAND2_X1_2618_ (
  .A1({ S18463 }),
  .A2({ S18339 }),
  .ZN({ S18464 })
);
OAI211_X1 #() 
OAI211_X1_947_ (
  .A({ S25957[150] }),
  .B({ S18464 }),
  .C1({ S18303 }),
  .C2({ S18462 }),
  .ZN({ S18465 })
);
NAND2_X1 #() 
NAND2_X1_2619_ (
  .A1({ S18460 }),
  .A2({ S18465 }),
  .ZN({ S18466 })
);
NAND2_X1 #() 
NAND2_X1_2620_ (
  .A1({ S18466 }),
  .A2({ S13688 }),
  .ZN({ S18467 })
);
NAND3_X1 #() 
NAND3_X1_2773_ (
  .A1({ S18455 }),
  .A2({ S25957[151] }),
  .A3({ S18467 }),
  .ZN({ S18468 })
);
AOI21_X1 #() 
AOI21_X1_1464_ (
  .A({ S25957[148] }),
  .B1({ S18392 }),
  .B2({ S18232 }),
  .ZN({ S18469 })
);
OAI21_X1 #() 
OAI21_X1_1368_ (
  .A({ S13688 }),
  .B1({ S18469 }),
  .B2({ S18415 }),
  .ZN({ S18471 })
);
NAND3_X1 #() 
NAND3_X1_2774_ (
  .A1({ S18311 }),
  .A2({ S18269 }),
  .A3({ S18178 }),
  .ZN({ S18472 })
);
NAND4_X1 #() 
NAND4_X1_331_ (
  .A1({ S18206 }),
  .A2({ S13895 }),
  .A3({ S18171 }),
  .A4({ S13898 }),
  .ZN({ S18473 })
);
OAI21_X1 #() 
OAI21_X1_1369_ (
  .A({ S44 }),
  .B1({ S18244 }),
  .B2({ S18429 }),
  .ZN({ S18474 })
);
NAND3_X1 #() 
NAND3_X1_2775_ (
  .A1({ S18474 }),
  .A2({ S25957[148] }),
  .A3({ S18473 }),
  .ZN({ S18475 })
);
NAND3_X1 #() 
NAND3_X1_2776_ (
  .A1({ S18475 }),
  .A2({ S25957[149] }),
  .A3({ S18472 }),
  .ZN({ S18476 })
);
NAND3_X1 #() 
NAND3_X1_2777_ (
  .A1({ S18471 }),
  .A2({ S18476 }),
  .A3({ S25957[150] }),
  .ZN({ S18477 })
);
AOI21_X1 #() 
AOI21_X1_1465_ (
  .A({ S18178 }),
  .B1({ S18422 }),
  .B2({ S18262 }),
  .ZN({ S18478 })
);
OAI21_X1 #() 
OAI21_X1_1370_ (
  .A({ S44 }),
  .B1({ S18461 }),
  .B2({ S18287 }),
  .ZN({ S18479 })
);
AOI21_X1 #() 
AOI21_X1_1466_ (
  .A({ S25957[148] }),
  .B1({ S18479 }),
  .B2({ S18387 }),
  .ZN({ S18480 })
);
OAI21_X1 #() 
OAI21_X1_1371_ (
  .A({ S25957[149] }),
  .B1({ S18480 }),
  .B2({ S18478 }),
  .ZN({ S18482 })
);
OAI21_X1 #() 
OAI21_X1_1372_ (
  .A({ S44 }),
  .B1({ S18244 }),
  .B2({ S18255 }),
  .ZN({ S18483 })
);
NOR2_X1 #() 
NOR2_X1_636_ (
  .A1({ S18287 }),
  .A2({ S18373 }),
  .ZN({ S18484 })
);
NAND2_X1 #() 
NAND2_X1_2621_ (
  .A1({ S18484 }),
  .A2({ S25957[147] }),
  .ZN({ S18485 })
);
NAND3_X1 #() 
NAND3_X1_2778_ (
  .A1({ S18485 }),
  .A2({ S18483 }),
  .A3({ S18178 }),
  .ZN({ S18486 })
);
NAND4_X1 #() 
NAND4_X1_332_ (
  .A1({ S18222 }),
  .A2({ S13899 }),
  .A3({ S18233 }),
  .A4({ S13900 }),
  .ZN({ S18487 })
);
INV_X1 #() 
INV_X1_812_ (
  .A({ S18487 }),
  .ZN({ S18488 })
);
OAI21_X1 #() 
OAI21_X1_1373_ (
  .A({ S25957[148] }),
  .B1({ S18341 }),
  .B2({ S18488 }),
  .ZN({ S18489 })
);
NAND3_X1 #() 
NAND3_X1_2779_ (
  .A1({ S18489 }),
  .A2({ S18486 }),
  .A3({ S13688 }),
  .ZN({ S18490 })
);
NAND2_X1 #() 
NAND2_X1_2622_ (
  .A1({ S18490 }),
  .A2({ S18482 }),
  .ZN({ S18491 })
);
OAI211_X1 #() 
OAI211_X1_948_ (
  .A({ S18477 }),
  .B({ S13526 }),
  .C1({ S18491 }),
  .C2({ S25957[150] }),
  .ZN({ S18493 })
);
NAND2_X1 #() 
NAND2_X1_2623_ (
  .A1({ S18468 }),
  .A2({ S18493 }),
  .ZN({ S18494 })
);
XNOR2_X1 #() 
XNOR2_X1_137_ (
  .A({ S18494 }),
  .B({ S25957[251] }),
  .ZN({ S25957[123] })
);
NAND2_X1 #() 
NAND2_X1_2624_ (
  .A1({ S18238 }),
  .A2({ S18178 }),
  .ZN({ S18495 })
);
NAND3_X1 #() 
NAND3_X1_2780_ (
  .A1({ S18232 }),
  .A2({ S18261 }),
  .A3({ S25957[148] }),
  .ZN({ S18496 })
);
OAI21_X1 #() 
OAI21_X1_1374_ (
  .A({ S18496 }),
  .B1({ S18495 }),
  .B2({ S18442 }),
  .ZN({ S18497 })
);
NAND2_X1 #() 
NAND2_X1_2625_ (
  .A1({ S25957[147] }),
  .A2({ S18234 }),
  .ZN({ S18498 })
);
AOI21_X1 #() 
AOI21_X1_1467_ (
  .A({ S25957[148] }),
  .B1({ S44 }),
  .B2({ S18160 }),
  .ZN({ S18499 })
);
AND2_X1 #() 
AND2_X1_171_ (
  .A1({ S18499 }),
  .A2({ S18498 }),
  .ZN({ S18500 })
);
NOR2_X1 #() 
NOR2_X1_637_ (
  .A1({ S18320 }),
  .A2({ S25957[147] }),
  .ZN({ S18501 })
);
NAND3_X1 #() 
NAND3_X1_2781_ (
  .A1({ S25957[148] }),
  .A2({ S18222 }),
  .A3({ S18233 }),
  .ZN({ S18503 })
);
AOI21_X1 #() 
AOI21_X1_1468_ (
  .A({ S18501 }),
  .B1({ S18300 }),
  .B2({ S18503 }),
  .ZN({ S18504 })
);
OAI21_X1 #() 
OAI21_X1_1375_ (
  .A({ S25957[149] }),
  .B1({ S18504 }),
  .B2({ S18500 }),
  .ZN({ S18505 })
);
OAI211_X1 #() 
OAI211_X1_949_ (
  .A({ S18505 }),
  .B({ S18185 }),
  .C1({ S25957[149] }),
  .C2({ S18497 }),
  .ZN({ S18506 })
);
AND2_X1 #() 
AND2_X1_172_ (
  .A1({ S18167 }),
  .A2({ S155 }),
  .ZN({ S18507 })
);
OAI211_X1 #() 
OAI211_X1_950_ (
  .A({ S18194 }),
  .B({ S18178 }),
  .C1({ S18292 }),
  .C2({ S18305 }),
  .ZN({ S18508 })
);
OAI211_X1 #() 
OAI211_X1_951_ (
  .A({ S18508 }),
  .B({ S25957[149] }),
  .C1({ S18178 }),
  .C2({ S18507 }),
  .ZN({ S18509 })
);
NAND2_X1 #() 
NAND2_X1_2626_ (
  .A1({ S18484 }),
  .A2({ S44 }),
  .ZN({ S18510 })
);
NAND2_X1 #() 
NAND2_X1_2627_ (
  .A1({ S18510 }),
  .A2({ S18463 }),
  .ZN({ S18511 })
);
NAND2_X1 #() 
NAND2_X1_2628_ (
  .A1({ S18286 }),
  .A2({ S18180 }),
  .ZN({ S18512 })
);
NAND3_X1 #() 
NAND3_X1_2782_ (
  .A1({ S44 }),
  .A2({ S18512 }),
  .A3({ S18233 }),
  .ZN({ S18514 })
);
NAND3_X1 #() 
NAND3_X1_2783_ (
  .A1({ S18514 }),
  .A2({ S18356 }),
  .A3({ S25957[148] }),
  .ZN({ S18515 })
);
NAND3_X1 #() 
NAND3_X1_2784_ (
  .A1({ S18511 }),
  .A2({ S13688 }),
  .A3({ S18515 }),
  .ZN({ S18516 })
);
NAND3_X1 #() 
NAND3_X1_2785_ (
  .A1({ S18509 }),
  .A2({ S18516 }),
  .A3({ S25957[150] }),
  .ZN({ S18517 })
);
NAND3_X1 #() 
NAND3_X1_2786_ (
  .A1({ S18506 }),
  .A2({ S13526 }),
  .A3({ S18517 }),
  .ZN({ S18518 })
);
NAND2_X1 #() 
NAND2_X1_2629_ (
  .A1({ S25957[148] }),
  .A2({ S18229 }),
  .ZN({ S18519 })
);
OAI21_X1 #() 
OAI21_X1_1376_ (
  .A({ S18359 }),
  .B1({ S18350 }),
  .B2({ S18345 }),
  .ZN({ S18520 })
);
OAI221_X1 #() 
OAI221_X1_66_ (
  .A({ S25957[149] }),
  .B1({ S18254 }),
  .B2({ S18519 }),
  .C1({ S18520 }),
  .C2({ S25957[148] }),
  .ZN({ S18521 })
);
NAND3_X1 #() 
NAND3_X1_2787_ (
  .A1({ S25957[147] }),
  .A2({ S18180 }),
  .A3({ S18208 }),
  .ZN({ S18522 })
);
NAND3_X1 #() 
NAND3_X1_2788_ (
  .A1({ S18357 }),
  .A2({ S18522 }),
  .A3({ S18178 }),
  .ZN({ S18523 })
);
NAND2_X1 #() 
NAND2_X1_2630_ (
  .A1({ S44 }),
  .A2({ S18188 }),
  .ZN({ S18525 })
);
OAI22_X1 #() 
OAI22_X1_64_ (
  .A1({ S18525 }),
  .A2({ S18417 }),
  .B1({ S44 }),
  .B2({ S18375 }),
  .ZN({ S18526 })
);
OAI211_X1 #() 
OAI211_X1_952_ (
  .A({ S18523 }),
  .B({ S13688 }),
  .C1({ S18526 }),
  .C2({ S18178 }),
  .ZN({ S18527 })
);
NAND3_X1 #() 
NAND3_X1_2789_ (
  .A1({ S18521 }),
  .A2({ S25957[150] }),
  .A3({ S18527 }),
  .ZN({ S18528 })
);
NAND4_X1 #() 
NAND4_X1_333_ (
  .A1({ S13895 }),
  .A2({ S13898 }),
  .A3({ S18179 }),
  .A4({ S18180 }),
  .ZN({ S18529 })
);
OAI211_X1 #() 
OAI211_X1_953_ (
  .A({ S18430 }),
  .B({ S25957[148] }),
  .C1({ S63 }),
  .C2({ S18529 }),
  .ZN({ S18530 })
);
OAI211_X1 #() 
OAI211_X1_954_ (
  .A({ S18321 }),
  .B({ S18178 }),
  .C1({ S44 }),
  .C2({ S18174 }),
  .ZN({ S18531 })
);
NAND3_X1 #() 
NAND3_X1_2790_ (
  .A1({ S18531 }),
  .A2({ S18530 }),
  .A3({ S13688 }),
  .ZN({ S18532 })
);
NOR2_X1 #() 
NOR2_X1_638_ (
  .A1({ S18322 }),
  .A2({ S25957[147] }),
  .ZN({ S18533 })
);
NAND3_X1 #() 
NAND3_X1_2791_ (
  .A1({ S25957[147] }),
  .A2({ S18246 }),
  .A3({ S18208 }),
  .ZN({ S18534 })
);
NAND3_X1 #() 
NAND3_X1_2792_ (
  .A1({ S18247 }),
  .A2({ S18534 }),
  .A3({ S25957[148] }),
  .ZN({ S18536 })
);
OAI211_X1 #() 
OAI211_X1_955_ (
  .A({ S18536 }),
  .B({ S25957[149] }),
  .C1({ S18533 }),
  .C2({ S18258 }),
  .ZN({ S18537 })
);
NAND3_X1 #() 
NAND3_X1_2793_ (
  .A1({ S18532 }),
  .A2({ S18537 }),
  .A3({ S18185 }),
  .ZN({ S18538 })
);
NAND3_X1 #() 
NAND3_X1_2794_ (
  .A1({ S18528 }),
  .A2({ S25957[151] }),
  .A3({ S18538 }),
  .ZN({ S18539 })
);
NAND2_X1 #() 
NAND2_X1_2631_ (
  .A1({ S18518 }),
  .A2({ S18539 }),
  .ZN({ S18540 })
);
XOR2_X1 #() 
XOR2_X1_58_ (
  .A({ S18540 }),
  .B({ S25957[252] }),
  .Z({ S25957[124] })
);
OAI221_X1 #() 
OAI221_X1_67_ (
  .A({ S25957[148] }),
  .B1({ S18529 }),
  .B2({ S18170 }),
  .C1({ S18182 }),
  .C2({ S63 }),
  .ZN({ S18541 })
);
OAI221_X1 #() 
OAI221_X1_68_ (
  .A({ S18178 }),
  .B1({ S25957[145] }),
  .B2({ S44 }),
  .C1({ S18525 }),
  .C2({ S18417 }),
  .ZN({ S18542 })
);
NAND3_X1 #() 
NAND3_X1_2795_ (
  .A1({ S18541 }),
  .A2({ S18542 }),
  .A3({ S25957[149] }),
  .ZN({ S18543 })
);
AOI21_X1 #() 
AOI21_X1_1469_ (
  .A({ S44 }),
  .B1({ S18205 }),
  .B2({ S18280 }),
  .ZN({ S18544 })
);
NAND3_X1 #() 
NAND3_X1_2796_ (
  .A1({ S18397 }),
  .A2({ S18315 }),
  .A3({ S18178 }),
  .ZN({ S18546 })
);
NAND3_X1 #() 
NAND3_X1_2797_ (
  .A1({ S18376 }),
  .A2({ S18498 }),
  .A3({ S25957[148] }),
  .ZN({ S18547 })
);
OAI211_X1 #() 
OAI211_X1_956_ (
  .A({ S18547 }),
  .B({ S13688 }),
  .C1({ S18546 }),
  .C2({ S18544 }),
  .ZN({ S18548 })
);
NAND3_X1 #() 
NAND3_X1_2798_ (
  .A1({ S18543 }),
  .A2({ S18548 }),
  .A3({ S18185 }),
  .ZN({ S18549 })
);
NAND3_X1 #() 
NAND3_X1_2799_ (
  .A1({ S25957[147] }),
  .A2({ S18246 }),
  .A3({ S18286 }),
  .ZN({ S18550 })
);
OAI21_X1 #() 
OAI21_X1_1377_ (
  .A({ S18550 }),
  .B1({ S25957[147] }),
  .B2({ S18257 }),
  .ZN({ S18551 })
);
NAND2_X1 #() 
NAND2_X1_2632_ (
  .A1({ S25957[147] }),
  .A2({ S18429 }),
  .ZN({ S18552 })
);
NAND3_X1 #() 
NAND3_X1_2800_ (
  .A1({ S18195 }),
  .A2({ S18240 }),
  .A3({ S18552 }),
  .ZN({ S18553 })
);
OAI211_X1 #() 
OAI211_X1_957_ (
  .A({ S18553 }),
  .B({ S25957[149] }),
  .C1({ S18551 }),
  .C2({ S18178 }),
  .ZN({ S18554 })
);
NAND2_X1 #() 
NAND2_X1_2633_ (
  .A1({ S18283 }),
  .A2({ S25957[148] }),
  .ZN({ S18555 })
);
NOR2_X1 #() 
NOR2_X1_639_ (
  .A1({ S25957[147] }),
  .A2({ S18210 }),
  .ZN({ S18557 })
);
NAND2_X1 #() 
NAND2_X1_2634_ (
  .A1({ S18473 }),
  .A2({ S18178 }),
  .ZN({ S18558 })
);
OAI221_X1 #() 
OAI221_X1_69_ (
  .A({ S13688 }),
  .B1({ S18558 }),
  .B2({ S18557 }),
  .C1({ S18555 }),
  .C2({ S18501 }),
  .ZN({ S18559 })
);
NAND3_X1 #() 
NAND3_X1_2801_ (
  .A1({ S18559 }),
  .A2({ S18554 }),
  .A3({ S25957[150] }),
  .ZN({ S18560 })
);
NAND3_X1 #() 
NAND3_X1_2802_ (
  .A1({ S18549 }),
  .A2({ S18560 }),
  .A3({ S25957[151] }),
  .ZN({ S18561 })
);
NAND3_X1 #() 
NAND3_X1_2803_ (
  .A1({ S18202 }),
  .A2({ S18191 }),
  .A3({ S18178 }),
  .ZN({ S18562 })
);
NAND2_X1 #() 
NAND2_X1_2635_ (
  .A1({ S18280 }),
  .A2({ S18282 }),
  .ZN({ S18563 })
);
OAI211_X1 #() 
OAI211_X1_958_ (
  .A({ S18487 }),
  .B({ S25957[148] }),
  .C1({ S18563 }),
  .C2({ S44 }),
  .ZN({ S18564 })
);
NAND3_X1 #() 
NAND3_X1_2804_ (
  .A1({ S18562 }),
  .A2({ S18564 }),
  .A3({ S25957[149] }),
  .ZN({ S18565 })
);
OAI21_X1 #() 
OAI21_X1_1378_ (
  .A({ S18194 }),
  .B1({ S18403 }),
  .B2({ S25957[147] }),
  .ZN({ S18566 })
);
OAI21_X1 #() 
OAI21_X1_1379_ (
  .A({ S44 }),
  .B1({ S18295 }),
  .B2({ S18373 }),
  .ZN({ S18568 })
);
NAND2_X1 #() 
NAND2_X1_2636_ (
  .A1({ S18300 }),
  .A2({ S18519 }),
  .ZN({ S18569 })
);
AOI22_X1 #() 
AOI22_X1_317_ (
  .A1({ S18566 }),
  .A2({ S18178 }),
  .B1({ S18568 }),
  .B2({ S18569 }),
  .ZN({ S18570 })
);
OAI21_X1 #() 
OAI21_X1_1380_ (
  .A({ S18565 }),
  .B1({ S18570 }),
  .B2({ S25957[149] }),
  .ZN({ S18571 })
);
OAI22_X1 #() 
OAI22_X1_65_ (
  .A1({ S18368 }),
  .A2({ S18170 }),
  .B1({ S25957[147] }),
  .B2({ S18361 }),
  .ZN({ S18572 })
);
NAND3_X1 #() 
NAND3_X1_2805_ (
  .A1({ S18249 }),
  .A2({ S18552 }),
  .A3({ S25957[148] }),
  .ZN({ S18573 })
);
OAI211_X1 #() 
OAI211_X1_959_ (
  .A({ S25957[149] }),
  .B({ S18573 }),
  .C1({ S18572 }),
  .C2({ S25957[148] }),
  .ZN({ S18574 })
);
OAI21_X1 #() 
OAI21_X1_1381_ (
  .A({ S18370 }),
  .B1({ S25957[147] }),
  .B2({ S18172 }),
  .ZN({ S18575 })
);
NAND3_X1 #() 
NAND3_X1_2806_ (
  .A1({ S25957[147] }),
  .A2({ S18229 }),
  .A3({ S18280 }),
  .ZN({ S18576 })
);
NAND3_X1 #() 
NAND3_X1_2807_ (
  .A1({ S18212 }),
  .A2({ S18576 }),
  .A3({ S25957[148] }),
  .ZN({ S18577 })
);
NAND3_X1 #() 
NAND3_X1_2808_ (
  .A1({ S18575 }),
  .A2({ S18577 }),
  .A3({ S13688 }),
  .ZN({ S18579 })
);
NAND3_X1 #() 
NAND3_X1_2809_ (
  .A1({ S18574 }),
  .A2({ S18185 }),
  .A3({ S18579 }),
  .ZN({ S18580 })
);
OAI211_X1 #() 
OAI211_X1_960_ (
  .A({ S13526 }),
  .B({ S18580 }),
  .C1({ S18571 }),
  .C2({ S18185 }),
  .ZN({ S18581 })
);
NAND2_X1 #() 
NAND2_X1_2637_ (
  .A1({ S18581 }),
  .A2({ S18561 }),
  .ZN({ S18582 })
);
XOR2_X1 #() 
XOR2_X1_59_ (
  .A({ S18582 }),
  .B({ S25957[253] }),
  .Z({ S25957[125] })
);
INV_X1 #() 
INV_X1_813_ (
  .A({ S25957[254] }),
  .ZN({ S18583 })
);
NAND4_X1 #() 
NAND4_X1_334_ (
  .A1({ S18291 }),
  .A2({ S18286 }),
  .A3({ S13900 }),
  .A4({ S13899 }),
  .ZN({ S18584 })
);
AOI21_X1 #() 
AOI21_X1_1470_ (
  .A({ S18178 }),
  .B1({ S18584 }),
  .B2({ S18473 }),
  .ZN({ S18585 })
);
NAND2_X1 #() 
NAND2_X1_2638_ (
  .A1({ S18388 }),
  .A2({ S18211 }),
  .ZN({ S18586 })
);
NAND2_X1 #() 
NAND2_X1_2639_ (
  .A1({ S18586 }),
  .A2({ S25957[147] }),
  .ZN({ S18587 })
);
AOI21_X1 #() 
AOI21_X1_1471_ (
  .A({ S25957[148] }),
  .B1({ S18587 }),
  .B2({ S18352 }),
  .ZN({ S18589 })
);
OAI21_X1 #() 
OAI21_X1_1382_ (
  .A({ S13688 }),
  .B1({ S18589 }),
  .B2({ S18585 }),
  .ZN({ S18590 })
);
NAND3_X1 #() 
NAND3_X1_2810_ (
  .A1({ S18207 }),
  .A2({ S18389 }),
  .A3({ S25957[148] }),
  .ZN({ S18591 })
);
NAND2_X1 #() 
NAND2_X1_2640_ (
  .A1({ S25957[147] }),
  .A2({ S18260 }),
  .ZN({ S18592 })
);
NAND3_X1 #() 
NAND3_X1_2811_ (
  .A1({ S18592 }),
  .A2({ S18178 }),
  .A3({ S18380 }),
  .ZN({ S18593 })
);
NAND3_X1 #() 
NAND3_X1_2812_ (
  .A1({ S18593 }),
  .A2({ S18591 }),
  .A3({ S25957[149] }),
  .ZN({ S18594 })
);
NAND3_X1 #() 
NAND3_X1_2813_ (
  .A1({ S18590 }),
  .A2({ S25957[150] }),
  .A3({ S18594 }),
  .ZN({ S18595 })
);
NAND4_X1 #() 
NAND4_X1_335_ (
  .A1({ S18406 }),
  .A2({ S13895 }),
  .A3({ S18160 }),
  .A4({ S13898 }),
  .ZN({ S18596 })
);
NAND4_X1 #() 
NAND4_X1_336_ (
  .A1({ S18210 }),
  .A2({ S18205 }),
  .A3({ S13900 }),
  .A4({ S13899 }),
  .ZN({ S18597 })
);
NAND3_X1 #() 
NAND3_X1_2814_ (
  .A1({ S18597 }),
  .A2({ S18596 }),
  .A3({ S18178 }),
  .ZN({ S18598 })
);
OAI211_X1 #() 
OAI211_X1_961_ (
  .A({ S25957[148] }),
  .B({ S18299 }),
  .C1({ S18563 }),
  .C2({ S25957[147] }),
  .ZN({ S18600 })
);
NAND3_X1 #() 
NAND3_X1_2815_ (
  .A1({ S18600 }),
  .A2({ S18598 }),
  .A3({ S25957[149] }),
  .ZN({ S18601 })
);
NAND4_X1 #() 
NAND4_X1_337_ (
  .A1({ S18267 }),
  .A2({ S18173 }),
  .A3({ S13898 }),
  .A4({ S13895 }),
  .ZN({ S18602 })
);
NAND3_X1 #() 
NAND3_X1_2816_ (
  .A1({ S18584 }),
  .A2({ S18602 }),
  .A3({ S18178 }),
  .ZN({ S18603 })
);
NAND3_X1 #() 
NAND3_X1_2817_ (
  .A1({ S13899 }),
  .A2({ S18229 }),
  .A3({ S13900 }),
  .ZN({ S18604 })
);
OAI211_X1 #() 
OAI211_X1_962_ (
  .A({ S25957[148] }),
  .B({ S18604 }),
  .C1({ S18355 }),
  .C2({ S44 }),
  .ZN({ S18605 })
);
NAND3_X1 #() 
NAND3_X1_2818_ (
  .A1({ S18603 }),
  .A2({ S13688 }),
  .A3({ S18605 }),
  .ZN({ S18606 })
);
NAND3_X1 #() 
NAND3_X1_2819_ (
  .A1({ S18601 }),
  .A2({ S18606 }),
  .A3({ S18185 }),
  .ZN({ S18607 })
);
NAND3_X1 #() 
NAND3_X1_2820_ (
  .A1({ S18595 }),
  .A2({ S25957[151] }),
  .A3({ S18607 }),
  .ZN({ S18608 })
);
NOR2_X1 #() 
NOR2_X1_640_ (
  .A1({ S18281 }),
  .A2({ S25957[147] }),
  .ZN({ S18609 })
);
NAND3_X1 #() 
NAND3_X1_2821_ (
  .A1({ S18168 }),
  .A2({ S13899 }),
  .A3({ S13900 }),
  .ZN({ S18611 })
);
NAND3_X1 #() 
NAND3_X1_2822_ (
  .A1({ S18611 }),
  .A2({ S25957[148] }),
  .A3({ S18326 }),
  .ZN({ S18612 })
);
OAI211_X1 #() 
OAI211_X1_963_ (
  .A({ S18612 }),
  .B({ S13688 }),
  .C1({ S18558 }),
  .C2({ S18609 }),
  .ZN({ S18613 })
);
NAND4_X1 #() 
NAND4_X1_338_ (
  .A1({ S13895 }),
  .A2({ S13898 }),
  .A3({ S18188 }),
  .A4({ S18173 }),
  .ZN({ S18614 })
);
OAI211_X1 #() 
OAI211_X1_964_ (
  .A({ S18614 }),
  .B({ S25957[148] }),
  .C1({ S25957[147] }),
  .C2({ S18193 }),
  .ZN({ S18615 })
);
INV_X1 #() 
INV_X1_814_ (
  .A({ S18360 }),
  .ZN({ S18616 })
);
OAI211_X1 #() 
OAI211_X1_965_ (
  .A({ S18616 }),
  .B({ S18178 }),
  .C1({ S44 }),
  .C2({ S18173 }),
  .ZN({ S18617 })
);
NAND3_X1 #() 
NAND3_X1_2823_ (
  .A1({ S18615 }),
  .A2({ S25957[149] }),
  .A3({ S18617 }),
  .ZN({ S18618 })
);
AOI21_X1 #() 
AOI21_X1_1472_ (
  .A({ S18185 }),
  .B1({ S18613 }),
  .B2({ S18618 }),
  .ZN({ S18619 })
);
AOI22_X1 #() 
AOI22_X1_318_ (
  .A1({ S18343 }),
  .A2({ S18262 }),
  .B1({ S18300 }),
  .B2({ S18301 }),
  .ZN({ S18620 })
);
AOI21_X1 #() 
AOI21_X1_1473_ (
  .A({ S25957[148] }),
  .B1({ S18487 }),
  .B2({ S18529 }),
  .ZN({ S18622 })
);
OAI21_X1 #() 
OAI21_X1_1383_ (
  .A({ S25957[149] }),
  .B1({ S18620 }),
  .B2({ S18622 }),
  .ZN({ S18623 })
);
NOR3_X1 #() 
NOR3_X1_91_ (
  .A1({ S44 }),
  .A2({ S18181 }),
  .A3({ S25957[148] }),
  .ZN({ S18624 })
);
AOI22_X1 #() 
AOI22_X1_319_ (
  .A1({ S18503 }),
  .A2({ S18300 }),
  .B1({ S44 }),
  .B2({ S18222 }),
  .ZN({ S18625 })
);
OAI21_X1 #() 
OAI21_X1_1384_ (
  .A({ S13688 }),
  .B1({ S18625 }),
  .B2({ S18624 }),
  .ZN({ S18626 })
);
AOI21_X1 #() 
AOI21_X1_1474_ (
  .A({ S25957[150] }),
  .B1({ S18623 }),
  .B2({ S18626 }),
  .ZN({ S18627 })
);
OAI21_X1 #() 
OAI21_X1_1385_ (
  .A({ S13526 }),
  .B1({ S18627 }),
  .B2({ S18619 }),
  .ZN({ S18628 })
);
NAND3_X1 #() 
NAND3_X1_2824_ (
  .A1({ S18628 }),
  .A2({ S18583 }),
  .A3({ S18608 }),
  .ZN({ S18629 })
);
NAND2_X1 #() 
NAND2_X1_2641_ (
  .A1({ S18613 }),
  .A2({ S18618 }),
  .ZN({ S18630 })
);
NAND2_X1 #() 
NAND2_X1_2642_ (
  .A1({ S18630 }),
  .A2({ S25957[150] }),
  .ZN({ S18631 })
);
NAND2_X1 #() 
NAND2_X1_2643_ (
  .A1({ S18343 }),
  .A2({ S18262 }),
  .ZN({ S18633 })
);
NAND2_X1 #() 
NAND2_X1_2644_ (
  .A1({ S18633 }),
  .A2({ S18302 }),
  .ZN({ S18634 })
);
INV_X1 #() 
INV_X1_815_ (
  .A({ S18622 }),
  .ZN({ S18635 })
);
NAND3_X1 #() 
NAND3_X1_2825_ (
  .A1({ S18635 }),
  .A2({ S18634 }),
  .A3({ S25957[149] }),
  .ZN({ S18636 })
);
NAND2_X1 #() 
NAND2_X1_2645_ (
  .A1({ S18503 }),
  .A2({ S18300 }),
  .ZN({ S18637 })
);
NAND3_X1 #() 
NAND3_X1_2826_ (
  .A1({ S18637 }),
  .A2({ S18343 }),
  .A3({ S18380 }),
  .ZN({ S18638 })
);
NAND3_X1 #() 
NAND3_X1_2827_ (
  .A1({ S18638 }),
  .A2({ S13688 }),
  .A3({ S18433 }),
  .ZN({ S18639 })
);
NAND3_X1 #() 
NAND3_X1_2828_ (
  .A1({ S18636 }),
  .A2({ S18639 }),
  .A3({ S18185 }),
  .ZN({ S18640 })
);
NAND3_X1 #() 
NAND3_X1_2829_ (
  .A1({ S18631 }),
  .A2({ S18640 }),
  .A3({ S13526 }),
  .ZN({ S18641 })
);
NAND2_X1 #() 
NAND2_X1_2646_ (
  .A1({ S18601 }),
  .A2({ S18606 }),
  .ZN({ S18642 })
);
NAND2_X1 #() 
NAND2_X1_2647_ (
  .A1({ S18642 }),
  .A2({ S18185 }),
  .ZN({ S18644 })
);
NAND2_X1 #() 
NAND2_X1_2648_ (
  .A1({ S18584 }),
  .A2({ S18473 }),
  .ZN({ S18645 })
);
NAND2_X1 #() 
NAND2_X1_2649_ (
  .A1({ S18645 }),
  .A2({ S25957[148] }),
  .ZN({ S18646 })
);
AOI22_X1 #() 
AOI22_X1_320_ (
  .A1({ S18391 }),
  .A2({ S25957[144] }),
  .B1({ S13895 }),
  .B2({ S13898 }),
  .ZN({ S18647 })
);
AOI22_X1 #() 
AOI22_X1_321_ (
  .A1({ S18211 }),
  .A2({ S18388 }),
  .B1({ S13899 }),
  .B2({ S13900 }),
  .ZN({ S18648 })
);
OAI21_X1 #() 
OAI21_X1_1386_ (
  .A({ S18178 }),
  .B1({ S18647 }),
  .B2({ S18648 }),
  .ZN({ S18649 })
);
AOI21_X1 #() 
AOI21_X1_1475_ (
  .A({ S25957[149] }),
  .B1({ S18646 }),
  .B2({ S18649 }),
  .ZN({ S18650 })
);
AND3_X1 #() 
AND3_X1_113_ (
  .A1({ S18593 }),
  .A2({ S18591 }),
  .A3({ S25957[149] }),
  .ZN({ S18651 })
);
OAI21_X1 #() 
OAI21_X1_1387_ (
  .A({ S25957[150] }),
  .B1({ S18650 }),
  .B2({ S18651 }),
  .ZN({ S18652 })
);
NAND3_X1 #() 
NAND3_X1_2830_ (
  .A1({ S18652 }),
  .A2({ S25957[151] }),
  .A3({ S18644 }),
  .ZN({ S18653 })
);
NAND3_X1 #() 
NAND3_X1_2831_ (
  .A1({ S18653 }),
  .A2({ S25957[254] }),
  .A3({ S18641 }),
  .ZN({ S18655 })
);
NAND2_X1 #() 
NAND2_X1_2650_ (
  .A1({ S18655 }),
  .A2({ S18629 }),
  .ZN({ S25957[126] })
);
AOI21_X1 #() 
AOI21_X1_1476_ (
  .A({ S18178 }),
  .B1({ S25957[147] }),
  .B2({ S18304 }),
  .ZN({ S18656 })
);
AND2_X1 #() 
AND2_X1_173_ (
  .A1({ S18474 }),
  .A2({ S18656 }),
  .ZN({ S18657 })
);
NAND2_X1 #() 
NAND2_X1_2651_ (
  .A1({ S25957[147] }),
  .A2({ S18294 }),
  .ZN({ S18658 })
);
AOI21_X1 #() 
AOI21_X1_1477_ (
  .A({ S25957[148] }),
  .B1({ S18658 }),
  .B2({ S18422 }),
  .ZN({ S18659 })
);
OAI21_X1 #() 
OAI21_X1_1388_ (
  .A({ S18185 }),
  .B1({ S18657 }),
  .B2({ S18659 }),
  .ZN({ S18660 })
);
AOI21_X1 #() 
AOI21_X1_1478_ (
  .A({ S44 }),
  .B1({ S18291 }),
  .B2({ S18294 }),
  .ZN({ S18661 })
);
NAND3_X1 #() 
NAND3_X1_2832_ (
  .A1({ S25957[147] }),
  .A2({ S18180 }),
  .A3({ S18173 }),
  .ZN({ S18662 })
);
NAND3_X1 #() 
NAND3_X1_2833_ (
  .A1({ S18662 }),
  .A2({ S18178 }),
  .A3({ S18352 }),
  .ZN({ S18663 })
);
NAND2_X1 #() 
NAND2_X1_2652_ (
  .A1({ S18483 }),
  .A2({ S25957[148] }),
  .ZN({ S18665 })
);
OAI211_X1 #() 
OAI211_X1_966_ (
  .A({ S25957[150] }),
  .B({ S18663 }),
  .C1({ S18665 }),
  .C2({ S18661 }),
  .ZN({ S18666 })
);
AOI21_X1 #() 
AOI21_X1_1479_ (
  .A({ S25957[151] }),
  .B1({ S18660 }),
  .B2({ S18666 }),
  .ZN({ S18667 })
);
AOI21_X1 #() 
AOI21_X1_1480_ (
  .A({ S18178 }),
  .B1({ S18525 }),
  .B2({ S18592 }),
  .ZN({ S18668 })
);
NOR2_X1 #() 
NOR2_X1_641_ (
  .A1({ S18262 }),
  .A2({ S18325 }),
  .ZN({ S18669 })
);
NOR2_X1 #() 
NOR2_X1_642_ (
  .A1({ S18495 }),
  .A2({ S18669 }),
  .ZN({ S18670 })
);
OAI21_X1 #() 
OAI21_X1_1389_ (
  .A({ S25957[150] }),
  .B1({ S18670 }),
  .B2({ S18668 }),
  .ZN({ S18671 })
);
OAI21_X1 #() 
OAI21_X1_1390_ (
  .A({ S44 }),
  .B1({ S18186 }),
  .B2({ S18255 }),
  .ZN({ S18672 })
);
AOI21_X1 #() 
AOI21_X1_1481_ (
  .A({ S18178 }),
  .B1({ S18672 }),
  .B2({ S18413 }),
  .ZN({ S18673 })
);
NAND3_X1 #() 
NAND3_X1_2834_ (
  .A1({ S44 }),
  .A2({ S18291 }),
  .A3({ S18206 }),
  .ZN({ S18674 })
);
AOI21_X1 #() 
AOI21_X1_1482_ (
  .A({ S25957[148] }),
  .B1({ S18674 }),
  .B2({ S18350 }),
  .ZN({ S18676 })
);
OAI21_X1 #() 
OAI21_X1_1391_ (
  .A({ S18185 }),
  .B1({ S18673 }),
  .B2({ S18676 }),
  .ZN({ S18677 })
);
AOI21_X1 #() 
AOI21_X1_1483_ (
  .A({ S13526 }),
  .B1({ S18671 }),
  .B2({ S18677 }),
  .ZN({ S18678 })
);
OAI21_X1 #() 
OAI21_X1_1392_ (
  .A({ S13688 }),
  .B1({ S18678 }),
  .B2({ S18667 }),
  .ZN({ S18679 })
);
NAND3_X1 #() 
NAND3_X1_2835_ (
  .A1({ S25957[147] }),
  .A2({ S18222 }),
  .A3({ S18280 }),
  .ZN({ S18680 })
);
NOR2_X1 #() 
NOR2_X1_643_ (
  .A1({ S18342 }),
  .A2({ S18373 }),
  .ZN({ S18681 })
);
NAND2_X1 #() 
NAND2_X1_2653_ (
  .A1({ S18681 }),
  .A2({ S44 }),
  .ZN({ S18682 })
);
NAND3_X1 #() 
NAND3_X1_2836_ (
  .A1({ S18682 }),
  .A2({ S18178 }),
  .A3({ S18680 }),
  .ZN({ S18683 })
);
NAND3_X1 #() 
NAND3_X1_2837_ (
  .A1({ S25957[147] }),
  .A2({ S18230 }),
  .A3({ S25957[148] }),
  .ZN({ S18684 })
);
NAND4_X1 #() 
NAND4_X1_339_ (
  .A1({ S44 }),
  .A2({ S25957[148] }),
  .A3({ S25957[145] }),
  .A4({ S18171 }),
  .ZN({ S18685 })
);
NAND3_X1 #() 
NAND3_X1_2838_ (
  .A1({ S18683 }),
  .A2({ S18684 }),
  .A3({ S18685 }),
  .ZN({ S18687 })
);
NAND2_X1 #() 
NAND2_X1_2654_ (
  .A1({ S18687 }),
  .A2({ S25957[150] }),
  .ZN({ S18688 })
);
NAND2_X1 #() 
NAND2_X1_2655_ (
  .A1({ S18333 }),
  .A2({ S18289 }),
  .ZN({ S18689 })
);
OAI211_X1 #() 
OAI211_X1_967_ (
  .A({ S18356 }),
  .B({ S25957[148] }),
  .C1({ S18345 }),
  .C2({ S18380 }),
  .ZN({ S18690 })
);
NAND3_X1 #() 
NAND3_X1_2839_ (
  .A1({ S18185 }),
  .A2({ S18690 }),
  .A3({ S18689 }),
  .ZN({ S18691 })
);
AOI21_X1 #() 
AOI21_X1_1484_ (
  .A({ S13526 }),
  .B1({ S18688 }),
  .B2({ S18691 }),
  .ZN({ S18692 })
);
OAI211_X1 #() 
OAI211_X1_968_ (
  .A({ S18522 }),
  .B({ S18178 }),
  .C1({ S18182 }),
  .C2({ S18391 }),
  .ZN({ S18693 })
);
OAI211_X1 #() 
OAI211_X1_969_ (
  .A({ S18315 }),
  .B({ S25957[148] }),
  .C1({ S44 }),
  .C2({ S18512 }),
  .ZN({ S18694 })
);
NAND3_X1 #() 
NAND3_X1_2840_ (
  .A1({ S18185 }),
  .A2({ S18693 }),
  .A3({ S18694 }),
  .ZN({ S18695 })
);
NOR2_X1 #() 
NOR2_X1_644_ (
  .A1({ S18681 }),
  .A2({ S44 }),
  .ZN({ S18696 })
);
NAND3_X1 #() 
NAND3_X1_2841_ (
  .A1({ S25957[147] }),
  .A2({ S18233 }),
  .A3({ S18222 }),
  .ZN({ S18698 })
);
NAND3_X1 #() 
NAND3_X1_2842_ (
  .A1({ S18698 }),
  .A2({ S18297 }),
  .A3({ S18178 }),
  .ZN({ S18699 })
);
OAI211_X1 #() 
OAI211_X1_970_ (
  .A({ S25957[150] }),
  .B({ S18699 }),
  .C1({ S18316 }),
  .C2({ S18696 }),
  .ZN({ S18700 })
);
AOI21_X1 #() 
AOI21_X1_1485_ (
  .A({ S25957[151] }),
  .B1({ S18700 }),
  .B2({ S18695 }),
  .ZN({ S18701 })
);
OAI21_X1 #() 
OAI21_X1_1393_ (
  .A({ S25957[149] }),
  .B1({ S18692 }),
  .B2({ S18701 }),
  .ZN({ S18702 })
);
NAND2_X1 #() 
NAND2_X1_2656_ (
  .A1({ S18702 }),
  .A2({ S18679 }),
  .ZN({ S18703 })
);
XNOR2_X1 #() 
XNOR2_X1_138_ (
  .A({ S18703 }),
  .B({ S25957[255] }),
  .ZN({ S25957[127] })
);
NAND3_X1 #() 
NAND3_X1_2843_ (
  .A1({ S16404 }),
  .A2({ S16455 }),
  .A3({ S25957[224] }),
  .ZN({ S18704 })
);
NAND3_X1 #() 
NAND3_X1_2844_ (
  .A1({ S16497 }),
  .A2({ S16336 }),
  .A3({ S16477 }),
  .ZN({ S18705 })
);
AOI21_X1 #() 
AOI21_X1_1486_ (
  .A({ S25957[192] }),
  .B1({ S18704 }),
  .B2({ S18705 }),
  .ZN({ S18706 })
);
INV_X1 #() 
INV_X1_816_ (
  .A({ S25957[192] }),
  .ZN({ S18708 })
);
AOI21_X1 #() 
AOI21_X1_1487_ (
  .A({ S18708 }),
  .B1({ S16456 }),
  .B2({ S16498 }),
  .ZN({ S18709 })
);
NOR2_X1 #() 
NOR2_X1_645_ (
  .A1({ S18706 }),
  .A2({ S18709 }),
  .ZN({ S25957[64] })
);
INV_X1 #() 
INV_X1_817_ (
  .A({ S25957[193] }),
  .ZN({ S18710 })
);
NAND3_X1 #() 
NAND3_X1_2845_ (
  .A1({ S16542 }),
  .A2({ S25957[225] }),
  .A3({ S16576 }),
  .ZN({ S18711 })
);
NAND3_X1 #() 
NAND3_X1_2846_ (
  .A1({ S16580 }),
  .A2({ S16579 }),
  .A3({ S16499 }),
  .ZN({ S18712 })
);
NAND3_X1 #() 
NAND3_X1_2847_ (
  .A1({ S18711 }),
  .A2({ S18712 }),
  .A3({ S18710 }),
  .ZN({ S18713 })
);
NAND3_X1 #() 
NAND3_X1_2848_ (
  .A1({ S16577 }),
  .A2({ S16581 }),
  .A3({ S25957[193] }),
  .ZN({ S18714 })
);
NAND2_X1 #() 
NAND2_X1_2657_ (
  .A1({ S18713 }),
  .A2({ S18714 }),
  .ZN({ S25957[65] })
);
NAND3_X1 #() 
NAND3_X1_2849_ (
  .A1({ S16644 }),
  .A2({ S16661 }),
  .A3({ S25957[194] }),
  .ZN({ S18715 })
);
NAND3_X1 #() 
NAND3_X1_2850_ (
  .A1({ S16643 }),
  .A2({ S16645 }),
  .A3({ S16612 }),
  .ZN({ S18717 })
);
NAND3_X1 #() 
NAND3_X1_2851_ (
  .A1({ S16656 }),
  .A2({ S16660 }),
  .A3({ S25957[226] }),
  .ZN({ S18718 })
);
NAND3_X1 #() 
NAND3_X1_2852_ (
  .A1({ S18717 }),
  .A2({ S18718 }),
  .A3({ S16299 }),
  .ZN({ S18719 })
);
NAND2_X1 #() 
NAND2_X1_2658_ (
  .A1({ S18715 }),
  .A2({ S18719 }),
  .ZN({ S25957[66] })
);
NAND3_X1 #() 
NAND3_X1_2853_ (
  .A1({ S16721 }),
  .A2({ S25957[195] }),
  .A3({ S16740 }),
  .ZN({ S18720 })
);
NAND3_X1 #() 
NAND3_X1_2854_ (
  .A1({ S16694 }),
  .A2({ S16720 }),
  .A3({ S25957[227] }),
  .ZN({ S18721 })
);
NAND3_X1 #() 
NAND3_X1_2855_ (
  .A1({ S16730 }),
  .A2({ S16739 }),
  .A3({ S16662 }),
  .ZN({ S18722 })
);
NAND3_X1 #() 
NAND3_X1_2856_ (
  .A1({ S18721 }),
  .A2({ S16300 }),
  .A3({ S18722 }),
  .ZN({ S18723 })
);
NAND2_X1 #() 
NAND2_X1_2659_ (
  .A1({ S18720 }),
  .A2({ S18723 }),
  .ZN({ S25957[67] })
);
NAND3_X1 #() 
NAND3_X1_2857_ (
  .A1({ S16795 }),
  .A2({ S16766 }),
  .A3({ S25957[324] }),
  .ZN({ S18724 })
);
NAND2_X1 #() 
NAND2_X1_2660_ (
  .A1({ S16751 }),
  .A2({ S25957[158] }),
  .ZN({ S18726 })
);
NOR2_X1 #() 
NOR2_X1_646_ (
  .A1({ S16757 }),
  .A2({ S25957[157] }),
  .ZN({ S18727 })
);
AOI21_X1 #() 
AOI21_X1_1488_ (
  .A({ S18727 }),
  .B1({ S16762 }),
  .B2({ S25957[157] }),
  .ZN({ S18728 })
);
OAI211_X1 #() 
OAI211_X1_971_ (
  .A({ S18726 }),
  .B({ S15640 }),
  .C1({ S18728 }),
  .C2({ S25957[158] }),
  .ZN({ S18729 })
);
OAI211_X1 #() 
OAI211_X1_972_ (
  .A({ S16781 }),
  .B({ S25957[159] }),
  .C1({ S16793 }),
  .C2({ S25957[158] }),
  .ZN({ S18730 })
);
NAND3_X1 #() 
NAND3_X1_2858_ (
  .A1({ S18729 }),
  .A2({ S15211 }),
  .A3({ S18730 }),
  .ZN({ S18731 })
);
NAND2_X1 #() 
NAND2_X1_2661_ (
  .A1({ S18731 }),
  .A2({ S18724 }),
  .ZN({ S18732 })
);
INV_X1 #() 
INV_X1_818_ (
  .A({ S18732 }),
  .ZN({ S25957[68] })
);
OAI211_X1 #() 
OAI211_X1_973_ (
  .A({ S16849 }),
  .B({ S25957[229] }),
  .C1({ S16825 }),
  .C2({ S16810 }),
  .ZN({ S18733 })
);
OAI21_X1 #() 
OAI21_X1_1394_ (
  .A({ S16285 }),
  .B1({ S16858 }),
  .B2({ S16859 }),
  .ZN({ S18734 })
);
AOI21_X1 #() 
AOI21_X1_1489_ (
  .A({ S25957[197] }),
  .B1({ S18734 }),
  .B2({ S18733 }),
  .ZN({ S18736 })
);
INV_X1 #() 
INV_X1_819_ (
  .A({ S25957[197] }),
  .ZN({ S18737 })
);
AOI21_X1 #() 
AOI21_X1_1490_ (
  .A({ S18737 }),
  .B1({ S16860 }),
  .B2({ S16850 }),
  .ZN({ S18738 })
);
NOR2_X1 #() 
NOR2_X1_647_ (
  .A1({ S18736 }),
  .A2({ S18738 }),
  .ZN({ S25957[69] })
);
AOI21_X1 #() 
AOI21_X1_1491_ (
  .A({ S25957[326] }),
  .B1({ S16881 }),
  .B2({ S16908 }),
  .ZN({ S18739 })
);
NAND3_X1 #() 
NAND3_X1_2859_ (
  .A1({ S16881 }),
  .A2({ S16908 }),
  .A3({ S25957[326] }),
  .ZN({ S18740 })
);
INV_X1 #() 
INV_X1_820_ (
  .A({ S18740 }),
  .ZN({ S18741 })
);
NOR2_X1 #() 
NOR2_X1_648_ (
  .A1({ S18741 }),
  .A2({ S18739 }),
  .ZN({ S25957[70] })
);
NOR2_X1 #() 
NOR2_X1_649_ (
  .A1({ S16953 }),
  .A2({ S16376 }),
  .ZN({ S18742 })
);
NOR2_X1 #() 
NOR2_X1_650_ (
  .A1({ S16956 }),
  .A2({ S16948 }),
  .ZN({ S18743 })
);
OAI21_X1 #() 
OAI21_X1_1395_ (
  .A({ S25957[158] }),
  .B1({ S18742 }),
  .B2({ S18743 }),
  .ZN({ S18745 })
);
OAI21_X1 #() 
OAI21_X1_1396_ (
  .A({ S16946 }),
  .B1({ S16941 }),
  .B2({ S16376 }),
  .ZN({ S18746 })
);
NAND2_X1 #() 
NAND2_X1_2662_ (
  .A1({ S18746 }),
  .A2({ S15729 }),
  .ZN({ S18747 })
);
NAND3_X1 #() 
NAND3_X1_2860_ (
  .A1({ S18747 }),
  .A2({ S18745 }),
  .A3({ S15640 }),
  .ZN({ S18748 })
);
OAI221_X1 #() 
OAI221_X1_70_ (
  .A({ S25957[158] }),
  .B1({ S16918 }),
  .B2({ S16920 }),
  .C1({ S16914 }),
  .C2({ S16376 }),
  .ZN({ S18749 })
);
OAI211_X1 #() 
OAI211_X1_974_ (
  .A({ S18749 }),
  .B({ S25957[159] }),
  .C1({ S25957[158] }),
  .C2({ S16933 }),
  .ZN({ S18750 })
);
AOI21_X1 #() 
AOI21_X1_1492_ (
  .A({ S16274 }),
  .B1({ S18748 }),
  .B2({ S18750 }),
  .ZN({ S18751 })
);
AOI21_X1 #() 
AOI21_X1_1493_ (
  .A({ S25957[327] }),
  .B1({ S16935 }),
  .B2({ S16958 }),
  .ZN({ S18752 })
);
NOR2_X1 #() 
NOR2_X1_651_ (
  .A1({ S18751 }),
  .A2({ S18752 }),
  .ZN({ S25957[71] })
);
XOR2_X1 #() 
XOR2_X1_60_ (
  .A({ S25957[104] }),
  .B({ S25957[200] }),
  .Z({ S25957[72] })
);
XNOR2_X1 #() 
XNOR2_X1_139_ (
  .A({ S25957[105] }),
  .B({ S16301 }),
  .ZN({ S25957[73] })
);
NAND3_X1 #() 
NAND3_X1_2861_ (
  .A1({ S17249 }),
  .A2({ S17218 }),
  .A3({ S25957[330] }),
  .ZN({ S18754 })
);
NAND2_X1 #() 
NAND2_X1_2663_ (
  .A1({ S17250 }),
  .A2({ S16302 }),
  .ZN({ S18755 })
);
NAND2_X1 #() 
NAND2_X1_2664_ (
  .A1({ S18755 }),
  .A2({ S18754 }),
  .ZN({ S18756 })
);
INV_X1 #() 
INV_X1_821_ (
  .A({ S18756 }),
  .ZN({ S25957[74] })
);
NAND3_X1 #() 
NAND3_X1_2862_ (
  .A1({ S17344 }),
  .A2({ S25957[203] }),
  .A3({ S17308 }),
  .ZN({ S18757 })
);
INV_X1 #() 
INV_X1_822_ (
  .A({ S25957[203] }),
  .ZN({ S18758 })
);
OAI211_X1 #() 
OAI211_X1_975_ (
  .A({ S17307 }),
  .B({ S25957[235] }),
  .C1({ S17282 }),
  .C2({ S16966 }),
  .ZN({ S18759 })
);
NAND3_X1 #() 
NAND3_X1_2863_ (
  .A1({ S17323 }),
  .A2({ S17343 }),
  .A3({ S17252 }),
  .ZN({ S18760 })
);
NAND3_X1 #() 
NAND3_X1_2864_ (
  .A1({ S18760 }),
  .A2({ S18758 }),
  .A3({ S18759 }),
  .ZN({ S18761 })
);
NAND2_X1 #() 
NAND2_X1_2665_ (
  .A1({ S18757 }),
  .A2({ S18761 }),
  .ZN({ S25957[75] })
);
XNOR2_X1 #() 
XNOR2_X1_140_ (
  .A({ S25957[108] }),
  .B({ S16304 }),
  .ZN({ S25957[76] })
);
XOR2_X1 #() 
XOR2_X1_61_ (
  .A({ S25957[109] }),
  .B({ S25957[205] }),
  .Z({ S25957[77] })
);
NAND3_X1 #() 
NAND3_X1_2865_ (
  .A1({ S17488 }),
  .A2({ S17507 }),
  .A3({ S25957[238] }),
  .ZN({ S18763 })
);
NAND3_X1 #() 
NAND3_X1_2866_ (
  .A1({ S17520 }),
  .A2({ S17512 }),
  .A3({ S17462 }),
  .ZN({ S18764 })
);
NAND3_X1 #() 
NAND3_X1_2867_ (
  .A1({ S18763 }),
  .A2({ S18764 }),
  .A3({ S14359 }),
  .ZN({ S18765 })
);
NAND3_X1 #() 
NAND3_X1_2868_ (
  .A1({ S17508 }),
  .A2({ S17521 }),
  .A3({ S25957[206] }),
  .ZN({ S18766 })
);
NAND2_X1 #() 
NAND2_X1_2666_ (
  .A1({ S18765 }),
  .A2({ S18766 }),
  .ZN({ S25957[78] })
);
NAND3_X1 #() 
NAND3_X1_2869_ (
  .A1({ S17130 }),
  .A2({ S17564 }),
  .A3({ S25957[132] }),
  .ZN({ S18767 })
);
NAND3_X1 #() 
NAND3_X1_2870_ (
  .A1({ S17562 }),
  .A2({ S17028 }),
  .A3({ S17377 }),
  .ZN({ S18768 })
);
AND2_X1 #() 
AND2_X1_174_ (
  .A1({ S18768 }),
  .A2({ S25957[133] }),
  .ZN({ S18770 })
);
NAND2_X1 #() 
NAND2_X1_2667_ (
  .A1({ S17553 }),
  .A2({ S17189 }),
  .ZN({ S18771 })
);
NAND2_X1 #() 
NAND2_X1_2668_ (
  .A1({ S17552 }),
  .A2({ S18771 }),
  .ZN({ S18772 })
);
AOI22_X1 #() 
AOI22_X1_322_ (
  .A1({ S18772 }),
  .A2({ S16967 }),
  .B1({ S18770 }),
  .B2({ S18767 }),
  .ZN({ S18773 })
);
NAND2_X1 #() 
NAND2_X1_2669_ (
  .A1({ S17549 }),
  .A2({ S17028 }),
  .ZN({ S18774 })
);
NAND3_X1 #() 
NAND3_X1_2871_ (
  .A1({ S18774 }),
  .A2({ S16967 }),
  .A3({ S17548 }),
  .ZN({ S18775 })
);
NAND3_X1 #() 
NAND3_X1_2872_ (
  .A1({ S17559 }),
  .A2({ S25957[133] }),
  .A3({ S17560 }),
  .ZN({ S18776 })
);
NAND3_X1 #() 
NAND3_X1_2873_ (
  .A1({ S18775 }),
  .A2({ S15041 }),
  .A3({ S18776 }),
  .ZN({ S18777 })
);
OAI211_X1 #() 
OAI211_X1_976_ (
  .A({ S16966 }),
  .B({ S18777 }),
  .C1({ S18773 }),
  .C2({ S15041 }),
  .ZN({ S18778 })
);
OAI21_X1 #() 
OAI21_X1_1397_ (
  .A({ S25957[134] }),
  .B1({ S17527 }),
  .B2({ S17533 }),
  .ZN({ S18779 })
);
OAI21_X1 #() 
OAI21_X1_1398_ (
  .A({ S17540 }),
  .B1({ S17536 }),
  .B2({ S17544 }),
  .ZN({ S18781 })
);
NAND2_X1 #() 
NAND2_X1_2670_ (
  .A1({ S18781 }),
  .A2({ S15041 }),
  .ZN({ S18782 })
);
NAND3_X1 #() 
NAND3_X1_2874_ (
  .A1({ S18782 }),
  .A2({ S18779 }),
  .A3({ S25957[135] }),
  .ZN({ S18783 })
);
AOI21_X1 #() 
AOI21_X1_1494_ (
  .A({ S16305 }),
  .B1({ S18783 }),
  .B2({ S18778 }),
  .ZN({ S18784 })
);
AOI21_X1 #() 
AOI21_X1_1495_ (
  .A({ S25957[335] }),
  .B1({ S17546 }),
  .B2({ S17569 }),
  .ZN({ S18785 })
);
NOR2_X1 #() 
NOR2_X1_652_ (
  .A1({ S18785 }),
  .A2({ S18784 }),
  .ZN({ S25957[79] })
);
NAND3_X1 #() 
NAND3_X1_2875_ (
  .A1({ S17717 }),
  .A2({ S25957[208] }),
  .A3({ S17690 }),
  .ZN({ S18786 })
);
NAND3_X1 #() 
NAND3_X1_2876_ (
  .A1({ S17689 }),
  .A2({ S17644 }),
  .A3({ S25957[240] }),
  .ZN({ S18787 })
);
OAI21_X1 #() 
OAI21_X1_1399_ (
  .A({ S17576 }),
  .B1({ S17708 }),
  .B2({ S17715 }),
  .ZN({ S18788 })
);
NAND3_X1 #() 
NAND3_X1_2877_ (
  .A1({ S18788 }),
  .A2({ S16308 }),
  .A3({ S18787 }),
  .ZN({ S18789 })
);
NAND2_X1 #() 
NAND2_X1_2671_ (
  .A1({ S18786 }),
  .A2({ S18789 }),
  .ZN({ S25957[80] })
);
NAND3_X1 #() 
NAND3_X1_2878_ (
  .A1({ S17818 }),
  .A2({ S17801 }),
  .A3({ S25957[209] }),
  .ZN({ S18791 })
);
NAND3_X1 #() 
NAND3_X1_2879_ (
  .A1({ S17762 }),
  .A2({ S17800 }),
  .A3({ S25957[241] }),
  .ZN({ S18792 })
);
NAND3_X1 #() 
NAND3_X1_2880_ (
  .A1({ S17817 }),
  .A2({ S17812 }),
  .A3({ S17718 }),
  .ZN({ S18793 })
);
NAND3_X1 #() 
NAND3_X1_2881_ (
  .A1({ S18793 }),
  .A2({ S18792 }),
  .A3({ S16310 }),
  .ZN({ S18794 })
);
NAND2_X1 #() 
NAND2_X1_2672_ (
  .A1({ S18791 }),
  .A2({ S18794 }),
  .ZN({ S25957[81] })
);
NAND3_X1 #() 
NAND3_X1_2882_ (
  .A1({ S17850 }),
  .A2({ S17886 }),
  .A3({ S25957[338] }),
  .ZN({ S18795 })
);
INV_X1 #() 
INV_X1_823_ (
  .A({ S18795 }),
  .ZN({ S18796 })
);
AOI21_X1 #() 
AOI21_X1_1496_ (
  .A({ S25957[338] }),
  .B1({ S17850 }),
  .B2({ S17886 }),
  .ZN({ S18797 })
);
NOR2_X1 #() 
NOR2_X1_653_ (
  .A1({ S18796 }),
  .A2({ S18797 }),
  .ZN({ S25957[82] })
);
NAND3_X1 #() 
NAND3_X1_2883_ (
  .A1({ S17919 }),
  .A2({ S25957[339] }),
  .A3({ S17949 }),
  .ZN({ S18799 })
);
INV_X1 #() 
INV_X1_824_ (
  .A({ S18799 }),
  .ZN({ S18800 })
);
AOI21_X1 #() 
AOI21_X1_1497_ (
  .A({ S25957[339] }),
  .B1({ S17919 }),
  .B2({ S17949 }),
  .ZN({ S18801 })
);
NOR2_X1 #() 
NOR2_X1_654_ (
  .A1({ S18800 }),
  .A2({ S18801 }),
  .ZN({ S25957[83] })
);
NAND3_X1 #() 
NAND3_X1_2884_ (
  .A1({ S18005 }),
  .A2({ S17979 }),
  .A3({ S16311 }),
  .ZN({ S18802 })
);
AOI21_X1 #() 
AOI21_X1_1498_ (
  .A({ S16311 }),
  .B1({ S18005 }),
  .B2({ S17979 }),
  .ZN({ S18803 })
);
INV_X1 #() 
INV_X1_825_ (
  .A({ S18803 }),
  .ZN({ S18804 })
);
NAND2_X1 #() 
NAND2_X1_2673_ (
  .A1({ S18804 }),
  .A2({ S18802 }),
  .ZN({ S25957[84] })
);
NAND3_X1 #() 
NAND3_X1_2885_ (
  .A1({ S18031 }),
  .A2({ S25957[341] }),
  .A3({ S18049 }),
  .ZN({ S18805 })
);
INV_X1 #() 
INV_X1_826_ (
  .A({ S18805 }),
  .ZN({ S18806 })
);
AOI21_X1 #() 
AOI21_X1_1499_ (
  .A({ S25957[341] }),
  .B1({ S18031 }),
  .B2({ S18049 }),
  .ZN({ S18808 })
);
NOR2_X1 #() 
NOR2_X1_655_ (
  .A1({ S18806 }),
  .A2({ S18808 }),
  .ZN({ S25957[85] })
);
XOR2_X1 #() 
XOR2_X1_62_ (
  .A({ S25957[118] }),
  .B({ S25957[214] }),
  .Z({ S25957[86] })
);
XNOR2_X1 #() 
XNOR2_X1_141_ (
  .A({ S25957[119] }),
  .B({ S13522 }),
  .ZN({ S25957[87] })
);
AND2_X1 #() 
AND2_X1_175_ (
  .A1({ S18226 }),
  .A2({ S18185 }),
  .ZN({ S18809 })
);
AOI22_X1 #() 
AOI22_X1_323_ (
  .A1({ S18809 }),
  .A2({ S18214 }),
  .B1({ S18199 }),
  .B2({ S18184 }),
  .ZN({ S18810 })
);
NAND3_X1 #() 
NAND3_X1_2886_ (
  .A1({ S18252 }),
  .A2({ S18276 }),
  .A3({ S25957[151] }),
  .ZN({ S18811 })
);
OAI211_X1 #() 
OAI211_X1_977_ (
  .A({ S16095 }),
  .B({ S18811 }),
  .C1({ S18810 }),
  .C2({ S25957[151] }),
  .ZN({ S18812 })
);
OAI21_X1 #() 
OAI21_X1_1400_ (
  .A({ S25957[344] }),
  .B1({ S18277 }),
  .B2({ S18228 }),
  .ZN({ S18813 })
);
NAND2_X1 #() 
NAND2_X1_2674_ (
  .A1({ S18813 }),
  .A2({ S18812 }),
  .ZN({ S25957[88] })
);
NAND3_X1 #() 
NAND3_X1_2887_ (
  .A1({ S18366 }),
  .A2({ S18331 }),
  .A3({ S16312 }),
  .ZN({ S18815 })
);
AOI21_X1 #() 
AOI21_X1_1500_ (
  .A({ S16312 }),
  .B1({ S18366 }),
  .B2({ S18331 }),
  .ZN({ S18816 })
);
INV_X1 #() 
INV_X1_827_ (
  .A({ S18816 }),
  .ZN({ S18817 })
);
NAND2_X1 #() 
NAND2_X1_2675_ (
  .A1({ S18817 }),
  .A2({ S18815 }),
  .ZN({ S25957[89] })
);
NAND3_X1 #() 
NAND3_X1_2888_ (
  .A1({ S18436 }),
  .A2({ S16244 }),
  .A3({ S18402 }),
  .ZN({ S18818 })
);
AOI21_X1 #() 
AOI21_X1_1501_ (
  .A({ S16244 }),
  .B1({ S18436 }),
  .B2({ S18402 }),
  .ZN({ S18819 })
);
INV_X1 #() 
INV_X1_828_ (
  .A({ S18819 }),
  .ZN({ S18820 })
);
NAND2_X1 #() 
NAND2_X1_2676_ (
  .A1({ S18820 }),
  .A2({ S18818 }),
  .ZN({ S25957[90] })
);
OAI211_X1 #() 
OAI211_X1_978_ (
  .A({ S18203 }),
  .B({ S25957[148] }),
  .C1({ S25957[147] }),
  .C2({ S18443 }),
  .ZN({ S18821 })
);
AOI22_X1 #() 
AOI22_X1_324_ (
  .A1({ S18169 }),
  .A2({ S18208 }),
  .B1({ S18409 }),
  .B2({ S25957[147] }),
  .ZN({ S18822 })
);
OAI211_X1 #() 
OAI211_X1_979_ (
  .A({ S25957[149] }),
  .B({ S18821 }),
  .C1({ S18822 }),
  .C2({ S25957[148] }),
  .ZN({ S18824 })
);
OAI211_X1 #() 
OAI211_X1_980_ (
  .A({ S18464 }),
  .B({ S13688 }),
  .C1({ S18303 }),
  .C2({ S18462 }),
  .ZN({ S18825 })
);
NAND3_X1 #() 
NAND3_X1_2889_ (
  .A1({ S18824 }),
  .A2({ S25957[150] }),
  .A3({ S18825 }),
  .ZN({ S18826 })
);
AOI21_X1 #() 
AOI21_X1_1502_ (
  .A({ S13688 }),
  .B1({ S18452 }),
  .B2({ S25957[148] }),
  .ZN({ S18827 })
);
AOI21_X1 #() 
AOI21_X1_1503_ (
  .A({ S25957[149] }),
  .B1({ S18457 }),
  .B2({ S18458 }),
  .ZN({ S18828 })
);
AOI21_X1 #() 
AOI21_X1_1504_ (
  .A({ S18828 }),
  .B1({ S18827 }),
  .B2({ S18449 }),
  .ZN({ S18829 })
);
OAI211_X1 #() 
OAI211_X1_981_ (
  .A({ S18826 }),
  .B({ S25957[151] }),
  .C1({ S18829 }),
  .C2({ S25957[150] }),
  .ZN({ S18830 })
);
OAI21_X1 #() 
OAI21_X1_1401_ (
  .A({ S18477 }),
  .B1({ S18491 }),
  .B2({ S25957[150] }),
  .ZN({ S18831 })
);
NAND2_X1 #() 
NAND2_X1_2677_ (
  .A1({ S18831 }),
  .A2({ S13526 }),
  .ZN({ S18832 })
);
AOI21_X1 #() 
AOI21_X1_1505_ (
  .A({ S15910 }),
  .B1({ S18832 }),
  .B2({ S18830 }),
  .ZN({ S18833 })
);
AOI21_X1 #() 
AOI21_X1_1506_ (
  .A({ S25957[347] }),
  .B1({ S18468 }),
  .B2({ S18493 }),
  .ZN({ S18835 })
);
NOR2_X1 #() 
NOR2_X1_656_ (
  .A1({ S18833 }),
  .A2({ S18835 }),
  .ZN({ S25957[91] })
);
NAND3_X1 #() 
NAND3_X1_2890_ (
  .A1({ S18518 }),
  .A2({ S25957[348] }),
  .A3({ S18539 }),
  .ZN({ S18836 })
);
NAND2_X1 #() 
NAND2_X1_2678_ (
  .A1({ S18540 }),
  .A2({ S16314 }),
  .ZN({ S18837 })
);
NAND2_X1 #() 
NAND2_X1_2679_ (
  .A1({ S18837 }),
  .A2({ S18836 }),
  .ZN({ S25957[92] })
);
NAND3_X1 #() 
NAND3_X1_2891_ (
  .A1({ S18581 }),
  .A2({ S18561 }),
  .A3({ S15818 }),
  .ZN({ S18838 })
);
NAND2_X1 #() 
NAND2_X1_2680_ (
  .A1({ S18582 }),
  .A2({ S25957[349] }),
  .ZN({ S18839 })
);
NAND2_X1 #() 
NAND2_X1_2681_ (
  .A1({ S18839 }),
  .A2({ S18838 }),
  .ZN({ S18840 })
);
INV_X1 #() 
INV_X1_829_ (
  .A({ S18840 }),
  .ZN({ S25957[93] })
);
NAND3_X1 #() 
NAND3_X1_2892_ (
  .A1({ S18655 }),
  .A2({ S25957[222] }),
  .A3({ S18629 }),
  .ZN({ S18841 })
);
INV_X1 #() 
INV_X1_830_ (
  .A({ S25957[222] }),
  .ZN({ S18843 })
);
NAND3_X1 #() 
NAND3_X1_2893_ (
  .A1({ S18653 }),
  .A2({ S18583 }),
  .A3({ S18641 }),
  .ZN({ S18844 })
);
NAND3_X1 #() 
NAND3_X1_2894_ (
  .A1({ S18628 }),
  .A2({ S25957[254] }),
  .A3({ S18608 }),
  .ZN({ S18845 })
);
NAND3_X1 #() 
NAND3_X1_2895_ (
  .A1({ S18844 }),
  .A2({ S18843 }),
  .A3({ S18845 }),
  .ZN({ S18846 })
);
NAND2_X1 #() 
NAND2_X1_2682_ (
  .A1({ S18841 }),
  .A2({ S18846 }),
  .ZN({ S25957[94] })
);
INV_X1 #() 
INV_X1_831_ (
  .A({ S18668 }),
  .ZN({ S18847 })
);
OAI21_X1 #() 
OAI21_X1_1402_ (
  .A({ S18847 }),
  .B1({ S18495 }),
  .B2({ S18669 }),
  .ZN({ S18848 })
);
NAND4_X1 #() 
NAND4_X1_340_ (
  .A1({ S18683 }),
  .A2({ S25957[149] }),
  .A3({ S18684 }),
  .A4({ S18685 }),
  .ZN({ S18849 })
);
OAI211_X1 #() 
OAI211_X1_982_ (
  .A({ S18849 }),
  .B({ S25957[150] }),
  .C1({ S18848 }),
  .C2({ S25957[149] }),
  .ZN({ S18850 })
);
OAI21_X1 #() 
OAI21_X1_1403_ (
  .A({ S13688 }),
  .B1({ S18673 }),
  .B2({ S18676 }),
  .ZN({ S18851 })
);
NAND3_X1 #() 
NAND3_X1_2896_ (
  .A1({ S18690 }),
  .A2({ S25957[149] }),
  .A3({ S18689 }),
  .ZN({ S18853 })
);
NAND2_X1 #() 
NAND2_X1_2683_ (
  .A1({ S18851 }),
  .A2({ S18853 }),
  .ZN({ S18854 })
);
NAND2_X1 #() 
NAND2_X1_2684_ (
  .A1({ S18854 }),
  .A2({ S18185 }),
  .ZN({ S18855 })
);
NAND3_X1 #() 
NAND3_X1_2897_ (
  .A1({ S18850 }),
  .A2({ S18855 }),
  .A3({ S25957[151] }),
  .ZN({ S18856 })
);
NOR2_X1 #() 
NOR2_X1_657_ (
  .A1({ S18343 }),
  .A2({ S18281 }),
  .ZN({ S18857 })
);
OAI21_X1 #() 
OAI21_X1_1404_ (
  .A({ S25957[148] }),
  .B1({ S18857 }),
  .B2({ S18661 }),
  .ZN({ S18858 })
);
NAND3_X1 #() 
NAND3_X1_2898_ (
  .A1({ S18382 }),
  .A2({ S18392 }),
  .A3({ S18178 }),
  .ZN({ S18859 })
);
NAND3_X1 #() 
NAND3_X1_2899_ (
  .A1({ S18858 }),
  .A2({ S13688 }),
  .A3({ S18859 }),
  .ZN({ S18860 })
);
OAI21_X1 #() 
OAI21_X1_1405_ (
  .A({ S18699 }),
  .B1({ S18316 }),
  .B2({ S18696 }),
  .ZN({ S18861 })
);
NAND2_X1 #() 
NAND2_X1_2685_ (
  .A1({ S18861 }),
  .A2({ S25957[149] }),
  .ZN({ S18862 })
);
NAND3_X1 #() 
NAND3_X1_2900_ (
  .A1({ S18862 }),
  .A2({ S25957[150] }),
  .A3({ S18860 }),
  .ZN({ S18864 })
);
AND3_X1 #() 
AND3_X1_114_ (
  .A1({ S18693 }),
  .A2({ S25957[149] }),
  .A3({ S18694 }),
  .ZN({ S18865 })
);
NAND2_X1 #() 
NAND2_X1_2686_ (
  .A1({ S18474 }),
  .A2({ S18656 }),
  .ZN({ S18866 })
);
NAND2_X1 #() 
NAND2_X1_2687_ (
  .A1({ S18658 }),
  .A2({ S18422 }),
  .ZN({ S18867 })
);
NAND2_X1 #() 
NAND2_X1_2688_ (
  .A1({ S18867 }),
  .A2({ S18178 }),
  .ZN({ S18868 })
);
AOI21_X1 #() 
AOI21_X1_1507_ (
  .A({ S25957[149] }),
  .B1({ S18868 }),
  .B2({ S18866 }),
  .ZN({ S18869 })
);
OAI21_X1 #() 
OAI21_X1_1406_ (
  .A({ S18185 }),
  .B1({ S18865 }),
  .B2({ S18869 }),
  .ZN({ S18870 })
);
NAND3_X1 #() 
NAND3_X1_2901_ (
  .A1({ S18870 }),
  .A2({ S18864 }),
  .A3({ S13526 }),
  .ZN({ S18871 })
);
NAND3_X1 #() 
NAND3_X1_2902_ (
  .A1({ S18856 }),
  .A2({ S18871 }),
  .A3({ S25957[351] }),
  .ZN({ S18872 })
);
INV_X1 #() 
INV_X1_832_ (
  .A({ S25957[351] }),
  .ZN({ S18873 })
);
NAND3_X1 #() 
NAND3_X1_2903_ (
  .A1({ S18702 }),
  .A2({ S18679 }),
  .A3({ S18873 }),
  .ZN({ S18875 })
);
NAND2_X1 #() 
NAND2_X1_2689_ (
  .A1({ S18875 }),
  .A2({ S18872 }),
  .ZN({ S25957[95] })
);
OAI21_X1 #() 
OAI21_X1_1407_ (
  .A({ S25957[160] }),
  .B1({ S18706 }),
  .B2({ S18709 }),
  .ZN({ S18876 })
);
INV_X1 #() 
INV_X1_833_ (
  .A({ S25957[160] }),
  .ZN({ S18877 })
);
NAND3_X1 #() 
NAND3_X1_2904_ (
  .A1({ S16456 }),
  .A2({ S16498 }),
  .A3({ S18708 }),
  .ZN({ S18878 })
);
NAND3_X1 #() 
NAND3_X1_2905_ (
  .A1({ S18704 }),
  .A2({ S18705 }),
  .A3({ S25957[192] }),
  .ZN({ S18879 })
);
NAND3_X1 #() 
NAND3_X1_2906_ (
  .A1({ S18878 }),
  .A2({ S18879 }),
  .A3({ S18877 }),
  .ZN({ S18880 })
);
NAND2_X1 #() 
NAND2_X1_2690_ (
  .A1({ S18876 }),
  .A2({ S18880 }),
  .ZN({ S25957[32] })
);
NAND3_X1 #() 
NAND3_X1_2907_ (
  .A1({ S18713 }),
  .A2({ S18714 }),
  .A3({ S25957[161] }),
  .ZN({ S18881 })
);
INV_X1 #() 
INV_X1_834_ (
  .A({ S25957[161] }),
  .ZN({ S18882 })
);
NAND3_X1 #() 
NAND3_X1_2908_ (
  .A1({ S16577 }),
  .A2({ S16581 }),
  .A3({ S18710 }),
  .ZN({ S18884 })
);
NAND3_X1 #() 
NAND3_X1_2909_ (
  .A1({ S18711 }),
  .A2({ S18712 }),
  .A3({ S25957[193] }),
  .ZN({ S18885 })
);
NAND3_X1 #() 
NAND3_X1_2910_ (
  .A1({ S18884 }),
  .A2({ S18885 }),
  .A3({ S18882 }),
  .ZN({ S18886 })
);
NAND2_X1 #() 
NAND2_X1_2691_ (
  .A1({ S18881 }),
  .A2({ S18886 }),
  .ZN({ S25957[33] })
);
INV_X1 #() 
INV_X1_835_ (
  .A({ S25957[162] }),
  .ZN({ S18887 })
);
NAND2_X1 #() 
NAND2_X1_2692_ (
  .A1({ S25957[66] }),
  .A2({ S18887 }),
  .ZN({ S18888 })
);
NAND3_X1 #() 
NAND3_X1_2911_ (
  .A1({ S18715 }),
  .A2({ S18719 }),
  .A3({ S25957[162] }),
  .ZN({ S18889 })
);
NAND2_X1 #() 
NAND2_X1_2693_ (
  .A1({ S18888 }),
  .A2({ S18889 }),
  .ZN({ S25957[34] })
);
NAND3_X1 #() 
NAND3_X1_2912_ (
  .A1({ S18720 }),
  .A2({ S18723 }),
  .A3({ S25957[163] }),
  .ZN({ S18890 })
);
NAND3_X1 #() 
NAND3_X1_2913_ (
  .A1({ S18721 }),
  .A2({ S25957[195] }),
  .A3({ S18722 }),
  .ZN({ S18891 })
);
NAND3_X1 #() 
NAND3_X1_2914_ (
  .A1({ S16721 }),
  .A2({ S16300 }),
  .A3({ S16740 }),
  .ZN({ S18893 })
);
NAND3_X1 #() 
NAND3_X1_2915_ (
  .A1({ S18891 }),
  .A2({ S18893 }),
  .A3({ S16316 }),
  .ZN({ S18894 })
);
NAND2_X1 #() 
NAND2_X1_2694_ (
  .A1({ S18890 }),
  .A2({ S18894 }),
  .ZN({ S25957[35] })
);
XNOR2_X1 #() 
XNOR2_X1_142_ (
  .A({ S18732 }),
  .B({ S25957[164] }),
  .ZN({ S25957[36] })
);
OAI21_X1 #() 
OAI21_X1_1408_ (
  .A({ S25957[165] }),
  .B1({ S18736 }),
  .B2({ S18738 }),
  .ZN({ S18895 })
);
NAND3_X1 #() 
NAND3_X1_2916_ (
  .A1({ S16860 }),
  .A2({ S18737 }),
  .A3({ S16850 }),
  .ZN({ S18896 })
);
NAND3_X1 #() 
NAND3_X1_2917_ (
  .A1({ S18734 }),
  .A2({ S25957[197] }),
  .A3({ S18733 }),
  .ZN({ S18897 })
);
NAND3_X1 #() 
NAND3_X1_2918_ (
  .A1({ S18896 }),
  .A2({ S18897 }),
  .A3({ S16317 }),
  .ZN({ S18898 })
);
NAND2_X1 #() 
NAND2_X1_2695_ (
  .A1({ S18895 }),
  .A2({ S18898 }),
  .ZN({ S25957[37] })
);
OAI21_X1 #() 
OAI21_X1_1409_ (
  .A({ S25957[166] }),
  .B1({ S18741 }),
  .B2({ S18739 }),
  .ZN({ S18899 })
);
INV_X1 #() 
INV_X1_836_ (
  .A({ S25957[166] }),
  .ZN({ S18901 })
);
NAND2_X1 #() 
NAND2_X1_2696_ (
  .A1({ S16909 }),
  .A2({ S12198 }),
  .ZN({ S18902 })
);
NAND3_X1 #() 
NAND3_X1_2919_ (
  .A1({ S18902 }),
  .A2({ S18901 }),
  .A3({ S18740 }),
  .ZN({ S18903 })
);
NAND2_X1 #() 
NAND2_X1_2697_ (
  .A1({ S18899 }),
  .A2({ S18903 }),
  .ZN({ S25957[38] })
);
OAI21_X1 #() 
OAI21_X1_1410_ (
  .A({ S25957[167] }),
  .B1({ S18751 }),
  .B2({ S18752 }),
  .ZN({ S18904 })
);
NAND3_X1 #() 
NAND3_X1_2920_ (
  .A1({ S16935 }),
  .A2({ S16958 }),
  .A3({ S25957[327] }),
  .ZN({ S18905 })
);
NAND3_X1 #() 
NAND3_X1_2921_ (
  .A1({ S18748 }),
  .A2({ S18750 }),
  .A3({ S16274 }),
  .ZN({ S18906 })
);
NAND3_X1 #() 
NAND3_X1_2922_ (
  .A1({ S18906 }),
  .A2({ S18905 }),
  .A3({ S14960 }),
  .ZN({ S18907 })
);
NAND2_X1 #() 
NAND2_X1_2698_ (
  .A1({ S18904 }),
  .A2({ S18907 }),
  .ZN({ S25957[39] })
);
NAND3_X1 #() 
NAND3_X1_2923_ (
  .A1({ S17043 }),
  .A2({ S17094 }),
  .A3({ S25957[232] }),
  .ZN({ S18908 })
);
NAND3_X1 #() 
NAND3_X1_2924_ (
  .A1({ S17099 }),
  .A2({ S17106 }),
  .A3({ S16965 }),
  .ZN({ S18910 })
);
AOI21_X1 #() 
AOI21_X1_1508_ (
  .A({ S25957[296] }),
  .B1({ S18908 }),
  .B2({ S18910 }),
  .ZN({ S18911 })
);
AOI21_X1 #() 
AOI21_X1_1509_ (
  .A({ S14666 }),
  .B1({ S17095 }),
  .B2({ S17107 }),
  .ZN({ S18912 })
);
NOR2_X1 #() 
NOR2_X1_658_ (
  .A1({ S18911 }),
  .A2({ S18912 }),
  .ZN({ S25957[40] })
);
INV_X1 #() 
INV_X1_837_ (
  .A({ S25957[297] }),
  .ZN({ S18913 })
);
NAND2_X1 #() 
NAND2_X1_2699_ (
  .A1({ S25957[105] }),
  .A2({ S18913 }),
  .ZN({ S18914 })
);
NAND3_X1 #() 
NAND3_X1_2925_ (
  .A1({ S17183 }),
  .A2({ S25957[297] }),
  .A3({ S17181 }),
  .ZN({ S18915 })
);
NAND2_X1 #() 
NAND2_X1_2700_ (
  .A1({ S18914 }),
  .A2({ S18915 }),
  .ZN({ S25957[41] })
);
XNOR2_X1 #() 
XNOR2_X1_143_ (
  .A({ S18756 }),
  .B({ S25957[170] }),
  .ZN({ S25957[42] })
);
INV_X1 #() 
INV_X1_838_ (
  .A({ S25957[171] }),
  .ZN({ S18916 })
);
NAND3_X1 #() 
NAND3_X1_2926_ (
  .A1({ S18760 }),
  .A2({ S25957[203] }),
  .A3({ S18759 }),
  .ZN({ S18918 })
);
NAND3_X1 #() 
NAND3_X1_2927_ (
  .A1({ S17344 }),
  .A2({ S18758 }),
  .A3({ S17308 }),
  .ZN({ S18919 })
);
NAND3_X1 #() 
NAND3_X1_2928_ (
  .A1({ S18918 }),
  .A2({ S18919 }),
  .A3({ S18916 }),
  .ZN({ S18920 })
);
NAND3_X1 #() 
NAND3_X1_2929_ (
  .A1({ S18757 }),
  .A2({ S18761 }),
  .A3({ S25957[171] }),
  .ZN({ S18921 })
);
NAND2_X1 #() 
NAND2_X1_2701_ (
  .A1({ S18920 }),
  .A2({ S18921 }),
  .ZN({ S25957[43] })
);
INV_X1 #() 
INV_X1_839_ (
  .A({ S25957[300] }),
  .ZN({ S18922 })
);
NAND3_X1 #() 
NAND3_X1_2930_ (
  .A1({ S17374 }),
  .A2({ S17398 }),
  .A3({ S25957[236] }),
  .ZN({ S18923 })
);
NAND3_X1 #() 
NAND3_X1_2931_ (
  .A1({ S17405 }),
  .A2({ S17401 }),
  .A3({ S17345 }),
  .ZN({ S18924 })
);
NAND3_X1 #() 
NAND3_X1_2932_ (
  .A1({ S18923 }),
  .A2({ S18924 }),
  .A3({ S18922 }),
  .ZN({ S18925 })
);
NAND3_X1 #() 
NAND3_X1_2933_ (
  .A1({ S17399 }),
  .A2({ S17406 }),
  .A3({ S25957[300] }),
  .ZN({ S18926 })
);
NAND2_X1 #() 
NAND2_X1_2702_ (
  .A1({ S18925 }),
  .A2({ S18926 }),
  .ZN({ S25957[44] })
);
NAND2_X1 #() 
NAND2_X1_2703_ (
  .A1({ S25957[109] }),
  .A2({ S16320 }),
  .ZN({ S18928 })
);
NAND3_X1 #() 
NAND3_X1_2934_ (
  .A1({ S17461 }),
  .A2({ S17451 }),
  .A3({ S25957[301] }),
  .ZN({ S18929 })
);
NAND2_X1 #() 
NAND2_X1_2704_ (
  .A1({ S18928 }),
  .A2({ S18929 }),
  .ZN({ S25957[45] })
);
NAND3_X1 #() 
NAND3_X1_2935_ (
  .A1({ S18765 }),
  .A2({ S18766 }),
  .A3({ S25957[174] }),
  .ZN({ S18930 })
);
INV_X1 #() 
INV_X1_840_ (
  .A({ S25957[174] }),
  .ZN({ S18931 })
);
NAND3_X1 #() 
NAND3_X1_2936_ (
  .A1({ S18763 }),
  .A2({ S18764 }),
  .A3({ S25957[206] }),
  .ZN({ S18932 })
);
NAND3_X1 #() 
NAND3_X1_2937_ (
  .A1({ S17508 }),
  .A2({ S17521 }),
  .A3({ S14359 }),
  .ZN({ S18933 })
);
NAND3_X1 #() 
NAND3_X1_2938_ (
  .A1({ S18932 }),
  .A2({ S18933 }),
  .A3({ S18931 }),
  .ZN({ S18934 })
);
NAND2_X1 #() 
NAND2_X1_2705_ (
  .A1({ S18930 }),
  .A2({ S18934 }),
  .ZN({ S25957[46] })
);
OAI21_X1 #() 
OAI21_X1_1411_ (
  .A({ S25957[175] }),
  .B1({ S18785 }),
  .B2({ S18784 }),
  .ZN({ S18936 })
);
INV_X1 #() 
INV_X1_841_ (
  .A({ S25957[175] }),
  .ZN({ S18937 })
);
NAND3_X1 #() 
NAND3_X1_2939_ (
  .A1({ S17546 }),
  .A2({ S25957[335] }),
  .A3({ S17569 }),
  .ZN({ S18938 })
);
NAND3_X1 #() 
NAND3_X1_2940_ (
  .A1({ S18783 }),
  .A2({ S18778 }),
  .A3({ S16305 }),
  .ZN({ S18939 })
);
NAND3_X1 #() 
NAND3_X1_2941_ (
  .A1({ S18938 }),
  .A2({ S18939 }),
  .A3({ S18937 }),
  .ZN({ S18940 })
);
NAND2_X1 #() 
NAND2_X1_2706_ (
  .A1({ S18936 }),
  .A2({ S18940 }),
  .ZN({ S25957[47] })
);
NAND3_X1 #() 
NAND3_X1_2942_ (
  .A1({ S18786 }),
  .A2({ S18789 }),
  .A3({ S25957[176] }),
  .ZN({ S18941 })
);
INV_X1 #() 
INV_X1_842_ (
  .A({ S25957[176] }),
  .ZN({ S18942 })
);
NAND3_X1 #() 
NAND3_X1_2943_ (
  .A1({ S18788 }),
  .A2({ S25957[208] }),
  .A3({ S18787 }),
  .ZN({ S18943 })
);
NAND3_X1 #() 
NAND3_X1_2944_ (
  .A1({ S17717 }),
  .A2({ S16308 }),
  .A3({ S17690 }),
  .ZN({ S18944 })
);
NAND3_X1 #() 
NAND3_X1_2945_ (
  .A1({ S18943 }),
  .A2({ S18944 }),
  .A3({ S18942 }),
  .ZN({ S18946 })
);
NAND2_X1 #() 
NAND2_X1_2707_ (
  .A1({ S18941 }),
  .A2({ S18946 }),
  .ZN({ S25957[48] })
);
INV_X1 #() 
INV_X1_843_ (
  .A({ S25957[305] }),
  .ZN({ S18947 })
);
XNOR2_X1 #() 
XNOR2_X1_144_ (
  .A({ S25957[113] }),
  .B({ S18947 }),
  .ZN({ S25957[49] })
);
NAND2_X1 #() 
NAND2_X1_2708_ (
  .A1({ S25957[82] }),
  .A2({ S16323 }),
  .ZN({ S18948 })
);
OAI21_X1 #() 
OAI21_X1_1412_ (
  .A({ S25957[178] }),
  .B1({ S18796 }),
  .B2({ S18797 }),
  .ZN({ S18949 })
);
NAND2_X1 #() 
NAND2_X1_2709_ (
  .A1({ S18948 }),
  .A2({ S18949 }),
  .ZN({ S25957[50] })
);
OAI21_X1 #() 
OAI21_X1_1413_ (
  .A({ S25957[179] }),
  .B1({ S18800 }),
  .B2({ S18801 }),
  .ZN({ S18950 })
);
INV_X1 #() 
INV_X1_844_ (
  .A({ S25957[179] }),
  .ZN({ S18951 })
);
INV_X1 #() 
INV_X1_845_ (
  .A({ S18801 }),
  .ZN({ S18952 })
);
NAND3_X1 #() 
NAND3_X1_2946_ (
  .A1({ S18952 }),
  .A2({ S18799 }),
  .A3({ S18951 }),
  .ZN({ S18954 })
);
NAND2_X1 #() 
NAND2_X1_2710_ (
  .A1({ S18950 }),
  .A2({ S18954 }),
  .ZN({ S25957[51] })
);
INV_X1 #() 
INV_X1_846_ (
  .A({ S18802 }),
  .ZN({ S18955 })
);
OAI22_X1 #() 
OAI22_X1_66_ (
  .A1({ S18955 }),
  .A2({ S18803 }),
  .B1({ S13770 }),
  .B2({ S13767 }),
  .ZN({ S18956 })
);
NAND3_X1 #() 
NAND3_X1_2947_ (
  .A1({ S18804 }),
  .A2({ S25957[180] }),
  .A3({ S18802 }),
  .ZN({ S18957 })
);
NAND2_X1 #() 
NAND2_X1_2711_ (
  .A1({ S18956 }),
  .A2({ S18957 }),
  .ZN({ S25957[52] })
);
OAI21_X1 #() 
OAI21_X1_1414_ (
  .A({ S25957[181] }),
  .B1({ S18806 }),
  .B2({ S18808 }),
  .ZN({ S18958 })
);
INV_X1 #() 
INV_X1_847_ (
  .A({ S25957[341] }),
  .ZN({ S18959 })
);
NAND2_X1 #() 
NAND2_X1_2712_ (
  .A1({ S18050 }),
  .A2({ S18959 }),
  .ZN({ S18960 })
);
NAND3_X1 #() 
NAND3_X1_2948_ (
  .A1({ S18960 }),
  .A2({ S18805 }),
  .A3({ S16325 }),
  .ZN({ S18961 })
);
NAND2_X1 #() 
NAND2_X1_2713_ (
  .A1({ S18958 }),
  .A2({ S18961 }),
  .ZN({ S25957[53] })
);
AND3_X1 #() 
AND3_X1_115_ (
  .A1({ S18104 }),
  .A2({ S18095 }),
  .A3({ S16326 }),
  .ZN({ S18963 })
);
AOI21_X1 #() 
AOI21_X1_1510_ (
  .A({ S16326 }),
  .B1({ S18095 }),
  .B2({ S18104 }),
  .ZN({ S18964 })
);
NOR2_X1 #() 
NOR2_X1_659_ (
  .A1({ S18963 }),
  .A2({ S18964 }),
  .ZN({ S25957[54] })
);
NAND3_X1 #() 
NAND3_X1_2949_ (
  .A1({ S18154 }),
  .A2({ S18149 }),
  .A3({ S25957[311] }),
  .ZN({ S18965 })
);
NAND3_X1 #() 
NAND3_X1_2950_ (
  .A1({ S18128 }),
  .A2({ S18148 }),
  .A3({ S13519 }),
  .ZN({ S18966 })
);
OAI211_X1 #() 
OAI211_X1_983_ (
  .A({ S18153 }),
  .B({ S25957[247] }),
  .C1({ S18150 }),
  .C2({ S25957[143] }),
  .ZN({ S18967 })
);
NAND3_X1 #() 
NAND3_X1_2951_ (
  .A1({ S18967 }),
  .A2({ S18966 }),
  .A3({ S10651 }),
  .ZN({ S18968 })
);
NAND2_X1 #() 
NAND2_X1_2714_ (
  .A1({ S18965 }),
  .A2({ S18968 }),
  .ZN({ S25957[55] })
);
INV_X1 #() 
INV_X1_848_ (
  .A({ S25957[184] }),
  .ZN({ S18969 })
);
NAND2_X1 #() 
NAND2_X1_2715_ (
  .A1({ S25957[88] }),
  .A2({ S18969 }),
  .ZN({ S18971 })
);
NAND3_X1 #() 
NAND3_X1_2952_ (
  .A1({ S18813 }),
  .A2({ S18812 }),
  .A3({ S25957[184] }),
  .ZN({ S18972 })
);
NAND2_X1 #() 
NAND2_X1_2716_ (
  .A1({ S18971 }),
  .A2({ S18972 }),
  .ZN({ S25957[56] })
);
NAND3_X1 #() 
NAND3_X1_2953_ (
  .A1({ S18817 }),
  .A2({ S25957[185] }),
  .A3({ S18815 }),
  .ZN({ S18973 })
);
INV_X1 #() 
INV_X1_849_ (
  .A({ S18815 }),
  .ZN({ S18974 })
);
OAI22_X1 #() 
OAI22_X1_67_ (
  .A1({ S18974 }),
  .A2({ S18816 }),
  .B1({ S16180 }),
  .B2({ S16176 }),
  .ZN({ S18975 })
);
NAND2_X1 #() 
NAND2_X1_2717_ (
  .A1({ S18975 }),
  .A2({ S18973 }),
  .ZN({ S25957[57] })
);
NAND2_X1 #() 
NAND2_X1_2718_ (
  .A1({ S25957[90] }),
  .A2({ S16328 }),
  .ZN({ S18976 })
);
NAND3_X1 #() 
NAND3_X1_2954_ (
  .A1({ S18820 }),
  .A2({ S18818 }),
  .A3({ S25957[186] }),
  .ZN({ S18977 })
);
NAND2_X1 #() 
NAND2_X1_2719_ (
  .A1({ S18976 }),
  .A2({ S18977 }),
  .ZN({ S25957[58] })
);
OAI21_X1 #() 
OAI21_X1_1415_ (
  .A({ S25957[187] }),
  .B1({ S18833 }),
  .B2({ S18835 }),
  .ZN({ S18979 })
);
INV_X1 #() 
INV_X1_850_ (
  .A({ S25957[187] }),
  .ZN({ S18980 })
);
NAND3_X1 #() 
NAND3_X1_2955_ (
  .A1({ S18468 }),
  .A2({ S25957[347] }),
  .A3({ S18493 }),
  .ZN({ S18981 })
);
NAND3_X1 #() 
NAND3_X1_2956_ (
  .A1({ S18832 }),
  .A2({ S18830 }),
  .A3({ S15910 }),
  .ZN({ S18982 })
);
NAND3_X1 #() 
NAND3_X1_2957_ (
  .A1({ S18982 }),
  .A2({ S18981 }),
  .A3({ S18980 }),
  .ZN({ S18983 })
);
NAND2_X1 #() 
NAND2_X1_2720_ (
  .A1({ S18979 }),
  .A2({ S18983 }),
  .ZN({ S25957[59] })
);
XNOR2_X1 #() 
XNOR2_X1_145_ (
  .A({ S25957[92] }),
  .B({ S16329 }),
  .ZN({ S25957[60] })
);
XNOR2_X1 #() 
XNOR2_X1_146_ (
  .A({ S18840 }),
  .B({ S25957[189] }),
  .ZN({ S25957[61] })
);
NAND3_X1 #() 
NAND3_X1_2958_ (
  .A1({ S18841 }),
  .A2({ S18846 }),
  .A3({ S25957[190] }),
  .ZN({ S18984 })
);
INV_X1 #() 
INV_X1_851_ (
  .A({ S25957[190] }),
  .ZN({ S18985 })
);
NAND3_X1 #() 
NAND3_X1_2959_ (
  .A1({ S18844 }),
  .A2({ S25957[222] }),
  .A3({ S18845 }),
  .ZN({ S18987 })
);
NAND3_X1 #() 
NAND3_X1_2960_ (
  .A1({ S18655 }),
  .A2({ S18843 }),
  .A3({ S18629 }),
  .ZN({ S18988 })
);
NAND3_X1 #() 
NAND3_X1_2961_ (
  .A1({ S18987 }),
  .A2({ S18988 }),
  .A3({ S18985 }),
  .ZN({ S18989 })
);
NAND2_X1 #() 
NAND2_X1_2721_ (
  .A1({ S18984 }),
  .A2({ S18989 }),
  .ZN({ S25957[62] })
);
NAND3_X1 #() 
NAND3_X1_2962_ (
  .A1({ S18875 }),
  .A2({ S25957[191] }),
  .A3({ S18872 }),
  .ZN({ S18990 })
);
INV_X1 #() 
INV_X1_852_ (
  .A({ S25957[191] }),
  .ZN({ S18991 })
);
AOI21_X1 #() 
AOI21_X1_1511_ (
  .A({ S18873 }),
  .B1({ S18702 }),
  .B2({ S18679 }),
  .ZN({ S18992 })
);
AOI21_X1 #() 
AOI21_X1_1512_ (
  .A({ S25957[351] }),
  .B1({ S18856 }),
  .B2({ S18871 }),
  .ZN({ S18993 })
);
OAI21_X1 #() 
OAI21_X1_1416_ (
  .A({ S18991 }),
  .B1({ S18992 }),
  .B2({ S18993 }),
  .ZN({ S18994 })
);
NAND2_X1 #() 
NAND2_X1_2722_ (
  .A1({ S18994 }),
  .A2({ S18990 }),
  .ZN({ S25957[63] })
);
NAND3_X1 #() 
NAND3_X1_2963_ (
  .A1({ S18876 }),
  .A2({ S25957[128] }),
  .A3({ S18880 }),
  .ZN({ S18996 })
);
OAI21_X1 #() 
OAI21_X1_1417_ (
  .A({ S18877 }),
  .B1({ S18706 }),
  .B2({ S18709 }),
  .ZN({ S18997 })
);
NAND3_X1 #() 
NAND3_X1_2964_ (
  .A1({ S18878 }),
  .A2({ S18879 }),
  .A3({ S25957[160] }),
  .ZN({ S18998 })
);
NAND3_X1 #() 
NAND3_X1_2965_ (
  .A1({ S18997 }),
  .A2({ S16964 }),
  .A3({ S18998 }),
  .ZN({ S18999 })
);
NAND2_X1 #() 
NAND2_X1_2723_ (
  .A1({ S18996 }),
  .A2({ S18999 }),
  .ZN({ S25957[0] })
);
NAND3_X1 #() 
NAND3_X1_2966_ (
  .A1({ S18713 }),
  .A2({ S18714 }),
  .A3({ S25957[257] }),
  .ZN({ S19000 })
);
NAND3_X1 #() 
NAND3_X1_2967_ (
  .A1({ S18884 }),
  .A2({ S18885 }),
  .A3({ S14141 }),
  .ZN({ S19001 })
);
NAND2_X1 #() 
NAND2_X1_2724_ (
  .A1({ S19000 }),
  .A2({ S19001 }),
  .ZN({ S25957[1] })
);
NAND3_X1 #() 
NAND3_X1_2968_ (
  .A1({ S18715 }),
  .A2({ S18719 }),
  .A3({ S14154 }),
  .ZN({ S19002 })
);
NAND3_X1 #() 
NAND3_X1_2969_ (
  .A1({ S18717 }),
  .A2({ S18718 }),
  .A3({ S25957[194] }),
  .ZN({ S19003 })
);
NAND3_X1 #() 
NAND3_X1_2970_ (
  .A1({ S16644 }),
  .A2({ S16661 }),
  .A3({ S16299 }),
  .ZN({ S19005 })
);
NAND3_X1 #() 
NAND3_X1_2971_ (
  .A1({ S19003 }),
  .A2({ S19005 }),
  .A3({ S25957[258] }),
  .ZN({ S19006 })
);
AND2_X1 #() 
AND2_X1_176_ (
  .A1({ S19006 }),
  .A2({ S19002 }),
  .ZN({ S25957[2] })
);
NAND3_X1 #() 
NAND3_X1_2972_ (
  .A1({ S18891 }),
  .A2({ S18893 }),
  .A3({ S38 }),
  .ZN({ S19007 })
);
NAND3_X1 #() 
NAND3_X1_2973_ (
  .A1({ S18720 }),
  .A2({ S18723 }),
  .A3({ S25957[259] }),
  .ZN({ S19008 })
);
NAND2_X1 #() 
NAND2_X1_2725_ (
  .A1({ S19007 }),
  .A2({ S19008 }),
  .ZN({ S25957[3] })
);
XNOR2_X1 #() 
XNOR2_X1_147_ (
  .A({ S18732 }),
  .B({ S25957[260] }),
  .ZN({ S25957[4] })
);
AOI21_X1 #() 
AOI21_X1_1513_ (
  .A({ S16317 }),
  .B1({ S18896 }),
  .B2({ S18897 }),
  .ZN({ S19009 })
);
AND3_X1 #() 
AND3_X1_116_ (
  .A1({ S18897 }),
  .A2({ S18896 }),
  .A3({ S16317 }),
  .ZN({ S19010 })
);
OAI21_X1 #() 
OAI21_X1_1418_ (
  .A({ S16967 }),
  .B1({ S19010 }),
  .B2({ S19009 }),
  .ZN({ S19011 })
);
NAND3_X1 #() 
NAND3_X1_2974_ (
  .A1({ S18895 }),
  .A2({ S25957[133] }),
  .A3({ S18898 }),
  .ZN({ S19013 })
);
NAND2_X1 #() 
NAND2_X1_2726_ (
  .A1({ S19011 }),
  .A2({ S19013 }),
  .ZN({ S25957[5] })
);
AOI21_X1 #() 
AOI21_X1_1514_ (
  .A({ S18901 }),
  .B1({ S18902 }),
  .B2({ S18740 }),
  .ZN({ S19014 })
);
NOR3_X1 #() 
NOR3_X1_92_ (
  .A1({ S18741 }),
  .A2({ S18739 }),
  .A3({ S25957[166] }),
  .ZN({ S19015 })
);
OAI21_X1 #() 
OAI21_X1_1419_ (
  .A({ S15041 }),
  .B1({ S19015 }),
  .B2({ S19014 }),
  .ZN({ S19016 })
);
NAND3_X1 #() 
NAND3_X1_2975_ (
  .A1({ S18899 }),
  .A2({ S18903 }),
  .A3({ S25957[134] }),
  .ZN({ S19017 })
);
NAND2_X1 #() 
NAND2_X1_2727_ (
  .A1({ S19016 }),
  .A2({ S19017 }),
  .ZN({ S25957[6] })
);
OAI21_X1 #() 
OAI21_X1_1420_ (
  .A({ S14960 }),
  .B1({ S18751 }),
  .B2({ S18752 }),
  .ZN({ S19018 })
);
NAND3_X1 #() 
NAND3_X1_2976_ (
  .A1({ S18906 }),
  .A2({ S18905 }),
  .A3({ S25957[167] }),
  .ZN({ S19019 })
);
NAND3_X1 #() 
NAND3_X1_2977_ (
  .A1({ S19018 }),
  .A2({ S16966 }),
  .A3({ S19019 }),
  .ZN({ S19020 })
);
NAND3_X1 #() 
NAND3_X1_2978_ (
  .A1({ S18904 }),
  .A2({ S25957[135] }),
  .A3({ S18907 }),
  .ZN({ S19022 })
);
NAND2_X1 #() 
NAND2_X1_2728_ (
  .A1({ S19020 }),
  .A2({ S19022 }),
  .ZN({ S25957[7] })
);
NAND3_X1 #() 
NAND3_X1_2979_ (
  .A1({ S17095 }),
  .A2({ S17107 }),
  .A3({ S14666 }),
  .ZN({ S19023 })
);
NAND3_X1 #() 
NAND3_X1_2980_ (
  .A1({ S18908 }),
  .A2({ S18910 }),
  .A3({ S25957[296] }),
  .ZN({ S19024 })
);
NAND3_X1 #() 
NAND3_X1_2981_ (
  .A1({ S19023 }),
  .A2({ S19024 }),
  .A3({ S17621 }),
  .ZN({ S19025 })
);
OAI21_X1 #() 
OAI21_X1_1421_ (
  .A({ S25957[136] }),
  .B1({ S18911 }),
  .B2({ S18912 }),
  .ZN({ S19026 })
);
NAND2_X1 #() 
NAND2_X1_2729_ (
  .A1({ S19026 }),
  .A2({ S19025 }),
  .ZN({ S25957[8] })
);
AOI21_X1 #() 
AOI21_X1_1515_ (
  .A({ S25957[297] }),
  .B1({ S17183 }),
  .B2({ S17181 }),
  .ZN({ S19027 })
);
NAND2_X1 #() 
NAND2_X1_2730_ (
  .A1({ S17182 }),
  .A2({ S17108 }),
  .ZN({ S19028 })
);
NAND3_X1 #() 
NAND3_X1_2982_ (
  .A1({ S17180 }),
  .A2({ S17148 }),
  .A3({ S25957[233] }),
  .ZN({ S19029 })
);
AOI21_X1 #() 
AOI21_X1_1516_ (
  .A({ S18913 }),
  .B1({ S19028 }),
  .B2({ S19029 }),
  .ZN({ S19031 })
);
OAI21_X1 #() 
OAI21_X1_1422_ (
  .A({ S17575 }),
  .B1({ S19027 }),
  .B2({ S19031 }),
  .ZN({ S19032 })
);
NAND3_X1 #() 
NAND3_X1_2983_ (
  .A1({ S18914 }),
  .A2({ S18915 }),
  .A3({ S25957[137] }),
  .ZN({ S19033 })
);
NAND2_X1 #() 
NAND2_X1_2731_ (
  .A1({ S19033 }),
  .A2({ S19032 }),
  .ZN({ S25957[9] })
);
XNOR2_X1 #() 
XNOR2_X1_148_ (
  .A({ S18756 }),
  .B({ S25957[266] }),
  .ZN({ S25957[10] })
);
AOI21_X1 #() 
AOI21_X1_1517_ (
  .A({ S25957[171] }),
  .B1({ S18757 }),
  .B2({ S18761 }),
  .ZN({ S19034 })
);
AOI21_X1 #() 
AOI21_X1_1518_ (
  .A({ S18916 }),
  .B1({ S18918 }),
  .B2({ S18919 }),
  .ZN({ S19035 })
);
OAI21_X1 #() 
OAI21_X1_1423_ (
  .A({ S47 }),
  .B1({ S19034 }),
  .B2({ S19035 }),
  .ZN({ S19036 })
);
NAND3_X1 #() 
NAND3_X1_2984_ (
  .A1({ S18920 }),
  .A2({ S18921 }),
  .A3({ S25957[139] }),
  .ZN({ S19037 })
);
NAND2_X1 #() 
NAND2_X1_2732_ (
  .A1({ S19036 }),
  .A2({ S19037 }),
  .ZN({ S25957[11] })
);
NAND3_X1 #() 
NAND3_X1_2985_ (
  .A1({ S18925 }),
  .A2({ S18926 }),
  .A3({ S25957[140] }),
  .ZN({ S19039 })
);
NAND3_X1 #() 
NAND3_X1_2986_ (
  .A1({ S17399 }),
  .A2({ S17406 }),
  .A3({ S18922 }),
  .ZN({ S19040 })
);
NAND3_X1 #() 
NAND3_X1_2987_ (
  .A1({ S18923 }),
  .A2({ S18924 }),
  .A3({ S25957[300] }),
  .ZN({ S19041 })
);
NAND3_X1 #() 
NAND3_X1_2988_ (
  .A1({ S19040 }),
  .A2({ S19041 }),
  .A3({ S17578 }),
  .ZN({ S19042 })
);
NAND2_X1 #() 
NAND2_X1_2733_ (
  .A1({ S19039 }),
  .A2({ S19042 }),
  .ZN({ S25957[12] })
);
AOI21_X1 #() 
AOI21_X1_1519_ (
  .A({ S25957[301] }),
  .B1({ S17461 }),
  .B2({ S17451 }),
  .ZN({ S19043 })
);
NAND3_X1 #() 
NAND3_X1_2989_ (
  .A1({ S17450 }),
  .A2({ S17426 }),
  .A3({ S25957[237] }),
  .ZN({ S19044 })
);
NAND3_X1 #() 
NAND3_X1_2990_ (
  .A1({ S17453 }),
  .A2({ S17460 }),
  .A3({ S14448 }),
  .ZN({ S19045 })
);
AOI21_X1 #() 
AOI21_X1_1520_ (
  .A({ S16320 }),
  .B1({ S19045 }),
  .B2({ S19044 }),
  .ZN({ S19046 })
);
OAI21_X1 #() 
OAI21_X1_1424_ (
  .A({ S17577 }),
  .B1({ S19043 }),
  .B2({ S19046 }),
  .ZN({ S19047 })
);
NAND3_X1 #() 
NAND3_X1_2991_ (
  .A1({ S18928 }),
  .A2({ S18929 }),
  .A3({ S25957[141] }),
  .ZN({ S19049 })
);
NAND2_X1 #() 
NAND2_X1_2734_ (
  .A1({ S19049 }),
  .A2({ S19047 }),
  .ZN({ S25957[13] })
);
NAND3_X1 #() 
NAND3_X1_2992_ (
  .A1({ S18932 }),
  .A2({ S18933 }),
  .A3({ S13391 }),
  .ZN({ S19050 })
);
NAND3_X1 #() 
NAND3_X1_2993_ (
  .A1({ S18765 }),
  .A2({ S18766 }),
  .A3({ S25957[270] }),
  .ZN({ S19051 })
);
NAND2_X1 #() 
NAND2_X1_2735_ (
  .A1({ S19050 }),
  .A2({ S19051 }),
  .ZN({ S25957[14] })
);
NAND3_X1 #() 
NAND3_X1_2994_ (
  .A1({ S18936 }),
  .A2({ S25957[143] }),
  .A3({ S18940 }),
  .ZN({ S19052 })
);
OAI21_X1 #() 
OAI21_X1_1425_ (
  .A({ S18937 }),
  .B1({ S18785 }),
  .B2({ S18784 }),
  .ZN({ S19053 })
);
NAND3_X1 #() 
NAND3_X1_2995_ (
  .A1({ S18938 }),
  .A2({ S18939 }),
  .A3({ S25957[175] }),
  .ZN({ S19054 })
);
NAND3_X1 #() 
NAND3_X1_2996_ (
  .A1({ S19053 }),
  .A2({ S14271 }),
  .A3({ S19054 }),
  .ZN({ S19055 })
);
NAND2_X1 #() 
NAND2_X1_2736_ (
  .A1({ S19052 }),
  .A2({ S19055 }),
  .ZN({ S25957[15] })
);
NAND3_X1 #() 
NAND3_X1_2997_ (
  .A1({ S18941 }),
  .A2({ S18946 }),
  .A3({ S25957[144] }),
  .ZN({ S19057 })
);
NAND3_X1 #() 
NAND3_X1_2998_ (
  .A1({ S18943 }),
  .A2({ S18944 }),
  .A3({ S25957[176] }),
  .ZN({ S19058 })
);
NAND3_X1 #() 
NAND3_X1_2999_ (
  .A1({ S18786 }),
  .A2({ S18789 }),
  .A3({ S18942 }),
  .ZN({ S19059 })
);
NAND3_X1 #() 
NAND3_X1_3000_ (
  .A1({ S19058 }),
  .A2({ S19059 }),
  .A3({ S18170 }),
  .ZN({ S19060 })
);
NAND2_X1 #() 
NAND2_X1_2737_ (
  .A1({ S19057 }),
  .A2({ S19060 }),
  .ZN({ S25957[16] })
);
NAND3_X1 #() 
NAND3_X1_3001_ (
  .A1({ S18791 }),
  .A2({ S18794 }),
  .A3({ S25957[273] }),
  .ZN({ S19061 })
);
NAND3_X1 #() 
NAND3_X1_3002_ (
  .A1({ S18793 }),
  .A2({ S18792 }),
  .A3({ S25957[209] }),
  .ZN({ S19062 })
);
NAND3_X1 #() 
NAND3_X1_3003_ (
  .A1({ S17818 }),
  .A2({ S17801 }),
  .A3({ S16310 }),
  .ZN({ S19063 })
);
NAND3_X1 #() 
NAND3_X1_3004_ (
  .A1({ S19062 }),
  .A2({ S19063 }),
  .A3({ S15527 }),
  .ZN({ S19064 })
);
NAND2_X1 #() 
NAND2_X1_2738_ (
  .A1({ S19061 }),
  .A2({ S19064 }),
  .ZN({ S25957[17] })
);
INV_X1 #() 
INV_X1_853_ (
  .A({ S18797 }),
  .ZN({ S19066 })
);
AOI21_X1 #() 
AOI21_X1_1521_ (
  .A({ S25957[274] }),
  .B1({ S19066 }),
  .B2({ S18795 }),
  .ZN({ S19067 })
);
NOR3_X1 #() 
NOR3_X1_93_ (
  .A1({ S18796 }),
  .A2({ S18797 }),
  .A3({ S15553 }),
  .ZN({ S19068 })
);
NOR2_X1 #() 
NOR2_X1_660_ (
  .A1({ S19067 }),
  .A2({ S19068 }),
  .ZN({ S25957[18] })
);
OAI21_X1 #() 
OAI21_X1_1426_ (
  .A({ S25957[275] }),
  .B1({ S18800 }),
  .B2({ S18801 }),
  .ZN({ S19069 })
);
NAND3_X1 #() 
NAND3_X1_3005_ (
  .A1({ S18952 }),
  .A2({ S18799 }),
  .A3({ S32 }),
  .ZN({ S19070 })
);
NAND2_X1 #() 
NAND2_X1_2739_ (
  .A1({ S19069 }),
  .A2({ S19070 }),
  .ZN({ S25957[19] })
);
OAI21_X1 #() 
OAI21_X1_1427_ (
  .A({ S13772 }),
  .B1({ S18955 }),
  .B2({ S18803 }),
  .ZN({ S19071 })
);
NAND3_X1 #() 
NAND3_X1_3006_ (
  .A1({ S18804 }),
  .A2({ S25957[276] }),
  .A3({ S18802 }),
  .ZN({ S19072 })
);
NAND2_X1 #() 
NAND2_X1_2740_ (
  .A1({ S19071 }),
  .A2({ S19072 }),
  .ZN({ S25957[20] })
);
AOI21_X1 #() 
AOI21_X1_1522_ (
  .A({ S25957[277] }),
  .B1({ S18960 }),
  .B2({ S18805 }),
  .ZN({ S19074 })
);
NOR3_X1 #() 
NOR3_X1_94_ (
  .A1({ S18806 }),
  .A2({ S18808 }),
  .A3({ S15621 }),
  .ZN({ S19075 })
);
NOR2_X1 #() 
NOR2_X1_661_ (
  .A1({ S19075 }),
  .A2({ S19074 }),
  .ZN({ S25957[21] })
);
NAND3_X1 #() 
NAND3_X1_3007_ (
  .A1({ S18095 }),
  .A2({ S18104 }),
  .A3({ S16326 }),
  .ZN({ S19076 })
);
NAND2_X1 #() 
NAND2_X1_2741_ (
  .A1({ S25957[118] }),
  .A2({ S25957[310] }),
  .ZN({ S19077 })
);
NAND3_X1 #() 
NAND3_X1_3008_ (
  .A1({ S19077 }),
  .A2({ S18185 }),
  .A3({ S19076 }),
  .ZN({ S19078 })
);
OAI21_X1 #() 
OAI21_X1_1428_ (
  .A({ S25957[150] }),
  .B1({ S18963 }),
  .B2({ S18964 }),
  .ZN({ S19079 })
);
NAND2_X1 #() 
NAND2_X1_2742_ (
  .A1({ S19079 }),
  .A2({ S19078 }),
  .ZN({ S25957[22] })
);
NAND3_X1 #() 
NAND3_X1_3009_ (
  .A1({ S18967 }),
  .A2({ S18966 }),
  .A3({ S25957[311] }),
  .ZN({ S19080 })
);
NAND3_X1 #() 
NAND3_X1_3010_ (
  .A1({ S18154 }),
  .A2({ S18149 }),
  .A3({ S10651 }),
  .ZN({ S19081 })
);
NAND3_X1 #() 
NAND3_X1_3011_ (
  .A1({ S19080 }),
  .A2({ S19081 }),
  .A3({ S13526 }),
  .ZN({ S19083 })
);
NAND3_X1 #() 
NAND3_X1_3012_ (
  .A1({ S18965 }),
  .A2({ S18968 }),
  .A3({ S25957[151] }),
  .ZN({ S19084 })
);
NAND2_X1 #() 
NAND2_X1_2743_ (
  .A1({ S19083 }),
  .A2({ S19084 }),
  .ZN({ S25957[23] })
);
AOI21_X1 #() 
AOI21_X1_1523_ (
  .A({ S25957[184] }),
  .B1({ S18813 }),
  .B2({ S18812 }),
  .ZN({ S19085 })
);
AND3_X1 #() 
AND3_X1_117_ (
  .A1({ S18813 }),
  .A2({ S18812 }),
  .A3({ S25957[184] }),
  .ZN({ S19086 })
);
OAI21_X1 #() 
OAI21_X1_1429_ (
  .A({ S16337 }),
  .B1({ S19086 }),
  .B2({ S19085 }),
  .ZN({ S19087 })
);
NAND3_X1 #() 
NAND3_X1_3013_ (
  .A1({ S18971 }),
  .A2({ S25957[152] }),
  .A3({ S18972 }),
  .ZN({ S19088 })
);
NAND2_X1 #() 
NAND2_X1_2744_ (
  .A1({ S19087 }),
  .A2({ S19088 }),
  .ZN({ S25957[24] })
);
NAND3_X1 #() 
NAND3_X1_3014_ (
  .A1({ S18817 }),
  .A2({ S25957[281] }),
  .A3({ S18815 }),
  .ZN({ S19089 })
);
OAI21_X1 #() 
OAI21_X1_1430_ (
  .A({ S14841 }),
  .B1({ S18974 }),
  .B2({ S18816 }),
  .ZN({ S19090 })
);
NAND2_X1 #() 
NAND2_X1_2745_ (
  .A1({ S19089 }),
  .A2({ S19090 }),
  .ZN({ S25957[25] })
);
NAND2_X1 #() 
NAND2_X1_2746_ (
  .A1({ S25957[90] }),
  .A2({ S14834 }),
  .ZN({ S19092 })
);
NAND3_X1 #() 
NAND3_X1_3015_ (
  .A1({ S18820 }),
  .A2({ S25957[282] }),
  .A3({ S18818 }),
  .ZN({ S19093 })
);
NAND2_X1 #() 
NAND2_X1_2747_ (
  .A1({ S19092 }),
  .A2({ S19093 }),
  .ZN({ S25957[26] })
);
NAND3_X1 #() 
NAND3_X1_3016_ (
  .A1({ S18979 }),
  .A2({ S25957[155] }),
  .A3({ S18983 }),
  .ZN({ S19094 })
);
OAI21_X1 #() 
OAI21_X1_1431_ (
  .A({ S18980 }),
  .B1({ S18833 }),
  .B2({ S18835 }),
  .ZN({ S19095 })
);
NAND3_X1 #() 
NAND3_X1_3017_ (
  .A1({ S18982 }),
  .A2({ S18981 }),
  .A3({ S25957[187] }),
  .ZN({ S19096 })
);
NAND3_X1 #() 
NAND3_X1_3018_ (
  .A1({ S19095 }),
  .A2({ S54 }),
  .A3({ S19096 }),
  .ZN({ S19097 })
);
NAND2_X1 #() 
NAND2_X1_2748_ (
  .A1({ S19094 }),
  .A2({ S19097 }),
  .ZN({ S25957[27] })
);
XNOR2_X1 #() 
XNOR2_X1_149_ (
  .A({ S25957[92] }),
  .B({ S14852 }),
  .ZN({ S25957[28] })
);
XNOR2_X1 #() 
XNOR2_X1_150_ (
  .A({ S18840 }),
  .B({ S25957[285] }),
  .ZN({ S25957[29] })
);
NAND3_X1 #() 
NAND3_X1_3019_ (
  .A1({ S18984 }),
  .A2({ S18989 }),
  .A3({ S25957[158] }),
  .ZN({ S19099 })
);
NAND3_X1 #() 
NAND3_X1_3020_ (
  .A1({ S18987 }),
  .A2({ S18988 }),
  .A3({ S25957[190] }),
  .ZN({ S19100 })
);
NAND3_X1 #() 
NAND3_X1_3021_ (
  .A1({ S18841 }),
  .A2({ S18846 }),
  .A3({ S18985 }),
  .ZN({ S19101 })
);
NAND3_X1 #() 
NAND3_X1_3022_ (
  .A1({ S19100 }),
  .A2({ S19101 }),
  .A3({ S15729 }),
  .ZN({ S19102 })
);
NAND2_X1 #() 
NAND2_X1_2749_ (
  .A1({ S19099 }),
  .A2({ S19102 }),
  .ZN({ S25957[30] })
);
OAI21_X1 #() 
OAI21_X1_1432_ (
  .A({ S25957[191] }),
  .B1({ S18992 }),
  .B2({ S18993 }),
  .ZN({ S19103 })
);
NAND3_X1 #() 
NAND3_X1_3023_ (
  .A1({ S18875 }),
  .A2({ S18991 }),
  .A3({ S18872 }),
  .ZN({ S19104 })
);
NAND3_X1 #() 
NAND3_X1_3024_ (
  .A1({ S19103 }),
  .A2({ S15640 }),
  .A3({ S19104 }),
  .ZN({ S19105 })
);
NAND3_X1 #() 
NAND3_X1_3025_ (
  .A1({ S18994 }),
  .A2({ S25957[159] }),
  .A3({ S18990 }),
  .ZN({ S19106 })
);
NAND2_X1 #() 
NAND2_X1_2750_ (
  .A1({ S19105 }),
  .A2({ S19106 }),
  .ZN({ S25957[31] })
);
INV_X1 #() 
INV_X1_854_ (
  .A({ S25956[9] }),
  .ZN({ S5628 })
);
INV_X1 #() 
INV_X1_855_ (
  .A({ S25956[8] }),
  .ZN({ S5639 })
);
NAND2_X1 #() 
NAND2_X1_2751_ (
  .A1({ S5628 }),
  .A2({ S5639 }),
  .ZN({ S27 })
);
NAND2_X1 #() 
NAND2_X1_2752_ (
  .A1({ S25956[9] }),
  .A2({ S25956[8] }),
  .ZN({ S5657 })
);
INV_X1 #() 
INV_X1_856_ (
  .A({ S5657 }),
  .ZN({ S29 })
);
INV_X1 #() 
INV_X1_857_ (
  .A({ S25956[23] }),
  .ZN({ S5675 })
);
INV_X1 #() 
INV_X1_858_ (
  .A({ S25956[15] }),
  .ZN({ S5686 })
);
INV_X1 #() 
INV_X1_859_ (
  .A({ S25956[13] }),
  .ZN({ S5697 })
);
INV_X1 #() 
INV_X1_860_ (
  .A({ S25956[12] }),
  .ZN({ S5708 })
);
INV_X1 #() 
INV_X1_861_ (
  .A({ S25956[11] }),
  .ZN({ S5719 })
);
INV_X1 #() 
INV_X1_862_ (
  .A({ S25956[10] }),
  .ZN({ S5730 })
);
NAND2_X1 #() 
NAND2_X1_2753_ (
  .A1({ S5730 }),
  .A2({ S5639 }),
  .ZN({ S5741 })
);
NAND2_X1 #() 
NAND2_X1_2754_ (
  .A1({ S5741 }),
  .A2({ S25956[9] }),
  .ZN({ S5749 })
);
INV_X1 #() 
INV_X1_863_ (
  .A({ S5749 }),
  .ZN({ S5760 })
);
NAND2_X1 #() 
NAND2_X1_2755_ (
  .A1({ S5730 }),
  .A2({ S25956[9] }),
  .ZN({ S5771 })
);
NAND2_X1 #() 
NAND2_X1_2756_ (
  .A1({ S5741 }),
  .A2({ S5771 }),
  .ZN({ S5782 })
);
NAND2_X1 #() 
NAND2_X1_2757_ (
  .A1({ S5782 }),
  .A2({ S25956[11] }),
  .ZN({ S5793 })
);
NAND2_X1 #() 
NAND2_X1_2758_ (
  .A1({ S25956[11] }),
  .A2({ S25956[10] }),
  .ZN({ S5804 })
);
INV_X1 #() 
INV_X1_864_ (
  .A({ S5804 }),
  .ZN({ S5815 })
);
NAND2_X1 #() 
NAND2_X1_2759_ (
  .A1({ S5815 }),
  .A2({ S25956[8] }),
  .ZN({ S5826 })
);
NAND2_X1 #() 
NAND2_X1_2760_ (
  .A1({ S5793 }),
  .A2({ S5826 }),
  .ZN({ S5837 })
);
AOI21_X1 #() 
AOI21_X1_1524_ (
  .A({ S5837 }),
  .B1({ S5760 }),
  .B2({ S5719 }),
  .ZN({ S5845 })
);
NAND2_X1 #() 
NAND2_X1_2761_ (
  .A1({ S25956[10] }),
  .A2({ S25956[9] }),
  .ZN({ S5856 })
);
INV_X1 #() 
INV_X1_865_ (
  .A({ S5856 }),
  .ZN({ S5867 })
);
NOR2_X1 #() 
NOR2_X1_662_ (
  .A1({ S5719 }),
  .A2({ S25956[8] }),
  .ZN({ S5878 })
);
INV_X1 #() 
INV_X1_866_ (
  .A({ S5878 }),
  .ZN({ S5889 })
);
NOR2_X1 #() 
NOR2_X1_663_ (
  .A1({ S5889 }),
  .A2({ S5867 }),
  .ZN({ S5900 })
);
NAND2_X1 #() 
NAND2_X1_2762_ (
  .A1({ S25956[10] }),
  .A2({ S25956[8] }),
  .ZN({ S5907 })
);
NAND2_X1 #() 
NAND2_X1_2763_ (
  .A1({ S5856 }),
  .A2({ S5907 }),
  .ZN({ S5918 })
);
INV_X1 #() 
INV_X1_867_ (
  .A({ S5918 }),
  .ZN({ S5929 })
);
NAND2_X1 #() 
NAND2_X1_2764_ (
  .A1({ S5657 }),
  .A2({ S5730 }),
  .ZN({ S5940 })
);
AOI21_X1 #() 
AOI21_X1_1525_ (
  .A({ S25956[11] }),
  .B1({ S5929 }),
  .B2({ S5940 }),
  .ZN({ S5951 })
);
AOI211_X1 #() 
AOI211_X1_33_ (
  .A({ S5900 }),
  .B({ S5951 }),
  .C1({ S29 }),
  .C2({ S25956[11] }),
  .ZN({ S5962 })
);
NAND2_X1 #() 
NAND2_X1_2765_ (
  .A1({ S5962 }),
  .A2({ S5708 }),
  .ZN({ S5973 })
);
OAI21_X1 #() 
OAI21_X1_1433_ (
  .A({ S5973 }),
  .B1({ S5708 }),
  .B2({ S5845 }),
  .ZN({ S5984 })
);
NAND2_X1 #() 
NAND2_X1_2766_ (
  .A1({ S5628 }),
  .A2({ S25956[10] }),
  .ZN({ S5995 })
);
INV_X1 #() 
INV_X1_868_ (
  .A({ S5995 }),
  .ZN({ S6006 })
);
NOR2_X1 #() 
NOR2_X1_664_ (
  .A1({ S6006 }),
  .A2({ S5719 }),
  .ZN({ S6015 })
);
NAND2_X1 #() 
NAND2_X1_2767_ (
  .A1({ S6015 }),
  .A2({ S5657 }),
  .ZN({ S6026 })
);
NOR2_X1 #() 
NOR2_X1_665_ (
  .A1({ S5628 }),
  .A2({ S25956[8] }),
  .ZN({ S6037 })
);
NOR2_X1 #() 
NOR2_X1_666_ (
  .A1({ S6037 }),
  .A2({ S25956[11] }),
  .ZN({ S6048 })
);
INV_X1 #() 
INV_X1_869_ (
  .A({ S6048 }),
  .ZN({ S6059 })
);
AOI21_X1 #() 
AOI21_X1_1526_ (
  .A({ S5708 }),
  .B1({ S6026 }),
  .B2({ S6059 }),
  .ZN({ S6070 })
);
NAND2_X1 #() 
NAND2_X1_2768_ (
  .A1({ S5730 }),
  .A2({ S5628 }),
  .ZN({ S6081 })
);
NOR2_X1 #() 
NOR2_X1_667_ (
  .A1({ S5639 }),
  .A2({ S25956[11] }),
  .ZN({ S6092 })
);
OAI211_X1 #() 
OAI211_X1_984_ (
  .A({ S5929 }),
  .B({ S5708 }),
  .C1({ S6081 }),
  .C2({ S6092 }),
  .ZN({ S6101 })
);
NAND2_X1 #() 
NAND2_X1_2769_ (
  .A1({ S6101 }),
  .A2({ S5697 }),
  .ZN({ S6110 })
);
OAI22_X1 #() 
OAI22_X1_68_ (
  .A1({ S5984 }),
  .A2({ S5697 }),
  .B1({ S6070 }),
  .B2({ S6110 }),
  .ZN({ S6121 })
);
INV_X1 #() 
INV_X1_870_ (
  .A({ S25956[14] }),
  .ZN({ S6132 })
);
NAND2_X1 #() 
NAND2_X1_2770_ (
  .A1({ S5628 }),
  .A2({ S25956[11] }),
  .ZN({ S6143 })
);
INV_X1 #() 
INV_X1_871_ (
  .A({ S6143 }),
  .ZN({ S6154 })
);
NAND2_X1 #() 
NAND2_X1_2771_ (
  .A1({ S6154 }),
  .A2({ S5730 }),
  .ZN({ S6165 })
);
INV_X1 #() 
INV_X1_872_ (
  .A({ S6165 }),
  .ZN({ S6176 })
);
NAND2_X1 #() 
NAND2_X1_2772_ (
  .A1({ S5639 }),
  .A2({ S25956[10] }),
  .ZN({ S6184 })
);
NAND2_X1 #() 
NAND2_X1_2773_ (
  .A1({ S6184 }),
  .A2({ S5856 }),
  .ZN({ S6194 })
);
NOR2_X1 #() 
NOR2_X1_668_ (
  .A1({ S25956[9] }),
  .A2({ S25956[8] }),
  .ZN({ S6204 })
);
NOR2_X1 #() 
NOR2_X1_669_ (
  .A1({ S5940 }),
  .A2({ S6204 }),
  .ZN({ S6215 })
);
NOR2_X1 #() 
NOR2_X1_670_ (
  .A1({ S6215 }),
  .A2({ S6194 }),
  .ZN({ S6226 })
);
AOI21_X1 #() 
AOI21_X1_1527_ (
  .A({ S6176 }),
  .B1({ S6226 }),
  .B2({ S5719 }),
  .ZN({ S6237 })
);
NOR2_X1 #() 
NOR2_X1_671_ (
  .A1({ S5639 }),
  .A2({ S25956[10] }),
  .ZN({ S6248 })
);
NOR2_X1 #() 
NOR2_X1_672_ (
  .A1({ S6248 }),
  .A2({ S25956[11] }),
  .ZN({ S6259 })
);
INV_X1 #() 
INV_X1_873_ (
  .A({ S6259 }),
  .ZN({ S6270 })
);
NAND2_X1 #() 
NAND2_X1_2774_ (
  .A1({ S5657 }),
  .A2({ S25956[10] }),
  .ZN({ S6281 })
);
NOR2_X1 #() 
NOR2_X1_673_ (
  .A1({ S6281 }),
  .A2({ S6204 }),
  .ZN({ S6292 })
);
NAND2_X1 #() 
NAND2_X1_2775_ (
  .A1({ S5628 }),
  .A2({ S25956[8] }),
  .ZN({ S6303 })
);
NAND2_X1 #() 
NAND2_X1_2776_ (
  .A1({ S6303 }),
  .A2({ S5730 }),
  .ZN({ S6314 })
);
NOR2_X1 #() 
NOR2_X1_674_ (
  .A1({ S6314 }),
  .A2({ S6037 }),
  .ZN({ S6325 })
);
OAI21_X1 #() 
OAI21_X1_1434_ (
  .A({ S25956[11] }),
  .B1({ S6325 }),
  .B2({ S6292 }),
  .ZN({ S6334 })
);
OAI211_X1 #() 
OAI211_X1_985_ (
  .A({ S6334 }),
  .B({ S25956[12] }),
  .C1({ S5867 }),
  .C2({ S6270 }),
  .ZN({ S6343 })
);
OAI211_X1 #() 
OAI211_X1_986_ (
  .A({ S6343 }),
  .B({ S5697 }),
  .C1({ S6237 }),
  .C2({ S25956[12] }),
  .ZN({ S6354 })
);
AOI21_X1 #() 
AOI21_X1_1528_ (
  .A({ S25956[12] }),
  .B1({ S5741 }),
  .B2({ S5719 }),
  .ZN({ S6365 })
);
OAI21_X1 #() 
OAI21_X1_1435_ (
  .A({ S6365 }),
  .B1({ S5628 }),
  .B2({ S5878 }),
  .ZN({ S6376 })
);
INV_X1 #() 
INV_X1_874_ (
  .A({ S5907 }),
  .ZN({ S6387 })
);
NOR2_X1 #() 
NOR2_X1_675_ (
  .A1({ S5628 }),
  .A2({ S25956[11] }),
  .ZN({ S6398 })
);
INV_X1 #() 
INV_X1_875_ (
  .A({ S6398 }),
  .ZN({ S6409 })
);
NAND2_X1 #() 
NAND2_X1_2777_ (
  .A1({ S5826 }),
  .A2({ S6143 }),
  .ZN({ S6417 })
);
NOR2_X1 #() 
NOR2_X1_676_ (
  .A1({ S6417 }),
  .A2({ S5708 }),
  .ZN({ S6425 })
);
OAI21_X1 #() 
OAI21_X1_1436_ (
  .A({ S6425 }),
  .B1({ S6387 }),
  .B2({ S6409 }),
  .ZN({ S6436 })
);
NAND3_X1 #() 
NAND3_X1_3026_ (
  .A1({ S6436 }),
  .A2({ S25956[13] }),
  .A3({ S6376 }),
  .ZN({ S6447 })
);
AND3_X1 #() 
AND3_X1_118_ (
  .A1({ S6354 }),
  .A2({ S6132 }),
  .A3({ S6447 }),
  .ZN({ S6458 })
);
AOI21_X1 #() 
AOI21_X1_1529_ (
  .A({ S6458 }),
  .B1({ S6121 }),
  .B2({ S25956[14] }),
  .ZN({ S6469 })
);
NAND2_X1 #() 
NAND2_X1_2778_ (
  .A1({ S5907 }),
  .A2({ S25956[11] }),
  .ZN({ S6480 })
);
INV_X1 #() 
INV_X1_876_ (
  .A({ S6480 }),
  .ZN({ S6491 })
);
NAND2_X1 #() 
NAND2_X1_2779_ (
  .A1({ S6491 }),
  .A2({ S5771 }),
  .ZN({ S6502 })
);
NAND2_X1 #() 
NAND2_X1_2780_ (
  .A1({ S6314 }),
  .A2({ S6281 }),
  .ZN({ S6511 })
);
AOI21_X1 #() 
AOI21_X1_1530_ (
  .A({ S25956[12] }),
  .B1({ S6511 }),
  .B2({ S5719 }),
  .ZN({ S6522 })
);
NAND2_X1 #() 
NAND2_X1_2781_ (
  .A1({ S5639 }),
  .A2({ S25956[9] }),
  .ZN({ S6533 })
);
NAND2_X1 #() 
NAND2_X1_2782_ (
  .A1({ S5782 }),
  .A2({ S6533 }),
  .ZN({ S6544 })
);
AOI21_X1 #() 
AOI21_X1_1531_ (
  .A({ S5719 }),
  .B1({ S6544 }),
  .B2({ S6281 }),
  .ZN({ S6555 })
);
INV_X1 #() 
INV_X1_877_ (
  .A({ S6555 }),
  .ZN({ S6566 })
);
INV_X1 #() 
INV_X1_878_ (
  .A({ S6092 }),
  .ZN({ S6576 })
);
NOR2_X1 #() 
NOR2_X1_677_ (
  .A1({ S6576 }),
  .A2({ S5856 }),
  .ZN({ S6583 })
);
NAND2_X1 #() 
NAND2_X1_2783_ (
  .A1({ S5856 }),
  .A2({ S5719 }),
  .ZN({ S6594 })
);
NOR2_X1 #() 
NOR2_X1_678_ (
  .A1({ S6594 }),
  .A2({ S25956[8] }),
  .ZN({ S6605 })
);
NOR3_X1 #() 
NOR3_X1_95_ (
  .A1({ S6583 }),
  .A2({ S6605 }),
  .A3({ S5708 }),
  .ZN({ S6616 })
);
AOI22_X1 #() 
AOI22_X1_325_ (
  .A1({ S6566 }),
  .A2({ S6616 }),
  .B1({ S6522 }),
  .B2({ S6502 }),
  .ZN({ S6627 })
);
INV_X1 #() 
INV_X1_879_ (
  .A({ S6281 }),
  .ZN({ S6638 })
);
NAND2_X1 #() 
NAND2_X1_2784_ (
  .A1({ S6638 }),
  .A2({ S5719 }),
  .ZN({ S6649 })
);
OAI21_X1 #() 
OAI21_X1_1437_ (
  .A({ S25956[11] }),
  .B1({ S5782 }),
  .B2({ S6006 }),
  .ZN({ S6656 })
);
AOI21_X1 #() 
AOI21_X1_1532_ (
  .A({ S25956[12] }),
  .B1({ S6656 }),
  .B2({ S6649 }),
  .ZN({ S6665 })
);
NAND2_X1 #() 
NAND2_X1_2785_ (
  .A1({ S29 }),
  .A2({ S5730 }),
  .ZN({ S6676 })
);
NOR2_X1 #() 
NOR2_X1_679_ (
  .A1({ S5995 }),
  .A2({ S25956[8] }),
  .ZN({ S6687 })
);
INV_X1 #() 
INV_X1_880_ (
  .A({ S6687 }),
  .ZN({ S6698 })
);
NAND2_X1 #() 
NAND2_X1_2786_ (
  .A1({ S6698 }),
  .A2({ S25956[11] }),
  .ZN({ S6709 })
);
INV_X1 #() 
INV_X1_881_ (
  .A({ S6709 }),
  .ZN({ S6720 })
);
NAND2_X1 #() 
NAND2_X1_2787_ (
  .A1({ S6720 }),
  .A2({ S6676 }),
  .ZN({ S6731 })
);
NOR2_X1 #() 
NOR2_X1_680_ (
  .A1({ S5856 }),
  .A2({ S25956[8] }),
  .ZN({ S6742 })
);
NOR2_X1 #() 
NOR2_X1_681_ (
  .A1({ S6742 }),
  .A2({ S25956[11] }),
  .ZN({ S6753 })
);
AOI21_X1 #() 
AOI21_X1_1533_ (
  .A({ S5708 }),
  .B1({ S6753 }),
  .B2({ S5741 }),
  .ZN({ S6763 })
);
AOI21_X1 #() 
AOI21_X1_1534_ (
  .A({ S6665 }),
  .B1({ S6731 }),
  .B2({ S6763 }),
  .ZN({ S6767 })
);
NAND2_X1 #() 
NAND2_X1_2788_ (
  .A1({ S6767 }),
  .A2({ S25956[13] }),
  .ZN({ S6778 })
);
OAI21_X1 #() 
OAI21_X1_1438_ (
  .A({ S6778 }),
  .B1({ S25956[13] }),
  .B2({ S6627 }),
  .ZN({ S6789 })
);
NAND2_X1 #() 
NAND2_X1_2789_ (
  .A1({ S6194 }),
  .A2({ S6533 }),
  .ZN({ S6800 })
);
NAND2_X1 #() 
NAND2_X1_2790_ (
  .A1({ S6800 }),
  .A2({ S5940 }),
  .ZN({ S6811 })
);
NAND2_X1 #() 
NAND2_X1_2791_ (
  .A1({ S6811 }),
  .A2({ S5719 }),
  .ZN({ S6822 })
);
OAI211_X1 #() 
OAI211_X1_987_ (
  .A({ S6822 }),
  .B({ S25956[12] }),
  .C1({ S6742 }),
  .C2({ S5719 }),
  .ZN({ S6832 })
);
INV_X1 #() 
INV_X1_882_ (
  .A({ S6800 }),
  .ZN({ S6838 })
);
NAND2_X1 #() 
NAND2_X1_2792_ (
  .A1({ S6838 }),
  .A2({ S5719 }),
  .ZN({ S6849 })
);
OAI211_X1 #() 
OAI211_X1_988_ (
  .A({ S6849 }),
  .B({ S5708 }),
  .C1({ S6281 }),
  .C2({ S5719 }),
  .ZN({ S6860 })
);
NAND3_X1 #() 
NAND3_X1_3027_ (
  .A1({ S6832 }),
  .A2({ S5697 }),
  .A3({ S6860 }),
  .ZN({ S6871 })
);
INV_X1 #() 
INV_X1_883_ (
  .A({ S6594 }),
  .ZN({ S6882 })
);
AOI21_X1 #() 
AOI21_X1_1535_ (
  .A({ S5719 }),
  .B1({ S27 }),
  .B2({ S5856 }),
  .ZN({ S6893 })
);
AOI21_X1 #() 
AOI21_X1_1536_ (
  .A({ S6893 }),
  .B1({ S6882 }),
  .B2({ S5940 }),
  .ZN({ S6904 })
);
NAND2_X1 #() 
NAND2_X1_2793_ (
  .A1({ S6491 }),
  .A2({ S6081 }),
  .ZN({ S6912 })
);
NAND3_X1 #() 
NAND3_X1_3028_ (
  .A1({ S6912 }),
  .A2({ S25956[12] }),
  .A3({ S6576 }),
  .ZN({ S6923 })
);
OAI211_X1 #() 
OAI211_X1_989_ (
  .A({ S6923 }),
  .B({ S25956[13] }),
  .C1({ S6904 }),
  .C2({ S25956[12] }),
  .ZN({ S6934 })
);
NAND3_X1 #() 
NAND3_X1_3029_ (
  .A1({ S6871 }),
  .A2({ S6132 }),
  .A3({ S6934 }),
  .ZN({ S6945 })
);
OAI211_X1 #() 
OAI211_X1_990_ (
  .A({ S6945 }),
  .B({ S5686 }),
  .C1({ S6789 }),
  .C2({ S6132 }),
  .ZN({ S6956 })
);
OAI21_X1 #() 
OAI21_X1_1439_ (
  .A({ S6956 }),
  .B1({ S6469 }),
  .B2({ S5686 }),
  .ZN({ S6967 })
);
XNOR2_X1 #() 
XNOR2_X1_151_ (
  .A({ S6967 }),
  .B({ S25956[119] }),
  .ZN({ S6978 })
);
XOR2_X1 #() 
XOR2_X1_63_ (
  .A({ S6978 }),
  .B({ S25956[87] }),
  .Z({ S6989 })
);
XNOR2_X1 #() 
XNOR2_X1_152_ (
  .A({ S6989 }),
  .B({ S25956[55] }),
  .ZN({ S25957[1207] })
);
XNOR2_X1 #() 
XNOR2_X1_153_ (
  .A({ S25957[1207] }),
  .B({ S5675 }),
  .ZN({ S25957[1175] })
);
NOR2_X1 #() 
NOR2_X1_682_ (
  .A1({ S6248 }),
  .A2({ S6143 }),
  .ZN({ S7020 })
);
NAND2_X1 #() 
NAND2_X1_2794_ (
  .A1({ S7020 }),
  .A2({ S6184 }),
  .ZN({ S7030 })
);
OAI211_X1 #() 
OAI211_X1_991_ (
  .A({ S7030 }),
  .B({ S25956[12] }),
  .C1({ S5929 }),
  .C2({ S25956[11] }),
  .ZN({ S7041 })
);
NAND2_X1 #() 
NAND2_X1_2795_ (
  .A1({ S6026 }),
  .A2({ S6409 }),
  .ZN({ S7052 })
);
AOI21_X1 #() 
AOI21_X1_1537_ (
  .A({ S5697 }),
  .B1({ S7052 }),
  .B2({ S5708 }),
  .ZN({ S7063 })
);
INV_X1 #() 
INV_X1_884_ (
  .A({ S5940 }),
  .ZN({ S7074 })
);
OAI21_X1 #() 
OAI21_X1_1440_ (
  .A({ S6522 }),
  .B1({ S7074 }),
  .B2({ S6709 }),
  .ZN({ S7085 })
);
OAI21_X1 #() 
OAI21_X1_1441_ (
  .A({ S5719 }),
  .B1({ S6215 }),
  .B2({ S6387 }),
  .ZN({ S7096 })
);
OAI21_X1 #() 
OAI21_X1_1442_ (
  .A({ S25956[11] }),
  .B1({ S6194 }),
  .B2({ S6248 }),
  .ZN({ S7107 })
);
AND2_X1 #() 
AND2_X1_177_ (
  .A1({ S7107 }),
  .A2({ S25956[12] }),
  .ZN({ S7113 })
);
NAND2_X1 #() 
NAND2_X1_2796_ (
  .A1({ S7113 }),
  .A2({ S7096 }),
  .ZN({ S7124 })
);
AOI21_X1 #() 
AOI21_X1_1538_ (
  .A({ S25956[13] }),
  .B1({ S7124 }),
  .B2({ S7085 }),
  .ZN({ S7135 })
);
AOI21_X1 #() 
AOI21_X1_1539_ (
  .A({ S7135 }),
  .B1({ S7063 }),
  .B2({ S7041 }),
  .ZN({ S7146 })
);
NAND2_X1 #() 
NAND2_X1_2797_ (
  .A1({ S27 }),
  .A2({ S5741 }),
  .ZN({ S7157 })
);
OAI21_X1 #() 
OAI21_X1_1443_ (
  .A({ S7096 }),
  .B1({ S7157 }),
  .B2({ S6480 }),
  .ZN({ S7168 })
);
NOR2_X1 #() 
NOR2_X1_683_ (
  .A1({ S7168 }),
  .A2({ S25956[12] }),
  .ZN({ S7179 })
);
AOI21_X1 #() 
AOI21_X1_1540_ (
  .A({ S6417 }),
  .B1({ S5782 }),
  .B2({ S5719 }),
  .ZN({ S7190 })
);
OAI21_X1 #() 
OAI21_X1_1444_ (
  .A({ S5697 }),
  .B1({ S7190 }),
  .B2({ S5708 }),
  .ZN({ S7201 })
);
NAND2_X1 #() 
NAND2_X1_2798_ (
  .A1({ S5730 }),
  .A2({ S25956[8] }),
  .ZN({ S7210 })
);
NAND2_X1 #() 
NAND2_X1_2799_ (
  .A1({ S6081 }),
  .A2({ S7210 }),
  .ZN({ S7221 })
);
INV_X1 #() 
INV_X1_885_ (
  .A({ S7221 }),
  .ZN({ S7232 })
);
OAI21_X1 #() 
OAI21_X1_1445_ (
  .A({ S5719 }),
  .B1({ S6281 }),
  .B2({ S6204 }),
  .ZN({ S7243 })
);
INV_X1 #() 
INV_X1_886_ (
  .A({ S7243 }),
  .ZN({ S7254 })
);
NAND2_X1 #() 
NAND2_X1_2800_ (
  .A1({ S7254 }),
  .A2({ S7232 }),
  .ZN({ S7265 })
);
NOR2_X1 #() 
NOR2_X1_684_ (
  .A1({ S5856 }),
  .A2({ S5719 }),
  .ZN({ S7275 })
);
NOR2_X1 #() 
NOR2_X1_685_ (
  .A1({ S7275 }),
  .A2({ S5708 }),
  .ZN({ S7286 })
);
INV_X1 #() 
INV_X1_887_ (
  .A({ S6015 }),
  .ZN({ S7297 })
);
NAND2_X1 #() 
NAND2_X1_2801_ (
  .A1({ S6037 }),
  .A2({ S5730 }),
  .ZN({ S7308 })
);
INV_X1 #() 
INV_X1_888_ (
  .A({ S7308 }),
  .ZN({ S7319 })
);
NOR2_X1 #() 
NOR2_X1_686_ (
  .A1({ S5907 }),
  .A2({ S5628 }),
  .ZN({ S7330 })
);
NOR2_X1 #() 
NOR2_X1_687_ (
  .A1({ S7330 }),
  .A2({ S6204 }),
  .ZN({ S7339 })
);
OAI22_X1 #() 
OAI22_X1_69_ (
  .A1({ S7297 }),
  .A2({ S7319 }),
  .B1({ S7339 }),
  .B2({ S25956[11] }),
  .ZN({ S7350 })
);
AOI22_X1 #() 
AOI22_X1_326_ (
  .A1({ S7350 }),
  .A2({ S5708 }),
  .B1({ S7265 }),
  .B2({ S7286 }),
  .ZN({ S7361 })
);
NAND2_X1 #() 
NAND2_X1_2802_ (
  .A1({ S7361 }),
  .A2({ S25956[13] }),
  .ZN({ S7372 })
);
OAI211_X1 #() 
OAI211_X1_992_ (
  .A({ S7372 }),
  .B({ S6132 }),
  .C1({ S7179 }),
  .C2({ S7201 }),
  .ZN({ S7383 })
);
OAI21_X1 #() 
OAI21_X1_1446_ (
  .A({ S7383 }),
  .B1({ S7146 }),
  .B2({ S6132 }),
  .ZN({ S7391 })
);
NOR2_X1 #() 
NOR2_X1_688_ (
  .A1({ S6638 }),
  .A2({ S6248 }),
  .ZN({ S7402 })
);
NOR2_X1 #() 
NOR2_X1_689_ (
  .A1({ S7402 }),
  .A2({ S25956[11] }),
  .ZN({ S7413 })
);
AOI211_X1 #() 
AOI211_X1_34_ (
  .A({ S5708 }),
  .B({ S7413 }),
  .C1({ S6533 }),
  .C2({ S6491 }),
  .ZN({ S7424 })
);
NAND2_X1 #() 
NAND2_X1_2803_ (
  .A1({ S6081 }),
  .A2({ S5639 }),
  .ZN({ S7435 })
);
NOR2_X1 #() 
NOR2_X1_690_ (
  .A1({ S7435 }),
  .A2({ S25956[11] }),
  .ZN({ S7446 })
);
NOR2_X1 #() 
NOR2_X1_691_ (
  .A1({ S5628 }),
  .A2({ S25956[10] }),
  .ZN({ S7457 })
);
NAND2_X1 #() 
NAND2_X1_2804_ (
  .A1({ S7457 }),
  .A2({ S25956[11] }),
  .ZN({ S7468 })
);
NAND2_X1 #() 
NAND2_X1_2805_ (
  .A1({ S7468 }),
  .A2({ S25956[12] }),
  .ZN({ S7475 })
);
NAND3_X1 #() 
NAND3_X1_3030_ (
  .A1({ S7107 }),
  .A2({ S7243 }),
  .A3({ S5708 }),
  .ZN({ S7486 })
);
OAI211_X1 #() 
OAI211_X1_993_ (
  .A({ S7486 }),
  .B({ S5697 }),
  .C1({ S7446 }),
  .C2({ S7475 }),
  .ZN({ S7497 })
);
NAND2_X1 #() 
NAND2_X1_2806_ (
  .A1({ S7210 }),
  .A2({ S25956[9] }),
  .ZN({ S7508 })
);
AOI22_X1 #() 
AOI22_X1_327_ (
  .A1({ S6491 }),
  .A2({ S6533 }),
  .B1({ S7508 }),
  .B2({ S5719 }),
  .ZN({ S7519 })
);
OAI21_X1 #() 
OAI21_X1_1447_ (
  .A({ S25956[13] }),
  .B1({ S7519 }),
  .B2({ S25956[12] }),
  .ZN({ S7530 })
);
OAI211_X1 #() 
OAI211_X1_994_ (
  .A({ S7497 }),
  .B({ S25956[14] }),
  .C1({ S7424 }),
  .C2({ S7530 }),
  .ZN({ S7541 })
);
NAND3_X1 #() 
NAND3_X1_3031_ (
  .A1({ S6184 }),
  .A2({ S25956[11] }),
  .A3({ S5657 }),
  .ZN({ S7552 })
);
NOR2_X1 #() 
NOR2_X1_692_ (
  .A1({ S6533 }),
  .A2({ S5719 }),
  .ZN({ S7560 })
);
INV_X1 #() 
INV_X1_889_ (
  .A({ S7560 }),
  .ZN({ S7570 })
);
NAND4_X1 #() 
NAND4_X1_341_ (
  .A1({ S6270 }),
  .A2({ S7570 }),
  .A3({ S25956[12] }),
  .A4({ S7552 }),
  .ZN({ S7581 })
);
AOI21_X1 #() 
AOI21_X1_1541_ (
  .A({ S6594 }),
  .B1({ S6248 }),
  .B2({ S5628 }),
  .ZN({ S7592 })
);
OAI21_X1 #() 
OAI21_X1_1448_ (
  .A({ S5708 }),
  .B1({ S7297 }),
  .B2({ S7457 }),
  .ZN({ S7603 })
);
OAI21_X1 #() 
OAI21_X1_1449_ (
  .A({ S7581 }),
  .B1({ S7603 }),
  .B2({ S7592 }),
  .ZN({ S7614 })
);
OAI21_X1 #() 
OAI21_X1_1450_ (
  .A({ S6081 }),
  .B1({ S5749 }),
  .B2({ S6387 }),
  .ZN({ S7625 })
);
AOI21_X1 #() 
AOI21_X1_1542_ (
  .A({ S25956[12] }),
  .B1({ S7625 }),
  .B2({ S25956[11] }),
  .ZN({ S7636 })
);
INV_X1 #() 
INV_X1_890_ (
  .A({ S7636 }),
  .ZN({ S7647 })
);
OAI211_X1 #() 
OAI211_X1_995_ (
  .A({ S6656 }),
  .B({ S25956[12] }),
  .C1({ S6081 }),
  .C2({ S6576 }),
  .ZN({ S7658 })
);
NAND3_X1 #() 
NAND3_X1_3032_ (
  .A1({ S7647 }),
  .A2({ S5697 }),
  .A3({ S7658 }),
  .ZN({ S7669 })
);
OAI21_X1 #() 
OAI21_X1_1451_ (
  .A({ S7669 }),
  .B1({ S7614 }),
  .B2({ S5697 }),
  .ZN({ S7680 })
);
OAI21_X1 #() 
OAI21_X1_1452_ (
  .A({ S7541 }),
  .B1({ S7680 }),
  .B2({ S25956[14] }),
  .ZN({ S7691 })
);
MUX2_X1 #() 
MUX2_X1_8_ (
  .A({ S7691 }),
  .B({ S7391 }),
  .S({ S25956[15] }),
  .Z({ S7702 })
);
XOR2_X1 #() 
XOR2_X1_64_ (
  .A({ S7702 }),
  .B({ S25956[118] }),
  .Z({ S25957[1270] })
);
XOR2_X1 #() 
XOR2_X1_65_ (
  .A({ S25957[1270] }),
  .B({ S25956[86] }),
  .Z({ S25957[1238] })
);
XOR2_X1 #() 
XOR2_X1_66_ (
  .A({ S25957[1238] }),
  .B({ S25956[54] }),
  .Z({ S25957[1206] })
);
XNOR2_X1 #() 
XNOR2_X1_154_ (
  .A({ S25957[1206] }),
  .B({ S25956[22] }),
  .ZN({ S7741 })
);
INV_X1 #() 
INV_X1_891_ (
  .A({ S7741 }),
  .ZN({ S25957[1174] })
);
INV_X1 #() 
INV_X1_892_ (
  .A({ S25956[21] }),
  .ZN({ S7762 })
);
INV_X1 #() 
INV_X1_893_ (
  .A({ S25956[85] }),
  .ZN({ S7773 })
);
NOR2_X1 #() 
NOR2_X1_693_ (
  .A1({ S6059 }),
  .A2({ S6248 }),
  .ZN({ S7782 })
);
OAI21_X1 #() 
OAI21_X1_1453_ (
  .A({ S5708 }),
  .B1({ S7782 }),
  .B2({ S5878 }),
  .ZN({ S7789 })
);
AOI21_X1 #() 
AOI21_X1_1543_ (
  .A({ S5719 }),
  .B1({ S6800 }),
  .B2({ S7308 }),
  .ZN({ S7800 })
);
OAI21_X1 #() 
OAI21_X1_1454_ (
  .A({ S25956[12] }),
  .B1({ S7800 }),
  .B2({ S7592 }),
  .ZN({ S7811 })
);
NAND3_X1 #() 
NAND3_X1_3033_ (
  .A1({ S7811 }),
  .A2({ S7789 }),
  .A3({ S25956[13] }),
  .ZN({ S7822 })
);
INV_X1 #() 
INV_X1_894_ (
  .A({ S5793 }),
  .ZN({ S7833 })
);
NOR2_X1 #() 
NOR2_X1_694_ (
  .A1({ S7833 }),
  .A2({ S5708 }),
  .ZN({ S7844 })
);
INV_X1 #() 
INV_X1_895_ (
  .A({ S7330 }),
  .ZN({ S7855 })
);
NAND3_X1 #() 
NAND3_X1_3034_ (
  .A1({ S7855 }),
  .A2({ S5719 }),
  .A3({ S5940 }),
  .ZN({ S7866 })
);
NAND3_X1 #() 
NAND3_X1_3035_ (
  .A1({ S7308 }),
  .A2({ S5719 }),
  .A3({ S5907 }),
  .ZN({ S7876 })
);
NAND2_X1 #() 
NAND2_X1_2807_ (
  .A1({ S7402 }),
  .A2({ S25956[11] }),
  .ZN({ S7882 })
);
AOI21_X1 #() 
AOI21_X1_1544_ (
  .A({ S25956[12] }),
  .B1({ S7882 }),
  .B2({ S7876 }),
  .ZN({ S7893 })
);
AOI21_X1 #() 
AOI21_X1_1545_ (
  .A({ S7893 }),
  .B1({ S7866 }),
  .B2({ S7844 }),
  .ZN({ S7904 })
);
AOI21_X1 #() 
AOI21_X1_1546_ (
  .A({ S6132 }),
  .B1({ S7904 }),
  .B2({ S5697 }),
  .ZN({ S7915 })
);
NAND2_X1 #() 
NAND2_X1_2808_ (
  .A1({ S6292 }),
  .A2({ S25956[11] }),
  .ZN({ S7926 })
);
NAND3_X1 #() 
NAND3_X1_3036_ (
  .A1({ S6048 }),
  .A2({ S5741 }),
  .A3({ S6303 }),
  .ZN({ S7937 })
);
NAND3_X1 #() 
NAND3_X1_3037_ (
  .A1({ S7844 }),
  .A2({ S7926 }),
  .A3({ S7937 }),
  .ZN({ S7948 })
);
NOR2_X1 #() 
NOR2_X1_695_ (
  .A1({ S6303 }),
  .A2({ S5719 }),
  .ZN({ S7959 })
);
OAI21_X1 #() 
OAI21_X1_1455_ (
  .A({ S5708 }),
  .B1({ S6583 }),
  .B2({ S7959 }),
  .ZN({ S7966 })
);
NAND3_X1 #() 
NAND3_X1_3038_ (
  .A1({ S7948 }),
  .A2({ S5697 }),
  .A3({ S7966 }),
  .ZN({ S7974 })
);
NAND2_X1 #() 
NAND2_X1_2809_ (
  .A1({ S5719 }),
  .A2({ S5730 }),
  .ZN({ S7985 })
);
NOR2_X1 #() 
NOR2_X1_696_ (
  .A1({ S7985 }),
  .A2({ S6533 }),
  .ZN({ S7996 })
);
INV_X1 #() 
INV_X1_896_ (
  .A({ S7996 }),
  .ZN({ S8007 })
);
OAI211_X1 #() 
OAI211_X1_996_ (
  .A({ S8007 }),
  .B({ S25956[12] }),
  .C1({ S7074 }),
  .C2({ S5719 }),
  .ZN({ S8018 })
);
NAND2_X1 #() 
NAND2_X1_2810_ (
  .A1({ S7855 }),
  .A2({ S7308 }),
  .ZN({ S8029 })
);
OAI211_X1 #() 
OAI211_X1_997_ (
  .A({ S5708 }),
  .B({ S6480 }),
  .C1({ S8029 }),
  .C2({ S25956[11] }),
  .ZN({ S8040 })
);
NAND3_X1 #() 
NAND3_X1_3039_ (
  .A1({ S8040 }),
  .A2({ S25956[13] }),
  .A3({ S8018 }),
  .ZN({ S8051 })
);
AND2_X1 #() 
AND2_X1_178_ (
  .A1({ S8051 }),
  .A2({ S6132 }),
  .ZN({ S8062 })
);
AOI22_X1 #() 
AOI22_X1_328_ (
  .A1({ S7915 }),
  .A2({ S7822 }),
  .B1({ S8062 }),
  .B2({ S7974 }),
  .ZN({ S8070 })
);
NAND2_X1 #() 
NAND2_X1_2811_ (
  .A1({ S6676 }),
  .A2({ S5719 }),
  .ZN({ S8080 })
);
NOR2_X1 #() 
NOR2_X1_697_ (
  .A1({ S6081 }),
  .A2({ S25956[8] }),
  .ZN({ S8091 })
);
OAI21_X1 #() 
OAI21_X1_1456_ (
  .A({ S25956[11] }),
  .B1({ S6292 }),
  .B2({ S8091 }),
  .ZN({ S8102 })
);
AOI21_X1 #() 
AOI21_X1_1547_ (
  .A({ S25956[12] }),
  .B1({ S8102 }),
  .B2({ S8080 }),
  .ZN({ S8113 })
);
OAI21_X1 #() 
OAI21_X1_1457_ (
  .A({ S25956[12] }),
  .B1({ S6270 }),
  .B2({ S25956[9] }),
  .ZN({ S8124 })
);
AOI21_X1 #() 
AOI21_X1_1548_ (
  .A({ S8124 }),
  .B1({ S6215 }),
  .B2({ S25956[11] }),
  .ZN({ S8133 })
);
OAI21_X1 #() 
OAI21_X1_1458_ (
  .A({ S5697 }),
  .B1({ S8133 }),
  .B2({ S8113 }),
  .ZN({ S8142 })
);
NAND3_X1 #() 
NAND3_X1_3040_ (
  .A1({ S5741 }),
  .A2({ S5719 }),
  .A3({ S5657 }),
  .ZN({ S8153 })
);
OAI21_X1 #() 
OAI21_X1_1459_ (
  .A({ S8153 }),
  .B1({ S6511 }),
  .B2({ S5719 }),
  .ZN({ S8164 })
);
NAND2_X1 #() 
NAND2_X1_2812_ (
  .A1({ S6048 }),
  .A2({ S6081 }),
  .ZN({ S8175 })
);
AOI21_X1 #() 
AOI21_X1_1549_ (
  .A({ S25956[12] }),
  .B1({ S8175 }),
  .B2({ S6143 }),
  .ZN({ S8186 })
);
AOI21_X1 #() 
AOI21_X1_1550_ (
  .A({ S8186 }),
  .B1({ S8164 }),
  .B2({ S25956[12] }),
  .ZN({ S8197 })
);
OAI21_X1 #() 
OAI21_X1_1460_ (
  .A({ S8142 }),
  .B1({ S5697 }),
  .B2({ S8197 }),
  .ZN({ S8205 })
);
AOI22_X1 #() 
AOI22_X1_329_ (
  .A1({ S6048 }),
  .A2({ S6314 }),
  .B1({ S6081 }),
  .B2({ S5878 }),
  .ZN({ S8216 })
);
NOR2_X1 #() 
NOR2_X1_698_ (
  .A1({ S5760 }),
  .A2({ S5719 }),
  .ZN({ S8227 })
);
NAND3_X1 #() 
NAND3_X1_3041_ (
  .A1({ S6409 }),
  .A2({ S5708 }),
  .A3({ S5907 }),
  .ZN({ S8238 })
);
OAI221_X1 #() 
OAI221_X1_71_ (
  .A({ S25956[13] }),
  .B1({ S8216 }),
  .B2({ S5708 }),
  .C1({ S8238 }),
  .C2({ S8227 }),
  .ZN({ S8249 })
);
NAND3_X1 #() 
NAND3_X1_3042_ (
  .A1({ S6849 }),
  .A2({ S5708 }),
  .A3({ S7107 }),
  .ZN({ S8260 })
);
NAND2_X1 #() 
NAND2_X1_2813_ (
  .A1({ S5995 }),
  .A2({ S5907 }),
  .ZN({ S8271 })
);
INV_X1 #() 
INV_X1_897_ (
  .A({ S8271 }),
  .ZN({ S8282 })
);
NAND3_X1 #() 
NAND3_X1_3043_ (
  .A1({ S7570 }),
  .A2({ S25956[12] }),
  .A3({ S8282 }),
  .ZN({ S8292 })
);
NAND3_X1 #() 
NAND3_X1_3044_ (
  .A1({ S8260 }),
  .A2({ S5697 }),
  .A3({ S8292 }),
  .ZN({ S8301 })
);
NAND3_X1 #() 
NAND3_X1_3045_ (
  .A1({ S8301 }),
  .A2({ S25956[14] }),
  .A3({ S8249 }),
  .ZN({ S8312 })
);
OAI211_X1 #() 
OAI211_X1_998_ (
  .A({ S8312 }),
  .B({ S25956[15] }),
  .C1({ S8205 }),
  .C2({ S25956[14] }),
  .ZN({ S8323 })
);
OAI21_X1 #() 
OAI21_X1_1461_ (
  .A({ S8323 }),
  .B1({ S8070 }),
  .B2({ S25956[15] }),
  .ZN({ S8334 })
);
XNOR2_X1 #() 
XNOR2_X1_155_ (
  .A({ S8334 }),
  .B({ S25956[117] }),
  .ZN({ S25957[1269] })
);
XNOR2_X1 #() 
XNOR2_X1_156_ (
  .A({ S25957[1269] }),
  .B({ S7773 }),
  .ZN({ S25957[1237] })
);
XOR2_X1 #() 
XOR2_X1_67_ (
  .A({ S25957[1237] }),
  .B({ S25956[53] }),
  .Z({ S25957[1205] })
);
XNOR2_X1 #() 
XNOR2_X1_157_ (
  .A({ S25957[1205] }),
  .B({ S7762 }),
  .ZN({ S25957[1173] })
);
INV_X1 #() 
INV_X1_898_ (
  .A({ S25956[20] }),
  .ZN({ S8385 })
);
INV_X1 #() 
INV_X1_899_ (
  .A({ S25956[84] }),
  .ZN({ S8396 })
);
INV_X1 #() 
INV_X1_900_ (
  .A({ S25956[116] }),
  .ZN({ S8407 })
);
NAND2_X1 #() 
NAND2_X1_2814_ (
  .A1({ S6154 }),
  .A2({ S5907 }),
  .ZN({ S8418 })
);
INV_X1 #() 
INV_X1_901_ (
  .A({ S8418 }),
  .ZN({ S8427 })
);
NAND2_X1 #() 
NAND2_X1_2815_ (
  .A1({ S8282 }),
  .A2({ S5719 }),
  .ZN({ S8437 })
);
OAI21_X1 #() 
OAI21_X1_1462_ (
  .A({ S5708 }),
  .B1({ S8437 }),
  .B2({ S7319 }),
  .ZN({ S8448 })
);
OAI21_X1 #() 
OAI21_X1_1463_ (
  .A({ S5719 }),
  .B1({ S5749 }),
  .B2({ S6387 }),
  .ZN({ S8459 })
);
OAI21_X1 #() 
OAI21_X1_1464_ (
  .A({ S8459 }),
  .B1({ S6006 }),
  .B2({ S6502 }),
  .ZN({ S8470 })
);
OAI22_X1 #() 
OAI22_X1_70_ (
  .A1({ S8448 }),
  .A2({ S8427 }),
  .B1({ S8470 }),
  .B2({ S5708 }),
  .ZN({ S8481 })
);
OAI21_X1 #() 
OAI21_X1_1465_ (
  .A({ S5719 }),
  .B1({ S6325 }),
  .B2({ S6638 }),
  .ZN({ S8492 })
);
NOR2_X1 #() 
NOR2_X1_699_ (
  .A1({ S7833 }),
  .A2({ S7560 }),
  .ZN({ S8503 })
);
AOI21_X1 #() 
AOI21_X1_1551_ (
  .A({ S25956[12] }),
  .B1({ S8503 }),
  .B2({ S8492 }),
  .ZN({ S8510 })
);
INV_X1 #() 
INV_X1_902_ (
  .A({ S6303 }),
  .ZN({ S8521 })
);
AOI211_X1 #() 
AOI211_X1_35_ (
  .A({ S5708 }),
  .B({ S7319 }),
  .C1({ S8521 }),
  .C2({ S7985 }),
  .ZN({ S8532 })
);
OAI21_X1 #() 
OAI21_X1_1466_ (
  .A({ S25956[13] }),
  .B1({ S8510 }),
  .B2({ S8532 }),
  .ZN({ S8543 })
);
OAI211_X1 #() 
OAI211_X1_999_ (
  .A({ S8543 }),
  .B({ S6132 }),
  .C1({ S8481 }),
  .C2({ S25956[13] }),
  .ZN({ S8554 })
);
NAND2_X1 #() 
NAND2_X1_2816_ (
  .A1({ S8175 }),
  .A2({ S25956[12] }),
  .ZN({ S8565 })
);
INV_X1 #() 
INV_X1_903_ (
  .A({ S6893 }),
  .ZN({ S8576 })
);
NAND3_X1 #() 
NAND3_X1_3046_ (
  .A1({ S6081 }),
  .A2({ S6184 }),
  .A3({ S5719 }),
  .ZN({ S8586 })
);
NAND3_X1 #() 
NAND3_X1_3047_ (
  .A1({ S8576 }),
  .A2({ S8586 }),
  .A3({ S5708 }),
  .ZN({ S8594 })
);
OAI21_X1 #() 
OAI21_X1_1467_ (
  .A({ S8594 }),
  .B1({ S8565 }),
  .B2({ S7020 }),
  .ZN({ S8605 })
);
NOR2_X1 #() 
NOR2_X1_700_ (
  .A1({ S6687 }),
  .A2({ S25956[11] }),
  .ZN({ S8616 })
);
INV_X1 #() 
INV_X1_904_ (
  .A({ S8616 }),
  .ZN({ S8627 })
);
NAND2_X1 #() 
NAND2_X1_2817_ (
  .A1({ S7844 }),
  .A2({ S8627 }),
  .ZN({ S8638 })
);
NOR2_X1 #() 
NOR2_X1_701_ (
  .A1({ S7457 }),
  .A2({ S25956[11] }),
  .ZN({ S8649 })
);
NAND2_X1 #() 
NAND2_X1_2818_ (
  .A1({ S8649 }),
  .A2({ S5639 }),
  .ZN({ S8660 })
);
NAND3_X1 #() 
NAND3_X1_3048_ (
  .A1({ S8660 }),
  .A2({ S5708 }),
  .A3({ S6912 }),
  .ZN({ S8671 })
);
NAND3_X1 #() 
NAND3_X1_3049_ (
  .A1({ S8638 }),
  .A2({ S25956[13] }),
  .A3({ S8671 }),
  .ZN({ S8682 })
);
OAI21_X1 #() 
OAI21_X1_1468_ (
  .A({ S8682 }),
  .B1({ S25956[13] }),
  .B2({ S8605 }),
  .ZN({ S8687 })
);
OAI21_X1 #() 
OAI21_X1_1469_ (
  .A({ S8554 }),
  .B1({ S6132 }),
  .B2({ S8687 }),
  .ZN({ S8698 })
);
NAND2_X1 #() 
NAND2_X1_2819_ (
  .A1({ S8698 }),
  .A2({ S25956[15] }),
  .ZN({ S8709 })
);
NAND3_X1 #() 
NAND3_X1_3050_ (
  .A1({ S6676 }),
  .A2({ S5719 }),
  .A3({ S6184 }),
  .ZN({ S8720 })
);
NOR2_X1 #() 
NOR2_X1_702_ (
  .A1({ S5815 }),
  .A2({ S25956[12] }),
  .ZN({ S8731 })
);
NOR2_X1 #() 
NOR2_X1_703_ (
  .A1({ S6594 }),
  .A2({ S6387 }),
  .ZN({ S8742 })
);
NAND2_X1 #() 
NAND2_X1_2820_ (
  .A1({ S8742 }),
  .A2({ S6081 }),
  .ZN({ S8753 })
);
AOI22_X1 #() 
AOI22_X1_330_ (
  .A1({ S6425 }),
  .A2({ S8753 }),
  .B1({ S8720 }),
  .B2({ S8731 }),
  .ZN({ S8763 })
);
NOR2_X1 #() 
NOR2_X1_704_ (
  .A1({ S6215 }),
  .A2({ S8271 }),
  .ZN({ S8770 })
);
OAI211_X1 #() 
OAI211_X1_1000_ (
  .A({ S7882 }),
  .B({ S5708 }),
  .C1({ S25956[11] }),
  .C2({ S8770 }),
  .ZN({ S8781 })
);
NAND2_X1 #() 
NAND2_X1_2821_ (
  .A1({ S5730 }),
  .A2({ S116 }),
  .ZN({ S8792 })
);
AOI21_X1 #() 
AOI21_X1_1552_ (
  .A({ S5697 }),
  .B1({ S8792 }),
  .B2({ S25956[12] }),
  .ZN({ S8803 })
);
AOI22_X1 #() 
AOI22_X1_331_ (
  .A1({ S8781 }),
  .A2({ S8803 }),
  .B1({ S8763 }),
  .B2({ S5697 }),
  .ZN({ S8814 })
);
NAND3_X1 #() 
NAND3_X1_3051_ (
  .A1({ S8437 }),
  .A2({ S6656 }),
  .A3({ S25956[12] }),
  .ZN({ S8825 })
);
MUX2_X1 #() 
MUX2_X1_9_ (
  .A({ S29 }),
  .B({ S6215 }),
  .S({ S25956[11] }),
  .Z({ S8836 })
);
OAI21_X1 #() 
OAI21_X1_1470_ (
  .A({ S8825 }),
  .B1({ S8836 }),
  .B2({ S25956[12] }),
  .ZN({ S8844 })
);
NAND3_X1 #() 
NAND3_X1_3052_ (
  .A1({ S8616 }),
  .A2({ S7210 }),
  .A3({ S5771 }),
  .ZN({ S8854 })
);
NOR2_X1 #() 
NOR2_X1_705_ (
  .A1({ S6480 }),
  .A2({ S6204 }),
  .ZN({ S8865 })
);
INV_X1 #() 
INV_X1_905_ (
  .A({ S8865 }),
  .ZN({ S8876 })
);
AOI21_X1 #() 
AOI21_X1_1553_ (
  .A({ S25956[12] }),
  .B1({ S8854 }),
  .B2({ S8876 }),
  .ZN({ S8887 })
);
AOI21_X1 #() 
AOI21_X1_1554_ (
  .A({ S8565 }),
  .B1({ S6491 }),
  .B2({ S6314 }),
  .ZN({ S8898 })
);
OAI21_X1 #() 
OAI21_X1_1471_ (
  .A({ S5697 }),
  .B1({ S8898 }),
  .B2({ S8887 }),
  .ZN({ S8909 })
);
OAI21_X1 #() 
OAI21_X1_1472_ (
  .A({ S8909 }),
  .B1({ S5697 }),
  .B2({ S8844 }),
  .ZN({ S8919 })
);
NAND2_X1 #() 
NAND2_X1_2822_ (
  .A1({ S8919 }),
  .A2({ S6132 }),
  .ZN({ S8930 })
);
OAI211_X1 #() 
OAI211_X1_1001_ (
  .A({ S8930 }),
  .B({ S5686 }),
  .C1({ S8814 }),
  .C2({ S6132 }),
  .ZN({ S8941 })
);
NAND2_X1 #() 
NAND2_X1_2823_ (
  .A1({ S8709 }),
  .A2({ S8941 }),
  .ZN({ S8948 })
);
NAND2_X1 #() 
NAND2_X1_2824_ (
  .A1({ S8948 }),
  .A2({ S8407 }),
  .ZN({ S8959 })
);
NAND3_X1 #() 
NAND3_X1_3053_ (
  .A1({ S8709 }),
  .A2({ S8941 }),
  .A3({ S25956[116] }),
  .ZN({ S8970 })
);
NAND2_X1 #() 
NAND2_X1_2825_ (
  .A1({ S8959 }),
  .A2({ S8970 }),
  .ZN({ S25957[1268] })
);
NAND2_X1 #() 
NAND2_X1_2826_ (
  .A1({ S25957[1268] }),
  .A2({ S8396 }),
  .ZN({ S8991 })
);
INV_X1 #() 
INV_X1_906_ (
  .A({ S25957[1268] }),
  .ZN({ S9002 })
);
NAND2_X1 #() 
NAND2_X1_2827_ (
  .A1({ S9002 }),
  .A2({ S25956[84] }),
  .ZN({ S9013 })
);
NAND2_X1 #() 
NAND2_X1_2828_ (
  .A1({ S9013 }),
  .A2({ S8991 }),
  .ZN({ S25957[1236] })
);
NOR2_X1 #() 
NOR2_X1_706_ (
  .A1({ S25957[1236] }),
  .A2({ S25956[52] }),
  .ZN({ S9034 })
);
INV_X1 #() 
INV_X1_907_ (
  .A({ S25956[52] }),
  .ZN({ S9042 })
);
AOI21_X1 #() 
AOI21_X1_1555_ (
  .A({ S9042 }),
  .B1({ S9013 }),
  .B2({ S8991 }),
  .ZN({ S9053 })
);
OAI21_X1 #() 
OAI21_X1_1473_ (
  .A({ S8385 }),
  .B1({ S9034 }),
  .B2({ S9053 }),
  .ZN({ S9064 })
);
INV_X1 #() 
INV_X1_908_ (
  .A({ S25957[1236] }),
  .ZN({ S9075 })
);
NAND2_X1 #() 
NAND2_X1_2829_ (
  .A1({ S9075 }),
  .A2({ S9042 }),
  .ZN({ S9086 })
);
INV_X1 #() 
INV_X1_909_ (
  .A({ S9053 }),
  .ZN({ S9097 })
);
NAND3_X1 #() 
NAND3_X1_3054_ (
  .A1({ S9086 }),
  .A2({ S9097 }),
  .A3({ S25956[20] }),
  .ZN({ S9108 })
);
NAND2_X1 #() 
NAND2_X1_2830_ (
  .A1({ S9108 }),
  .A2({ S9064 }),
  .ZN({ S9119 })
);
INV_X1 #() 
INV_X1_910_ (
  .A({ S9119 }),
  .ZN({ S25957[1172] })
);
INV_X1 #() 
INV_X1_911_ (
  .A({ S25956[51] }),
  .ZN({ S9140 })
);
INV_X1 #() 
INV_X1_912_ (
  .A({ S25956[83] }),
  .ZN({ S9151 })
);
OAI221_X1 #() 
OAI221_X1_72_ (
  .A({ S25956[12] }),
  .B1({ S5749 }),
  .B2({ S5719 }),
  .C1({ S7243 }),
  .C2({ S5782 }),
  .ZN({ S9162 })
);
NAND3_X1 #() 
NAND3_X1_3055_ (
  .A1({ S8731 }),
  .A2({ S27 }),
  .A3({ S7210 }),
  .ZN({ S9173 })
);
AND2_X1 #() 
AND2_X1_179_ (
  .A1({ S9162 }),
  .A2({ S9173 }),
  .ZN({ S9183 })
);
NAND3_X1 #() 
NAND3_X1_3056_ (
  .A1({ S7435 }),
  .A2({ S5719 }),
  .A3({ S6303 }),
  .ZN({ S9190 })
);
NOR2_X1 #() 
NOR2_X1_707_ (
  .A1({ S7221 }),
  .A2({ S6194 }),
  .ZN({ S9201 })
);
NAND2_X1 #() 
NAND2_X1_2831_ (
  .A1({ S9201 }),
  .A2({ S25956[11] }),
  .ZN({ S9212 })
);
AOI21_X1 #() 
AOI21_X1_1556_ (
  .A({ S25956[12] }),
  .B1({ S9212 }),
  .B2({ S9190 }),
  .ZN({ S9223 })
);
OAI21_X1 #() 
OAI21_X1_1474_ (
  .A({ S25956[12] }),
  .B1({ S6594 }),
  .B2({ S25956[8] }),
  .ZN({ S9234 })
);
AOI211_X1 #() 
AOI211_X1_36_ (
  .A({ S8865 }),
  .B({ S9234 }),
  .C1({ S29 }),
  .C2({ S5719 }),
  .ZN({ S9245 })
);
OAI21_X1 #() 
OAI21_X1_1475_ (
  .A({ S25956[13] }),
  .B1({ S9223 }),
  .B2({ S9245 }),
  .ZN({ S9256 })
);
OAI211_X1 #() 
OAI211_X1_1002_ (
  .A({ S9256 }),
  .B({ S25956[14] }),
  .C1({ S9183 }),
  .C2({ S25956[13] }),
  .ZN({ S9266 })
);
NAND2_X1 #() 
NAND2_X1_2832_ (
  .A1({ S7254 }),
  .A2({ S6081 }),
  .ZN({ S9276 })
);
NAND2_X1 #() 
NAND2_X1_2833_ (
  .A1({ S8029 }),
  .A2({ S25956[11] }),
  .ZN({ S9287 })
);
NAND3_X1 #() 
NAND3_X1_3057_ (
  .A1({ S9276 }),
  .A2({ S5708 }),
  .A3({ S9287 }),
  .ZN({ S9298 })
);
OAI21_X1 #() 
OAI21_X1_1476_ (
  .A({ S5719 }),
  .B1({ S6194 }),
  .B2({ S6248 }),
  .ZN({ S9309 })
);
OAI211_X1 #() 
OAI211_X1_1003_ (
  .A({ S25956[12] }),
  .B({ S9309 }),
  .C1({ S6709 }),
  .C2({ S6215 }),
  .ZN({ S9320 })
);
NAND3_X1 #() 
NAND3_X1_3058_ (
  .A1({ S9298 }),
  .A2({ S9320 }),
  .A3({ S25956[13] }),
  .ZN({ S9331 })
);
NAND2_X1 #() 
NAND2_X1_2834_ (
  .A1({ S5815 }),
  .A2({ S6533 }),
  .ZN({ S9340 })
);
NOR2_X1 #() 
NOR2_X1_708_ (
  .A1({ S9340 }),
  .A2({ S8521 }),
  .ZN({ S9349 })
);
OAI21_X1 #() 
OAI21_X1_1477_ (
  .A({ S6165 }),
  .B1({ S6270 }),
  .B2({ S6204 }),
  .ZN({ S9360 })
);
OAI21_X1 #() 
OAI21_X1_1478_ (
  .A({ S5708 }),
  .B1({ S9360 }),
  .B2({ S9349 }),
  .ZN({ S9371 })
);
OAI211_X1 #() 
OAI211_X1_1004_ (
  .A({ S8586 }),
  .B({ S25956[12] }),
  .C1({ S6325 }),
  .C2({ S5719 }),
  .ZN({ S9382 })
);
NAND3_X1 #() 
NAND3_X1_3059_ (
  .A1({ S9371 }),
  .A2({ S5697 }),
  .A3({ S9382 }),
  .ZN({ S9393 })
);
AND2_X1 #() 
AND2_X1_180_ (
  .A1({ S9393 }),
  .A2({ S9331 }),
  .ZN({ S9404 })
);
OAI211_X1 #() 
OAI211_X1_1005_ (
  .A({ S9266 }),
  .B({ S25956[15] }),
  .C1({ S9404 }),
  .C2({ S25956[14] }),
  .ZN({ S9414 })
);
NAND2_X1 #() 
NAND2_X1_2835_ (
  .A1({ S8649 }),
  .A2({ S6303 }),
  .ZN({ S9422 })
);
NOR2_X1 #() 
NOR2_X1_709_ (
  .A1({ S5900 }),
  .A2({ S25956[12] }),
  .ZN({ S9433 })
);
AOI22_X1 #() 
AOI22_X1_332_ (
  .A1({ S7113 }),
  .A2({ S6822 }),
  .B1({ S9422 }),
  .B2({ S9433 }),
  .ZN({ S9444 })
);
NOR2_X1 #() 
NOR2_X1_710_ (
  .A1({ S6511 }),
  .A2({ S25956[11] }),
  .ZN({ S9455 })
);
OAI21_X1 #() 
OAI21_X1_1479_ (
  .A({ S5708 }),
  .B1({ S9455 }),
  .B2({ S5837 }),
  .ZN({ S9466 })
);
NAND2_X1 #() 
NAND2_X1_2836_ (
  .A1({ S6081 }),
  .A2({ S25956[8] }),
  .ZN({ S9477 })
);
NAND2_X1 #() 
NAND2_X1_2837_ (
  .A1({ S9477 }),
  .A2({ S5719 }),
  .ZN({ S9488 })
);
OAI211_X1 #() 
OAI211_X1_1006_ (
  .A({ S9466 }),
  .B({ S5697 }),
  .C1({ S5708 }),
  .C2({ S9488 }),
  .ZN({ S9499 })
);
OAI21_X1 #() 
OAI21_X1_1480_ (
  .A({ S9499 }),
  .B1({ S9444 }),
  .B2({ S5697 }),
  .ZN({ S9510 })
);
NAND2_X1 #() 
NAND2_X1_2838_ (
  .A1({ S9510 }),
  .A2({ S25956[14] }),
  .ZN({ S9520 })
);
NOR2_X1 #() 
NOR2_X1_711_ (
  .A1({ S6583 }),
  .A2({ S6605 }),
  .ZN({ S9529 })
);
NAND3_X1 #() 
NAND3_X1_3060_ (
  .A1({ S9529 }),
  .A2({ S5826 }),
  .A3({ S7552 }),
  .ZN({ S9540 })
);
AOI21_X1 #() 
AOI21_X1_1557_ (
  .A({ S6480 }),
  .B1({ S5657 }),
  .B2({ S27 }),
  .ZN({ S9551 })
);
NOR3_X1 #() 
NOR3_X1_96_ (
  .A1({ S7592 }),
  .A2({ S9551 }),
  .A3({ S5708 }),
  .ZN({ S9562 })
);
AOI21_X1 #() 
AOI21_X1_1558_ (
  .A({ S9562 }),
  .B1({ S9540 }),
  .B2({ S5708 }),
  .ZN({ S9573 })
);
NAND3_X1 #() 
NAND3_X1_3061_ (
  .A1({ S7297 }),
  .A2({ S25956[8] }),
  .A3({ S5771 }),
  .ZN({ S9584 })
);
NAND3_X1 #() 
NAND3_X1_3062_ (
  .A1({ S6709 }),
  .A2({ S25956[12] }),
  .A3({ S6838 }),
  .ZN({ S9595 })
);
OAI211_X1 #() 
OAI211_X1_1007_ (
  .A({ S9595 }),
  .B({ S25956[13] }),
  .C1({ S9584 }),
  .C2({ S25956[12] }),
  .ZN({ S9606 })
);
OAI21_X1 #() 
OAI21_X1_1481_ (
  .A({ S9606 }),
  .B1({ S9573 }),
  .B2({ S25956[13] }),
  .ZN({ S9616 })
);
OAI211_X1 #() 
OAI211_X1_1008_ (
  .A({ S9520 }),
  .B({ S5686 }),
  .C1({ S25956[14] }),
  .C2({ S9616 }),
  .ZN({ S9627 })
);
NAND2_X1 #() 
NAND2_X1_2839_ (
  .A1({ S9627 }),
  .A2({ S9414 }),
  .ZN({ S9638 })
);
OR2_X1 #() 
OR2_X1_37_ (
  .A1({ S9638 }),
  .A2({ S25956[115] }),
  .ZN({ S9649 })
);
NAND2_X1 #() 
NAND2_X1_2840_ (
  .A1({ S9638 }),
  .A2({ S25956[115] }),
  .ZN({ S9660 })
);
NAND2_X1 #() 
NAND2_X1_2841_ (
  .A1({ S9649 }),
  .A2({ S9660 }),
  .ZN({ S25957[1267] })
);
NAND2_X1 #() 
NAND2_X1_2842_ (
  .A1({ S25957[1267] }),
  .A2({ S9151 }),
  .ZN({ S9681 })
);
NAND3_X1 #() 
NAND3_X1_3063_ (
  .A1({ S9649 }),
  .A2({ S25956[83] }),
  .A3({ S9660 }),
  .ZN({ S9692 })
);
NAND3_X1 #() 
NAND3_X1_3064_ (
  .A1({ S9681 }),
  .A2({ S9692 }),
  .A3({ S9140 }),
  .ZN({ S9703 })
);
INV_X1 #() 
INV_X1_913_ (
  .A({ S9703 }),
  .ZN({ S9713 })
);
AOI21_X1 #() 
AOI21_X1_1559_ (
  .A({ S9140 }),
  .B1({ S9681 }),
  .B2({ S9692 }),
  .ZN({ S9724 })
);
OAI21_X1 #() 
OAI21_X1_1482_ (
  .A({ S25956[19] }),
  .B1({ S9713 }),
  .B2({ S9724 }),
  .ZN({ S9735 })
);
INV_X1 #() 
INV_X1_914_ (
  .A({ S25956[19] }),
  .ZN({ S9746 })
);
INV_X1 #() 
INV_X1_915_ (
  .A({ S9724 }),
  .ZN({ S9757 })
);
NAND3_X1 #() 
NAND3_X1_3065_ (
  .A1({ S9757 }),
  .A2({ S9746 }),
  .A3({ S9703 }),
  .ZN({ S9768 })
);
NAND2_X1 #() 
NAND2_X1_2843_ (
  .A1({ S9735 }),
  .A2({ S9768 }),
  .ZN({ S25957[1171] })
);
INV_X1 #() 
INV_X1_916_ (
  .A({ S25957[1171] }),
  .ZN({ S50 })
);
INV_X1 #() 
INV_X1_917_ (
  .A({ S25956[48] }),
  .ZN({ S9792 })
);
INV_X1 #() 
INV_X1_918_ (
  .A({ S25956[80] }),
  .ZN({ S9803 })
);
INV_X1 #() 
INV_X1_919_ (
  .A({ S25956[112] }),
  .ZN({ S9814 })
);
NAND3_X1 #() 
NAND3_X1_3066_ (
  .A1({ S7937 }),
  .A2({ S5708 }),
  .A3({ S7030 }),
  .ZN({ S9825 })
);
INV_X1 #() 
INV_X1_920_ (
  .A({ S6081 }),
  .ZN({ S9836 })
);
NOR2_X1 #() 
NOR2_X1_712_ (
  .A1({ S9836 }),
  .A2({ S25956[11] }),
  .ZN({ S9847 })
);
AOI21_X1 #() 
AOI21_X1_1560_ (
  .A({ S5708 }),
  .B1({ S9847 }),
  .B2({ S7339 }),
  .ZN({ S9858 })
);
OAI21_X1 #() 
OAI21_X1_1483_ (
  .A({ S9858 }),
  .B1({ S5719 }),
  .B2({ S6544 }),
  .ZN({ S9869 })
);
INV_X1 #() 
INV_X1_921_ (
  .A({ S8742 }),
  .ZN({ S9880 })
);
OAI22_X1 #() 
OAI22_X1_71_ (
  .A1({ S9880 }),
  .A2({ S5782 }),
  .B1({ S7339 }),
  .B2({ S5719 }),
  .ZN({ S9891 })
);
NAND2_X1 #() 
NAND2_X1_2844_ (
  .A1({ S9891 }),
  .A2({ S5708 }),
  .ZN({ S9901 })
);
AOI21_X1 #() 
AOI21_X1_1561_ (
  .A({ S25956[13] }),
  .B1({ S9901 }),
  .B2({ S9869 }),
  .ZN({ S9911 })
);
NOR2_X1 #() 
NOR2_X1_713_ (
  .A1({ S7782 }),
  .A2({ S5708 }),
  .ZN({ S9917 })
);
AOI21_X1 #() 
AOI21_X1_1562_ (
  .A({ S5697 }),
  .B1({ S9917 }),
  .B2({ S8876 }),
  .ZN({ S9928 })
);
AOI21_X1 #() 
AOI21_X1_1563_ (
  .A({ S9911 }),
  .B1({ S9825 }),
  .B2({ S9928 }),
  .ZN({ S9939 })
);
NAND2_X1 #() 
NAND2_X1_2845_ (
  .A1({ S7625 }),
  .A2({ S25956[11] }),
  .ZN({ S9950 })
);
NAND2_X1 #() 
NAND2_X1_2846_ (
  .A1({ S6811 }),
  .A2({ S25956[11] }),
  .ZN({ S9961 })
);
OAI21_X1 #() 
OAI21_X1_1484_ (
  .A({ S9961 }),
  .B1({ S25956[11] }),
  .B2({ S7435 }),
  .ZN({ S9972 })
);
AOI22_X1 #() 
AOI22_X1_333_ (
  .A1({ S9972 }),
  .A2({ S25956[12] }),
  .B1({ S6365 }),
  .B2({ S9950 }),
  .ZN({ S9983 })
);
NAND2_X1 #() 
NAND2_X1_2847_ (
  .A1({ S9847 }),
  .A2({ S27 }),
  .ZN({ S9993 })
);
NAND3_X1 #() 
NAND3_X1_3067_ (
  .A1({ S7882 }),
  .A2({ S5708 }),
  .A3({ S9993 }),
  .ZN({ S10004 })
);
NAND4_X1 #() 
NAND4_X1_342_ (
  .A1({ S7308 }),
  .A2({ S5889 }),
  .A3({ S5995 }),
  .A4({ S25956[12] }),
  .ZN({ S10012 })
);
NAND3_X1 #() 
NAND3_X1_3068_ (
  .A1({ S10004 }),
  .A2({ S5697 }),
  .A3({ S10012 }),
  .ZN({ S10022 })
);
OAI21_X1 #() 
OAI21_X1_1485_ (
  .A({ S10022 }),
  .B1({ S9983 }),
  .B2({ S5697 }),
  .ZN({ S10033 })
);
NAND2_X1 #() 
NAND2_X1_2848_ (
  .A1({ S10033 }),
  .A2({ S25956[14] }),
  .ZN({ S10044 })
);
OAI21_X1 #() 
OAI21_X1_1486_ (
  .A({ S10044 }),
  .B1({ S25956[14] }),
  .B2({ S9939 }),
  .ZN({ S10055 })
);
NAND2_X1 #() 
NAND2_X1_2849_ (
  .A1({ S10055 }),
  .A2({ S5686 }),
  .ZN({ S10066 })
);
OAI21_X1 #() 
OAI21_X1_1487_ (
  .A({ S7882 }),
  .B1({ S25956[11] }),
  .B2({ S7319 }),
  .ZN({ S10077 })
);
NOR2_X1 #() 
NOR2_X1_714_ (
  .A1({ S9201 }),
  .A2({ S25956[11] }),
  .ZN({ S10087 })
);
OR3_X1 #() 
OR3_X1_16_ (
  .A1({ S10087 }),
  .A2({ S9349 }),
  .A3({ S5708 }),
  .ZN({ S10096 })
);
OAI211_X1 #() 
OAI211_X1_1009_ (
  .A({ S10096 }),
  .B({ S5697 }),
  .C1({ S10077 }),
  .C2({ S25956[12] }),
  .ZN({ S10107 })
);
NAND3_X1 #() 
NAND3_X1_3069_ (
  .A1({ S8854 }),
  .A2({ S25956[12] }),
  .A3({ S9340 }),
  .ZN({ S10118 })
);
NOR2_X1 #() 
NOR2_X1_715_ (
  .A1({ S6215 }),
  .A2({ S6594 }),
  .ZN({ S10129 })
);
OAI21_X1 #() 
OAI21_X1_1488_ (
  .A({ S5708 }),
  .B1({ S5837 }),
  .B2({ S10129 }),
  .ZN({ S10140 })
);
NAND3_X1 #() 
NAND3_X1_3070_ (
  .A1({ S10118 }),
  .A2({ S10140 }),
  .A3({ S25956[13] }),
  .ZN({ S10151 })
);
NAND3_X1 #() 
NAND3_X1_3071_ (
  .A1({ S10107 }),
  .A2({ S25956[14] }),
  .A3({ S10151 }),
  .ZN({ S10160 })
);
NAND2_X1 #() 
NAND2_X1_2850_ (
  .A1({ S8503 }),
  .A2({ S8627 }),
  .ZN({ S10169 })
);
AOI21_X1 #() 
AOI21_X1_1564_ (
  .A({ S9234 }),
  .B1({ S6709 }),
  .B2({ S9488 }),
  .ZN({ S10180 })
);
AOI21_X1 #() 
AOI21_X1_1565_ (
  .A({ S10180 }),
  .B1({ S10169 }),
  .B2({ S5708 }),
  .ZN({ S10191 })
);
AOI21_X1 #() 
AOI21_X1_1566_ (
  .A({ S7157 }),
  .B1({ S5719 }),
  .B2({ S5907 }),
  .ZN({ S10202 })
);
NOR3_X1 #() 
NOR3_X1_97_ (
  .A1({ S10202 }),
  .A2({ S6605 }),
  .A3({ S25956[12] }),
  .ZN({ S10213 })
);
NAND2_X1 #() 
NAND2_X1_2851_ (
  .A1({ S6215 }),
  .A2({ S5719 }),
  .ZN({ S10224 })
);
AND2_X1 #() 
AND2_X1_181_ (
  .A1({ S10224 }),
  .A2({ S7286 }),
  .ZN({ S10235 })
);
OAI21_X1 #() 
OAI21_X1_1489_ (
  .A({ S5697 }),
  .B1({ S10213 }),
  .B2({ S10235 }),
  .ZN({ S10246 })
);
OAI211_X1 #() 
OAI211_X1_1010_ (
  .A({ S10246 }),
  .B({ S6132 }),
  .C1({ S10191 }),
  .C2({ S5697 }),
  .ZN({ S10253 })
);
AND2_X1 #() 
AND2_X1_182_ (
  .A1({ S10160 }),
  .A2({ S10253 }),
  .ZN({ S10262 })
);
NAND2_X1 #() 
NAND2_X1_2852_ (
  .A1({ S10262 }),
  .A2({ S25956[15] }),
  .ZN({ S10273 })
);
NAND3_X1 #() 
NAND3_X1_3072_ (
  .A1({ S10066 }),
  .A2({ S9814 }),
  .A3({ S10273 }),
  .ZN({ S10284 })
);
NAND2_X1 #() 
NAND2_X1_2853_ (
  .A1({ S10066 }),
  .A2({ S10273 }),
  .ZN({ S10295 })
);
NAND2_X1 #() 
NAND2_X1_2854_ (
  .A1({ S10295 }),
  .A2({ S25956[112] }),
  .ZN({ S10306 })
);
NAND2_X1 #() 
NAND2_X1_2855_ (
  .A1({ S10306 }),
  .A2({ S10284 }),
  .ZN({ S25957[1264] })
);
NAND2_X1 #() 
NAND2_X1_2856_ (
  .A1({ S25957[1264] }),
  .A2({ S9803 }),
  .ZN({ S10327 })
);
NAND3_X1 #() 
NAND3_X1_3073_ (
  .A1({ S10306 }),
  .A2({ S25956[80] }),
  .A3({ S10284 }),
  .ZN({ S10338 })
);
NAND3_X1 #() 
NAND3_X1_3074_ (
  .A1({ S10327 }),
  .A2({ S10338 }),
  .A3({ S9792 }),
  .ZN({ S10346 })
);
INV_X1 #() 
INV_X1_922_ (
  .A({ S10346 }),
  .ZN({ S10357 })
);
AOI21_X1 #() 
AOI21_X1_1567_ (
  .A({ S9792 }),
  .B1({ S10327 }),
  .B2({ S10338 }),
  .ZN({ S10368 })
);
OAI21_X1 #() 
OAI21_X1_1490_ (
  .A({ S25956[16] }),
  .B1({ S10357 }),
  .B2({ S10368 }),
  .ZN({ S10379 })
);
INV_X1 #() 
INV_X1_923_ (
  .A({ S25956[16] }),
  .ZN({ S10390 })
);
NAND2_X1 #() 
NAND2_X1_2857_ (
  .A1({ S10327 }),
  .A2({ S10338 }),
  .ZN({ S25957[1232] })
);
NAND2_X1 #() 
NAND2_X1_2858_ (
  .A1({ S25957[1232] }),
  .A2({ S25956[48] }),
  .ZN({ S10407 })
);
NAND3_X1 #() 
NAND3_X1_3075_ (
  .A1({ S10407 }),
  .A2({ S10390 }),
  .A3({ S10346 }),
  .ZN({ S10417 })
);
NAND2_X1 #() 
NAND2_X1_2859_ (
  .A1({ S10379 }),
  .A2({ S10417 }),
  .ZN({ S25957[1168] })
);
INV_X1 #() 
INV_X1_924_ (
  .A({ S25956[49] }),
  .ZN({ S10438 })
);
INV_X1 #() 
INV_X1_925_ (
  .A({ S25956[81] }),
  .ZN({ S10449 })
);
INV_X1 #() 
INV_X1_926_ (
  .A({ S25956[113] }),
  .ZN({ S10460 })
);
AOI21_X1 #() 
AOI21_X1_1568_ (
  .A({ S9349 }),
  .B1({ S7402 }),
  .B2({ S5719 }),
  .ZN({ S10471 })
);
AOI21_X1 #() 
AOI21_X1_1569_ (
  .A({ S6398 }),
  .B1({ S8418 }),
  .B2({ S5741 }),
  .ZN({ S10482 })
);
NAND2_X1 #() 
NAND2_X1_2860_ (
  .A1({ S7855 }),
  .A2({ S25956[12] }),
  .ZN({ S10493 })
);
OAI22_X1 #() 
OAI22_X1_72_ (
  .A1({ S10471 }),
  .A2({ S25956[12] }),
  .B1({ S10482 }),
  .B2({ S10493 }),
  .ZN({ S10504 })
);
AOI21_X1 #() 
AOI21_X1_1570_ (
  .A({ S9551 }),
  .B1({ S8616 }),
  .B2({ S7210 }),
  .ZN({ S10512 })
);
AOI22_X1 #() 
AOI22_X1_334_ (
  .A1({ S6365 }),
  .A2({ S5628 }),
  .B1({ S5708 }),
  .B2({ S6387 }),
  .ZN({ S10522 })
);
OAI211_X1 #() 
OAI211_X1_1011_ (
  .A({ S10522 }),
  .B({ S25956[13] }),
  .C1({ S10512 }),
  .C2({ S5708 }),
  .ZN({ S10533 })
);
OAI21_X1 #() 
OAI21_X1_1491_ (
  .A({ S10533 }),
  .B1({ S10504 }),
  .B2({ S25956[13] }),
  .ZN({ S10544 })
);
NOR3_X1 #() 
NOR3_X1_98_ (
  .A1({ S9455 }),
  .A2({ S6176 }),
  .A3({ S25956[12] }),
  .ZN({ S10555 })
);
AOI21_X1 #() 
AOI21_X1_1571_ (
  .A({ S10555 }),
  .B1({ S8586 }),
  .B2({ S6425 }),
  .ZN({ S10566 })
);
AOI21_X1 #() 
AOI21_X1_1572_ (
  .A({ S5708 }),
  .B1({ S9287 }),
  .B2({ S8660 }),
  .ZN({ S10577 })
);
OR2_X1 #() 
OR2_X1_38_ (
  .A1({ S6522 }),
  .A2({ S5697 }),
  .ZN({ S10588 })
);
OAI221_X1 #() 
OAI221_X1_73_ (
  .A({ S6132 }),
  .B1({ S10588 }),
  .B2({ S10577 }),
  .C1({ S10566 }),
  .C2({ S25956[13] }),
  .ZN({ S10599 })
);
OAI21_X1 #() 
OAI21_X1_1492_ (
  .A({ S10599 }),
  .B1({ S10544 }),
  .B2({ S6132 }),
  .ZN({ S10610 })
);
NAND2_X1 #() 
NAND2_X1_2861_ (
  .A1({ S10610 }),
  .A2({ S5686 }),
  .ZN({ S10621 })
);
NOR2_X1 #() 
NOR2_X1_716_ (
  .A1({ S6709 }),
  .A2({ S8029 }),
  .ZN({ S10632 })
);
OAI211_X1 #() 
OAI211_X1_1012_ (
  .A({ S5708 }),
  .B({ S7552 }),
  .C1({ S9488 }),
  .C2({ S8091 }),
  .ZN({ S10643 })
);
OAI21_X1 #() 
OAI21_X1_1493_ (
  .A({ S10643 }),
  .B1({ S10632 }),
  .B2({ S9234 }),
  .ZN({ S10653 })
);
NOR2_X1 #() 
NOR2_X1_717_ (
  .A1({ S6638 }),
  .A2({ S25956[11] }),
  .ZN({ S10662 })
);
NOR3_X1 #() 
NOR3_X1_99_ (
  .A1({ S8227 }),
  .A2({ S10662 }),
  .A3({ S5708 }),
  .ZN({ S10673 })
);
NOR2_X1 #() 
NOR2_X1_718_ (
  .A1({ S6811 }),
  .A2({ S5719 }),
  .ZN({ S10684 })
);
OAI21_X1 #() 
OAI21_X1_1494_ (
  .A({ S5708 }),
  .B1({ S6742 }),
  .B2({ S25956[11] }),
  .ZN({ S10695 })
);
OAI21_X1 #() 
OAI21_X1_1495_ (
  .A({ S25956[13] }),
  .B1({ S10684 }),
  .B2({ S10695 }),
  .ZN({ S10706 })
);
OAI221_X1 #() 
OAI221_X1_74_ (
  .A({ S25956[14] }),
  .B1({ S10653 }),
  .B2({ S25956[13] }),
  .C1({ S10706 }),
  .C2({ S10673 }),
  .ZN({ S10717 })
);
INV_X1 #() 
INV_X1_927_ (
  .A({ S6763 }),
  .ZN({ S10727 })
);
NAND3_X1 #() 
NAND3_X1_3076_ (
  .A1({ S9422 }),
  .A2({ S7570 }),
  .A3({ S8731 }),
  .ZN({ S10738 })
);
NOR3_X1 #() 
NOR3_X1_100_ (
  .A1({ S6292 }),
  .A2({ S6248 }),
  .A3({ S5719 }),
  .ZN({ S10749 })
);
OAI21_X1 #() 
OAI21_X1_1496_ (
  .A({ S10738 }),
  .B1({ S10727 }),
  .B2({ S10749 }),
  .ZN({ S10760 })
);
NOR2_X1 #() 
NOR2_X1_719_ (
  .A1({ S8448 }),
  .A2({ S6555 }),
  .ZN({ S10771 })
);
AOI21_X1 #() 
AOI21_X1_1573_ (
  .A({ S25956[11] }),
  .B1({ S5749 }),
  .B2({ S6081 }),
  .ZN({ S10782 })
);
OAI21_X1 #() 
OAI21_X1_1497_ (
  .A({ S5697 }),
  .B1({ S10782 }),
  .B2({ S7475 }),
  .ZN({ S10793 })
);
OAI221_X1 #() 
OAI221_X1_75_ (
  .A({ S6132 }),
  .B1({ S10771 }),
  .B2({ S10793 }),
  .C1({ S10760 }),
  .C2({ S5697 }),
  .ZN({ S10803 })
);
NAND3_X1 #() 
NAND3_X1_3077_ (
  .A1({ S10803 }),
  .A2({ S10717 }),
  .A3({ S25956[15] }),
  .ZN({ S10812 })
);
NAND3_X1 #() 
NAND3_X1_3078_ (
  .A1({ S10621 }),
  .A2({ S10460 }),
  .A3({ S10812 }),
  .ZN({ S10819 })
);
NAND2_X1 #() 
NAND2_X1_2862_ (
  .A1({ S10621 }),
  .A2({ S10812 }),
  .ZN({ S10830 })
);
NAND2_X1 #() 
NAND2_X1_2863_ (
  .A1({ S10830 }),
  .A2({ S25956[113] }),
  .ZN({ S10841 })
);
NAND2_X1 #() 
NAND2_X1_2864_ (
  .A1({ S10841 }),
  .A2({ S10819 }),
  .ZN({ S25957[1265] })
);
NAND2_X1 #() 
NAND2_X1_2865_ (
  .A1({ S25957[1265] }),
  .A2({ S10449 }),
  .ZN({ S10862 })
);
NAND3_X1 #() 
NAND3_X1_3079_ (
  .A1({ S10841 }),
  .A2({ S25956[81] }),
  .A3({ S10819 }),
  .ZN({ S10873 })
);
NAND3_X1 #() 
NAND3_X1_3080_ (
  .A1({ S10862 }),
  .A2({ S10873 }),
  .A3({ S10438 }),
  .ZN({ S10884 })
);
INV_X1 #() 
INV_X1_928_ (
  .A({ S10884 }),
  .ZN({ S10895 })
);
AOI21_X1 #() 
AOI21_X1_1574_ (
  .A({ S10438 }),
  .B1({ S10862 }),
  .B2({ S10873 }),
  .ZN({ S10904 })
);
OAI21_X1 #() 
OAI21_X1_1498_ (
  .A({ S25956[17] }),
  .B1({ S10895 }),
  .B2({ S10904 }),
  .ZN({ S10915 })
);
INV_X1 #() 
INV_X1_929_ (
  .A({ S25956[17] }),
  .ZN({ S10926 })
);
INV_X1 #() 
INV_X1_930_ (
  .A({ S10904 }),
  .ZN({ S10937 })
);
NAND3_X1 #() 
NAND3_X1_3081_ (
  .A1({ S10937 }),
  .A2({ S10926 }),
  .A3({ S10884 }),
  .ZN({ S10948 })
);
NAND2_X1 #() 
NAND2_X1_2866_ (
  .A1({ S10915 }),
  .A2({ S10948 }),
  .ZN({ S25957[1169] })
);
INV_X1 #() 
INV_X1_931_ (
  .A({ S25956[50] }),
  .ZN({ S10969 })
);
INV_X1 #() 
INV_X1_932_ (
  .A({ S25956[82] }),
  .ZN({ S10980 })
);
INV_X1 #() 
INV_X1_933_ (
  .A({ S25956[114] }),
  .ZN({ S10990 })
);
NAND3_X1 #() 
NAND3_X1_3082_ (
  .A1({ S8459 }),
  .A2({ S7286 }),
  .A3({ S7570 }),
  .ZN({ S10997 })
);
OAI211_X1 #() 
OAI211_X1_1013_ (
  .A({ S5697 }),
  .B({ S10997 }),
  .C1({ S7647 }),
  .C2({ S10129 }),
  .ZN({ S11006 })
);
NOR3_X1 #() 
NOR3_X1_101_ (
  .A1({ S7074 }),
  .A2({ S7330 }),
  .A3({ S5719 }),
  .ZN({ S11017 })
);
NAND2_X1 #() 
NAND2_X1_2867_ (
  .A1({ S8007 }),
  .A2({ S5708 }),
  .ZN({ S11028 })
);
OAI211_X1 #() 
OAI211_X1_1014_ (
  .A({ S9276 }),
  .B({ S25956[12] }),
  .C1({ S8091 }),
  .C2({ S6480 }),
  .ZN({ S11039 })
);
OAI211_X1 #() 
OAI211_X1_1015_ (
  .A({ S11039 }),
  .B({ S25956[13] }),
  .C1({ S11017 }),
  .C2({ S11028 }),
  .ZN({ S11050 })
);
AOI21_X1 #() 
AOI21_X1_1575_ (
  .A({ S25956[14] }),
  .B1({ S11050 }),
  .B2({ S11006 }),
  .ZN({ S11061 })
);
NAND2_X1 #() 
NAND2_X1_2868_ (
  .A1({ S5867 }),
  .A2({ S5719 }),
  .ZN({ S11072 })
);
NAND3_X1 #() 
NAND3_X1_3083_ (
  .A1({ S9488 }),
  .A2({ S25956[12] }),
  .A3({ S11072 }),
  .ZN({ S11083 })
);
AOI21_X1 #() 
AOI21_X1_1576_ (
  .A({ S11083 }),
  .B1({ S7308 }),
  .B2({ S6491 }),
  .ZN({ S11093 })
);
AOI21_X1 #() 
AOI21_X1_1577_ (
  .A({ S10087 }),
  .B1({ S7508 }),
  .B2({ S25956[11] }),
  .ZN({ S11104 })
);
AOI21_X1 #() 
AOI21_X1_1578_ (
  .A({ S11093 }),
  .B1({ S11104 }),
  .B2({ S5708 }),
  .ZN({ S11115 })
);
NOR2_X1 #() 
NOR2_X1_720_ (
  .A1({ S11115 }),
  .A2({ S25956[13] }),
  .ZN({ S11126 })
);
AOI21_X1 #() 
AOI21_X1_1579_ (
  .A({ S25956[12] }),
  .B1({ S8649 }),
  .B2({ S25956[8] }),
  .ZN({ S11136 })
);
OAI21_X1 #() 
OAI21_X1_1499_ (
  .A({ S7435 }),
  .B1({ S9847 }),
  .B2({ S6154 }),
  .ZN({ S11147 })
);
AOI22_X1 #() 
AOI22_X1_335_ (
  .A1({ S11136 }),
  .A2({ S6334 }),
  .B1({ S11147 }),
  .B2({ S25956[12] }),
  .ZN({ S11158 })
);
AOI211_X1 #() 
AOI211_X1_37_ (
  .A({ S6132 }),
  .B({ S11126 }),
  .C1({ S25956[13] }),
  .C2({ S11158 }),
  .ZN({ S11169 })
);
OAI21_X1 #() 
OAI21_X1_1500_ (
  .A({ S5686 }),
  .B1({ S11169 }),
  .B2({ S11061 }),
  .ZN({ S11180 })
);
NOR4_X1 #() 
NOR4_X1_2_ (
  .A1({ S8649 }),
  .A2({ S7560 }),
  .A3({ S7275 }),
  .A4({ S5708 }),
  .ZN({ S11188 })
);
OAI21_X1 #() 
OAI21_X1_1501_ (
  .A({ S5697 }),
  .B1({ S11028 }),
  .B2({ S7275 }),
  .ZN({ S11198 })
);
INV_X1 #() 
INV_X1_934_ (
  .A({ S9477 }),
  .ZN({ S11209 })
);
AOI211_X1 #() 
AOI211_X1_38_ (
  .A({ S5708 }),
  .B({ S9455 }),
  .C1({ S25956[11] }),
  .C2({ S11209 }),
  .ZN({ S11220 })
);
OAI211_X1 #() 
OAI211_X1_1016_ (
  .A({ S9880 }),
  .B({ S8418 }),
  .C1({ S5657 }),
  .C2({ S5719 }),
  .ZN({ S11231 })
);
OAI21_X1 #() 
OAI21_X1_1502_ (
  .A({ S25956[13] }),
  .B1({ S11231 }),
  .B2({ S25956[12] }),
  .ZN({ S11242 })
);
OAI22_X1 #() 
OAI22_X1_73_ (
  .A1({ S11220 }),
  .A2({ S11242 }),
  .B1({ S11198 }),
  .B2({ S11188 }),
  .ZN({ S11253 })
);
AND3_X1 #() 
AND3_X1_119_ (
  .A1({ S10224 }),
  .A2({ S6502 }),
  .A3({ S11072 }),
  .ZN({ S11264 })
);
AOI211_X1 #() 
AOI211_X1_39_ (
  .A({ S6882 }),
  .B({ S25956[12] }),
  .C1({ S8770 }),
  .C2({ S25956[11] }),
  .ZN({ S11275 })
);
AOI211_X1 #() 
AOI211_X1_40_ (
  .A({ S5697 }),
  .B({ S11275 }),
  .C1({ S11264 }),
  .C2({ S25956[12] }),
  .ZN({ S11285 })
);
AOI21_X1 #() 
AOI21_X1_1580_ (
  .A({ S8124 }),
  .B1({ S6226 }),
  .B2({ S25956[11] }),
  .ZN({ S11294 })
);
AOI211_X1 #() 
AOI211_X1_41_ (
  .A({ S25956[12] }),
  .B({ S6893 }),
  .C1({ S9836 }),
  .C2({ S5719 }),
  .ZN({ S11305 })
);
OR2_X1 #() 
OR2_X1_39_ (
  .A1({ S11305 }),
  .A2({ S25956[13] }),
  .ZN({ S11316 })
);
OAI21_X1 #() 
OAI21_X1_1503_ (
  .A({ S25956[14] }),
  .B1({ S11316 }),
  .B2({ S11294 }),
  .ZN({ S11327 })
);
OAI221_X1 #() 
OAI221_X1_76_ (
  .A({ S25956[15] }),
  .B1({ S11253 }),
  .B2({ S25956[14] }),
  .C1({ S11285 }),
  .C2({ S11327 }),
  .ZN({ S11338 })
);
AND2_X1 #() 
AND2_X1_183_ (
  .A1({ S11180 }),
  .A2({ S11338 }),
  .ZN({ S11349 })
);
NAND2_X1 #() 
NAND2_X1_2869_ (
  .A1({ S11349 }),
  .A2({ S10990 }),
  .ZN({ S11360 })
);
NAND2_X1 #() 
NAND2_X1_2870_ (
  .A1({ S11180 }),
  .A2({ S11338 }),
  .ZN({ S11371 })
);
NAND2_X1 #() 
NAND2_X1_2871_ (
  .A1({ S11371 }),
  .A2({ S25956[114] }),
  .ZN({ S11382 })
);
NAND3_X1 #() 
NAND3_X1_3084_ (
  .A1({ S11360 }),
  .A2({ S10980 }),
  .A3({ S11382 }),
  .ZN({ S11393 })
);
NAND2_X1 #() 
NAND2_X1_2872_ (
  .A1({ S11371 }),
  .A2({ S10990 }),
  .ZN({ S11404 })
);
NAND2_X1 #() 
NAND2_X1_2873_ (
  .A1({ S11349 }),
  .A2({ S25956[114] }),
  .ZN({ S11414 })
);
NAND3_X1 #() 
NAND3_X1_3085_ (
  .A1({ S11414 }),
  .A2({ S25956[82] }),
  .A3({ S11404 }),
  .ZN({ S11421 })
);
NAND3_X1 #() 
NAND3_X1_3086_ (
  .A1({ S11393 }),
  .A2({ S11421 }),
  .A3({ S10969 }),
  .ZN({ S11432 })
);
NAND3_X1 #() 
NAND3_X1_3087_ (
  .A1({ S11414 }),
  .A2({ S10980 }),
  .A3({ S11404 }),
  .ZN({ S11443 })
);
NAND3_X1 #() 
NAND3_X1_3088_ (
  .A1({ S11360 }),
  .A2({ S25956[82] }),
  .A3({ S11382 }),
  .ZN({ S11454 })
);
NAND3_X1 #() 
NAND3_X1_3089_ (
  .A1({ S11443 }),
  .A2({ S11454 }),
  .A3({ S25956[50] }),
  .ZN({ S11465 })
);
NAND3_X1 #() 
NAND3_X1_3090_ (
  .A1({ S11432 }),
  .A2({ S11465 }),
  .A3({ S25956[18] }),
  .ZN({ S11476 })
);
INV_X1 #() 
INV_X1_935_ (
  .A({ S25956[18] }),
  .ZN({ S11487 })
);
NAND3_X1 #() 
NAND3_X1_3091_ (
  .A1({ S11443 }),
  .A2({ S11454 }),
  .A3({ S10969 }),
  .ZN({ S11498 })
);
NAND3_X1 #() 
NAND3_X1_3092_ (
  .A1({ S11393 }),
  .A2({ S11421 }),
  .A3({ S25956[50] }),
  .ZN({ S11507 })
);
NAND3_X1 #() 
NAND3_X1_3093_ (
  .A1({ S11498 }),
  .A2({ S11507 }),
  .A3({ S11487 }),
  .ZN({ S11518 })
);
NAND2_X1 #() 
NAND2_X1_2874_ (
  .A1({ S11476 }),
  .A2({ S11518 }),
  .ZN({ S25957[1170] })
);
INV_X1 #() 
INV_X1_936_ (
  .A({ S25956[1] }),
  .ZN({ S11539 })
);
INV_X1 #() 
INV_X1_937_ (
  .A({ S25956[0] }),
  .ZN({ S11550 })
);
NAND2_X1 #() 
NAND2_X1_2875_ (
  .A1({ S11539 }),
  .A2({ S11550 }),
  .ZN({ S56 })
);
AND2_X1 #() 
AND2_X1_184_ (
  .A1({ S25956[0] }),
  .A2({ S25956[1] }),
  .ZN({ S58 })
);
INV_X1 #() 
INV_X1_938_ (
  .A({ S25956[47] }),
  .ZN({ S11581 })
);
INV_X1 #() 
INV_X1_939_ (
  .A({ S25956[79] }),
  .ZN({ S11590 })
);
INV_X1 #() 
INV_X1_940_ (
  .A({ S25956[111] }),
  .ZN({ S11598 })
);
INV_X1 #() 
INV_X1_941_ (
  .A({ S25956[7] }),
  .ZN({ S11609 })
);
INV_X1 #() 
INV_X1_942_ (
  .A({ S25956[6] }),
  .ZN({ S11620 })
);
INV_X1 #() 
INV_X1_943_ (
  .A({ S25956[5] }),
  .ZN({ S11631 })
);
INV_X1 #() 
INV_X1_944_ (
  .A({ S25956[2] }),
  .ZN({ S11642 })
);
NAND2_X1 #() 
NAND2_X1_2876_ (
  .A1({ S11642 }),
  .A2({ S25956[1] }),
  .ZN({ S11653 })
);
INV_X1 #() 
INV_X1_945_ (
  .A({ S25956[3] }),
  .ZN({ S11664 })
);
AOI21_X1 #() 
AOI21_X1_1581_ (
  .A({ S11664 }),
  .B1({ S25956[2] }),
  .B2({ S25956[0] }),
  .ZN({ S11672 })
);
NAND2_X1 #() 
NAND2_X1_2877_ (
  .A1({ S11672 }),
  .A2({ S11653 }),
  .ZN({ S11683 })
);
INV_X1 #() 
INV_X1_946_ (
  .A({ S11683 }),
  .ZN({ S11694 })
);
AOI21_X1 #() 
AOI21_X1_1582_ (
  .A({ S11642 }),
  .B1({ S25956[1] }),
  .B2({ S25956[0] }),
  .ZN({ S11705 })
);
NAND2_X1 #() 
NAND2_X1_2878_ (
  .A1({ S11705 }),
  .A2({ S11664 }),
  .ZN({ S11716 })
);
NAND2_X1 #() 
NAND2_X1_2879_ (
  .A1({ S11539 }),
  .A2({ S25956[0] }),
  .ZN({ S11727 })
);
NOR2_X1 #() 
NOR2_X1_721_ (
  .A1({ S25956[3] }),
  .A2({ S25956[2] }),
  .ZN({ S11736 })
);
AOI21_X1 #() 
AOI21_X1_1583_ (
  .A({ S25956[4] }),
  .B1({ S11727 }),
  .B2({ S11736 }),
  .ZN({ S11744 })
);
NAND2_X1 #() 
NAND2_X1_2880_ (
  .A1({ S11716 }),
  .A2({ S11744 }),
  .ZN({ S11755 })
);
NAND2_X1 #() 
NAND2_X1_2881_ (
  .A1({ S25956[1] }),
  .A2({ S25956[0] }),
  .ZN({ S11766 })
);
NAND2_X1 #() 
NAND2_X1_2882_ (
  .A1({ S11766 }),
  .A2({ S25956[2] }),
  .ZN({ S11777 })
);
NAND2_X1 #() 
NAND2_X1_2883_ (
  .A1({ S11550 }),
  .A2({ S25956[1] }),
  .ZN({ S11788 })
);
NAND3_X1 #() 
NAND3_X1_3094_ (
  .A1({ S11727 }),
  .A2({ S11788 }),
  .A3({ S11642 }),
  .ZN({ S11799 })
);
AOI21_X1 #() 
AOI21_X1_1584_ (
  .A({ S11664 }),
  .B1({ S11799 }),
  .B2({ S11777 }),
  .ZN({ S11810 })
);
AND2_X1 #() 
AND2_X1_185_ (
  .A1({ S25956[0] }),
  .A2({ S25956[2] }),
  .ZN({ S11821 })
);
NOR2_X1 #() 
NOR2_X1_722_ (
  .A1({ S11539 }),
  .A2({ S25956[3] }),
  .ZN({ S11832 })
);
NAND2_X1 #() 
NAND2_X1_2884_ (
  .A1({ S11832 }),
  .A2({ S11821 }),
  .ZN({ S11842 })
);
NAND2_X1 #() 
NAND2_X1_2885_ (
  .A1({ S25956[2] }),
  .A2({ S25956[1] }),
  .ZN({ S11853 })
);
NAND3_X1 #() 
NAND3_X1_3095_ (
  .A1({ S11853 }),
  .A2({ S11664 }),
  .A3({ S11550 }),
  .ZN({ S11864 })
);
NAND3_X1 #() 
NAND3_X1_3096_ (
  .A1({ S11842 }),
  .A2({ S25956[4] }),
  .A3({ S11864 }),
  .ZN({ S11875 })
);
OAI22_X1 #() 
OAI22_X1_74_ (
  .A1({ S11810 }),
  .A2({ S11875 }),
  .B1({ S11755 }),
  .B2({ S11694 }),
  .ZN({ S11886 })
);
NAND2_X1 #() 
NAND2_X1_2886_ (
  .A1({ S11886 }),
  .A2({ S11631 }),
  .ZN({ S11895 })
);
NAND3_X1 #() 
NAND3_X1_3097_ (
  .A1({ S11539 }),
  .A2({ S11550 }),
  .A3({ S25956[2] }),
  .ZN({ S11906 })
);
NAND2_X1 #() 
NAND2_X1_2887_ (
  .A1({ S11906 }),
  .A2({ S25956[3] }),
  .ZN({ S11917 })
);
AOI21_X1 #() 
AOI21_X1_1585_ (
  .A({ S11917 }),
  .B1({ S58 }),
  .B2({ S11642 }),
  .ZN({ S11928 })
);
NAND2_X1 #() 
NAND2_X1_2888_ (
  .A1({ S11642 }),
  .A2({ S11550 }),
  .ZN({ S11939 })
);
NAND3_X1 #() 
NAND3_X1_3098_ (
  .A1({ S11550 }),
  .A2({ S25956[2] }),
  .A3({ S25956[1] }),
  .ZN({ S11950 })
);
NAND3_X1 #() 
NAND3_X1_3099_ (
  .A1({ S11950 }),
  .A2({ S11939 }),
  .A3({ S11664 }),
  .ZN({ S11961 })
);
NAND2_X1 #() 
NAND2_X1_2889_ (
  .A1({ S11961 }),
  .A2({ S25956[4] }),
  .ZN({ S11971 })
);
NOR2_X1 #() 
NOR2_X1_723_ (
  .A1({ S11642 }),
  .A2({ S25956[1] }),
  .ZN({ S11978 })
);
AOI21_X1 #() 
AOI21_X1_1586_ (
  .A({ S25956[2] }),
  .B1({ S11539 }),
  .B2({ S25956[0] }),
  .ZN({ S11987 })
);
OAI21_X1 #() 
OAI21_X1_1504_ (
  .A({ S25956[3] }),
  .B1({ S11987 }),
  .B2({ S11978 }),
  .ZN({ S11998 })
);
AND2_X1 #() 
AND2_X1_186_ (
  .A1({ S11998 }),
  .A2({ S11716 }),
  .ZN({ S12009 })
);
OAI221_X1 #() 
OAI221_X1_77_ (
  .A({ S25956[5] }),
  .B1({ S11928 }),
  .B2({ S11971 }),
  .C1({ S12009 }),
  .C2({ S25956[4] }),
  .ZN({ S12020 })
);
AOI21_X1 #() 
AOI21_X1_1587_ (
  .A({ S11620 }),
  .B1({ S12020 }),
  .B2({ S11895 }),
  .ZN({ S12031 })
);
NAND2_X1 #() 
NAND2_X1_2890_ (
  .A1({ S11766 }),
  .A2({ S11642 }),
  .ZN({ S12042 })
);
AOI21_X1 #() 
AOI21_X1_1588_ (
  .A({ S25956[3] }),
  .B1({ S25956[2] }),
  .B2({ S25956[1] }),
  .ZN({ S12053 })
);
NAND2_X1 #() 
NAND2_X1_2891_ (
  .A1({ S12042 }),
  .A2({ S12053 }),
  .ZN({ S12064 })
);
NAND3_X1 #() 
NAND3_X1_3100_ (
  .A1({ S11727 }),
  .A2({ S11653 }),
  .A3({ S25956[3] }),
  .ZN({ S12075 })
);
AOI21_X1 #() 
AOI21_X1_1589_ (
  .A({ S25956[4] }),
  .B1({ S12075 }),
  .B2({ S12064 }),
  .ZN({ S12086 })
);
NAND2_X1 #() 
NAND2_X1_2892_ (
  .A1({ S11642 }),
  .A2({ S11539 }),
  .ZN({ S12097 })
);
NAND2_X1 #() 
NAND2_X1_2893_ (
  .A1({ S11672 }),
  .A2({ S12097 }),
  .ZN({ S12108 })
);
INV_X1 #() 
INV_X1_947_ (
  .A({ S25956[4] }),
  .ZN({ S12118 })
);
NOR2_X1 #() 
NOR2_X1_724_ (
  .A1({ S11550 }),
  .A2({ S25956[3] }),
  .ZN({ S12127 })
);
NOR2_X1 #() 
NOR2_X1_725_ (
  .A1({ S12127 }),
  .A2({ S12118 }),
  .ZN({ S12138 })
);
AOI21_X1 #() 
AOI21_X1_1590_ (
  .A({ S12086 }),
  .B1({ S12108 }),
  .B2({ S12138 }),
  .ZN({ S12149 })
);
OAI21_X1 #() 
OAI21_X1_1505_ (
  .A({ S25956[2] }),
  .B1({ S25956[1] }),
  .B2({ S25956[0] }),
  .ZN({ S12160 })
);
NAND3_X1 #() 
NAND3_X1_3101_ (
  .A1({ S11642 }),
  .A2({ S25956[1] }),
  .A3({ S25956[0] }),
  .ZN({ S12171 })
);
OAI211_X1 #() 
OAI211_X1_1017_ (
  .A({ S12171 }),
  .B({ S11664 }),
  .C1({ S12160 }),
  .C2({ S58 }),
  .ZN({ S12182 })
);
AOI21_X1 #() 
AOI21_X1_1591_ (
  .A({ S12118 }),
  .B1({ S11950 }),
  .B2({ S25956[3] }),
  .ZN({ S12193 })
);
NOR3_X1 #() 
NOR3_X1_102_ (
  .A1({ S11642 }),
  .A2({ S25956[1] }),
  .A3({ S25956[0] }),
  .ZN({ S12201 })
);
AND3_X1 #() 
AND3_X1_120_ (
  .A1({ S25956[0] }),
  .A2({ S25956[1] }),
  .A3({ S25956[2] }),
  .ZN({ S12210 })
);
NOR2_X1 #() 
NOR2_X1_726_ (
  .A1({ S12201 }),
  .A2({ S12210 }),
  .ZN({ S12221 })
);
NOR2_X1 #() 
NOR2_X1_727_ (
  .A1({ S12221 }),
  .A2({ S25956[3] }),
  .ZN({ S12232 })
);
NOR2_X1 #() 
NOR2_X1_728_ (
  .A1({ S11777 }),
  .A2({ S11664 }),
  .ZN({ S12243 })
);
NOR3_X1 #() 
NOR3_X1_103_ (
  .A1({ S12232 }),
  .A2({ S12243 }),
  .A3({ S25956[4] }),
  .ZN({ S12254 })
);
AOI21_X1 #() 
AOI21_X1_1592_ (
  .A({ S12254 }),
  .B1({ S12193 }),
  .B2({ S12182 }),
  .ZN({ S12265 })
);
MUX2_X1 #() 
MUX2_X1_10_ (
  .A({ S12149 }),
  .B({ S12265 }),
  .S({ S11631 }),
  .Z({ S12276 })
);
AOI21_X1 #() 
AOI21_X1_1593_ (
  .A({ S12031 }),
  .B1({ S12276 }),
  .B2({ S11620 }),
  .ZN({ S12283 })
);
NAND2_X1 #() 
NAND2_X1_2894_ (
  .A1({ S12283 }),
  .A2({ S11609 }),
  .ZN({ S12292 })
);
AOI21_X1 #() 
AOI21_X1_1594_ (
  .A({ S25956[0] }),
  .B1({ S25956[1] }),
  .B2({ S25956[2] }),
  .ZN({ S12303 })
);
OAI21_X1 #() 
OAI21_X1_1506_ (
  .A({ S25956[3] }),
  .B1({ S12303 }),
  .B2({ S58 }),
  .ZN({ S12314 })
);
NAND3_X1 #() 
NAND3_X1_3102_ (
  .A1({ S11906 }),
  .A2({ S12171 }),
  .A3({ S11664 }),
  .ZN({ S12325 })
);
AOI21_X1 #() 
AOI21_X1_1595_ (
  .A({ S25956[4] }),
  .B1({ S12325 }),
  .B2({ S12314 }),
  .ZN({ S12336 })
);
OAI21_X1 #() 
OAI21_X1_1507_ (
  .A({ S25956[1] }),
  .B1({ S25956[2] }),
  .B2({ S25956[0] }),
  .ZN({ S12347 })
);
OAI21_X1 #() 
OAI21_X1_1508_ (
  .A({ S25956[3] }),
  .B1({ S11987 }),
  .B2({ S11821 }),
  .ZN({ S12357 })
);
OAI21_X1 #() 
OAI21_X1_1509_ (
  .A({ S12357 }),
  .B1({ S25956[3] }),
  .B2({ S12347 }),
  .ZN({ S12366 })
);
OAI21_X1 #() 
OAI21_X1_1510_ (
  .A({ S25956[5] }),
  .B1({ S12366 }),
  .B2({ S12118 }),
  .ZN({ S12377 })
);
NAND2_X1 #() 
NAND2_X1_2895_ (
  .A1({ S11539 }),
  .A2({ S25956[2] }),
  .ZN({ S12388 })
);
NAND3_X1 #() 
NAND3_X1_3103_ (
  .A1({ S12388 }),
  .A2({ S25956[3] }),
  .A3({ S11766 }),
  .ZN({ S12399 })
);
NAND2_X1 #() 
NAND2_X1_2896_ (
  .A1({ S11788 }),
  .A2({ S11664 }),
  .ZN({ S12410 })
);
AOI21_X1 #() 
AOI21_X1_1596_ (
  .A({ S12118 }),
  .B1({ S12399 }),
  .B2({ S12410 }),
  .ZN({ S12421 })
);
INV_X1 #() 
INV_X1_948_ (
  .A({ S12160 }),
  .ZN({ S12432 })
);
NOR2_X1 #() 
NOR2_X1_729_ (
  .A1({ S25956[2] }),
  .A2({ S25956[1] }),
  .ZN({ S12442 })
);
INV_X1 #() 
INV_X1_949_ (
  .A({ S12127 }),
  .ZN({ S12449 })
);
AOI211_X1 #() 
AOI211_X1_42_ (
  .A({ S25956[4] }),
  .B({ S12432 }),
  .C1({ S12442 }),
  .C2({ S12449 }),
  .ZN({ S12457 })
);
OAI21_X1 #() 
OAI21_X1_1511_ (
  .A({ S11631 }),
  .B1({ S12457 }),
  .B2({ S12421 }),
  .ZN({ S12468 })
);
OAI21_X1 #() 
OAI21_X1_1512_ (
  .A({ S12468 }),
  .B1({ S12336 }),
  .B2({ S12377 }),
  .ZN({ S12479 })
);
NOR3_X1 #() 
NOR3_X1_104_ (
  .A1({ S11664 }),
  .A2({ S25956[2] }),
  .A3({ S25956[1] }),
  .ZN({ S12490 })
);
OAI21_X1 #() 
OAI21_X1_1513_ (
  .A({ S25956[2] }),
  .B1({ S11550 }),
  .B2({ S25956[1] }),
  .ZN({ S12501 })
);
AOI21_X1 #() 
AOI21_X1_1597_ (
  .A({ S25956[2] }),
  .B1({ S25956[1] }),
  .B2({ S25956[0] }),
  .ZN({ S12512 })
);
NAND2_X1 #() 
NAND2_X1_2897_ (
  .A1({ S56 }),
  .A2({ S12512 }),
  .ZN({ S12520 })
);
AND2_X1 #() 
AND2_X1_187_ (
  .A1({ S12520 }),
  .A2({ S12501 }),
  .ZN({ S12530 })
);
AOI21_X1 #() 
AOI21_X1_1598_ (
  .A({ S12490 }),
  .B1({ S12530 }),
  .B2({ S11664 }),
  .ZN({ S12541 })
);
NAND3_X1 #() 
NAND3_X1_3104_ (
  .A1({ S11987 }),
  .A2({ S25956[3] }),
  .A3({ S11788 }),
  .ZN({ S12552 })
);
AOI21_X1 #() 
AOI21_X1_1599_ (
  .A({ S25956[3] }),
  .B1({ S11642 }),
  .B2({ S25956[0] }),
  .ZN({ S12563 })
);
NAND2_X1 #() 
NAND2_X1_2898_ (
  .A1({ S12563 }),
  .A2({ S11853 }),
  .ZN({ S12574 })
);
NAND3_X1 #() 
NAND3_X1_3105_ (
  .A1({ S12432 }),
  .A2({ S25956[3] }),
  .A3({ S11766 }),
  .ZN({ S12581 })
);
NAND4_X1 #() 
NAND4_X1_343_ (
  .A1({ S12581 }),
  .A2({ S12552 }),
  .A3({ S12574 }),
  .A4({ S25956[4] }),
  .ZN({ S12589 })
);
OAI211_X1 #() 
OAI211_X1_1018_ (
  .A({ S12589 }),
  .B({ S11631 }),
  .C1({ S12541 }),
  .C2({ S25956[4] }),
  .ZN({ S12600 })
);
NOR2_X1 #() 
NOR2_X1_730_ (
  .A1({ S11664 }),
  .A2({ S25956[0] }),
  .ZN({ S12611 })
);
AOI21_X1 #() 
AOI21_X1_1600_ (
  .A({ S25956[4] }),
  .B1({ S11939 }),
  .B2({ S11664 }),
  .ZN({ S12622 })
);
OAI21_X1 #() 
OAI21_X1_1514_ (
  .A({ S12622 }),
  .B1({ S11539 }),
  .B2({ S12611 }),
  .ZN({ S12633 })
);
NAND2_X1 #() 
NAND2_X1_2899_ (
  .A1({ S11664 }),
  .A2({ S25956[1] }),
  .ZN({ S12644 })
);
NAND2_X1 #() 
NAND2_X1_2900_ (
  .A1({ S25956[2] }),
  .A2({ S25956[0] }),
  .ZN({ S12655 })
);
AOI21_X1 #() 
AOI21_X1_1601_ (
  .A({ S11664 }),
  .B1({ S12655 }),
  .B2({ S25956[1] }),
  .ZN({ S12666 })
);
NOR2_X1 #() 
NOR2_X1_731_ (
  .A1({ S12666 }),
  .A2({ S12118 }),
  .ZN({ S12676 })
);
OAI21_X1 #() 
OAI21_X1_1515_ (
  .A({ S12676 }),
  .B1({ S11821 }),
  .B2({ S12644 }),
  .ZN({ S12684 })
);
NAND3_X1 #() 
NAND3_X1_3106_ (
  .A1({ S12684 }),
  .A2({ S25956[5] }),
  .A3({ S12633 }),
  .ZN({ S12695 })
);
NAND3_X1 #() 
NAND3_X1_3107_ (
  .A1({ S12600 }),
  .A2({ S11620 }),
  .A3({ S12695 }),
  .ZN({ S12706 })
);
OAI211_X1 #() 
OAI211_X1_1019_ (
  .A({ S12706 }),
  .B({ S25956[7] }),
  .C1({ S12479 }),
  .C2({ S11620 }),
  .ZN({ S12717 })
);
NAND2_X1 #() 
NAND2_X1_2901_ (
  .A1({ S12292 }),
  .A2({ S12717 }),
  .ZN({ S12728 })
);
NAND2_X1 #() 
NAND2_X1_2902_ (
  .A1({ S12728 }),
  .A2({ S11598 }),
  .ZN({ S12739 })
);
NAND3_X1 #() 
NAND3_X1_3108_ (
  .A1({ S12292 }),
  .A2({ S25956[111] }),
  .A3({ S12717 }),
  .ZN({ S12750 })
);
NAND2_X1 #() 
NAND2_X1_2903_ (
  .A1({ S12739 }),
  .A2({ S12750 }),
  .ZN({ S12761 })
);
NAND2_X1 #() 
NAND2_X1_2904_ (
  .A1({ S12761 }),
  .A2({ S11590 }),
  .ZN({ S12772 })
);
INV_X1 #() 
INV_X1_950_ (
  .A({ S12761 }),
  .ZN({ S25957[1263] })
);
NAND2_X1 #() 
NAND2_X1_2905_ (
  .A1({ S25957[1263] }),
  .A2({ S25956[79] }),
  .ZN({ S12793 })
);
NAND2_X1 #() 
NAND2_X1_2906_ (
  .A1({ S12793 }),
  .A2({ S12772 }),
  .ZN({ S12802 })
);
NAND2_X1 #() 
NAND2_X1_2907_ (
  .A1({ S12802 }),
  .A2({ S11581 }),
  .ZN({ S12811 })
);
NAND3_X1 #() 
NAND3_X1_3109_ (
  .A1({ S12793 }),
  .A2({ S25956[47] }),
  .A3({ S12772 }),
  .ZN({ S12822 })
);
NAND3_X1 #() 
NAND3_X1_3110_ (
  .A1({ S12811 }),
  .A2({ S12822 }),
  .A3({ S5686 }),
  .ZN({ S12833 })
);
NAND3_X1 #() 
NAND3_X1_3111_ (
  .A1({ S12793 }),
  .A2({ S11581 }),
  .A3({ S12772 }),
  .ZN({ S12844 })
);
NAND2_X1 #() 
NAND2_X1_2908_ (
  .A1({ S12802 }),
  .A2({ S25956[47] }),
  .ZN({ S12855 })
);
NAND3_X1 #() 
NAND3_X1_3112_ (
  .A1({ S12855 }),
  .A2({ S25956[15] }),
  .A3({ S12844 }),
  .ZN({ S12866 })
);
NAND2_X1 #() 
NAND2_X1_2909_ (
  .A1({ S12833 }),
  .A2({ S12866 }),
  .ZN({ S25957[1167] })
);
INV_X1 #() 
INV_X1_951_ (
  .A({ S25956[46] }),
  .ZN({ S12886 })
);
INV_X1 #() 
INV_X1_952_ (
  .A({ S25956[78] }),
  .ZN({ S12895 })
);
INV_X1 #() 
INV_X1_953_ (
  .A({ S25956[110] }),
  .ZN({ S12906 })
);
NOR2_X1 #() 
NOR2_X1_732_ (
  .A1({ S11550 }),
  .A2({ S25956[2] }),
  .ZN({ S12917 })
);
OAI21_X1 #() 
OAI21_X1_1516_ (
  .A({ S11664 }),
  .B1({ S11705 }),
  .B2({ S12917 }),
  .ZN({ S12928 })
);
NAND2_X1 #() 
NAND2_X1_2910_ (
  .A1({ S11672 }),
  .A2({ S11788 }),
  .ZN({ S12939 })
);
NAND3_X1 #() 
NAND3_X1_3113_ (
  .A1({ S12928 }),
  .A2({ S25956[4] }),
  .A3({ S12939 }),
  .ZN({ S12950 })
);
NAND2_X1 #() 
NAND2_X1_2911_ (
  .A1({ S11642 }),
  .A2({ S25956[0] }),
  .ZN({ S12961 })
);
AOI21_X1 #() 
AOI21_X1_1602_ (
  .A({ S25956[3] }),
  .B1({ S12961 }),
  .B2({ S25956[1] }),
  .ZN({ S12970 })
);
AOI21_X1 #() 
AOI21_X1_1603_ (
  .A({ S12970 }),
  .B1({ S11672 }),
  .B2({ S11788 }),
  .ZN({ S12978 })
);
OAI21_X1 #() 
OAI21_X1_1517_ (
  .A({ S12950 }),
  .B1({ S12978 }),
  .B2({ S25956[4] }),
  .ZN({ S12989 })
);
NAND3_X1 #() 
NAND3_X1_3114_ (
  .A1({ S11853 }),
  .A2({ S12655 }),
  .A3({ S11664 }),
  .ZN({ S13000 })
);
NAND2_X1 #() 
NAND2_X1_2912_ (
  .A1({ S12501 }),
  .A2({ S12961 }),
  .ZN({ S13011 })
);
NAND2_X1 #() 
NAND2_X1_2913_ (
  .A1({ S13011 }),
  .A2({ S25956[3] }),
  .ZN({ S13022 })
);
NAND3_X1 #() 
NAND3_X1_3115_ (
  .A1({ S11664 }),
  .A2({ S25956[1] }),
  .A3({ S25956[0] }),
  .ZN({ S13033 })
);
AND4_X1 #() 
AND4_X1_8_ (
  .A1({ S12118 }),
  .A2({ S13022 }),
  .A3({ S13033 }),
  .A4({ S13000 }),
  .ZN({ S13044 })
);
OAI21_X1 #() 
OAI21_X1_1518_ (
  .A({ S11550 }),
  .B1({ S25956[2] }),
  .B2({ S25956[1] }),
  .ZN({ S13055 })
);
NOR2_X1 #() 
NOR2_X1_733_ (
  .A1({ S13055 }),
  .A2({ S25956[3] }),
  .ZN({ S13066 })
);
OAI21_X1 #() 
OAI21_X1_1519_ (
  .A({ S25956[4] }),
  .B1({ S11653 }),
  .B2({ S11664 }),
  .ZN({ S13077 })
);
OAI21_X1 #() 
OAI21_X1_1520_ (
  .A({ S11631 }),
  .B1({ S13066 }),
  .B2({ S13077 }),
  .ZN({ S13087 })
);
OAI22_X1 #() 
OAI22_X1_75_ (
  .A1({ S12989 }),
  .A2({ S11631 }),
  .B1({ S13044 }),
  .B2({ S13087 }),
  .ZN({ S13098 })
);
NAND2_X1 #() 
NAND2_X1_2914_ (
  .A1({ S11550 }),
  .A2({ S25956[2] }),
  .ZN({ S13109 })
);
NAND3_X1 #() 
NAND3_X1_3116_ (
  .A1({ S13109 }),
  .A2({ S25956[3] }),
  .A3({ S11766 }),
  .ZN({ S13120 })
);
NOR2_X1 #() 
NOR2_X1_734_ (
  .A1({ S12563 }),
  .A2({ S12118 }),
  .ZN({ S13131 })
);
NAND3_X1 #() 
NAND3_X1_3117_ (
  .A1({ S11550 }),
  .A2({ S25956[3] }),
  .A3({ S25956[1] }),
  .ZN({ S13142 })
);
AND3_X1 #() 
AND3_X1_121_ (
  .A1({ S13131 }),
  .A2({ S13120 }),
  .A3({ S13142 }),
  .ZN({ S13153 })
);
OAI21_X1 #() 
OAI21_X1_1521_ (
  .A({ S11642 }),
  .B1({ S11539 }),
  .B2({ S25956[0] }),
  .ZN({ S13161 })
);
AOI21_X1 #() 
AOI21_X1_1604_ (
  .A({ S11664 }),
  .B1({ S13161 }),
  .B2({ S11950 }),
  .ZN({ S13172 })
);
OAI211_X1 #() 
OAI211_X1_1020_ (
  .A({ S11998 }),
  .B({ S25956[4] }),
  .C1({ S12097 }),
  .C2({ S12449 }),
  .ZN({ S13183 })
);
OAI21_X1 #() 
OAI21_X1_1522_ (
  .A({ S13183 }),
  .B1({ S25956[4] }),
  .B2({ S13172 }),
  .ZN({ S13194 })
);
OAI21_X1 #() 
OAI21_X1_1523_ (
  .A({ S11642 }),
  .B1({ S11550 }),
  .B2({ S25956[1] }),
  .ZN({ S13205 })
);
AOI21_X1 #() 
AOI21_X1_1605_ (
  .A({ S25956[3] }),
  .B1({ S13205 }),
  .B2({ S12388 }),
  .ZN({ S13216 })
);
INV_X1 #() 
INV_X1_954_ (
  .A({ S11653 }),
  .ZN({ S13227 })
);
NAND2_X1 #() 
NAND2_X1_2915_ (
  .A1({ S12388 }),
  .A2({ S25956[3] }),
  .ZN({ S13238 })
);
OAI21_X1 #() 
OAI21_X1_1524_ (
  .A({ S12118 }),
  .B1({ S13238 }),
  .B2({ S13227 }),
  .ZN({ S13248 })
);
OAI21_X1 #() 
OAI21_X1_1525_ (
  .A({ S25956[5] }),
  .B1({ S13248 }),
  .B2({ S13216 }),
  .ZN({ S13259 })
);
OAI221_X1 #() 
OAI221_X1_78_ (
  .A({ S11620 }),
  .B1({ S13153 }),
  .B2({ S13259 }),
  .C1({ S13194 }),
  .C2({ S25956[5] }),
  .ZN({ S13270 })
);
OAI21_X1 #() 
OAI21_X1_1526_ (
  .A({ S13270 }),
  .B1({ S11620 }),
  .B2({ S13098 }),
  .ZN({ S13281 })
);
NOR2_X1 #() 
NOR2_X1_735_ (
  .A1({ S11664 }),
  .A2({ S25956[1] }),
  .ZN({ S13292 })
);
NAND3_X1 #() 
NAND3_X1_3118_ (
  .A1({ S13292 }),
  .A2({ S13109 }),
  .A3({ S12961 }),
  .ZN({ S13302 })
);
OAI211_X1 #() 
OAI211_X1_1021_ (
  .A({ S13302 }),
  .B({ S25956[4] }),
  .C1({ S12160 }),
  .C2({ S25956[3] }),
  .ZN({ S13313 })
);
NAND2_X1 #() 
NAND2_X1_2916_ (
  .A1({ S12399 }),
  .A2({ S12644 }),
  .ZN({ S13323 })
);
AOI21_X1 #() 
AOI21_X1_1606_ (
  .A({ S11631 }),
  .B1({ S13323 }),
  .B2({ S12118 }),
  .ZN({ S13334 })
);
NOR2_X1 #() 
NOR2_X1_736_ (
  .A1({ S11917 }),
  .A2({ S12512 }),
  .ZN({ S13345 })
);
NAND4_X1 #() 
NAND4_X1_344_ (
  .A1({ S12171 }),
  .A2({ S56 }),
  .A3({ S13109 }),
  .A4({ S11664 }),
  .ZN({ S13356 })
);
NAND3_X1 #() 
NAND3_X1_3119_ (
  .A1({ S13022 }),
  .A2({ S25956[4] }),
  .A3({ S13356 }),
  .ZN({ S13367 })
);
OAI21_X1 #() 
OAI21_X1_1527_ (
  .A({ S13367 }),
  .B1({ S11755 }),
  .B2({ S13345 }),
  .ZN({ S13378 })
);
AOI22_X1 #() 
AOI22_X1_336_ (
  .A1({ S13378 }),
  .A2({ S11631 }),
  .B1({ S13334 }),
  .B2({ S13313 }),
  .ZN({ S13387 })
);
NOR2_X1 #() 
NOR2_X1_737_ (
  .A1({ S25956[1] }),
  .A2({ S25956[0] }),
  .ZN({ S13395 })
);
OAI21_X1 #() 
OAI21_X1_1528_ (
  .A({ S11664 }),
  .B1({ S12210 }),
  .B2({ S13395 }),
  .ZN({ S13406 })
);
NAND3_X1 #() 
NAND3_X1_3120_ (
  .A1({ S11550 }),
  .A2({ S11642 }),
  .A3({ S25956[1] }),
  .ZN({ S13417 })
);
NAND3_X1 #() 
NAND3_X1_3121_ (
  .A1({ S13417 }),
  .A2({ S25956[3] }),
  .A3({ S12388 }),
  .ZN({ S13428 })
);
AOI21_X1 #() 
AOI21_X1_1607_ (
  .A({ S25956[4] }),
  .B1({ S13406 }),
  .B2({ S13428 }),
  .ZN({ S13439 })
);
NAND2_X1 #() 
NAND2_X1_2917_ (
  .A1({ S12655 }),
  .A2({ S25956[3] }),
  .ZN({ S13450 })
);
OAI21_X1 #() 
OAI21_X1_1529_ (
  .A({ S13356 }),
  .B1({ S12303 }),
  .B2({ S13450 }),
  .ZN({ S13461 })
);
NOR2_X1 #() 
NOR2_X1_738_ (
  .A1({ S13461 }),
  .A2({ S25956[4] }),
  .ZN({ S13472 })
);
AOI21_X1 #() 
AOI21_X1_1608_ (
  .A({ S12666 }),
  .B1({ S11987 }),
  .B2({ S11664 }),
  .ZN({ S13483 })
);
OAI21_X1 #() 
OAI21_X1_1530_ (
  .A({ S11631 }),
  .B1({ S13483 }),
  .B2({ S12118 }),
  .ZN({ S13494 })
);
AOI21_X1 #() 
AOI21_X1_1609_ (
  .A({ S25956[3] }),
  .B1({ S12221 }),
  .B2({ S13417 }),
  .ZN({ S13505 })
);
NAND3_X1 #() 
NAND3_X1_3122_ (
  .A1({ S25956[3] }),
  .A2({ S25956[2] }),
  .A3({ S25956[1] }),
  .ZN({ S13516 })
);
NAND2_X1 #() 
NAND2_X1_2918_ (
  .A1({ S13516 }),
  .A2({ S25956[4] }),
  .ZN({ S13525 })
);
OAI21_X1 #() 
OAI21_X1_1531_ (
  .A({ S25956[5] }),
  .B1({ S13505 }),
  .B2({ S13525 }),
  .ZN({ S13533 })
);
OAI22_X1 #() 
OAI22_X1_76_ (
  .A1({ S13533 }),
  .A2({ S13439 }),
  .B1({ S13472 }),
  .B2({ S13494 }),
  .ZN({ S13544 })
);
MUX2_X1 #() 
MUX2_X1_11_ (
  .A({ S13387 }),
  .B({ S13544 }),
  .S({ S11620 }),
  .Z({ S13555 })
);
NAND2_X1 #() 
NAND2_X1_2919_ (
  .A1({ S13555 }),
  .A2({ S25956[7] }),
  .ZN({ S13566 })
);
OAI211_X1 #() 
OAI211_X1_1022_ (
  .A({ S13566 }),
  .B({ S12906 }),
  .C1({ S13281 }),
  .C2({ S25956[7] }),
  .ZN({ S13577 })
);
OR2_X1 #() 
OR2_X1_40_ (
  .A1({ S13555 }),
  .A2({ S11609 }),
  .ZN({ S13588 })
);
NAND2_X1 #() 
NAND2_X1_2920_ (
  .A1({ S13281 }),
  .A2({ S11609 }),
  .ZN({ S13599 })
);
NAND3_X1 #() 
NAND3_X1_3123_ (
  .A1({ S13588 }),
  .A2({ S25956[110] }),
  .A3({ S13599 }),
  .ZN({ S13610 })
);
NAND2_X1 #() 
NAND2_X1_2921_ (
  .A1({ S13610 }),
  .A2({ S13577 }),
  .ZN({ S25957[1262] })
);
NAND2_X1 #() 
NAND2_X1_2922_ (
  .A1({ S25957[1262] }),
  .A2({ S12895 }),
  .ZN({ S13629 })
);
INV_X1 #() 
INV_X1_955_ (
  .A({ S25957[1262] }),
  .ZN({ S13640 })
);
NAND2_X1 #() 
NAND2_X1_2923_ (
  .A1({ S13640 }),
  .A2({ S25956[78] }),
  .ZN({ S13651 })
);
NAND3_X1 #() 
NAND3_X1_3124_ (
  .A1({ S13651 }),
  .A2({ S12886 }),
  .A3({ S13629 }),
  .ZN({ S13662 })
);
INV_X1 #() 
INV_X1_956_ (
  .A({ S13662 }),
  .ZN({ S13673 })
);
AOI21_X1 #() 
AOI21_X1_1610_ (
  .A({ S12886 }),
  .B1({ S13651 }),
  .B2({ S13629 }),
  .ZN({ S13684 })
);
OAI21_X1 #() 
OAI21_X1_1532_ (
  .A({ S25956[14] }),
  .B1({ S13673 }),
  .B2({ S13684 }),
  .ZN({ S13691 })
);
NAND2_X1 #() 
NAND2_X1_2924_ (
  .A1({ S13651 }),
  .A2({ S13629 }),
  .ZN({ S25957[1230] })
);
NAND2_X1 #() 
NAND2_X1_2925_ (
  .A1({ S25957[1230] }),
  .A2({ S25956[46] }),
  .ZN({ S13712 })
);
NAND3_X1 #() 
NAND3_X1_3125_ (
  .A1({ S13712 }),
  .A2({ S6132 }),
  .A3({ S13662 }),
  .ZN({ S13723 })
);
NAND2_X1 #() 
NAND2_X1_2926_ (
  .A1({ S13691 }),
  .A2({ S13723 }),
  .ZN({ S25957[1166] })
);
INV_X1 #() 
INV_X1_957_ (
  .A({ S25956[45] }),
  .ZN({ S13744 })
);
INV_X1 #() 
INV_X1_958_ (
  .A({ S25956[109] }),
  .ZN({ S13755 })
);
NAND2_X1 #() 
NAND2_X1_2927_ (
  .A1({ S12171 }),
  .A2({ S11664 }),
  .ZN({ S13766 })
);
OAI21_X1 #() 
OAI21_X1_1533_ (
  .A({ S11642 }),
  .B1({ S25956[1] }),
  .B2({ S25956[0] }),
  .ZN({ S13776 })
);
NAND3_X1 #() 
NAND3_X1_3126_ (
  .A1({ S12221 }),
  .A2({ S25956[3] }),
  .A3({ S13776 }),
  .ZN({ S13784 })
);
AOI21_X1 #() 
AOI21_X1_1611_ (
  .A({ S25956[4] }),
  .B1({ S13784 }),
  .B2({ S13766 }),
  .ZN({ S13795 })
);
NAND3_X1 #() 
NAND3_X1_3127_ (
  .A1({ S56 }),
  .A2({ S12512 }),
  .A3({ S25956[3] }),
  .ZN({ S13806 })
);
AOI21_X1 #() 
AOI21_X1_1612_ (
  .A({ S12118 }),
  .B1({ S12563 }),
  .B2({ S11539 }),
  .ZN({ S13817 })
);
AOI211_X1 #() 
AOI211_X1_43_ (
  .A({ S25956[5] }),
  .B({ S13795 }),
  .C1({ S13806 }),
  .C2({ S13817 }),
  .ZN({ S13828 })
);
AND2_X1 #() 
AND2_X1_188_ (
  .A1({ S25956[2] }),
  .A2({ S25956[3] }),
  .ZN({ S13839 })
);
AOI21_X1 #() 
AOI21_X1_1613_ (
  .A({ S13839 }),
  .B1({ S11939 }),
  .B2({ S11766 }),
  .ZN({ S13850 })
);
OAI21_X1 #() 
OAI21_X1_1534_ (
  .A({ S25956[4] }),
  .B1({ S13850 }),
  .B2({ S12243 }),
  .ZN({ S13861 })
);
NAND2_X1 #() 
NAND2_X1_2928_ (
  .A1({ S11539 }),
  .A2({ S25956[3] }),
  .ZN({ S13872 })
);
AOI21_X1 #() 
AOI21_X1_1614_ (
  .A({ S25956[3] }),
  .B1({ S11550 }),
  .B2({ S25956[1] }),
  .ZN({ S13883 })
);
NAND2_X1 #() 
NAND2_X1_2929_ (
  .A1({ S13883 }),
  .A2({ S12097 }),
  .ZN({ S13893 })
);
NAND3_X1 #() 
NAND3_X1_3128_ (
  .A1({ S13893 }),
  .A2({ S12118 }),
  .A3({ S13872 }),
  .ZN({ S13902 })
);
AOI21_X1 #() 
AOI21_X1_1615_ (
  .A({ S11631 }),
  .B1({ S13861 }),
  .B2({ S13902 }),
  .ZN({ S13913 })
);
OR2_X1 #() 
OR2_X1_41_ (
  .A1({ S13913 }),
  .A2({ S25956[6] }),
  .ZN({ S13924 })
);
NAND2_X1 #() 
NAND2_X1_2930_ (
  .A1({ S12347 }),
  .A2({ S25956[3] }),
  .ZN({ S13935 })
);
AND3_X1 #() 
AND3_X1_122_ (
  .A1({ S13935 }),
  .A2({ S12644 }),
  .A3({ S12655 }),
  .ZN({ S13946 })
);
OAI221_X1 #() 
OAI221_X1_79_ (
  .A({ S25956[4] }),
  .B1({ S13055 }),
  .B2({ S11664 }),
  .C1({ S12410 }),
  .C2({ S11987 }),
  .ZN({ S13957 })
);
OAI211_X1 #() 
OAI211_X1_1023_ (
  .A({ S13957 }),
  .B({ S25956[5] }),
  .C1({ S13946 }),
  .C2({ S25956[4] }),
  .ZN({ S13968 })
);
NAND2_X1 #() 
NAND2_X1_2931_ (
  .A1({ S13022 }),
  .A2({ S12118 }),
  .ZN({ S13979 })
);
NAND2_X1 #() 
NAND2_X1_2932_ (
  .A1({ S11788 }),
  .A2({ S25956[2] }),
  .ZN({ S13987 })
);
NAND3_X1 #() 
NAND3_X1_3129_ (
  .A1({ S13987 }),
  .A2({ S25956[4] }),
  .A3({ S13142 }),
  .ZN({ S13998 })
);
OAI21_X1 #() 
OAI21_X1_1535_ (
  .A({ S13998 }),
  .B1({ S13979 }),
  .B2({ S12232 }),
  .ZN({ S14009 })
);
NAND2_X1 #() 
NAND2_X1_2933_ (
  .A1({ S14009 }),
  .A2({ S11631 }),
  .ZN({ S14020 })
);
NAND3_X1 #() 
NAND3_X1_3130_ (
  .A1({ S14020 }),
  .A2({ S25956[6] }),
  .A3({ S13968 }),
  .ZN({ S14031 })
);
OAI211_X1 #() 
OAI211_X1_1024_ (
  .A({ S14031 }),
  .B({ S25956[7] }),
  .C1({ S13828 }),
  .C2({ S13924 }),
  .ZN({ S14042 })
);
NAND3_X1 #() 
NAND3_X1_3131_ (
  .A1({ S25956[2] }),
  .A2({ S25956[1] }),
  .A3({ S25956[0] }),
  .ZN({ S14053 })
);
NAND4_X1 #() 
NAND4_X1_345_ (
  .A1({ S13417 }),
  .A2({ S11906 }),
  .A3({ S14053 }),
  .A4({ S25956[3] }),
  .ZN({ S14064 })
);
NAND3_X1 #() 
NAND3_X1_3132_ (
  .A1({ S13205 }),
  .A2({ S11664 }),
  .A3({ S12388 }),
  .ZN({ S14073 })
);
AND2_X1 #() 
AND2_X1_189_ (
  .A1({ S14073 }),
  .A2({ S25956[4] }),
  .ZN({ S14084 })
);
INV_X1 #() 
INV_X1_959_ (
  .A({ S12611 }),
  .ZN({ S14095 })
);
NAND2_X1 #() 
NAND2_X1_2934_ (
  .A1({ S13883 }),
  .A2({ S12961 }),
  .ZN({ S14106 })
);
AOI21_X1 #() 
AOI21_X1_1616_ (
  .A({ S25956[4] }),
  .B1({ S14106 }),
  .B2({ S14095 }),
  .ZN({ S14117 })
);
AOI211_X1 #() 
AOI211_X1_44_ (
  .A({ S11631 }),
  .B({ S14117 }),
  .C1({ S14064 }),
  .C2({ S14084 }),
  .ZN({ S14128 })
);
AOI21_X1 #() 
AOI21_X1_1617_ (
  .A({ S12118 }),
  .B1({ S11987 }),
  .B2({ S25956[3] }),
  .ZN({ S14138 })
);
NAND3_X1 #() 
NAND3_X1_3133_ (
  .A1({ S13883 }),
  .A2({ S11939 }),
  .A3({ S11727 }),
  .ZN({ S14146 })
);
NAND3_X1 #() 
NAND3_X1_3134_ (
  .A1({ S12581 }),
  .A2({ S14138 }),
  .A3({ S14146 }),
  .ZN({ S14157 })
);
AOI22_X1 #() 
AOI22_X1_337_ (
  .A1({ S11832 }),
  .A2({ S11821 }),
  .B1({ S13292 }),
  .B2({ S25956[0] }),
  .ZN({ S14168 })
);
OAI211_X1 #() 
OAI211_X1_1025_ (
  .A({ S14157 }),
  .B({ S11631 }),
  .C1({ S25956[4] }),
  .C2({ S14168 }),
  .ZN({ S14179 })
);
NAND3_X1 #() 
NAND3_X1_3135_ (
  .A1({ S13417 }),
  .A2({ S11664 }),
  .A3({ S14053 }),
  .ZN({ S14190 })
);
NAND3_X1 #() 
NAND3_X1_3136_ (
  .A1({ S14190 }),
  .A2({ S12118 }),
  .A3({ S13450 }),
  .ZN({ S14201 })
);
OAI221_X1 #() 
OAI221_X1_80_ (
  .A({ S25956[4] }),
  .B1({ S12512 }),
  .B2({ S11664 }),
  .C1({ S11939 }),
  .C2({ S12644 }),
  .ZN({ S14212 })
);
NAND3_X1 #() 
NAND3_X1_3137_ (
  .A1({ S14201 }),
  .A2({ S14212 }),
  .A3({ S25956[5] }),
  .ZN({ S14223 })
);
NAND3_X1 #() 
NAND3_X1_3138_ (
  .A1({ S14179 }),
  .A2({ S11620 }),
  .A3({ S14223 }),
  .ZN({ S14234 })
);
NAND3_X1 #() 
NAND3_X1_3139_ (
  .A1({ S13417 }),
  .A2({ S11664 }),
  .A3({ S12655 }),
  .ZN({ S14245 })
);
NAND3_X1 #() 
NAND3_X1_3140_ (
  .A1({ S11777 }),
  .A2({ S25956[3] }),
  .A3({ S12961 }),
  .ZN({ S14256 })
);
AND2_X1 #() 
AND2_X1_190_ (
  .A1({ S14245 }),
  .A2({ S14256 }),
  .ZN({ S14267 })
);
NAND3_X1 #() 
NAND3_X1_3141_ (
  .A1({ S12042 }),
  .A2({ S11664 }),
  .A3({ S14053 }),
  .ZN({ S14275 })
);
NAND2_X1 #() 
NAND2_X1_2935_ (
  .A1({ S14138 }),
  .A2({ S14275 }),
  .ZN({ S14286 })
);
OAI21_X1 #() 
OAI21_X1_1536_ (
  .A({ S14286 }),
  .B1({ S14267 }),
  .B2({ S25956[4] }),
  .ZN({ S14297 })
);
OAI21_X1 #() 
OAI21_X1_1537_ (
  .A({ S25956[6] }),
  .B1({ S14297 }),
  .B2({ S25956[5] }),
  .ZN({ S14308 })
);
OAI211_X1 #() 
OAI211_X1_1026_ (
  .A({ S14234 }),
  .B({ S11609 }),
  .C1({ S14308 }),
  .C2({ S14128 }),
  .ZN({ S14319 })
);
AOI21_X1 #() 
AOI21_X1_1618_ (
  .A({ S13755 }),
  .B1({ S14042 }),
  .B2({ S14319 }),
  .ZN({ S14330 })
);
NAND3_X1 #() 
NAND3_X1_3142_ (
  .A1({ S14042 }),
  .A2({ S14319 }),
  .A3({ S13755 }),
  .ZN({ S14341 })
);
INV_X1 #() 
INV_X1_960_ (
  .A({ S14341 }),
  .ZN({ S14352 })
);
OAI21_X1 #() 
OAI21_X1_1538_ (
  .A({ S25956[77] }),
  .B1({ S14352 }),
  .B2({ S14330 }),
  .ZN({ S14362 })
);
INV_X1 #() 
INV_X1_961_ (
  .A({ S25956[77] }),
  .ZN({ S14369 })
);
INV_X1 #() 
INV_X1_962_ (
  .A({ S14330 }),
  .ZN({ S14380 })
);
NAND3_X1 #() 
NAND3_X1_3143_ (
  .A1({ S14380 }),
  .A2({ S14369 }),
  .A3({ S14341 }),
  .ZN({ S14391 })
);
NAND3_X1 #() 
NAND3_X1_3144_ (
  .A1({ S14362 }),
  .A2({ S14391 }),
  .A3({ S13744 }),
  .ZN({ S14402 })
);
OAI21_X1 #() 
OAI21_X1_1539_ (
  .A({ S14369 }),
  .B1({ S14352 }),
  .B2({ S14330 }),
  .ZN({ S14413 })
);
NAND3_X1 #() 
NAND3_X1_3145_ (
  .A1({ S14380 }),
  .A2({ S25956[77] }),
  .A3({ S14341 }),
  .ZN({ S14424 })
);
NAND3_X1 #() 
NAND3_X1_3146_ (
  .A1({ S14413 }),
  .A2({ S14424 }),
  .A3({ S25956[45] }),
  .ZN({ S14435 })
);
NAND3_X1 #() 
NAND3_X1_3147_ (
  .A1({ S14402 }),
  .A2({ S14435 }),
  .A3({ S25956[13] }),
  .ZN({ S14446 })
);
NAND3_X1 #() 
NAND3_X1_3148_ (
  .A1({ S14362 }),
  .A2({ S14391 }),
  .A3({ S25956[45] }),
  .ZN({ S14453 })
);
NAND3_X1 #() 
NAND3_X1_3149_ (
  .A1({ S14413 }),
  .A2({ S14424 }),
  .A3({ S13744 }),
  .ZN({ S14461 })
);
NAND3_X1 #() 
NAND3_X1_3150_ (
  .A1({ S14453 }),
  .A2({ S14461 }),
  .A3({ S5697 }),
  .ZN({ S14472 })
);
NAND2_X1 #() 
NAND2_X1_2936_ (
  .A1({ S14446 }),
  .A2({ S14472 }),
  .ZN({ S14483 })
);
INV_X1 #() 
INV_X1_963_ (
  .A({ S14483 }),
  .ZN({ S25957[1165] })
);
INV_X1 #() 
INV_X1_964_ (
  .A({ S25956[76] }),
  .ZN({ S14504 })
);
INV_X1 #() 
INV_X1_965_ (
  .A({ S25956[108] }),
  .ZN({ S14515 })
);
NAND3_X1 #() 
NAND3_X1_3151_ (
  .A1({ S12171 }),
  .A2({ S11664 }),
  .A3({ S13109 }),
  .ZN({ S14526 })
);
AOI21_X1 #() 
AOI21_X1_1619_ (
  .A({ S25956[4] }),
  .B1({ S25956[2] }),
  .B2({ S25956[3] }),
  .ZN({ S14534 })
);
NAND2_X1 #() 
NAND2_X1_2937_ (
  .A1({ S14526 }),
  .A2({ S14534 }),
  .ZN({ S14545 })
);
OAI21_X1 #() 
OAI21_X1_1540_ (
  .A({ S12676 }),
  .B1({ S12442 }),
  .B2({ S13000 }),
  .ZN({ S14556 })
);
NAND2_X1 #() 
NAND2_X1_2938_ (
  .A1({ S14556 }),
  .A2({ S14545 }),
  .ZN({ S14567 })
);
INV_X1 #() 
INV_X1_966_ (
  .A({ S117 }),
  .ZN({ S14578 })
);
OAI21_X1 #() 
OAI21_X1_1541_ (
  .A({ S25956[4] }),
  .B1({ S14578 }),
  .B2({ S25956[2] }),
  .ZN({ S14589 })
);
AOI21_X1 #() 
AOI21_X1_1620_ (
  .A({ S25956[3] }),
  .B1({ S12520 }),
  .B2({ S13987 }),
  .ZN({ S14595 })
);
NAND2_X1 #() 
NAND2_X1_2939_ (
  .A1({ S14256 }),
  .A2({ S12118 }),
  .ZN({ S14606 })
);
OAI211_X1 #() 
OAI211_X1_1027_ (
  .A({ S14589 }),
  .B({ S25956[5] }),
  .C1({ S14595 }),
  .C2({ S14606 }),
  .ZN({ S14617 })
);
OAI211_X1 #() 
OAI211_X1_1028_ (
  .A({ S14617 }),
  .B({ S25956[6] }),
  .C1({ S14567 }),
  .C2({ S25956[5] }),
  .ZN({ S14628 })
);
NAND3_X1 #() 
NAND3_X1_3152_ (
  .A1({ S11906 }),
  .A2({ S13776 }),
  .A3({ S11664 }),
  .ZN({ S14639 })
);
NAND3_X1 #() 
NAND3_X1_3153_ (
  .A1({ S56 }),
  .A2({ S25956[3] }),
  .A3({ S12655 }),
  .ZN({ S14650 })
);
AOI21_X1 #() 
AOI21_X1_1621_ (
  .A({ S25956[4] }),
  .B1({ S14639 }),
  .B2({ S14650 }),
  .ZN({ S14661 })
);
NAND4_X1 #() 
NAND4_X1_346_ (
  .A1({ S11939 }),
  .A2({ S11653 }),
  .A3({ S25956[3] }),
  .A4({ S12655 }),
  .ZN({ S14671 })
);
NAND3_X1 #() 
NAND3_X1_3154_ (
  .A1({ S14671 }),
  .A2({ S13893 }),
  .A3({ S25956[4] }),
  .ZN({ S14678 })
);
INV_X1 #() 
INV_X1_967_ (
  .A({ S14678 }),
  .ZN({ S14689 })
);
OAI21_X1 #() 
OAI21_X1_1542_ (
  .A({ S11631 }),
  .B1({ S14689 }),
  .B2({ S14661 }),
  .ZN({ S14700 })
);
NAND3_X1 #() 
NAND3_X1_3155_ (
  .A1({ S12388 }),
  .A2({ S11664 }),
  .A3({ S12655 }),
  .ZN({ S14711 })
);
NAND3_X1 #() 
NAND3_X1_3156_ (
  .A1({ S11998 }),
  .A2({ S25956[4] }),
  .A3({ S14711 }),
  .ZN({ S14722 })
);
NAND3_X1 #() 
NAND3_X1_3157_ (
  .A1({ S13806 }),
  .A2({ S12118 }),
  .A3({ S13033 }),
  .ZN({ S14733 })
);
NAND3_X1 #() 
NAND3_X1_3158_ (
  .A1({ S14722 }),
  .A2({ S25956[5] }),
  .A3({ S14733 }),
  .ZN({ S14742 })
);
NAND3_X1 #() 
NAND3_X1_3159_ (
  .A1({ S14700 }),
  .A2({ S11620 }),
  .A3({ S14742 }),
  .ZN({ S14752 })
);
NAND3_X1 #() 
NAND3_X1_3160_ (
  .A1({ S14752 }),
  .A2({ S14628 }),
  .A3({ S11609 }),
  .ZN({ S14763 })
);
NOR2_X1 #() 
NOR2_X1_739_ (
  .A1({ S13872 }),
  .A2({ S11821 }),
  .ZN({ S14774 })
);
NOR3_X1 #() 
NOR3_X1_105_ (
  .A1({ S11539 }),
  .A2({ S25956[0] }),
  .A3({ S25956[2] }),
  .ZN({ S14785 })
);
OAI21_X1 #() 
OAI21_X1_1543_ (
  .A({ S12118 }),
  .B1({ S14711 }),
  .B2({ S14785 }),
  .ZN({ S14796 })
);
NAND2_X1 #() 
NAND2_X1_2940_ (
  .A1({ S11653 }),
  .A2({ S12655 }),
  .ZN({ S14807 })
);
OAI21_X1 #() 
OAI21_X1_1544_ (
  .A({ S11664 }),
  .B1({ S12347 }),
  .B2({ S11821 }),
  .ZN({ S14817 })
);
OAI21_X1 #() 
OAI21_X1_1545_ (
  .A({ S14817 }),
  .B1({ S14807 }),
  .B2({ S13238 }),
  .ZN({ S14824 })
);
OAI22_X1 #() 
OAI22_X1_77_ (
  .A1({ S14824 }),
  .A2({ S12118 }),
  .B1({ S14796 }),
  .B2({ S14774 }),
  .ZN({ S14835 })
);
AOI21_X1 #() 
AOI21_X1_1622_ (
  .A({ S25956[3] }),
  .B1({ S11799 }),
  .B2({ S11777 }),
  .ZN({ S14846 })
);
NAND3_X1 #() 
NAND3_X1_3161_ (
  .A1({ S11727 }),
  .A2({ S25956[3] }),
  .A3({ S11642 }),
  .ZN({ S14857 })
);
NAND2_X1 #() 
NAND2_X1_2941_ (
  .A1({ S14857 }),
  .A2({ S13142 }),
  .ZN({ S14868 })
);
OAI21_X1 #() 
OAI21_X1_1546_ (
  .A({ S12118 }),
  .B1({ S14846 }),
  .B2({ S14868 }),
  .ZN({ S14879 })
);
OAI211_X1 #() 
OAI211_X1_1029_ (
  .A({ S13417 }),
  .B({ S25956[4] }),
  .C1({ S11727 }),
  .C2({ S11736 }),
  .ZN({ S14890 })
);
AND2_X1 #() 
AND2_X1_191_ (
  .A1({ S14890 }),
  .A2({ S25956[5] }),
  .ZN({ S14901 })
);
AOI22_X1 #() 
AOI22_X1_338_ (
  .A1({ S14835 }),
  .A2({ S11631 }),
  .B1({ S14879 }),
  .B2({ S14901 }),
  .ZN({ S14912 })
);
NOR2_X1 #() 
NOR2_X1_740_ (
  .A1({ S12917 }),
  .A2({ S13872 }),
  .ZN({ S14923 })
);
NAND2_X1 #() 
NAND2_X1_2942_ (
  .A1({ S13893 }),
  .A2({ S25956[4] }),
  .ZN({ S14934 })
);
NAND2_X1 #() 
NAND2_X1_2943_ (
  .A1({ S14807 }),
  .A2({ S11664 }),
  .ZN({ S14945 })
);
NAND3_X1 #() 
NAND3_X1_3162_ (
  .A1({ S14945 }),
  .A2({ S12118 }),
  .A3({ S12075 }),
  .ZN({ S14956 })
);
OAI21_X1 #() 
OAI21_X1_1547_ (
  .A({ S14956 }),
  .B1({ S14923 }),
  .B2({ S14934 }),
  .ZN({ S14964 })
);
NAND2_X1 #() 
NAND2_X1_2944_ (
  .A1({ S11906 }),
  .A2({ S11664 }),
  .ZN({ S14975 })
);
NAND2_X1 #() 
NAND2_X1_2945_ (
  .A1({ S14138 }),
  .A2({ S14975 }),
  .ZN({ S14986 })
);
OAI21_X1 #() 
OAI21_X1_1548_ (
  .A({ S11664 }),
  .B1({ S11539 }),
  .B2({ S25956[2] }),
  .ZN({ S14997 })
);
OAI211_X1 #() 
OAI211_X1_1030_ (
  .A({ S12108 }),
  .B({ S12118 }),
  .C1({ S25956[0] }),
  .C2({ S14997 }),
  .ZN({ S15008 })
);
NAND3_X1 #() 
NAND3_X1_3163_ (
  .A1({ S15008 }),
  .A2({ S25956[5] }),
  .A3({ S14986 }),
  .ZN({ S15019 })
);
OAI211_X1 #() 
OAI211_X1_1031_ (
  .A({ S15019 }),
  .B({ S25956[6] }),
  .C1({ S14964 }),
  .C2({ S25956[5] }),
  .ZN({ S15030 })
);
OAI211_X1 #() 
OAI211_X1_1032_ (
  .A({ S15030 }),
  .B({ S25956[7] }),
  .C1({ S14912 }),
  .C2({ S25956[6] }),
  .ZN({ S15040 })
);
NAND3_X1 #() 
NAND3_X1_3164_ (
  .A1({ S15040 }),
  .A2({ S14763 }),
  .A3({ S14515 }),
  .ZN({ S15049 })
);
NAND2_X1 #() 
NAND2_X1_2946_ (
  .A1({ S14835 }),
  .A2({ S11631 }),
  .ZN({ S15060 })
);
NAND2_X1 #() 
NAND2_X1_2947_ (
  .A1({ S14879 }),
  .A2({ S14901 }),
  .ZN({ S15071 })
);
NAND3_X1 #() 
NAND3_X1_3165_ (
  .A1({ S15060 }),
  .A2({ S15071 }),
  .A3({ S11620 }),
  .ZN({ S15082 })
);
OAI21_X1 #() 
OAI21_X1_1549_ (
  .A({ S15019 }),
  .B1({ S14964 }),
  .B2({ S25956[5] }),
  .ZN({ S15093 })
);
NAND2_X1 #() 
NAND2_X1_2948_ (
  .A1({ S15093 }),
  .A2({ S25956[6] }),
  .ZN({ S15104 })
);
NAND3_X1 #() 
NAND3_X1_3166_ (
  .A1({ S15104 }),
  .A2({ S15082 }),
  .A3({ S25956[7] }),
  .ZN({ S15115 })
);
NAND2_X1 #() 
NAND2_X1_2949_ (
  .A1({ S14752 }),
  .A2({ S14628 }),
  .ZN({ S15126 })
);
NAND2_X1 #() 
NAND2_X1_2950_ (
  .A1({ S15126 }),
  .A2({ S11609 }),
  .ZN({ S15135 })
);
NAND3_X1 #() 
NAND3_X1_3167_ (
  .A1({ S15135 }),
  .A2({ S15115 }),
  .A3({ S25956[108] }),
  .ZN({ S15143 })
);
NAND3_X1 #() 
NAND3_X1_3168_ (
  .A1({ S15143 }),
  .A2({ S15049 }),
  .A3({ S14504 }),
  .ZN({ S15154 })
);
NAND3_X1 #() 
NAND3_X1_3169_ (
  .A1({ S15040 }),
  .A2({ S14763 }),
  .A3({ S25956[108] }),
  .ZN({ S15165 })
);
NAND3_X1 #() 
NAND3_X1_3170_ (
  .A1({ S15135 }),
  .A2({ S15115 }),
  .A3({ S14515 }),
  .ZN({ S15176 })
);
NAND3_X1 #() 
NAND3_X1_3171_ (
  .A1({ S15176 }),
  .A2({ S15165 }),
  .A3({ S25956[76] }),
  .ZN({ S15187 })
);
AOI21_X1 #() 
AOI21_X1_1623_ (
  .A({ S25956[44] }),
  .B1({ S15154 }),
  .B2({ S15187 }),
  .ZN({ S15198 })
);
INV_X1 #() 
INV_X1_968_ (
  .A({ S25956[44] }),
  .ZN({ S15209 })
);
NAND3_X1 #() 
NAND3_X1_3172_ (
  .A1({ S15176 }),
  .A2({ S15165 }),
  .A3({ S14504 }),
  .ZN({ S15219 })
);
NAND3_X1 #() 
NAND3_X1_3173_ (
  .A1({ S15143 }),
  .A2({ S15049 }),
  .A3({ S25956[76] }),
  .ZN({ S15228 })
);
AOI21_X1 #() 
AOI21_X1_1624_ (
  .A({ S15209 }),
  .B1({ S15219 }),
  .B2({ S15228 }),
  .ZN({ S15239 })
);
OAI21_X1 #() 
OAI21_X1_1550_ (
  .A({ S25956[12] }),
  .B1({ S15198 }),
  .B2({ S15239 }),
  .ZN({ S15250 })
);
NAND3_X1 #() 
NAND3_X1_3174_ (
  .A1({ S15219 }),
  .A2({ S15228 }),
  .A3({ S15209 }),
  .ZN({ S15261 })
);
NAND3_X1 #() 
NAND3_X1_3175_ (
  .A1({ S15154 }),
  .A2({ S15187 }),
  .A3({ S25956[44] }),
  .ZN({ S15272 })
);
NAND3_X1 #() 
NAND3_X1_3176_ (
  .A1({ S15261 }),
  .A2({ S15272 }),
  .A3({ S5708 }),
  .ZN({ S15283 })
);
NAND2_X1 #() 
NAND2_X1_2951_ (
  .A1({ S15250 }),
  .A2({ S15283 }),
  .ZN({ S25957[1164] })
);
INV_X1 #() 
INV_X1_969_ (
  .A({ S25956[75] }),
  .ZN({ S15304 })
);
INV_X1 #() 
INV_X1_970_ (
  .A({ S25956[107] }),
  .ZN({ S15313 })
);
OAI211_X1 #() 
OAI211_X1_1033_ (
  .A({ S56 }),
  .B({ S25956[3] }),
  .C1({ S25956[2] }),
  .C2({ S11766 }),
  .ZN({ S15324 })
);
NAND3_X1 #() 
NAND3_X1_3177_ (
  .A1({ S15324 }),
  .A2({ S14073 }),
  .A3({ S25956[4] }),
  .ZN({ S15335 })
);
AOI21_X1 #() 
AOI21_X1_1625_ (
  .A({ S25956[4] }),
  .B1({ S13839 }),
  .B2({ S25956[0] }),
  .ZN({ S15346 })
);
NAND4_X1 #() 
NAND4_X1_347_ (
  .A1({ S15346 }),
  .A2({ S13120 }),
  .A3({ S11842 }),
  .A4({ S11864 }),
  .ZN({ S15357 })
);
NAND3_X1 #() 
NAND3_X1_3178_ (
  .A1({ S15335 }),
  .A2({ S15357 }),
  .A3({ S11631 }),
  .ZN({ S15368 })
);
NAND2_X1 #() 
NAND2_X1_2952_ (
  .A1({ S11917 }),
  .A2({ S25956[4] }),
  .ZN({ S15379 })
);
NAND4_X1 #() 
NAND4_X1_348_ (
  .A1({ S13238 }),
  .A2({ S11653 }),
  .A3({ S12118 }),
  .A4({ S25956[0] }),
  .ZN({ S15390 })
);
OAI211_X1 #() 
OAI211_X1_1034_ (
  .A({ S15390 }),
  .B({ S25956[5] }),
  .C1({ S15379 }),
  .C2({ S12221 }),
  .ZN({ S15397 })
);
NAND3_X1 #() 
NAND3_X1_3179_ (
  .A1({ S15368 }),
  .A2({ S11620 }),
  .A3({ S15397 }),
  .ZN({ S15408 })
);
NAND3_X1 #() 
NAND3_X1_3180_ (
  .A1({ S13022 }),
  .A2({ S25956[4] }),
  .A3({ S12182 }),
  .ZN({ S15419 })
);
AOI21_X1 #() 
AOI21_X1_1626_ (
  .A({ S25956[3] }),
  .B1({ S11642 }),
  .B2({ S25956[1] }),
  .ZN({ S15430 })
);
AOI22_X1 #() 
AOI22_X1_339_ (
  .A1({ S15430 }),
  .A2({ S11727 }),
  .B1({ S12303 }),
  .B2({ S25956[3] }),
  .ZN({ S15441 })
);
AOI21_X1 #() 
AOI21_X1_1627_ (
  .A({ S11631 }),
  .B1({ S15441 }),
  .B2({ S12118 }),
  .ZN({ S15452 })
);
NAND2_X1 #() 
NAND2_X1_2953_ (
  .A1({ S15419 }),
  .A2({ S15452 }),
  .ZN({ S15462 })
);
NAND3_X1 #() 
NAND3_X1_3181_ (
  .A1({ S11766 }),
  .A2({ S12655 }),
  .A3({ S11664 }),
  .ZN({ S15473 })
);
NAND2_X1 #() 
NAND2_X1_2954_ (
  .A1({ S15473 }),
  .A2({ S25956[4] }),
  .ZN({ S15484 })
);
AOI21_X1 #() 
AOI21_X1_1628_ (
  .A({ S25956[3] }),
  .B1({ S11766 }),
  .B2({ S25956[2] }),
  .ZN({ S15495 })
);
NAND2_X1 #() 
NAND2_X1_2955_ (
  .A1({ S15495 }),
  .A2({ S13205 }),
  .ZN({ S15506 })
);
NAND3_X1 #() 
NAND3_X1_3182_ (
  .A1({ S12357 }),
  .A2({ S15506 }),
  .A3({ S12118 }),
  .ZN({ S15516 })
);
NAND3_X1 #() 
NAND3_X1_3183_ (
  .A1({ S15516 }),
  .A2({ S11631 }),
  .A3({ S15484 }),
  .ZN({ S15525 })
);
NAND3_X1 #() 
NAND3_X1_3184_ (
  .A1({ S15462 }),
  .A2({ S25956[6] }),
  .A3({ S15525 }),
  .ZN({ S15536 })
);
NAND3_X1 #() 
NAND3_X1_3185_ (
  .A1({ S15536 }),
  .A2({ S11609 }),
  .A3({ S15408 }),
  .ZN({ S15547 })
);
INV_X1 #() 
INV_X1_971_ (
  .A({ S12490 }),
  .ZN({ S15558 })
);
NAND2_X1 #() 
NAND2_X1_2956_ (
  .A1({ S12563 }),
  .A2({ S56 }),
  .ZN({ S15569 })
);
NAND3_X1 #() 
NAND3_X1_3186_ (
  .A1({ S11727 }),
  .A2({ S11788 }),
  .A3({ S13839 }),
  .ZN({ S15580 })
);
NAND3_X1 #() 
NAND3_X1_3187_ (
  .A1({ S15569 }),
  .A2({ S15558 }),
  .A3({ S15580 }),
  .ZN({ S15591 })
);
NAND2_X1 #() 
NAND2_X1_2957_ (
  .A1({ S15591 }),
  .A2({ S12118 }),
  .ZN({ S15602 })
);
NAND2_X1 #() 
NAND2_X1_2958_ (
  .A1({ S11799 }),
  .A2({ S25956[3] }),
  .ZN({ S15613 })
);
NAND3_X1 #() 
NAND3_X1_3188_ (
  .A1({ S15613 }),
  .A2({ S25956[4] }),
  .A3({ S14945 }),
  .ZN({ S15624 })
);
NAND3_X1 #() 
NAND3_X1_3189_ (
  .A1({ S15602 }),
  .A2({ S15624 }),
  .A3({ S11631 }),
  .ZN({ S15635 })
);
NAND2_X1 #() 
NAND2_X1_2959_ (
  .A1({ S13011 }),
  .A2({ S11664 }),
  .ZN({ S15643 })
);
NAND3_X1 #() 
NAND3_X1_3190_ (
  .A1({ S12520 }),
  .A2({ S25956[3] }),
  .A3({ S11906 }),
  .ZN({ S15654 })
);
NAND3_X1 #() 
NAND3_X1_3191_ (
  .A1({ S15643 }),
  .A2({ S15654 }),
  .A3({ S25956[4] }),
  .ZN({ S15665 })
);
OAI211_X1 #() 
OAI211_X1_1035_ (
  .A({ S11664 }),
  .B({ S12097 }),
  .C1({ S12160 }),
  .C2({ S58 }),
  .ZN({ S15676 })
);
NAND3_X1 #() 
NAND3_X1_3192_ (
  .A1({ S13161 }),
  .A2({ S11777 }),
  .A3({ S25956[3] }),
  .ZN({ S15687 })
);
NAND3_X1 #() 
NAND3_X1_3193_ (
  .A1({ S15676 }),
  .A2({ S15687 }),
  .A3({ S12118 }),
  .ZN({ S15698 })
);
NAND3_X1 #() 
NAND3_X1_3194_ (
  .A1({ S15665 }),
  .A2({ S25956[5] }),
  .A3({ S15698 }),
  .ZN({ S15709 })
);
NAND3_X1 #() 
NAND3_X1_3195_ (
  .A1({ S15635 }),
  .A2({ S15709 }),
  .A3({ S11620 }),
  .ZN({ S15720 })
);
NAND2_X1 #() 
NAND2_X1_2960_ (
  .A1({ S11766 }),
  .A2({ S11853 }),
  .ZN({ S15730 })
);
AOI21_X1 #() 
AOI21_X1_1629_ (
  .A({ S25956[1] }),
  .B1({ S25956[2] }),
  .B2({ S25956[0] }),
  .ZN({ S15737 })
);
NOR2_X1 #() 
NOR2_X1_741_ (
  .A1({ S15730 }),
  .A2({ S15737 }),
  .ZN({ S15748 })
);
NOR2_X1 #() 
NOR2_X1_742_ (
  .A1({ S11550 }),
  .A2({ S25956[1] }),
  .ZN({ S15759 })
);
NOR2_X1 #() 
NOR2_X1_743_ (
  .A1({ S15759 }),
  .A2({ S25956[3] }),
  .ZN({ S15770 })
);
AOI22_X1 #() 
AOI22_X1_340_ (
  .A1({ S15748 }),
  .A2({ S25956[3] }),
  .B1({ S15770 }),
  .B2({ S13055 }),
  .ZN({ S15781 })
);
NAND3_X1 #() 
NAND3_X1_3196_ (
  .A1({ S11950 }),
  .A2({ S11664 }),
  .A3({ S11727 }),
  .ZN({ S15792 })
);
NAND3_X1 #() 
NAND3_X1_3197_ (
  .A1({ S15792 }),
  .A2({ S14650 }),
  .A3({ S25956[4] }),
  .ZN({ S15803 })
);
OAI211_X1 #() 
OAI211_X1_1036_ (
  .A({ S15803 }),
  .B({ S25956[5] }),
  .C1({ S15781 }),
  .C2({ S25956[4] }),
  .ZN({ S15814 })
);
OAI211_X1 #() 
OAI211_X1_1037_ (
  .A({ S13205 }),
  .B({ S11664 }),
  .C1({ S11777 }),
  .C2({ S13395 }),
  .ZN({ S15825 })
);
AOI21_X1 #() 
AOI21_X1_1630_ (
  .A({ S12118 }),
  .B1({ S15730 }),
  .B2({ S25956[3] }),
  .ZN({ S15833 })
);
NAND2_X1 #() 
NAND2_X1_2961_ (
  .A1({ S15825 }),
  .A2({ S15833 }),
  .ZN({ S15844 })
);
NAND2_X1 #() 
NAND2_X1_2962_ (
  .A1({ S11788 }),
  .A2({ S12655 }),
  .ZN({ S15855 })
);
AOI21_X1 #() 
AOI21_X1_1631_ (
  .A({ S25956[5] }),
  .B1({ S15855 }),
  .B2({ S14534 }),
  .ZN({ S15866 })
);
AOI21_X1 #() 
AOI21_X1_1632_ (
  .A({ S11620 }),
  .B1({ S15844 }),
  .B2({ S15866 }),
  .ZN({ S15877 })
);
NAND2_X1 #() 
NAND2_X1_2963_ (
  .A1({ S15814 }),
  .A2({ S15877 }),
  .ZN({ S15888 })
);
NAND2_X1 #() 
NAND2_X1_2964_ (
  .A1({ S15720 }),
  .A2({ S15888 }),
  .ZN({ S15899 })
);
NAND2_X1 #() 
NAND2_X1_2965_ (
  .A1({ S15899 }),
  .A2({ S25956[7] }),
  .ZN({ S15908 })
);
NAND3_X1 #() 
NAND3_X1_3198_ (
  .A1({ S15908 }),
  .A2({ S15313 }),
  .A3({ S15547 }),
  .ZN({ S15915 })
);
AND3_X1 #() 
AND3_X1_123_ (
  .A1({ S15536 }),
  .A2({ S15408 }),
  .A3({ S11609 }),
  .ZN({ S15926 })
);
AOI21_X1 #() 
AOI21_X1_1633_ (
  .A({ S11609 }),
  .B1({ S15720 }),
  .B2({ S15888 }),
  .ZN({ S15937 })
);
OAI21_X1 #() 
OAI21_X1_1551_ (
  .A({ S25956[107] }),
  .B1({ S15937 }),
  .B2({ S15926 }),
  .ZN({ S15948 })
);
NAND3_X1 #() 
NAND3_X1_3199_ (
  .A1({ S15915 }),
  .A2({ S15948 }),
  .A3({ S15304 }),
  .ZN({ S15959 })
);
NAND3_X1 #() 
NAND3_X1_3200_ (
  .A1({ S15908 }),
  .A2({ S25956[107] }),
  .A3({ S15547 }),
  .ZN({ S15970 })
);
OAI21_X1 #() 
OAI21_X1_1552_ (
  .A({ S15313 }),
  .B1({ S15937 }),
  .B2({ S15926 }),
  .ZN({ S15981 })
);
NAND3_X1 #() 
NAND3_X1_3201_ (
  .A1({ S15970 }),
  .A2({ S15981 }),
  .A3({ S25956[75] }),
  .ZN({ S15992 })
);
AOI21_X1 #() 
AOI21_X1_1634_ (
  .A({ S25956[43] }),
  .B1({ S15959 }),
  .B2({ S15992 }),
  .ZN({ S16000 })
);
INV_X1 #() 
INV_X1_972_ (
  .A({ S25956[43] }),
  .ZN({ S16009 })
);
NAND3_X1 #() 
NAND3_X1_3202_ (
  .A1({ S15970 }),
  .A2({ S15981 }),
  .A3({ S15304 }),
  .ZN({ S16020 })
);
NAND3_X1 #() 
NAND3_X1_3203_ (
  .A1({ S15915 }),
  .A2({ S15948 }),
  .A3({ S25956[75] }),
  .ZN({ S16031 })
);
AOI21_X1 #() 
AOI21_X1_1635_ (
  .A({ S16009 }),
  .B1({ S16020 }),
  .B2({ S16031 }),
  .ZN({ S16042 })
);
OAI21_X1 #() 
OAI21_X1_1553_ (
  .A({ S5719 }),
  .B1({ S16000 }),
  .B2({ S16042 }),
  .ZN({ S16053 })
);
NAND3_X1 #() 
NAND3_X1_3204_ (
  .A1({ S16020 }),
  .A2({ S16031 }),
  .A3({ S16009 }),
  .ZN({ S16064 })
);
NAND3_X1 #() 
NAND3_X1_3205_ (
  .A1({ S15959 }),
  .A2({ S15992 }),
  .A3({ S25956[43] }),
  .ZN({ S16075 })
);
NAND3_X1 #() 
NAND3_X1_3206_ (
  .A1({ S16064 }),
  .A2({ S16075 }),
  .A3({ S25956[11] }),
  .ZN({ S16086 })
);
NAND2_X1 #() 
NAND2_X1_2966_ (
  .A1({ S16053 }),
  .A2({ S16086 }),
  .ZN({ S65 })
);
OAI21_X1 #() 
OAI21_X1_1554_ (
  .A({ S25956[11] }),
  .B1({ S16000 }),
  .B2({ S16042 }),
  .ZN({ S16104 })
);
NAND3_X1 #() 
NAND3_X1_3207_ (
  .A1({ S16064 }),
  .A2({ S16075 }),
  .A3({ S5719 }),
  .ZN({ S16114 })
);
NAND2_X1 #() 
NAND2_X1_2967_ (
  .A1({ S16104 }),
  .A2({ S16114 }),
  .ZN({ S25957[1163] })
);
INV_X1 #() 
INV_X1_973_ (
  .A({ S25956[72] }),
  .ZN({ S16135 })
);
INV_X1 #() 
INV_X1_974_ (
  .A({ S25956[104] }),
  .ZN({ S16146 })
);
NAND2_X1 #() 
NAND2_X1_2968_ (
  .A1({ S13417 }),
  .A2({ S11664 }),
  .ZN({ S16157 })
);
NAND3_X1 #() 
NAND3_X1_3208_ (
  .A1({ S14256 }),
  .A2({ S16157 }),
  .A3({ S12118 }),
  .ZN({ S16168 })
);
OAI21_X1 #() 
OAI21_X1_1555_ (
  .A({ S11664 }),
  .B1({ S15730 }),
  .B2({ S15737 }),
  .ZN({ S16178 })
);
NAND3_X1 #() 
NAND3_X1_3209_ (
  .A1({ S16178 }),
  .A2({ S25956[4] }),
  .A3({ S15580 }),
  .ZN({ S16186 })
);
NAND3_X1 #() 
NAND3_X1_3210_ (
  .A1({ S16186 }),
  .A2({ S11631 }),
  .A3({ S16168 }),
  .ZN({ S16193 })
);
NAND3_X1 #() 
NAND3_X1_3211_ (
  .A1({ S56 }),
  .A2({ S11766 }),
  .A3({ S11736 }),
  .ZN({ S16204 })
);
AND2_X1 #() 
AND2_X1_192_ (
  .A1({ S25956[1] }),
  .A2({ S25956[2] }),
  .ZN({ S16215 })
);
NAND2_X1 #() 
NAND2_X1_2969_ (
  .A1({ S16215 }),
  .A2({ S11664 }),
  .ZN({ S16226 })
);
NAND4_X1 #() 
NAND4_X1_349_ (
  .A1({ S14671 }),
  .A2({ S16204 }),
  .A3({ S12118 }),
  .A4({ S16226 }),
  .ZN({ S16237 })
);
AOI21_X1 #() 
AOI21_X1_1636_ (
  .A({ S12118 }),
  .B1({ S11788 }),
  .B2({ S13839 }),
  .ZN({ S16248 })
);
AOI21_X1 #() 
AOI21_X1_1637_ (
  .A({ S11631 }),
  .B1({ S14639 }),
  .B2({ S16248 }),
  .ZN({ S16257 })
);
NAND2_X1 #() 
NAND2_X1_2970_ (
  .A1({ S16257 }),
  .A2({ S16237 }),
  .ZN({ S16258 })
);
NAND3_X1 #() 
NAND3_X1_3212_ (
  .A1({ S16193 }),
  .A2({ S25956[6] }),
  .A3({ S16258 }),
  .ZN({ S16259 })
);
NAND3_X1 #() 
NAND3_X1_3213_ (
  .A1({ S14975 }),
  .A2({ S14857 }),
  .A3({ S13142 }),
  .ZN({ S16261 })
);
OAI21_X1 #() 
OAI21_X1_1556_ (
  .A({ S15473 }),
  .B1({ S12201 }),
  .B2({ S11664 }),
  .ZN({ S16263 })
);
AOI21_X1 #() 
AOI21_X1_1638_ (
  .A({ S12118 }),
  .B1({ S12053 }),
  .B2({ S11550 }),
  .ZN({ S16264 })
);
AOI22_X1 #() 
AOI22_X1_341_ (
  .A1({ S16261 }),
  .A2({ S12118 }),
  .B1({ S16263 }),
  .B2({ S16264 }),
  .ZN({ S16265 })
);
AOI22_X1 #() 
AOI22_X1_342_ (
  .A1({ S11853 }),
  .A2({ S11550 }),
  .B1({ S12655 }),
  .B2({ S11664 }),
  .ZN({ S16267 })
);
NAND2_X1 #() 
NAND2_X1_2971_ (
  .A1({ S11864 }),
  .A2({ S12118 }),
  .ZN({ S16268 })
);
NOR2_X1 #() 
NOR2_X1_744_ (
  .A1({ S16268 }),
  .A2({ S16267 }),
  .ZN({ S16270 })
);
NOR2_X1 #() 
NOR2_X1_745_ (
  .A1({ S58 }),
  .A2({ S13395 }),
  .ZN({ S16273 })
);
AOI21_X1 #() 
AOI21_X1_1639_ (
  .A({ S13525 }),
  .B1({ S16273 }),
  .B2({ S11736 }),
  .ZN({ S16276 })
);
OAI21_X1 #() 
OAI21_X1_1557_ (
  .A({ S11631 }),
  .B1({ S16270 }),
  .B2({ S16276 }),
  .ZN({ S16277 })
);
OAI211_X1 #() 
OAI211_X1_1038_ (
  .A({ S16277 }),
  .B({ S11620 }),
  .C1({ S16265 }),
  .C2({ S11631 }),
  .ZN({ S16280 })
);
NAND3_X1 #() 
NAND3_X1_3214_ (
  .A1({ S16280 }),
  .A2({ S25956[7] }),
  .A3({ S16259 }),
  .ZN({ S16283 })
);
NAND2_X1 #() 
NAND2_X1_2972_ (
  .A1({ S13161 }),
  .A2({ S11950 }),
  .ZN({ S16288 })
);
NAND2_X1 #() 
NAND2_X1_2973_ (
  .A1({ S16288 }),
  .A2({ S25956[3] }),
  .ZN({ S16292 })
);
NAND4_X1 #() 
NAND4_X1_350_ (
  .A1({ S11906 }),
  .A2({ S12042 }),
  .A3({ S25956[3] }),
  .A4({ S14053 }),
  .ZN({ S16297 })
);
AOI21_X1 #() 
AOI21_X1_1640_ (
  .A({ S12118 }),
  .B1({ S13055 }),
  .B2({ S11664 }),
  .ZN({ S16298 })
);
AOI22_X1 #() 
AOI22_X1_343_ (
  .A1({ S16292 }),
  .A2({ S12622 }),
  .B1({ S16297 }),
  .B2({ S16298 }),
  .ZN({ S16303 })
);
OAI21_X1 #() 
OAI21_X1_1558_ (
  .A({ S11664 }),
  .B1({ S11821 }),
  .B2({ S25956[1] }),
  .ZN({ S16309 })
);
NAND3_X1 #() 
NAND3_X1_3215_ (
  .A1({ S14256 }),
  .A2({ S12118 }),
  .A3({ S16309 }),
  .ZN({ S16313 })
);
NAND4_X1 #() 
NAND4_X1_351_ (
  .A1({ S14095 }),
  .A2({ S13417 }),
  .A3({ S25956[4] }),
  .A4({ S12388 }),
  .ZN({ S16315 })
);
NAND3_X1 #() 
NAND3_X1_3216_ (
  .A1({ S16313 }),
  .A2({ S11631 }),
  .A3({ S16315 }),
  .ZN({ S16319 })
);
OAI211_X1 #() 
OAI211_X1_1039_ (
  .A({ S16319 }),
  .B({ S25956[6] }),
  .C1({ S16303 }),
  .C2({ S11631 }),
  .ZN({ S16324 })
);
NAND3_X1 #() 
NAND3_X1_3217_ (
  .A1({ S13205 }),
  .A2({ S11664 }),
  .A3({ S12160 }),
  .ZN({ S16327 })
);
OAI211_X1 #() 
OAI211_X1_1040_ (
  .A({ S11788 }),
  .B({ S25956[3] }),
  .C1({ S16215 }),
  .C2({ S13395 }),
  .ZN({ S16332 })
);
NAND2_X1 #() 
NAND2_X1_2974_ (
  .A1({ S16327 }),
  .A2({ S16332 }),
  .ZN({ S16341 })
);
AOI21_X1 #() 
AOI21_X1_1641_ (
  .A({ S25956[3] }),
  .B1({ S12655 }),
  .B2({ S11539 }),
  .ZN({ S16352 })
);
AOI21_X1 #() 
AOI21_X1_1642_ (
  .A({ S12118 }),
  .B1({ S16352 }),
  .B2({ S14053 }),
  .ZN({ S16363 })
);
AOI22_X1 #() 
AOI22_X1_344_ (
  .A1({ S16341 }),
  .A2({ S12118 }),
  .B1({ S16363 }),
  .B2({ S12552 }),
  .ZN({ S16374 })
);
NAND3_X1 #() 
NAND3_X1_3218_ (
  .A1({ S14106 }),
  .A2({ S14650 }),
  .A3({ S25956[4] }),
  .ZN({ S16385 })
);
NAND3_X1 #() 
NAND3_X1_3219_ (
  .A1({ S14146 }),
  .A2({ S12118 }),
  .A3({ S13302 }),
  .ZN({ S16396 })
);
NAND3_X1 #() 
NAND3_X1_3220_ (
  .A1({ S16396 }),
  .A2({ S16385 }),
  .A3({ S25956[5] }),
  .ZN({ S16407 })
);
OAI211_X1 #() 
OAI211_X1_1041_ (
  .A({ S16407 }),
  .B({ S11620 }),
  .C1({ S16374 }),
  .C2({ S25956[5] }),
  .ZN({ S16418 })
);
NAND3_X1 #() 
NAND3_X1_3221_ (
  .A1({ S16418 }),
  .A2({ S11609 }),
  .A3({ S16324 }),
  .ZN({ S16429 })
);
NAND3_X1 #() 
NAND3_X1_3222_ (
  .A1({ S16429 }),
  .A2({ S16283 }),
  .A3({ S16146 }),
  .ZN({ S16440 })
);
NAND2_X1 #() 
NAND2_X1_2975_ (
  .A1({ S16429 }),
  .A2({ S16283 }),
  .ZN({ S16451 })
);
NAND2_X1 #() 
NAND2_X1_2976_ (
  .A1({ S16451 }),
  .A2({ S25956[104] }),
  .ZN({ S16462 })
);
NAND3_X1 #() 
NAND3_X1_3223_ (
  .A1({ S16462 }),
  .A2({ S16135 }),
  .A3({ S16440 }),
  .ZN({ S16473 })
);
NAND3_X1 #() 
NAND3_X1_3224_ (
  .A1({ S16429 }),
  .A2({ S16283 }),
  .A3({ S25956[104] }),
  .ZN({ S16484 })
);
NAND2_X1 #() 
NAND2_X1_2977_ (
  .A1({ S16451 }),
  .A2({ S16146 }),
  .ZN({ S16495 })
);
NAND3_X1 #() 
NAND3_X1_3225_ (
  .A1({ S16495 }),
  .A2({ S25956[72] }),
  .A3({ S16484 }),
  .ZN({ S16505 })
);
AOI21_X1 #() 
AOI21_X1_1643_ (
  .A({ S25956[40] }),
  .B1({ S16473 }),
  .B2({ S16505 }),
  .ZN({ S16516 })
);
INV_X1 #() 
INV_X1_975_ (
  .A({ S25956[40] }),
  .ZN({ S16527 })
);
NAND3_X1 #() 
NAND3_X1_3226_ (
  .A1({ S16495 }),
  .A2({ S16135 }),
  .A3({ S16484 }),
  .ZN({ S16538 })
);
NAND3_X1 #() 
NAND3_X1_3227_ (
  .A1({ S16462 }),
  .A2({ S25956[72] }),
  .A3({ S16440 }),
  .ZN({ S16549 })
);
AOI21_X1 #() 
AOI21_X1_1644_ (
  .A({ S16527 }),
  .B1({ S16538 }),
  .B2({ S16549 }),
  .ZN({ S16560 })
);
OAI21_X1 #() 
OAI21_X1_1559_ (
  .A({ S25956[8] }),
  .B1({ S16516 }),
  .B2({ S16560 }),
  .ZN({ S16571 })
);
NAND3_X1 #() 
NAND3_X1_3228_ (
  .A1({ S16538 }),
  .A2({ S16549 }),
  .A3({ S16527 }),
  .ZN({ S16582 })
);
NAND3_X1 #() 
NAND3_X1_3229_ (
  .A1({ S16473 }),
  .A2({ S16505 }),
  .A3({ S25956[40] }),
  .ZN({ S16592 })
);
NAND3_X1 #() 
NAND3_X1_3230_ (
  .A1({ S16582 }),
  .A2({ S16592 }),
  .A3({ S5639 }),
  .ZN({ S16603 })
);
NAND2_X1 #() 
NAND2_X1_2978_ (
  .A1({ S16571 }),
  .A2({ S16603 }),
  .ZN({ S25957[1160] })
);
INV_X1 #() 
INV_X1_976_ (
  .A({ S25956[73] }),
  .ZN({ S16624 })
);
INV_X1 #() 
INV_X1_977_ (
  .A({ S25956[105] }),
  .ZN({ S16635 })
);
NAND3_X1 #() 
NAND3_X1_3231_ (
  .A1({ S11906 }),
  .A2({ S25956[3] }),
  .A3({ S14053 }),
  .ZN({ S16646 })
);
NAND3_X1 #() 
NAND3_X1_3232_ (
  .A1({ S12928 }),
  .A2({ S12118 }),
  .A3({ S16646 }),
  .ZN({ S16657 })
);
NOR2_X1 #() 
NOR2_X1_746_ (
  .A1({ S25956[2] }),
  .A2({ S25956[0] }),
  .ZN({ S16667 })
);
AOI21_X1 #() 
AOI21_X1_1645_ (
  .A({ S16667 }),
  .B1({ S15737 }),
  .B2({ S25956[3] }),
  .ZN({ S16678 })
);
OAI211_X1 #() 
OAI211_X1_1042_ (
  .A({ S25956[4] }),
  .B({ S14053 }),
  .C1({ S16678 }),
  .C2({ S11832 }),
  .ZN({ S16689 })
);
NAND3_X1 #() 
NAND3_X1_3233_ (
  .A1({ S16657 }),
  .A2({ S11631 }),
  .A3({ S16689 }),
  .ZN({ S16700 })
);
NOR2_X1 #() 
NOR2_X1_747_ (
  .A1({ S16273 }),
  .A2({ S13450 }),
  .ZN({ S16711 })
);
AOI21_X1 #() 
AOI21_X1_1646_ (
  .A({ S25956[3] }),
  .B1({ S11939 }),
  .B2({ S12160 }),
  .ZN({ S16722 })
);
OAI21_X1 #() 
OAI21_X1_1560_ (
  .A({ S25956[4] }),
  .B1({ S16711 }),
  .B2({ S16722 }),
  .ZN({ S16733 })
);
OAI21_X1 #() 
OAI21_X1_1561_ (
  .A({ S25956[5] }),
  .B1({ S12655 }),
  .B2({ S25956[4] }),
  .ZN({ S16743 })
);
AOI21_X1 #() 
AOI21_X1_1647_ (
  .A({ S16743 }),
  .B1({ S12622 }),
  .B2({ S11539 }),
  .ZN({ S16754 })
);
AOI21_X1 #() 
AOI21_X1_1648_ (
  .A({ S11620 }),
  .B1({ S16733 }),
  .B2({ S16754 }),
  .ZN({ S16765 })
);
AOI21_X1 #() 
AOI21_X1_1649_ (
  .A({ S12490 }),
  .B1({ S15495 }),
  .B2({ S13205 }),
  .ZN({ S16776 })
);
OAI211_X1 #() 
OAI211_X1_1043_ (
  .A({ S13872 }),
  .B({ S12655 }),
  .C1({ S11653 }),
  .C2({ S25956[3] }),
  .ZN({ S16787 })
);
NAND2_X1 #() 
NAND2_X1_2979_ (
  .A1({ S16787 }),
  .A2({ S25956[4] }),
  .ZN({ S16797 })
);
OAI211_X1 #() 
OAI211_X1_1044_ (
  .A({ S16797 }),
  .B({ S11631 }),
  .C1({ S16776 }),
  .C2({ S25956[4] }),
  .ZN({ S16808 })
);
NOR2_X1 #() 
NOR2_X1_748_ (
  .A1({ S14997 }),
  .A2({ S25956[0] }),
  .ZN({ S16819 })
);
AOI21_X1 #() 
AOI21_X1_1650_ (
  .A({ S11664 }),
  .B1({ S13417 }),
  .B2({ S14053 }),
  .ZN({ S16830 })
);
OAI21_X1 #() 
OAI21_X1_1562_ (
  .A({ S25956[4] }),
  .B1({ S16830 }),
  .B2({ S16819 }),
  .ZN({ S16841 })
);
AOI21_X1 #() 
AOI21_X1_1651_ (
  .A({ S11631 }),
  .B1({ S11716 }),
  .B2({ S11744 }),
  .ZN({ S16852 })
);
AOI21_X1 #() 
AOI21_X1_1652_ (
  .A({ S25956[6] }),
  .B1({ S16841 }),
  .B2({ S16852 }),
  .ZN({ S16862 })
);
AOI22_X1 #() 
AOI22_X1_345_ (
  .A1({ S16765 }),
  .A2({ S16700 }),
  .B1({ S16862 }),
  .B2({ S16808 }),
  .ZN({ S16873 })
);
INV_X1 #() 
INV_X1_978_ (
  .A({ S12303 }),
  .ZN({ S16884 })
);
AOI21_X1 #() 
AOI21_X1_1653_ (
  .A({ S11664 }),
  .B1({ S16884 }),
  .B2({ S14053 }),
  .ZN({ S16895 })
);
OAI211_X1 #() 
OAI211_X1_1045_ (
  .A({ S14534 }),
  .B({ S13142 }),
  .C1({ S14997 }),
  .C2({ S15759 }),
  .ZN({ S16906 })
);
OAI211_X1 #() 
OAI211_X1_1046_ (
  .A({ S16906 }),
  .B({ S25956[5] }),
  .C1({ S11971 }),
  .C2({ S16895 }),
  .ZN({ S16916 })
);
NOR2_X1 #() 
NOR2_X1_749_ (
  .A1({ S11810 }),
  .A2({ S14796 }),
  .ZN({ S16927 })
);
AOI21_X1 #() 
AOI21_X1_1654_ (
  .A({ S25956[3] }),
  .B1({ S12097 }),
  .B2({ S12347 }),
  .ZN({ S16938 })
);
OAI21_X1 #() 
OAI21_X1_1563_ (
  .A({ S11631 }),
  .B1({ S16938 }),
  .B2({ S13077 }),
  .ZN({ S16949 })
);
OAI211_X1 #() 
OAI211_X1_1047_ (
  .A({ S16916 }),
  .B({ S11620 }),
  .C1({ S16927 }),
  .C2({ S16949 }),
  .ZN({ S16960 })
);
OAI211_X1 #() 
OAI211_X1_1048_ (
  .A({ S13935 }),
  .B({ S25956[4] }),
  .C1({ S11705 }),
  .C2({ S25956[3] }),
  .ZN({ S16968 })
);
AOI21_X1 #() 
AOI21_X1_1655_ (
  .A({ S25956[4] }),
  .B1({ S11950 }),
  .B2({ S11664 }),
  .ZN({ S16979 })
);
NAND2_X1 #() 
NAND2_X1_2980_ (
  .A1({ S16297 }),
  .A2({ S16979 }),
  .ZN({ S16990 })
);
NAND3_X1 #() 
NAND3_X1_3234_ (
  .A1({ S16990 }),
  .A2({ S25956[5] }),
  .A3({ S16968 }),
  .ZN({ S17001 })
);
NOR3_X1 #() 
NOR3_X1_106_ (
  .A1({ S25956[2] }),
  .A2({ S25956[1] }),
  .A3({ S25956[0] }),
  .ZN({ S17012 })
);
OAI211_X1 #() 
OAI211_X1_1049_ (
  .A({ S13120 }),
  .B({ S12118 }),
  .C1({ S15473 }),
  .C2({ S17012 }),
  .ZN({ S17023 })
);
NAND2_X1 #() 
NAND2_X1_2981_ (
  .A1({ S14064 }),
  .A2({ S16264 }),
  .ZN({ S17034 })
);
NAND3_X1 #() 
NAND3_X1_3235_ (
  .A1({ S17034 }),
  .A2({ S17023 }),
  .A3({ S11631 }),
  .ZN({ S17045 })
);
NAND3_X1 #() 
NAND3_X1_3236_ (
  .A1({ S17045 }),
  .A2({ S17001 }),
  .A3({ S25956[6] }),
  .ZN({ S17056 })
);
NAND3_X1 #() 
NAND3_X1_3237_ (
  .A1({ S16960 }),
  .A2({ S25956[7] }),
  .A3({ S17056 }),
  .ZN({ S17067 })
);
OAI211_X1 #() 
OAI211_X1_1050_ (
  .A({ S17067 }),
  .B({ S16635 }),
  .C1({ S16873 }),
  .C2({ S25956[7] }),
  .ZN({ S17078 })
);
XNOR2_X1 #() 
XNOR2_X1_158_ (
  .A({ S25956[1] }),
  .B({ S25956[0] }),
  .ZN({ S17089 })
);
NAND2_X1 #() 
NAND2_X1_2982_ (
  .A1({ S11939 }),
  .A2({ S12160 }),
  .ZN({ S17100 })
);
AOI22_X1 #() 
AOI22_X1_346_ (
  .A1({ S17100 }),
  .A2({ S11664 }),
  .B1({ S17089 }),
  .B2({ S11672 }),
  .ZN({ S17110 })
);
OAI21_X1 #() 
OAI21_X1_1564_ (
  .A({ S16754 }),
  .B1({ S17110 }),
  .B2({ S12118 }),
  .ZN({ S17121 })
);
NAND3_X1 #() 
NAND3_X1_3238_ (
  .A1({ S16700 }),
  .A2({ S17121 }),
  .A3({ S25956[6] }),
  .ZN({ S17132 })
);
NAND2_X1 #() 
NAND2_X1_2983_ (
  .A1({ S16841 }),
  .A2({ S16852 }),
  .ZN({ S17143 })
);
NAND3_X1 #() 
NAND3_X1_3239_ (
  .A1({ S17143 }),
  .A2({ S16808 }),
  .A3({ S11620 }),
  .ZN({ S17154 })
);
AOI21_X1 #() 
AOI21_X1_1656_ (
  .A({ S25956[7] }),
  .B1({ S17132 }),
  .B2({ S17154 }),
  .ZN({ S17165 })
);
AND3_X1 #() 
AND3_X1_124_ (
  .A1({ S16960 }),
  .A2({ S25956[7] }),
  .A3({ S17056 }),
  .ZN({ S17176 })
);
OAI21_X1 #() 
OAI21_X1_1565_ (
  .A({ S25956[105] }),
  .B1({ S17176 }),
  .B2({ S17165 }),
  .ZN({ S17186 })
);
NAND3_X1 #() 
NAND3_X1_3240_ (
  .A1({ S17186 }),
  .A2({ S16624 }),
  .A3({ S17078 }),
  .ZN({ S17197 })
);
OAI211_X1 #() 
OAI211_X1_1051_ (
  .A({ S17067 }),
  .B({ S25956[105] }),
  .C1({ S16873 }),
  .C2({ S25956[7] }),
  .ZN({ S17208 })
);
OAI21_X1 #() 
OAI21_X1_1566_ (
  .A({ S16635 }),
  .B1({ S17176 }),
  .B2({ S17165 }),
  .ZN({ S17219 })
);
NAND3_X1 #() 
NAND3_X1_3241_ (
  .A1({ S17219 }),
  .A2({ S25956[73] }),
  .A3({ S17208 }),
  .ZN({ S17230 })
);
AOI21_X1 #() 
AOI21_X1_1657_ (
  .A({ S25956[41] }),
  .B1({ S17197 }),
  .B2({ S17230 }),
  .ZN({ S17241 })
);
INV_X1 #() 
INV_X1_979_ (
  .A({ S25956[41] }),
  .ZN({ S17251 })
);
NAND3_X1 #() 
NAND3_X1_3242_ (
  .A1({ S17219 }),
  .A2({ S16624 }),
  .A3({ S17208 }),
  .ZN({ S17262 })
);
NAND3_X1 #() 
NAND3_X1_3243_ (
  .A1({ S17186 }),
  .A2({ S25956[73] }),
  .A3({ S17078 }),
  .ZN({ S17273 })
);
AOI21_X1 #() 
AOI21_X1_1658_ (
  .A({ S17251 }),
  .B1({ S17262 }),
  .B2({ S17273 }),
  .ZN({ S17284 })
);
OAI21_X1 #() 
OAI21_X1_1567_ (
  .A({ S25956[9] }),
  .B1({ S17241 }),
  .B2({ S17284 }),
  .ZN({ S17295 })
);
NAND3_X1 #() 
NAND3_X1_3244_ (
  .A1({ S17262 }),
  .A2({ S17273 }),
  .A3({ S17251 }),
  .ZN({ S17306 })
);
NAND3_X1 #() 
NAND3_X1_3245_ (
  .A1({ S17197 }),
  .A2({ S17230 }),
  .A3({ S25956[41] }),
  .ZN({ S17317 })
);
NAND3_X1 #() 
NAND3_X1_3246_ (
  .A1({ S17306 }),
  .A2({ S17317 }),
  .A3({ S5628 }),
  .ZN({ S17328 })
);
NAND2_X1 #() 
NAND2_X1_2984_ (
  .A1({ S17295 }),
  .A2({ S17328 }),
  .ZN({ S25957[1161] })
);
INV_X1 #() 
INV_X1_980_ (
  .A({ S25956[42] }),
  .ZN({ S17348 })
);
INV_X1 #() 
INV_X1_981_ (
  .A({ S25956[74] }),
  .ZN({ S17359 })
);
INV_X1 #() 
INV_X1_982_ (
  .A({ S25956[106] }),
  .ZN({ S17370 })
);
NAND3_X1 #() 
NAND3_X1_3247_ (
  .A1({ S12961 }),
  .A2({ S25956[3] }),
  .A3({ S25956[1] }),
  .ZN({ S17381 })
);
NAND3_X1 #() 
NAND3_X1_3248_ (
  .A1({ S12501 }),
  .A2({ S13161 }),
  .A3({ S11664 }),
  .ZN({ S17392 })
);
NAND3_X1 #() 
NAND3_X1_3249_ (
  .A1({ S17392 }),
  .A2({ S12118 }),
  .A3({ S17381 }),
  .ZN({ S17403 })
);
OAI211_X1 #() 
OAI211_X1_1052_ (
  .A({ S16226 }),
  .B({ S15473 }),
  .C1({ S14785 }),
  .C2({ S13450 }),
  .ZN({ S17413 })
);
NAND2_X1 #() 
NAND2_X1_2985_ (
  .A1({ S17413 }),
  .A2({ S25956[4] }),
  .ZN({ S17424 })
);
NAND3_X1 #() 
NAND3_X1_3250_ (
  .A1({ S17424 }),
  .A2({ S17403 }),
  .A3({ S25956[6] }),
  .ZN({ S17435 })
);
AND2_X1 #() 
AND2_X1_193_ (
  .A1({ S14817 }),
  .A2({ S17381 }),
  .ZN({ S17446 })
);
NAND2_X1 #() 
NAND2_X1_2986_ (
  .A1({ S11853 }),
  .A2({ S11664 }),
  .ZN({ S17457 })
);
AOI21_X1 #() 
AOI21_X1_1659_ (
  .A({ S17457 }),
  .B1({ S12512 }),
  .B2({ S56 }),
  .ZN({ S17467 })
);
OAI21_X1 #() 
OAI21_X1_1568_ (
  .A({ S12118 }),
  .B1({ S17467 }),
  .B2({ S13172 }),
  .ZN({ S17478 })
);
OAI211_X1 #() 
OAI211_X1_1053_ (
  .A({ S17478 }),
  .B({ S11620 }),
  .C1({ S17446 }),
  .C2({ S12118 }),
  .ZN({ S17489 })
);
AOI21_X1 #() 
AOI21_X1_1660_ (
  .A({ S25956[5] }),
  .B1({ S17489 }),
  .B2({ S17435 }),
  .ZN({ S17500 })
);
AOI21_X1 #() 
AOI21_X1_1661_ (
  .A({ S12442 }),
  .B1({ S13000 }),
  .B2({ S13033 }),
  .ZN({ S17511 })
);
NOR3_X1 #() 
NOR3_X1_107_ (
  .A1({ S12210 }),
  .A2({ S12512 }),
  .A3({ S11664 }),
  .ZN({ S17522 })
);
OAI21_X1 #() 
OAI21_X1_1569_ (
  .A({ S12118 }),
  .B1({ S11939 }),
  .B2({ S12644 }),
  .ZN({ S17532 })
);
OAI21_X1 #() 
OAI21_X1_1570_ (
  .A({ S25956[4] }),
  .B1({ S17012 }),
  .B2({ S13450 }),
  .ZN({ S17543 })
);
OAI22_X1 #() 
OAI22_X1_78_ (
  .A1({ S17511 }),
  .A2({ S17543 }),
  .B1({ S17522 }),
  .B2({ S17532 }),
  .ZN({ S17554 })
);
AOI21_X1 #() 
AOI21_X1_1662_ (
  .A({ S25956[4] }),
  .B1({ S15430 }),
  .B2({ S25956[0] }),
  .ZN({ S17565 })
);
NAND3_X1 #() 
NAND3_X1_3251_ (
  .A1({ S12581 }),
  .A2({ S17565 }),
  .A3({ S12552 }),
  .ZN({ S17574 })
);
OAI211_X1 #() 
OAI211_X1_1054_ (
  .A({ S12097 }),
  .B({ S25956[0] }),
  .C1({ S11539 }),
  .C2({ S11664 }),
  .ZN({ S17584 })
);
AOI21_X1 #() 
AOI21_X1_1663_ (
  .A({ S12118 }),
  .B1({ S12442 }),
  .B2({ S25956[3] }),
  .ZN({ S17595 })
);
AOI21_X1 #() 
AOI21_X1_1664_ (
  .A({ S11620 }),
  .B1({ S17584 }),
  .B2({ S17595 }),
  .ZN({ S17606 })
);
AOI22_X1 #() 
AOI22_X1_347_ (
  .A1({ S17554 }),
  .A2({ S11620 }),
  .B1({ S17574 }),
  .B2({ S17606 }),
  .ZN({ S17617 })
);
OAI21_X1 #() 
OAI21_X1_1571_ (
  .A({ S11609 }),
  .B1({ S17617 }),
  .B2({ S11631 }),
  .ZN({ S17628 })
);
INV_X1 #() 
INV_X1_983_ (
  .A({ S13516 }),
  .ZN({ S17639 })
);
NAND3_X1 #() 
NAND3_X1_3252_ (
  .A1({ S17381 }),
  .A2({ S25956[4] }),
  .A3({ S14997 }),
  .ZN({ S17650 })
);
OAI211_X1 #() 
OAI211_X1_1055_ (
  .A({ S17650 }),
  .B({ S11631 }),
  .C1({ S17639 }),
  .C2({ S17532 }),
  .ZN({ S17661 })
);
NAND3_X1 #() 
NAND3_X1_3253_ (
  .A1({ S12097 }),
  .A2({ S25956[3] }),
  .A3({ S25956[0] }),
  .ZN({ S17672 })
);
AND3_X1 #() 
AND3_X1_125_ (
  .A1({ S15506 }),
  .A2({ S25956[4] }),
  .A3({ S17672 }),
  .ZN({ S17683 })
);
NAND2_X1 #() 
NAND2_X1_2987_ (
  .A1({ S58 }),
  .A2({ S25956[3] }),
  .ZN({ S17694 })
);
OAI211_X1 #() 
OAI211_X1_1056_ (
  .A({ S17694 }),
  .B({ S13000 }),
  .C1({ S11821 }),
  .C2({ S13872 }),
  .ZN({ S17705 })
);
OAI21_X1 #() 
OAI21_X1_1572_ (
  .A({ S25956[5] }),
  .B1({ S17705 }),
  .B2({ S25956[4] }),
  .ZN({ S17716 })
);
OAI211_X1 #() 
OAI211_X1_1057_ (
  .A({ S17661 }),
  .B({ S11620 }),
  .C1({ S17716 }),
  .C2({ S17683 }),
  .ZN({ S17726 })
);
NAND3_X1 #() 
NAND3_X1_3254_ (
  .A1({ S12520 }),
  .A2({ S13987 }),
  .A3({ S25956[3] }),
  .ZN({ S17737 })
);
NOR2_X1 #() 
NOR2_X1_750_ (
  .A1({ S12053 }),
  .A2({ S25956[4] }),
  .ZN({ S17748 })
);
NAND2_X1 #() 
NAND2_X1_2988_ (
  .A1({ S17737 }),
  .A2({ S17748 }),
  .ZN({ S17759 })
);
NAND4_X1 #() 
NAND4_X1_352_ (
  .A1({ S11683 }),
  .A2({ S25956[4] }),
  .A3({ S16204 }),
  .A4({ S16226 }),
  .ZN({ S17770 })
);
NAND3_X1 #() 
NAND3_X1_3255_ (
  .A1({ S17759 }),
  .A2({ S17770 }),
  .A3({ S25956[5] }),
  .ZN({ S17781 })
);
NAND3_X1 #() 
NAND3_X1_3256_ (
  .A1({ S12520 }),
  .A2({ S25956[3] }),
  .A3({ S12501 }),
  .ZN({ S17792 })
);
NAND2_X1 #() 
NAND2_X1_2989_ (
  .A1({ S17792 }),
  .A2({ S13817 }),
  .ZN({ S17803 })
);
AOI21_X1 #() 
AOI21_X1_1665_ (
  .A({ S25956[4] }),
  .B1({ S12442 }),
  .B2({ S11664 }),
  .ZN({ S17814 })
);
AOI21_X1 #() 
AOI21_X1_1666_ (
  .A({ S25956[5] }),
  .B1({ S12075 }),
  .B2({ S17814 }),
  .ZN({ S17824 })
);
AOI21_X1 #() 
AOI21_X1_1667_ (
  .A({ S11620 }),
  .B1({ S17803 }),
  .B2({ S17824 }),
  .ZN({ S17835 })
);
NAND2_X1 #() 
NAND2_X1_2990_ (
  .A1({ S17835 }),
  .A2({ S17781 }),
  .ZN({ S17846 })
);
NAND3_X1 #() 
NAND3_X1_3257_ (
  .A1({ S17846 }),
  .A2({ S17726 }),
  .A3({ S25956[7] }),
  .ZN({ S17857 })
);
OAI211_X1 #() 
OAI211_X1_1058_ (
  .A({ S17857 }),
  .B({ S17370 }),
  .C1({ S17628 }),
  .C2({ S17500 }),
  .ZN({ S17868 })
);
OAI21_X1 #() 
OAI21_X1_1573_ (
  .A({ S17857 }),
  .B1({ S17628 }),
  .B2({ S17500 }),
  .ZN({ S17879 })
);
NAND2_X1 #() 
NAND2_X1_2991_ (
  .A1({ S17879 }),
  .A2({ S25956[106] }),
  .ZN({ S17889 })
);
NAND3_X1 #() 
NAND3_X1_3258_ (
  .A1({ S17889 }),
  .A2({ S17359 }),
  .A3({ S17868 }),
  .ZN({ S17900 })
);
NAND2_X1 #() 
NAND2_X1_2992_ (
  .A1({ S17879 }),
  .A2({ S17370 }),
  .ZN({ S17911 })
);
OAI211_X1 #() 
OAI211_X1_1059_ (
  .A({ S17857 }),
  .B({ S25956[106] }),
  .C1({ S17628 }),
  .C2({ S17500 }),
  .ZN({ S17922 })
);
NAND3_X1 #() 
NAND3_X1_3259_ (
  .A1({ S17911 }),
  .A2({ S25956[74] }),
  .A3({ S17922 }),
  .ZN({ S17933 })
);
NAND3_X1 #() 
NAND3_X1_3260_ (
  .A1({ S17900 }),
  .A2({ S17933 }),
  .A3({ S17348 }),
  .ZN({ S17944 })
);
NAND3_X1 #() 
NAND3_X1_3261_ (
  .A1({ S17911 }),
  .A2({ S17359 }),
  .A3({ S17922 }),
  .ZN({ S17954 })
);
NAND3_X1 #() 
NAND3_X1_3262_ (
  .A1({ S17889 }),
  .A2({ S25956[74] }),
  .A3({ S17868 }),
  .ZN({ S17965 })
);
NAND3_X1 #() 
NAND3_X1_3263_ (
  .A1({ S17954 }),
  .A2({ S17965 }),
  .A3({ S25956[42] }),
  .ZN({ S17976 })
);
NAND3_X1 #() 
NAND3_X1_3264_ (
  .A1({ S17944 }),
  .A2({ S17976 }),
  .A3({ S25956[10] }),
  .ZN({ S17987 })
);
NAND3_X1 #() 
NAND3_X1_3265_ (
  .A1({ S17954 }),
  .A2({ S17965 }),
  .A3({ S17348 }),
  .ZN({ S17998 })
);
NAND3_X1 #() 
NAND3_X1_3266_ (
  .A1({ S17900 }),
  .A2({ S17933 }),
  .A3({ S25956[42] }),
  .ZN({ S18008 })
);
NAND3_X1 #() 
NAND3_X1_3267_ (
  .A1({ S17998 }),
  .A2({ S18008 }),
  .A3({ S5730 }),
  .ZN({ S18019 })
);
NAND2_X1 #() 
NAND2_X1_2993_ (
  .A1({ S17987 }),
  .A2({ S18019 }),
  .ZN({ S25957[1162] })
);
NOR2_X1 #() 
NOR2_X1_751_ (
  .A1({ S25956[25] }),
  .A2({ S25956[24] }),
  .ZN({ S18040 })
);
INV_X1 #() 
INV_X1_984_ (
  .A({ S18040 }),
  .ZN({ S66 })
);
NAND2_X1 #() 
NAND2_X1_2994_ (
  .A1({ S25956[25] }),
  .A2({ S25956[24] }),
  .ZN({ S18060 })
);
INV_X1 #() 
INV_X1_985_ (
  .A({ S18060 }),
  .ZN({ S67 })
);
INV_X1 #() 
INV_X1_986_ (
  .A({ S25956[31] }),
  .ZN({ S18081 })
);
INV_X1 #() 
INV_X1_987_ (
  .A({ S25956[30] }),
  .ZN({ S18092 })
);
INV_X1 #() 
INV_X1_988_ (
  .A({ S25956[29] }),
  .ZN({ S18103 })
);
INV_X1 #() 
INV_X1_989_ (
  .A({ S25956[28] }),
  .ZN({ S18113 })
);
INV_X1 #() 
INV_X1_990_ (
  .A({ S25956[27] }),
  .ZN({ S18124 })
);
NOR2_X1 #() 
NOR2_X1_752_ (
  .A1({ S18060 }),
  .A2({ S18124 }),
  .ZN({ S18135 })
);
INV_X1 #() 
INV_X1_991_ (
  .A({ S18135 }),
  .ZN({ S18146 })
);
NAND2_X1 #() 
NAND2_X1_2995_ (
  .A1({ S25956[26] }),
  .A2({ S25956[25] }),
  .ZN({ S18156 })
);
NOR2_X1 #() 
NOR2_X1_753_ (
  .A1({ S18124 }),
  .A2({ S25956[24] }),
  .ZN({ S18165 })
);
NAND2_X1 #() 
NAND2_X1_2996_ (
  .A1({ S18165 }),
  .A2({ S18156 }),
  .ZN({ S18176 })
);
NAND2_X1 #() 
NAND2_X1_2997_ (
  .A1({ S18040 }),
  .A2({ S25956[26] }),
  .ZN({ S18187 })
);
INV_X1 #() 
INV_X1_992_ (
  .A({ S25956[26] }),
  .ZN({ S18198 })
);
NAND2_X1 #() 
NAND2_X1_2998_ (
  .A1({ S67 }),
  .A2({ S18198 }),
  .ZN({ S18209 })
);
NAND3_X1 #() 
NAND3_X1_3268_ (
  .A1({ S18209 }),
  .A2({ S18124 }),
  .A3({ S18187 }),
  .ZN({ S18220 })
);
NAND3_X1 #() 
NAND3_X1_3269_ (
  .A1({ S18220 }),
  .A2({ S18146 }),
  .A3({ S18176 }),
  .ZN({ S18231 })
);
INV_X1 #() 
INV_X1_993_ (
  .A({ S25956[24] }),
  .ZN({ S18242 })
);
NAND2_X1 #() 
NAND2_X1_2999_ (
  .A1({ S18198 }),
  .A2({ S18242 }),
  .ZN({ S18253 })
);
NAND2_X1 #() 
NAND2_X1_3000_ (
  .A1({ S18198 }),
  .A2({ S25956[25] }),
  .ZN({ S18264 })
);
NAND2_X1 #() 
NAND2_X1_3001_ (
  .A1({ S18253 }),
  .A2({ S18264 }),
  .ZN({ S18275 })
);
NAND2_X1 #() 
NAND2_X1_3002_ (
  .A1({ S18275 }),
  .A2({ S25956[27] }),
  .ZN({ S18285 })
);
INV_X1 #() 
INV_X1_994_ (
  .A({ S18285 }),
  .ZN({ S18296 })
);
NOR2_X1 #() 
NOR2_X1_754_ (
  .A1({ S18296 }),
  .A2({ S18113 }),
  .ZN({ S18307 })
);
NAND2_X1 #() 
NAND2_X1_3003_ (
  .A1({ S25956[26] }),
  .A2({ S25956[24] }),
  .ZN({ S18318 })
);
NOR2_X1 #() 
NOR2_X1_755_ (
  .A1({ S18318 }),
  .A2({ S18124 }),
  .ZN({ S18329 })
);
NAND2_X1 #() 
NAND2_X1_3004_ (
  .A1({ S18253 }),
  .A2({ S25956[25] }),
  .ZN({ S18340 })
);
INV_X1 #() 
INV_X1_995_ (
  .A({ S18340 }),
  .ZN({ S18351 })
);
AOI21_X1 #() 
AOI21_X1_1668_ (
  .A({ S18329 }),
  .B1({ S18351 }),
  .B2({ S18124 }),
  .ZN({ S18362 })
);
AOI22_X1 #() 
AOI22_X1_348_ (
  .A1({ S18307 }),
  .A2({ S18362 }),
  .B1({ S18231 }),
  .B2({ S18113 }),
  .ZN({ S18372 })
);
INV_X1 #() 
INV_X1_996_ (
  .A({ S25956[25] }),
  .ZN({ S18383 })
);
NAND2_X1 #() 
NAND2_X1_3005_ (
  .A1({ S18383 }),
  .A2({ S25956[26] }),
  .ZN({ S18394 })
);
NAND3_X1 #() 
NAND3_X1_3270_ (
  .A1({ S18394 }),
  .A2({ S25956[27] }),
  .A3({ S18060 }),
  .ZN({ S18405 })
);
NAND2_X1 #() 
NAND2_X1_3006_ (
  .A1({ S18242 }),
  .A2({ S25956[25] }),
  .ZN({ S18416 })
);
NAND2_X1 #() 
NAND2_X1_3007_ (
  .A1({ S18416 }),
  .A2({ S18124 }),
  .ZN({ S18427 })
);
AOI21_X1 #() 
AOI21_X1_1669_ (
  .A({ S18113 }),
  .B1({ S18405 }),
  .B2({ S18427 }),
  .ZN({ S18438 })
);
NAND2_X1 #() 
NAND2_X1_3008_ (
  .A1({ S18156 }),
  .A2({ S18318 }),
  .ZN({ S18448 })
);
INV_X1 #() 
INV_X1_997_ (
  .A({ S18448 }),
  .ZN({ S18459 })
);
NOR2_X1 #() 
NOR2_X1_756_ (
  .A1({ S25956[26] }),
  .A2({ S25956[25] }),
  .ZN({ S18470 })
);
INV_X1 #() 
INV_X1_998_ (
  .A({ S18470 }),
  .ZN({ S18481 })
);
NAND2_X1 #() 
NAND2_X1_3009_ (
  .A1({ S18124 }),
  .A2({ S25956[24] }),
  .ZN({ S18492 })
);
INV_X1 #() 
INV_X1_999_ (
  .A({ S18492 }),
  .ZN({ S18502 })
);
OAI211_X1 #() 
OAI211_X1_1060_ (
  .A({ S18459 }),
  .B({ S18113 }),
  .C1({ S18481 }),
  .C2({ S18502 }),
  .ZN({ S18513 })
);
NAND2_X1 #() 
NAND2_X1_3010_ (
  .A1({ S18513 }),
  .A2({ S18103 }),
  .ZN({ S18524 })
);
OAI22_X1 #() 
OAI22_X1_79_ (
  .A1({ S18372 }),
  .A2({ S18103 }),
  .B1({ S18438 }),
  .B2({ S18524 }),
  .ZN({ S18535 })
);
NAND2_X1 #() 
NAND2_X1_3011_ (
  .A1({ S18383 }),
  .A2({ S25956[27] }),
  .ZN({ S18545 })
);
NOR2_X1 #() 
NOR2_X1_757_ (
  .A1({ S18545 }),
  .A2({ S25956[26] }),
  .ZN({ S18556 })
);
NAND2_X1 #() 
NAND2_X1_3012_ (
  .A1({ S18383 }),
  .A2({ S25956[24] }),
  .ZN({ S18567 })
);
NAND2_X1 #() 
NAND2_X1_3013_ (
  .A1({ S18567 }),
  .A2({ S25956[26] }),
  .ZN({ S18578 })
);
INV_X1 #() 
INV_X1_1000_ (
  .A({ S18578 }),
  .ZN({ S18588 })
);
NAND2_X1 #() 
NAND2_X1_3014_ (
  .A1({ S18060 }),
  .A2({ S18198 }),
  .ZN({ S18599 })
);
NOR2_X1 #() 
NOR2_X1_758_ (
  .A1({ S18599 }),
  .A2({ S18040 }),
  .ZN({ S18610 })
);
NOR2_X1 #() 
NOR2_X1_759_ (
  .A1({ S18588 }),
  .A2({ S18610 }),
  .ZN({ S18621 })
);
AOI21_X1 #() 
AOI21_X1_1670_ (
  .A({ S18556 }),
  .B1({ S18621 }),
  .B2({ S18124 }),
  .ZN({ S18632 })
);
NAND2_X1 #() 
NAND2_X1_3015_ (
  .A1({ S18296 }),
  .A2({ S18416 }),
  .ZN({ S18643 })
);
NAND2_X1 #() 
NAND2_X1_3016_ (
  .A1({ S18643 }),
  .A2({ S25956[28] }),
  .ZN({ S18654 })
);
INV_X1 #() 
INV_X1_1001_ (
  .A({ S18156 }),
  .ZN({ S18664 })
);
NOR2_X1 #() 
NOR2_X1_760_ (
  .A1({ S18242 }),
  .A2({ S25956[26] }),
  .ZN({ S18675 })
);
INV_X1 #() 
INV_X1_1002_ (
  .A({ S18675 }),
  .ZN({ S18686 })
);
NAND2_X1 #() 
NAND2_X1_3017_ (
  .A1({ S18686 }),
  .A2({ S18124 }),
  .ZN({ S18697 })
);
NAND2_X1 #() 
NAND2_X1_3018_ (
  .A1({ S18060 }),
  .A2({ S25956[26] }),
  .ZN({ S18707 })
);
NOR2_X1 #() 
NOR2_X1_761_ (
  .A1({ S18707 }),
  .A2({ S18040 }),
  .ZN({ S18716 })
);
NAND2_X1 #() 
NAND2_X1_3019_ (
  .A1({ S18716 }),
  .A2({ S25956[27] }),
  .ZN({ S18725 })
);
OAI21_X1 #() 
OAI21_X1_1574_ (
  .A({ S18725 }),
  .B1({ S18664 }),
  .B2({ S18697 }),
  .ZN({ S18735 })
);
OAI22_X1 #() 
OAI22_X1_80_ (
  .A1({ S18654 }),
  .A2({ S18735 }),
  .B1({ S18632 }),
  .B2({ S25956[28] }),
  .ZN({ S18744 })
);
AOI21_X1 #() 
AOI21_X1_1671_ (
  .A({ S25956[28] }),
  .B1({ S18253 }),
  .B2({ S18124 }),
  .ZN({ S18753 })
);
OAI21_X1 #() 
OAI21_X1_1575_ (
  .A({ S18753 }),
  .B1({ S18383 }),
  .B2({ S18165 }),
  .ZN({ S18762 })
);
INV_X1 #() 
INV_X1_1003_ (
  .A({ S18318 }),
  .ZN({ S18769 })
);
NAND2_X1 #() 
NAND2_X1_3020_ (
  .A1({ S18124 }),
  .A2({ S25956[25] }),
  .ZN({ S18780 })
);
INV_X1 #() 
INV_X1_1004_ (
  .A({ S18329 }),
  .ZN({ S18790 })
);
NAND2_X1 #() 
NAND2_X1_3021_ (
  .A1({ S18790 }),
  .A2({ S18545 }),
  .ZN({ S18798 })
);
NOR2_X1 #() 
NOR2_X1_762_ (
  .A1({ S18798 }),
  .A2({ S18113 }),
  .ZN({ S18807 })
);
OAI21_X1 #() 
OAI21_X1_1576_ (
  .A({ S18807 }),
  .B1({ S18769 }),
  .B2({ S18780 }),
  .ZN({ S18814 })
);
NAND3_X1 #() 
NAND3_X1_3271_ (
  .A1({ S18814 }),
  .A2({ S25956[29] }),
  .A3({ S18762 }),
  .ZN({ S18823 })
);
OAI21_X1 #() 
OAI21_X1_1577_ (
  .A({ S18823 }),
  .B1({ S18744 }),
  .B2({ S25956[29] }),
  .ZN({ S18834 })
);
NAND2_X1 #() 
NAND2_X1_3022_ (
  .A1({ S18834 }),
  .A2({ S18092 }),
  .ZN({ S18842 })
);
OAI21_X1 #() 
OAI21_X1_1578_ (
  .A({ S18842 }),
  .B1({ S18092 }),
  .B2({ S18535 }),
  .ZN({ S18852 })
);
NOR2_X1 #() 
NOR2_X1_763_ (
  .A1({ S18383 }),
  .A2({ S25956[26] }),
  .ZN({ S18863 })
);
NAND2_X1 #() 
NAND2_X1_3023_ (
  .A1({ S18318 }),
  .A2({ S25956[27] }),
  .ZN({ S18874 })
);
NOR2_X1 #() 
NOR2_X1_764_ (
  .A1({ S18874 }),
  .A2({ S18863 }),
  .ZN({ S18883 })
);
INV_X1 #() 
INV_X1_1005_ (
  .A({ S18707 }),
  .ZN({ S18892 })
);
NAND2_X1 #() 
NAND2_X1_3024_ (
  .A1({ S18892 }),
  .A2({ S18124 }),
  .ZN({ S18900 })
);
NOR2_X1 #() 
NOR2_X1_765_ (
  .A1({ S25956[27] }),
  .A2({ S25956[26] }),
  .ZN({ S18909 })
);
NAND2_X1 #() 
NAND2_X1_3025_ (
  .A1({ S18567 }),
  .A2({ S18909 }),
  .ZN({ S18917 })
);
NAND3_X1 #() 
NAND3_X1_3272_ (
  .A1({ S18900 }),
  .A2({ S18113 }),
  .A3({ S18917 }),
  .ZN({ S18927 })
);
NAND2_X1 #() 
NAND2_X1_3026_ (
  .A1({ S18275 }),
  .A2({ S18416 }),
  .ZN({ S18935 })
);
AOI21_X1 #() 
AOI21_X1_1672_ (
  .A({ S18124 }),
  .B1({ S18935 }),
  .B2({ S18707 }),
  .ZN({ S18945 })
);
NOR2_X1 #() 
NOR2_X1_766_ (
  .A1({ S18492 }),
  .A2({ S18156 }),
  .ZN({ S18953 })
);
NAND2_X1 #() 
NAND2_X1_3027_ (
  .A1({ S18156 }),
  .A2({ S18124 }),
  .ZN({ S18962 })
);
NOR2_X1 #() 
NOR2_X1_767_ (
  .A1({ S18962 }),
  .A2({ S25956[24] }),
  .ZN({ S18970 })
);
NOR2_X1 #() 
NOR2_X1_768_ (
  .A1({ S18970 }),
  .A2({ S18953 }),
  .ZN({ S18978 })
);
NAND2_X1 #() 
NAND2_X1_3028_ (
  .A1({ S18978 }),
  .A2({ S25956[28] }),
  .ZN({ S18986 })
);
OAI22_X1 #() 
OAI22_X1_81_ (
  .A1({ S18986 }),
  .A2({ S18945 }),
  .B1({ S18927 }),
  .B2({ S18883 }),
  .ZN({ S18995 })
);
NAND3_X1 #() 
NAND3_X1_3273_ (
  .A1({ S18209 }),
  .A2({ S25956[27] }),
  .A3({ S18187 }),
  .ZN({ S19004 })
);
NAND2_X1 #() 
NAND2_X1_3029_ (
  .A1({ S18962 }),
  .A2({ S18492 }),
  .ZN({ S19012 })
);
AOI21_X1 #() 
AOI21_X1_1673_ (
  .A({ S18113 }),
  .B1({ S19012 }),
  .B2({ S18253 }),
  .ZN({ S19021 })
);
NAND2_X1 #() 
NAND2_X1_3030_ (
  .A1({ S18567 }),
  .A2({ S18198 }),
  .ZN({ S19030 })
);
AOI21_X1 #() 
AOI21_X1_1674_ (
  .A({ S18124 }),
  .B1({ S19030 }),
  .B2({ S18394 }),
  .ZN({ S19038 })
);
INV_X1 #() 
INV_X1_1006_ (
  .A({ S19038 }),
  .ZN({ S19048 })
);
AOI21_X1 #() 
AOI21_X1_1675_ (
  .A({ S25956[28] }),
  .B1({ S19048 }),
  .B2({ S18900 }),
  .ZN({ S19056 })
);
AOI21_X1 #() 
AOI21_X1_1676_ (
  .A({ S19056 }),
  .B1({ S19021 }),
  .B2({ S19004 }),
  .ZN({ S19065 })
);
MUX2_X1 #() 
MUX2_X1_12_ (
  .A({ S18995 }),
  .B({ S19065 }),
  .S({ S25956[29] }),
  .Z({ S19073 })
);
NOR2_X1 #() 
NOR2_X1_769_ (
  .A1({ S18156 }),
  .A2({ S25956[24] }),
  .ZN({ S19082 })
);
NAND2_X1 #() 
NAND2_X1_3031_ (
  .A1({ S66 }),
  .A2({ S18060 }),
  .ZN({ S19091 })
);
NAND2_X1 #() 
NAND2_X1_3032_ (
  .A1({ S19091 }),
  .A2({ S25956[26] }),
  .ZN({ S19098 })
);
NAND2_X1 #() 
NAND2_X1_3033_ (
  .A1({ S19098 }),
  .A2({ S18599 }),
  .ZN({ S19107 })
);
NAND2_X1 #() 
NAND2_X1_3034_ (
  .A1({ S19107 }),
  .A2({ S18124 }),
  .ZN({ S19108 })
);
OAI211_X1 #() 
OAI211_X1_1061_ (
  .A({ S19108 }),
  .B({ S25956[28] }),
  .C1({ S19082 }),
  .C2({ S18124 }),
  .ZN({ S19109 })
);
INV_X1 #() 
INV_X1_1007_ (
  .A({ S19098 }),
  .ZN({ S19110 })
);
NAND2_X1 #() 
NAND2_X1_3035_ (
  .A1({ S19110 }),
  .A2({ S18124 }),
  .ZN({ S19111 })
);
OAI211_X1 #() 
OAI211_X1_1062_ (
  .A({ S19111 }),
  .B({ S18113 }),
  .C1({ S18707 }),
  .C2({ S18124 }),
  .ZN({ S19112 })
);
NAND3_X1 #() 
NAND3_X1_3274_ (
  .A1({ S19109 }),
  .A2({ S18103 }),
  .A3({ S19112 }),
  .ZN({ S19113 })
);
INV_X1 #() 
INV_X1_1008_ (
  .A({ S18962 }),
  .ZN({ S19114 })
);
AOI21_X1 #() 
AOI21_X1_1677_ (
  .A({ S18124 }),
  .B1({ S66 }),
  .B2({ S18156 }),
  .ZN({ S19115 })
);
AOI21_X1 #() 
AOI21_X1_1678_ (
  .A({ S19115 }),
  .B1({ S19114 }),
  .B2({ S18599 }),
  .ZN({ S19116 })
);
INV_X1 #() 
INV_X1_1009_ (
  .A({ S18874 }),
  .ZN({ S19117 })
);
NAND2_X1 #() 
NAND2_X1_3036_ (
  .A1({ S19117 }),
  .A2({ S18481 }),
  .ZN({ S19118 })
);
NAND3_X1 #() 
NAND3_X1_3275_ (
  .A1({ S19118 }),
  .A2({ S25956[28] }),
  .A3({ S18492 }),
  .ZN({ S19119 })
);
OAI211_X1 #() 
OAI211_X1_1063_ (
  .A({ S19119 }),
  .B({ S25956[29] }),
  .C1({ S19116 }),
  .C2({ S25956[28] }),
  .ZN({ S19120 })
);
NAND3_X1 #() 
NAND3_X1_3276_ (
  .A1({ S19113 }),
  .A2({ S18092 }),
  .A3({ S19120 }),
  .ZN({ S19121 })
);
OAI211_X1 #() 
OAI211_X1_1064_ (
  .A({ S19121 }),
  .B({ S18081 }),
  .C1({ S19073 }),
  .C2({ S18092 }),
  .ZN({ S19122 })
);
OAI21_X1 #() 
OAI21_X1_1579_ (
  .A({ S19122 }),
  .B1({ S18852 }),
  .B2({ S18081 }),
  .ZN({ S19123 })
);
XNOR2_X1 #() 
XNOR2_X1_159_ (
  .A({ S19123 }),
  .B({ S25956[103] }),
  .ZN({ S19124 })
);
XOR2_X1 #() 
XOR2_X1_68_ (
  .A({ S19124 }),
  .B({ S25956[71] }),
  .Z({ S19125 })
);
XNOR2_X1 #() 
XNOR2_X1_160_ (
  .A({ S19125 }),
  .B({ S25956[39] }),
  .ZN({ S25957[1191] })
);
XNOR2_X1 #() 
XNOR2_X1_161_ (
  .A({ S25957[1191] }),
  .B({ S25956[7] }),
  .ZN({ S19126 })
);
INV_X1 #() 
INV_X1_1010_ (
  .A({ S19126 }),
  .ZN({ S25957[1159] })
);
INV_X1 #() 
INV_X1_1011_ (
  .A({ S25956[70] }),
  .ZN({ S19127 })
);
NOR2_X1 #() 
NOR2_X1_770_ (
  .A1({ S18664 }),
  .A2({ S25956[24] }),
  .ZN({ S19128 })
);
OAI21_X1 #() 
OAI21_X1_1580_ (
  .A({ S18124 }),
  .B1({ S18610 }),
  .B2({ S18769 }),
  .ZN({ S19129 })
);
OAI21_X1 #() 
OAI21_X1_1581_ (
  .A({ S19129 }),
  .B1({ S19128 }),
  .B2({ S18874 }),
  .ZN({ S19130 })
);
NAND2_X1 #() 
NAND2_X1_3037_ (
  .A1({ S19130 }),
  .A2({ S18113 }),
  .ZN({ S19131 })
);
NAND2_X1 #() 
NAND2_X1_3038_ (
  .A1({ S18917 }),
  .A2({ S25956[28] }),
  .ZN({ S19132 })
);
OAI211_X1 #() 
OAI211_X1_1065_ (
  .A({ S19131 }),
  .B({ S18103 }),
  .C1({ S18798 }),
  .C2({ S19132 }),
  .ZN({ S19133 })
);
NAND2_X1 #() 
NAND2_X1_3039_ (
  .A1({ S18416 }),
  .A2({ S18198 }),
  .ZN({ S19134 })
);
OAI21_X1 #() 
OAI21_X1_1582_ (
  .A({ S18124 }),
  .B1({ S18707 }),
  .B2({ S18040 }),
  .ZN({ S19135 })
);
INV_X1 #() 
INV_X1_1012_ (
  .A({ S19135 }),
  .ZN({ S19136 })
);
NAND2_X1 #() 
NAND2_X1_3040_ (
  .A1({ S25956[27] }),
  .A2({ S25956[26] }),
  .ZN({ S19137 })
);
INV_X1 #() 
INV_X1_1013_ (
  .A({ S19137 }),
  .ZN({ S19138 })
);
NAND2_X1 #() 
NAND2_X1_3041_ (
  .A1({ S19138 }),
  .A2({ S25956[25] }),
  .ZN({ S19139 })
);
NAND2_X1 #() 
NAND2_X1_3042_ (
  .A1({ S19139 }),
  .A2({ S25956[28] }),
  .ZN({ S19140 })
);
AOI21_X1 #() 
AOI21_X1_1679_ (
  .A({ S19140 }),
  .B1({ S19136 }),
  .B2({ S19134 }),
  .ZN({ S19141 })
);
NAND2_X1 #() 
NAND2_X1_3043_ (
  .A1({ S18394 }),
  .A2({ S25956[27] }),
  .ZN({ S19142 })
);
NOR2_X1 #() 
NOR2_X1_771_ (
  .A1({ S18383 }),
  .A2({ S25956[24] }),
  .ZN({ S19143 })
);
NAND2_X1 #() 
NAND2_X1_3044_ (
  .A1({ S19143 }),
  .A2({ S18198 }),
  .ZN({ S19144 })
);
INV_X1 #() 
INV_X1_1014_ (
  .A({ S19144 }),
  .ZN({ S19145 })
);
NOR2_X1 #() 
NOR2_X1_772_ (
  .A1({ S18318 }),
  .A2({ S18383 }),
  .ZN({ S19146 })
);
NOR2_X1 #() 
NOR2_X1_773_ (
  .A1({ S19146 }),
  .A2({ S18040 }),
  .ZN({ S19147 })
);
OAI22_X1 #() 
OAI22_X1_82_ (
  .A1({ S19145 }),
  .A2({ S19142 }),
  .B1({ S19147 }),
  .B2({ S25956[27] }),
  .ZN({ S19148 })
);
AOI21_X1 #() 
AOI21_X1_1680_ (
  .A({ S19141 }),
  .B1({ S18113 }),
  .B2({ S19148 }),
  .ZN({ S19149 })
);
OAI211_X1 #() 
OAI211_X1_1066_ (
  .A({ S19133 }),
  .B({ S18092 }),
  .C1({ S18103 }),
  .C2({ S19149 }),
  .ZN({ S19150 })
);
NAND2_X1 #() 
NAND2_X1_3045_ (
  .A1({ S18242 }),
  .A2({ S25956[26] }),
  .ZN({ S19151 })
);
NOR2_X1 #() 
NOR2_X1_774_ (
  .A1({ S18675 }),
  .A2({ S18545 }),
  .ZN({ S19152 })
);
NAND2_X1 #() 
NAND2_X1_3046_ (
  .A1({ S19152 }),
  .A2({ S19151 }),
  .ZN({ S19153 })
);
OAI211_X1 #() 
OAI211_X1_1067_ (
  .A({ S19153 }),
  .B({ S25956[28] }),
  .C1({ S18459 }),
  .C2({ S25956[27] }),
  .ZN({ S19154 })
);
NAND2_X1 #() 
NAND2_X1_3047_ (
  .A1({ S18405 }),
  .A2({ S18780 }),
  .ZN({ S19155 })
);
AOI21_X1 #() 
AOI21_X1_1681_ (
  .A({ S18103 }),
  .B1({ S19155 }),
  .B2({ S18113 }),
  .ZN({ S19156 })
);
INV_X1 #() 
INV_X1_1015_ (
  .A({ S18599 }),
  .ZN({ S19157 })
);
NAND2_X1 #() 
NAND2_X1_3048_ (
  .A1({ S18187 }),
  .A2({ S25956[27] }),
  .ZN({ S19158 })
);
NOR2_X1 #() 
NOR2_X1_775_ (
  .A1({ S19158 }),
  .A2({ S19157 }),
  .ZN({ S19159 })
);
OAI21_X1 #() 
OAI21_X1_1583_ (
  .A({ S25956[27] }),
  .B1({ S18588 }),
  .B2({ S18675 }),
  .ZN({ S19160 })
);
NAND3_X1 #() 
NAND3_X1_3277_ (
  .A1({ S19160 }),
  .A2({ S19129 }),
  .A3({ S25956[28] }),
  .ZN({ S19161 })
);
OAI21_X1 #() 
OAI21_X1_1584_ (
  .A({ S19161 }),
  .B1({ S18927 }),
  .B2({ S19159 }),
  .ZN({ S19162 })
);
AOI22_X1 #() 
AOI22_X1_349_ (
  .A1({ S19162 }),
  .A2({ S18103 }),
  .B1({ S19154 }),
  .B2({ S19156 }),
  .ZN({ S19163 })
);
NAND2_X1 #() 
NAND2_X1_3049_ (
  .A1({ S19163 }),
  .A2({ S25956[30] }),
  .ZN({ S19164 })
);
NAND3_X1 #() 
NAND3_X1_3278_ (
  .A1({ S19150 }),
  .A2({ S25956[31] }),
  .A3({ S19164 }),
  .ZN({ S19165 })
);
NOR2_X1 #() 
NOR2_X1_776_ (
  .A1({ S18892 }),
  .A2({ S18675 }),
  .ZN({ S19166 })
);
NOR2_X1 #() 
NOR2_X1_777_ (
  .A1({ S19166 }),
  .A2({ S25956[27] }),
  .ZN({ S19167 })
);
AOI211_X1 #() 
AOI211_X1_45_ (
  .A({ S18113 }),
  .B({ S19167 }),
  .C1({ S18416 }),
  .C2({ S19117 }),
  .ZN({ S19168 })
);
NOR2_X1 #() 
NOR2_X1_778_ (
  .A1({ S18470 }),
  .A2({ S25956[24] }),
  .ZN({ S19169 })
);
NAND2_X1 #() 
NAND2_X1_3050_ (
  .A1({ S19169 }),
  .A2({ S18124 }),
  .ZN({ S19170 })
);
NAND2_X1 #() 
NAND2_X1_3051_ (
  .A1({ S18863 }),
  .A2({ S25956[27] }),
  .ZN({ S19171 })
);
NAND3_X1 #() 
NAND3_X1_3279_ (
  .A1({ S19170 }),
  .A2({ S25956[28] }),
  .A3({ S19171 }),
  .ZN({ S19172 })
);
NAND3_X1 #() 
NAND3_X1_3280_ (
  .A1({ S19160 }),
  .A2({ S19135 }),
  .A3({ S18113 }),
  .ZN({ S19173 })
);
NAND3_X1 #() 
NAND3_X1_3281_ (
  .A1({ S19173 }),
  .A2({ S18103 }),
  .A3({ S19172 }),
  .ZN({ S19174 })
);
NAND2_X1 #() 
NAND2_X1_3052_ (
  .A1({ S18416 }),
  .A2({ S18156 }),
  .ZN({ S19175 })
);
INV_X1 #() 
INV_X1_1016_ (
  .A({ S19175 }),
  .ZN({ S19176 })
);
AOI22_X1 #() 
AOI22_X1_350_ (
  .A1({ S19176 }),
  .A2({ S18124 }),
  .B1({ S19117 }),
  .B2({ S18416 }),
  .ZN({ S19177 })
);
OAI21_X1 #() 
OAI21_X1_1585_ (
  .A({ S25956[29] }),
  .B1({ S19177 }),
  .B2({ S25956[28] }),
  .ZN({ S19178 })
);
OAI211_X1 #() 
OAI211_X1_1068_ (
  .A({ S19174 }),
  .B({ S25956[30] }),
  .C1({ S19168 }),
  .C2({ S19178 }),
  .ZN({ S19179 })
);
NAND3_X1 #() 
NAND3_X1_3282_ (
  .A1({ S19151 }),
  .A2({ S25956[27] }),
  .A3({ S18060 }),
  .ZN({ S19180 })
);
NAND2_X1 #() 
NAND2_X1_3053_ (
  .A1({ S19143 }),
  .A2({ S25956[27] }),
  .ZN({ S19181 })
);
NAND4_X1 #() 
NAND4_X1_353_ (
  .A1({ S18697 }),
  .A2({ S25956[28] }),
  .A3({ S19180 }),
  .A4({ S19181 }),
  .ZN({ S19182 })
);
AOI21_X1 #() 
AOI21_X1_1682_ (
  .A({ S18962 }),
  .B1({ S18675 }),
  .B2({ S18383 }),
  .ZN({ S19183 })
);
OAI21_X1 #() 
OAI21_X1_1586_ (
  .A({ S18113 }),
  .B1({ S19142 }),
  .B2({ S18863 }),
  .ZN({ S19184 })
);
OAI21_X1 #() 
OAI21_X1_1587_ (
  .A({ S19182 }),
  .B1({ S19183 }),
  .B2({ S19184 }),
  .ZN({ S19185 })
);
AOI211_X1 #() 
AOI211_X1_46_ (
  .A({ S18113 }),
  .B({ S19038 }),
  .C1({ S18470 }),
  .C2({ S18502 }),
  .ZN({ S19186 })
);
INV_X1 #() 
INV_X1_1017_ (
  .A({ S19134 }),
  .ZN({ S19187 })
);
OAI21_X1 #() 
OAI21_X1_1588_ (
  .A({ S25956[27] }),
  .B1({ S19187 }),
  .B2({ S19082 }),
  .ZN({ S19188 })
);
NAND2_X1 #() 
NAND2_X1_3054_ (
  .A1({ S19188 }),
  .A2({ S18113 }),
  .ZN({ S19189 })
);
NAND2_X1 #() 
NAND2_X1_3055_ (
  .A1({ S19189 }),
  .A2({ S18103 }),
  .ZN({ S19190 })
);
OAI221_X1 #() 
OAI221_X1_81_ (
  .A({ S18092 }),
  .B1({ S19185 }),
  .B2({ S18103 }),
  .C1({ S19186 }),
  .C2({ S19190 }),
  .ZN({ S19191 })
);
AND2_X1 #() 
AND2_X1_194_ (
  .A1({ S19179 }),
  .A2({ S19191 }),
  .ZN({ S19192 })
);
OAI21_X1 #() 
OAI21_X1_1589_ (
  .A({ S19165 }),
  .B1({ S19192 }),
  .B2({ S25956[31] }),
  .ZN({ S19193 })
);
XOR2_X1 #() 
XOR2_X1_69_ (
  .A({ S19193 }),
  .B({ S25956[102] }),
  .Z({ S25957[1254] })
);
XNOR2_X1 #() 
XNOR2_X1_162_ (
  .A({ S25957[1254] }),
  .B({ S19127 }),
  .ZN({ S25957[1222] })
);
XOR2_X1 #() 
XOR2_X1_70_ (
  .A({ S25957[1222] }),
  .B({ S25956[38] }),
  .Z({ S25957[1190] })
);
XNOR2_X1 #() 
XNOR2_X1_163_ (
  .A({ S25957[1190] }),
  .B({ S25956[6] }),
  .ZN({ S19194 })
);
INV_X1 #() 
INV_X1_1018_ (
  .A({ S19194 }),
  .ZN({ S25957[1158] })
);
INV_X1 #() 
INV_X1_1019_ (
  .A({ S25956[69] }),
  .ZN({ S19195 })
);
NOR2_X1 #() 
NOR2_X1_779_ (
  .A1({ S18427 }),
  .A2({ S18675 }),
  .ZN({ S19196 })
);
OAI21_X1 #() 
OAI21_X1_1590_ (
  .A({ S18113 }),
  .B1({ S19196 }),
  .B2({ S18165 }),
  .ZN({ S19197 })
);
NAND3_X1 #() 
NAND3_X1_3283_ (
  .A1({ S19030 }),
  .A2({ S18124 }),
  .A3({ S18394 }),
  .ZN({ S19198 })
);
NAND3_X1 #() 
NAND3_X1_3284_ (
  .A1({ S19098 }),
  .A2({ S25956[27] }),
  .A3({ S19144 }),
  .ZN({ S19199 })
);
NAND3_X1 #() 
NAND3_X1_3285_ (
  .A1({ S19199 }),
  .A2({ S25956[28] }),
  .A3({ S19198 }),
  .ZN({ S19200 })
);
NAND3_X1 #() 
NAND3_X1_3286_ (
  .A1({ S19200 }),
  .A2({ S25956[29] }),
  .A3({ S19197 }),
  .ZN({ S19201 })
);
INV_X1 #() 
INV_X1_1020_ (
  .A({ S19146 }),
  .ZN({ S19202 })
);
NAND3_X1 #() 
NAND3_X1_3287_ (
  .A1({ S19202 }),
  .A2({ S18124 }),
  .A3({ S18599 }),
  .ZN({ S19203 })
);
NAND3_X1 #() 
NAND3_X1_3288_ (
  .A1({ S19144 }),
  .A2({ S18124 }),
  .A3({ S18318 }),
  .ZN({ S19204 })
);
NAND2_X1 #() 
NAND2_X1_3056_ (
  .A1({ S19166 }),
  .A2({ S25956[27] }),
  .ZN({ S19205 })
);
AOI21_X1 #() 
AOI21_X1_1683_ (
  .A({ S25956[28] }),
  .B1({ S19205 }),
  .B2({ S19204 }),
  .ZN({ S19206 })
);
AOI21_X1 #() 
AOI21_X1_1684_ (
  .A({ S19206 }),
  .B1({ S19203 }),
  .B2({ S18307 }),
  .ZN({ S19207 })
);
AOI21_X1 #() 
AOI21_X1_1685_ (
  .A({ S18092 }),
  .B1({ S19207 }),
  .B2({ S18103 }),
  .ZN({ S19208 })
);
INV_X1 #() 
INV_X1_1021_ (
  .A({ S18427 }),
  .ZN({ S19209 })
);
NAND3_X1 #() 
NAND3_X1_3289_ (
  .A1({ S19209 }),
  .A2({ S18253 }),
  .A3({ S18567 }),
  .ZN({ S19210 })
);
NAND3_X1 #() 
NAND3_X1_3290_ (
  .A1({ S18307 }),
  .A2({ S18725 }),
  .A3({ S19210 }),
  .ZN({ S19211 })
);
NOR2_X1 #() 
NOR2_X1_780_ (
  .A1({ S18567 }),
  .A2({ S18124 }),
  .ZN({ S19212 })
);
OAI21_X1 #() 
OAI21_X1_1591_ (
  .A({ S18113 }),
  .B1({ S18953 }),
  .B2({ S19212 }),
  .ZN({ S19213 })
);
NAND3_X1 #() 
NAND3_X1_3291_ (
  .A1({ S19211 }),
  .A2({ S18103 }),
  .A3({ S19213 }),
  .ZN({ S19214 })
);
OAI221_X1 #() 
OAI221_X1_82_ (
  .A({ S25956[28] }),
  .B1({ S18253 }),
  .B2({ S18780 }),
  .C1({ S19157 }),
  .C2({ S18124 }),
  .ZN({ S19215 })
);
NAND2_X1 #() 
NAND2_X1_3057_ (
  .A1({ S19202 }),
  .A2({ S19144 }),
  .ZN({ S19216 })
);
AOI21_X1 #() 
AOI21_X1_1686_ (
  .A({ S18329 }),
  .B1({ S19216 }),
  .B2({ S18124 }),
  .ZN({ S19217 })
);
OAI21_X1 #() 
OAI21_X1_1592_ (
  .A({ S19215 }),
  .B1({ S19217 }),
  .B2({ S25956[28] }),
  .ZN({ S19218 })
);
NOR2_X1 #() 
NOR2_X1_781_ (
  .A1({ S19218 }),
  .A2({ S18103 }),
  .ZN({ S19219 })
);
NOR2_X1 #() 
NOR2_X1_782_ (
  .A1({ S19219 }),
  .A2({ S25956[30] }),
  .ZN({ S19220 })
);
AOI22_X1 #() 
AOI22_X1_351_ (
  .A1({ S19201 }),
  .A2({ S19208 }),
  .B1({ S19220 }),
  .B2({ S19214 }),
  .ZN({ S19221 })
);
NAND2_X1 #() 
NAND2_X1_3058_ (
  .A1({ S18209 }),
  .A2({ S18124 }),
  .ZN({ S19222 })
);
NOR2_X1 #() 
NOR2_X1_783_ (
  .A1({ S18253 }),
  .A2({ S25956[25] }),
  .ZN({ S19223 })
);
OAI21_X1 #() 
OAI21_X1_1593_ (
  .A({ S25956[27] }),
  .B1({ S18716 }),
  .B2({ S19223 }),
  .ZN({ S19224 })
);
AOI21_X1 #() 
AOI21_X1_1687_ (
  .A({ S25956[28] }),
  .B1({ S19224 }),
  .B2({ S19222 }),
  .ZN({ S19225 })
);
OAI21_X1 #() 
OAI21_X1_1594_ (
  .A({ S25956[28] }),
  .B1({ S18697 }),
  .B2({ S25956[25] }),
  .ZN({ S19226 })
);
AOI21_X1 #() 
AOI21_X1_1688_ (
  .A({ S19226 }),
  .B1({ S18610 }),
  .B2({ S25956[27] }),
  .ZN({ S19227 })
);
OAI21_X1 #() 
OAI21_X1_1595_ (
  .A({ S18103 }),
  .B1({ S19227 }),
  .B2({ S19225 }),
  .ZN({ S19228 })
);
AOI21_X1 #() 
AOI21_X1_1689_ (
  .A({ S19138 }),
  .B1({ S18253 }),
  .B2({ S18060 }),
  .ZN({ S19229 })
);
AOI21_X1 #() 
AOI21_X1_1690_ (
  .A({ S19229 }),
  .B1({ S19138 }),
  .B2({ S18060 }),
  .ZN({ S19230 })
);
NAND2_X1 #() 
NAND2_X1_3059_ (
  .A1({ S19209 }),
  .A2({ S18481 }),
  .ZN({ S19231 })
);
AOI21_X1 #() 
AOI21_X1_1691_ (
  .A({ S25956[28] }),
  .B1({ S19231 }),
  .B2({ S18545 }),
  .ZN({ S19232 })
);
AOI21_X1 #() 
AOI21_X1_1692_ (
  .A({ S19232 }),
  .B1({ S19230 }),
  .B2({ S25956[28] }),
  .ZN({ S19233 })
);
OAI21_X1 #() 
OAI21_X1_1596_ (
  .A({ S19228 }),
  .B1({ S19233 }),
  .B2({ S18103 }),
  .ZN({ S19234 })
);
AOI22_X1 #() 
AOI22_X1_352_ (
  .A1({ S19209 }),
  .A2({ S19030 }),
  .B1({ S18481 }),
  .B2({ S18165 }),
  .ZN({ S19235 })
);
NOR2_X1 #() 
NOR2_X1_784_ (
  .A1({ S18351 }),
  .A2({ S18124 }),
  .ZN({ S19236 })
);
NAND3_X1 #() 
NAND3_X1_3292_ (
  .A1({ S18780 }),
  .A2({ S18113 }),
  .A3({ S18318 }),
  .ZN({ S19237 })
);
OAI221_X1 #() 
OAI221_X1_83_ (
  .A({ S25956[29] }),
  .B1({ S19236 }),
  .B2({ S19237 }),
  .C1({ S19235 }),
  .C2({ S18113 }),
  .ZN({ S19238 })
);
NAND3_X1 #() 
NAND3_X1_3293_ (
  .A1({ S19111 }),
  .A2({ S18113 }),
  .A3({ S19160 }),
  .ZN({ S19239 })
);
NAND2_X1 #() 
NAND2_X1_3060_ (
  .A1({ S18416 }),
  .A2({ S25956[26] }),
  .ZN({ S19240 })
);
NAND3_X1 #() 
NAND3_X1_3294_ (
  .A1({ S19181 }),
  .A2({ S25956[28] }),
  .A3({ S19240 }),
  .ZN({ S19241 })
);
NAND3_X1 #() 
NAND3_X1_3295_ (
  .A1({ S19239 }),
  .A2({ S18103 }),
  .A3({ S19241 }),
  .ZN({ S19242 })
);
NAND3_X1 #() 
NAND3_X1_3296_ (
  .A1({ S19242 }),
  .A2({ S25956[30] }),
  .A3({ S19238 }),
  .ZN({ S19243 })
);
OAI211_X1 #() 
OAI211_X1_1069_ (
  .A({ S19243 }),
  .B({ S25956[31] }),
  .C1({ S19234 }),
  .C2({ S25956[30] }),
  .ZN({ S19244 })
);
OAI21_X1 #() 
OAI21_X1_1597_ (
  .A({ S19244 }),
  .B1({ S19221 }),
  .B2({ S25956[31] }),
  .ZN({ S19245 })
);
XNOR2_X1 #() 
XNOR2_X1_164_ (
  .A({ S19245 }),
  .B({ S25956[101] }),
  .ZN({ S25957[1253] })
);
XNOR2_X1 #() 
XNOR2_X1_165_ (
  .A({ S25957[1253] }),
  .B({ S19195 }),
  .ZN({ S25957[1221] })
);
XNOR2_X1 #() 
XNOR2_X1_166_ (
  .A({ S25957[1221] }),
  .B({ S25956[37] }),
  .ZN({ S19246 })
);
NAND2_X1 #() 
NAND2_X1_3061_ (
  .A1({ S19246 }),
  .A2({ S11631 }),
  .ZN({ S19247 })
);
INV_X1 #() 
INV_X1_1022_ (
  .A({ S19246 }),
  .ZN({ S25957[1189] })
);
NAND2_X1 #() 
NAND2_X1_3062_ (
  .A1({ S25957[1189] }),
  .A2({ S25956[5] }),
  .ZN({ S19248 })
);
AND2_X1 #() 
AND2_X1_195_ (
  .A1({ S19248 }),
  .A2({ S19247 }),
  .ZN({ S25957[1157] })
);
INV_X1 #() 
INV_X1_1023_ (
  .A({ S25956[68] }),
  .ZN({ S19249 })
);
INV_X1 #() 
INV_X1_1024_ (
  .A({ S25956[100] }),
  .ZN({ S19250 })
);
NOR2_X1 #() 
NOR2_X1_785_ (
  .A1({ S18863 }),
  .A2({ S25956[27] }),
  .ZN({ S19251 })
);
NAND2_X1 #() 
NAND2_X1_3063_ (
  .A1({ S19251 }),
  .A2({ S18242 }),
  .ZN({ S19252 })
);
NAND3_X1 #() 
NAND3_X1_3297_ (
  .A1({ S19252 }),
  .A2({ S18113 }),
  .A3({ S19118 }),
  .ZN({ S19253 })
);
INV_X1 #() 
INV_X1_1025_ (
  .A({ S19152 }),
  .ZN({ S19254 })
);
AOI21_X1 #() 
AOI21_X1_1693_ (
  .A({ S18113 }),
  .B1({ S19209 }),
  .B2({ S18481 }),
  .ZN({ S19255 })
);
NAND2_X1 #() 
NAND2_X1_3064_ (
  .A1({ S18264 }),
  .A2({ S18318 }),
  .ZN({ S19256 })
);
NAND2_X1 #() 
NAND2_X1_3065_ (
  .A1({ S19256 }),
  .A2({ S18124 }),
  .ZN({ S19257 })
);
NOR2_X1 #() 
NOR2_X1_786_ (
  .A1({ S19115 }),
  .A2({ S25956[28] }),
  .ZN({ S19258 })
);
AOI22_X1 #() 
AOI22_X1_353_ (
  .A1({ S19254 }),
  .A2({ S19255 }),
  .B1({ S19258 }),
  .B2({ S19257 }),
  .ZN({ S19259 })
);
NAND2_X1 #() 
NAND2_X1_3066_ (
  .A1({ S18187 }),
  .A2({ S18124 }),
  .ZN({ S19260 })
);
AOI21_X1 #() 
AOI21_X1_1694_ (
  .A({ S18103 }),
  .B1({ S18307 }),
  .B2({ S19260 }),
  .ZN({ S19261 })
);
AOI22_X1 #() 
AOI22_X1_354_ (
  .A1({ S19261 }),
  .A2({ S19253 }),
  .B1({ S19259 }),
  .B2({ S18103 }),
  .ZN({ S19262 })
);
AOI21_X1 #() 
AOI21_X1_1695_ (
  .A({ S25956[27] }),
  .B1({ S18935 }),
  .B2({ S18707 }),
  .ZN({ S19263 })
);
OAI21_X1 #() 
OAI21_X1_1598_ (
  .A({ S25956[27] }),
  .B1({ S18275 }),
  .B2({ S19082 }),
  .ZN({ S19264 })
);
INV_X1 #() 
INV_X1_1026_ (
  .A({ S19264 }),
  .ZN({ S19265 })
);
OAI21_X1 #() 
OAI21_X1_1599_ (
  .A({ S18113 }),
  .B1({ S19263 }),
  .B2({ S19265 }),
  .ZN({ S19266 })
);
OAI211_X1 #() 
OAI211_X1_1070_ (
  .A({ S19144 }),
  .B({ S25956[28] }),
  .C1({ S18567 }),
  .C2({ S18909 }),
  .ZN({ S19267 })
);
AOI21_X1 #() 
AOI21_X1_1696_ (
  .A({ S18103 }),
  .B1({ S19266 }),
  .B2({ S19267 }),
  .ZN({ S19268 })
);
NAND2_X1 #() 
NAND2_X1_3067_ (
  .A1({ S19117 }),
  .A2({ S18383 }),
  .ZN({ S19269 })
);
NAND2_X1 #() 
NAND2_X1_3068_ (
  .A1({ S19240 }),
  .A2({ S18124 }),
  .ZN({ S19270 })
);
NOR2_X1 #() 
NOR2_X1_787_ (
  .A1({ S19270 }),
  .A2({ S19145 }),
  .ZN({ S19271 })
);
NOR2_X1 #() 
NOR2_X1_788_ (
  .A1({ S19271 }),
  .A2({ S25956[28] }),
  .ZN({ S19272 })
);
OAI21_X1 #() 
OAI21_X1_1600_ (
  .A({ S18124 }),
  .B1({ S18340 }),
  .B2({ S18769 }),
  .ZN({ S19273 })
);
OAI21_X1 #() 
OAI21_X1_1601_ (
  .A({ S19273 }),
  .B1({ S19256 }),
  .B2({ S19142 }),
  .ZN({ S19274 })
);
OAI21_X1 #() 
OAI21_X1_1602_ (
  .A({ S18103 }),
  .B1({ S19274 }),
  .B2({ S18113 }),
  .ZN({ S19275 })
);
AOI21_X1 #() 
AOI21_X1_1697_ (
  .A({ S19275 }),
  .B1({ S19272 }),
  .B2({ S19269 }),
  .ZN({ S19276 })
);
OAI21_X1 #() 
OAI21_X1_1603_ (
  .A({ S18092 }),
  .B1({ S19276 }),
  .B2({ S19268 }),
  .ZN({ S19277 })
);
OAI211_X1 #() 
OAI211_X1_1071_ (
  .A({ S19277 }),
  .B({ S25956[31] }),
  .C1({ S19262 }),
  .C2({ S18092 }),
  .ZN({ S19278 })
);
NAND3_X1 #() 
NAND3_X1_3298_ (
  .A1({ S19048 }),
  .A2({ S25956[28] }),
  .A3({ S19270 }),
  .ZN({ S19279 })
);
NOR3_X1 #() 
NOR3_X1_108_ (
  .A1({ S19260 }),
  .A2({ S18863 }),
  .A3({ S18675 }),
  .ZN({ S19280 })
);
NOR2_X1 #() 
NOR2_X1_789_ (
  .A1({ S18874 }),
  .A2({ S18040 }),
  .ZN({ S19281 })
);
OAI21_X1 #() 
OAI21_X1_1604_ (
  .A({ S18113 }),
  .B1({ S19280 }),
  .B2({ S19281 }),
  .ZN({ S19282 })
);
OAI21_X1 #() 
OAI21_X1_1605_ (
  .A({ S19255 }),
  .B1({ S18275 }),
  .B2({ S18874 }),
  .ZN({ S19283 })
);
AOI21_X1 #() 
AOI21_X1_1698_ (
  .A({ S25956[29] }),
  .B1({ S19282 }),
  .B2({ S19283 }),
  .ZN({ S19284 })
);
AOI22_X1 #() 
AOI22_X1_355_ (
  .A1({ S18610 }),
  .A2({ S25956[27] }),
  .B1({ S25956[25] }),
  .B2({ S18502 }),
  .ZN({ S19285 })
);
AOI21_X1 #() 
AOI21_X1_1699_ (
  .A({ S18103 }),
  .B1({ S19285 }),
  .B2({ S18113 }),
  .ZN({ S19286 })
);
AOI21_X1 #() 
AOI21_X1_1700_ (
  .A({ S19284 }),
  .B1({ S19286 }),
  .B2({ S19279 }),
  .ZN({ S19287 })
);
NAND3_X1 #() 
NAND3_X1_3299_ (
  .A1({ S18209 }),
  .A2({ S18124 }),
  .A3({ S19151 }),
  .ZN({ S19288 })
);
NOR2_X1 #() 
NOR2_X1_790_ (
  .A1({ S19138 }),
  .A2({ S25956[28] }),
  .ZN({ S19289 })
);
NAND3_X1 #() 
NAND3_X1_3300_ (
  .A1({ S19114 }),
  .A2({ S18318 }),
  .A3({ S18481 }),
  .ZN({ S19290 })
);
AOI22_X1 #() 
AOI22_X1_356_ (
  .A1({ S18807 }),
  .A2({ S19290 }),
  .B1({ S19288 }),
  .B2({ S19289 }),
  .ZN({ S19291 })
);
NAND2_X1 #() 
NAND2_X1_3069_ (
  .A1({ S18394 }),
  .A2({ S18318 }),
  .ZN({ S19292 })
);
NOR2_X1 #() 
NOR2_X1_791_ (
  .A1({ S18610 }),
  .A2({ S19292 }),
  .ZN({ S19293 })
);
OAI211_X1 #() 
OAI211_X1_1072_ (
  .A({ S19205 }),
  .B({ S18113 }),
  .C1({ S25956[27] }),
  .C2({ S19293 }),
  .ZN({ S19294 })
);
NAND2_X1 #() 
NAND2_X1_3070_ (
  .A1({ S18198 }),
  .A2({ S118 }),
  .ZN({ S19295 })
);
AOI21_X1 #() 
AOI21_X1_1701_ (
  .A({ S18103 }),
  .B1({ S19295 }),
  .B2({ S25956[28] }),
  .ZN({ S19296 })
);
AOI22_X1 #() 
AOI22_X1_357_ (
  .A1({ S19291 }),
  .A2({ S18103 }),
  .B1({ S19294 }),
  .B2({ S19296 }),
  .ZN({ S19297 })
);
OR2_X1 #() 
OR2_X1_42_ (
  .A1({ S19297 }),
  .A2({ S18092 }),
  .ZN({ S19298 })
);
OAI211_X1 #() 
OAI211_X1_1073_ (
  .A({ S19298 }),
  .B({ S18081 }),
  .C1({ S19287 }),
  .C2({ S25956[30] }),
  .ZN({ S19299 })
);
NAND2_X1 #() 
NAND2_X1_3071_ (
  .A1({ S19299 }),
  .A2({ S19278 }),
  .ZN({ S19300 })
);
NAND2_X1 #() 
NAND2_X1_3072_ (
  .A1({ S19300 }),
  .A2({ S19250 }),
  .ZN({ S19301 })
);
NAND3_X1 #() 
NAND3_X1_3301_ (
  .A1({ S19299 }),
  .A2({ S19278 }),
  .A3({ S25956[100] }),
  .ZN({ S19302 })
);
NAND2_X1 #() 
NAND2_X1_3073_ (
  .A1({ S19301 }),
  .A2({ S19302 }),
  .ZN({ S25957[1252] })
);
NAND2_X1 #() 
NAND2_X1_3074_ (
  .A1({ S25957[1252] }),
  .A2({ S19249 }),
  .ZN({ S19303 })
);
INV_X1 #() 
INV_X1_1027_ (
  .A({ S25957[1252] }),
  .ZN({ S19304 })
);
NAND2_X1 #() 
NAND2_X1_3075_ (
  .A1({ S19304 }),
  .A2({ S25956[68] }),
  .ZN({ S19305 })
);
NAND2_X1 #() 
NAND2_X1_3076_ (
  .A1({ S19305 }),
  .A2({ S19303 }),
  .ZN({ S25957[1220] })
);
NOR2_X1 #() 
NOR2_X1_792_ (
  .A1({ S25957[1220] }),
  .A2({ S25956[36] }),
  .ZN({ S19306 })
);
NAND2_X1 #() 
NAND2_X1_3077_ (
  .A1({ S25957[1220] }),
  .A2({ S25956[36] }),
  .ZN({ S19307 })
);
INV_X1 #() 
INV_X1_1028_ (
  .A({ S19307 }),
  .ZN({ S19308 })
);
OAI21_X1 #() 
OAI21_X1_1606_ (
  .A({ S25956[4] }),
  .B1({ S19308 }),
  .B2({ S19306 }),
  .ZN({ S19309 })
);
INV_X1 #() 
INV_X1_1029_ (
  .A({ S25956[36] }),
  .ZN({ S19310 })
);
INV_X1 #() 
INV_X1_1030_ (
  .A({ S25957[1220] }),
  .ZN({ S19311 })
);
NAND2_X1 #() 
NAND2_X1_3078_ (
  .A1({ S19311 }),
  .A2({ S19310 }),
  .ZN({ S19312 })
);
NAND3_X1 #() 
NAND3_X1_3302_ (
  .A1({ S19312 }),
  .A2({ S12118 }),
  .A3({ S19307 }),
  .ZN({ S19313 })
);
NAND2_X1 #() 
NAND2_X1_3079_ (
  .A1({ S19309 }),
  .A2({ S19313 }),
  .ZN({ S25957[1156] })
);
INV_X1 #() 
INV_X1_1031_ (
  .A({ S25956[35] }),
  .ZN({ S19314 })
);
INV_X1 #() 
INV_X1_1032_ (
  .A({ S25956[67] }),
  .ZN({ S19315 })
);
INV_X1 #() 
INV_X1_1033_ (
  .A({ S25956[99] }),
  .ZN({ S19316 })
);
AND4_X1 #() 
AND4_X1_9_ (
  .A1({ S25956[24] }),
  .A2({ S19142 }),
  .A3({ S18113 }),
  .A4({ S18264 }),
  .ZN({ S19317 })
);
NAND2_X1 #() 
NAND2_X1_3080_ (
  .A1({ S19091 }),
  .A2({ S19117 }),
  .ZN({ S19318 })
);
NAND3_X1 #() 
NAND3_X1_3303_ (
  .A1({ S18978 }),
  .A2({ S18790 }),
  .A3({ S19180 }),
  .ZN({ S19319 })
);
NOR2_X1 #() 
NOR2_X1_793_ (
  .A1({ S19183 }),
  .A2({ S18113 }),
  .ZN({ S19320 })
);
AOI22_X1 #() 
AOI22_X1_358_ (
  .A1({ S19319 }),
  .A2({ S18113 }),
  .B1({ S19320 }),
  .B2({ S19318 }),
  .ZN({ S19321 })
);
NAND2_X1 #() 
NAND2_X1_3081_ (
  .A1({ S19158 }),
  .A2({ S25956[28] }),
  .ZN({ S19322 })
);
OAI21_X1 #() 
OAI21_X1_1607_ (
  .A({ S25956[29] }),
  .B1({ S19322 }),
  .B2({ S19098 }),
  .ZN({ S19323 })
);
OAI221_X1 #() 
OAI221_X1_84_ (
  .A({ S18092 }),
  .B1({ S19317 }),
  .B2({ S19323 }),
  .C1({ S19321 }),
  .C2({ S25956[29] }),
  .ZN({ S19324 })
);
NAND3_X1 #() 
NAND3_X1_3304_ (
  .A1({ S19108 }),
  .A2({ S25956[28] }),
  .A3({ S19160 }),
  .ZN({ S19325 })
);
NAND2_X1 #() 
NAND2_X1_3082_ (
  .A1({ S19251 }),
  .A2({ S18567 }),
  .ZN({ S19326 })
);
NAND3_X1 #() 
NAND3_X1_3305_ (
  .A1({ S19326 }),
  .A2({ S18113 }),
  .A3({ S18176 }),
  .ZN({ S19327 })
);
NAND3_X1 #() 
NAND3_X1_3306_ (
  .A1({ S19325 }),
  .A2({ S25956[29] }),
  .A3({ S19327 }),
  .ZN({ S19328 })
);
NAND3_X1 #() 
NAND3_X1_3307_ (
  .A1({ S18060 }),
  .A2({ S18318 }),
  .A3({ S18124 }),
  .ZN({ S19329 })
);
NAND2_X1 #() 
NAND2_X1_3083_ (
  .A1({ S19329 }),
  .A2({ S25956[28] }),
  .ZN({ S19330 })
);
NOR2_X1 #() 
NOR2_X1_794_ (
  .A1({ S18296 }),
  .A2({ S18329 }),
  .ZN({ S19331 })
);
NOR2_X1 #() 
NOR2_X1_795_ (
  .A1({ S18892 }),
  .A2({ S25956[27] }),
  .ZN({ S19332 })
);
NAND2_X1 #() 
NAND2_X1_3084_ (
  .A1({ S19332 }),
  .A2({ S19030 }),
  .ZN({ S19333 })
);
NAND3_X1 #() 
NAND3_X1_3308_ (
  .A1({ S19331 }),
  .A2({ S19333 }),
  .A3({ S18113 }),
  .ZN({ S19334 })
);
NAND3_X1 #() 
NAND3_X1_3309_ (
  .A1({ S19334 }),
  .A2({ S18103 }),
  .A3({ S19330 }),
  .ZN({ S19335 })
);
NAND3_X1 #() 
NAND3_X1_3310_ (
  .A1({ S19328 }),
  .A2({ S25956[30] }),
  .A3({ S19335 }),
  .ZN({ S19336 })
);
NAND3_X1 #() 
NAND3_X1_3311_ (
  .A1({ S19336 }),
  .A2({ S19324 }),
  .A3({ S18081 }),
  .ZN({ S19337 })
);
OAI21_X1 #() 
OAI21_X1_1608_ (
  .A({ S18124 }),
  .B1({ S18588 }),
  .B2({ S18675 }),
  .ZN({ S19338 })
);
OAI21_X1 #() 
OAI21_X1_1609_ (
  .A({ S19338 }),
  .B1({ S18610 }),
  .B2({ S19158 }),
  .ZN({ S19339 })
);
NAND2_X1 #() 
NAND2_X1_3085_ (
  .A1({ S19136 }),
  .A2({ S18481 }),
  .ZN({ S19340 })
);
NAND2_X1 #() 
NAND2_X1_3086_ (
  .A1({ S19216 }),
  .A2({ S25956[27] }),
  .ZN({ S19341 })
);
NAND3_X1 #() 
NAND3_X1_3312_ (
  .A1({ S19340 }),
  .A2({ S18113 }),
  .A3({ S19341 }),
  .ZN({ S19342 })
);
OAI21_X1 #() 
OAI21_X1_1610_ (
  .A({ S19342 }),
  .B1({ S19339 }),
  .B2({ S18113 }),
  .ZN({ S19343 })
);
NAND2_X1 #() 
NAND2_X1_3087_ (
  .A1({ S19091 }),
  .A2({ S19138 }),
  .ZN({ S19344 })
);
OAI21_X1 #() 
OAI21_X1_1611_ (
  .A({ S19344 }),
  .B1({ S18040 }),
  .B2({ S18697 }),
  .ZN({ S19345 })
);
OAI21_X1 #() 
OAI21_X1_1612_ (
  .A({ S18113 }),
  .B1({ S19345 }),
  .B2({ S18556 }),
  .ZN({ S19346 })
);
NAND2_X1 #() 
NAND2_X1_3088_ (
  .A1({ S18935 }),
  .A2({ S25956[27] }),
  .ZN({ S19347 })
);
NAND3_X1 #() 
NAND3_X1_3313_ (
  .A1({ S19347 }),
  .A2({ S25956[28] }),
  .A3({ S19257 }),
  .ZN({ S19348 })
);
NAND3_X1 #() 
NAND3_X1_3314_ (
  .A1({ S19346 }),
  .A2({ S18103 }),
  .A3({ S19348 }),
  .ZN({ S19349 })
);
OAI211_X1 #() 
OAI211_X1_1074_ (
  .A({ S19349 }),
  .B({ S18092 }),
  .C1({ S19343 }),
  .C2({ S18103 }),
  .ZN({ S19350 })
);
NAND2_X1 #() 
NAND2_X1_3089_ (
  .A1({ S18567 }),
  .A2({ S18124 }),
  .ZN({ S19351 })
);
NAND3_X1 #() 
NAND3_X1_3315_ (
  .A1({ S18578 }),
  .A2({ S19134 }),
  .A3({ S25956[27] }),
  .ZN({ S19352 })
);
OAI21_X1 #() 
OAI21_X1_1613_ (
  .A({ S19352 }),
  .B1({ S19169 }),
  .B2({ S19351 }),
  .ZN({ S19353 })
);
NAND2_X1 #() 
NAND2_X1_3090_ (
  .A1({ S19353 }),
  .A2({ S18113 }),
  .ZN({ S19354 })
);
NAND2_X1 #() 
NAND2_X1_3091_ (
  .A1({ S19012 }),
  .A2({ S18567 }),
  .ZN({ S19355 })
);
OAI211_X1 #() 
OAI211_X1_1075_ (
  .A({ S19355 }),
  .B({ S25956[28] }),
  .C1({ S18040 }),
  .C2({ S18874 }),
  .ZN({ S19356 })
);
NAND3_X1 #() 
NAND3_X1_3316_ (
  .A1({ S19354 }),
  .A2({ S25956[29] }),
  .A3({ S19356 }),
  .ZN({ S19357 })
);
OAI221_X1 #() 
OAI221_X1_85_ (
  .A({ S25956[28] }),
  .B1({ S18340 }),
  .B2({ S18124 }),
  .C1({ S19135 }),
  .C2({ S18275 }),
  .ZN({ S19358 })
);
NAND3_X1 #() 
NAND3_X1_3317_ (
  .A1({ S19289 }),
  .A2({ S66 }),
  .A3({ S18686 }),
  .ZN({ S19359 })
);
NAND3_X1 #() 
NAND3_X1_3318_ (
  .A1({ S19358 }),
  .A2({ S18103 }),
  .A3({ S19359 }),
  .ZN({ S19360 })
);
NAND3_X1 #() 
NAND3_X1_3319_ (
  .A1({ S19357 }),
  .A2({ S25956[30] }),
  .A3({ S19360 }),
  .ZN({ S19361 })
);
NAND2_X1 #() 
NAND2_X1_3092_ (
  .A1({ S19350 }),
  .A2({ S19361 }),
  .ZN({ S19362 })
);
NAND2_X1 #() 
NAND2_X1_3093_ (
  .A1({ S19362 }),
  .A2({ S25956[31] }),
  .ZN({ S19363 })
);
NAND3_X1 #() 
NAND3_X1_3320_ (
  .A1({ S19363 }),
  .A2({ S19316 }),
  .A3({ S19337 }),
  .ZN({ S19364 })
);
NAND2_X1 #() 
NAND2_X1_3094_ (
  .A1({ S19363 }),
  .A2({ S19337 }),
  .ZN({ S19365 })
);
NAND2_X1 #() 
NAND2_X1_3095_ (
  .A1({ S19365 }),
  .A2({ S25956[99] }),
  .ZN({ S19366 })
);
NAND2_X1 #() 
NAND2_X1_3096_ (
  .A1({ S19366 }),
  .A2({ S19364 }),
  .ZN({ S25957[1251] })
);
NAND2_X1 #() 
NAND2_X1_3097_ (
  .A1({ S25957[1251] }),
  .A2({ S19315 }),
  .ZN({ S19367 })
);
INV_X1 #() 
INV_X1_1034_ (
  .A({ S25957[1251] }),
  .ZN({ S19368 })
);
NAND2_X1 #() 
NAND2_X1_3098_ (
  .A1({ S19368 }),
  .A2({ S25956[67] }),
  .ZN({ S19369 })
);
NAND3_X1 #() 
NAND3_X1_3321_ (
  .A1({ S19369 }),
  .A2({ S19314 }),
  .A3({ S19367 }),
  .ZN({ S19370 })
);
INV_X1 #() 
INV_X1_1035_ (
  .A({ S19370 }),
  .ZN({ S19371 })
);
AOI21_X1 #() 
AOI21_X1_1702_ (
  .A({ S19314 }),
  .B1({ S19369 }),
  .B2({ S19367 }),
  .ZN({ S19372 })
);
OAI21_X1 #() 
OAI21_X1_1614_ (
  .A({ S11664 }),
  .B1({ S19371 }),
  .B2({ S19372 }),
  .ZN({ S19373 })
);
INV_X1 #() 
INV_X1_1036_ (
  .A({ S19372 }),
  .ZN({ S19374 })
);
NAND3_X1 #() 
NAND3_X1_3322_ (
  .A1({ S19374 }),
  .A2({ S25956[3] }),
  .A3({ S19370 }),
  .ZN({ S19375 })
);
NAND2_X1 #() 
NAND2_X1_3099_ (
  .A1({ S19373 }),
  .A2({ S19375 }),
  .ZN({ S68 })
);
INV_X1 #() 
INV_X1_1037_ (
  .A({ S68 }),
  .ZN({ S25957[1155] })
);
INV_X1 #() 
INV_X1_1038_ (
  .A({ S25956[32] }),
  .ZN({ S19376 })
);
INV_X1 #() 
INV_X1_1039_ (
  .A({ S25956[64] }),
  .ZN({ S19377 })
);
INV_X1 #() 
INV_X1_1040_ (
  .A({ S25956[96] }),
  .ZN({ S19378 })
);
AOI21_X1 #() 
AOI21_X1_1703_ (
  .A({ S19280 }),
  .B1({ S19292 }),
  .B2({ S25956[27] }),
  .ZN({ S19379 })
);
INV_X1 #() 
INV_X1_1041_ (
  .A({ S18610 }),
  .ZN({ S19380 })
);
NAND2_X1 #() 
NAND2_X1_3100_ (
  .A1({ S19380 }),
  .A2({ S19114 }),
  .ZN({ S19381 })
);
NAND3_X1 #() 
NAND3_X1_3323_ (
  .A1({ S19331 }),
  .A2({ S18113 }),
  .A3({ S19381 }),
  .ZN({ S19382 })
);
OAI21_X1 #() 
OAI21_X1_1615_ (
  .A({ S19382 }),
  .B1({ S19379 }),
  .B2({ S18113 }),
  .ZN({ S19383 })
);
NAND2_X1 #() 
NAND2_X1_3101_ (
  .A1({ S19383 }),
  .A2({ S25956[29] }),
  .ZN({ S19384 })
);
AOI21_X1 #() 
AOI21_X1_1704_ (
  .A({ S25956[27] }),
  .B1({ S18578 }),
  .B2({ S19134 }),
  .ZN({ S19385 })
);
AOI21_X1 #() 
AOI21_X1_1705_ (
  .A({ S19385 }),
  .B1({ S19138 }),
  .B2({ S19091 }),
  .ZN({ S19386 })
);
AOI21_X1 #() 
AOI21_X1_1706_ (
  .A({ S25956[28] }),
  .B1({ S19143 }),
  .B2({ S18909 }),
  .ZN({ S19387 })
);
OAI21_X1 #() 
OAI21_X1_1616_ (
  .A({ S19387 }),
  .B1({ S19166 }),
  .B2({ S18124 }),
  .ZN({ S19388 })
);
OAI21_X1 #() 
OAI21_X1_1617_ (
  .A({ S19388 }),
  .B1({ S19386 }),
  .B2({ S18113 }),
  .ZN({ S19389 })
);
NAND2_X1 #() 
NAND2_X1_3102_ (
  .A1({ S19389 }),
  .A2({ S18103 }),
  .ZN({ S19390 })
);
NAND3_X1 #() 
NAND3_X1_3324_ (
  .A1({ S19384 }),
  .A2({ S19390 }),
  .A3({ S25956[30] }),
  .ZN({ S19391 })
);
INV_X1 #() 
INV_X1_1042_ (
  .A({ S18970 }),
  .ZN({ S19392 })
);
AOI21_X1 #() 
AOI21_X1_1707_ (
  .A({ S25956[28] }),
  .B1({ S19264 }),
  .B2({ S19260 }),
  .ZN({ S19393 })
);
AOI21_X1 #() 
AOI21_X1_1708_ (
  .A({ S18113 }),
  .B1({ S19158 }),
  .B2({ S19329 }),
  .ZN({ S19394 })
);
AOI21_X1 #() 
AOI21_X1_1709_ (
  .A({ S19393 }),
  .B1({ S19392 }),
  .B2({ S19394 }),
  .ZN({ S19395 })
);
OAI21_X1 #() 
OAI21_X1_1618_ (
  .A({ S18124 }),
  .B1({ S19082 }),
  .B2({ S18675 }),
  .ZN({ S19396 })
);
AOI21_X1 #() 
AOI21_X1_1710_ (
  .A({ S25956[28] }),
  .B1({ S19396 }),
  .B2({ S18176 }),
  .ZN({ S19397 })
);
AOI21_X1 #() 
AOI21_X1_1711_ (
  .A({ S19140 }),
  .B1({ S18610 }),
  .B2({ S18124 }),
  .ZN({ S19398 })
);
OAI21_X1 #() 
OAI21_X1_1619_ (
  .A({ S18103 }),
  .B1({ S19398 }),
  .B2({ S19397 }),
  .ZN({ S19399 })
);
OAI21_X1 #() 
OAI21_X1_1620_ (
  .A({ S19399 }),
  .B1({ S19395 }),
  .B2({ S18103 }),
  .ZN({ S19400 })
);
OAI21_X1 #() 
OAI21_X1_1621_ (
  .A({ S19391 }),
  .B1({ S19400 }),
  .B2({ S25956[30] }),
  .ZN({ S19401 })
);
NAND2_X1 #() 
NAND2_X1_3103_ (
  .A1({ S19401 }),
  .A2({ S25956[31] }),
  .ZN({ S19402 })
);
NAND2_X1 #() 
NAND2_X1_3104_ (
  .A1({ S19107 }),
  .A2({ S25956[27] }),
  .ZN({ S19403 })
);
NAND2_X1 #() 
NAND2_X1_3105_ (
  .A1({ S19403 }),
  .A2({ S19170 }),
  .ZN({ S19404 })
);
AOI22_X1 #() 
AOI22_X1_359_ (
  .A1({ S19404 }),
  .A2({ S25956[28] }),
  .B1({ S18753 }),
  .B2({ S19188 }),
  .ZN({ S19405 })
);
AOI21_X1 #() 
AOI21_X1_1712_ (
  .A({ S25956[27] }),
  .B1({ S18318 }),
  .B2({ S18383 }),
  .ZN({ S19406 })
);
NAND2_X1 #() 
NAND2_X1_3106_ (
  .A1({ S19205 }),
  .A2({ S18113 }),
  .ZN({ S19407 })
);
INV_X1 #() 
INV_X1_1043_ (
  .A({ S18165 }),
  .ZN({ S19408 })
);
NAND4_X1 #() 
NAND4_X1_354_ (
  .A1({ S19144 }),
  .A2({ S19408 }),
  .A3({ S18394 }),
  .A4({ S25956[28] }),
  .ZN({ S19409 })
);
OAI211_X1 #() 
OAI211_X1_1076_ (
  .A({ S18103 }),
  .B({ S19409 }),
  .C1({ S19407 }),
  .C2({ S19406 }),
  .ZN({ S19410 })
);
OAI21_X1 #() 
OAI21_X1_1622_ (
  .A({ S19410 }),
  .B1({ S19405 }),
  .B2({ S18103 }),
  .ZN({ S19411 })
);
AND3_X1 #() 
AND3_X1_126_ (
  .A1({ S19210 }),
  .A2({ S19153 }),
  .A3({ S18113 }),
  .ZN({ S19412 })
);
AOI21_X1 #() 
AOI21_X1_1713_ (
  .A({ S18113 }),
  .B1({ S19202 }),
  .B2({ S19406 }),
  .ZN({ S19413 })
);
NAND3_X1 #() 
NAND3_X1_3325_ (
  .A1({ S19114 }),
  .A2({ S19030 }),
  .A3({ S18318 }),
  .ZN({ S19414 })
);
OAI21_X1 #() 
OAI21_X1_1623_ (
  .A({ S19414 }),
  .B1({ S18124 }),
  .B2({ S19147 }),
  .ZN({ S19415 })
);
AOI22_X1 #() 
AOI22_X1_360_ (
  .A1({ S19413 }),
  .A2({ S18643 }),
  .B1({ S19415 }),
  .B2({ S18113 }),
  .ZN({ S19416 })
);
NOR3_X1 #() 
NOR3_X1_109_ (
  .A1({ S19196 }),
  .A2({ S19281 }),
  .A3({ S18113 }),
  .ZN({ S19417 })
);
OR2_X1 #() 
OR2_X1_43_ (
  .A1({ S19417 }),
  .A2({ S18103 }),
  .ZN({ S19418 })
);
OAI221_X1 #() 
OAI221_X1_86_ (
  .A({ S18092 }),
  .B1({ S19418 }),
  .B2({ S19412 }),
  .C1({ S19416 }),
  .C2({ S25956[29] }),
  .ZN({ S19419 })
);
OAI21_X1 #() 
OAI21_X1_1624_ (
  .A({ S19419 }),
  .B1({ S19411 }),
  .B2({ S18092 }),
  .ZN({ S19420 })
);
NAND2_X1 #() 
NAND2_X1_3107_ (
  .A1({ S19420 }),
  .A2({ S18081 }),
  .ZN({ S19421 })
);
NAND2_X1 #() 
NAND2_X1_3108_ (
  .A1({ S19402 }),
  .A2({ S19421 }),
  .ZN({ S19422 })
);
NAND2_X1 #() 
NAND2_X1_3109_ (
  .A1({ S19422 }),
  .A2({ S19378 }),
  .ZN({ S19423 })
);
NAND3_X1 #() 
NAND3_X1_3326_ (
  .A1({ S19402 }),
  .A2({ S25956[96] }),
  .A3({ S19421 }),
  .ZN({ S19424 })
);
NAND2_X1 #() 
NAND2_X1_3110_ (
  .A1({ S19423 }),
  .A2({ S19424 }),
  .ZN({ S25957[1248] })
);
NAND2_X1 #() 
NAND2_X1_3111_ (
  .A1({ S25957[1248] }),
  .A2({ S19377 }),
  .ZN({ S19425 })
);
NAND3_X1 #() 
NAND3_X1_3327_ (
  .A1({ S19423 }),
  .A2({ S25956[64] }),
  .A3({ S19424 }),
  .ZN({ S19426 })
);
NAND3_X1 #() 
NAND3_X1_3328_ (
  .A1({ S19425 }),
  .A2({ S19426 }),
  .A3({ S19376 }),
  .ZN({ S19427 })
);
INV_X1 #() 
INV_X1_1044_ (
  .A({ S19427 }),
  .ZN({ S19428 })
);
AOI21_X1 #() 
AOI21_X1_1714_ (
  .A({ S19376 }),
  .B1({ S19425 }),
  .B2({ S19426 }),
  .ZN({ S19429 })
);
OAI21_X1 #() 
OAI21_X1_1625_ (
  .A({ S25956[0] }),
  .B1({ S19428 }),
  .B2({ S19429 }),
  .ZN({ S19430 })
);
INV_X1 #() 
INV_X1_1045_ (
  .A({ S19429 }),
  .ZN({ S19431 })
);
NAND3_X1 #() 
NAND3_X1_3329_ (
  .A1({ S19431 }),
  .A2({ S11550 }),
  .A3({ S19427 }),
  .ZN({ S19432 })
);
NAND2_X1 #() 
NAND2_X1_3112_ (
  .A1({ S19430 }),
  .A2({ S19432 }),
  .ZN({ S25957[1152] })
);
INV_X1 #() 
INV_X1_1046_ (
  .A({ S25956[65] }),
  .ZN({ S19433 })
);
INV_X1 #() 
INV_X1_1047_ (
  .A({ S25956[97] }),
  .ZN({ S19434 })
);
AOI211_X1 #() 
AOI211_X1_47_ (
  .A({ S25956[28] }),
  .B({ S19167 }),
  .C1({ S19098 }),
  .C2({ S25956[27] }),
  .ZN({ S19435 })
);
NAND2_X1 #() 
NAND2_X1_3113_ (
  .A1({ S19269 }),
  .A2({ S18253 }),
  .ZN({ S19436 })
);
AOI211_X1 #() 
AOI211_X1_48_ (
  .A({ S19146 }),
  .B({ S18113 }),
  .C1({ S19436 }),
  .C2({ S18780 }),
  .ZN({ S19437 })
);
OR2_X1 #() 
OR2_X1_44_ (
  .A1({ S19437 }),
  .A2({ S25956[29] }),
  .ZN({ S19438 })
);
NOR2_X1 #() 
NOR2_X1_796_ (
  .A1({ S19260 }),
  .A2({ S18675 }),
  .ZN({ S19439 })
);
AOI21_X1 #() 
AOI21_X1_1715_ (
  .A({ S19439 }),
  .B1({ S19117 }),
  .B2({ S19091 }),
  .ZN({ S19440 })
);
AOI22_X1 #() 
AOI22_X1_361_ (
  .A1({ S18753 }),
  .A2({ S18383 }),
  .B1({ S18113 }),
  .B2({ S18769 }),
  .ZN({ S19441 })
);
OAI211_X1 #() 
OAI211_X1_1077_ (
  .A({ S19441 }),
  .B({ S25956[29] }),
  .C1({ S19440 }),
  .C2({ S18113 }),
  .ZN({ S19442 })
);
OAI21_X1 #() 
OAI21_X1_1626_ (
  .A({ S19442 }),
  .B1({ S19438 }),
  .B2({ S19435 }),
  .ZN({ S19443 })
);
NOR2_X1 #() 
NOR2_X1_797_ (
  .A1({ S18556 }),
  .A2({ S25956[28] }),
  .ZN({ S19444 })
);
AOI22_X1 #() 
AOI22_X1_362_ (
  .A1({ S18807 }),
  .A2({ S19257 }),
  .B1({ S19333 }),
  .B2({ S19444 }),
  .ZN({ S19445 })
);
AOI21_X1 #() 
AOI21_X1_1716_ (
  .A({ S18113 }),
  .B1({ S19341 }),
  .B2({ S19252 }),
  .ZN({ S19446 })
);
NAND2_X1 #() 
NAND2_X1_3114_ (
  .A1({ S18927 }),
  .A2({ S25956[29] }),
  .ZN({ S19447 })
);
OAI221_X1 #() 
OAI221_X1_87_ (
  .A({ S18092 }),
  .B1({ S19446 }),
  .B2({ S19447 }),
  .C1({ S19445 }),
  .C2({ S25956[29] }),
  .ZN({ S19448 })
);
OAI21_X1 #() 
OAI21_X1_1627_ (
  .A({ S19448 }),
  .B1({ S19443 }),
  .B2({ S18092 }),
  .ZN({ S19449 })
);
NAND2_X1 #() 
NAND2_X1_3115_ (
  .A1({ S19449 }),
  .A2({ S18081 }),
  .ZN({ S19450 })
);
NAND3_X1 #() 
NAND3_X1_3330_ (
  .A1({ S19199 }),
  .A2({ S25956[28] }),
  .A3({ S19392 }),
  .ZN({ S19451 })
);
OAI21_X1 #() 
OAI21_X1_1628_ (
  .A({ S19180 }),
  .B1({ S19223 }),
  .B2({ S19329 }),
  .ZN({ S19452 })
);
OAI21_X1 #() 
OAI21_X1_1629_ (
  .A({ S19451 }),
  .B1({ S25956[28] }),
  .B2({ S19452 }),
  .ZN({ S19453 })
);
NOR3_X1 #() 
NOR3_X1_110_ (
  .A1({ S19236 }),
  .A2({ S19332 }),
  .A3({ S18113 }),
  .ZN({ S19454 })
);
NOR2_X1 #() 
NOR2_X1_798_ (
  .A1({ S19107 }),
  .A2({ S18124 }),
  .ZN({ S19455 })
);
NAND3_X1 #() 
NAND3_X1_3331_ (
  .A1({ S18962 }),
  .A2({ S18113 }),
  .A3({ S18492 }),
  .ZN({ S19456 })
);
OAI21_X1 #() 
OAI21_X1_1630_ (
  .A({ S25956[29] }),
  .B1({ S19455 }),
  .B2({ S19456 }),
  .ZN({ S19457 })
);
OAI221_X1 #() 
OAI221_X1_88_ (
  .A({ S25956[30] }),
  .B1({ S19457 }),
  .B2({ S19454 }),
  .C1({ S19453 }),
  .C2({ S25956[29] }),
  .ZN({ S19458 })
);
NAND3_X1 #() 
NAND3_X1_3332_ (
  .A1({ S19326 }),
  .A2({ S19181 }),
  .A3({ S19289 }),
  .ZN({ S19459 })
);
NOR3_X1 #() 
NOR3_X1_111_ (
  .A1({ S18945 }),
  .A2({ S19271 }),
  .A3({ S25956[28] }),
  .ZN({ S19460 })
);
NAND2_X1 #() 
NAND2_X1_3116_ (
  .A1({ S19171 }),
  .A2({ S25956[28] }),
  .ZN({ S19461 })
);
NOR2_X1 #() 
NOR2_X1_799_ (
  .A1({ S18481 }),
  .A2({ S25956[27] }),
  .ZN({ S19462 })
);
AOI211_X1 #() 
AOI211_X1_49_ (
  .A({ S19462 }),
  .B({ S19461 }),
  .C1({ S18351 }),
  .C2({ S18124 }),
  .ZN({ S19463 })
);
NOR3_X1 #() 
NOR3_X1_112_ (
  .A1({ S19460 }),
  .A2({ S19463 }),
  .A3({ S25956[29] }),
  .ZN({ S19464 })
);
OAI21_X1 #() 
OAI21_X1_1631_ (
  .A({ S25956[27] }),
  .B1({ S19128 }),
  .B2({ S19146 }),
  .ZN({ S19465 })
);
AOI21_X1 #() 
AOI21_X1_1717_ (
  .A({ S18103 }),
  .B1({ S19021 }),
  .B2({ S19465 }),
  .ZN({ S19466 })
);
AOI21_X1 #() 
AOI21_X1_1718_ (
  .A({ S19464 }),
  .B1({ S19459 }),
  .B2({ S19466 }),
  .ZN({ S19467 })
);
NAND2_X1 #() 
NAND2_X1_3117_ (
  .A1({ S19467 }),
  .A2({ S18092 }),
  .ZN({ S19468 })
);
NAND3_X1 #() 
NAND3_X1_3333_ (
  .A1({ S19468 }),
  .A2({ S25956[31] }),
  .A3({ S19458 }),
  .ZN({ S19469 })
);
NAND3_X1 #() 
NAND3_X1_3334_ (
  .A1({ S19469 }),
  .A2({ S19450 }),
  .A3({ S19434 }),
  .ZN({ S19470 })
);
NAND2_X1 #() 
NAND2_X1_3118_ (
  .A1({ S19468 }),
  .A2({ S19458 }),
  .ZN({ S19471 })
);
NAND2_X1 #() 
NAND2_X1_3119_ (
  .A1({ S19471 }),
  .A2({ S25956[31] }),
  .ZN({ S19472 })
);
OAI211_X1 #() 
OAI211_X1_1078_ (
  .A({ S19472 }),
  .B({ S25956[97] }),
  .C1({ S25956[31] }),
  .C2({ S19449 }),
  .ZN({ S19473 })
);
NAND3_X1 #() 
NAND3_X1_3335_ (
  .A1({ S19473 }),
  .A2({ S19433 }),
  .A3({ S19470 }),
  .ZN({ S19474 })
);
NAND3_X1 #() 
NAND3_X1_3336_ (
  .A1({ S19469 }),
  .A2({ S19450 }),
  .A3({ S25956[97] }),
  .ZN({ S19475 })
);
OAI211_X1 #() 
OAI211_X1_1079_ (
  .A({ S19472 }),
  .B({ S19434 }),
  .C1({ S25956[31] }),
  .C2({ S19449 }),
  .ZN({ S19476 })
);
NAND3_X1 #() 
NAND3_X1_3337_ (
  .A1({ S19476 }),
  .A2({ S25956[65] }),
  .A3({ S19475 }),
  .ZN({ S19477 })
);
AOI21_X1 #() 
AOI21_X1_1719_ (
  .A({ S25956[33] }),
  .B1({ S19477 }),
  .B2({ S19474 }),
  .ZN({ S19478 })
);
INV_X1 #() 
INV_X1_1048_ (
  .A({ S25956[33] }),
  .ZN({ S19479 })
);
NAND3_X1 #() 
NAND3_X1_3338_ (
  .A1({ S19476 }),
  .A2({ S19433 }),
  .A3({ S19475 }),
  .ZN({ S19480 })
);
NAND3_X1 #() 
NAND3_X1_3339_ (
  .A1({ S19473 }),
  .A2({ S25956[65] }),
  .A3({ S19470 }),
  .ZN({ S19481 })
);
AOI21_X1 #() 
AOI21_X1_1720_ (
  .A({ S19479 }),
  .B1({ S19480 }),
  .B2({ S19481 }),
  .ZN({ S19482 })
);
OAI21_X1 #() 
OAI21_X1_1632_ (
  .A({ S25956[1] }),
  .B1({ S19478 }),
  .B2({ S19482 }),
  .ZN({ S19483 })
);
NAND3_X1 #() 
NAND3_X1_3340_ (
  .A1({ S19480 }),
  .A2({ S19481 }),
  .A3({ S19479 }),
  .ZN({ S19484 })
);
NAND3_X1 #() 
NAND3_X1_3341_ (
  .A1({ S19474 }),
  .A2({ S19477 }),
  .A3({ S25956[33] }),
  .ZN({ S19485 })
);
NAND3_X1 #() 
NAND3_X1_3342_ (
  .A1({ S19484 }),
  .A2({ S19485 }),
  .A3({ S11539 }),
  .ZN({ S19486 })
);
NAND2_X1 #() 
NAND2_X1_3120_ (
  .A1({ S19483 }),
  .A2({ S19486 }),
  .ZN({ S25957[1153] })
);
INV_X1 #() 
INV_X1_1049_ (
  .A({ S25956[34] }),
  .ZN({ S19487 })
);
INV_X1 #() 
INV_X1_1050_ (
  .A({ S25956[66] }),
  .ZN({ S19488 })
);
INV_X1 #() 
INV_X1_1051_ (
  .A({ S25956[98] }),
  .ZN({ S19489 })
);
NAND2_X1 #() 
NAND2_X1_3121_ (
  .A1({ S19175 }),
  .A2({ S25956[27] }),
  .ZN({ S19490 })
);
NOR2_X1 #() 
NOR2_X1_800_ (
  .A1({ S19251 }),
  .A2({ S18113 }),
  .ZN({ S19491 })
);
AOI22_X1 #() 
AOI22_X1_363_ (
  .A1({ S19491 }),
  .A2({ S19490 }),
  .B1({ S19387 }),
  .B2({ S19139 }),
  .ZN({ S19492 })
);
AOI21_X1 #() 
AOI21_X1_1721_ (
  .A({ S18113 }),
  .B1({ S19333 }),
  .B2({ S18790 }),
  .ZN({ S19493 })
);
OAI21_X1 #() 
OAI21_X1_1633_ (
  .A({ S18459 }),
  .B1({ S18124 }),
  .B2({ S18264 }),
  .ZN({ S19494 })
);
OAI211_X1 #() 
OAI211_X1_1080_ (
  .A({ S25956[29] }),
  .B({ S18146 }),
  .C1({ S19494 }),
  .C2({ S25956[28] }),
  .ZN({ S19495 })
);
OAI22_X1 #() 
OAI22_X1_83_ (
  .A1({ S19493 }),
  .A2({ S19495 }),
  .B1({ S19492 }),
  .B2({ S25956[29] }),
  .ZN({ S19496 })
);
AOI21_X1 #() 
AOI21_X1_1722_ (
  .A({ S19226 }),
  .B1({ S18621 }),
  .B2({ S25956[27] }),
  .ZN({ S19497 })
);
NAND2_X1 #() 
NAND2_X1_3122_ (
  .A1({ S18664 }),
  .A2({ S18124 }),
  .ZN({ S19498 })
);
OAI221_X1 #() 
OAI221_X1_89_ (
  .A({ S19498 }),
  .B1({ S18863 }),
  .B2({ S18874 }),
  .C1({ S19380 }),
  .C2({ S25956[27] }),
  .ZN({ S19499 })
);
AOI21_X1 #() 
AOI21_X1_1723_ (
  .A({ S19114 }),
  .B1({ S19293 }),
  .B2({ S25956[27] }),
  .ZN({ S19500 })
);
AOI21_X1 #() 
AOI21_X1_1724_ (
  .A({ S18103 }),
  .B1({ S19500 }),
  .B2({ S18113 }),
  .ZN({ S19501 })
);
OAI21_X1 #() 
OAI21_X1_1634_ (
  .A({ S19501 }),
  .B1({ S18113 }),
  .B2({ S19499 }),
  .ZN({ S19502 })
);
OAI21_X1 #() 
OAI21_X1_1635_ (
  .A({ S19258 }),
  .B1({ S25956[27] }),
  .B2({ S18481 }),
  .ZN({ S19503 })
);
NAND2_X1 #() 
NAND2_X1_3123_ (
  .A1({ S19503 }),
  .A2({ S18103 }),
  .ZN({ S19504 })
);
OAI21_X1 #() 
OAI21_X1_1636_ (
  .A({ S19502 }),
  .B1({ S19497 }),
  .B2({ S19504 }),
  .ZN({ S19505 })
);
NAND2_X1 #() 
NAND2_X1_3124_ (
  .A1({ S19505 }),
  .A2({ S25956[30] }),
  .ZN({ S19506 })
);
OAI211_X1 #() 
OAI211_X1_1081_ (
  .A({ S19506 }),
  .B({ S25956[31] }),
  .C1({ S19496 }),
  .C2({ S25956[30] }),
  .ZN({ S19507 })
);
NAND3_X1 #() 
NAND3_X1_3343_ (
  .A1({ S19381 }),
  .A2({ S19188 }),
  .A3({ S18113 }),
  .ZN({ S19508 })
);
NAND3_X1 #() 
NAND3_X1_3344_ (
  .A1({ S19273 }),
  .A2({ S25956[28] }),
  .A3({ S19490 }),
  .ZN({ S19509 })
);
AOI21_X1 #() 
AOI21_X1_1725_ (
  .A({ S25956[29] }),
  .B1({ S19508 }),
  .B2({ S19509 }),
  .ZN({ S19510 })
);
NAND3_X1 #() 
NAND3_X1_3345_ (
  .A1({ S19202 }),
  .A2({ S25956[27] }),
  .A3({ S18599 }),
  .ZN({ S19511 })
);
NAND2_X1 #() 
NAND2_X1_3125_ (
  .A1({ S19511 }),
  .A2({ S19387 }),
  .ZN({ S19512 })
);
OAI211_X1 #() 
OAI211_X1_1082_ (
  .A({ S19340 }),
  .B({ S25956[28] }),
  .C1({ S19223 }),
  .C2({ S18874 }),
  .ZN({ S19513 })
);
AOI21_X1 #() 
AOI21_X1_1726_ (
  .A({ S18103 }),
  .B1({ S19513 }),
  .B2({ S19512 }),
  .ZN({ S19514 })
);
OR2_X1 #() 
OR2_X1_45_ (
  .A1({ S19514 }),
  .A2({ S19510 }),
  .ZN({ S19515 })
);
OAI21_X1 #() 
OAI21_X1_1637_ (
  .A({ S18113 }),
  .B1({ S19175 }),
  .B2({ S18124 }),
  .ZN({ S19516 })
);
OAI211_X1 #() 
OAI211_X1_1083_ (
  .A({ S19498 }),
  .B({ S19329 }),
  .C1({ S19145 }),
  .C2({ S18874 }),
  .ZN({ S19517 })
);
OAI22_X1 #() 
OAI22_X1_84_ (
  .A1({ S19517 }),
  .A2({ S18113 }),
  .B1({ S19385 }),
  .B2({ S19516 }),
  .ZN({ S19518 })
);
NOR2_X1 #() 
NOR2_X1_801_ (
  .A1({ S19518 }),
  .A2({ S25956[29] }),
  .ZN({ S19519 })
);
AOI21_X1 #() 
AOI21_X1_1727_ (
  .A({ S25956[28] }),
  .B1({ S19251 }),
  .B2({ S25956[24] }),
  .ZN({ S19520 })
);
NAND3_X1 #() 
NAND3_X1_3346_ (
  .A1({ S18643 }),
  .A2({ S18725 }),
  .A3({ S19520 }),
  .ZN({ S19521 })
);
AOI21_X1 #() 
AOI21_X1_1728_ (
  .A({ S18502 }),
  .B1({ S18578 }),
  .B2({ S18264 }),
  .ZN({ S19522 })
);
OAI21_X1 #() 
OAI21_X1_1638_ (
  .A({ S25956[28] }),
  .B1({ S19522 }),
  .B2({ S19462 }),
  .ZN({ S19523 })
);
AOI21_X1 #() 
AOI21_X1_1729_ (
  .A({ S18103 }),
  .B1({ S19521 }),
  .B2({ S19523 }),
  .ZN({ S19524 })
);
OAI21_X1 #() 
OAI21_X1_1639_ (
  .A({ S25956[30] }),
  .B1({ S19519 }),
  .B2({ S19524 }),
  .ZN({ S19525 })
);
OAI211_X1 #() 
OAI211_X1_1084_ (
  .A({ S19525 }),
  .B({ S18081 }),
  .C1({ S19515 }),
  .C2({ S25956[30] }),
  .ZN({ S19526 })
);
NAND3_X1 #() 
NAND3_X1_3347_ (
  .A1({ S19507 }),
  .A2({ S19489 }),
  .A3({ S19526 }),
  .ZN({ S19527 })
);
NAND2_X1 #() 
NAND2_X1_3126_ (
  .A1({ S19507 }),
  .A2({ S19526 }),
  .ZN({ S19528 })
);
NAND2_X1 #() 
NAND2_X1_3127_ (
  .A1({ S19528 }),
  .A2({ S25956[98] }),
  .ZN({ S19529 })
);
NAND2_X1 #() 
NAND2_X1_3128_ (
  .A1({ S19529 }),
  .A2({ S19527 }),
  .ZN({ S19530 })
);
NAND2_X1 #() 
NAND2_X1_3129_ (
  .A1({ S19530 }),
  .A2({ S19488 }),
  .ZN({ S19531 })
);
NAND3_X1 #() 
NAND3_X1_3348_ (
  .A1({ S19529 }),
  .A2({ S19527 }),
  .A3({ S25956[66] }),
  .ZN({ S19532 })
);
NAND3_X1 #() 
NAND3_X1_3349_ (
  .A1({ S19531 }),
  .A2({ S19532 }),
  .A3({ S19487 }),
  .ZN({ S19533 })
);
NAND2_X1 #() 
NAND2_X1_3130_ (
  .A1({ S19531 }),
  .A2({ S19532 }),
  .ZN({ S19534 })
);
NAND2_X1 #() 
NAND2_X1_3131_ (
  .A1({ S19534 }),
  .A2({ S25956[34] }),
  .ZN({ S19535 })
);
NAND3_X1 #() 
NAND3_X1_3350_ (
  .A1({ S19535 }),
  .A2({ S25956[2] }),
  .A3({ S19533 }),
  .ZN({ S19536 })
);
NAND2_X1 #() 
NAND2_X1_3132_ (
  .A1({ S19534 }),
  .A2({ S19487 }),
  .ZN({ S19537 })
);
NAND3_X1 #() 
NAND3_X1_3351_ (
  .A1({ S19531 }),
  .A2({ S19532 }),
  .A3({ S25956[34] }),
  .ZN({ S19538 })
);
NAND3_X1 #() 
NAND3_X1_3352_ (
  .A1({ S19537 }),
  .A2({ S19538 }),
  .A3({ S11642 }),
  .ZN({ S19539 })
);
NAND2_X1 #() 
NAND2_X1_3133_ (
  .A1({ S19536 }),
  .A2({ S19539 }),
  .ZN({ S25957[1154] })
);
NAND2_X1 #() 
NAND2_X1_3134_ (
  .A1({ S10390 }),
  .A2({ S10926 }),
  .ZN({ S69 })
);
NAND2_X1 #() 
NAND2_X1_3135_ (
  .A1({ S25956[16] }),
  .A2({ S25956[17] }),
  .ZN({ S19540 })
);
INV_X1 #() 
INV_X1_1052_ (
  .A({ S19540 }),
  .ZN({ S70 })
);
INV_X1 #() 
INV_X1_1053_ (
  .A({ S25956[22] }),
  .ZN({ S19541 })
);
NAND2_X1 #() 
NAND2_X1_3136_ (
  .A1({ S10390 }),
  .A2({ S25956[17] }),
  .ZN({ S19542 })
);
NAND2_X1 #() 
NAND2_X1_3137_ (
  .A1({ S19542 }),
  .A2({ S9746 }),
  .ZN({ S19543 })
);
NAND2_X1 #() 
NAND2_X1_3138_ (
  .A1({ S10926 }),
  .A2({ S25956[18] }),
  .ZN({ S19544 })
);
NAND2_X1 #() 
NAND2_X1_3139_ (
  .A1({ S19540 }),
  .A2({ S25956[19] }),
  .ZN({ S19545 })
);
INV_X1 #() 
INV_X1_1054_ (
  .A({ S19545 }),
  .ZN({ S19546 })
);
NAND2_X1 #() 
NAND2_X1_3140_ (
  .A1({ S19546 }),
  .A2({ S19544 }),
  .ZN({ S19547 })
);
AOI21_X1 #() 
AOI21_X1_1730_ (
  .A({ S8385 }),
  .B1({ S19547 }),
  .B2({ S19543 }),
  .ZN({ S19548 })
);
NOR2_X1 #() 
NOR2_X1_802_ (
  .A1({ S25956[17] }),
  .A2({ S25956[18] }),
  .ZN({ S19549 })
);
NAND2_X1 #() 
NAND2_X1_3141_ (
  .A1({ S9746 }),
  .A2({ S25956[16] }),
  .ZN({ S19550 })
);
NAND2_X1 #() 
NAND2_X1_3142_ (
  .A1({ S25956[16] }),
  .A2({ S25956[18] }),
  .ZN({ S19551 })
);
NAND2_X1 #() 
NAND2_X1_3143_ (
  .A1({ S25956[17] }),
  .A2({ S25956[18] }),
  .ZN({ S19552 })
);
NAND2_X1 #() 
NAND2_X1_3144_ (
  .A1({ S19551 }),
  .A2({ S19552 }),
  .ZN({ S19553 })
);
AOI211_X1 #() 
AOI211_X1_50_ (
  .A({ S25956[20] }),
  .B({ S19553 }),
  .C1({ S19549 }),
  .C2({ S19550 }),
  .ZN({ S19554 })
);
NOR3_X1 #() 
NOR3_X1_113_ (
  .A1({ S19548 }),
  .A2({ S19554 }),
  .A3({ S25956[21] }),
  .ZN({ S19555 })
);
NAND2_X1 #() 
NAND2_X1_3145_ (
  .A1({ S10926 }),
  .A2({ S25956[16] }),
  .ZN({ S19556 })
);
INV_X1 #() 
INV_X1_1055_ (
  .A({ S19556 }),
  .ZN({ S19557 })
);
INV_X1 #() 
INV_X1_1056_ (
  .A({ S19552 }),
  .ZN({ S19558 })
);
NAND2_X1 #() 
NAND2_X1_3146_ (
  .A1({ S19558 }),
  .A2({ S10390 }),
  .ZN({ S19559 })
);
NAND2_X1 #() 
NAND2_X1_3147_ (
  .A1({ S19559 }),
  .A2({ S25956[19] }),
  .ZN({ S19560 })
);
NOR2_X1 #() 
NOR2_X1_803_ (
  .A1({ S19540 }),
  .A2({ S25956[18] }),
  .ZN({ S19561 })
);
NOR2_X1 #() 
NOR2_X1_804_ (
  .A1({ S25956[16] }),
  .A2({ S25956[17] }),
  .ZN({ S19562 })
);
NAND2_X1 #() 
NAND2_X1_3148_ (
  .A1({ S19562 }),
  .A2({ S25956[18] }),
  .ZN({ S19563 })
);
NAND2_X1 #() 
NAND2_X1_3149_ (
  .A1({ S19563 }),
  .A2({ S9746 }),
  .ZN({ S19564 })
);
OAI22_X1 #() 
OAI22_X1_85_ (
  .A1({ S19560 }),
  .A2({ S19557 }),
  .B1({ S19564 }),
  .B2({ S19561 }),
  .ZN({ S19565 })
);
NAND2_X1 #() 
NAND2_X1_3150_ (
  .A1({ S19565 }),
  .A2({ S8385 }),
  .ZN({ S19566 })
);
NAND2_X1 #() 
NAND2_X1_3151_ (
  .A1({ S10390 }),
  .A2({ S11487 }),
  .ZN({ S19567 })
);
NAND2_X1 #() 
NAND2_X1_3152_ (
  .A1({ S19567 }),
  .A2({ S9746 }),
  .ZN({ S19568 })
);
NAND2_X1 #() 
NAND2_X1_3153_ (
  .A1({ S11487 }),
  .A2({ S25956[17] }),
  .ZN({ S19569 })
);
NAND2_X1 #() 
NAND2_X1_3154_ (
  .A1({ S19567 }),
  .A2({ S19569 }),
  .ZN({ S19570 })
);
NAND2_X1 #() 
NAND2_X1_3155_ (
  .A1({ S19570 }),
  .A2({ S25956[19] }),
  .ZN({ S19571 })
);
NOR2_X1 #() 
NOR2_X1_805_ (
  .A1({ S19551 }),
  .A2({ S9746 }),
  .ZN({ S19572 })
);
INV_X1 #() 
INV_X1_1057_ (
  .A({ S19572 }),
  .ZN({ S19573 })
);
NAND2_X1 #() 
NAND2_X1_3156_ (
  .A1({ S19571 }),
  .A2({ S19573 }),
  .ZN({ S19574 })
);
INV_X1 #() 
INV_X1_1058_ (
  .A({ S19574 }),
  .ZN({ S19575 })
);
OAI21_X1 #() 
OAI21_X1_1640_ (
  .A({ S19575 }),
  .B1({ S10926 }),
  .B2({ S19568 }),
  .ZN({ S19576 })
);
OAI21_X1 #() 
OAI21_X1_1641_ (
  .A({ S19566 }),
  .B1({ S19576 }),
  .B2({ S8385 }),
  .ZN({ S19577 })
);
AOI21_X1 #() 
AOI21_X1_1731_ (
  .A({ S19555 }),
  .B1({ S19577 }),
  .B2({ S25956[21] }),
  .ZN({ S19578 })
);
NOR2_X1 #() 
NOR2_X1_806_ (
  .A1({ S19578 }),
  .A2({ S19541 }),
  .ZN({ S19579 })
);
NAND2_X1 #() 
NAND2_X1_3157_ (
  .A1({ S19551 }),
  .A2({ S25956[19] }),
  .ZN({ S19580 })
);
INV_X1 #() 
INV_X1_1059_ (
  .A({ S19580 }),
  .ZN({ S19581 })
);
NAND2_X1 #() 
NAND2_X1_3158_ (
  .A1({ S19581 }),
  .A2({ S19569 }),
  .ZN({ S19582 })
);
NAND2_X1 #() 
NAND2_X1_3159_ (
  .A1({ S19540 }),
  .A2({ S25956[18] }),
  .ZN({ S19583 })
);
NAND2_X1 #() 
NAND2_X1_3160_ (
  .A1({ S19556 }),
  .A2({ S11487 }),
  .ZN({ S19584 })
);
NAND2_X1 #() 
NAND2_X1_3161_ (
  .A1({ S19584 }),
  .A2({ S19583 }),
  .ZN({ S19585 })
);
AOI21_X1 #() 
AOI21_X1_1732_ (
  .A({ S25956[20] }),
  .B1({ S19585 }),
  .B2({ S9746 }),
  .ZN({ S19586 })
);
NAND2_X1 #() 
NAND2_X1_3162_ (
  .A1({ S19586 }),
  .A2({ S19582 }),
  .ZN({ S19587 })
);
NAND2_X1 #() 
NAND2_X1_3163_ (
  .A1({ S19570 }),
  .A2({ S19542 }),
  .ZN({ S19588 })
);
AOI21_X1 #() 
AOI21_X1_1733_ (
  .A({ S9746 }),
  .B1({ S19588 }),
  .B2({ S19583 }),
  .ZN({ S19589 })
);
NOR2_X1 #() 
NOR2_X1_807_ (
  .A1({ S25956[16] }),
  .A2({ S25956[18] }),
  .ZN({ S19590 })
);
INV_X1 #() 
INV_X1_1060_ (
  .A({ S19551 }),
  .ZN({ S19591 })
);
NAND2_X1 #() 
NAND2_X1_3164_ (
  .A1({ S19591 }),
  .A2({ S25956[17] }),
  .ZN({ S19592 })
);
NAND2_X1 #() 
NAND2_X1_3165_ (
  .A1({ S19592 }),
  .A2({ S19563 }),
  .ZN({ S19593 })
);
OAI21_X1 #() 
OAI21_X1_1642_ (
  .A({ S9746 }),
  .B1({ S19593 }),
  .B2({ S19590 }),
  .ZN({ S19594 })
);
NAND2_X1 #() 
NAND2_X1_3166_ (
  .A1({ S19594 }),
  .A2({ S25956[20] }),
  .ZN({ S19595 })
);
OAI21_X1 #() 
OAI21_X1_1643_ (
  .A({ S19587 }),
  .B1({ S19595 }),
  .B2({ S19589 }),
  .ZN({ S19596 })
);
NAND2_X1 #() 
NAND2_X1_3167_ (
  .A1({ S19563 }),
  .A2({ S25956[19] }),
  .ZN({ S19597 })
);
NAND2_X1 #() 
NAND2_X1_3168_ (
  .A1({ S19552 }),
  .A2({ S9746 }),
  .ZN({ S19598 })
);
NAND2_X1 #() 
NAND2_X1_3169_ (
  .A1({ S19598 }),
  .A2({ S19550 }),
  .ZN({ S19599 })
);
AOI21_X1 #() 
AOI21_X1_1734_ (
  .A({ S8385 }),
  .B1({ S19599 }),
  .B2({ S19567 }),
  .ZN({ S19600 })
);
OAI21_X1 #() 
OAI21_X1_1644_ (
  .A({ S19600 }),
  .B1({ S19561 }),
  .B2({ S19597 }),
  .ZN({ S19601 })
);
INV_X1 #() 
INV_X1_1061_ (
  .A({ S19583 }),
  .ZN({ S19602 })
);
NAND2_X1 #() 
NAND2_X1_3170_ (
  .A1({ S19602 }),
  .A2({ S9746 }),
  .ZN({ S19603 })
);
INV_X1 #() 
INV_X1_1062_ (
  .A({ S19544 }),
  .ZN({ S19604 })
);
OAI21_X1 #() 
OAI21_X1_1645_ (
  .A({ S25956[19] }),
  .B1({ S19570 }),
  .B2({ S19604 }),
  .ZN({ S19605 })
);
AND2_X1 #() 
AND2_X1_196_ (
  .A1({ S19605 }),
  .A2({ S19603 }),
  .ZN({ S19606 })
);
OAI21_X1 #() 
OAI21_X1_1646_ (
  .A({ S19601 }),
  .B1({ S19606 }),
  .B2({ S25956[20] }),
  .ZN({ S19607 })
);
NAND2_X1 #() 
NAND2_X1_3171_ (
  .A1({ S19607 }),
  .A2({ S25956[21] }),
  .ZN({ S19608 })
);
OAI211_X1 #() 
OAI211_X1_1085_ (
  .A({ S19608 }),
  .B({ S25956[22] }),
  .C1({ S25956[21] }),
  .C2({ S19596 }),
  .ZN({ S19609 })
);
NAND2_X1 #() 
NAND2_X1_3172_ (
  .A1({ S19593 }),
  .A2({ S9746 }),
  .ZN({ S19610 })
);
OAI211_X1 #() 
OAI211_X1_1086_ (
  .A({ S19610 }),
  .B({ S8385 }),
  .C1({ S11487 }),
  .C2({ S19545 }),
  .ZN({ S19611 })
);
NAND2_X1 #() 
NAND2_X1_3173_ (
  .A1({ S19553 }),
  .A2({ S19540 }),
  .ZN({ S19612 })
);
INV_X1 #() 
INV_X1_1063_ (
  .A({ S19561 }),
  .ZN({ S19613 })
);
NAND3_X1 #() 
NAND3_X1_3353_ (
  .A1({ S19612 }),
  .A2({ S19613 }),
  .A3({ S9746 }),
  .ZN({ S19614 })
);
AOI21_X1 #() 
AOI21_X1_1735_ (
  .A({ S8385 }),
  .B1({ S19559 }),
  .B2({ S25956[19] }),
  .ZN({ S19615 })
);
AOI21_X1 #() 
AOI21_X1_1736_ (
  .A({ S25956[21] }),
  .B1({ S19614 }),
  .B2({ S19615 }),
  .ZN({ S19616 })
);
NAND2_X1 #() 
NAND2_X1_3174_ (
  .A1({ S19540 }),
  .A2({ S11487 }),
  .ZN({ S19617 })
);
INV_X1 #() 
INV_X1_1064_ (
  .A({ S19598 }),
  .ZN({ S19618 })
);
NAND2_X1 #() 
NAND2_X1_3175_ (
  .A1({ S19618 }),
  .A2({ S19617 }),
  .ZN({ S19619 })
);
NAND3_X1 #() 
NAND3_X1_3354_ (
  .A1({ S19569 }),
  .A2({ S19556 }),
  .A3({ S25956[19] }),
  .ZN({ S19620 })
);
AOI21_X1 #() 
AOI21_X1_1737_ (
  .A({ S25956[20] }),
  .B1({ S19619 }),
  .B2({ S19620 }),
  .ZN({ S19621 })
);
NAND2_X1 #() 
NAND2_X1_3176_ (
  .A1({ S10926 }),
  .A2({ S11487 }),
  .ZN({ S19622 })
);
NAND2_X1 #() 
NAND2_X1_3177_ (
  .A1({ S19581 }),
  .A2({ S19622 }),
  .ZN({ S19623 })
);
INV_X1 #() 
INV_X1_1065_ (
  .A({ S19550 }),
  .ZN({ S19624 })
);
NOR2_X1 #() 
NOR2_X1_808_ (
  .A1({ S19624 }),
  .A2({ S8385 }),
  .ZN({ S19625 })
);
AOI21_X1 #() 
AOI21_X1_1738_ (
  .A({ S19621 }),
  .B1({ S19623 }),
  .B2({ S19625 }),
  .ZN({ S19626 })
);
AOI22_X1 #() 
AOI22_X1_364_ (
  .A1({ S19626 }),
  .A2({ S25956[21] }),
  .B1({ S19611 }),
  .B2({ S19616 }),
  .ZN({ S19627 })
);
OAI211_X1 #() 
OAI211_X1_1087_ (
  .A({ S19609 }),
  .B({ S5675 }),
  .C1({ S25956[22] }),
  .C2({ S19627 }),
  .ZN({ S19628 })
);
NOR2_X1 #() 
NOR2_X1_809_ (
  .A1({ S10926 }),
  .A2({ S25956[19] }),
  .ZN({ S19629 })
);
NAND2_X1 #() 
NAND2_X1_3178_ (
  .A1({ S10926 }),
  .A2({ S25956[19] }),
  .ZN({ S19630 })
);
NAND2_X1 #() 
NAND2_X1_3179_ (
  .A1({ S19573 }),
  .A2({ S19630 }),
  .ZN({ S19631 })
);
AOI211_X1 #() 
AOI211_X1_51_ (
  .A({ S8385 }),
  .B({ S19631 }),
  .C1({ S19551 }),
  .C2({ S19629 }),
  .ZN({ S19632 })
);
NAND2_X1 #() 
NAND2_X1_3180_ (
  .A1({ S19556 }),
  .A2({ S25956[18] }),
  .ZN({ S19633 })
);
NOR2_X1 #() 
NOR2_X1_810_ (
  .A1({ S19617 }),
  .A2({ S19562 }),
  .ZN({ S19634 })
);
INV_X1 #() 
INV_X1_1066_ (
  .A({ S19634 }),
  .ZN({ S19635 })
);
NAND2_X1 #() 
NAND2_X1_3181_ (
  .A1({ S19635 }),
  .A2({ S19633 }),
  .ZN({ S19636 })
);
NAND2_X1 #() 
NAND2_X1_3182_ (
  .A1({ S19636 }),
  .A2({ S9746 }),
  .ZN({ S19637 })
);
NAND2_X1 #() 
NAND2_X1_3183_ (
  .A1({ S19622 }),
  .A2({ S25956[19] }),
  .ZN({ S19638 })
);
NAND3_X1 #() 
NAND3_X1_3355_ (
  .A1({ S19637 }),
  .A2({ S8385 }),
  .A3({ S19638 }),
  .ZN({ S19639 })
);
AOI21_X1 #() 
AOI21_X1_1739_ (
  .A({ S9746 }),
  .B1({ S19588 }),
  .B2({ S19612 }),
  .ZN({ S19640 })
);
NAND2_X1 #() 
NAND2_X1_3184_ (
  .A1({ S11487 }),
  .A2({ S25956[16] }),
  .ZN({ S19641 })
);
NAND2_X1 #() 
NAND2_X1_3185_ (
  .A1({ S19641 }),
  .A2({ S9746 }),
  .ZN({ S19642 })
);
OAI21_X1 #() 
OAI21_X1_1647_ (
  .A({ S25956[20] }),
  .B1({ S19642 }),
  .B2({ S19558 }),
  .ZN({ S19643 })
);
OAI21_X1 #() 
OAI21_X1_1648_ (
  .A({ S19639 }),
  .B1({ S19640 }),
  .B2({ S19643 }),
  .ZN({ S19644 })
);
AOI21_X1 #() 
AOI21_X1_1740_ (
  .A({ S25956[20] }),
  .B1({ S19567 }),
  .B2({ S9746 }),
  .ZN({ S19645 })
);
NOR2_X1 #() 
NOR2_X1_811_ (
  .A1({ S9746 }),
  .A2({ S25956[16] }),
  .ZN({ S19646 })
);
OAI21_X1 #() 
OAI21_X1_1649_ (
  .A({ S19645 }),
  .B1({ S10926 }),
  .B2({ S19646 }),
  .ZN({ S19647 })
);
NAND2_X1 #() 
NAND2_X1_3186_ (
  .A1({ S19647 }),
  .A2({ S25956[21] }),
  .ZN({ S19648 })
);
OAI22_X1 #() 
OAI22_X1_86_ (
  .A1({ S19644 }),
  .A2({ S25956[21] }),
  .B1({ S19632 }),
  .B2({ S19648 }),
  .ZN({ S19649 })
);
OAI21_X1 #() 
OAI21_X1_1650_ (
  .A({ S25956[23] }),
  .B1({ S19649 }),
  .B2({ S25956[22] }),
  .ZN({ S19650 })
);
OAI21_X1 #() 
OAI21_X1_1651_ (
  .A({ S19628 }),
  .B1({ S19650 }),
  .B2({ S19579 }),
  .ZN({ S19651 })
);
XNOR2_X1 #() 
XNOR2_X1_167_ (
  .A({ S19651 }),
  .B({ S25956[127] }),
  .ZN({ S25957[1279] })
);
INV_X1 #() 
INV_X1_1067_ (
  .A({ S25957[1279] }),
  .ZN({ S19652 })
);
OR2_X1 #() 
OR2_X1_46_ (
  .A1({ S19652 }),
  .A2({ S25956[95] }),
  .ZN({ S19653 })
);
NAND2_X1 #() 
NAND2_X1_3187_ (
  .A1({ S19652 }),
  .A2({ S25956[95] }),
  .ZN({ S19654 })
);
NAND2_X1 #() 
NAND2_X1_3188_ (
  .A1({ S19653 }),
  .A2({ S19654 }),
  .ZN({ S25957[1247] })
);
NOR2_X1 #() 
NOR2_X1_812_ (
  .A1({ S25957[1247] }),
  .A2({ S25956[63] }),
  .ZN({ S19655 })
);
NAND2_X1 #() 
NAND2_X1_3189_ (
  .A1({ S25957[1247] }),
  .A2({ S25956[63] }),
  .ZN({ S19656 })
);
INV_X1 #() 
INV_X1_1068_ (
  .A({ S19656 }),
  .ZN({ S19657 })
);
OAI21_X1 #() 
OAI21_X1_1652_ (
  .A({ S25956[31] }),
  .B1({ S19657 }),
  .B2({ S19655 }),
  .ZN({ S19658 })
);
NOR2_X1 #() 
NOR2_X1_813_ (
  .A1({ S19657 }),
  .A2({ S19655 }),
  .ZN({ S25957[1215] })
);
NAND2_X1 #() 
NAND2_X1_3190_ (
  .A1({ S25957[1215] }),
  .A2({ S18081 }),
  .ZN({ S19659 })
);
NAND2_X1 #() 
NAND2_X1_3191_ (
  .A1({ S19659 }),
  .A2({ S19658 }),
  .ZN({ S25957[1183] })
);
INV_X1 #() 
INV_X1_1069_ (
  .A({ S25956[62] }),
  .ZN({ S19660 })
);
INV_X1 #() 
INV_X1_1070_ (
  .A({ S25956[94] }),
  .ZN({ S19661 })
);
NAND3_X1 #() 
NAND3_X1_3356_ (
  .A1({ S19563 }),
  .A2({ S25956[19] }),
  .A3({ S19617 }),
  .ZN({ S19662 })
);
OAI21_X1 #() 
OAI21_X1_1653_ (
  .A({ S9746 }),
  .B1({ S19634 }),
  .B2({ S19591 }),
  .ZN({ S19663 })
);
NAND2_X1 #() 
NAND2_X1_3192_ (
  .A1({ S19633 }),
  .A2({ S19641 }),
  .ZN({ S19664 })
);
AOI21_X1 #() 
AOI21_X1_1741_ (
  .A({ S8385 }),
  .B1({ S19664 }),
  .B2({ S25956[19] }),
  .ZN({ S19665 })
);
AOI22_X1 #() 
AOI22_X1_365_ (
  .A1({ S19586 }),
  .A2({ S19662 }),
  .B1({ S19665 }),
  .B2({ S19663 }),
  .ZN({ S19666 })
);
NAND2_X1 #() 
NAND2_X1_3193_ (
  .A1({ S10390 }),
  .A2({ S25956[18] }),
  .ZN({ S19667 })
);
NOR2_X1 #() 
NOR2_X1_814_ (
  .A1({ S10390 }),
  .A2({ S25956[18] }),
  .ZN({ S19668 })
);
NOR2_X1 #() 
NOR2_X1_815_ (
  .A1({ S19668 }),
  .A2({ S19630 }),
  .ZN({ S19669 })
);
NAND2_X1 #() 
NAND2_X1_3194_ (
  .A1({ S19669 }),
  .A2({ S19667 }),
  .ZN({ S19670 })
);
NAND2_X1 #() 
NAND2_X1_3195_ (
  .A1({ S19553 }),
  .A2({ S9746 }),
  .ZN({ S19671 })
);
AOI21_X1 #() 
AOI21_X1_1742_ (
  .A({ S8385 }),
  .B1({ S19670 }),
  .B2({ S19671 }),
  .ZN({ S19672 })
);
NOR2_X1 #() 
NOR2_X1_816_ (
  .A1({ S19629 }),
  .A2({ S25956[20] }),
  .ZN({ S19673 })
);
AOI21_X1 #() 
AOI21_X1_1743_ (
  .A({ S19672 }),
  .B1({ S19547 }),
  .B2({ S19673 }),
  .ZN({ S19674 })
);
MUX2_X1 #() 
MUX2_X1_13_ (
  .A({ S19666 }),
  .B({ S19674 }),
  .S({ S25956[21] }),
  .Z({ S19675 })
);
NOR2_X1 #() 
NOR2_X1_817_ (
  .A1({ S19552 }),
  .A2({ S25956[16] }),
  .ZN({ S19676 })
);
OAI21_X1 #() 
OAI21_X1_1654_ (
  .A({ S25956[19] }),
  .B1({ S19676 }),
  .B2({ S19668 }),
  .ZN({ S19677 })
);
NAND3_X1 #() 
NAND3_X1_3357_ (
  .A1({ S19663 }),
  .A2({ S8385 }),
  .A3({ S19677 }),
  .ZN({ S19678 })
);
NOR2_X1 #() 
NOR2_X1_818_ (
  .A1({ S19584 }),
  .A2({ S25956[19] }),
  .ZN({ S19679 })
);
OAI21_X1 #() 
OAI21_X1_1655_ (
  .A({ S25956[20] }),
  .B1({ S19631 }),
  .B2({ S19679 }),
  .ZN({ S19680 })
);
NAND3_X1 #() 
NAND3_X1_3358_ (
  .A1({ S19678 }),
  .A2({ S7762 }),
  .A3({ S19680 }),
  .ZN({ S19681 })
);
NOR2_X1 #() 
NOR2_X1_819_ (
  .A1({ S10926 }),
  .A2({ S25956[16] }),
  .ZN({ S19682 })
);
NAND2_X1 #() 
NAND2_X1_3196_ (
  .A1({ S19682 }),
  .A2({ S11487 }),
  .ZN({ S19683 })
);
INV_X1 #() 
INV_X1_1071_ (
  .A({ S19683 }),
  .ZN({ S19684 })
);
NOR2_X1 #() 
NOR2_X1_820_ (
  .A1({ S19593 }),
  .A2({ S19684 }),
  .ZN({ S19685 })
);
NOR2_X1 #() 
NOR2_X1_821_ (
  .A1({ S19685 }),
  .A2({ S25956[19] }),
  .ZN({ S19686 })
);
NAND2_X1 #() 
NAND2_X1_3197_ (
  .A1({ S19558 }),
  .A2({ S25956[19] }),
  .ZN({ S19687 })
);
NAND2_X1 #() 
NAND2_X1_3198_ (
  .A1({ S19687 }),
  .A2({ S25956[20] }),
  .ZN({ S19688 })
);
NAND2_X1 #() 
NAND2_X1_3199_ (
  .A1({ S19552 }),
  .A2({ S25956[16] }),
  .ZN({ S19689 })
);
NAND2_X1 #() 
NAND2_X1_3200_ (
  .A1({ S19689 }),
  .A2({ S19542 }),
  .ZN({ S19690 })
);
NAND2_X1 #() 
NAND2_X1_3201_ (
  .A1({ S19690 }),
  .A2({ S9746 }),
  .ZN({ S19691 })
);
OAI21_X1 #() 
OAI21_X1_1656_ (
  .A({ S25956[19] }),
  .B1({ S19684 }),
  .B2({ S19604 }),
  .ZN({ S19692 })
);
NAND3_X1 #() 
NAND3_X1_3359_ (
  .A1({ S19692 }),
  .A2({ S8385 }),
  .A3({ S19691 }),
  .ZN({ S19693 })
);
OAI211_X1 #() 
OAI211_X1_1088_ (
  .A({ S19693 }),
  .B({ S25956[21] }),
  .C1({ S19686 }),
  .C2({ S19688 }),
  .ZN({ S19694 })
);
NAND3_X1 #() 
NAND3_X1_3360_ (
  .A1({ S19694 }),
  .A2({ S19541 }),
  .A3({ S19681 }),
  .ZN({ S19695 })
);
OAI21_X1 #() 
OAI21_X1_1657_ (
  .A({ S19695 }),
  .B1({ S19675 }),
  .B2({ S19541 }),
  .ZN({ S19696 })
);
NOR2_X1 #() 
NOR2_X1_822_ (
  .A1({ S19602 }),
  .A2({ S19668 }),
  .ZN({ S19697 })
);
OAI221_X1 #() 
OAI221_X1_90_ (
  .A({ S25956[20] }),
  .B1({ S19682 }),
  .B2({ S19580 }),
  .C1({ S19697 }),
  .C2({ S25956[19] }),
  .ZN({ S19698 })
);
AOI22_X1 #() 
AOI22_X1_366_ (
  .A1({ S19542 }),
  .A2({ S19551 }),
  .B1({ S10926 }),
  .B2({ S9746 }),
  .ZN({ S19699 })
);
OAI21_X1 #() 
OAI21_X1_1658_ (
  .A({ S19698 }),
  .B1({ S25956[20] }),
  .B2({ S19699 }),
  .ZN({ S19700 })
);
NOR2_X1 #() 
NOR2_X1_823_ (
  .A1({ S19549 }),
  .A2({ S25956[19] }),
  .ZN({ S19701 })
);
INV_X1 #() 
INV_X1_1072_ (
  .A({ S19701 }),
  .ZN({ S19702 })
);
OAI221_X1 #() 
OAI221_X1_91_ (
  .A({ S25956[20] }),
  .B1({ S19569 }),
  .B2({ S9746 }),
  .C1({ S19702 }),
  .C2({ S25956[16] }),
  .ZN({ S19703 })
);
NAND2_X1 #() 
NAND2_X1_3202_ (
  .A1({ S19664 }),
  .A2({ S25956[19] }),
  .ZN({ S19704 })
);
NAND2_X1 #() 
NAND2_X1_3203_ (
  .A1({ S19618 }),
  .A2({ S19551 }),
  .ZN({ S19705 })
);
NAND2_X1 #() 
NAND2_X1_3204_ (
  .A1({ S70 }),
  .A2({ S9746 }),
  .ZN({ S19706 })
);
NAND4_X1 #() 
NAND4_X1_355_ (
  .A1({ S19704 }),
  .A2({ S8385 }),
  .A3({ S19705 }),
  .A4({ S19706 }),
  .ZN({ S19707 })
);
NAND3_X1 #() 
NAND3_X1_3361_ (
  .A1({ S19707 }),
  .A2({ S7762 }),
  .A3({ S19703 }),
  .ZN({ S19708 })
);
OAI21_X1 #() 
OAI21_X1_1659_ (
  .A({ S19708 }),
  .B1({ S19700 }),
  .B2({ S7762 }),
  .ZN({ S19709 })
);
INV_X1 #() 
INV_X1_1073_ (
  .A({ S19563 }),
  .ZN({ S19710 })
);
OAI211_X1 #() 
OAI211_X1_1089_ (
  .A({ S25956[20] }),
  .B({ S19642 }),
  .C1({ S19710 }),
  .C2({ S19545 }),
  .ZN({ S19711 })
);
NAND2_X1 #() 
NAND2_X1_3205_ (
  .A1({ S19544 }),
  .A2({ S25956[19] }),
  .ZN({ S19712 })
);
NOR2_X1 #() 
NOR2_X1_824_ (
  .A1({ S10926 }),
  .A2({ S25956[18] }),
  .ZN({ S19713 })
);
NAND2_X1 #() 
NAND2_X1_3206_ (
  .A1({ S19668 }),
  .A2({ S10926 }),
  .ZN({ S19714 })
);
NAND2_X1 #() 
NAND2_X1_3207_ (
  .A1({ S19714 }),
  .A2({ S19618 }),
  .ZN({ S19715 })
);
OAI211_X1 #() 
OAI211_X1_1090_ (
  .A({ S19715 }),
  .B({ S8385 }),
  .C1({ S19712 }),
  .C2({ S19713 }),
  .ZN({ S19716 })
);
AOI21_X1 #() 
AOI21_X1_1744_ (
  .A({ S7762 }),
  .B1({ S19716 }),
  .B2({ S19711 }),
  .ZN({ S19717 })
);
NAND2_X1 #() 
NAND2_X1_3208_ (
  .A1({ S19542 }),
  .A2({ S11487 }),
  .ZN({ S19718 })
);
NAND2_X1 #() 
NAND2_X1_3209_ (
  .A1({ S19559 }),
  .A2({ S19718 }),
  .ZN({ S19719 })
);
NAND2_X1 #() 
NAND2_X1_3210_ (
  .A1({ S19719 }),
  .A2({ S25956[19] }),
  .ZN({ S19720 })
);
NAND2_X1 #() 
NAND2_X1_3211_ (
  .A1({ S19720 }),
  .A2({ S8385 }),
  .ZN({ S19721 })
);
OAI211_X1 #() 
OAI211_X1_1091_ (
  .A({ S19605 }),
  .B({ S25956[20] }),
  .C1({ S19622 }),
  .C2({ S19550 }),
  .ZN({ S19722 })
);
AOI21_X1 #() 
AOI21_X1_1745_ (
  .A({ S25956[21] }),
  .B1({ S19722 }),
  .B2({ S19721 }),
  .ZN({ S19723 })
);
OAI21_X1 #() 
OAI21_X1_1660_ (
  .A({ S19541 }),
  .B1({ S19717 }),
  .B2({ S19723 }),
  .ZN({ S19724 })
);
OAI21_X1 #() 
OAI21_X1_1661_ (
  .A({ S19724 }),
  .B1({ S19709 }),
  .B2({ S19541 }),
  .ZN({ S19725 })
);
MUX2_X1 #() 
MUX2_X1_14_ (
  .A({ S19725 }),
  .B({ S19696 }),
  .S({ S25956[23] }),
  .Z({ S19726 })
);
XNOR2_X1 #() 
XNOR2_X1_168_ (
  .A({ S19726 }),
  .B({ S25956[126] }),
  .ZN({ S19727 })
);
INV_X1 #() 
INV_X1_1074_ (
  .A({ S19727 }),
  .ZN({ S25957[1278] })
);
NAND2_X1 #() 
NAND2_X1_3212_ (
  .A1({ S25957[1278] }),
  .A2({ S19661 }),
  .ZN({ S19728 })
);
NAND2_X1 #() 
NAND2_X1_3213_ (
  .A1({ S19727 }),
  .A2({ S25956[94] }),
  .ZN({ S19729 })
);
NAND3_X1 #() 
NAND3_X1_3362_ (
  .A1({ S19728 }),
  .A2({ S19729 }),
  .A3({ S19660 }),
  .ZN({ S19730 })
);
INV_X1 #() 
INV_X1_1075_ (
  .A({ S19730 }),
  .ZN({ S19731 })
);
AOI21_X1 #() 
AOI21_X1_1746_ (
  .A({ S19660 }),
  .B1({ S19728 }),
  .B2({ S19729 }),
  .ZN({ S19732 })
);
OAI21_X1 #() 
OAI21_X1_1662_ (
  .A({ S25956[30] }),
  .B1({ S19731 }),
  .B2({ S19732 }),
  .ZN({ S19733 })
);
INV_X1 #() 
INV_X1_1076_ (
  .A({ S19732 }),
  .ZN({ S19734 })
);
NAND3_X1 #() 
NAND3_X1_3363_ (
  .A1({ S19734 }),
  .A2({ S18092 }),
  .A3({ S19730 }),
  .ZN({ S19735 })
);
NAND2_X1 #() 
NAND2_X1_3214_ (
  .A1({ S19733 }),
  .A2({ S19735 }),
  .ZN({ S25957[1182] })
);
INV_X1 #() 
INV_X1_1077_ (
  .A({ S25956[93] }),
  .ZN({ S19736 })
);
AOI22_X1 #() 
AOI22_X1_367_ (
  .A1({ S19557 }),
  .A2({ S25956[19] }),
  .B1({ S19629 }),
  .B2({ S19591 }),
  .ZN({ S19737 })
);
NAND3_X1 #() 
NAND3_X1_3364_ (
  .A1({ S19714 }),
  .A2({ S19592 }),
  .A3({ S19563 }),
  .ZN({ S19738 })
);
NOR2_X1 #() 
NOR2_X1_825_ (
  .A1({ S19738 }),
  .A2({ S9746 }),
  .ZN({ S19739 })
);
NAND4_X1 #() 
NAND4_X1_356_ (
  .A1({ S19567 }),
  .A2({ S19556 }),
  .A3({ S19542 }),
  .A4({ S9746 }),
  .ZN({ S19740 })
);
NAND2_X1 #() 
NAND2_X1_3215_ (
  .A1({ S19740 }),
  .A2({ S25956[20] }),
  .ZN({ S19741 })
);
OAI221_X1 #() 
OAI221_X1_92_ (
  .A({ S7762 }),
  .B1({ S25956[20] }),
  .B2({ S19737 }),
  .C1({ S19739 }),
  .C2({ S19741 }),
  .ZN({ S19742 })
);
NAND2_X1 #() 
NAND2_X1_3216_ (
  .A1({ S19629 }),
  .A2({ S19590 }),
  .ZN({ S19743 })
);
AOI21_X1 #() 
AOI21_X1_1747_ (
  .A({ S8385 }),
  .B1({ S19617 }),
  .B2({ S25956[19] }),
  .ZN({ S19744 })
);
NAND2_X1 #() 
NAND2_X1_3217_ (
  .A1({ S19683 }),
  .A2({ S19592 }),
  .ZN({ S19745 })
);
INV_X1 #() 
INV_X1_1078_ (
  .A({ S19745 }),
  .ZN({ S19746 })
);
AOI21_X1 #() 
AOI21_X1_1748_ (
  .A({ S19581 }),
  .B1({ S19746 }),
  .B2({ S9746 }),
  .ZN({ S19747 })
);
AOI22_X1 #() 
AOI22_X1_368_ (
  .A1({ S19747 }),
  .A2({ S8385 }),
  .B1({ S19743 }),
  .B2({ S19744 }),
  .ZN({ S19748 })
);
AOI21_X1 #() 
AOI21_X1_1749_ (
  .A({ S25956[22] }),
  .B1({ S19748 }),
  .B2({ S25956[21] }),
  .ZN({ S19749 })
);
INV_X1 #() 
INV_X1_1079_ (
  .A({ S19646 }),
  .ZN({ S19750 })
);
NOR2_X1 #() 
NOR2_X1_826_ (
  .A1({ S19682 }),
  .A2({ S25956[19] }),
  .ZN({ S19751 })
);
NAND2_X1 #() 
NAND2_X1_3218_ (
  .A1({ S19751 }),
  .A2({ S19641 }),
  .ZN({ S19752 })
);
AOI21_X1 #() 
AOI21_X1_1750_ (
  .A({ S25956[20] }),
  .B1({ S19752 }),
  .B2({ S19750 }),
  .ZN({ S19753 })
);
OAI21_X1 #() 
OAI21_X1_1663_ (
  .A({ S19715 }),
  .B1({ S19685 }),
  .B2({ S9746 }),
  .ZN({ S19754 })
);
AOI21_X1 #() 
AOI21_X1_1751_ (
  .A({ S19753 }),
  .B1({ S19754 }),
  .B2({ S25956[20] }),
  .ZN({ S19755 })
);
NAND2_X1 #() 
NAND2_X1_3219_ (
  .A1({ S19755 }),
  .A2({ S25956[21] }),
  .ZN({ S19756 })
);
INV_X1 #() 
INV_X1_1080_ (
  .A({ S19571 }),
  .ZN({ S19757 })
);
NOR2_X1 #() 
NOR2_X1_827_ (
  .A1({ S19757 }),
  .A2({ S8385 }),
  .ZN({ S19758 })
);
AND2_X1 #() 
AND2_X1_197_ (
  .A1({ S19592 }),
  .A2({ S19617 }),
  .ZN({ S19759 })
);
NAND2_X1 #() 
NAND2_X1_3220_ (
  .A1({ S19759 }),
  .A2({ S9746 }),
  .ZN({ S19760 })
);
NAND2_X1 #() 
NAND2_X1_3221_ (
  .A1({ S19542 }),
  .A2({ S19551 }),
  .ZN({ S19761 })
);
NAND2_X1 #() 
NAND2_X1_3222_ (
  .A1({ S19761 }),
  .A2({ S19667 }),
  .ZN({ S19762 })
);
INV_X1 #() 
INV_X1_1081_ (
  .A({ S19762 }),
  .ZN({ S19763 })
);
NAND2_X1 #() 
NAND2_X1_3223_ (
  .A1({ S19697 }),
  .A2({ S25956[19] }),
  .ZN({ S19764 })
);
OAI21_X1 #() 
OAI21_X1_1664_ (
  .A({ S19764 }),
  .B1({ S25956[19] }),
  .B2({ S19763 }),
  .ZN({ S19765 })
);
AOI22_X1 #() 
AOI22_X1_369_ (
  .A1({ S19765 }),
  .A2({ S8385 }),
  .B1({ S19758 }),
  .B2({ S19760 }),
  .ZN({ S19766 })
);
AOI21_X1 #() 
AOI21_X1_1752_ (
  .A({ S19541 }),
  .B1({ S19766 }),
  .B2({ S7762 }),
  .ZN({ S19767 })
);
AOI22_X1 #() 
AOI22_X1_370_ (
  .A1({ S19767 }),
  .A2({ S19756 }),
  .B1({ S19749 }),
  .B2({ S19742 }),
  .ZN({ S19768 })
);
NAND2_X1 #() 
NAND2_X1_3224_ (
  .A1({ S19768 }),
  .A2({ S5675 }),
  .ZN({ S19769 })
);
NAND3_X1 #() 
NAND3_X1_3365_ (
  .A1({ S19610 }),
  .A2({ S19704 }),
  .A3({ S8385 }),
  .ZN({ S19770 })
);
INV_X1 #() 
INV_X1_1082_ (
  .A({ S19718 }),
  .ZN({ S19771 })
);
AOI21_X1 #() 
AOI21_X1_1753_ (
  .A({ S19771 }),
  .B1({ S19682 }),
  .B2({ S9746 }),
  .ZN({ S19772 })
);
OAI211_X1 #() 
OAI211_X1_1092_ (
  .A({ S19770 }),
  .B({ S7762 }),
  .C1({ S8385 }),
  .C2({ S19772 }),
  .ZN({ S19773 })
);
OAI21_X1 #() 
OAI21_X1_1665_ (
  .A({ S9746 }),
  .B1({ S19591 }),
  .B2({ S25956[17] }),
  .ZN({ S19774 })
);
NAND2_X1 #() 
NAND2_X1_3225_ (
  .A1({ S19546 }),
  .A2({ S19552 }),
  .ZN({ S19775 })
);
NAND3_X1 #() 
NAND3_X1_3366_ (
  .A1({ S19775 }),
  .A2({ S19573 }),
  .A3({ S19774 }),
  .ZN({ S19776 })
);
OAI221_X1 #() 
OAI221_X1_93_ (
  .A({ S25956[20] }),
  .B1({ S19638 }),
  .B2({ S25956[16] }),
  .C1({ S19570 }),
  .C2({ S19543 }),
  .ZN({ S19777 })
);
INV_X1 #() 
INV_X1_1083_ (
  .A({ S19777 }),
  .ZN({ S19778 })
);
AOI21_X1 #() 
AOI21_X1_1754_ (
  .A({ S19778 }),
  .B1({ S19776 }),
  .B2({ S8385 }),
  .ZN({ S19779 })
);
OAI21_X1 #() 
OAI21_X1_1666_ (
  .A({ S19773 }),
  .B1({ S19779 }),
  .B2({ S7762 }),
  .ZN({ S19780 })
);
NAND2_X1 #() 
NAND2_X1_3226_ (
  .A1({ S19613 }),
  .A2({ S9746 }),
  .ZN({ S19781 })
);
NOR2_X1 #() 
NOR2_X1_828_ (
  .A1({ S19583 }),
  .A2({ S19562 }),
  .ZN({ S19782 })
);
NAND2_X1 #() 
NAND2_X1_3227_ (
  .A1({ S19549 }),
  .A2({ S10390 }),
  .ZN({ S19783 })
);
INV_X1 #() 
INV_X1_1084_ (
  .A({ S19783 }),
  .ZN({ S19784 })
);
OAI21_X1 #() 
OAI21_X1_1667_ (
  .A({ S25956[19] }),
  .B1({ S19782 }),
  .B2({ S19784 }),
  .ZN({ S19785 })
);
AOI21_X1 #() 
AOI21_X1_1755_ (
  .A({ S25956[20] }),
  .B1({ S19785 }),
  .B2({ S19781 }),
  .ZN({ S19786 })
);
NAND3_X1 #() 
NAND3_X1_3367_ (
  .A1({ S19641 }),
  .A2({ S9746 }),
  .A3({ S10926 }),
  .ZN({ S19787 })
);
NOR2_X1 #() 
NOR2_X1_829_ (
  .A1({ S19562 }),
  .A2({ S25956[18] }),
  .ZN({ S19788 })
);
AOI21_X1 #() 
AOI21_X1_1756_ (
  .A({ S8385 }),
  .B1({ S19546 }),
  .B2({ S19788 }),
  .ZN({ S19789 })
);
AOI21_X1 #() 
AOI21_X1_1757_ (
  .A({ S19786 }),
  .B1({ S19787 }),
  .B2({ S19789 }),
  .ZN({ S19790 })
);
NOR2_X1 #() 
NOR2_X1_830_ (
  .A1({ S9746 }),
  .A2({ S11487 }),
  .ZN({ S19791 })
);
NAND2_X1 #() 
NAND2_X1_3228_ (
  .A1({ S19667 }),
  .A2({ S19556 }),
  .ZN({ S19792 })
);
OAI22_X1 #() 
OAI22_X1_87_ (
  .A1({ S19792 }),
  .A2({ S19791 }),
  .B1({ S19545 }),
  .B2({ S11487 }),
  .ZN({ S19793 })
);
INV_X1 #() 
INV_X1_1085_ (
  .A({ S19630 }),
  .ZN({ S19794 })
);
NOR2_X1 #() 
NOR2_X1_831_ (
  .A1({ S19543 }),
  .A2({ S19549 }),
  .ZN({ S19795 })
);
OAI21_X1 #() 
OAI21_X1_1668_ (
  .A({ S8385 }),
  .B1({ S19795 }),
  .B2({ S19794 }),
  .ZN({ S19796 })
);
OAI21_X1 #() 
OAI21_X1_1669_ (
  .A({ S19796 }),
  .B1({ S19793 }),
  .B2({ S8385 }),
  .ZN({ S19797 })
);
NAND2_X1 #() 
NAND2_X1_3229_ (
  .A1({ S19797 }),
  .A2({ S25956[21] }),
  .ZN({ S19798 })
);
OAI21_X1 #() 
OAI21_X1_1670_ (
  .A({ S19798 }),
  .B1({ S19790 }),
  .B2({ S25956[21] }),
  .ZN({ S19799 })
);
MUX2_X1 #() 
MUX2_X1_15_ (
  .A({ S19799 }),
  .B({ S19780 }),
  .S({ S25956[22] }),
  .Z({ S19800 })
);
OAI211_X1 #() 
OAI211_X1_1093_ (
  .A({ S19769 }),
  .B({ S25956[125] }),
  .C1({ S19800 }),
  .C2({ S5675 }),
  .ZN({ S19801 })
);
INV_X1 #() 
INV_X1_1086_ (
  .A({ S25956[125] }),
  .ZN({ S19802 })
);
NAND2_X1 #() 
NAND2_X1_3230_ (
  .A1({ S19800 }),
  .A2({ S25956[23] }),
  .ZN({ S19803 })
);
OAI211_X1 #() 
OAI211_X1_1094_ (
  .A({ S19803 }),
  .B({ S19802 }),
  .C1({ S19768 }),
  .C2({ S25956[23] }),
  .ZN({ S19804 })
);
NAND3_X1 #() 
NAND3_X1_3368_ (
  .A1({ S19804 }),
  .A2({ S19736 }),
  .A3({ S19801 }),
  .ZN({ S19805 })
);
INV_X1 #() 
INV_X1_1087_ (
  .A({ S19805 }),
  .ZN({ S19806 })
);
AOI21_X1 #() 
AOI21_X1_1758_ (
  .A({ S19736 }),
  .B1({ S19804 }),
  .B2({ S19801 }),
  .ZN({ S19807 })
);
OAI21_X1 #() 
OAI21_X1_1671_ (
  .A({ S25956[61] }),
  .B1({ S19806 }),
  .B2({ S19807 }),
  .ZN({ S19808 })
);
INV_X1 #() 
INV_X1_1088_ (
  .A({ S25956[61] }),
  .ZN({ S19809 })
);
INV_X1 #() 
INV_X1_1089_ (
  .A({ S19807 }),
  .ZN({ S19810 })
);
NAND3_X1 #() 
NAND3_X1_3369_ (
  .A1({ S19810 }),
  .A2({ S19809 }),
  .A3({ S19805 }),
  .ZN({ S19811 })
);
NAND2_X1 #() 
NAND2_X1_3231_ (
  .A1({ S19808 }),
  .A2({ S19811 }),
  .ZN({ S25957[1213] })
);
NAND2_X1 #() 
NAND2_X1_3232_ (
  .A1({ S25957[1213] }),
  .A2({ S18103 }),
  .ZN({ S19812 })
);
NAND3_X1 #() 
NAND3_X1_3370_ (
  .A1({ S19808 }),
  .A2({ S19811 }),
  .A3({ S25956[29] }),
  .ZN({ S19813 })
);
NAND2_X1 #() 
NAND2_X1_3233_ (
  .A1({ S19812 }),
  .A2({ S19813 }),
  .ZN({ S25957[1181] })
);
INV_X1 #() 
INV_X1_1090_ (
  .A({ S25956[92] }),
  .ZN({ S19814 })
);
INV_X1 #() 
INV_X1_1091_ (
  .A({ S25956[124] }),
  .ZN({ S19815 })
);
AND2_X1 #() 
AND2_X1_198_ (
  .A1({ S11487 }),
  .A2({ S119 }),
  .ZN({ S19816 })
);
NAND2_X1 #() 
NAND2_X1_3234_ (
  .A1({ S19544 }),
  .A2({ S19551 }),
  .ZN({ S19817 })
);
OAI21_X1 #() 
OAI21_X1_1672_ (
  .A({ S9746 }),
  .B1({ S19634 }),
  .B2({ S19817 }),
  .ZN({ S19818 })
);
NAND3_X1 #() 
NAND3_X1_3371_ (
  .A1({ S19764 }),
  .A2({ S19818 }),
  .A3({ S8385 }),
  .ZN({ S19819 })
);
OAI211_X1 #() 
OAI211_X1_1095_ (
  .A({ S19819 }),
  .B({ S25956[21] }),
  .C1({ S8385 }),
  .C2({ S19816 }),
  .ZN({ S19820 })
);
NAND3_X1 #() 
NAND3_X1_3372_ (
  .A1({ S19613 }),
  .A2({ S9746 }),
  .A3({ S19667 }),
  .ZN({ S19821 })
);
NOR2_X1 #() 
NOR2_X1_832_ (
  .A1({ S19791 }),
  .A2({ S25956[20] }),
  .ZN({ S19822 })
);
NOR2_X1 #() 
NOR2_X1_833_ (
  .A1({ S19705 }),
  .A2({ S19549 }),
  .ZN({ S19823 })
);
NOR2_X1 #() 
NOR2_X1_834_ (
  .A1({ S19823 }),
  .A2({ S19631 }),
  .ZN({ S19824 })
);
AOI22_X1 #() 
AOI22_X1_371_ (
  .A1({ S19824 }),
  .A2({ S25956[20] }),
  .B1({ S19821 }),
  .B2({ S19822 }),
  .ZN({ S19825 })
);
NAND2_X1 #() 
NAND2_X1_3235_ (
  .A1({ S19825 }),
  .A2({ S7762 }),
  .ZN({ S19826 })
);
NAND2_X1 #() 
NAND2_X1_3236_ (
  .A1({ S19826 }),
  .A2({ S19820 }),
  .ZN({ S19827 })
);
OAI211_X1 #() 
OAI211_X1_1096_ (
  .A({ S19605 }),
  .B({ S25956[20] }),
  .C1({ S25956[19] }),
  .C2({ S19817 }),
  .ZN({ S19828 })
);
OAI211_X1 #() 
OAI211_X1_1097_ (
  .A({ S8385 }),
  .B({ S19706 }),
  .C1({ S19635 }),
  .C2({ S9746 }),
  .ZN({ S19829 })
);
AND2_X1 #() 
AND2_X1_199_ (
  .A1({ S19828 }),
  .A2({ S19829 }),
  .ZN({ S19830 })
);
NOR2_X1 #() 
NOR2_X1_835_ (
  .A1({ S19564 }),
  .A2({ S19788 }),
  .ZN({ S19831 })
);
NOR2_X1 #() 
NOR2_X1_836_ (
  .A1({ S19580 }),
  .A2({ S19562 }),
  .ZN({ S19832 })
);
OAI21_X1 #() 
OAI21_X1_1673_ (
  .A({ S8385 }),
  .B1({ S19831 }),
  .B2({ S19832 }),
  .ZN({ S19833 })
);
OAI221_X1 #() 
OAI221_X1_94_ (
  .A({ S25956[20] }),
  .B1({ S19543 }),
  .B2({ S19549 }),
  .C1({ S19570 }),
  .C2({ S19580 }),
  .ZN({ S19834 })
);
AOI21_X1 #() 
AOI21_X1_1759_ (
  .A({ S25956[21] }),
  .B1({ S19833 }),
  .B2({ S19834 }),
  .ZN({ S19835 })
);
AOI21_X1 #() 
AOI21_X1_1760_ (
  .A({ S19835 }),
  .B1({ S19830 }),
  .B2({ S25956[21] }),
  .ZN({ S19836 })
);
NAND2_X1 #() 
NAND2_X1_3237_ (
  .A1({ S19836 }),
  .A2({ S19541 }),
  .ZN({ S19837 })
);
OAI211_X1 #() 
OAI211_X1_1098_ (
  .A({ S19837 }),
  .B({ S5675 }),
  .C1({ S19827 }),
  .C2({ S19541 }),
  .ZN({ S19838 })
);
NOR2_X1 #() 
NOR2_X1_837_ (
  .A1({ S19713 }),
  .A2({ S25956[19] }),
  .ZN({ S19839 })
);
NAND2_X1 #() 
NAND2_X1_3238_ (
  .A1({ S19839 }),
  .A2({ S10390 }),
  .ZN({ S19840 })
);
AOI21_X1 #() 
AOI21_X1_1761_ (
  .A({ S25956[20] }),
  .B1({ S19840 }),
  .B2({ S19623 }),
  .ZN({ S19841 })
);
AOI21_X1 #() 
AOI21_X1_1762_ (
  .A({ S8385 }),
  .B1({ S19571 }),
  .B2({ S19564 }),
  .ZN({ S19842 })
);
OR3_X1 #() 
OR3_X1_17_ (
  .A1({ S19841 }),
  .A2({ S19842 }),
  .A3({ S19541 }),
  .ZN({ S19843 })
);
AOI21_X1 #() 
AOI21_X1_1763_ (
  .A({ S25956[19] }),
  .B1({ S19588 }),
  .B2({ S19583 }),
  .ZN({ S19844 })
);
OAI21_X1 #() 
OAI21_X1_1674_ (
  .A({ S25956[19] }),
  .B1({ S19570 }),
  .B2({ S19682 }),
  .ZN({ S19845 })
);
INV_X1 #() 
INV_X1_1092_ (
  .A({ S19845 }),
  .ZN({ S19846 })
);
OAI21_X1 #() 
OAI21_X1_1675_ (
  .A({ S8385 }),
  .B1({ S19844 }),
  .B2({ S19846 }),
  .ZN({ S19847 })
);
NOR2_X1 #() 
NOR2_X1_838_ (
  .A1({ S25956[19] }),
  .A2({ S25956[18] }),
  .ZN({ S19848 })
);
OAI211_X1 #() 
OAI211_X1_1099_ (
  .A({ S19683 }),
  .B({ S25956[20] }),
  .C1({ S19556 }),
  .C2({ S19848 }),
  .ZN({ S19849 })
);
NAND3_X1 #() 
NAND3_X1_3373_ (
  .A1({ S19847 }),
  .A2({ S19541 }),
  .A3({ S19849 }),
  .ZN({ S19850 })
);
AOI21_X1 #() 
AOI21_X1_1764_ (
  .A({ S7762 }),
  .B1({ S19850 }),
  .B2({ S19843 }),
  .ZN({ S19851 })
);
NAND2_X1 #() 
NAND2_X1_3239_ (
  .A1({ S19701 }),
  .A2({ S19667 }),
  .ZN({ S19852 })
);
AND2_X1 #() 
AND2_X1_200_ (
  .A1({ S19852 }),
  .A2({ S19620 }),
  .ZN({ S19853 })
);
OAI21_X1 #() 
OAI21_X1_1676_ (
  .A({ S25956[20] }),
  .B1({ S19795 }),
  .B2({ S19669 }),
  .ZN({ S19854 })
);
OAI211_X1 #() 
OAI211_X1_1100_ (
  .A({ S19854 }),
  .B({ S25956[22] }),
  .C1({ S19853 }),
  .C2({ S25956[20] }),
  .ZN({ S19855 })
);
NOR2_X1 #() 
NOR2_X1_839_ (
  .A1({ S19591 }),
  .A2({ S19630 }),
  .ZN({ S19856 })
);
NAND2_X1 #() 
NAND2_X1_3240_ (
  .A1({ S19719 }),
  .A2({ S9746 }),
  .ZN({ S19857 })
);
NAND2_X1 #() 
NAND2_X1_3241_ (
  .A1({ S19857 }),
  .A2({ S8385 }),
  .ZN({ S19858 })
);
NOR2_X1 #() 
NOR2_X1_840_ (
  .A1({ S19858 }),
  .A2({ S19856 }),
  .ZN({ S19859 })
);
INV_X1 #() 
INV_X1_1093_ (
  .A({ S19617 }),
  .ZN({ S19860 })
);
OAI21_X1 #() 
OAI21_X1_1677_ (
  .A({ S9746 }),
  .B1({ S19860 }),
  .B2({ S19817 }),
  .ZN({ S19861 })
);
OAI21_X1 #() 
OAI21_X1_1678_ (
  .A({ S19861 }),
  .B1({ S19604 }),
  .B2({ S19582 }),
  .ZN({ S19862 })
);
NOR2_X1 #() 
NOR2_X1_841_ (
  .A1({ S19862 }),
  .A2({ S8385 }),
  .ZN({ S19863 })
);
OAI21_X1 #() 
OAI21_X1_1679_ (
  .A({ S19541 }),
  .B1({ S19859 }),
  .B2({ S19863 }),
  .ZN({ S19864 })
);
AOI21_X1 #() 
AOI21_X1_1765_ (
  .A({ S25956[21] }),
  .B1({ S19864 }),
  .B2({ S19855 }),
  .ZN({ S19865 })
);
OR3_X1 #() 
OR3_X1_18_ (
  .A1({ S19865 }),
  .A2({ S19851 }),
  .A3({ S5675 }),
  .ZN({ S19866 })
);
NAND3_X1 #() 
NAND3_X1_3374_ (
  .A1({ S19866 }),
  .A2({ S19815 }),
  .A3({ S19838 }),
  .ZN({ S19867 })
);
OAI21_X1 #() 
OAI21_X1_1680_ (
  .A({ S25956[23] }),
  .B1({ S19865 }),
  .B2({ S19851 }),
  .ZN({ S19868 })
);
NAND2_X1 #() 
NAND2_X1_3242_ (
  .A1({ S19827 }),
  .A2({ S25956[22] }),
  .ZN({ S19869 })
);
OAI21_X1 #() 
OAI21_X1_1681_ (
  .A({ S19869 }),
  .B1({ S25956[22] }),
  .B2({ S19836 }),
  .ZN({ S19870 })
);
OAI211_X1 #() 
OAI211_X1_1101_ (
  .A({ S25956[124] }),
  .B({ S19868 }),
  .C1({ S19870 }),
  .C2({ S25956[23] }),
  .ZN({ S19871 })
);
NAND3_X1 #() 
NAND3_X1_3375_ (
  .A1({ S19871 }),
  .A2({ S19867 }),
  .A3({ S19814 }),
  .ZN({ S19872 })
);
NAND3_X1 #() 
NAND3_X1_3376_ (
  .A1({ S19866 }),
  .A2({ S25956[124] }),
  .A3({ S19838 }),
  .ZN({ S19873 })
);
OAI211_X1 #() 
OAI211_X1_1102_ (
  .A({ S19815 }),
  .B({ S19868 }),
  .C1({ S19870 }),
  .C2({ S25956[23] }),
  .ZN({ S19874 })
);
NAND3_X1 #() 
NAND3_X1_3377_ (
  .A1({ S19874 }),
  .A2({ S19873 }),
  .A3({ S25956[92] }),
  .ZN({ S19875 })
);
AOI21_X1 #() 
AOI21_X1_1766_ (
  .A({ S25956[60] }),
  .B1({ S19875 }),
  .B2({ S19872 }),
  .ZN({ S19876 })
);
INV_X1 #() 
INV_X1_1094_ (
  .A({ S25956[60] }),
  .ZN({ S19877 })
);
NAND3_X1 #() 
NAND3_X1_3378_ (
  .A1({ S19874 }),
  .A2({ S19873 }),
  .A3({ S19814 }),
  .ZN({ S19878 })
);
NAND3_X1 #() 
NAND3_X1_3379_ (
  .A1({ S19871 }),
  .A2({ S19867 }),
  .A3({ S25956[92] }),
  .ZN({ S19879 })
);
AOI21_X1 #() 
AOI21_X1_1767_ (
  .A({ S19877 }),
  .B1({ S19878 }),
  .B2({ S19879 }),
  .ZN({ S19880 })
);
OAI21_X1 #() 
OAI21_X1_1682_ (
  .A({ S25956[28] }),
  .B1({ S19876 }),
  .B2({ S19880 }),
  .ZN({ S19881 })
);
NAND3_X1 #() 
NAND3_X1_3380_ (
  .A1({ S19878 }),
  .A2({ S19879 }),
  .A3({ S19877 }),
  .ZN({ S19882 })
);
NAND3_X1 #() 
NAND3_X1_3381_ (
  .A1({ S19875 }),
  .A2({ S19872 }),
  .A3({ S25956[60] }),
  .ZN({ S19883 })
);
NAND3_X1 #() 
NAND3_X1_3382_ (
  .A1({ S19882 }),
  .A2({ S19883 }),
  .A3({ S18113 }),
  .ZN({ S19884 })
);
NAND2_X1 #() 
NAND2_X1_3243_ (
  .A1({ S19881 }),
  .A2({ S19884 }),
  .ZN({ S25957[1180] })
);
INV_X1 #() 
INV_X1_1095_ (
  .A({ S25956[91] }),
  .ZN({ S19885 })
);
INV_X1 #() 
INV_X1_1096_ (
  .A({ S25956[123] }),
  .ZN({ S19886 })
);
NAND2_X1 #() 
NAND2_X1_3244_ (
  .A1({ S19633 }),
  .A2({ S19718 }),
  .ZN({ S19887 })
);
OAI22_X1 #() 
OAI22_X1_88_ (
  .A1({ S19887 }),
  .A2({ S9746 }),
  .B1({ S19543 }),
  .B2({ S19792 }),
  .ZN({ S19888 })
);
NAND2_X1 #() 
NAND2_X1_3245_ (
  .A1({ S19888 }),
  .A2({ S8385 }),
  .ZN({ S19889 })
);
INV_X1 #() 
INV_X1_1097_ (
  .A({ S19599 }),
  .ZN({ S19890 })
);
INV_X1 #() 
INV_X1_1098_ (
  .A({ S19832 }),
  .ZN({ S19891 })
);
OAI211_X1 #() 
OAI211_X1_1103_ (
  .A({ S19891 }),
  .B({ S25956[20] }),
  .C1({ S19890 }),
  .C2({ S19557 }),
  .ZN({ S19892 })
);
NAND3_X1 #() 
NAND3_X1_3383_ (
  .A1({ S19889 }),
  .A2({ S25956[21] }),
  .A3({ S19892 }),
  .ZN({ S19893 })
);
OAI21_X1 #() 
OAI21_X1_1683_ (
  .A({ S19775 }),
  .B1({ S19738 }),
  .B2({ S25956[19] }),
  .ZN({ S19894 })
);
NAND2_X1 #() 
NAND2_X1_3246_ (
  .A1({ S19894 }),
  .A2({ S25956[20] }),
  .ZN({ S19895 })
);
AOI21_X1 #() 
AOI21_X1_1768_ (
  .A({ S25956[21] }),
  .B1({ S19822 }),
  .B2({ S19761 }),
  .ZN({ S19896 })
);
NAND2_X1 #() 
NAND2_X1_3247_ (
  .A1({ S19895 }),
  .A2({ S19896 }),
  .ZN({ S19897 })
);
NAND2_X1 #() 
NAND2_X1_3248_ (
  .A1({ S19897 }),
  .A2({ S19893 }),
  .ZN({ S19898 })
);
NAND2_X1 #() 
NAND2_X1_3249_ (
  .A1({ S19898 }),
  .A2({ S25956[22] }),
  .ZN({ S19899 })
);
NAND2_X1 #() 
NAND2_X1_3250_ (
  .A1({ S19593 }),
  .A2({ S25956[19] }),
  .ZN({ S19900 })
);
AOI22_X1 #() 
AOI22_X1_372_ (
  .A1({ S19761 }),
  .A2({ S9746 }),
  .B1({ S19794 }),
  .B2({ S11487 }),
  .ZN({ S19901 })
);
NAND2_X1 #() 
NAND2_X1_3251_ (
  .A1({ S19900 }),
  .A2({ S19901 }),
  .ZN({ S19902 })
);
NAND2_X1 #() 
NAND2_X1_3252_ (
  .A1({ S19902 }),
  .A2({ S8385 }),
  .ZN({ S19903 })
);
NAND2_X1 #() 
NAND2_X1_3253_ (
  .A1({ S19588 }),
  .A2({ S25956[19] }),
  .ZN({ S19904 })
);
NAND3_X1 #() 
NAND3_X1_3384_ (
  .A1({ S19904 }),
  .A2({ S25956[20] }),
  .A3({ S19852 }),
  .ZN({ S19905 })
);
AND2_X1 #() 
AND2_X1_201_ (
  .A1({ S19903 }),
  .A2({ S19905 }),
  .ZN({ S19906 })
);
NAND2_X1 #() 
NAND2_X1_3254_ (
  .A1({ S19745 }),
  .A2({ S25956[19] }),
  .ZN({ S19907 })
);
NAND2_X1 #() 
NAND2_X1_3255_ (
  .A1({ S19612 }),
  .A2({ S19701 }),
  .ZN({ S19908 })
);
NAND2_X1 #() 
NAND2_X1_3256_ (
  .A1({ S19907 }),
  .A2({ S19908 }),
  .ZN({ S19909 })
);
NAND2_X1 #() 
NAND2_X1_3257_ (
  .A1({ S19909 }),
  .A2({ S8385 }),
  .ZN({ S19910 })
);
OAI22_X1 #() 
OAI22_X1_89_ (
  .A1({ S19904 }),
  .A2({ S19553 }),
  .B1({ S19664 }),
  .B2({ S25956[19] }),
  .ZN({ S19911 })
);
OAI211_X1 #() 
OAI211_X1_1104_ (
  .A({ S19910 }),
  .B({ S25956[21] }),
  .C1({ S19911 }),
  .C2({ S8385 }),
  .ZN({ S19912 })
);
OAI211_X1 #() 
OAI211_X1_1105_ (
  .A({ S19912 }),
  .B({ S19541 }),
  .C1({ S19906 }),
  .C2({ S25956[21] }),
  .ZN({ S19913 })
);
NAND3_X1 #() 
NAND3_X1_3385_ (
  .A1({ S19913 }),
  .A2({ S19899 }),
  .A3({ S25956[23] }),
  .ZN({ S19914 })
);
NAND2_X1 #() 
NAND2_X1_3258_ (
  .A1({ S19665 }),
  .A2({ S19614 }),
  .ZN({ S19915 })
);
NAND2_X1 #() 
NAND2_X1_3259_ (
  .A1({ S19839 }),
  .A2({ S19556 }),
  .ZN({ S19916 })
);
NAND2_X1 #() 
NAND2_X1_3260_ (
  .A1({ S19646 }),
  .A2({ S19552 }),
  .ZN({ S19917 })
);
NAND2_X1 #() 
NAND2_X1_3261_ (
  .A1({ S19916 }),
  .A2({ S19917 }),
  .ZN({ S19918 })
);
OAI211_X1 #() 
OAI211_X1_1106_ (
  .A({ S19915 }),
  .B({ S25956[21] }),
  .C1({ S25956[20] }),
  .C2({ S19918 }),
  .ZN({ S19919 })
);
AOI21_X1 #() 
AOI21_X1_1769_ (
  .A({ S25956[19] }),
  .B1({ S19622 }),
  .B2({ S25956[16] }),
  .ZN({ S19920 })
);
NAND3_X1 #() 
NAND3_X1_3386_ (
  .A1({ S19584 }),
  .A2({ S9746 }),
  .A3({ S19583 }),
  .ZN({ S19921 })
);
NAND2_X1 #() 
NAND2_X1_3262_ (
  .A1({ S19921 }),
  .A2({ S8385 }),
  .ZN({ S19922 })
);
OAI221_X1 #() 
OAI221_X1_95_ (
  .A({ S7762 }),
  .B1({ S19920 }),
  .B2({ S8385 }),
  .C1({ S19922 }),
  .C2({ S19574 }),
  .ZN({ S19923 })
);
NAND3_X1 #() 
NAND3_X1_3387_ (
  .A1({ S19919 }),
  .A2({ S25956[22] }),
  .A3({ S19923 }),
  .ZN({ S19924 })
);
NAND3_X1 #() 
NAND3_X1_3388_ (
  .A1({ S19593 }),
  .A2({ S19597 }),
  .A3({ S25956[20] }),
  .ZN({ S19925 })
);
NAND3_X1 #() 
NAND3_X1_3389_ (
  .A1({ S19712 }),
  .A2({ S25956[16] }),
  .A3({ S19569 }),
  .ZN({ S19926 })
);
OAI21_X1 #() 
OAI21_X1_1684_ (
  .A({ S19925 }),
  .B1({ S25956[20] }),
  .B2({ S19926 }),
  .ZN({ S19927 })
);
AOI21_X1 #() 
AOI21_X1_1770_ (
  .A({ S9746 }),
  .B1({ S19567 }),
  .B2({ S19556 }),
  .ZN({ S19928 })
);
NOR3_X1 #() 
NOR3_X1_114_ (
  .A1({ S19928 }),
  .A2({ S19572 }),
  .A3({ S25956[20] }),
  .ZN({ S19929 })
);
NAND2_X1 #() 
NAND2_X1_3263_ (
  .A1({ S19594 }),
  .A2({ S19929 }),
  .ZN({ S19930 })
);
INV_X1 #() 
INV_X1_1099_ (
  .A({ S19715 }),
  .ZN({ S19931 })
);
NOR3_X1 #() 
NOR3_X1_115_ (
  .A1({ S19634 }),
  .A2({ S19553 }),
  .A3({ S9746 }),
  .ZN({ S19932 })
);
OAI21_X1 #() 
OAI21_X1_1685_ (
  .A({ S25956[20] }),
  .B1({ S19932 }),
  .B2({ S19931 }),
  .ZN({ S19933 })
);
NAND3_X1 #() 
NAND3_X1_3390_ (
  .A1({ S19933 }),
  .A2({ S19930 }),
  .A3({ S7762 }),
  .ZN({ S19934 })
);
OAI211_X1 #() 
OAI211_X1_1107_ (
  .A({ S19934 }),
  .B({ S19541 }),
  .C1({ S7762 }),
  .C2({ S19927 }),
  .ZN({ S19935 })
);
NAND3_X1 #() 
NAND3_X1_3391_ (
  .A1({ S19935 }),
  .A2({ S5675 }),
  .A3({ S19924 }),
  .ZN({ S19936 })
);
NAND3_X1 #() 
NAND3_X1_3392_ (
  .A1({ S19914 }),
  .A2({ S19936 }),
  .A3({ S19886 }),
  .ZN({ S19937 })
);
NAND2_X1 #() 
NAND2_X1_3264_ (
  .A1({ S19911 }),
  .A2({ S25956[20] }),
  .ZN({ S19938 })
);
OAI211_X1 #() 
OAI211_X1_1108_ (
  .A({ S19938 }),
  .B({ S25956[21] }),
  .C1({ S25956[20] }),
  .C2({ S19909 }),
  .ZN({ S19939 })
);
NAND3_X1 #() 
NAND3_X1_3393_ (
  .A1({ S19903 }),
  .A2({ S7762 }),
  .A3({ S19905 }),
  .ZN({ S19940 })
);
NAND3_X1 #() 
NAND3_X1_3394_ (
  .A1({ S19939 }),
  .A2({ S19541 }),
  .A3({ S19940 }),
  .ZN({ S19941 })
);
OAI211_X1 #() 
OAI211_X1_1109_ (
  .A({ S19941 }),
  .B({ S25956[23] }),
  .C1({ S19541 }),
  .C2({ S19898 }),
  .ZN({ S19942 })
);
NAND2_X1 #() 
NAND2_X1_3265_ (
  .A1({ S19935 }),
  .A2({ S19924 }),
  .ZN({ S19943 })
);
NAND2_X1 #() 
NAND2_X1_3266_ (
  .A1({ S19943 }),
  .A2({ S5675 }),
  .ZN({ S19944 })
);
NAND3_X1 #() 
NAND3_X1_3395_ (
  .A1({ S19942 }),
  .A2({ S19944 }),
  .A3({ S25956[123] }),
  .ZN({ S19945 })
);
NAND3_X1 #() 
NAND3_X1_3396_ (
  .A1({ S19945 }),
  .A2({ S19937 }),
  .A3({ S19885 }),
  .ZN({ S19946 })
);
NAND3_X1 #() 
NAND3_X1_3397_ (
  .A1({ S19914 }),
  .A2({ S19936 }),
  .A3({ S25956[123] }),
  .ZN({ S19947 })
);
NAND3_X1 #() 
NAND3_X1_3398_ (
  .A1({ S19942 }),
  .A2({ S19944 }),
  .A3({ S19886 }),
  .ZN({ S19948 })
);
NAND3_X1 #() 
NAND3_X1_3399_ (
  .A1({ S19948 }),
  .A2({ S19947 }),
  .A3({ S25956[91] }),
  .ZN({ S19949 })
);
AOI21_X1 #() 
AOI21_X1_1771_ (
  .A({ S25956[59] }),
  .B1({ S19946 }),
  .B2({ S19949 }),
  .ZN({ S19950 })
);
INV_X1 #() 
INV_X1_1100_ (
  .A({ S25956[59] }),
  .ZN({ S19951 })
);
NAND3_X1 #() 
NAND3_X1_3400_ (
  .A1({ S19948 }),
  .A2({ S19947 }),
  .A3({ S19885 }),
  .ZN({ S19952 })
);
NAND3_X1 #() 
NAND3_X1_3401_ (
  .A1({ S19945 }),
  .A2({ S19937 }),
  .A3({ S25956[91] }),
  .ZN({ S19953 })
);
AOI21_X1 #() 
AOI21_X1_1772_ (
  .A({ S19951 }),
  .B1({ S19952 }),
  .B2({ S19953 }),
  .ZN({ S19954 })
);
OAI21_X1 #() 
OAI21_X1_1686_ (
  .A({ S18124 }),
  .B1({ S19950 }),
  .B2({ S19954 }),
  .ZN({ S19955 })
);
NAND3_X1 #() 
NAND3_X1_3402_ (
  .A1({ S19952 }),
  .A2({ S19953 }),
  .A3({ S19951 }),
  .ZN({ S19956 })
);
NAND3_X1 #() 
NAND3_X1_3403_ (
  .A1({ S19946 }),
  .A2({ S19949 }),
  .A3({ S25956[59] }),
  .ZN({ S19957 })
);
NAND3_X1 #() 
NAND3_X1_3404_ (
  .A1({ S19956 }),
  .A2({ S19957 }),
  .A3({ S25956[27] }),
  .ZN({ S19958 })
);
NAND2_X1 #() 
NAND2_X1_3267_ (
  .A1({ S19955 }),
  .A2({ S19958 }),
  .ZN({ S71 })
);
OAI21_X1 #() 
OAI21_X1_1687_ (
  .A({ S25956[27] }),
  .B1({ S19950 }),
  .B2({ S19954 }),
  .ZN({ S19959 })
);
NAND3_X1 #() 
NAND3_X1_3405_ (
  .A1({ S19956 }),
  .A2({ S19957 }),
  .A3({ S18124 }),
  .ZN({ S19960 })
);
NAND2_X1 #() 
NAND2_X1_3268_ (
  .A1({ S19959 }),
  .A2({ S19960 }),
  .ZN({ S25957[1179] })
);
INV_X1 #() 
INV_X1_1101_ (
  .A({ S25956[120] }),
  .ZN({ S19961 })
);
OAI21_X1 #() 
OAI21_X1_1688_ (
  .A({ S25956[19] }),
  .B1({ S19782 }),
  .B2({ S19561 }),
  .ZN({ S19962 })
);
AOI21_X1 #() 
AOI21_X1_1773_ (
  .A({ S8385 }),
  .B1({ S19751 }),
  .B2({ S19667 }),
  .ZN({ S19963 })
);
AOI22_X1 #() 
AOI22_X1_373_ (
  .A1({ S19962 }),
  .A2({ S19963 }),
  .B1({ S19720 }),
  .B2({ S19645 }),
  .ZN({ S19964 })
);
NAND3_X1 #() 
NAND3_X1_3406_ (
  .A1({ S19764 }),
  .A2({ S8385 }),
  .A3({ S19774 }),
  .ZN({ S19965 })
);
NAND4_X1 #() 
NAND4_X1_357_ (
  .A1({ S19683 }),
  .A2({ S19750 }),
  .A3({ S19544 }),
  .A4({ S25956[20] }),
  .ZN({ S19966 })
);
NAND3_X1 #() 
NAND3_X1_3407_ (
  .A1({ S19965 }),
  .A2({ S7762 }),
  .A3({ S19966 }),
  .ZN({ S19967 })
);
OAI21_X1 #() 
OAI21_X1_1689_ (
  .A({ S19967 }),
  .B1({ S7762 }),
  .B2({ S19964 }),
  .ZN({ S19968 })
);
OAI22_X1 #() 
OAI22_X1_90_ (
  .A1({ S19705 }),
  .A2({ S19570 }),
  .B1({ S9746 }),
  .B2({ S19690 }),
  .ZN({ S19969 })
);
NAND2_X1 #() 
NAND2_X1_3269_ (
  .A1({ S19549 }),
  .A2({ S9746 }),
  .ZN({ S19970 })
);
NAND4_X1 #() 
NAND4_X1_358_ (
  .A1({ S19610 }),
  .A2({ S19904 }),
  .A3({ S25956[20] }),
  .A4({ S19970 }),
  .ZN({ S19971 })
);
OAI211_X1 #() 
OAI211_X1_1110_ (
  .A({ S19971 }),
  .B({ S7762 }),
  .C1({ S25956[20] }),
  .C2({ S19969 }),
  .ZN({ S19972 })
);
NAND3_X1 #() 
NAND3_X1_3408_ (
  .A1({ S19752 }),
  .A2({ S19891 }),
  .A3({ S25956[20] }),
  .ZN({ S19973 })
);
NAND3_X1 #() 
NAND3_X1_3409_ (
  .A1({ S19670 }),
  .A2({ S19740 }),
  .A3({ S8385 }),
  .ZN({ S19974 })
);
NAND3_X1 #() 
NAND3_X1_3410_ (
  .A1({ S19973 }),
  .A2({ S19974 }),
  .A3({ S25956[21] }),
  .ZN({ S19975 })
);
NAND3_X1 #() 
NAND3_X1_3411_ (
  .A1({ S19972 }),
  .A2({ S19541 }),
  .A3({ S19975 }),
  .ZN({ S19976 })
);
OAI211_X1 #() 
OAI211_X1_1111_ (
  .A({ S19976 }),
  .B({ S5675 }),
  .C1({ S19541 }),
  .C2({ S19968 }),
  .ZN({ S19977 })
);
NAND2_X1 #() 
NAND2_X1_3270_ (
  .A1({ S19542 }),
  .A2({ S25956[18] }),
  .ZN({ S19978 })
);
NOR2_X1 #() 
NOR2_X1_842_ (
  .A1({ S19978 }),
  .A2({ S9746 }),
  .ZN({ S19979 })
);
OAI21_X1 #() 
OAI21_X1_1690_ (
  .A({ S25956[21] }),
  .B1({ S19831 }),
  .B2({ S19979 }),
  .ZN({ S19980 })
);
NAND3_X1 #() 
NAND3_X1_3412_ (
  .A1({ S19887 }),
  .A2({ S7762 }),
  .A3({ S9746 }),
  .ZN({ S19981 })
);
AND3_X1 #() 
AND3_X1_127_ (
  .A1({ S19981 }),
  .A2({ S19900 }),
  .A3({ S25956[20] }),
  .ZN({ S19982 })
);
NOR2_X1 #() 
NOR2_X1_843_ (
  .A1({ S19634 }),
  .A2({ S19598 }),
  .ZN({ S19983 })
);
NOR3_X1 #() 
NOR3_X1_116_ (
  .A1({ S19574 }),
  .A2({ S19983 }),
  .A3({ S7762 }),
  .ZN({ S19984 })
);
OAI211_X1 #() 
OAI211_X1_1112_ (
  .A({ S7762 }),
  .B({ S19743 }),
  .C1({ S19697 }),
  .C2({ S9746 }),
  .ZN({ S19985 })
);
NAND2_X1 #() 
NAND2_X1_3271_ (
  .A1({ S19985 }),
  .A2({ S8385 }),
  .ZN({ S19986 })
);
NOR2_X1 #() 
NOR2_X1_844_ (
  .A1({ S19986 }),
  .A2({ S19984 }),
  .ZN({ S19987 })
);
AOI21_X1 #() 
AOI21_X1_1774_ (
  .A({ S19987 }),
  .B1({ S19982 }),
  .B2({ S19980 }),
  .ZN({ S19988 })
);
AOI21_X1 #() 
AOI21_X1_1775_ (
  .A({ S25956[20] }),
  .B1({ S19845 }),
  .B2({ S19564 }),
  .ZN({ S19989 })
);
NAND2_X1 #() 
NAND2_X1_3272_ (
  .A1({ S19714 }),
  .A2({ S19559 }),
  .ZN({ S19990 })
);
NAND2_X1 #() 
NAND2_X1_3273_ (
  .A1({ S19990 }),
  .A2({ S9746 }),
  .ZN({ S19991 })
);
NAND2_X1 #() 
NAND2_X1_3274_ (
  .A1({ S19991 }),
  .A2({ S19597 }),
  .ZN({ S19992 })
);
AOI21_X1 #() 
AOI21_X1_1776_ (
  .A({ S19989 }),
  .B1({ S25956[20] }),
  .B2({ S19992 }),
  .ZN({ S19993 })
);
AOI21_X1 #() 
AOI21_X1_1777_ (
  .A({ S19688 }),
  .B1({ S19634 }),
  .B2({ S9746 }),
  .ZN({ S19994 })
);
OAI21_X1 #() 
OAI21_X1_1691_ (
  .A({ S9746 }),
  .B1({ S19676 }),
  .B2({ S19668 }),
  .ZN({ S19995 })
);
AOI21_X1 #() 
AOI21_X1_1778_ (
  .A({ S25956[20] }),
  .B1({ S19995 }),
  .B2({ S19917 }),
  .ZN({ S19996 })
);
OAI21_X1 #() 
OAI21_X1_1692_ (
  .A({ S7762 }),
  .B1({ S19994 }),
  .B2({ S19996 }),
  .ZN({ S19997 })
);
OAI211_X1 #() 
OAI211_X1_1113_ (
  .A({ S19541 }),
  .B({ S19997 }),
  .C1({ S19993 }),
  .C2({ S7762 }),
  .ZN({ S19998 })
);
OAI211_X1 #() 
OAI211_X1_1114_ (
  .A({ S19998 }),
  .B({ S25956[23] }),
  .C1({ S19988 }),
  .C2({ S19541 }),
  .ZN({ S19999 })
);
NAND3_X1 #() 
NAND3_X1_3413_ (
  .A1({ S19999 }),
  .A2({ S19961 }),
  .A3({ S19977 }),
  .ZN({ S20000 })
);
AND2_X1 #() 
AND2_X1_202_ (
  .A1({ S19972 }),
  .A2({ S19975 }),
  .ZN({ S20001 })
);
NAND2_X1 #() 
NAND2_X1_3275_ (
  .A1({ S19968 }),
  .A2({ S25956[22] }),
  .ZN({ S20002 })
);
OAI211_X1 #() 
OAI211_X1_1115_ (
  .A({ S20002 }),
  .B({ S5675 }),
  .C1({ S20001 }),
  .C2({ S25956[22] }),
  .ZN({ S20003 })
);
OAI21_X1 #() 
OAI21_X1_1693_ (
  .A({ S19997 }),
  .B1({ S19993 }),
  .B2({ S7762 }),
  .ZN({ S20004 })
);
NAND2_X1 #() 
NAND2_X1_3276_ (
  .A1({ S20004 }),
  .A2({ S19541 }),
  .ZN({ S20005 })
);
NAND4_X1 #() 
NAND4_X1_359_ (
  .A1({ S19980 }),
  .A2({ S19981 }),
  .A3({ S25956[20] }),
  .A4({ S19900 }),
  .ZN({ S20006 })
);
OAI211_X1 #() 
OAI211_X1_1116_ (
  .A({ S20006 }),
  .B({ S25956[22] }),
  .C1({ S19984 }),
  .C2({ S19986 }),
  .ZN({ S20007 })
);
NAND3_X1 #() 
NAND3_X1_3414_ (
  .A1({ S20005 }),
  .A2({ S25956[23] }),
  .A3({ S20007 }),
  .ZN({ S20008 })
);
NAND3_X1 #() 
NAND3_X1_3415_ (
  .A1({ S20003 }),
  .A2({ S25956[120] }),
  .A3({ S20008 }),
  .ZN({ S20009 })
);
AOI21_X1 #() 
AOI21_X1_1779_ (
  .A({ S25956[88] }),
  .B1({ S20009 }),
  .B2({ S20000 }),
  .ZN({ S20010 })
);
INV_X1 #() 
INV_X1_1102_ (
  .A({ S25956[88] }),
  .ZN({ S20011 })
);
NAND3_X1 #() 
NAND3_X1_3416_ (
  .A1({ S19999 }),
  .A2({ S25956[120] }),
  .A3({ S19977 }),
  .ZN({ S20012 })
);
NAND3_X1 #() 
NAND3_X1_3417_ (
  .A1({ S20003 }),
  .A2({ S19961 }),
  .A3({ S20008 }),
  .ZN({ S20013 })
);
AOI21_X1 #() 
AOI21_X1_1780_ (
  .A({ S20011 }),
  .B1({ S20013 }),
  .B2({ S20012 }),
  .ZN({ S20014 })
);
OAI21_X1 #() 
OAI21_X1_1694_ (
  .A({ S25956[56] }),
  .B1({ S20010 }),
  .B2({ S20014 }),
  .ZN({ S20015 })
);
INV_X1 #() 
INV_X1_1103_ (
  .A({ S25956[56] }),
  .ZN({ S20016 })
);
NAND3_X1 #() 
NAND3_X1_3418_ (
  .A1({ S20013 }),
  .A2({ S20012 }),
  .A3({ S20011 }),
  .ZN({ S20017 })
);
NAND3_X1 #() 
NAND3_X1_3419_ (
  .A1({ S20009 }),
  .A2({ S20000 }),
  .A3({ S25956[88] }),
  .ZN({ S20018 })
);
NAND3_X1 #() 
NAND3_X1_3420_ (
  .A1({ S20017 }),
  .A2({ S20018 }),
  .A3({ S20016 }),
  .ZN({ S20019 })
);
NAND3_X1 #() 
NAND3_X1_3421_ (
  .A1({ S20015 }),
  .A2({ S25956[24] }),
  .A3({ S20019 }),
  .ZN({ S20020 })
);
OAI21_X1 #() 
OAI21_X1_1695_ (
  .A({ S20016 }),
  .B1({ S20010 }),
  .B2({ S20014 }),
  .ZN({ S20021 })
);
NAND3_X1 #() 
NAND3_X1_3422_ (
  .A1({ S20017 }),
  .A2({ S20018 }),
  .A3({ S25956[56] }),
  .ZN({ S20022 })
);
NAND3_X1 #() 
NAND3_X1_3423_ (
  .A1({ S20021 }),
  .A2({ S18242 }),
  .A3({ S20022 }),
  .ZN({ S20023 })
);
NAND2_X1 #() 
NAND2_X1_3277_ (
  .A1({ S20020 }),
  .A2({ S20023 }),
  .ZN({ S25957[1176] })
);
INV_X1 #() 
INV_X1_1104_ (
  .A({ S25956[57] }),
  .ZN({ S20024 })
);
INV_X1 #() 
INV_X1_1105_ (
  .A({ S25956[89] }),
  .ZN({ S20025 })
);
NAND3_X1 #() 
NAND3_X1_3424_ (
  .A1({ S19783 }),
  .A2({ S19551 }),
  .A3({ S19630 }),
  .ZN({ S20026 })
);
OAI21_X1 #() 
OAI21_X1_1696_ (
  .A({ S25956[20] }),
  .B1({ S19710 }),
  .B2({ S19642 }),
  .ZN({ S20027 })
);
OAI221_X1 #() 
OAI221_X1_96_ (
  .A({ S25956[21] }),
  .B1({ S25956[20] }),
  .B2({ S20026 }),
  .C1({ S19932 }),
  .C2({ S20027 }),
  .ZN({ S20028 })
);
NAND2_X1 #() 
NAND2_X1_3278_ (
  .A1({ S19697 }),
  .A2({ S9746 }),
  .ZN({ S20029 })
);
NAND3_X1 #() 
NAND3_X1_3425_ (
  .A1({ S20029 }),
  .A2({ S19900 }),
  .A3({ S8385 }),
  .ZN({ S20030 })
);
OAI21_X1 #() 
OAI21_X1_1697_ (
  .A({ S9746 }),
  .B1({ S19602 }),
  .B2({ S19788 }),
  .ZN({ S20031 })
);
NAND3_X1 #() 
NAND3_X1_3426_ (
  .A1({ S19962 }),
  .A2({ S25956[20] }),
  .A3({ S20031 }),
  .ZN({ S20032 })
);
NAND3_X1 #() 
NAND3_X1_3427_ (
  .A1({ S20030 }),
  .A2({ S7762 }),
  .A3({ S20032 }),
  .ZN({ S20033 })
);
NAND3_X1 #() 
NAND3_X1_3428_ (
  .A1({ S20033 }),
  .A2({ S20028 }),
  .A3({ S25956[22] }),
  .ZN({ S20034 })
);
AOI21_X1 #() 
AOI21_X1_1781_ (
  .A({ S8385 }),
  .B1({ S19907 }),
  .B2({ S19840 }),
  .ZN({ S20035 })
);
OAI21_X1 #() 
OAI21_X1_1698_ (
  .A({ S25956[21] }),
  .B1({ S20035 }),
  .B2({ S19586 }),
  .ZN({ S20036 })
);
NAND2_X1 #() 
NAND2_X1_3279_ (
  .A1({ S19852 }),
  .A2({ S25956[20] }),
  .ZN({ S20037 })
);
OAI211_X1 #() 
OAI211_X1_1117_ (
  .A({ S19921 }),
  .B({ S8385 }),
  .C1({ S25956[18] }),
  .C2({ S19630 }),
  .ZN({ S20038 })
);
OAI211_X1 #() 
OAI211_X1_1118_ (
  .A({ S20038 }),
  .B({ S7762 }),
  .C1({ S19631 }),
  .C2({ S20037 }),
  .ZN({ S20039 })
);
NAND3_X1 #() 
NAND3_X1_3429_ (
  .A1({ S20036 }),
  .A2({ S19541 }),
  .A3({ S20039 }),
  .ZN({ S20040 })
);
NAND3_X1 #() 
NAND3_X1_3430_ (
  .A1({ S20040 }),
  .A2({ S20034 }),
  .A3({ S5675 }),
  .ZN({ S20041 })
);
OAI221_X1 #() 
OAI221_X1_97_ (
  .A({ S19970 }),
  .B1({ S9746 }),
  .B2({ S19569 }),
  .C1({ S19568 }),
  .C2({ S10926 }),
  .ZN({ S20042 })
);
OAI22_X1 #() 
OAI22_X1_91_ (
  .A1({ S19858 }),
  .A2({ S19589 }),
  .B1({ S8385 }),
  .B2({ S20042 }),
  .ZN({ S20043 })
);
OAI21_X1 #() 
OAI21_X1_1699_ (
  .A({ S19916 }),
  .B1({ S9746 }),
  .B2({ S19771 }),
  .ZN({ S20044 })
);
NAND3_X1 #() 
NAND3_X1_3431_ (
  .A1({ S19559 }),
  .A2({ S25956[19] }),
  .A3({ S19689 }),
  .ZN({ S20045 })
);
AOI21_X1 #() 
AOI21_X1_1782_ (
  .A({ S7762 }),
  .B1({ S19600 }),
  .B2({ S20045 }),
  .ZN({ S20046 })
);
OAI21_X1 #() 
OAI21_X1_1700_ (
  .A({ S20046 }),
  .B1({ S25956[20] }),
  .B2({ S20044 }),
  .ZN({ S20047 })
);
OAI211_X1 #() 
OAI211_X1_1119_ (
  .A({ S19541 }),
  .B({ S20047 }),
  .C1({ S20043 }),
  .C2({ S25956[21] }),
  .ZN({ S20048 })
);
OAI21_X1 #() 
OAI21_X1_1701_ (
  .A({ S19775 }),
  .B1({ S19602 }),
  .B2({ S25956[19] }),
  .ZN({ S20049 })
);
NAND3_X1 #() 
NAND3_X1_3432_ (
  .A1({ S19962 }),
  .A2({ S8385 }),
  .A3({ S19890 }),
  .ZN({ S20050 })
);
OAI21_X1 #() 
OAI21_X1_1702_ (
  .A({ S20050 }),
  .B1({ S8385 }),
  .B2({ S20049 }),
  .ZN({ S20051 })
);
OAI221_X1 #() 
OAI221_X1_98_ (
  .A({ S25956[20] }),
  .B1({ S19598 }),
  .B2({ S25956[16] }),
  .C1({ S19745 }),
  .C2({ S19597 }),
  .ZN({ S20052 })
);
AOI21_X1 #() 
AOI21_X1_1783_ (
  .A({ S19928 }),
  .B1({ S19920 }),
  .B2({ S19783 }),
  .ZN({ S20053 })
);
NAND2_X1 #() 
NAND2_X1_3280_ (
  .A1({ S20053 }),
  .A2({ S8385 }),
  .ZN({ S20054 })
);
NAND3_X1 #() 
NAND3_X1_3433_ (
  .A1({ S20052 }),
  .A2({ S20054 }),
  .A3({ S7762 }),
  .ZN({ S20055 })
);
OAI211_X1 #() 
OAI211_X1_1120_ (
  .A({ S20055 }),
  .B({ S25956[22] }),
  .C1({ S20051 }),
  .C2({ S7762 }),
  .ZN({ S20056 })
);
NAND3_X1 #() 
NAND3_X1_3434_ (
  .A1({ S20056 }),
  .A2({ S20048 }),
  .A3({ S25956[23] }),
  .ZN({ S20057 })
);
NAND3_X1 #() 
NAND3_X1_3435_ (
  .A1({ S20057 }),
  .A2({ S20041 }),
  .A3({ S25956[121] }),
  .ZN({ S20058 })
);
INV_X1 #() 
INV_X1_1106_ (
  .A({ S25956[121] }),
  .ZN({ S20059 })
);
NAND2_X1 #() 
NAND2_X1_3281_ (
  .A1({ S20057 }),
  .A2({ S20041 }),
  .ZN({ S20060 })
);
NAND2_X1 #() 
NAND2_X1_3282_ (
  .A1({ S20060 }),
  .A2({ S20059 }),
  .ZN({ S20061 })
);
NAND3_X1 #() 
NAND3_X1_3436_ (
  .A1({ S20061 }),
  .A2({ S20025 }),
  .A3({ S20058 }),
  .ZN({ S20062 })
);
NAND3_X1 #() 
NAND3_X1_3437_ (
  .A1({ S20057 }),
  .A2({ S20041 }),
  .A3({ S20059 }),
  .ZN({ S20063 })
);
NAND2_X1 #() 
NAND2_X1_3283_ (
  .A1({ S20060 }),
  .A2({ S25956[121] }),
  .ZN({ S20064 })
);
NAND3_X1 #() 
NAND3_X1_3438_ (
  .A1({ S20064 }),
  .A2({ S25956[89] }),
  .A3({ S20063 }),
  .ZN({ S20065 })
);
AND3_X1 #() 
AND3_X1_128_ (
  .A1({ S20065 }),
  .A2({ S20062 }),
  .A3({ S20024 }),
  .ZN({ S20066 })
);
AOI21_X1 #() 
AOI21_X1_1784_ (
  .A({ S20024 }),
  .B1({ S20062 }),
  .B2({ S20065 }),
  .ZN({ S20067 })
);
OAI21_X1 #() 
OAI21_X1_1703_ (
  .A({ S25956[25] }),
  .B1({ S20066 }),
  .B2({ S20067 }),
  .ZN({ S20068 })
);
NAND3_X1 #() 
NAND3_X1_3439_ (
  .A1({ S20062 }),
  .A2({ S20065 }),
  .A3({ S20024 }),
  .ZN({ S20069 })
);
NAND2_X1 #() 
NAND2_X1_3284_ (
  .A1({ S20062 }),
  .A2({ S20065 }),
  .ZN({ S25957[1241] })
);
NAND2_X1 #() 
NAND2_X1_3285_ (
  .A1({ S25957[1241] }),
  .A2({ S25956[57] }),
  .ZN({ S20070 })
);
NAND3_X1 #() 
NAND3_X1_3440_ (
  .A1({ S20070 }),
  .A2({ S18383 }),
  .A3({ S20069 }),
  .ZN({ S20071 })
);
NAND2_X1 #() 
NAND2_X1_3286_ (
  .A1({ S20068 }),
  .A2({ S20071 }),
  .ZN({ S25957[1177] })
);
INV_X1 #() 
INV_X1_1107_ (
  .A({ S25956[90] }),
  .ZN({ S20072 })
);
INV_X1 #() 
INV_X1_1108_ (
  .A({ S25956[122] }),
  .ZN({ S20073 })
);
NOR3_X1 #() 
NOR3_X1_117_ (
  .A1({ S19557 }),
  .A2({ S19549 }),
  .A3({ S9746 }),
  .ZN({ S20074 })
);
OAI21_X1 #() 
OAI21_X1_1704_ (
  .A({ S25956[20] }),
  .B1({ S20074 }),
  .B2({ S19920 }),
  .ZN({ S20075 })
);
INV_X1 #() 
INV_X1_1109_ (
  .A({ S19839 }),
  .ZN({ S20076 })
);
OAI21_X1 #() 
OAI21_X1_1705_ (
  .A({ S8385 }),
  .B1({ S20076 }),
  .B2({ S10390 }),
  .ZN({ S20077 })
);
OAI211_X1 #() 
OAI211_X1_1121_ (
  .A({ S20075 }),
  .B({ S25956[21] }),
  .C1({ S20077 }),
  .C2({ S19640 }),
  .ZN({ S20078 })
);
OAI22_X1 #() 
OAI22_X1_92_ (
  .A1({ S19762 }),
  .A2({ S9746 }),
  .B1({ S19702 }),
  .B2({ S19689 }),
  .ZN({ S20079 })
);
NAND3_X1 #() 
NAND3_X1_3441_ (
  .A1({ S19641 }),
  .A2({ S25956[19] }),
  .A3({ S25956[17] }),
  .ZN({ S20080 })
);
OAI211_X1 #() 
OAI211_X1_1122_ (
  .A({ S20080 }),
  .B({ S8385 }),
  .C1({ S19887 }),
  .C2({ S25956[19] }),
  .ZN({ S20081 })
);
OAI211_X1 #() 
OAI211_X1_1123_ (
  .A({ S20081 }),
  .B({ S7762 }),
  .C1({ S20079 }),
  .C2({ S8385 }),
  .ZN({ S20082 })
);
AOI21_X1 #() 
AOI21_X1_1785_ (
  .A({ S19541 }),
  .B1({ S20078 }),
  .B2({ S20082 }),
  .ZN({ S20083 })
);
NAND2_X1 #() 
NAND2_X1_3287_ (
  .A1({ S19861 }),
  .A2({ S20080 }),
  .ZN({ S20084 })
);
OAI22_X1 #() 
OAI22_X1_93_ (
  .A1({ S19721 }),
  .A2({ S19983 }),
  .B1({ S20084 }),
  .B2({ S8385 }),
  .ZN({ S20085 })
);
NAND2_X1 #() 
NAND2_X1_3288_ (
  .A1({ S19759 }),
  .A2({ S25956[19] }),
  .ZN({ S20086 })
);
NAND3_X1 #() 
NAND3_X1_3442_ (
  .A1({ S20086 }),
  .A2({ S8385 }),
  .A3({ S19743 }),
  .ZN({ S20087 })
);
OAI211_X1 #() 
OAI211_X1_1124_ (
  .A({ S19908 }),
  .B({ S25956[20] }),
  .C1({ S19784 }),
  .C2({ S19580 }),
  .ZN({ S20088 })
);
NAND3_X1 #() 
NAND3_X1_3443_ (
  .A1({ S20087 }),
  .A2({ S25956[21] }),
  .A3({ S20088 }),
  .ZN({ S20089 })
);
OAI21_X1 #() 
OAI21_X1_1706_ (
  .A({ S20089 }),
  .B1({ S25956[21] }),
  .B2({ S20085 }),
  .ZN({ S20090 })
);
OAI21_X1 #() 
OAI21_X1_1707_ (
  .A({ S5675 }),
  .B1({ S20090 }),
  .B2({ S25956[22] }),
  .ZN({ S20091 })
);
AOI22_X1 #() 
AOI22_X1_374_ (
  .A1({ S19546 }),
  .A2({ S19761 }),
  .B1({ S19553 }),
  .B2({ S9746 }),
  .ZN({ S20092 })
);
OAI211_X1 #() 
OAI211_X1_1125_ (
  .A({ S19921 }),
  .B({ S25956[20] }),
  .C1({ S10390 }),
  .C2({ S19638 }),
  .ZN({ S20093 })
);
OAI21_X1 #() 
OAI21_X1_1708_ (
  .A({ S20093 }),
  .B1({ S25956[20] }),
  .B2({ S20092 }),
  .ZN({ S20094 })
);
NAND3_X1 #() 
NAND3_X1_3444_ (
  .A1({ S19743 }),
  .A2({ S19687 }),
  .A3({ S8385 }),
  .ZN({ S20095 })
);
NAND3_X1 #() 
NAND3_X1_3445_ (
  .A1({ S20076 }),
  .A2({ S25956[20] }),
  .A3({ S20080 }),
  .ZN({ S20096 })
);
NAND3_X1 #() 
NAND3_X1_3446_ (
  .A1({ S20096 }),
  .A2({ S7762 }),
  .A3({ S20095 }),
  .ZN({ S20097 })
);
OAI211_X1 #() 
OAI211_X1_1126_ (
  .A({ S19541 }),
  .B({ S20097 }),
  .C1({ S20094 }),
  .C2({ S7762 }),
  .ZN({ S20098 })
);
OAI21_X1 #() 
OAI21_X1_1709_ (
  .A({ S9746 }),
  .B1({ S19634 }),
  .B2({ S19558 }),
  .ZN({ S20099 })
);
NAND3_X1 #() 
NAND3_X1_3447_ (
  .A1({ S20099 }),
  .A2({ S25956[20] }),
  .A3({ S19582 }),
  .ZN({ S20100 })
);
NAND3_X1 #() 
NAND3_X1_3448_ (
  .A1({ S19635 }),
  .A2({ S25956[19] }),
  .A3({ S19978 }),
  .ZN({ S20101 })
);
NAND3_X1 #() 
NAND3_X1_3449_ (
  .A1({ S20101 }),
  .A2({ S8385 }),
  .A3({ S19598 }),
  .ZN({ S20102 })
);
NAND3_X1 #() 
NAND3_X1_3450_ (
  .A1({ S20102 }),
  .A2({ S20100 }),
  .A3({ S25956[21] }),
  .ZN({ S20103 })
);
OAI211_X1 #() 
OAI211_X1_1127_ (
  .A({ S25956[20] }),
  .B({ S19787 }),
  .C1({ S19636 }),
  .C2({ S9746 }),
  .ZN({ S20104 })
);
NAND3_X1 #() 
NAND3_X1_3451_ (
  .A1({ S19620 }),
  .A2({ S8385 }),
  .A3({ S19970 }),
  .ZN({ S20105 })
);
NAND3_X1 #() 
NAND3_X1_3452_ (
  .A1({ S20104 }),
  .A2({ S7762 }),
  .A3({ S20105 }),
  .ZN({ S20106 })
);
NAND3_X1 #() 
NAND3_X1_3453_ (
  .A1({ S20106 }),
  .A2({ S20103 }),
  .A3({ S25956[22] }),
  .ZN({ S20107 })
);
NAND3_X1 #() 
NAND3_X1_3454_ (
  .A1({ S20107 }),
  .A2({ S20098 }),
  .A3({ S25956[23] }),
  .ZN({ S20108 })
);
OAI211_X1 #() 
OAI211_X1_1128_ (
  .A({ S20073 }),
  .B({ S20108 }),
  .C1({ S20091 }),
  .C2({ S20083 }),
  .ZN({ S20109 })
);
OAI21_X1 #() 
OAI21_X1_1710_ (
  .A({ S20108 }),
  .B1({ S20091 }),
  .B2({ S20083 }),
  .ZN({ S20110 })
);
NAND2_X1 #() 
NAND2_X1_3289_ (
  .A1({ S20110 }),
  .A2({ S25956[122] }),
  .ZN({ S20111 })
);
NAND3_X1 #() 
NAND3_X1_3455_ (
  .A1({ S20111 }),
  .A2({ S20072 }),
  .A3({ S20109 }),
  .ZN({ S20112 })
);
OAI211_X1 #() 
OAI211_X1_1129_ (
  .A({ S25956[122] }),
  .B({ S20108 }),
  .C1({ S20091 }),
  .C2({ S20083 }),
  .ZN({ S20113 })
);
NAND2_X1 #() 
NAND2_X1_3290_ (
  .A1({ S20110 }),
  .A2({ S20073 }),
  .ZN({ S20114 })
);
NAND3_X1 #() 
NAND3_X1_3456_ (
  .A1({ S20114 }),
  .A2({ S25956[90] }),
  .A3({ S20113 }),
  .ZN({ S20115 })
);
AOI21_X1 #() 
AOI21_X1_1786_ (
  .A({ S25956[58] }),
  .B1({ S20112 }),
  .B2({ S20115 }),
  .ZN({ S20116 })
);
INV_X1 #() 
INV_X1_1110_ (
  .A({ S25956[58] }),
  .ZN({ S20117 })
);
NAND3_X1 #() 
NAND3_X1_3457_ (
  .A1({ S20114 }),
  .A2({ S20072 }),
  .A3({ S20113 }),
  .ZN({ S20118 })
);
NAND3_X1 #() 
NAND3_X1_3458_ (
  .A1({ S20111 }),
  .A2({ S25956[90] }),
  .A3({ S20109 }),
  .ZN({ S20119 })
);
AOI21_X1 #() 
AOI21_X1_1787_ (
  .A({ S20117 }),
  .B1({ S20118 }),
  .B2({ S20119 }),
  .ZN({ S20120 })
);
OAI21_X1 #() 
OAI21_X1_1711_ (
  .A({ S25956[26] }),
  .B1({ S20116 }),
  .B2({ S20120 }),
  .ZN({ S20121 })
);
NAND3_X1 #() 
NAND3_X1_3459_ (
  .A1({ S20118 }),
  .A2({ S20119 }),
  .A3({ S20117 }),
  .ZN({ S20122 })
);
NAND3_X1 #() 
NAND3_X1_3460_ (
  .A1({ S20112 }),
  .A2({ S20115 }),
  .A3({ S25956[58] }),
  .ZN({ S20123 })
);
NAND3_X1 #() 
NAND3_X1_3461_ (
  .A1({ S20122 }),
  .A2({ S20123 }),
  .A3({ S18198 }),
  .ZN({ S20124 })
);
NAND2_X1 #() 
NAND2_X1_3291_ (
  .A1({ S20121 }),
  .A2({ S20124 }),
  .ZN({ S25957[1178] })
);
OAI21_X1 #() 
OAI21_X1_1712_ (
  .A({ S5639 }),
  .B1({ S16516 }),
  .B2({ S16560 }),
  .ZN({ S20125 })
);
NAND3_X1 #() 
NAND3_X1_3462_ (
  .A1({ S16582 }),
  .A2({ S16592 }),
  .A3({ S25956[8] }),
  .ZN({ S20126 })
);
OAI21_X1 #() 
OAI21_X1_1713_ (
  .A({ S5628 }),
  .B1({ S17241 }),
  .B2({ S17284 }),
  .ZN({ S20127 })
);
NAND3_X1 #() 
NAND3_X1_3463_ (
  .A1({ S17306 }),
  .A2({ S17317 }),
  .A3({ S25956[9] }),
  .ZN({ S20128 })
);
NAND4_X1 #() 
NAND4_X1_360_ (
  .A1({ S20125 }),
  .A2({ S20127 }),
  .A3({ S20126 }),
  .A4({ S20128 }),
  .ZN({ S20129 })
);
INV_X1 #() 
INV_X1_1111_ (
  .A({ S20129 }),
  .ZN({ S72 })
);
NAND4_X1 #() 
NAND4_X1_361_ (
  .A1({ S16571 }),
  .A2({ S17295 }),
  .A3({ S16603 }),
  .A4({ S17328 }),
  .ZN({ S73 })
);
INV_X1 #() 
INV_X1_1112_ (
  .A({ S6989 }),
  .ZN({ S25957[1239] })
);
AND2_X1 #() 
AND2_X1_203_ (
  .A1({ S13691 }),
  .A2({ S13723 }),
  .ZN({ S20130 })
);
AND2_X1 #() 
AND2_X1_204_ (
  .A1({ S15250 }),
  .A2({ S15283 }),
  .ZN({ S20131 })
);
NAND4_X1 #() 
NAND4_X1_362_ (
  .A1({ S16571 }),
  .A2({ S16603 }),
  .A3({ S17987 }),
  .A4({ S18019 }),
  .ZN({ S20132 })
);
INV_X1 #() 
INV_X1_1113_ (
  .A({ S20132 }),
  .ZN({ S20133 })
);
NAND3_X1 #() 
NAND3_X1_3464_ (
  .A1({ S17998 }),
  .A2({ S18008 }),
  .A3({ S25956[10] }),
  .ZN({ S20134 })
);
NAND3_X1 #() 
NAND3_X1_3465_ (
  .A1({ S17944 }),
  .A2({ S17976 }),
  .A3({ S5730 }),
  .ZN({ S20135 })
);
NAND4_X1 #() 
NAND4_X1_363_ (
  .A1({ S16571 }),
  .A2({ S16603 }),
  .A3({ S20134 }),
  .A4({ S20135 }),
  .ZN({ S20136 })
);
NAND2_X1 #() 
NAND2_X1_3292_ (
  .A1({ S20127 }),
  .A2({ S20128 }),
  .ZN({ S20137 })
);
NAND2_X1 #() 
NAND2_X1_3293_ (
  .A1({ S20134 }),
  .A2({ S20135 }),
  .ZN({ S20138 })
);
NAND3_X1 #() 
NAND3_X1_3466_ (
  .A1({ S25957[1160] }),
  .A2({ S20137 }),
  .A3({ S20138 }),
  .ZN({ S20139 })
);
NAND3_X1 #() 
NAND3_X1_3467_ (
  .A1({ S20139 }),
  .A2({ S25957[1163] }),
  .A3({ S20136 }),
  .ZN({ S20140 })
);
NAND2_X1 #() 
NAND2_X1_3294_ (
  .A1({ S65 }),
  .A2({ S25957[1161] }),
  .ZN({ S20141 })
);
OAI21_X1 #() 
OAI21_X1_1714_ (
  .A({ S20140 }),
  .B1({ S20133 }),
  .B2({ S20141 }),
  .ZN({ S20142 })
);
NAND3_X1 #() 
NAND3_X1_3468_ (
  .A1({ S25957[1160] }),
  .A2({ S25957[1161] }),
  .A3({ S20138 }),
  .ZN({ S20143 })
);
NAND2_X1 #() 
NAND2_X1_3295_ (
  .A1({ S20125 }),
  .A2({ S20126 }),
  .ZN({ S20144 })
);
NAND3_X1 #() 
NAND3_X1_3469_ (
  .A1({ S20144 }),
  .A2({ S20137 }),
  .A3({ S25957[1162] }),
  .ZN({ S20145 })
);
NAND2_X1 #() 
NAND2_X1_3296_ (
  .A1({ S20143 }),
  .A2({ S20145 }),
  .ZN({ S20146 })
);
NAND2_X1 #() 
NAND2_X1_3297_ (
  .A1({ S20146 }),
  .A2({ S65 }),
  .ZN({ S20147 })
);
NAND4_X1 #() 
NAND4_X1_364_ (
  .A1({ S20125 }),
  .A2({ S17295 }),
  .A3({ S20126 }),
  .A4({ S17328 }),
  .ZN({ S20148 })
);
INV_X1 #() 
INV_X1_1114_ (
  .A({ S20148 }),
  .ZN({ S20149 })
);
NAND4_X1 #() 
NAND4_X1_365_ (
  .A1({ S20127 }),
  .A2({ S20134 }),
  .A3({ S20135 }),
  .A4({ S20128 }),
  .ZN({ S20150 })
);
NOR2_X1 #() 
NOR2_X1_845_ (
  .A1({ S20150 }),
  .A2({ S25957[1160] }),
  .ZN({ S20151 })
);
OAI21_X1 #() 
OAI21_X1_1715_ (
  .A({ S25957[1163] }),
  .B1({ S20151 }),
  .B2({ S20149 }),
  .ZN({ S20152 })
);
NAND3_X1 #() 
NAND3_X1_3470_ (
  .A1({ S20147 }),
  .A2({ S20131 }),
  .A3({ S20152 }),
  .ZN({ S20153 })
);
OAI21_X1 #() 
OAI21_X1_1716_ (
  .A({ S20153 }),
  .B1({ S20131 }),
  .B2({ S20142 }),
  .ZN({ S20154 })
);
NAND4_X1 #() 
NAND4_X1_366_ (
  .A1({ S17295 }),
  .A2({ S20134 }),
  .A3({ S20135 }),
  .A4({ S17328 }),
  .ZN({ S20155 })
);
NAND2_X1 #() 
NAND2_X1_3298_ (
  .A1({ S20155 }),
  .A2({ S25957[1163] }),
  .ZN({ S20156 })
);
NOR2_X1 #() 
NOR2_X1_846_ (
  .A1({ S20156 }),
  .A2({ S72 }),
  .ZN({ S20157 })
);
AOI22_X1 #() 
AOI22_X1_375_ (
  .A1({ S20144 }),
  .A2({ S25957[1161] }),
  .B1({ S16086 }),
  .B2({ S16053 }),
  .ZN({ S20158 })
);
OAI21_X1 #() 
OAI21_X1_1717_ (
  .A({ S25957[1164] }),
  .B1({ S20157 }),
  .B2({ S20158 }),
  .ZN({ S20159 })
);
NAND4_X1 #() 
NAND4_X1_367_ (
  .A1({ S20125 }),
  .A2({ S20126 }),
  .A3({ S20134 }),
  .A4({ S20135 }),
  .ZN({ S20160 })
);
NAND4_X1 #() 
NAND4_X1_368_ (
  .A1({ S17295 }),
  .A2({ S17987 }),
  .A3({ S18019 }),
  .A4({ S17328 }),
  .ZN({ S20161 })
);
OAI211_X1 #() 
OAI211_X1_1130_ (
  .A({ S20160 }),
  .B({ S20150 }),
  .C1({ S20161 }),
  .C2({ S25957[1160] }),
  .ZN({ S20162 })
);
NAND3_X1 #() 
NAND3_X1_3471_ (
  .A1({ S25957[1163] }),
  .A2({ S25957[1160] }),
  .A3({ S20137 }),
  .ZN({ S20163 })
);
INV_X1 #() 
INV_X1_1115_ (
  .A({ S20163 }),
  .ZN({ S20164 })
);
NOR3_X1 #() 
NOR3_X1_118_ (
  .A1({ S20164 }),
  .A2({ S20162 }),
  .A3({ S25957[1164] }),
  .ZN({ S20165 })
);
NOR2_X1 #() 
NOR2_X1_847_ (
  .A1({ S20165 }),
  .A2({ S25957[1165] }),
  .ZN({ S20166 })
);
AOI22_X1 #() 
AOI22_X1_376_ (
  .A1({ S20154 }),
  .A2({ S25957[1165] }),
  .B1({ S20166 }),
  .B2({ S20159 }),
  .ZN({ S20167 })
);
AOI22_X1 #() 
AOI22_X1_377_ (
  .A1({ S16603 }),
  .A2({ S16571 }),
  .B1({ S17987 }),
  .B2({ S18019 }),
  .ZN({ S20168 })
);
OAI21_X1 #() 
OAI21_X1_1718_ (
  .A({ S25957[1163] }),
  .B1({ S20168 }),
  .B2({ S20137 }),
  .ZN({ S20169 })
);
OAI21_X1 #() 
OAI21_X1_1719_ (
  .A({ S20169 }),
  .B1({ S20168 }),
  .B2({ S20141 }),
  .ZN({ S20170 })
);
OAI21_X1 #() 
OAI21_X1_1720_ (
  .A({ S65 }),
  .B1({ S20161 }),
  .B2({ S25957[1160] }),
  .ZN({ S20171 })
);
NAND3_X1 #() 
NAND3_X1_3472_ (
  .A1({ S20171 }),
  .A2({ S20131 }),
  .A3({ S20129 }),
  .ZN({ S20172 })
);
OAI211_X1 #() 
OAI211_X1_1131_ (
  .A({ S25957[1165] }),
  .B({ S20172 }),
  .C1({ S20170 }),
  .C2({ S20131 }),
  .ZN({ S20173 })
);
NAND2_X1 #() 
NAND2_X1_3299_ (
  .A1({ S20148 }),
  .A2({ S20138 }),
  .ZN({ S20174 })
);
NAND2_X1 #() 
NAND2_X1_3300_ (
  .A1({ S20129 }),
  .A2({ S25957[1162] }),
  .ZN({ S20175 })
);
AOI21_X1 #() 
AOI21_X1_1788_ (
  .A({ S25957[1163] }),
  .B1({ S20174 }),
  .B2({ S20175 }),
  .ZN({ S20176 })
);
INV_X1 #() 
INV_X1_1116_ (
  .A({ S20161 }),
  .ZN({ S20177 })
);
AOI21_X1 #() 
AOI21_X1_1789_ (
  .A({ S25957[1164] }),
  .B1({ S20177 }),
  .B2({ S25957[1163] }),
  .ZN({ S20178 })
);
INV_X1 #() 
INV_X1_1117_ (
  .A({ S20178 }),
  .ZN({ S20179 })
);
NAND2_X1 #() 
NAND2_X1_3301_ (
  .A1({ S20161 }),
  .A2({ S20144 }),
  .ZN({ S20180 })
);
AOI21_X1 #() 
AOI21_X1_1790_ (
  .A({ S20179 }),
  .B1({ S20176 }),
  .B2({ S20180 }),
  .ZN({ S20181 })
);
NAND4_X1 #() 
NAND4_X1_369_ (
  .A1({ S16571 }),
  .A2({ S20127 }),
  .A3({ S16603 }),
  .A4({ S20128 }),
  .ZN({ S20182 })
);
NAND3_X1 #() 
NAND3_X1_3473_ (
  .A1({ S20148 }),
  .A2({ S20182 }),
  .A3({ S25957[1162] }),
  .ZN({ S20183 })
);
NAND3_X1 #() 
NAND3_X1_3474_ (
  .A1({ S20129 }),
  .A2({ S73 }),
  .A3({ S20138 }),
  .ZN({ S20184 })
);
NAND3_X1 #() 
NAND3_X1_3475_ (
  .A1({ S20183 }),
  .A2({ S20184 }),
  .A3({ S25957[1163] }),
  .ZN({ S20185 })
);
AOI21_X1 #() 
AOI21_X1_1791_ (
  .A({ S25957[1163] }),
  .B1({ S25957[1160] }),
  .B2({ S20138 }),
  .ZN({ S20186 })
);
NAND2_X1 #() 
NAND2_X1_3302_ (
  .A1({ S20186 }),
  .A2({ S20150 }),
  .ZN({ S20187 })
);
AOI21_X1 #() 
AOI21_X1_1792_ (
  .A({ S20131 }),
  .B1({ S20185 }),
  .B2({ S20187 }),
  .ZN({ S20188 })
);
OAI21_X1 #() 
OAI21_X1_1721_ (
  .A({ S14483 }),
  .B1({ S20181 }),
  .B2({ S20188 }),
  .ZN({ S20189 })
);
NAND3_X1 #() 
NAND3_X1_3476_ (
  .A1({ S20189 }),
  .A2({ S20130 }),
  .A3({ S20173 }),
  .ZN({ S20190 })
);
OAI211_X1 #() 
OAI211_X1_1132_ (
  .A({ S20190 }),
  .B({ S25957[1167] }),
  .C1({ S20167 }),
  .C2({ S20130 }),
  .ZN({ S20191 })
);
INV_X1 #() 
INV_X1_1118_ (
  .A({ S25957[1167] }),
  .ZN({ S20192 })
);
NAND4_X1 #() 
NAND4_X1_370_ (
  .A1({ S20127 }),
  .A2({ S17987 }),
  .A3({ S18019 }),
  .A4({ S20128 }),
  .ZN({ S20193 })
);
AOI22_X1 #() 
AOI22_X1_378_ (
  .A1({ S25957[1160] }),
  .A2({ S25957[1162] }),
  .B1({ S16114 }),
  .B2({ S16104 }),
  .ZN({ S20194 })
);
NAND2_X1 #() 
NAND2_X1_3303_ (
  .A1({ S20194 }),
  .A2({ S20193 }),
  .ZN({ S20195 })
);
NAND3_X1 #() 
NAND3_X1_3477_ (
  .A1({ S20193 }),
  .A2({ S20155 }),
  .A3({ S25957[1160] }),
  .ZN({ S20196 })
);
AOI21_X1 #() 
AOI21_X1_1793_ (
  .A({ S25957[1164] }),
  .B1({ S20196 }),
  .B2({ S65 }),
  .ZN({ S20197 })
);
NAND2_X1 #() 
NAND2_X1_3304_ (
  .A1({ S20197 }),
  .A2({ S20195 }),
  .ZN({ S20198 })
);
AOI21_X1 #() 
AOI21_X1_1794_ (
  .A({ S25957[1163] }),
  .B1({ S20183 }),
  .B2({ S20132 }),
  .ZN({ S20199 })
);
NAND3_X1 #() 
NAND3_X1_3478_ (
  .A1({ S20148 }),
  .A2({ S20182 }),
  .A3({ S20138 }),
  .ZN({ S20200 })
);
AOI21_X1 #() 
AOI21_X1_1795_ (
  .A({ S65 }),
  .B1({ S20200 }),
  .B2({ S20175 }),
  .ZN({ S20201 })
);
OR3_X1 #() 
OR3_X1_19_ (
  .A1({ S20201 }),
  .A2({ S20199 }),
  .A3({ S20131 }),
  .ZN({ S20202 })
);
AOI21_X1 #() 
AOI21_X1_1796_ (
  .A({ S25957[1165] }),
  .B1({ S20202 }),
  .B2({ S20198 }),
  .ZN({ S20203 })
);
NOR2_X1 #() 
NOR2_X1_848_ (
  .A1({ S20146 }),
  .A2({ S65 }),
  .ZN({ S20204 })
);
AOI21_X1 #() 
AOI21_X1_1797_ (
  .A({ S25957[1160] }),
  .B1({ S20137 }),
  .B2({ S25957[1162] }),
  .ZN({ S20205 })
);
OAI21_X1 #() 
OAI21_X1_1722_ (
  .A({ S25957[1164] }),
  .B1({ S20205 }),
  .B2({ S25957[1163] }),
  .ZN({ S20206 })
);
NAND4_X1 #() 
NAND4_X1_371_ (
  .A1({ S20155 }),
  .A2({ S20132 }),
  .A3({ S20193 }),
  .A4({ S25957[1163] }),
  .ZN({ S20207 })
);
NAND3_X1 #() 
NAND3_X1_3479_ (
  .A1({ S20136 }),
  .A2({ S20155 }),
  .A3({ S65 }),
  .ZN({ S20208 })
);
NAND3_X1 #() 
NAND3_X1_3480_ (
  .A1({ S20207 }),
  .A2({ S20131 }),
  .A3({ S20208 }),
  .ZN({ S20209 })
);
OAI21_X1 #() 
OAI21_X1_1723_ (
  .A({ S20209 }),
  .B1({ S20204 }),
  .B2({ S20206 }),
  .ZN({ S20210 })
);
OAI21_X1 #() 
OAI21_X1_1724_ (
  .A({ S25957[1166] }),
  .B1({ S20210 }),
  .B2({ S14483 }),
  .ZN({ S20211 })
);
AOI22_X1 #() 
AOI22_X1_379_ (
  .A1({ S20136 }),
  .A2({ S20150 }),
  .B1({ S20144 }),
  .B2({ S25957[1161] }),
  .ZN({ S20212 })
);
NOR2_X1 #() 
NOR2_X1_849_ (
  .A1({ S20212 }),
  .A2({ S25957[1163] }),
  .ZN({ S20213 })
);
AOI21_X1 #() 
AOI21_X1_1798_ (
  .A({ S20213 }),
  .B1({ S20175 }),
  .B2({ S25957[1163] }),
  .ZN({ S20214 })
);
NOR2_X1 #() 
NOR2_X1_850_ (
  .A1({ S20214 }),
  .A2({ S25957[1164] }),
  .ZN({ S20215 })
);
NAND3_X1 #() 
NAND3_X1_3481_ (
  .A1({ S20144 }),
  .A2({ S25957[1161] }),
  .A3({ S25957[1162] }),
  .ZN({ S20216 })
);
NAND3_X1 #() 
NAND3_X1_3482_ (
  .A1({ S25957[1160] }),
  .A2({ S20137 }),
  .A3({ S25957[1162] }),
  .ZN({ S20217 })
);
NAND2_X1 #() 
NAND2_X1_3305_ (
  .A1({ S20216 }),
  .A2({ S20217 }),
  .ZN({ S20218 })
);
NAND2_X1 #() 
NAND2_X1_3306_ (
  .A1({ S20143 }),
  .A2({ S65 }),
  .ZN({ S20219 })
);
OAI22_X1 #() 
OAI22_X1_94_ (
  .A1({ S20218 }),
  .A2({ S20219 }),
  .B1({ S20151 }),
  .B2({ S65 }),
  .ZN({ S20220 })
);
OAI21_X1 #() 
OAI21_X1_1725_ (
  .A({ S14483 }),
  .B1({ S20220 }),
  .B2({ S20131 }),
  .ZN({ S20221 })
);
NAND2_X1 #() 
NAND2_X1_3307_ (
  .A1({ S20129 }),
  .A2({ S20138 }),
  .ZN({ S20222 })
);
AND2_X1 #() 
AND2_X1_205_ (
  .A1({ S20193 }),
  .A2({ S25957[1163] }),
  .ZN({ S20223 })
);
NAND2_X1 #() 
NAND2_X1_3308_ (
  .A1({ S20150 }),
  .A2({ S65 }),
  .ZN({ S20224 })
);
INV_X1 #() 
INV_X1_1119_ (
  .A({ S20224 }),
  .ZN({ S20225 })
);
AOI22_X1 #() 
AOI22_X1_380_ (
  .A1({ S20225 }),
  .A2({ S20222 }),
  .B1({ S20223 }),
  .B2({ S20148 }),
  .ZN({ S20226 })
);
NAND2_X1 #() 
NAND2_X1_3309_ (
  .A1({ S65 }),
  .A2({ S25957[1160] }),
  .ZN({ S20227 })
);
NAND3_X1 #() 
NAND3_X1_3483_ (
  .A1({ S20160 }),
  .A2({ S20161 }),
  .A3({ S25957[1163] }),
  .ZN({ S20228 })
);
NAND3_X1 #() 
NAND3_X1_3484_ (
  .A1({ S20228 }),
  .A2({ S25957[1164] }),
  .A3({ S20227 }),
  .ZN({ S20229 })
);
OAI211_X1 #() 
OAI211_X1_1133_ (
  .A({ S25957[1165] }),
  .B({ S20229 }),
  .C1({ S20226 }),
  .C2({ S25957[1164] }),
  .ZN({ S20230 })
);
OAI211_X1 #() 
OAI211_X1_1134_ (
  .A({ S20130 }),
  .B({ S20230 }),
  .C1({ S20215 }),
  .C2({ S20221 }),
  .ZN({ S20231 })
);
OAI21_X1 #() 
OAI21_X1_1726_ (
  .A({ S20231 }),
  .B1({ S20203 }),
  .B2({ S20211 }),
  .ZN({ S20232 })
);
NAND2_X1 #() 
NAND2_X1_3310_ (
  .A1({ S20232 }),
  .A2({ S20192 }),
  .ZN({ S20233 })
);
NAND3_X1 #() 
NAND3_X1_3485_ (
  .A1({ S20233 }),
  .A2({ S6978 }),
  .A3({ S20191 }),
  .ZN({ S20234 })
);
INV_X1 #() 
INV_X1_1120_ (
  .A({ S6978 }),
  .ZN({ S25957[1271] })
);
NAND2_X1 #() 
NAND2_X1_3311_ (
  .A1({ S20233 }),
  .A2({ S20191 }),
  .ZN({ S20235 })
);
NAND2_X1 #() 
NAND2_X1_3312_ (
  .A1({ S20235 }),
  .A2({ S25957[1271] }),
  .ZN({ S20236 })
);
NAND3_X1 #() 
NAND3_X1_3486_ (
  .A1({ S20236 }),
  .A2({ S25957[1239] }),
  .A3({ S20234 }),
  .ZN({ S20237 })
);
NAND2_X1 #() 
NAND2_X1_3313_ (
  .A1({ S20236 }),
  .A2({ S20234 }),
  .ZN({ S25957[1143] })
);
NAND2_X1 #() 
NAND2_X1_3314_ (
  .A1({ S25957[1143] }),
  .A2({ S6989 }),
  .ZN({ S20238 })
);
NAND2_X1 #() 
NAND2_X1_3315_ (
  .A1({ S20238 }),
  .A2({ S20237 }),
  .ZN({ S25957[1111] })
);
INV_X1 #() 
INV_X1_1121_ (
  .A({ S25957[1111] }),
  .ZN({ S20239 })
);
NAND2_X1 #() 
NAND2_X1_3316_ (
  .A1({ S20239 }),
  .A2({ S5675 }),
  .ZN({ S20240 })
);
NAND2_X1 #() 
NAND2_X1_3317_ (
  .A1({ S25957[1111] }),
  .A2({ S25956[23] }),
  .ZN({ S20241 })
);
NAND2_X1 #() 
NAND2_X1_3318_ (
  .A1({ S20240 }),
  .A2({ S20241 }),
  .ZN({ S20242 })
);
INV_X1 #() 
INV_X1_1122_ (
  .A({ S20242 }),
  .ZN({ S25957[1047] })
);
NAND2_X1 #() 
NAND2_X1_3319_ (
  .A1({ S73 }),
  .A2({ S25957[1162] }),
  .ZN({ S20243 })
);
NAND4_X1 #() 
NAND4_X1_372_ (
  .A1({ S20125 }),
  .A2({ S20126 }),
  .A3({ S17987 }),
  .A4({ S18019 }),
  .ZN({ S20244 })
);
NAND4_X1 #() 
NAND4_X1_373_ (
  .A1({ S20136 }),
  .A2({ S20244 }),
  .A3({ S25957[1163] }),
  .A4({ S20137 }),
  .ZN({ S20245 })
);
OAI211_X1 #() 
OAI211_X1_1135_ (
  .A({ S20245 }),
  .B({ S25957[1164] }),
  .C1({ S25957[1163] }),
  .C2({ S20243 }),
  .ZN({ S20246 })
);
INV_X1 #() 
INV_X1_1123_ (
  .A({ S20141 }),
  .ZN({ S20247 })
);
OAI21_X1 #() 
OAI21_X1_1727_ (
  .A({ S20131 }),
  .B1({ S20157 }),
  .B2({ S20247 }),
  .ZN({ S20248 })
);
NAND3_X1 #() 
NAND3_X1_3487_ (
  .A1({ S20248 }),
  .A2({ S25957[1165] }),
  .A3({ S20246 }),
  .ZN({ S20249 })
);
INV_X1 #() 
INV_X1_1124_ (
  .A({ S20200 }),
  .ZN({ S20250 })
);
NAND2_X1 #() 
NAND2_X1_3320_ (
  .A1({ S20136 }),
  .A2({ S65 }),
  .ZN({ S20251 })
);
NAND2_X1 #() 
NAND2_X1_3321_ (
  .A1({ S20182 }),
  .A2({ S25957[1162] }),
  .ZN({ S20252 })
);
NAND3_X1 #() 
NAND3_X1_3488_ (
  .A1({ S20252 }),
  .A2({ S25957[1163] }),
  .A3({ S20132 }),
  .ZN({ S20253 })
);
OAI21_X1 #() 
OAI21_X1_1728_ (
  .A({ S20253 }),
  .B1({ S20250 }),
  .B2({ S20251 }),
  .ZN({ S20254 })
);
OAI21_X1 #() 
OAI21_X1_1729_ (
  .A({ S20169 }),
  .B1({ S25957[1163] }),
  .B2({ S20174 }),
  .ZN({ S20255 })
);
AOI21_X1 #() 
AOI21_X1_1799_ (
  .A({ S25957[1165] }),
  .B1({ S20255 }),
  .B2({ S25957[1164] }),
  .ZN({ S20256 })
);
OAI21_X1 #() 
OAI21_X1_1730_ (
  .A({ S20256 }),
  .B1({ S25957[1164] }),
  .B2({ S20254 }),
  .ZN({ S20257 })
);
OAI21_X1 #() 
OAI21_X1_1731_ (
  .A({ S73 }),
  .B1({ S20160 }),
  .B2({ S20137 }),
  .ZN({ S20258 })
);
INV_X1 #() 
INV_X1_1125_ (
  .A({ S20155 }),
  .ZN({ S20259 })
);
NAND3_X1 #() 
NAND3_X1_3489_ (
  .A1({ S20144 }),
  .A2({ S25957[1161] }),
  .A3({ S20138 }),
  .ZN({ S20260 })
);
INV_X1 #() 
INV_X1_1126_ (
  .A({ S20260 }),
  .ZN({ S20261 })
);
OAI21_X1 #() 
OAI21_X1_1732_ (
  .A({ S25957[1163] }),
  .B1({ S20261 }),
  .B2({ S20259 }),
  .ZN({ S20262 })
);
OAI211_X1 #() 
OAI211_X1_1136_ (
  .A({ S20262 }),
  .B({ S20131 }),
  .C1({ S25957[1163] }),
  .C2({ S20258 }),
  .ZN({ S20263 })
);
NAND2_X1 #() 
NAND2_X1_3322_ (
  .A1({ S20212 }),
  .A2({ S65 }),
  .ZN({ S20264 })
);
NAND3_X1 #() 
NAND3_X1_3490_ (
  .A1({ S20133 }),
  .A2({ S65 }),
  .A3({ S25957[1161] }),
  .ZN({ S20265 })
);
INV_X1 #() 
INV_X1_1127_ (
  .A({ S20150 }),
  .ZN({ S20266 })
);
AOI21_X1 #() 
AOI21_X1_1800_ (
  .A({ S20131 }),
  .B1({ S20266 }),
  .B2({ S25957[1163] }),
  .ZN({ S20267 })
);
NAND3_X1 #() 
NAND3_X1_3491_ (
  .A1({ S20264 }),
  .A2({ S20265 }),
  .A3({ S20267 }),
  .ZN({ S20268 })
);
NAND3_X1 #() 
NAND3_X1_3492_ (
  .A1({ S20263 }),
  .A2({ S25957[1165] }),
  .A3({ S20268 }),
  .ZN({ S20269 })
);
AOI21_X1 #() 
AOI21_X1_1801_ (
  .A({ S25957[1166] }),
  .B1({ S20257 }),
  .B2({ S20269 }),
  .ZN({ S20270 })
);
AOI21_X1 #() 
AOI21_X1_1802_ (
  .A({ S65 }),
  .B1({ S20259 }),
  .B2({ S20144 }),
  .ZN({ S20271 })
);
NAND3_X1 #() 
NAND3_X1_3493_ (
  .A1({ S20129 }),
  .A2({ S25957[1163] }),
  .A3({ S20138 }),
  .ZN({ S20272 })
);
OAI211_X1 #() 
OAI211_X1_1137_ (
  .A({ S20131 }),
  .B({ S20272 }),
  .C1({ S20176 }),
  .C2({ S20271 }),
  .ZN({ S20273 })
);
NAND3_X1 #() 
NAND3_X1_3494_ (
  .A1({ S20244 }),
  .A2({ S20136 }),
  .A3({ S20150 }),
  .ZN({ S20274 })
);
NAND2_X1 #() 
NAND2_X1_3323_ (
  .A1({ S20274 }),
  .A2({ S25957[1163] }),
  .ZN({ S20275 })
);
OAI21_X1 #() 
OAI21_X1_1733_ (
  .A({ S20275 }),
  .B1({ S20250 }),
  .B2({ S20251 }),
  .ZN({ S20276 })
);
AOI21_X1 #() 
AOI21_X1_1803_ (
  .A({ S25957[1165] }),
  .B1({ S20276 }),
  .B2({ S25957[1164] }),
  .ZN({ S20277 })
);
AOI21_X1 #() 
AOI21_X1_1804_ (
  .A({ S20130 }),
  .B1({ S20277 }),
  .B2({ S20273 }),
  .ZN({ S20278 })
);
AOI21_X1 #() 
AOI21_X1_1805_ (
  .A({ S20270 }),
  .B1({ S20249 }),
  .B2({ S20278 }),
  .ZN({ S20279 })
);
NAND2_X1 #() 
NAND2_X1_3324_ (
  .A1({ S20182 }),
  .A2({ S20160 }),
  .ZN({ S20280 })
);
NAND4_X1 #() 
NAND4_X1_374_ (
  .A1({ S20136 }),
  .A2({ S20244 }),
  .A3({ S20155 }),
  .A4({ S65 }),
  .ZN({ S20281 })
);
NAND2_X1 #() 
NAND2_X1_3325_ (
  .A1({ S20281 }),
  .A2({ S25957[1164] }),
  .ZN({ S20282 })
);
AOI21_X1 #() 
AOI21_X1_1806_ (
  .A({ S20282 }),
  .B1({ S20280 }),
  .B2({ S25957[1163] }),
  .ZN({ S20283 })
);
NOR2_X1 #() 
NOR2_X1_851_ (
  .A1({ S20160 }),
  .A2({ S65 }),
  .ZN({ S20284 })
);
NAND2_X1 #() 
NAND2_X1_3326_ (
  .A1({ S20182 }),
  .A2({ S20150 }),
  .ZN({ S20285 })
);
NOR2_X1 #() 
NOR2_X1_852_ (
  .A1({ S20284 }),
  .A2({ S20285 }),
  .ZN({ S20286 })
);
NOR2_X1 #() 
NOR2_X1_853_ (
  .A1({ S20286 }),
  .A2({ S25957[1164] }),
  .ZN({ S20287 })
);
OAI21_X1 #() 
OAI21_X1_1734_ (
  .A({ S25957[1165] }),
  .B1({ S20283 }),
  .B2({ S20287 }),
  .ZN({ S20288 })
);
INV_X1 #() 
INV_X1_1128_ (
  .A({ S20193 }),
  .ZN({ S20289 })
);
NAND2_X1 #() 
NAND2_X1_3327_ (
  .A1({ S20289 }),
  .A2({ S25957[1163] }),
  .ZN({ S20290 })
);
OAI211_X1 #() 
OAI211_X1_1138_ (
  .A({ S20290 }),
  .B({ S25957[1164] }),
  .C1({ S25957[1163] }),
  .C2({ S20180 }),
  .ZN({ S20291 })
);
AOI21_X1 #() 
AOI21_X1_1807_ (
  .A({ S25957[1164] }),
  .B1({ S20274 }),
  .B2({ S25957[1163] }),
  .ZN({ S20292 })
);
OAI21_X1 #() 
OAI21_X1_1735_ (
  .A({ S20292 }),
  .B1({ S25957[1163] }),
  .B2({ S20218 }),
  .ZN({ S20293 })
);
NAND3_X1 #() 
NAND3_X1_3495_ (
  .A1({ S20293 }),
  .A2({ S14483 }),
  .A3({ S20291 }),
  .ZN({ S20294 })
);
NAND3_X1 #() 
NAND3_X1_3496_ (
  .A1({ S20288 }),
  .A2({ S25957[1166] }),
  .A3({ S20294 }),
  .ZN({ S20295 })
);
AOI21_X1 #() 
AOI21_X1_1808_ (
  .A({ S20131 }),
  .B1({ S20139 }),
  .B2({ S65 }),
  .ZN({ S20296 })
);
NAND2_X1 #() 
NAND2_X1_3328_ (
  .A1({ S20182 }),
  .A2({ S20138 }),
  .ZN({ S20297 })
);
NAND2_X1 #() 
NAND2_X1_3329_ (
  .A1({ S20297 }),
  .A2({ S20216 }),
  .ZN({ S20298 })
);
NAND2_X1 #() 
NAND2_X1_3330_ (
  .A1({ S20298 }),
  .A2({ S25957[1163] }),
  .ZN({ S20299 })
);
NOR2_X1 #() 
NOR2_X1_854_ (
  .A1({ S20299 }),
  .A2({ S25957[1164] }),
  .ZN({ S20300 })
);
AOI21_X1 #() 
AOI21_X1_1809_ (
  .A({ S20300 }),
  .B1({ S20296 }),
  .B2({ S20207 }),
  .ZN({ S20301 })
);
NOR2_X1 #() 
NOR2_X1_855_ (
  .A1({ S20186 }),
  .A2({ S20131 }),
  .ZN({ S20302 })
);
NOR2_X1 #() 
NOR2_X1_856_ (
  .A1({ S20157 }),
  .A2({ S20164 }),
  .ZN({ S20303 })
);
AOI22_X1 #() 
AOI22_X1_381_ (
  .A1({ S20225 }),
  .A2({ S20139 }),
  .B1({ S20223 }),
  .B2({ S20155 }),
  .ZN({ S20304 })
);
AOI22_X1 #() 
AOI22_X1_382_ (
  .A1({ S20304 }),
  .A2({ S20131 }),
  .B1({ S20303 }),
  .B2({ S20302 }),
  .ZN({ S20305 })
);
NAND2_X1 #() 
NAND2_X1_3331_ (
  .A1({ S20305 }),
  .A2({ S25957[1165] }),
  .ZN({ S20306 })
);
OAI211_X1 #() 
OAI211_X1_1139_ (
  .A({ S20306 }),
  .B({ S20130 }),
  .C1({ S25957[1165] }),
  .C2({ S20301 }),
  .ZN({ S20307 })
);
NAND3_X1 #() 
NAND3_X1_3497_ (
  .A1({ S20307 }),
  .A2({ S20192 }),
  .A3({ S20295 }),
  .ZN({ S20308 })
);
OAI21_X1 #() 
OAI21_X1_1736_ (
  .A({ S20308 }),
  .B1({ S20279 }),
  .B2({ S20192 }),
  .ZN({ S20309 })
);
NAND2_X1 #() 
NAND2_X1_3332_ (
  .A1({ S20309 }),
  .A2({ S25957[1270] }),
  .ZN({ S20310 })
);
INV_X1 #() 
INV_X1_1129_ (
  .A({ S25957[1270] }),
  .ZN({ S20311 })
);
OAI211_X1 #() 
OAI211_X1_1140_ (
  .A({ S20311 }),
  .B({ S20308 }),
  .C1({ S20279 }),
  .C2({ S20192 }),
  .ZN({ S20312 })
);
NAND2_X1 #() 
NAND2_X1_3333_ (
  .A1({ S20310 }),
  .A2({ S20312 }),
  .ZN({ S25957[1142] })
);
NOR2_X1 #() 
NOR2_X1_857_ (
  .A1({ S25957[1142] }),
  .A2({ S25957[1238] }),
  .ZN({ S20313 })
);
NAND2_X1 #() 
NAND2_X1_3334_ (
  .A1({ S25957[1142] }),
  .A2({ S25957[1238] }),
  .ZN({ S20314 })
);
INV_X1 #() 
INV_X1_1130_ (
  .A({ S20314 }),
  .ZN({ S20315 })
);
OAI21_X1 #() 
OAI21_X1_1737_ (
  .A({ S25956[22] }),
  .B1({ S20315 }),
  .B2({ S20313 }),
  .ZN({ S20316 })
);
NOR2_X1 #() 
NOR2_X1_858_ (
  .A1({ S20315 }),
  .A2({ S20313 }),
  .ZN({ S25957[1110] })
);
NAND2_X1 #() 
NAND2_X1_3335_ (
  .A1({ S25957[1110] }),
  .A2({ S19541 }),
  .ZN({ S20317 })
);
NAND2_X1 #() 
NAND2_X1_3336_ (
  .A1({ S20317 }),
  .A2({ S20316 }),
  .ZN({ S25957[1046] })
);
INV_X1 #() 
INV_X1_1131_ (
  .A({ S25957[1269] }),
  .ZN({ S20318 })
);
NAND3_X1 #() 
NAND3_X1_3498_ (
  .A1({ S20244 }),
  .A2({ S20161 }),
  .A3({ S25957[1163] }),
  .ZN({ S20319 })
);
AOI21_X1 #() 
AOI21_X1_1810_ (
  .A({ S20131 }),
  .B1({ S20158 }),
  .B2({ S25957[1162] }),
  .ZN({ S20320 })
);
AOI22_X1 #() 
AOI22_X1_383_ (
  .A1({ S20292 }),
  .A2({ S20264 }),
  .B1({ S20320 }),
  .B2({ S20319 }),
  .ZN({ S20321 })
);
NAND2_X1 #() 
NAND2_X1_3337_ (
  .A1({ S25957[1163] }),
  .A2({ S20144 }),
  .ZN({ S20322 })
);
NAND3_X1 #() 
NAND3_X1_3499_ (
  .A1({ S20174 }),
  .A2({ S65 }),
  .A3({ S20216 }),
  .ZN({ S20323 })
);
OAI21_X1 #() 
OAI21_X1_1738_ (
  .A({ S20323 }),
  .B1({ S20177 }),
  .B2({ S20322 }),
  .ZN({ S20324 })
);
NAND3_X1 #() 
NAND3_X1_3500_ (
  .A1({ S20129 }),
  .A2({ S20150 }),
  .A3({ S25957[1163] }),
  .ZN({ S20325 })
);
NAND3_X1 #() 
NAND3_X1_3501_ (
  .A1({ S20325 }),
  .A2({ S20160 }),
  .A3({ S20141 }),
  .ZN({ S20326 })
);
NAND3_X1 #() 
NAND3_X1_3502_ (
  .A1({ S20326 }),
  .A2({ S15250 }),
  .A3({ S15283 }),
  .ZN({ S20327 })
);
OAI211_X1 #() 
OAI211_X1_1141_ (
  .A({ S20327 }),
  .B({ S25957[1165] }),
  .C1({ S20324 }),
  .C2({ S20131 }),
  .ZN({ S20328 })
);
OAI211_X1 #() 
OAI211_X1_1142_ (
  .A({ S20328 }),
  .B({ S25957[1166] }),
  .C1({ S25957[1165] }),
  .C2({ S20321 }),
  .ZN({ S20329 })
);
AOI21_X1 #() 
AOI21_X1_1811_ (
  .A({ S25957[1163] }),
  .B1({ S20289 }),
  .B2({ S25957[1160] }),
  .ZN({ S20330 })
);
NAND3_X1 #() 
NAND3_X1_3503_ (
  .A1({ S20129 }),
  .A2({ S73 }),
  .A3({ S25957[1162] }),
  .ZN({ S20331 })
);
NAND3_X1 #() 
NAND3_X1_3504_ (
  .A1({ S20144 }),
  .A2({ S20137 }),
  .A3({ S20138 }),
  .ZN({ S20332 })
);
AOI21_X1 #() 
AOI21_X1_1812_ (
  .A({ S65 }),
  .B1({ S20331 }),
  .B2({ S20332 }),
  .ZN({ S20333 })
);
NOR3_X1 #() 
NOR3_X1_119_ (
  .A1({ S20333 }),
  .A2({ S20330 }),
  .A3({ S25957[1164] }),
  .ZN({ S20334 })
);
AOI21_X1 #() 
AOI21_X1_1813_ (
  .A({ S25957[1162] }),
  .B1({ S20148 }),
  .B2({ S20182 }),
  .ZN({ S20335 })
);
AOI22_X1 #() 
AOI22_X1_384_ (
  .A1({ S20335 }),
  .A2({ S25957[1163] }),
  .B1({ S20186 }),
  .B2({ S20137 }),
  .ZN({ S20336 })
);
OAI21_X1 #() 
OAI21_X1_1739_ (
  .A({ S14483 }),
  .B1({ S20336 }),
  .B2({ S20131 }),
  .ZN({ S20337 })
);
NAND3_X1 #() 
NAND3_X1_3505_ (
  .A1({ S20182 }),
  .A2({ S20161 }),
  .A3({ S65 }),
  .ZN({ S20338 })
);
AOI21_X1 #() 
AOI21_X1_1814_ (
  .A({ S25957[1164] }),
  .B1({ S25957[1163] }),
  .B2({ S20137 }),
  .ZN({ S20339 })
);
NAND2_X1 #() 
NAND2_X1_3338_ (
  .A1({ S20339 }),
  .A2({ S20338 }),
  .ZN({ S20340 })
);
AOI21_X1 #() 
AOI21_X1_1815_ (
  .A({ S25957[1163] }),
  .B1({ S20144 }),
  .B2({ S20138 }),
  .ZN({ S20341 })
);
AOI21_X1 #() 
AOI21_X1_1816_ (
  .A({ S20131 }),
  .B1({ S20341 }),
  .B2({ S20129 }),
  .ZN({ S20342 })
);
OAI21_X1 #() 
OAI21_X1_1740_ (
  .A({ S20342 }),
  .B1({ S65 }),
  .B2({ S20196 }),
  .ZN({ S20343 })
);
NAND3_X1 #() 
NAND3_X1_3506_ (
  .A1({ S20343 }),
  .A2({ S25957[1165] }),
  .A3({ S20340 }),
  .ZN({ S20344 })
);
OAI21_X1 #() 
OAI21_X1_1741_ (
  .A({ S20344 }),
  .B1({ S20334 }),
  .B2({ S20337 }),
  .ZN({ S20345 })
);
NAND2_X1 #() 
NAND2_X1_3339_ (
  .A1({ S20345 }),
  .A2({ S20130 }),
  .ZN({ S20346 })
);
NAND3_X1 #() 
NAND3_X1_3507_ (
  .A1({ S20346 }),
  .A2({ S25957[1167] }),
  .A3({ S20329 }),
  .ZN({ S20347 })
);
NAND3_X1 #() 
NAND3_X1_3508_ (
  .A1({ S25957[1160] }),
  .A2({ S25957[1161] }),
  .A3({ S25957[1162] }),
  .ZN({ S20348 })
);
NAND2_X1 #() 
NAND2_X1_3340_ (
  .A1({ S20348 }),
  .A2({ S20260 }),
  .ZN({ S20349 })
);
AOI21_X1 #() 
AOI21_X1_1817_ (
  .A({ S20284 }),
  .B1({ S20349 }),
  .B2({ S65 }),
  .ZN({ S20350 })
);
OAI21_X1 #() 
OAI21_X1_1742_ (
  .A({ S65 }),
  .B1({ S20193 }),
  .B2({ S25957[1160] }),
  .ZN({ S20351 })
);
NAND2_X1 #() 
NAND2_X1_3341_ (
  .A1({ S20351 }),
  .A2({ S20272 }),
  .ZN({ S20352 })
);
AOI21_X1 #() 
AOI21_X1_1818_ (
  .A({ S14483 }),
  .B1({ S20352 }),
  .B2({ S25957[1164] }),
  .ZN({ S20353 })
);
OAI21_X1 #() 
OAI21_X1_1743_ (
  .A({ S20353 }),
  .B1({ S25957[1164] }),
  .B2({ S20350 }),
  .ZN({ S20354 })
);
NAND4_X1 #() 
NAND4_X1_375_ (
  .A1({ S20182 }),
  .A2({ S20148 }),
  .A3({ S20132 }),
  .A4({ S65 }),
  .ZN({ S20355 })
);
NAND3_X1 #() 
NAND3_X1_3509_ (
  .A1({ S20183 }),
  .A2({ S25957[1163] }),
  .A3({ S20139 }),
  .ZN({ S20356 })
);
NAND3_X1 #() 
NAND3_X1_3510_ (
  .A1({ S20356 }),
  .A2({ S25957[1164] }),
  .A3({ S20355 }),
  .ZN({ S20357 })
);
NOR2_X1 #() 
NOR2_X1_859_ (
  .A1({ S20160 }),
  .A2({ S20137 }),
  .ZN({ S20358 })
);
AOI21_X1 #() 
AOI21_X1_1819_ (
  .A({ S20164 }),
  .B1({ S65 }),
  .B2({ S20358 }),
  .ZN({ S20359 })
);
OAI21_X1 #() 
OAI21_X1_1744_ (
  .A({ S20357 }),
  .B1({ S25957[1164] }),
  .B2({ S20359 }),
  .ZN({ S20360 })
);
OAI21_X1 #() 
OAI21_X1_1745_ (
  .A({ S20354 }),
  .B1({ S20360 }),
  .B2({ S25957[1165] }),
  .ZN({ S20361 })
);
NAND4_X1 #() 
NAND4_X1_376_ (
  .A1({ S20155 }),
  .A2({ S20132 }),
  .A3({ S20193 }),
  .A4({ S65 }),
  .ZN({ S20362 })
);
NAND3_X1 #() 
NAND3_X1_3511_ (
  .A1({ S20183 }),
  .A2({ S25957[1163] }),
  .A3({ S20260 }),
  .ZN({ S20363 })
);
AOI21_X1 #() 
AOI21_X1_1820_ (
  .A({ S20131 }),
  .B1({ S20363 }),
  .B2({ S20362 }),
  .ZN({ S20364 })
);
NAND3_X1 #() 
NAND3_X1_3512_ (
  .A1({ S20182 }),
  .A2({ S20244 }),
  .A3({ S65 }),
  .ZN({ S20365 })
);
NAND3_X1 #() 
NAND3_X1_3513_ (
  .A1({ S20365 }),
  .A2({ S20131 }),
  .A3({ S20322 }),
  .ZN({ S20366 })
);
NAND2_X1 #() 
NAND2_X1_3342_ (
  .A1({ S20366 }),
  .A2({ S25957[1165] }),
  .ZN({ S20367 })
);
NAND4_X1 #() 
NAND4_X1_377_ (
  .A1({ S20136 }),
  .A2({ S20244 }),
  .A3({ S20155 }),
  .A4({ S25957[1163] }),
  .ZN({ S20368 })
);
NAND3_X1 #() 
NAND3_X1_3514_ (
  .A1({ S20260 }),
  .A2({ S65 }),
  .A3({ S20160 }),
  .ZN({ S20369 })
);
AOI21_X1 #() 
AOI21_X1_1821_ (
  .A({ S25957[1164] }),
  .B1({ S20369 }),
  .B2({ S20368 }),
  .ZN({ S20370 })
);
AOI21_X1 #() 
AOI21_X1_1822_ (
  .A({ S25957[1163] }),
  .B1({ S20175 }),
  .B2({ S20143 }),
  .ZN({ S20371 })
);
NAND3_X1 #() 
NAND3_X1_3515_ (
  .A1({ S20148 }),
  .A2({ S25957[1163] }),
  .A3({ S20138 }),
  .ZN({ S20372 })
);
NAND2_X1 #() 
NAND2_X1_3343_ (
  .A1({ S20372 }),
  .A2({ S25957[1164] }),
  .ZN({ S20373 })
);
NOR2_X1 #() 
NOR2_X1_860_ (
  .A1({ S20371 }),
  .A2({ S20373 }),
  .ZN({ S20374 })
);
OAI21_X1 #() 
OAI21_X1_1746_ (
  .A({ S14483 }),
  .B1({ S20374 }),
  .B2({ S20370 }),
  .ZN({ S20375 })
);
OAI21_X1 #() 
OAI21_X1_1747_ (
  .A({ S20375 }),
  .B1({ S20364 }),
  .B2({ S20367 }),
  .ZN({ S20376 })
);
NAND2_X1 #() 
NAND2_X1_3344_ (
  .A1({ S20376 }),
  .A2({ S25957[1166] }),
  .ZN({ S20377 })
);
OAI211_X1 #() 
OAI211_X1_1143_ (
  .A({ S20377 }),
  .B({ S20192 }),
  .C1({ S25957[1166] }),
  .C2({ S20361 }),
  .ZN({ S20378 })
);
NAND3_X1 #() 
NAND3_X1_3516_ (
  .A1({ S20378 }),
  .A2({ S20347 }),
  .A3({ S20318 }),
  .ZN({ S20379 })
);
NAND2_X1 #() 
NAND2_X1_3345_ (
  .A1({ S20346 }),
  .A2({ S20329 }),
  .ZN({ S20380 })
);
NAND2_X1 #() 
NAND2_X1_3346_ (
  .A1({ S20380 }),
  .A2({ S25957[1167] }),
  .ZN({ S20381 })
);
AOI21_X1 #() 
AOI21_X1_1823_ (
  .A({ S25957[1167] }),
  .B1({ S20361 }),
  .B2({ S20130 }),
  .ZN({ S20382 })
);
OAI21_X1 #() 
OAI21_X1_1748_ (
  .A({ S20382 }),
  .B1({ S20130 }),
  .B2({ S20376 }),
  .ZN({ S20383 })
);
NAND3_X1 #() 
NAND3_X1_3517_ (
  .A1({ S20381 }),
  .A2({ S20383 }),
  .A3({ S25957[1269] }),
  .ZN({ S20384 })
);
NAND3_X1 #() 
NAND3_X1_3518_ (
  .A1({ S20384 }),
  .A2({ S25957[1237] }),
  .A3({ S20379 }),
  .ZN({ S20385 })
);
INV_X1 #() 
INV_X1_1132_ (
  .A({ S25957[1237] }),
  .ZN({ S20386 })
);
NAND3_X1 #() 
NAND3_X1_3519_ (
  .A1({ S20381 }),
  .A2({ S20383 }),
  .A3({ S20318 }),
  .ZN({ S20387 })
);
NAND3_X1 #() 
NAND3_X1_3520_ (
  .A1({ S20378 }),
  .A2({ S20347 }),
  .A3({ S25957[1269] }),
  .ZN({ S20388 })
);
NAND3_X1 #() 
NAND3_X1_3521_ (
  .A1({ S20387 }),
  .A2({ S20386 }),
  .A3({ S20388 }),
  .ZN({ S20389 })
);
NAND3_X1 #() 
NAND3_X1_3522_ (
  .A1({ S20385 }),
  .A2({ S20389 }),
  .A3({ S7762 }),
  .ZN({ S20390 })
);
NAND3_X1 #() 
NAND3_X1_3523_ (
  .A1({ S20384 }),
  .A2({ S20386 }),
  .A3({ S20379 }),
  .ZN({ S20391 })
);
NAND3_X1 #() 
NAND3_X1_3524_ (
  .A1({ S20387 }),
  .A2({ S25957[1237] }),
  .A3({ S20388 }),
  .ZN({ S20392 })
);
NAND3_X1 #() 
NAND3_X1_3525_ (
  .A1({ S20391 }),
  .A2({ S20392 }),
  .A3({ S25956[21] }),
  .ZN({ S20393 })
);
NAND2_X1 #() 
NAND2_X1_3347_ (
  .A1({ S20390 }),
  .A2({ S20393 }),
  .ZN({ S25957[1045] })
);
NOR2_X1 #() 
NOR2_X1_861_ (
  .A1({ S9034 }),
  .A2({ S9053 }),
  .ZN({ S25957[1204] })
);
OAI21_X1 #() 
OAI21_X1_1749_ (
  .A({ S25957[1163] }),
  .B1({ S20151 }),
  .B2({ S20177 }),
  .ZN({ S20394 })
);
NAND3_X1 #() 
NAND3_X1_3526_ (
  .A1({ S20143 }),
  .A2({ S20216 }),
  .A3({ S65 }),
  .ZN({ S20395 })
);
NAND3_X1 #() 
NAND3_X1_3527_ (
  .A1({ S20394 }),
  .A2({ S25957[1164] }),
  .A3({ S20395 }),
  .ZN({ S20396 })
);
NAND3_X1 #() 
NAND3_X1_3528_ (
  .A1({ S20160 }),
  .A2({ S25957[1163] }),
  .A3({ S20137 }),
  .ZN({ S20397 })
);
NAND2_X1 #() 
NAND2_X1_3348_ (
  .A1({ S20298 }),
  .A2({ S65 }),
  .ZN({ S20398 })
);
NAND3_X1 #() 
NAND3_X1_3529_ (
  .A1({ S20398 }),
  .A2({ S20131 }),
  .A3({ S20397 }),
  .ZN({ S20399 })
);
NAND3_X1 #() 
NAND3_X1_3530_ (
  .A1({ S20399 }),
  .A2({ S14483 }),
  .A3({ S20396 }),
  .ZN({ S20400 })
);
NAND2_X1 #() 
NAND2_X1_3349_ (
  .A1({ S20244 }),
  .A2({ S20161 }),
  .ZN({ S20401 })
);
AOI22_X1 #() 
AOI22_X1_385_ (
  .A1({ S20401 }),
  .A2({ S20148 }),
  .B1({ S20129 }),
  .B2({ S25957[1162] }),
  .ZN({ S20402 })
);
NAND4_X1 #() 
NAND4_X1_378_ (
  .A1({ S20148 }),
  .A2({ S20160 }),
  .A3({ S20155 }),
  .A4({ S25957[1163] }),
  .ZN({ S20403 })
);
OAI211_X1 #() 
OAI211_X1_1144_ (
  .A({ S20131 }),
  .B({ S20403 }),
  .C1({ S20402 }),
  .C2({ S25957[1163] }),
  .ZN({ S20404 })
);
NAND2_X1 #() 
NAND2_X1_3350_ (
  .A1({ S20148 }),
  .A2({ S25957[1162] }),
  .ZN({ S20405 })
);
NAND2_X1 #() 
NAND2_X1_3351_ (
  .A1({ S20405 }),
  .A2({ S20297 }),
  .ZN({ S20406 })
);
NAND2_X1 #() 
NAND2_X1_3352_ (
  .A1({ S20406 }),
  .A2({ S20163 }),
  .ZN({ S20407 })
);
AOI21_X1 #() 
AOI21_X1_1824_ (
  .A({ S14483 }),
  .B1({ S20407 }),
  .B2({ S25957[1164] }),
  .ZN({ S20408 })
);
NAND2_X1 #() 
NAND2_X1_3353_ (
  .A1({ S20408 }),
  .A2({ S20404 }),
  .ZN({ S20409 })
);
NAND3_X1 #() 
NAND3_X1_3531_ (
  .A1({ S20409 }),
  .A2({ S20400 }),
  .A3({ S20130 }),
  .ZN({ S20410 })
);
NAND3_X1 #() 
NAND3_X1_3532_ (
  .A1({ S20193 }),
  .A2({ S65 }),
  .A3({ S20144 }),
  .ZN({ S20411 })
);
NAND3_X1 #() 
NAND3_X1_3533_ (
  .A1({ S20228 }),
  .A2({ S20411 }),
  .A3({ S20131 }),
  .ZN({ S20412 })
);
OAI21_X1 #() 
OAI21_X1_1750_ (
  .A({ S65 }),
  .B1({ S20155 }),
  .B2({ S25957[1160] }),
  .ZN({ S20413 })
);
NAND3_X1 #() 
NAND3_X1_3534_ (
  .A1({ S20413 }),
  .A2({ S20372 }),
  .A3({ S25957[1164] }),
  .ZN({ S20414 })
);
NAND3_X1 #() 
NAND3_X1_3535_ (
  .A1({ S20414 }),
  .A2({ S20412 }),
  .A3({ S25957[1165] }),
  .ZN({ S20415 })
);
NAND2_X1 #() 
NAND2_X1_3354_ (
  .A1({ S20148 }),
  .A2({ S20193 }),
  .ZN({ S20416 })
);
NAND3_X1 #() 
NAND3_X1_3536_ (
  .A1({ S20136 }),
  .A2({ S20161 }),
  .A3({ S65 }),
  .ZN({ S20417 })
);
OAI211_X1 #() 
OAI211_X1_1145_ (
  .A({ S20417 }),
  .B({ S20131 }),
  .C1({ S20416 }),
  .C2({ S65 }),
  .ZN({ S20418 })
);
NAND3_X1 #() 
NAND3_X1_3537_ (
  .A1({ S20244 }),
  .A2({ S25957[1163] }),
  .A3({ S20137 }),
  .ZN({ S20419 })
);
NAND3_X1 #() 
NAND3_X1_3538_ (
  .A1({ S20338 }),
  .A2({ S20419 }),
  .A3({ S25957[1164] }),
  .ZN({ S20420 })
);
NAND3_X1 #() 
NAND3_X1_3539_ (
  .A1({ S20418 }),
  .A2({ S20420 }),
  .A3({ S14483 }),
  .ZN({ S20421 })
);
NAND3_X1 #() 
NAND3_X1_3540_ (
  .A1({ S20421 }),
  .A2({ S20415 }),
  .A3({ S25957[1166] }),
  .ZN({ S20422 })
);
NAND3_X1 #() 
NAND3_X1_3541_ (
  .A1({ S20410 }),
  .A2({ S25957[1167] }),
  .A3({ S20422 }),
  .ZN({ S20423 })
);
NAND4_X1 #() 
NAND4_X1_379_ (
  .A1({ S20150 }),
  .A2({ S20160 }),
  .A3({ S20161 }),
  .A4({ S65 }),
  .ZN({ S20424 })
);
NAND3_X1 #() 
NAND3_X1_3542_ (
  .A1({ S20169 }),
  .A2({ S20424 }),
  .A3({ S25957[1164] }),
  .ZN({ S20425 })
);
NOR2_X1 #() 
NOR2_X1_862_ (
  .A1({ S20193 }),
  .A2({ S20144 }),
  .ZN({ S20426 })
);
AOI21_X1 #() 
AOI21_X1_1825_ (
  .A({ S25957[1164] }),
  .B1({ S25957[1163] }),
  .B2({ S25957[1162] }),
  .ZN({ S20427 })
);
OAI21_X1 #() 
OAI21_X1_1751_ (
  .A({ S20427 }),
  .B1({ S20426 }),
  .B2({ S20251 }),
  .ZN({ S20428 })
);
NAND3_X1 #() 
NAND3_X1_3543_ (
  .A1({ S20425 }),
  .A2({ S20428 }),
  .A3({ S14483 }),
  .ZN({ S20429 })
);
NAND3_X1 #() 
NAND3_X1_3544_ (
  .A1({ S20182 }),
  .A2({ S65 }),
  .A3({ S25957[1162] }),
  .ZN({ S20430 })
);
NAND4_X1 #() 
NAND4_X1_380_ (
  .A1({ S20129 }),
  .A2({ S73 }),
  .A3({ S65 }),
  .A4({ S20138 }),
  .ZN({ S20431 })
);
NAND2_X1 #() 
NAND2_X1_3355_ (
  .A1({ S20431 }),
  .A2({ S20430 }),
  .ZN({ S20432 })
);
NAND2_X1 #() 
NAND2_X1_3356_ (
  .A1({ S20368 }),
  .A2({ S20131 }),
  .ZN({ S20433 })
);
INV_X1 #() 
INV_X1_1133_ (
  .A({ S120 }),
  .ZN({ S20434 })
);
OAI21_X1 #() 
OAI21_X1_1752_ (
  .A({ S25957[1164] }),
  .B1({ S20434 }),
  .B2({ S25957[1162] }),
  .ZN({ S20435 })
);
OAI211_X1 #() 
OAI211_X1_1146_ (
  .A({ S25957[1165] }),
  .B({ S20435 }),
  .C1({ S20432 }),
  .C2({ S20433 }),
  .ZN({ S20436 })
);
AOI21_X1 #() 
AOI21_X1_1826_ (
  .A({ S20130 }),
  .B1({ S20436 }),
  .B2({ S20429 }),
  .ZN({ S20437 })
);
NAND4_X1 #() 
NAND4_X1_381_ (
  .A1({ S20129 }),
  .A2({ S73 }),
  .A3({ S25957[1163] }),
  .A4({ S20138 }),
  .ZN({ S20438 })
);
NAND2_X1 #() 
NAND2_X1_3357_ (
  .A1({ S72 }),
  .A2({ S65 }),
  .ZN({ S20439 })
);
AND2_X1 #() 
AND2_X1_206_ (
  .A1({ S20439 }),
  .A2({ S20438 }),
  .ZN({ S20440 })
);
NAND3_X1 #() 
NAND3_X1_3545_ (
  .A1({ S20207 }),
  .A2({ S25957[1164] }),
  .A3({ S20430 }),
  .ZN({ S20441 })
);
OAI211_X1 #() 
OAI211_X1_1147_ (
  .A({ S25957[1165] }),
  .B({ S20441 }),
  .C1({ S20440 }),
  .C2({ S25957[1164] }),
  .ZN({ S20442 })
);
NAND4_X1 #() 
NAND4_X1_382_ (
  .A1({ S20132 }),
  .A2({ S20160 }),
  .A3({ S20193 }),
  .A4({ S25957[1163] }),
  .ZN({ S20443 })
);
NAND3_X1 #() 
NAND3_X1_3546_ (
  .A1({ S20443 }),
  .A2({ S25957[1164] }),
  .A3({ S20338 }),
  .ZN({ S20444 })
);
AOI22_X1 #() 
AOI22_X1_386_ (
  .A1({ S20162 }),
  .A2({ S65 }),
  .B1({ S20194 }),
  .B2({ S73 }),
  .ZN({ S20445 })
);
OAI211_X1 #() 
OAI211_X1_1148_ (
  .A({ S14483 }),
  .B({ S20444 }),
  .C1({ S20445 }),
  .C2({ S25957[1164] }),
  .ZN({ S20446 })
);
AND3_X1 #() 
AND3_X1_129_ (
  .A1({ S20442 }),
  .A2({ S20446 }),
  .A3({ S20130 }),
  .ZN({ S20447 })
);
OAI21_X1 #() 
OAI21_X1_1753_ (
  .A({ S20192 }),
  .B1({ S20447 }),
  .B2({ S20437 }),
  .ZN({ S20448 })
);
NAND3_X1 #() 
NAND3_X1_3547_ (
  .A1({ S20448 }),
  .A2({ S20423 }),
  .A3({ S9002 }),
  .ZN({ S20449 })
);
AOI21_X1 #() 
AOI21_X1_1827_ (
  .A({ S25957[1163] }),
  .B1({ S20297 }),
  .B2({ S20216 }),
  .ZN({ S20450 })
);
NOR2_X1 #() 
NOR2_X1_863_ (
  .A1({ S20450 }),
  .A2({ S25957[1164] }),
  .ZN({ S20451 })
);
AOI21_X1 #() 
AOI21_X1_1828_ (
  .A({ S25957[1165] }),
  .B1({ S20451 }),
  .B2({ S20397 }),
  .ZN({ S20452 })
);
AOI22_X1 #() 
AOI22_X1_387_ (
  .A1({ S20452 }),
  .A2({ S20396 }),
  .B1({ S20404 }),
  .B2({ S20408 }),
  .ZN({ S20453 })
);
NAND2_X1 #() 
NAND2_X1_3358_ (
  .A1({ S20422 }),
  .A2({ S25957[1167] }),
  .ZN({ S20454 })
);
AOI21_X1 #() 
AOI21_X1_1829_ (
  .A({ S20454 }),
  .B1({ S20453 }),
  .B2({ S20130 }),
  .ZN({ S20455 })
);
NAND2_X1 #() 
NAND2_X1_3359_ (
  .A1({ S20436 }),
  .A2({ S20429 }),
  .ZN({ S20456 })
);
NAND2_X1 #() 
NAND2_X1_3360_ (
  .A1({ S20456 }),
  .A2({ S25957[1166] }),
  .ZN({ S20457 })
);
NAND3_X1 #() 
NAND3_X1_3548_ (
  .A1({ S20442 }),
  .A2({ S20446 }),
  .A3({ S20130 }),
  .ZN({ S20458 })
);
AOI21_X1 #() 
AOI21_X1_1830_ (
  .A({ S25957[1167] }),
  .B1({ S20457 }),
  .B2({ S20458 }),
  .ZN({ S20459 })
);
OAI21_X1 #() 
OAI21_X1_1754_ (
  .A({ S25957[1268] }),
  .B1({ S20455 }),
  .B2({ S20459 }),
  .ZN({ S20460 })
);
NAND3_X1 #() 
NAND3_X1_3549_ (
  .A1({ S20460 }),
  .A2({ S20449 }),
  .A3({ S9075 }),
  .ZN({ S20461 })
);
OAI21_X1 #() 
OAI21_X1_1755_ (
  .A({ S9002 }),
  .B1({ S20455 }),
  .B2({ S20459 }),
  .ZN({ S20462 })
);
NAND3_X1 #() 
NAND3_X1_3550_ (
  .A1({ S20448 }),
  .A2({ S20423 }),
  .A3({ S25957[1268] }),
  .ZN({ S20463 })
);
NAND3_X1 #() 
NAND3_X1_3551_ (
  .A1({ S20462 }),
  .A2({ S20463 }),
  .A3({ S25957[1236] }),
  .ZN({ S20464 })
);
AOI21_X1 #() 
AOI21_X1_1831_ (
  .A({ S25957[1204] }),
  .B1({ S20461 }),
  .B2({ S20464 }),
  .ZN({ S20465 })
);
AND3_X1 #() 
AND3_X1_130_ (
  .A1({ S20464 }),
  .A2({ S20461 }),
  .A3({ S25957[1204] }),
  .ZN({ S20466 })
);
OAI21_X1 #() 
OAI21_X1_1756_ (
  .A({ S25957[1172] }),
  .B1({ S20466 }),
  .B2({ S20465 }),
  .ZN({ S20467 })
);
INV_X1 #() 
INV_X1_1134_ (
  .A({ S25957[1204] }),
  .ZN({ S20468 })
);
AOI21_X1 #() 
AOI21_X1_1832_ (
  .A({ S25957[1236] }),
  .B1({ S20462 }),
  .B2({ S20463 }),
  .ZN({ S20469 })
);
AOI21_X1 #() 
AOI21_X1_1833_ (
  .A({ S9075 }),
  .B1({ S20460 }),
  .B2({ S20449 }),
  .ZN({ S20470 })
);
OAI21_X1 #() 
OAI21_X1_1757_ (
  .A({ S20468 }),
  .B1({ S20469 }),
  .B2({ S20470 }),
  .ZN({ S20471 })
);
NAND3_X1 #() 
NAND3_X1_3552_ (
  .A1({ S20461 }),
  .A2({ S20464 }),
  .A3({ S25957[1204] }),
  .ZN({ S20472 })
);
NAND3_X1 #() 
NAND3_X1_3553_ (
  .A1({ S20471 }),
  .A2({ S9119 }),
  .A3({ S20472 }),
  .ZN({ S20473 })
);
NAND2_X1 #() 
NAND2_X1_3361_ (
  .A1({ S20467 }),
  .A2({ S20473 }),
  .ZN({ S25957[1044] })
);
NOR2_X1 #() 
NOR2_X1_864_ (
  .A1({ S9713 }),
  .A2({ S9724 }),
  .ZN({ S25957[1203] })
);
NAND2_X1 #() 
NAND2_X1_3362_ (
  .A1({ S9681 }),
  .A2({ S9692 }),
  .ZN({ S25957[1235] })
);
NAND3_X1 #() 
NAND3_X1_3554_ (
  .A1({ S20180 }),
  .A2({ S65 }),
  .A3({ S20148 }),
  .ZN({ S20474 })
);
NAND3_X1 #() 
NAND3_X1_3555_ (
  .A1({ S20405 }),
  .A2({ S20297 }),
  .A3({ S25957[1163] }),
  .ZN({ S20475 })
);
AOI21_X1 #() 
AOI21_X1_1834_ (
  .A({ S25957[1164] }),
  .B1({ S20475 }),
  .B2({ S20474 }),
  .ZN({ S20476 })
);
NAND3_X1 #() 
NAND3_X1_3556_ (
  .A1({ S73 }),
  .A2({ S20160 }),
  .A3({ S25957[1163] }),
  .ZN({ S20477 })
);
NAND3_X1 #() 
NAND3_X1_3557_ (
  .A1({ S20216 }),
  .A2({ S65 }),
  .A3({ S20148 }),
  .ZN({ S20478 })
);
NAND3_X1 #() 
NAND3_X1_3558_ (
  .A1({ S20478 }),
  .A2({ S25957[1164] }),
  .A3({ S20477 }),
  .ZN({ S20479 })
);
NAND2_X1 #() 
NAND2_X1_3363_ (
  .A1({ S20479 }),
  .A2({ S25957[1165] }),
  .ZN({ S20480 })
);
NAND3_X1 #() 
NAND3_X1_3559_ (
  .A1({ S20183 }),
  .A2({ S65 }),
  .A3({ S20139 }),
  .ZN({ S20481 })
);
AOI21_X1 #() 
AOI21_X1_1835_ (
  .A({ S20131 }),
  .B1({ S20481 }),
  .B2({ S20325 }),
  .ZN({ S20482 })
);
NAND2_X1 #() 
NAND2_X1_3364_ (
  .A1({ S20427 }),
  .A2({ S20280 }),
  .ZN({ S20483 })
);
NAND2_X1 #() 
NAND2_X1_3365_ (
  .A1({ S20483 }),
  .A2({ S14483 }),
  .ZN({ S20484 })
);
OAI22_X1 #() 
OAI22_X1_95_ (
  .A1({ S20480 }),
  .A2({ S20476 }),
  .B1({ S20482 }),
  .B2({ S20484 }),
  .ZN({ S20485 })
);
AND2_X1 #() 
AND2_X1_207_ (
  .A1({ S20485 }),
  .A2({ S25957[1166] }),
  .ZN({ S20486 })
);
AOI22_X1 #() 
AOI22_X1_388_ (
  .A1({ S20223 }),
  .A2({ S20331 }),
  .B1({ S20280 }),
  .B2({ S65 }),
  .ZN({ S20487 })
);
NAND4_X1 #() 
NAND4_X1_383_ (
  .A1({ S20319 }),
  .A2({ S20417 }),
  .A3({ S25957[1164] }),
  .A4({ S20163 }),
  .ZN({ S20488 })
);
OAI211_X1 #() 
OAI211_X1_1149_ (
  .A({ S14483 }),
  .B({ S20488 }),
  .C1({ S20487 }),
  .C2({ S25957[1164] }),
  .ZN({ S20489 })
);
NAND2_X1 #() 
NAND2_X1_3366_ (
  .A1({ S20161 }),
  .A2({ S65 }),
  .ZN({ S20490 })
);
NAND4_X1 #() 
NAND4_X1_384_ (
  .A1({ S20136 }),
  .A2({ S20244 }),
  .A3({ S25957[1163] }),
  .A4({ S25957[1161] }),
  .ZN({ S20491 })
);
OAI211_X1 #() 
OAI211_X1_1150_ (
  .A({ S20131 }),
  .B({ S20491 }),
  .C1({ S20218 }),
  .C2({ S20490 }),
  .ZN({ S20492 })
);
NAND2_X1 #() 
NAND2_X1_3367_ (
  .A1({ S20145 }),
  .A2({ S25957[1163] }),
  .ZN({ S20493 })
);
NAND3_X1 #() 
NAND3_X1_3560_ (
  .A1({ S20217 }),
  .A2({ S65 }),
  .A3({ S20132 }),
  .ZN({ S20494 })
);
OAI211_X1 #() 
OAI211_X1_1151_ (
  .A({ S20494 }),
  .B({ S25957[1164] }),
  .C1({ S20493 }),
  .C2({ S20335 }),
  .ZN({ S20495 })
);
NAND3_X1 #() 
NAND3_X1_3561_ (
  .A1({ S20495 }),
  .A2({ S20492 }),
  .A3({ S25957[1165] }),
  .ZN({ S20496 })
);
AND2_X1 #() 
AND2_X1_208_ (
  .A1({ S20496 }),
  .A2({ S20489 }),
  .ZN({ S20497 })
);
OAI21_X1 #() 
OAI21_X1_1758_ (
  .A({ S25957[1167] }),
  .B1({ S20497 }),
  .B2({ S25957[1166] }),
  .ZN({ S20498 })
);
OAI211_X1 #() 
OAI211_X1_1152_ (
  .A({ S20275 }),
  .B({ S25957[1164] }),
  .C1({ S20218 }),
  .C2({ S20219 }),
  .ZN({ S20499 })
);
INV_X1 #() 
INV_X1_1135_ (
  .A({ S20499 }),
  .ZN({ S20500 })
);
NAND3_X1 #() 
NAND3_X1_3562_ (
  .A1({ S20150 }),
  .A2({ S25957[1163] }),
  .A3({ S20144 }),
  .ZN({ S20501 })
);
OAI21_X1 #() 
OAI21_X1_1759_ (
  .A({ S20501 }),
  .B1({ S20416 }),
  .B2({ S25957[1163] }),
  .ZN({ S20502 })
);
OAI21_X1 #() 
OAI21_X1_1760_ (
  .A({ S25957[1165] }),
  .B1({ S20502 }),
  .B2({ S25957[1164] }),
  .ZN({ S20503 })
);
NAND4_X1 #() 
NAND4_X1_385_ (
  .A1({ S20193 }),
  .A2({ S20155 }),
  .A3({ S65 }),
  .A4({ S25957[1160] }),
  .ZN({ S20504 })
);
AOI21_X1 #() 
AOI21_X1_1836_ (
  .A({ S25957[1164] }),
  .B1({ S20140 }),
  .B2({ S20504 }),
  .ZN({ S20505 })
);
NAND2_X1 #() 
NAND2_X1_3368_ (
  .A1({ S20160 }),
  .A2({ S65 }),
  .ZN({ S20506 })
);
NOR3_X1 #() 
NOR3_X1_120_ (
  .A1({ S20506 }),
  .A2({ S72 }),
  .A3({ S20131 }),
  .ZN({ S20507 })
);
OAI21_X1 #() 
OAI21_X1_1761_ (
  .A({ S14483 }),
  .B1({ S20505 }),
  .B2({ S20507 }),
  .ZN({ S20508 })
);
OAI211_X1 #() 
OAI211_X1_1153_ (
  .A({ S20508 }),
  .B({ S25957[1166] }),
  .C1({ S20500 }),
  .C2({ S20503 }),
  .ZN({ S20509 })
);
OAI21_X1 #() 
OAI21_X1_1762_ (
  .A({ S73 }),
  .B1({ S20129 }),
  .B2({ S25957[1162] }),
  .ZN({ S20510 })
);
OAI211_X1 #() 
OAI211_X1_1154_ (
  .A({ S20362 }),
  .B({ S25957[1164] }),
  .C1({ S20510 }),
  .C2({ S65 }),
  .ZN({ S20511 })
);
NAND2_X1 #() 
NAND2_X1_3369_ (
  .A1({ S25957[1163] }),
  .A2({ S25957[1162] }),
  .ZN({ S20512 })
);
OAI211_X1 #() 
OAI211_X1_1155_ (
  .A({ S20272 }),
  .B({ S20131 }),
  .C1({ S20144 }),
  .C2({ S20512 }),
  .ZN({ S20513 })
);
OAI21_X1 #() 
OAI21_X1_1763_ (
  .A({ S20511 }),
  .B1({ S20199 }),
  .B2({ S20513 }),
  .ZN({ S20514 })
);
NAND3_X1 #() 
NAND3_X1_3563_ (
  .A1({ S20148 }),
  .A2({ S20160 }),
  .A3({ S65 }),
  .ZN({ S20515 })
);
NAND4_X1 #() 
NAND4_X1_386_ (
  .A1({ S20515 }),
  .A2({ S20322 }),
  .A3({ S20156 }),
  .A4({ S20131 }),
  .ZN({ S20516 })
);
NAND2_X1 #() 
NAND2_X1_3370_ (
  .A1({ S20493 }),
  .A2({ S25957[1164] }),
  .ZN({ S20517 })
);
OAI211_X1 #() 
OAI211_X1_1156_ (
  .A({ S25957[1165] }),
  .B({ S20516 }),
  .C1({ S20213 }),
  .C2({ S20517 }),
  .ZN({ S20518 })
);
OAI211_X1 #() 
OAI211_X1_1157_ (
  .A({ S20518 }),
  .B({ S20130 }),
  .C1({ S20514 }),
  .C2({ S25957[1165] }),
  .ZN({ S20519 })
);
NAND3_X1 #() 
NAND3_X1_3564_ (
  .A1({ S20509 }),
  .A2({ S20519 }),
  .A3({ S20192 }),
  .ZN({ S20520 })
);
OAI211_X1 #() 
OAI211_X1_1158_ (
  .A({ S20520 }),
  .B({ S25957[1267] }),
  .C1({ S20498 }),
  .C2({ S20486 }),
  .ZN({ S20521 })
);
INV_X1 #() 
INV_X1_1136_ (
  .A({ S25957[1267] }),
  .ZN({ S20522 })
);
NAND3_X1 #() 
NAND3_X1_3565_ (
  .A1({ S20496 }),
  .A2({ S20489 }),
  .A3({ S20130 }),
  .ZN({ S20523 })
);
OAI211_X1 #() 
OAI211_X1_1159_ (
  .A({ S20523 }),
  .B({ S25957[1167] }),
  .C1({ S20485 }),
  .C2({ S20130 }),
  .ZN({ S20524 })
);
AOI22_X1 #() 
AOI22_X1_389_ (
  .A1({ S20330 }),
  .A2({ S20331 }),
  .B1({ S20274 }),
  .B2({ S25957[1163] }),
  .ZN({ S20525 })
);
NAND2_X1 #() 
NAND2_X1_3371_ (
  .A1({ S20502 }),
  .A2({ S20131 }),
  .ZN({ S20526 })
);
OAI211_X1 #() 
OAI211_X1_1160_ (
  .A({ S25957[1165] }),
  .B({ S20526 }),
  .C1({ S20525 }),
  .C2({ S20131 }),
  .ZN({ S20527 })
);
NAND2_X1 #() 
NAND2_X1_3372_ (
  .A1({ S20197 }),
  .A2({ S20443 }),
  .ZN({ S20528 })
);
NOR2_X1 #() 
NOR2_X1_865_ (
  .A1({ S20507 }),
  .A2({ S25957[1165] }),
  .ZN({ S20529 })
);
NAND2_X1 #() 
NAND2_X1_3373_ (
  .A1({ S20529 }),
  .A2({ S20528 }),
  .ZN({ S20530 })
);
NAND3_X1 #() 
NAND3_X1_3566_ (
  .A1({ S20527 }),
  .A2({ S20530 }),
  .A3({ S25957[1166] }),
  .ZN({ S20531 })
);
OAI21_X1 #() 
OAI21_X1_1764_ (
  .A({ S20518 }),
  .B1({ S20514 }),
  .B2({ S25957[1165] }),
  .ZN({ S20532 })
);
NAND2_X1 #() 
NAND2_X1_3374_ (
  .A1({ S20532 }),
  .A2({ S20130 }),
  .ZN({ S20533 })
);
NAND3_X1 #() 
NAND3_X1_3567_ (
  .A1({ S20533 }),
  .A2({ S20531 }),
  .A3({ S20192 }),
  .ZN({ S20534 })
);
NAND3_X1 #() 
NAND3_X1_3568_ (
  .A1({ S20534 }),
  .A2({ S20524 }),
  .A3({ S20522 }),
  .ZN({ S20535 })
);
NAND3_X1 #() 
NAND3_X1_3569_ (
  .A1({ S20521 }),
  .A2({ S20535 }),
  .A3({ S25957[1235] }),
  .ZN({ S20536 })
);
INV_X1 #() 
INV_X1_1137_ (
  .A({ S25957[1235] }),
  .ZN({ S20537 })
);
NAND3_X1 #() 
NAND3_X1_3570_ (
  .A1({ S20534 }),
  .A2({ S20524 }),
  .A3({ S25957[1267] }),
  .ZN({ S20538 })
);
OAI211_X1 #() 
OAI211_X1_1161_ (
  .A({ S20520 }),
  .B({ S20522 }),
  .C1({ S20498 }),
  .C2({ S20486 }),
  .ZN({ S20539 })
);
NAND3_X1 #() 
NAND3_X1_3571_ (
  .A1({ S20539 }),
  .A2({ S20538 }),
  .A3({ S20537 }),
  .ZN({ S20540 })
);
NAND3_X1 #() 
NAND3_X1_3572_ (
  .A1({ S20536 }),
  .A2({ S20540 }),
  .A3({ S25957[1203] }),
  .ZN({ S20541 })
);
INV_X1 #() 
INV_X1_1138_ (
  .A({ S25957[1203] }),
  .ZN({ S20542 })
);
NAND3_X1 #() 
NAND3_X1_3573_ (
  .A1({ S20521 }),
  .A2({ S20535 }),
  .A3({ S20537 }),
  .ZN({ S20543 })
);
NAND3_X1 #() 
NAND3_X1_3574_ (
  .A1({ S20539 }),
  .A2({ S20538 }),
  .A3({ S25957[1235] }),
  .ZN({ S20544 })
);
NAND3_X1 #() 
NAND3_X1_3575_ (
  .A1({ S20543 }),
  .A2({ S20544 }),
  .A3({ S20542 }),
  .ZN({ S20545 })
);
NAND3_X1 #() 
NAND3_X1_3576_ (
  .A1({ S20541 }),
  .A2({ S20545 }),
  .A3({ S25957[1171] }),
  .ZN({ S20546 })
);
NAND3_X1 #() 
NAND3_X1_3577_ (
  .A1({ S20536 }),
  .A2({ S20540 }),
  .A3({ S20542 }),
  .ZN({ S20547 })
);
NAND3_X1 #() 
NAND3_X1_3578_ (
  .A1({ S20543 }),
  .A2({ S20544 }),
  .A3({ S25957[1203] }),
  .ZN({ S20548 })
);
NAND3_X1 #() 
NAND3_X1_3579_ (
  .A1({ S20547 }),
  .A2({ S20548 }),
  .A3({ S50 }),
  .ZN({ S20549 })
);
NAND2_X1 #() 
NAND2_X1_3375_ (
  .A1({ S20546 }),
  .A2({ S20549 }),
  .ZN({ S74 })
);
AND2_X1 #() 
AND2_X1_209_ (
  .A1({ S20549 }),
  .A2({ S20546 }),
  .ZN({ S25957[1043] })
);
INV_X1 #() 
INV_X1_1139_ (
  .A({ S25957[1264] }),
  .ZN({ S20550 })
);
AOI21_X1 #() 
AOI21_X1_1837_ (
  .A({ S25957[1163] }),
  .B1({ S20243 }),
  .B2({ S20332 }),
  .ZN({ S20551 })
);
NAND3_X1 #() 
NAND3_X1_3580_ (
  .A1({ S20182 }),
  .A2({ S25957[1163] }),
  .A3({ S25957[1162] }),
  .ZN({ S20552 })
);
INV_X1 #() 
INV_X1_1140_ (
  .A({ S20552 }),
  .ZN({ S20553 })
);
OAI21_X1 #() 
OAI21_X1_1765_ (
  .A({ S25957[1164] }),
  .B1({ S20551 }),
  .B2({ S20553 }),
  .ZN({ S20554 })
);
AOI21_X1 #() 
AOI21_X1_1838_ (
  .A({ S25957[1164] }),
  .B1({ S20196 }),
  .B2({ S20158 }),
  .ZN({ S20555 })
);
NAND2_X1 #() 
NAND2_X1_3376_ (
  .A1({ S20555 }),
  .A2({ S20140 }),
  .ZN({ S20556 })
);
AOI21_X1 #() 
AOI21_X1_1839_ (
  .A({ S14483 }),
  .B1({ S20554 }),
  .B2({ S20556 }),
  .ZN({ S20557 })
);
NOR2_X1 #() 
NOR2_X1_866_ (
  .A1({ S20160 }),
  .A2({ S25957[1161] }),
  .ZN({ S20558 })
);
NAND4_X1 #() 
NAND4_X1_387_ (
  .A1({ S20148 }),
  .A2({ S20182 }),
  .A3({ S25957[1163] }),
  .A4({ S25957[1162] }),
  .ZN({ S20559 })
);
OAI211_X1 #() 
OAI211_X1_1162_ (
  .A({ S20559 }),
  .B({ S25957[1164] }),
  .C1({ S20351 }),
  .C2({ S20558 }),
  .ZN({ S20560 })
);
NAND3_X1 #() 
NAND3_X1_3581_ (
  .A1({ S20368 }),
  .A2({ S20351 }),
  .A3({ S20131 }),
  .ZN({ S20561 })
);
AND3_X1 #() 
AND3_X1_131_ (
  .A1({ S20560 }),
  .A2({ S14483 }),
  .A3({ S20561 }),
  .ZN({ S20562 })
);
OAI21_X1 #() 
OAI21_X1_1766_ (
  .A({ S25957[1166] }),
  .B1({ S20557 }),
  .B2({ S20562 }),
  .ZN({ S20563 })
);
NOR2_X1 #() 
NOR2_X1_867_ (
  .A1({ S20506 }),
  .A2({ S72 }),
  .ZN({ S20564 })
);
NAND3_X1 #() 
NAND3_X1_3582_ (
  .A1({ S20150 }),
  .A2({ S65 }),
  .A3({ S20144 }),
  .ZN({ S20565 })
);
OAI21_X1 #() 
OAI21_X1_1767_ (
  .A({ S20565 }),
  .B1({ S20564 }),
  .B2({ S20271 }),
  .ZN({ S20566 })
);
NAND2_X1 #() 
NAND2_X1_3377_ (
  .A1({ S20403 }),
  .A2({ S20413 }),
  .ZN({ S20567 })
);
NAND2_X1 #() 
NAND2_X1_3378_ (
  .A1({ S20567 }),
  .A2({ S20131 }),
  .ZN({ S20568 })
);
OAI211_X1 #() 
OAI211_X1_1163_ (
  .A({ S25957[1165] }),
  .B({ S20568 }),
  .C1({ S20566 }),
  .C2({ S20131 }),
  .ZN({ S20569 })
);
NAND4_X1 #() 
NAND4_X1_388_ (
  .A1({ S20132 }),
  .A2({ S20160 }),
  .A3({ S20155 }),
  .A4({ S65 }),
  .ZN({ S20570 })
);
NAND2_X1 #() 
NAND2_X1_3379_ (
  .A1({ S20570 }),
  .A2({ S20501 }),
  .ZN({ S20571 })
);
AOI22_X1 #() 
AOI22_X1_390_ (
  .A1({ S20571 }),
  .A2({ S20131 }),
  .B1({ S20267 }),
  .B2({ S20431 }),
  .ZN({ S20572 })
);
AOI21_X1 #() 
AOI21_X1_1840_ (
  .A({ S25957[1166] }),
  .B1({ S20572 }),
  .B2({ S14483 }),
  .ZN({ S20573 })
);
NAND2_X1 #() 
NAND2_X1_3380_ (
  .A1({ S20573 }),
  .A2({ S20569 }),
  .ZN({ S20574 })
);
AOI21_X1 #() 
AOI21_X1_1841_ (
  .A({ S20192 }),
  .B1({ S20563 }),
  .B2({ S20574 }),
  .ZN({ S20575 })
);
NAND2_X1 #() 
NAND2_X1_3381_ (
  .A1({ S20193 }),
  .A2({ S65 }),
  .ZN({ S20576 })
);
NOR2_X1 #() 
NOR2_X1_868_ (
  .A1({ S20218 }),
  .A2({ S20576 }),
  .ZN({ S20577 })
);
NAND3_X1 #() 
NAND3_X1_3583_ (
  .A1({ S20319 }),
  .A2({ S25957[1164] }),
  .A3({ S20163 }),
  .ZN({ S20578 })
);
NOR2_X1 #() 
NOR2_X1_869_ (
  .A1({ S20577 }),
  .A2({ S20578 }),
  .ZN({ S20579 })
);
AOI21_X1 #() 
AOI21_X1_1842_ (
  .A({ S25957[1163] }),
  .B1({ S20139 }),
  .B2({ S20145 }),
  .ZN({ S20580 })
);
NAND4_X1 #() 
NAND4_X1_389_ (
  .A1({ S20182 }),
  .A2({ S20148 }),
  .A3({ S20193 }),
  .A4({ S25957[1163] }),
  .ZN({ S20581 })
);
NAND2_X1 #() 
NAND2_X1_3382_ (
  .A1({ S20581 }),
  .A2({ S20131 }),
  .ZN({ S20582 })
);
OAI21_X1 #() 
OAI21_X1_1768_ (
  .A({ S14483 }),
  .B1({ S20582 }),
  .B2({ S20580 }),
  .ZN({ S20583 })
);
NAND3_X1 #() 
NAND3_X1_3584_ (
  .A1({ S20355 }),
  .A2({ S20245 }),
  .A3({ S20131 }),
  .ZN({ S20584 })
);
NAND3_X1 #() 
NAND3_X1_3585_ (
  .A1({ S20365 }),
  .A2({ S20477 }),
  .A3({ S25957[1164] }),
  .ZN({ S20585 })
);
NAND3_X1 #() 
NAND3_X1_3586_ (
  .A1({ S20584 }),
  .A2({ S20585 }),
  .A3({ S25957[1165] }),
  .ZN({ S20586 })
);
OAI211_X1 #() 
OAI211_X1_1164_ (
  .A({ S20130 }),
  .B({ S20586 }),
  .C1({ S20579 }),
  .C2({ S20583 }),
  .ZN({ S20587 })
);
NAND2_X1 #() 
NAND2_X1_3383_ (
  .A1({ S20160 }),
  .A2({ S20137 }),
  .ZN({ S20588 })
);
NAND2_X1 #() 
NAND2_X1_3384_ (
  .A1({ S20588 }),
  .A2({ S65 }),
  .ZN({ S20589 })
);
INV_X1 #() 
INV_X1_1141_ (
  .A({ S20589 }),
  .ZN({ S20590 })
);
NAND4_X1 #() 
NAND4_X1_390_ (
  .A1({ S20322 }),
  .A2({ S20260 }),
  .A3({ S20155 }),
  .A4({ S25957[1164] }),
  .ZN({ S20591 })
);
OAI211_X1 #() 
OAI211_X1_1165_ (
  .A({ S14483 }),
  .B({ S20591 }),
  .C1({ S20590 }),
  .C2({ S20433 }),
  .ZN({ S20592 })
);
NOR2_X1 #() 
NOR2_X1_870_ (
  .A1({ S20341 }),
  .A2({ S25957[1164] }),
  .ZN({ S20593 })
);
NAND4_X1 #() 
NAND4_X1_391_ (
  .A1({ S20588 }),
  .A2({ S20348 }),
  .A3({ S20132 }),
  .A4({ S25957[1163] }),
  .ZN({ S20594 })
);
AOI21_X1 #() 
AOI21_X1_1843_ (
  .A({ S20131 }),
  .B1({ S20180 }),
  .B2({ S65 }),
  .ZN({ S20595 })
);
AOI22_X1 #() 
AOI22_X1_391_ (
  .A1({ S20299 }),
  .A2({ S20593 }),
  .B1({ S20594 }),
  .B2({ S20595 }),
  .ZN({ S20596 })
);
OAI211_X1 #() 
OAI211_X1_1166_ (
  .A({ S20592 }),
  .B({ S25957[1166] }),
  .C1({ S20596 }),
  .C2({ S14483 }),
  .ZN({ S20597 })
);
AND3_X1 #() 
AND3_X1_132_ (
  .A1({ S20597 }),
  .A2({ S20587 }),
  .A3({ S20192 }),
  .ZN({ S20598 })
);
OAI21_X1 #() 
OAI21_X1_1769_ (
  .A({ S20550 }),
  .B1({ S20575 }),
  .B2({ S20598 }),
  .ZN({ S20599 })
);
NAND2_X1 #() 
NAND2_X1_3385_ (
  .A1({ S73 }),
  .A2({ S20138 }),
  .ZN({ S20600 })
);
NAND3_X1 #() 
NAND3_X1_3587_ (
  .A1({ S20600 }),
  .A2({ S65 }),
  .A3({ S20145 }),
  .ZN({ S20601 })
);
NAND2_X1 #() 
NAND2_X1_3386_ (
  .A1({ S20601 }),
  .A2({ S20552 }),
  .ZN({ S20602 })
);
AOI22_X1 #() 
AOI22_X1_392_ (
  .A1({ S20602 }),
  .A2({ S25957[1164] }),
  .B1({ S20555 }),
  .B2({ S20140 }),
  .ZN({ S20603 })
);
NAND3_X1 #() 
NAND3_X1_3588_ (
  .A1({ S20560 }),
  .A2({ S14483 }),
  .A3({ S20561 }),
  .ZN({ S20604 })
);
OAI21_X1 #() 
OAI21_X1_1770_ (
  .A({ S20604 }),
  .B1({ S20603 }),
  .B2({ S14483 }),
  .ZN({ S20605 })
);
AOI22_X1 #() 
AOI22_X1_393_ (
  .A1({ S20605 }),
  .A2({ S25957[1166] }),
  .B1({ S20569 }),
  .B2({ S20573 }),
  .ZN({ S20606 })
);
NAND3_X1 #() 
NAND3_X1_3589_ (
  .A1({ S20597 }),
  .A2({ S20587 }),
  .A3({ S20192 }),
  .ZN({ S20607 })
);
OAI211_X1 #() 
OAI211_X1_1167_ (
  .A({ S25957[1264] }),
  .B({ S20607 }),
  .C1({ S20606 }),
  .C2({ S20192 }),
  .ZN({ S20608 })
);
AOI21_X1 #() 
AOI21_X1_1844_ (
  .A({ S25956[48] }),
  .B1({ S20599 }),
  .B2({ S20608 }),
  .ZN({ S20609 })
);
OAI21_X1 #() 
OAI21_X1_1771_ (
  .A({ S25957[1264] }),
  .B1({ S20575 }),
  .B2({ S20598 }),
  .ZN({ S20610 })
);
OAI211_X1 #() 
OAI211_X1_1168_ (
  .A({ S20550 }),
  .B({ S20607 }),
  .C1({ S20606 }),
  .C2({ S20192 }),
  .ZN({ S20611 })
);
AOI21_X1 #() 
AOI21_X1_1845_ (
  .A({ S9792 }),
  .B1({ S20610 }),
  .B2({ S20611 }),
  .ZN({ S20612 })
);
OAI21_X1 #() 
OAI21_X1_1772_ (
  .A({ S25957[1168] }),
  .B1({ S20609 }),
  .B2({ S20612 }),
  .ZN({ S20613 })
);
OAI21_X1 #() 
OAI21_X1_1773_ (
  .A({ S10390 }),
  .B1({ S10357 }),
  .B2({ S10368 }),
  .ZN({ S20614 })
);
NAND3_X1 #() 
NAND3_X1_3590_ (
  .A1({ S10407 }),
  .A2({ S25956[16] }),
  .A3({ S10346 }),
  .ZN({ S20615 })
);
NAND2_X1 #() 
NAND2_X1_3387_ (
  .A1({ S20614 }),
  .A2({ S20615 }),
  .ZN({ S20616 })
);
NAND3_X1 #() 
NAND3_X1_3591_ (
  .A1({ S20610 }),
  .A2({ S20611 }),
  .A3({ S9792 }),
  .ZN({ S20617 })
);
NAND3_X1 #() 
NAND3_X1_3592_ (
  .A1({ S20599 }),
  .A2({ S20608 }),
  .A3({ S25956[48] }),
  .ZN({ S20618 })
);
NAND3_X1 #() 
NAND3_X1_3593_ (
  .A1({ S20617 }),
  .A2({ S20618 }),
  .A3({ S20616 }),
  .ZN({ S20619 })
);
NAND2_X1 #() 
NAND2_X1_3388_ (
  .A1({ S20613 }),
  .A2({ S20619 }),
  .ZN({ S25957[1040] })
);
NOR2_X1 #() 
NOR2_X1_871_ (
  .A1({ S10895 }),
  .A2({ S10904 }),
  .ZN({ S25957[1201] })
);
INV_X1 #() 
INV_X1_1142_ (
  .A({ S25957[1201] }),
  .ZN({ S20620 })
);
NAND2_X1 #() 
NAND2_X1_3389_ (
  .A1({ S10862 }),
  .A2({ S10873 }),
  .ZN({ S25957[1233] })
);
INV_X1 #() 
INV_X1_1143_ (
  .A({ S25957[1233] }),
  .ZN({ S20621 })
);
AOI21_X1 #() 
AOI21_X1_1846_ (
  .A({ S65 }),
  .B1({ S20183 }),
  .B2({ S20132 }),
  .ZN({ S20622 })
);
OAI211_X1 #() 
OAI211_X1_1169_ (
  .A({ S20319 }),
  .B({ S20131 }),
  .C1({ S20149 }),
  .C2({ S20576 }),
  .ZN({ S20623 })
);
OAI21_X1 #() 
OAI21_X1_1774_ (
  .A({ S20623 }),
  .B1({ S20622 }),
  .B2({ S20206 }),
  .ZN({ S20624 })
);
NAND2_X1 #() 
NAND2_X1_3390_ (
  .A1({ S20624 }),
  .A2({ S25957[1165] }),
  .ZN({ S20625 })
);
NOR2_X1 #() 
NOR2_X1_872_ (
  .A1({ S20141 }),
  .A2({ S20133 }),
  .ZN({ S20626 })
);
NAND2_X1 #() 
NAND2_X1_3391_ (
  .A1({ S20177 }),
  .A2({ S65 }),
  .ZN({ S20627 })
);
NAND2_X1 #() 
NAND2_X1_3392_ (
  .A1({ S20290 }),
  .A2({ S20627 }),
  .ZN({ S20628 })
);
OAI21_X1 #() 
OAI21_X1_1775_ (
  .A({ S25957[1164] }),
  .B1({ S20628 }),
  .B2({ S20626 }),
  .ZN({ S20629 })
);
OAI21_X1 #() 
OAI21_X1_1776_ (
  .A({ S20131 }),
  .B1({ S20201 }),
  .B2({ S20450 }),
  .ZN({ S20630 })
);
NAND3_X1 #() 
NAND3_X1_3594_ (
  .A1({ S20630 }),
  .A2({ S20629 }),
  .A3({ S14483 }),
  .ZN({ S20631 })
);
AOI21_X1 #() 
AOI21_X1_1847_ (
  .A({ S25957[1166] }),
  .B1({ S20631 }),
  .B2({ S20625 }),
  .ZN({ S20632 })
);
OAI21_X1 #() 
OAI21_X1_1777_ (
  .A({ S25957[1163] }),
  .B1({ S20132 }),
  .B2({ S20137 }),
  .ZN({ S20633 })
);
OAI211_X1 #() 
OAI211_X1_1170_ (
  .A({ S25957[1164] }),
  .B({ S20565 }),
  .C1({ S20212 }),
  .C2({ S20633 }),
  .ZN({ S20634 })
);
NAND2_X1 #() 
NAND2_X1_3393_ (
  .A1({ S20129 }),
  .A2({ S20160 }),
  .ZN({ S20635 })
);
NAND3_X1 #() 
NAND3_X1_3595_ (
  .A1({ S20129 }),
  .A2({ S20136 }),
  .A3({ S25957[1163] }),
  .ZN({ S20636 })
);
OAI211_X1 #() 
OAI211_X1_1171_ (
  .A({ S20131 }),
  .B({ S20636 }),
  .C1({ S20171 }),
  .C2({ S20635 }),
  .ZN({ S20637 })
);
NAND3_X1 #() 
NAND3_X1_3596_ (
  .A1({ S20634 }),
  .A2({ S14483 }),
  .A3({ S20637 }),
  .ZN({ S20638 })
);
NAND3_X1 #() 
NAND3_X1_3597_ (
  .A1({ S20132 }),
  .A2({ S20161 }),
  .A3({ S25957[1163] }),
  .ZN({ S20639 })
);
NOR2_X1 #() 
NOR2_X1_873_ (
  .A1({ S20258 }),
  .A2({ S20639 }),
  .ZN({ S20640 })
);
NAND3_X1 #() 
NAND3_X1_3598_ (
  .A1({ S20224 }),
  .A2({ S20227 }),
  .A3({ S20131 }),
  .ZN({ S20641 })
);
NAND3_X1 #() 
NAND3_X1_3599_ (
  .A1({ S20208 }),
  .A2({ S20325 }),
  .A3({ S25957[1164] }),
  .ZN({ S20642 })
);
OAI211_X1 #() 
OAI211_X1_1172_ (
  .A({ S25957[1165] }),
  .B({ S20642 }),
  .C1({ S20640 }),
  .C2({ S20641 }),
  .ZN({ S20643 })
);
NAND3_X1 #() 
NAND3_X1_3600_ (
  .A1({ S20638 }),
  .A2({ S25957[1166] }),
  .A3({ S20643 }),
  .ZN({ S20644 })
);
NAND2_X1 #() 
NAND2_X1_3394_ (
  .A1({ S20644 }),
  .A2({ S25957[1167] }),
  .ZN({ S20645 })
);
AOI21_X1 #() 
AOI21_X1_1848_ (
  .A({ S20131 }),
  .B1({ S20491 }),
  .B2({ S20411 }),
  .ZN({ S20646 })
);
OAI21_X1 #() 
OAI21_X1_1778_ (
  .A({ S25957[1165] }),
  .B1({ S20646 }),
  .B2({ S20197 }),
  .ZN({ S20647 })
);
NAND2_X1 #() 
NAND2_X1_3395_ (
  .A1({ S20178 }),
  .A2({ S20504 }),
  .ZN({ S20648 })
);
NAND3_X1 #() 
NAND3_X1_3601_ (
  .A1({ S20169 }),
  .A2({ S25957[1164] }),
  .A3({ S20417 }),
  .ZN({ S20649 })
);
NAND3_X1 #() 
NAND3_X1_3602_ (
  .A1({ S20648 }),
  .A2({ S20649 }),
  .A3({ S14483 }),
  .ZN({ S20650 })
);
NAND3_X1 #() 
NAND3_X1_3603_ (
  .A1({ S20647 }),
  .A2({ S20650 }),
  .A3({ S20130 }),
  .ZN({ S20651 })
);
NAND3_X1 #() 
NAND3_X1_3604_ (
  .A1({ S20559 }),
  .A2({ S20281 }),
  .A3({ S20131 }),
  .ZN({ S20652 })
);
OAI21_X1 #() 
OAI21_X1_1779_ (
  .A({ S25957[1164] }),
  .B1({ S20171 }),
  .B2({ S20358 }),
  .ZN({ S20653 })
);
OAI211_X1 #() 
OAI211_X1_1173_ (
  .A({ S20652 }),
  .B({ S14483 }),
  .C1({ S20653 }),
  .C2({ S20640 }),
  .ZN({ S20654 })
);
AND2_X1 #() 
AND2_X1_210_ (
  .A1({ S20510 }),
  .A2({ S25957[1163] }),
  .ZN({ S20655 })
);
OAI211_X1 #() 
OAI211_X1_1174_ (
  .A({ S20244 }),
  .B({ S65 }),
  .C1({ S20155 }),
  .C2({ S25957[1160] }),
  .ZN({ S20656 })
);
NAND2_X1 #() 
NAND2_X1_3396_ (
  .A1({ S20656 }),
  .A2({ S25957[1164] }),
  .ZN({ S20657 })
);
NAND2_X1 #() 
NAND2_X1_3397_ (
  .A1({ S20180 }),
  .A2({ S20244 }),
  .ZN({ S20658 })
);
AOI21_X1 #() 
AOI21_X1_1849_ (
  .A({ S14483 }),
  .B1({ S20658 }),
  .B2({ S20339 }),
  .ZN({ S20659 })
);
OAI21_X1 #() 
OAI21_X1_1780_ (
  .A({ S20659 }),
  .B1({ S20655 }),
  .B2({ S20657 }),
  .ZN({ S20660 })
);
NAND3_X1 #() 
NAND3_X1_3605_ (
  .A1({ S20654 }),
  .A2({ S20660 }),
  .A3({ S25957[1166] }),
  .ZN({ S20661 })
);
NAND3_X1 #() 
NAND3_X1_3606_ (
  .A1({ S20661 }),
  .A2({ S20192 }),
  .A3({ S20651 }),
  .ZN({ S20662 })
);
OAI211_X1 #() 
OAI211_X1_1175_ (
  .A({ S20662 }),
  .B({ S25957[1265] }),
  .C1({ S20632 }),
  .C2({ S20645 }),
  .ZN({ S20663 })
);
INV_X1 #() 
INV_X1_1144_ (
  .A({ S25957[1265] }),
  .ZN({ S20664 })
);
OAI21_X1 #() 
OAI21_X1_1781_ (
  .A({ S20662 }),
  .B1({ S20632 }),
  .B2({ S20645 }),
  .ZN({ S20665 })
);
NAND2_X1 #() 
NAND2_X1_3398_ (
  .A1({ S20665 }),
  .A2({ S20664 }),
  .ZN({ S20666 })
);
NAND3_X1 #() 
NAND3_X1_3607_ (
  .A1({ S20666 }),
  .A2({ S20621 }),
  .A3({ S20663 }),
  .ZN({ S20667 })
);
OAI211_X1 #() 
OAI211_X1_1176_ (
  .A({ S20662 }),
  .B({ S20664 }),
  .C1({ S20632 }),
  .C2({ S20645 }),
  .ZN({ S20668 })
);
NAND2_X1 #() 
NAND2_X1_3399_ (
  .A1({ S20665 }),
  .A2({ S25957[1265] }),
  .ZN({ S20669 })
);
NAND3_X1 #() 
NAND3_X1_3608_ (
  .A1({ S20669 }),
  .A2({ S25957[1233] }),
  .A3({ S20668 }),
  .ZN({ S20670 })
);
AOI21_X1 #() 
AOI21_X1_1850_ (
  .A({ S20620 }),
  .B1({ S20667 }),
  .B2({ S20670 }),
  .ZN({ S20671 })
);
NAND3_X1 #() 
NAND3_X1_3609_ (
  .A1({ S20666 }),
  .A2({ S25957[1233] }),
  .A3({ S20663 }),
  .ZN({ S20672 })
);
NAND3_X1 #() 
NAND3_X1_3610_ (
  .A1({ S20669 }),
  .A2({ S20621 }),
  .A3({ S20668 }),
  .ZN({ S20673 })
);
AOI21_X1 #() 
AOI21_X1_1851_ (
  .A({ S25957[1201] }),
  .B1({ S20672 }),
  .B2({ S20673 }),
  .ZN({ S20674 })
);
OAI21_X1 #() 
OAI21_X1_1782_ (
  .A({ S25957[1169] }),
  .B1({ S20671 }),
  .B2({ S20674 }),
  .ZN({ S20675 })
);
INV_X1 #() 
INV_X1_1145_ (
  .A({ S25957[1169] }),
  .ZN({ S20676 })
);
NAND3_X1 #() 
NAND3_X1_3611_ (
  .A1({ S20672 }),
  .A2({ S20673 }),
  .A3({ S25957[1201] }),
  .ZN({ S20677 })
);
NAND3_X1 #() 
NAND3_X1_3612_ (
  .A1({ S20667 }),
  .A2({ S20670 }),
  .A3({ S20620 }),
  .ZN({ S20678 })
);
NAND3_X1 #() 
NAND3_X1_3613_ (
  .A1({ S20677 }),
  .A2({ S20678 }),
  .A3({ S20676 }),
  .ZN({ S20679 })
);
NAND2_X1 #() 
NAND2_X1_3400_ (
  .A1({ S20675 }),
  .A2({ S20679 }),
  .ZN({ S25957[1041] })
);
NAND3_X1 #() 
NAND3_X1_3614_ (
  .A1({ S11498 }),
  .A2({ S11507 }),
  .A3({ S25956[18] }),
  .ZN({ S20680 })
);
NAND3_X1 #() 
NAND3_X1_3615_ (
  .A1({ S11432 }),
  .A2({ S11465 }),
  .A3({ S11487 }),
  .ZN({ S20681 })
);
NAND2_X1 #() 
NAND2_X1_3401_ (
  .A1({ S20680 }),
  .A2({ S20681 }),
  .ZN({ S20682 })
);
NAND2_X1 #() 
NAND2_X1_3402_ (
  .A1({ S11414 }),
  .A2({ S11404 }),
  .ZN({ S20683 })
);
INV_X1 #() 
INV_X1_1146_ (
  .A({ S20683 }),
  .ZN({ S25957[1266] })
);
OAI21_X1 #() 
OAI21_X1_1783_ (
  .A({ S65 }),
  .B1({ S20335 }),
  .B2({ S20266 }),
  .ZN({ S20684 })
);
NAND3_X1 #() 
NAND3_X1_3616_ (
  .A1({ S20684 }),
  .A2({ S25957[1164] }),
  .A3({ S20195 }),
  .ZN({ S20685 })
);
NAND3_X1 #() 
NAND3_X1_3617_ (
  .A1({ S20184 }),
  .A2({ S25957[1163] }),
  .A3({ S20252 }),
  .ZN({ S20686 })
);
NOR2_X1 #() 
NOR2_X1_874_ (
  .A1({ S20225 }),
  .A2({ S25957[1164] }),
  .ZN({ S20687 })
);
AOI21_X1 #() 
AOI21_X1_1852_ (
  .A({ S14483 }),
  .B1({ S20687 }),
  .B2({ S20686 }),
  .ZN({ S20688 })
);
OAI211_X1 #() 
OAI211_X1_1177_ (
  .A({ S20627 }),
  .B({ S20131 }),
  .C1({ S65 }),
  .C2({ S20416 }),
  .ZN({ S20689 })
);
NAND3_X1 #() 
NAND3_X1_3618_ (
  .A1({ S20196 }),
  .A2({ S25957[1163] }),
  .A3({ S20180 }),
  .ZN({ S20690 })
);
AOI21_X1 #() 
AOI21_X1_1853_ (
  .A({ S20131 }),
  .B1({ S20186 }),
  .B2({ S20137 }),
  .ZN({ S20691 })
);
AOI21_X1 #() 
AOI21_X1_1854_ (
  .A({ S25957[1165] }),
  .B1({ S20691 }),
  .B2({ S20690 }),
  .ZN({ S20692 })
);
AOI22_X1 #() 
AOI22_X1_394_ (
  .A1({ S20685 }),
  .A2({ S20688 }),
  .B1({ S20692 }),
  .B2({ S20689 }),
  .ZN({ S20693 })
);
NAND3_X1 #() 
NAND3_X1_3619_ (
  .A1({ S20244 }),
  .A2({ S25957[1163] }),
  .A3({ S25957[1161] }),
  .ZN({ S20694 })
);
NAND3_X1 #() 
NAND3_X1_3620_ (
  .A1({ S20694 }),
  .A2({ S25957[1164] }),
  .A3({ S20576 }),
  .ZN({ S20695 })
);
OAI221_X1 #() 
OAI221_X1_99_ (
  .A({ S20131 }),
  .B1({ S20150 }),
  .B2({ S65 }),
  .C1({ S20141 }),
  .C2({ S20132 }),
  .ZN({ S20696 })
);
NAND3_X1 #() 
NAND3_X1_3621_ (
  .A1({ S20696 }),
  .A2({ S14483 }),
  .A3({ S20695 }),
  .ZN({ S20697 })
);
NAND3_X1 #() 
NAND3_X1_3622_ (
  .A1({ S20161 }),
  .A2({ S25957[1163] }),
  .A3({ S25957[1160] }),
  .ZN({ S20698 })
);
NAND3_X1 #() 
NAND3_X1_3623_ (
  .A1({ S20504 }),
  .A2({ S25957[1164] }),
  .A3({ S20698 }),
  .ZN({ S20699 })
);
NAND3_X1 #() 
NAND3_X1_3624_ (
  .A1({ S20160 }),
  .A2({ S20150 }),
  .A3({ S65 }),
  .ZN({ S20700 })
);
NAND3_X1 #() 
NAND3_X1_3625_ (
  .A1({ S20217 }),
  .A2({ S25957[1163] }),
  .A3({ S20182 }),
  .ZN({ S20701 })
);
NAND3_X1 #() 
NAND3_X1_3626_ (
  .A1({ S20701 }),
  .A2({ S20131 }),
  .A3({ S20700 }),
  .ZN({ S20702 })
);
NAND3_X1 #() 
NAND3_X1_3627_ (
  .A1({ S20702 }),
  .A2({ S25957[1165] }),
  .A3({ S20699 }),
  .ZN({ S20703 })
);
NAND2_X1 #() 
NAND2_X1_3403_ (
  .A1({ S20703 }),
  .A2({ S20697 }),
  .ZN({ S20704 })
);
NAND2_X1 #() 
NAND2_X1_3404_ (
  .A1({ S20704 }),
  .A2({ S20130 }),
  .ZN({ S20705 })
);
OAI211_X1 #() 
OAI211_X1_1178_ (
  .A({ S20705 }),
  .B({ S25957[1167] }),
  .C1({ S20693 }),
  .C2({ S20130 }),
  .ZN({ S20706 })
);
AOI21_X1 #() 
AOI21_X1_1855_ (
  .A({ S65 }),
  .B1({ S20405 }),
  .B2({ S20193 }),
  .ZN({ S20707 })
);
OAI21_X1 #() 
OAI21_X1_1784_ (
  .A({ S25957[1164] }),
  .B1({ S20707 }),
  .B2({ S20564 }),
  .ZN({ S20708 })
);
OAI211_X1 #() 
OAI211_X1_1179_ (
  .A({ S20185 }),
  .B({ S20131 }),
  .C1({ S20144 }),
  .C2({ S20576 }),
  .ZN({ S20709 })
);
NAND3_X1 #() 
NAND3_X1_3628_ (
  .A1({ S20709 }),
  .A2({ S20708 }),
  .A3({ S25957[1165] }),
  .ZN({ S20710 })
);
NAND3_X1 #() 
NAND3_X1_3629_ (
  .A1({ S20161 }),
  .A2({ S20150 }),
  .A3({ S25957[1160] }),
  .ZN({ S20711 })
);
AOI22_X1 #() 
AOI22_X1_395_ (
  .A1({ S20711 }),
  .A2({ S65 }),
  .B1({ S20194 }),
  .B2({ S20260 }),
  .ZN({ S20712 })
);
OAI211_X1 #() 
OAI211_X1_1180_ (
  .A({ S20131 }),
  .B({ S20694 }),
  .C1({ S20406 }),
  .C2({ S25957[1163] }),
  .ZN({ S20713 })
);
OAI211_X1 #() 
OAI211_X1_1181_ (
  .A({ S20713 }),
  .B({ S14483 }),
  .C1({ S20131 }),
  .C2({ S20712 }),
  .ZN({ S20714 })
);
NAND3_X1 #() 
NAND3_X1_3630_ (
  .A1({ S20710 }),
  .A2({ S20714 }),
  .A3({ S25957[1166] }),
  .ZN({ S20715 })
);
NAND2_X1 #() 
NAND2_X1_3405_ (
  .A1({ S20194 }),
  .A2({ S20332 }),
  .ZN({ S20716 })
);
OAI211_X1 #() 
OAI211_X1_1182_ (
  .A({ S20716 }),
  .B({ S25957[1164] }),
  .C1({ S20218 }),
  .C2({ S20490 }),
  .ZN({ S20717 })
);
NAND3_X1 #() 
NAND3_X1_3631_ (
  .A1({ S20222 }),
  .A2({ S25957[1163] }),
  .A3({ S20348 }),
  .ZN({ S20718 })
);
NAND3_X1 #() 
NAND3_X1_3632_ (
  .A1({ S20718 }),
  .A2({ S20131 }),
  .A3({ S20265 }),
  .ZN({ S20719 })
);
NAND3_X1 #() 
NAND3_X1_3633_ (
  .A1({ S20717 }),
  .A2({ S20719 }),
  .A3({ S25957[1165] }),
  .ZN({ S20720 })
);
NAND2_X1 #() 
NAND2_X1_3406_ (
  .A1({ S20299 }),
  .A2({ S20555 }),
  .ZN({ S20721 })
);
AOI21_X1 #() 
AOI21_X1_1856_ (
  .A({ S20131 }),
  .B1({ S20285 }),
  .B2({ S25957[1163] }),
  .ZN({ S20722 })
);
AOI21_X1 #() 
AOI21_X1_1857_ (
  .A({ S25957[1165] }),
  .B1({ S20722 }),
  .B2({ S20395 }),
  .ZN({ S20723 })
);
NAND2_X1 #() 
NAND2_X1_3407_ (
  .A1({ S20723 }),
  .A2({ S20721 }),
  .ZN({ S20724 })
);
NAND2_X1 #() 
NAND2_X1_3408_ (
  .A1({ S20724 }),
  .A2({ S20720 }),
  .ZN({ S20725 })
);
NAND2_X1 #() 
NAND2_X1_3409_ (
  .A1({ S20725 }),
  .A2({ S20130 }),
  .ZN({ S20726 })
);
NAND3_X1 #() 
NAND3_X1_3634_ (
  .A1({ S20726 }),
  .A2({ S20715 }),
  .A3({ S20192 }),
  .ZN({ S20727 })
);
NAND3_X1 #() 
NAND3_X1_3635_ (
  .A1({ S20727 }),
  .A2({ S20706 }),
  .A3({ S25957[1266] }),
  .ZN({ S20728 })
);
NAND2_X1 #() 
NAND2_X1_3410_ (
  .A1({ S20685 }),
  .A2({ S20688 }),
  .ZN({ S20729 })
);
NAND2_X1 #() 
NAND2_X1_3411_ (
  .A1({ S20692 }),
  .A2({ S20689 }),
  .ZN({ S20730 })
);
NAND3_X1 #() 
NAND3_X1_3636_ (
  .A1({ S20730 }),
  .A2({ S20729 }),
  .A3({ S25957[1166] }),
  .ZN({ S20731 })
);
NAND3_X1 #() 
NAND3_X1_3637_ (
  .A1({ S20703 }),
  .A2({ S20130 }),
  .A3({ S20697 }),
  .ZN({ S20732 })
);
NAND3_X1 #() 
NAND3_X1_3638_ (
  .A1({ S20731 }),
  .A2({ S25957[1167] }),
  .A3({ S20732 }),
  .ZN({ S20733 })
);
NAND3_X1 #() 
NAND3_X1_3639_ (
  .A1({ S20331 }),
  .A2({ S20200 }),
  .A3({ S25957[1163] }),
  .ZN({ S20734 })
);
NAND3_X1 #() 
NAND3_X1_3640_ (
  .A1({ S20734 }),
  .A2({ S25957[1165] }),
  .A3({ S20515 }),
  .ZN({ S20735 })
);
OAI221_X1 #() 
OAI221_X1_100_ (
  .A({ S14483 }),
  .B1({ S20285 }),
  .B2({ S65 }),
  .C1({ S20351 }),
  .C2({ S20558 }),
  .ZN({ S20736 })
);
NAND3_X1 #() 
NAND3_X1_3641_ (
  .A1({ S20735 }),
  .A2({ S20736 }),
  .A3({ S20131 }),
  .ZN({ S20737 })
);
AOI21_X1 #() 
AOI21_X1_1858_ (
  .A({ S25957[1163] }),
  .B1({ S20635 }),
  .B2({ S20150 }),
  .ZN({ S20738 })
);
NAND2_X1 #() 
NAND2_X1_3412_ (
  .A1({ S20194 }),
  .A2({ S20260 }),
  .ZN({ S20739 })
);
NAND2_X1 #() 
NAND2_X1_3413_ (
  .A1({ S20739 }),
  .A2({ S14483 }),
  .ZN({ S20740 })
);
NAND2_X1 #() 
NAND2_X1_3414_ (
  .A1({ S20227 }),
  .A2({ S25957[1161] }),
  .ZN({ S20741 })
);
NAND4_X1 #() 
NAND4_X1_392_ (
  .A1({ S25957[1165] }),
  .A2({ S20741 }),
  .A3({ S20627 }),
  .A4({ S20136 }),
  .ZN({ S20742 })
);
OAI211_X1 #() 
OAI211_X1_1183_ (
  .A({ S20742 }),
  .B({ S25957[1164] }),
  .C1({ S20740 }),
  .C2({ S20738 }),
  .ZN({ S20743 })
);
AOI21_X1 #() 
AOI21_X1_1859_ (
  .A({ S20130 }),
  .B1({ S20737 }),
  .B2({ S20743 }),
  .ZN({ S20744 })
);
AOI21_X1 #() 
AOI21_X1_1860_ (
  .A({ S25957[1166] }),
  .B1({ S20724 }),
  .B2({ S20720 }),
  .ZN({ S20745 })
);
OAI21_X1 #() 
OAI21_X1_1785_ (
  .A({ S20192 }),
  .B1({ S20744 }),
  .B2({ S20745 }),
  .ZN({ S20746 })
);
NAND3_X1 #() 
NAND3_X1_3642_ (
  .A1({ S20746 }),
  .A2({ S20733 }),
  .A3({ S20683 }),
  .ZN({ S20747 })
);
AOI21_X1 #() 
AOI21_X1_1861_ (
  .A({ S25956[50] }),
  .B1({ S20728 }),
  .B2({ S20747 }),
  .ZN({ S20748 })
);
NAND3_X1 #() 
NAND3_X1_3643_ (
  .A1({ S20746 }),
  .A2({ S20733 }),
  .A3({ S25957[1266] }),
  .ZN({ S20749 })
);
NAND3_X1 #() 
NAND3_X1_3644_ (
  .A1({ S20727 }),
  .A2({ S20706 }),
  .A3({ S20683 }),
  .ZN({ S20750 })
);
AOI21_X1 #() 
AOI21_X1_1862_ (
  .A({ S10969 }),
  .B1({ S20750 }),
  .B2({ S20749 }),
  .ZN({ S20751 })
);
OAI21_X1 #() 
OAI21_X1_1786_ (
  .A({ S20682 }),
  .B1({ S20748 }),
  .B2({ S20751 }),
  .ZN({ S20752 })
);
NAND3_X1 #() 
NAND3_X1_3645_ (
  .A1({ S20750 }),
  .A2({ S20749 }),
  .A3({ S10969 }),
  .ZN({ S20753 })
);
NAND3_X1 #() 
NAND3_X1_3646_ (
  .A1({ S20728 }),
  .A2({ S20747 }),
  .A3({ S25956[50] }),
  .ZN({ S20754 })
);
NAND3_X1 #() 
NAND3_X1_3647_ (
  .A1({ S20753 }),
  .A2({ S20754 }),
  .A3({ S25957[1170] }),
  .ZN({ S20755 })
);
NAND2_X1 #() 
NAND2_X1_3415_ (
  .A1({ S20752 }),
  .A2({ S20755 }),
  .ZN({ S25957[1042] })
);
NAND2_X1 #() 
NAND2_X1_3416_ (
  .A1({ S12855 }),
  .A2({ S12844 }),
  .ZN({ S25957[1199] })
);
OAI21_X1 #() 
OAI21_X1_1787_ (
  .A({ S11550 }),
  .B1({ S19428 }),
  .B2({ S19429 }),
  .ZN({ S20756 })
);
NAND3_X1 #() 
NAND3_X1_3648_ (
  .A1({ S19431 }),
  .A2({ S25956[0] }),
  .A3({ S19427 }),
  .ZN({ S20757 })
);
NAND3_X1 #() 
NAND3_X1_3649_ (
  .A1({ S25957[1153] }),
  .A2({ S20756 }),
  .A3({ S20757 }),
  .ZN({ S20758 })
);
INV_X1 #() 
INV_X1_1147_ (
  .A({ S20758 }),
  .ZN({ S75 })
);
OAI21_X1 #() 
OAI21_X1_1788_ (
  .A({ S11539 }),
  .B1({ S19478 }),
  .B2({ S19482 }),
  .ZN({ S20759 })
);
NAND3_X1 #() 
NAND3_X1_3650_ (
  .A1({ S19484 }),
  .A2({ S19485 }),
  .A3({ S25956[1] }),
  .ZN({ S20760 })
);
NAND2_X1 #() 
NAND2_X1_3417_ (
  .A1({ S20759 }),
  .A2({ S20760 }),
  .ZN({ S20761 })
);
NAND3_X1 #() 
NAND3_X1_3651_ (
  .A1({ S20761 }),
  .A2({ S19430 }),
  .A3({ S19432 }),
  .ZN({ S76 })
);
INV_X1 #() 
INV_X1_1148_ (
  .A({ S12802 }),
  .ZN({ S25957[1231] })
);
NAND4_X1 #() 
NAND4_X1_393_ (
  .A1({ S19536 }),
  .A2({ S19539 }),
  .A3({ S19483 }),
  .A4({ S19486 }),
  .ZN({ S20762 })
);
NAND4_X1 #() 
NAND4_X1_394_ (
  .A1({ S20756 }),
  .A2({ S20757 }),
  .A3({ S19536 }),
  .A4({ S19539 }),
  .ZN({ S20763 })
);
NAND2_X1 #() 
NAND2_X1_3418_ (
  .A1({ S76 }),
  .A2({ S20763 }),
  .ZN({ S20764 })
);
NAND2_X1 #() 
NAND2_X1_3419_ (
  .A1({ S20764 }),
  .A2({ S20762 }),
  .ZN({ S20765 })
);
NAND4_X1 #() 
NAND4_X1_395_ (
  .A1({ S19430 }),
  .A2({ S19432 }),
  .A3({ S19536 }),
  .A4({ S19539 }),
  .ZN({ S20766 })
);
INV_X1 #() 
INV_X1_1149_ (
  .A({ S20766 }),
  .ZN({ S20767 })
);
NAND3_X1 #() 
NAND3_X1_3652_ (
  .A1({ S19537 }),
  .A2({ S19538 }),
  .A3({ S25956[2] }),
  .ZN({ S20768 })
);
NAND3_X1 #() 
NAND3_X1_3653_ (
  .A1({ S19535 }),
  .A2({ S11642 }),
  .A3({ S19533 }),
  .ZN({ S20769 })
);
NAND4_X1 #() 
NAND4_X1_396_ (
  .A1({ S20768 }),
  .A2({ S20769 }),
  .A3({ S20759 }),
  .A4({ S20760 }),
  .ZN({ S20770 })
);
OAI21_X1 #() 
OAI21_X1_1789_ (
  .A({ S68 }),
  .B1({ S20770 }),
  .B2({ S25957[1152] }),
  .ZN({ S20771 })
);
OAI21_X1 #() 
OAI21_X1_1790_ (
  .A({ S25957[1156] }),
  .B1({ S20771 }),
  .B2({ S20767 }),
  .ZN({ S20772 })
);
AOI21_X1 #() 
AOI21_X1_1863_ (
  .A({ S20772 }),
  .B1({ S20765 }),
  .B2({ S25957[1155] }),
  .ZN({ S20773 })
);
INV_X1 #() 
INV_X1_1150_ (
  .A({ S25957[1156] }),
  .ZN({ S20774 })
);
NAND2_X1 #() 
NAND2_X1_3420_ (
  .A1({ S20768 }),
  .A2({ S20769 }),
  .ZN({ S20775 })
);
NAND3_X1 #() 
NAND3_X1_3654_ (
  .A1({ S20761 }),
  .A2({ S20756 }),
  .A3({ S20757 }),
  .ZN({ S20776 })
);
NAND2_X1 #() 
NAND2_X1_3421_ (
  .A1({ S20776 }),
  .A2({ S20775 }),
  .ZN({ S20777 })
);
NAND2_X1 #() 
NAND2_X1_3422_ (
  .A1({ S25957[1154] }),
  .A2({ S20761 }),
  .ZN({ S20778 })
);
NAND3_X1 #() 
NAND3_X1_3655_ (
  .A1({ S20777 }),
  .A2({ S25957[1155] }),
  .A3({ S20778 }),
  .ZN({ S20779 })
);
NAND4_X1 #() 
NAND4_X1_397_ (
  .A1({ S19430 }),
  .A2({ S19432 }),
  .A3({ S20768 }),
  .A4({ S20769 }),
  .ZN({ S20780 })
);
NAND3_X1 #() 
NAND3_X1_3656_ (
  .A1({ S20778 }),
  .A2({ S20780 }),
  .A3({ S68 }),
  .ZN({ S20781 })
);
AND3_X1 #() 
AND3_X1_133_ (
  .A1({ S20779 }),
  .A2({ S20774 }),
  .A3({ S20781 }),
  .ZN({ S20782 })
);
OAI21_X1 #() 
OAI21_X1_1791_ (
  .A({ S25957[1157] }),
  .B1({ S20773 }),
  .B2({ S20782 }),
  .ZN({ S20783 })
);
NAND2_X1 #() 
NAND2_X1_3423_ (
  .A1({ S19248 }),
  .A2({ S19247 }),
  .ZN({ S20784 })
);
NAND4_X1 #() 
NAND4_X1_398_ (
  .A1({ S19536 }),
  .A2({ S19539 }),
  .A3({ S20759 }),
  .A4({ S20760 }),
  .ZN({ S20785 })
);
INV_X1 #() 
INV_X1_1151_ (
  .A({ S20785 }),
  .ZN({ S20786 })
);
NAND4_X1 #() 
NAND4_X1_399_ (
  .A1({ S20756 }),
  .A2({ S20757 }),
  .A3({ S20768 }),
  .A4({ S20769 }),
  .ZN({ S20787 })
);
NAND2_X1 #() 
NAND2_X1_3424_ (
  .A1({ S20787 }),
  .A2({ S25957[1155] }),
  .ZN({ S20788 })
);
NAND4_X1 #() 
NAND4_X1_400_ (
  .A1({ S20778 }),
  .A2({ S20766 }),
  .A3({ S20780 }),
  .A4({ S20785 }),
  .ZN({ S20789 })
);
AOI21_X1 #() 
AOI21_X1_1864_ (
  .A({ S25957[1156] }),
  .B1({ S20789 }),
  .B2({ S68 }),
  .ZN({ S20790 })
);
OAI21_X1 #() 
OAI21_X1_1792_ (
  .A({ S20790 }),
  .B1({ S20786 }),
  .B2({ S20788 }),
  .ZN({ S20791 })
);
NAND2_X1 #() 
NAND2_X1_3425_ (
  .A1({ S20758 }),
  .A2({ S25957[1154] }),
  .ZN({ S20792 })
);
NAND3_X1 #() 
NAND3_X1_3657_ (
  .A1({ S25957[1153] }),
  .A2({ S19430 }),
  .A3({ S19432 }),
  .ZN({ S20793 })
);
NAND3_X1 #() 
NAND3_X1_3658_ (
  .A1({ S20776 }),
  .A2({ S20793 }),
  .A3({ S20775 }),
  .ZN({ S20794 })
);
AOI21_X1 #() 
AOI21_X1_1865_ (
  .A({ S68 }),
  .B1({ S20794 }),
  .B2({ S20792 }),
  .ZN({ S20795 })
);
NAND3_X1 #() 
NAND3_X1_3659_ (
  .A1({ S20758 }),
  .A2({ S76 }),
  .A3({ S25957[1154] }),
  .ZN({ S20796 })
);
NAND3_X1 #() 
NAND3_X1_3660_ (
  .A1({ S20796 }),
  .A2({ S68 }),
  .A3({ S20763 }),
  .ZN({ S20797 })
);
NAND2_X1 #() 
NAND2_X1_3426_ (
  .A1({ S20797 }),
  .A2({ S25957[1156] }),
  .ZN({ S20798 })
);
OAI211_X1 #() 
OAI211_X1_1184_ (
  .A({ S20791 }),
  .B({ S20784 }),
  .C1({ S20795 }),
  .C2({ S20798 }),
  .ZN({ S20799 })
);
AND3_X1 #() 
AND3_X1_134_ (
  .A1({ S20799 }),
  .A2({ S20783 }),
  .A3({ S19126 }),
  .ZN({ S20800 })
);
OAI21_X1 #() 
OAI21_X1_1793_ (
  .A({ S25957[1156] }),
  .B1({ S20777 }),
  .B2({ S68 }),
  .ZN({ S20801 })
);
NAND2_X1 #() 
NAND2_X1_3427_ (
  .A1({ S20766 }),
  .A2({ S25957[1153] }),
  .ZN({ S20802 })
);
AOI22_X1 #() 
AOI22_X1_396_ (
  .A1({ S19430 }),
  .A2({ S19432 }),
  .B1({ S19539 }),
  .B2({ S19536 }),
  .ZN({ S20803 })
);
NAND2_X1 #() 
NAND2_X1_3428_ (
  .A1({ S20803 }),
  .A2({ S25957[1155] }),
  .ZN({ S20804 })
);
OAI21_X1 #() 
OAI21_X1_1794_ (
  .A({ S20804 }),
  .B1({ S20802 }),
  .B2({ S25957[1155] }),
  .ZN({ S20805 })
);
AOI21_X1 #() 
AOI21_X1_1866_ (
  .A({ S20775 }),
  .B1({ S20776 }),
  .B2({ S20793 }),
  .ZN({ S20806 })
);
INV_X1 #() 
INV_X1_1152_ (
  .A({ S20762 }),
  .ZN({ S20807 })
);
NAND2_X1 #() 
NAND2_X1_3429_ (
  .A1({ S20807 }),
  .A2({ S25957[1152] }),
  .ZN({ S20808 })
);
INV_X1 #() 
INV_X1_1153_ (
  .A({ S20808 }),
  .ZN({ S20809 })
);
OAI21_X1 #() 
OAI21_X1_1795_ (
  .A({ S25957[1155] }),
  .B1({ S20806 }),
  .B2({ S20809 }),
  .ZN({ S20810 })
);
OAI21_X1 #() 
OAI21_X1_1796_ (
  .A({ S20810 }),
  .B1({ S25957[1155] }),
  .B2({ S20765 }),
  .ZN({ S20811 })
);
OAI22_X1 #() 
OAI22_X1_96_ (
  .A1({ S20811 }),
  .A2({ S25957[1156] }),
  .B1({ S20801 }),
  .B2({ S20805 }),
  .ZN({ S20812 })
);
NAND2_X1 #() 
NAND2_X1_3430_ (
  .A1({ S20793 }),
  .A2({ S68 }),
  .ZN({ S20813 })
);
NAND2_X1 #() 
NAND2_X1_3431_ (
  .A1({ S20793 }),
  .A2({ S20762 }),
  .ZN({ S20814 })
);
NAND2_X1 #() 
NAND2_X1_3432_ (
  .A1({ S20814 }),
  .A2({ S25957[1155] }),
  .ZN({ S20815 })
);
AOI21_X1 #() 
AOI21_X1_1867_ (
  .A({ S20774 }),
  .B1({ S20815 }),
  .B2({ S20813 }),
  .ZN({ S20816 })
);
NOR2_X1 #() 
NOR2_X1_875_ (
  .A1({ S68 }),
  .A2({ S25957[1153] }),
  .ZN({ S20817 })
);
NAND2_X1 #() 
NAND2_X1_3433_ (
  .A1({ S76 }),
  .A2({ S25957[1154] }),
  .ZN({ S20818 })
);
NAND2_X1 #() 
NAND2_X1_3434_ (
  .A1({ S20756 }),
  .A2({ S20757 }),
  .ZN({ S20819 })
);
NAND3_X1 #() 
NAND3_X1_3661_ (
  .A1({ S20819 }),
  .A2({ S20761 }),
  .A3({ S20775 }),
  .ZN({ S20820 })
);
NAND2_X1 #() 
NAND2_X1_3435_ (
  .A1({ S20818 }),
  .A2({ S20820 }),
  .ZN({ S20821 })
);
AOI21_X1 #() 
AOI21_X1_1868_ (
  .A({ S20821 }),
  .B1({ S20817 }),
  .B2({ S25957[1152] }),
  .ZN({ S20822 })
);
AOI211_X1 #() 
AOI211_X1_52_ (
  .A({ S25957[1157] }),
  .B({ S20816 }),
  .C1({ S20774 }),
  .C2({ S20822 }),
  .ZN({ S20823 })
);
AOI21_X1 #() 
AOI21_X1_1869_ (
  .A({ S20823 }),
  .B1({ S20812 }),
  .B2({ S25957[1157] }),
  .ZN({ S20824 })
);
NOR2_X1 #() 
NOR2_X1_876_ (
  .A1({ S20824 }),
  .A2({ S19126 }),
  .ZN({ S20825 })
);
OAI21_X1 #() 
OAI21_X1_1797_ (
  .A({ S25957[1158] }),
  .B1({ S20825 }),
  .B2({ S20800 }),
  .ZN({ S20826 })
);
NAND2_X1 #() 
NAND2_X1_3436_ (
  .A1({ S25957[1155] }),
  .A2({ S20785 }),
  .ZN({ S20827 })
);
INV_X1 #() 
INV_X1_1154_ (
  .A({ S20827 }),
  .ZN({ S20828 })
);
INV_X1 #() 
INV_X1_1155_ (
  .A({ S20770 }),
  .ZN({ S20829 })
);
NOR2_X1 #() 
NOR2_X1_877_ (
  .A1({ S20829 }),
  .A2({ S25957[1155] }),
  .ZN({ S20830 })
);
NAND2_X1 #() 
NAND2_X1_3437_ (
  .A1({ S20758 }),
  .A2({ S20775 }),
  .ZN({ S20831 })
);
AOI22_X1 #() 
AOI22_X1_397_ (
  .A1({ S20776 }),
  .A2({ S20828 }),
  .B1({ S20830 }),
  .B2({ S20831 }),
  .ZN({ S20832 })
);
NOR2_X1 #() 
NOR2_X1_878_ (
  .A1({ S20803 }),
  .A2({ S68 }),
  .ZN({ S20833 })
);
NAND2_X1 #() 
NAND2_X1_3438_ (
  .A1({ S20833 }),
  .A2({ S20762 }),
  .ZN({ S20834 })
);
OAI211_X1 #() 
OAI211_X1_1185_ (
  .A({ S20834 }),
  .B({ S25957[1156] }),
  .C1({ S25957[1155] }),
  .C2({ S20819 }),
  .ZN({ S20835 })
);
OAI211_X1 #() 
OAI211_X1_1186_ (
  .A({ S20835 }),
  .B({ S25957[1157] }),
  .C1({ S25957[1156] }),
  .C2({ S20832 }),
  .ZN({ S20836 })
);
AOI21_X1 #() 
AOI21_X1_1870_ (
  .A({ S68 }),
  .B1({ S20829 }),
  .B2({ S20819 }),
  .ZN({ S20837 })
);
OAI21_X1 #() 
OAI21_X1_1798_ (
  .A({ S68 }),
  .B1({ S20785 }),
  .B2({ S20819 }),
  .ZN({ S20838 })
);
OAI21_X1 #() 
OAI21_X1_1799_ (
  .A({ S25957[1156] }),
  .B1({ S20806 }),
  .B2({ S20838 }),
  .ZN({ S20839 })
);
NAND2_X1 #() 
NAND2_X1_3439_ (
  .A1({ S20776 }),
  .A2({ S25957[1154] }),
  .ZN({ S20840 })
);
NOR2_X1 #() 
NOR2_X1_879_ (
  .A1({ S20840 }),
  .A2({ S20813 }),
  .ZN({ S20841 })
);
NOR2_X1 #() 
NOR2_X1_880_ (
  .A1({ S68 }),
  .A2({ S20775 }),
  .ZN({ S20842 })
);
NAND2_X1 #() 
NAND2_X1_3440_ (
  .A1({ S20842 }),
  .A2({ S20758 }),
  .ZN({ S20843 })
);
NAND2_X1 #() 
NAND2_X1_3441_ (
  .A1({ S20843 }),
  .A2({ S20774 }),
  .ZN({ S20844 })
);
OAI221_X1 #() 
OAI221_X1_101_ (
  .A({ S20784 }),
  .B1({ S20841 }),
  .B2({ S20844 }),
  .C1({ S20839 }),
  .C2({ S20837 }),
  .ZN({ S20845 })
);
AOI21_X1 #() 
AOI21_X1_1871_ (
  .A({ S25957[1159] }),
  .B1({ S20836 }),
  .B2({ S20845 }),
  .ZN({ S20846 })
);
NAND2_X1 #() 
NAND2_X1_3442_ (
  .A1({ S20780 }),
  .A2({ S68 }),
  .ZN({ S20847 })
);
INV_X1 #() 
INV_X1_1156_ (
  .A({ S20847 }),
  .ZN({ S20848 })
);
NAND3_X1 #() 
NAND3_X1_3662_ (
  .A1({ S20762 }),
  .A2({ S20770 }),
  .A3({ S25957[1152] }),
  .ZN({ S20849 })
);
NAND2_X1 #() 
NAND2_X1_3443_ (
  .A1({ S20849 }),
  .A2({ S76 }),
  .ZN({ S20850 })
);
NAND2_X1 #() 
NAND2_X1_3444_ (
  .A1({ S20850 }),
  .A2({ S20848 }),
  .ZN({ S20851 })
);
NAND2_X1 #() 
NAND2_X1_3445_ (
  .A1({ S20817 }),
  .A2({ S20775 }),
  .ZN({ S20852 })
);
NAND3_X1 #() 
NAND3_X1_3663_ (
  .A1({ S20851 }),
  .A2({ S20774 }),
  .A3({ S20852 }),
  .ZN({ S20853 })
);
AOI21_X1 #() 
AOI21_X1_1872_ (
  .A({ S68 }),
  .B1({ S20794 }),
  .B2({ S20796 }),
  .ZN({ S20854 })
);
NAND2_X1 #() 
NAND2_X1_3446_ (
  .A1({ S20763 }),
  .A2({ S68 }),
  .ZN({ S20855 })
);
NOR2_X1 #() 
NOR2_X1_881_ (
  .A1({ S20855 }),
  .A2({ S20829 }),
  .ZN({ S20856 })
);
OAI21_X1 #() 
OAI21_X1_1800_ (
  .A({ S25957[1156] }),
  .B1({ S20854 }),
  .B2({ S20856 }),
  .ZN({ S20857 })
);
AOI21_X1 #() 
AOI21_X1_1873_ (
  .A({ S25957[1157] }),
  .B1({ S20857 }),
  .B2({ S20853 }),
  .ZN({ S20858 })
);
NOR2_X1 #() 
NOR2_X1_882_ (
  .A1({ S25957[1155] }),
  .A2({ S20761 }),
  .ZN({ S20859 })
);
INV_X1 #() 
INV_X1_1157_ (
  .A({ S20817 }),
  .ZN({ S20860 })
);
NAND2_X1 #() 
NAND2_X1_3447_ (
  .A1({ S20804 }),
  .A2({ S20860 }),
  .ZN({ S20861 })
);
AOI211_X1 #() 
AOI211_X1_53_ (
  .A({ S20774 }),
  .B({ S20861 }),
  .C1({ S20787 }),
  .C2({ S20859 }),
  .ZN({ S20862 })
);
AOI21_X1 #() 
AOI21_X1_1874_ (
  .A({ S25957[1156] }),
  .B1({ S20766 }),
  .B2({ S68 }),
  .ZN({ S20863 })
);
NOR2_X1 #() 
NOR2_X1_883_ (
  .A1({ S20859 }),
  .A2({ S75 }),
  .ZN({ S20864 })
);
AOI211_X1 #() 
AOI211_X1_54_ (
  .A({ S20784 }),
  .B({ S20862 }),
  .C1({ S20863 }),
  .C2({ S20864 }),
  .ZN({ S20865 })
);
NOR3_X1 #() 
NOR3_X1_121_ (
  .A1({ S20865 }),
  .A2({ S20858 }),
  .A3({ S19126 }),
  .ZN({ S20866 })
);
OAI21_X1 #() 
OAI21_X1_1801_ (
  .A({ S19194 }),
  .B1({ S20866 }),
  .B2({ S20846 }),
  .ZN({ S20867 })
);
NAND2_X1 #() 
NAND2_X1_3448_ (
  .A1({ S20867 }),
  .A2({ S20826 }),
  .ZN({ S20868 })
);
NAND2_X1 #() 
NAND2_X1_3449_ (
  .A1({ S20868 }),
  .A2({ S12761 }),
  .ZN({ S20869 })
);
NAND3_X1 #() 
NAND3_X1_3664_ (
  .A1({ S20867 }),
  .A2({ S20826 }),
  .A3({ S25957[1263] }),
  .ZN({ S20870 })
);
NAND3_X1 #() 
NAND3_X1_3665_ (
  .A1({ S20869 }),
  .A2({ S20870 }),
  .A3({ S25957[1231] }),
  .ZN({ S20871 })
);
NAND2_X1 #() 
NAND2_X1_3450_ (
  .A1({ S20869 }),
  .A2({ S20870 }),
  .ZN({ S25957[1135] })
);
NAND2_X1 #() 
NAND2_X1_3451_ (
  .A1({ S25957[1135] }),
  .A2({ S12802 }),
  .ZN({ S20872 })
);
NAND2_X1 #() 
NAND2_X1_3452_ (
  .A1({ S20872 }),
  .A2({ S20871 }),
  .ZN({ S25957[1103] })
);
INV_X1 #() 
INV_X1_1158_ (
  .A({ S25957[1103] }),
  .ZN({ S20873 })
);
NAND2_X1 #() 
NAND2_X1_3453_ (
  .A1({ S20873 }),
  .A2({ S5686 }),
  .ZN({ S20874 })
);
NAND2_X1 #() 
NAND2_X1_3454_ (
  .A1({ S25957[1103] }),
  .A2({ S25956[15] }),
  .ZN({ S20875 })
);
AND2_X1 #() 
AND2_X1_211_ (
  .A1({ S20874 }),
  .A2({ S20875 }),
  .ZN({ S25957[1039] })
);
NOR2_X1 #() 
NOR2_X1_884_ (
  .A1({ S13673 }),
  .A2({ S13684 }),
  .ZN({ S25957[1198] })
);
INV_X1 #() 
INV_X1_1159_ (
  .A({ S25957[1230] }),
  .ZN({ S20876 })
);
AOI21_X1 #() 
AOI21_X1_1875_ (
  .A({ S20859 }),
  .B1({ S20814 }),
  .B2({ S25957[1155] }),
  .ZN({ S20877 })
);
NAND3_X1 #() 
NAND3_X1_3666_ (
  .A1({ S20817 }),
  .A2({ S20780 }),
  .A3({ S20763 }),
  .ZN({ S20878 })
);
OAI211_X1 #() 
OAI211_X1_1187_ (
  .A({ S20878 }),
  .B({ S25957[1156] }),
  .C1({ S25957[1155] }),
  .C2({ S20818 }),
  .ZN({ S20879 })
);
OAI211_X1 #() 
OAI211_X1_1188_ (
  .A({ S20879 }),
  .B({ S25957[1157] }),
  .C1({ S25957[1156] }),
  .C2({ S20877 }),
  .ZN({ S20880 })
);
NAND3_X1 #() 
NAND3_X1_3667_ (
  .A1({ S20780 }),
  .A2({ S20763 }),
  .A3({ S20770 }),
  .ZN({ S20881 })
);
NAND2_X1 #() 
NAND2_X1_3455_ (
  .A1({ S20881 }),
  .A2({ S25957[1155] }),
  .ZN({ S20882 })
);
INV_X1 #() 
INV_X1_1160_ (
  .A({ S20882 }),
  .ZN({ S20883 })
);
AOI21_X1 #() 
AOI21_X1_1876_ (
  .A({ S20883 }),
  .B1({ S20848 }),
  .B2({ S20794 }),
  .ZN({ S20884 })
);
NAND3_X1 #() 
NAND3_X1_3668_ (
  .A1({ S20819 }),
  .A2({ S20761 }),
  .A3({ S25957[1154] }),
  .ZN({ S20885 })
);
AND2_X1 #() 
AND2_X1_212_ (
  .A1({ S20885 }),
  .A2({ S25957[1155] }),
  .ZN({ S20886 })
);
AOI21_X1 #() 
AOI21_X1_1877_ (
  .A({ S20886 }),
  .B1({ S20789 }),
  .B2({ S68 }),
  .ZN({ S20887 })
);
OAI21_X1 #() 
OAI21_X1_1802_ (
  .A({ S20774 }),
  .B1({ S20831 }),
  .B2({ S68 }),
  .ZN({ S20888 })
);
OAI221_X1 #() 
OAI221_X1_102_ (
  .A({ S20784 }),
  .B1({ S20887 }),
  .B2({ S20888 }),
  .C1({ S20884 }),
  .C2({ S20774 }),
  .ZN({ S20889 })
);
NAND3_X1 #() 
NAND3_X1_3669_ (
  .A1({ S20889 }),
  .A2({ S25957[1158] }),
  .A3({ S20880 }),
  .ZN({ S20890 })
);
NAND3_X1 #() 
NAND3_X1_3670_ (
  .A1({ S20819 }),
  .A2({ S25957[1153] }),
  .A3({ S20775 }),
  .ZN({ S20891 })
);
NAND2_X1 #() 
NAND2_X1_3456_ (
  .A1({ S20891 }),
  .A2({ S20778 }),
  .ZN({ S20892 })
);
NOR2_X1 #() 
NOR2_X1_885_ (
  .A1({ S20892 }),
  .A2({ S68 }),
  .ZN({ S20893 })
);
INV_X1 #() 
INV_X1_1161_ (
  .A({ S76 }),
  .ZN({ S20894 })
);
NAND3_X1 #() 
NAND3_X1_3671_ (
  .A1({ S25957[1152] }),
  .A2({ S25957[1153] }),
  .A3({ S25957[1154] }),
  .ZN({ S20895 })
);
INV_X1 #() 
INV_X1_1162_ (
  .A({ S20895 }),
  .ZN({ S20896 })
);
OAI21_X1 #() 
OAI21_X1_1803_ (
  .A({ S68 }),
  .B1({ S20896 }),
  .B2({ S20894 }),
  .ZN({ S20897 })
);
NAND2_X1 #() 
NAND2_X1_3457_ (
  .A1({ S20897 }),
  .A2({ S20774 }),
  .ZN({ S20898 })
);
NAND2_X1 #() 
NAND2_X1_3458_ (
  .A1({ S20829 }),
  .A2({ S25957[1155] }),
  .ZN({ S20899 })
);
NAND2_X1 #() 
NAND2_X1_3459_ (
  .A1({ S20859 }),
  .A2({ S20767 }),
  .ZN({ S20900 })
);
NAND2_X1 #() 
NAND2_X1_3460_ (
  .A1({ S20900 }),
  .A2({ S20899 }),
  .ZN({ S20901 })
);
OAI21_X1 #() 
OAI21_X1_1804_ (
  .A({ S25957[1156] }),
  .B1({ S20901 }),
  .B2({ S20841 }),
  .ZN({ S20902 })
);
OAI211_X1 #() 
OAI211_X1_1189_ (
  .A({ S20902 }),
  .B({ S25957[1157] }),
  .C1({ S20893 }),
  .C2({ S20898 }),
  .ZN({ S20903 })
);
NAND3_X1 #() 
NAND3_X1_3672_ (
  .A1({ S76 }),
  .A2({ S20787 }),
  .A3({ S25957[1155] }),
  .ZN({ S20904 })
);
INV_X1 #() 
INV_X1_1163_ (
  .A({ S20904 }),
  .ZN({ S20905 })
);
AOI22_X1 #() 
AOI22_X1_398_ (
  .A1({ S20905 }),
  .A2({ S20766 }),
  .B1({ S20848 }),
  .B2({ S20794 }),
  .ZN({ S20906 })
);
OAI21_X1 #() 
OAI21_X1_1805_ (
  .A({ S25957[1156] }),
  .B1({ S20777 }),
  .B2({ S25957[1155] }),
  .ZN({ S20907 })
);
OAI221_X1 #() 
OAI221_X1_103_ (
  .A({ S20784 }),
  .B1({ S20907 }),
  .B2({ S20861 }),
  .C1({ S20906 }),
  .C2({ S25957[1156] }),
  .ZN({ S20908 })
);
AND2_X1 #() 
AND2_X1_213_ (
  .A1({ S20903 }),
  .A2({ S20908 }),
  .ZN({ S20909 })
);
NAND2_X1 #() 
NAND2_X1_3461_ (
  .A1({ S20909 }),
  .A2({ S19194 }),
  .ZN({ S20910 })
);
AOI21_X1 #() 
AOI21_X1_1878_ (
  .A({ S19126 }),
  .B1({ S20890 }),
  .B2({ S20910 }),
  .ZN({ S20911 })
);
NAND4_X1 #() 
NAND4_X1_401_ (
  .A1({ S20763 }),
  .A2({ S20778 }),
  .A3({ S20780 }),
  .A4({ S68 }),
  .ZN({ S20912 })
);
OAI211_X1 #() 
OAI211_X1_1190_ (
  .A({ S20912 }),
  .B({ S25957[1156] }),
  .C1({ S68 }),
  .C2({ S20764 }),
  .ZN({ S20913 })
);
NAND2_X1 #() 
NAND2_X1_3462_ (
  .A1({ S20793 }),
  .A2({ S20770 }),
  .ZN({ S20914 })
);
INV_X1 #() 
INV_X1_1164_ (
  .A({ S20914 }),
  .ZN({ S20915 })
);
AOI21_X1 #() 
AOI21_X1_1879_ (
  .A({ S25957[1156] }),
  .B1({ S20915 }),
  .B2({ S20804 }),
  .ZN({ S20916 })
);
INV_X1 #() 
INV_X1_1165_ (
  .A({ S20916 }),
  .ZN({ S20917 })
);
AOI21_X1 #() 
AOI21_X1_1880_ (
  .A({ S20784 }),
  .B1({ S20917 }),
  .B2({ S20913 }),
  .ZN({ S20918 })
);
NAND2_X1 #() 
NAND2_X1_3463_ (
  .A1({ S20762 }),
  .A2({ S20819 }),
  .ZN({ S20919 })
);
NAND2_X1 #() 
NAND2_X1_3464_ (
  .A1({ S20919 }),
  .A2({ S68 }),
  .ZN({ S20920 })
);
AOI21_X1 #() 
AOI21_X1_1881_ (
  .A({ S20774 }),
  .B1({ S20920 }),
  .B2({ S20827 }),
  .ZN({ S20921 })
);
AOI21_X1 #() 
AOI21_X1_1882_ (
  .A({ S25957[1156] }),
  .B1({ S20796 }),
  .B2({ S68 }),
  .ZN({ S20922 })
);
AOI211_X1 #() 
AOI211_X1_55_ (
  .A({ S25957[1157] }),
  .B({ S20921 }),
  .C1({ S20882 }),
  .C2({ S20922 }),
  .ZN({ S20923 })
);
OAI21_X1 #() 
OAI21_X1_1806_ (
  .A({ S25957[1158] }),
  .B1({ S20923 }),
  .B2({ S20918 }),
  .ZN({ S20924 })
);
OAI211_X1 #() 
OAI211_X1_1191_ (
  .A({ S20779 }),
  .B({ S25957[1156] }),
  .C1({ S20809 }),
  .C2({ S25957[1155] }),
  .ZN({ S20925 })
);
OAI211_X1 #() 
OAI211_X1_1192_ (
  .A({ S20763 }),
  .B({ S20762 }),
  .C1({ S20770 }),
  .C2({ S25957[1152] }),
  .ZN({ S20926 })
);
NAND3_X1 #() 
NAND3_X1_3673_ (
  .A1({ S20926 }),
  .A2({ S20774 }),
  .A3({ S25957[1155] }),
  .ZN({ S20927 })
);
NAND3_X1 #() 
NAND3_X1_3674_ (
  .A1({ S20925 }),
  .A2({ S20784 }),
  .A3({ S20927 }),
  .ZN({ S20928 })
);
NAND2_X1 #() 
NAND2_X1_3465_ (
  .A1({ S20885 }),
  .A2({ S25957[1155] }),
  .ZN({ S20929 })
);
OAI211_X1 #() 
OAI211_X1_1193_ (
  .A({ S25957[1156] }),
  .B({ S20855 }),
  .C1({ S20929 }),
  .C2({ S75 }),
  .ZN({ S20930 })
);
INV_X1 #() 
INV_X1_1166_ (
  .A({ S20830 }),
  .ZN({ S20931 })
);
NAND2_X1 #() 
NAND2_X1_3466_ (
  .A1({ S20778 }),
  .A2({ S25957[1155] }),
  .ZN({ S20932 })
);
OAI221_X1 #() 
OAI221_X1_104_ (
  .A({ S20774 }),
  .B1({ S20932 }),
  .B2({ S20786 }),
  .C1({ S20809 }),
  .C2({ S20931 }),
  .ZN({ S20933 })
);
AND2_X1 #() 
AND2_X1_214_ (
  .A1({ S20933 }),
  .A2({ S20930 }),
  .ZN({ S20934 })
);
OAI211_X1 #() 
OAI211_X1_1194_ (
  .A({ S19194 }),
  .B({ S20928 }),
  .C1({ S20934 }),
  .C2({ S20784 }),
  .ZN({ S20935 })
);
AOI21_X1 #() 
AOI21_X1_1883_ (
  .A({ S25957[1159] }),
  .B1({ S20935 }),
  .B2({ S20924 }),
  .ZN({ S20936 })
);
OAI21_X1 #() 
OAI21_X1_1807_ (
  .A({ S25957[1262] }),
  .B1({ S20911 }),
  .B2({ S20936 }),
  .ZN({ S20937 })
);
OR3_X1 #() 
OR3_X1_20_ (
  .A1({ S20911 }),
  .A2({ S20936 }),
  .A3({ S25957[1262] }),
  .ZN({ S20938 })
);
NAND2_X1 #() 
NAND2_X1_3467_ (
  .A1({ S20938 }),
  .A2({ S20937 }),
  .ZN({ S25957[1134] })
);
NAND2_X1 #() 
NAND2_X1_3468_ (
  .A1({ S25957[1134] }),
  .A2({ S20876 }),
  .ZN({ S20939 })
);
NAND3_X1 #() 
NAND3_X1_3675_ (
  .A1({ S20938 }),
  .A2({ S25957[1230] }),
  .A3({ S20937 }),
  .ZN({ S20940 })
);
NAND2_X1 #() 
NAND2_X1_3469_ (
  .A1({ S20939 }),
  .A2({ S20940 }),
  .ZN({ S25957[1102] })
);
NAND2_X1 #() 
NAND2_X1_3470_ (
  .A1({ S25957[1102] }),
  .A2({ S25956[14] }),
  .ZN({ S20941 })
);
NAND3_X1 #() 
NAND3_X1_3676_ (
  .A1({ S20939 }),
  .A2({ S20940 }),
  .A3({ S6132 }),
  .ZN({ S20942 })
);
AND2_X1 #() 
AND2_X1_215_ (
  .A1({ S20941 }),
  .A2({ S20942 }),
  .ZN({ S25957[1038] })
);
NAND2_X1 #() 
NAND2_X1_3471_ (
  .A1({ S14453 }),
  .A2({ S14461 }),
  .ZN({ S25957[1197] })
);
NOR2_X1 #() 
NOR2_X1_886_ (
  .A1({ S14352 }),
  .A2({ S14330 }),
  .ZN({ S25957[1261] })
);
INV_X1 #() 
INV_X1_1167_ (
  .A({ S25957[1261] }),
  .ZN({ S20943 })
);
AOI22_X1 #() 
AOI22_X1_399_ (
  .A1({ S20780 }),
  .A2({ S20770 }),
  .B1({ S20819 }),
  .B2({ S25957[1153] }),
  .ZN({ S20944 })
);
NAND4_X1 #() 
NAND4_X1_402_ (
  .A1({ S20778 }),
  .A2({ S20766 }),
  .A3({ S20785 }),
  .A4({ S68 }),
  .ZN({ S20945 })
);
NAND2_X1 #() 
NAND2_X1_3472_ (
  .A1({ S20891 }),
  .A2({ S25957[1155] }),
  .ZN({ S20946 })
);
OAI211_X1 #() 
OAI211_X1_1195_ (
  .A({ S25957[1156] }),
  .B({ S20945 }),
  .C1({ S20946 }),
  .C2({ S20944 }),
  .ZN({ S20947 })
);
NOR2_X1 #() 
NOR2_X1_887_ (
  .A1({ S25957[1152] }),
  .A2({ S68 }),
  .ZN({ S20948 })
);
INV_X1 #() 
INV_X1_1168_ (
  .A({ S20948 }),
  .ZN({ S20949 })
);
NAND3_X1 #() 
NAND3_X1_3677_ (
  .A1({ S20793 }),
  .A2({ S20763 }),
  .A3({ S68 }),
  .ZN({ S20950 })
);
AND2_X1 #() 
AND2_X1_216_ (
  .A1({ S20949 }),
  .A2({ S20950 }),
  .ZN({ S20951 })
);
OAI211_X1 #() 
OAI211_X1_1196_ (
  .A({ S20947 }),
  .B({ S25957[1157] }),
  .C1({ S25957[1156] }),
  .C2({ S20951 }),
  .ZN({ S20952 })
);
NAND4_X1 #() 
NAND4_X1_403_ (
  .A1({ S20763 }),
  .A2({ S20778 }),
  .A3({ S20780 }),
  .A4({ S25957[1155] }),
  .ZN({ S20953 })
);
NAND3_X1 #() 
NAND3_X1_3678_ (
  .A1({ S20891 }),
  .A2({ S68 }),
  .A3({ S20787 }),
  .ZN({ S20954 })
);
AOI21_X1 #() 
AOI21_X1_1884_ (
  .A({ S25957[1156] }),
  .B1({ S20954 }),
  .B2({ S20953 }),
  .ZN({ S20955 })
);
NAND2_X1 #() 
NAND2_X1_3473_ (
  .A1({ S20786 }),
  .A2({ S25957[1152] }),
  .ZN({ S20956 })
);
AOI21_X1 #() 
AOI21_X1_1885_ (
  .A({ S25957[1155] }),
  .B1({ S20956 }),
  .B2({ S20792 }),
  .ZN({ S20957 })
);
OAI21_X1 #() 
OAI21_X1_1808_ (
  .A({ S20784 }),
  .B1({ S20957 }),
  .B2({ S20801 }),
  .ZN({ S20958 })
);
OAI211_X1 #() 
OAI211_X1_1197_ (
  .A({ S20952 }),
  .B({ S25957[1158] }),
  .C1({ S20955 }),
  .C2({ S20958 }),
  .ZN({ S20959 })
);
NAND2_X1 #() 
NAND2_X1_3474_ (
  .A1({ S20804 }),
  .A2({ S20847 }),
  .ZN({ S20960 })
);
NAND2_X1 #() 
NAND2_X1_3475_ (
  .A1({ S20916 }),
  .A2({ S20960 }),
  .ZN({ S20961 })
);
NOR2_X1 #() 
NOR2_X1_888_ (
  .A1({ S20831 }),
  .A2({ S68 }),
  .ZN({ S20962 })
);
NAND2_X1 #() 
NAND2_X1_3476_ (
  .A1({ S20891 }),
  .A2({ S68 }),
  .ZN({ S20963 })
);
INV_X1 #() 
INV_X1_1169_ (
  .A({ S20963 }),
  .ZN({ S20964 })
);
OAI21_X1 #() 
OAI21_X1_1809_ (
  .A({ S25957[1156] }),
  .B1({ S20964 }),
  .B2({ S20962 }),
  .ZN({ S20965 })
);
NAND3_X1 #() 
NAND3_X1_3679_ (
  .A1({ S20961 }),
  .A2({ S20965 }),
  .A3({ S25957[1157] }),
  .ZN({ S20966 })
);
NAND3_X1 #() 
NAND3_X1_3680_ (
  .A1({ S20776 }),
  .A2({ S20793 }),
  .A3({ S25957[1154] }),
  .ZN({ S20967 })
);
NAND3_X1 #() 
NAND3_X1_3681_ (
  .A1({ S20967 }),
  .A2({ S20808 }),
  .A3({ S25957[1155] }),
  .ZN({ S20968 })
);
NAND4_X1 #() 
NAND4_X1_404_ (
  .A1({ S20793 }),
  .A2({ S20776 }),
  .A3({ S20766 }),
  .A4({ S68 }),
  .ZN({ S20969 })
);
NAND3_X1 #() 
NAND3_X1_3682_ (
  .A1({ S20968 }),
  .A2({ S25957[1156] }),
  .A3({ S20969 }),
  .ZN({ S20970 })
);
AOI22_X1 #() 
AOI22_X1_400_ (
  .A1({ S20896 }),
  .A2({ S68 }),
  .B1({ S25957[1152] }),
  .B2({ S20817 }),
  .ZN({ S20971 })
);
OAI211_X1 #() 
OAI211_X1_1198_ (
  .A({ S20970 }),
  .B({ S20784 }),
  .C1({ S25957[1156] }),
  .C2({ S20971 }),
  .ZN({ S20972 })
);
NAND3_X1 #() 
NAND3_X1_3683_ (
  .A1({ S20972 }),
  .A2({ S19194 }),
  .A3({ S20966 }),
  .ZN({ S20973 })
);
NAND3_X1 #() 
NAND3_X1_3684_ (
  .A1({ S20973 }),
  .A2({ S20959 }),
  .A3({ S19126 }),
  .ZN({ S20974 })
);
NAND2_X1 #() 
NAND2_X1_3477_ (
  .A1({ S20787 }),
  .A2({ S20761 }),
  .ZN({ S20975 })
);
NAND2_X1 #() 
NAND2_X1_3478_ (
  .A1({ S20975 }),
  .A2({ S68 }),
  .ZN({ S20976 })
);
NAND3_X1 #() 
NAND3_X1_3685_ (
  .A1({ S20758 }),
  .A2({ S25957[1155] }),
  .A3({ S20770 }),
  .ZN({ S20977 })
);
AND3_X1 #() 
AND3_X1_135_ (
  .A1({ S20976 }),
  .A2({ S20804 }),
  .A3({ S20977 }),
  .ZN({ S20978 })
);
NAND3_X1 #() 
NAND3_X1_3686_ (
  .A1({ S20793 }),
  .A2({ S20766 }),
  .A3({ S20785 }),
  .ZN({ S20979 })
);
OAI221_X1 #() 
OAI221_X1_105_ (
  .A({ S25957[1156] }),
  .B1({ S20949 }),
  .B2({ S20807 }),
  .C1({ S20979 }),
  .C2({ S25957[1155] }),
  .ZN({ S20980 })
);
OAI21_X1 #() 
OAI21_X1_1810_ (
  .A({ S20980 }),
  .B1({ S25957[1156] }),
  .B2({ S20978 }),
  .ZN({ S20981 })
);
OAI21_X1 #() 
OAI21_X1_1811_ (
  .A({ S20774 }),
  .B1({ S20883 }),
  .B2({ S20944 }),
  .ZN({ S20982 })
);
NAND2_X1 #() 
NAND2_X1_3479_ (
  .A1({ S20778 }),
  .A2({ S20787 }),
  .ZN({ S20983 })
);
NAND2_X1 #() 
NAND2_X1_3480_ (
  .A1({ S20983 }),
  .A2({ S68 }),
  .ZN({ S20984 })
);
NAND3_X1 #() 
NAND3_X1_3687_ (
  .A1({ S20763 }),
  .A2({ S25957[1155] }),
  .A3({ S20762 }),
  .ZN({ S20985 })
);
AND2_X1 #() 
AND2_X1_217_ (
  .A1({ S20984 }),
  .A2({ S20985 }),
  .ZN({ S20986 })
);
OAI211_X1 #() 
OAI211_X1_1199_ (
  .A({ S20982 }),
  .B({ S20784 }),
  .C1({ S20774 }),
  .C2({ S20986 }),
  .ZN({ S20987 })
);
OAI21_X1 #() 
OAI21_X1_1812_ (
  .A({ S20987 }),
  .B1({ S20981 }),
  .B2({ S20784 }),
  .ZN({ S20988 })
);
NAND2_X1 #() 
NAND2_X1_3481_ (
  .A1({ S20796 }),
  .A2({ S20820 }),
  .ZN({ S20989 })
);
NAND2_X1 #() 
NAND2_X1_3482_ (
  .A1({ S20989 }),
  .A2({ S25957[1155] }),
  .ZN({ S20990 })
);
AOI21_X1 #() 
AOI21_X1_1886_ (
  .A({ S25957[1156] }),
  .B1({ S20990 }),
  .B2({ S20838 }),
  .ZN({ S20991 })
);
AOI21_X1 #() 
AOI21_X1_1887_ (
  .A({ S25957[1154] }),
  .B1({ S20776 }),
  .B2({ S20793 }),
  .ZN({ S20992 })
);
NAND2_X1 #() 
NAND2_X1_3483_ (
  .A1({ S20992 }),
  .A2({ S25957[1155] }),
  .ZN({ S20993 })
);
AOI21_X1 #() 
AOI21_X1_1888_ (
  .A({ S25957[1153] }),
  .B1({ S25957[1152] }),
  .B2({ S20775 }),
  .ZN({ S20994 })
);
AOI21_X1 #() 
AOI21_X1_1889_ (
  .A({ S20774 }),
  .B1({ S20994 }),
  .B2({ S68 }),
  .ZN({ S20995 })
);
NAND2_X1 #() 
NAND2_X1_3484_ (
  .A1({ S20993 }),
  .A2({ S20995 }),
  .ZN({ S20996 })
);
NAND2_X1 #() 
NAND2_X1_3485_ (
  .A1({ S20996 }),
  .A2({ S20784 }),
  .ZN({ S20997 })
);
NAND2_X1 #() 
NAND2_X1_3486_ (
  .A1({ S20758 }),
  .A2({ S20778 }),
  .ZN({ S20998 })
);
AOI21_X1 #() 
AOI21_X1_1890_ (
  .A({ S20817 }),
  .B1({ S20998 }),
  .B2({ S68 }),
  .ZN({ S20999 })
);
INV_X1 #() 
INV_X1_1170_ (
  .A({ S20842 }),
  .ZN({ S21000 })
);
NAND3_X1 #() 
NAND3_X1_3688_ (
  .A1({ S21000 }),
  .A2({ S20780 }),
  .A3({ S20776 }),
  .ZN({ S21001 })
);
NAND3_X1 #() 
NAND3_X1_3689_ (
  .A1({ S21001 }),
  .A2({ S25957[1156] }),
  .A3({ S20843 }),
  .ZN({ S21002 })
);
OAI211_X1 #() 
OAI211_X1_1200_ (
  .A({ S21002 }),
  .B({ S25957[1157] }),
  .C1({ S25957[1156] }),
  .C2({ S20999 }),
  .ZN({ S21003 })
);
OAI211_X1 #() 
OAI211_X1_1201_ (
  .A({ S21003 }),
  .B({ S19194 }),
  .C1({ S20991 }),
  .C2({ S20997 }),
  .ZN({ S21004 })
);
OAI211_X1 #() 
OAI211_X1_1202_ (
  .A({ S21004 }),
  .B({ S25957[1159] }),
  .C1({ S20988 }),
  .C2({ S19194 }),
  .ZN({ S21005 })
);
NAND2_X1 #() 
NAND2_X1_3487_ (
  .A1({ S21005 }),
  .A2({ S20974 }),
  .ZN({ S21006 })
);
NAND2_X1 #() 
NAND2_X1_3488_ (
  .A1({ S21006 }),
  .A2({ S20943 }),
  .ZN({ S21007 })
);
NAND3_X1 #() 
NAND3_X1_3690_ (
  .A1({ S21005 }),
  .A2({ S25957[1261] }),
  .A3({ S20974 }),
  .ZN({ S21008 })
);
NAND3_X1 #() 
NAND3_X1_3691_ (
  .A1({ S21007 }),
  .A2({ S25956[45] }),
  .A3({ S21008 }),
  .ZN({ S21009 })
);
NAND2_X1 #() 
NAND2_X1_3489_ (
  .A1({ S21007 }),
  .A2({ S21008 }),
  .ZN({ S25957[1133] })
);
NAND2_X1 #() 
NAND2_X1_3490_ (
  .A1({ S25957[1133] }),
  .A2({ S13744 }),
  .ZN({ S21010 })
);
NAND3_X1 #() 
NAND3_X1_3692_ (
  .A1({ S21010 }),
  .A2({ S14483 }),
  .A3({ S21009 }),
  .ZN({ S21011 })
);
NAND2_X1 #() 
NAND2_X1_3491_ (
  .A1({ S25957[1133] }),
  .A2({ S25956[45] }),
  .ZN({ S21012 })
);
NAND3_X1 #() 
NAND3_X1_3693_ (
  .A1({ S21007 }),
  .A2({ S13744 }),
  .A3({ S21008 }),
  .ZN({ S21013 })
);
NAND3_X1 #() 
NAND3_X1_3694_ (
  .A1({ S21012 }),
  .A2({ S21013 }),
  .A3({ S25957[1165] }),
  .ZN({ S21014 })
);
NAND2_X1 #() 
NAND2_X1_3492_ (
  .A1({ S21011 }),
  .A2({ S21014 }),
  .ZN({ S21015 })
);
INV_X1 #() 
INV_X1_1171_ (
  .A({ S21015 }),
  .ZN({ S25957[1037] })
);
NOR2_X1 #() 
NOR2_X1_889_ (
  .A1({ S15198 }),
  .A2({ S15239 }),
  .ZN({ S25957[1196] })
);
NAND2_X1 #() 
NAND2_X1_3493_ (
  .A1({ S15219 }),
  .A2({ S15228 }),
  .ZN({ S25957[1228] })
);
NAND2_X1 #() 
NAND2_X1_3494_ (
  .A1({ S15143 }),
  .A2({ S15049 }),
  .ZN({ S25957[1260] })
);
NAND2_X1 #() 
NAND2_X1_3495_ (
  .A1({ S20885 }),
  .A2({ S68 }),
  .ZN({ S21016 })
);
INV_X1 #() 
INV_X1_1172_ (
  .A({ S21016 }),
  .ZN({ S21017 })
);
NOR2_X1 #() 
NOR2_X1_890_ (
  .A1({ S20801 }),
  .A2({ S21017 }),
  .ZN({ S21018 })
);
NAND3_X1 #() 
NAND3_X1_3695_ (
  .A1({ S20785 }),
  .A2({ S20819 }),
  .A3({ S68 }),
  .ZN({ S21019 })
);
AND3_X1 #() 
AND3_X1_136_ (
  .A1({ S20834 }),
  .A2({ S20774 }),
  .A3({ S21019 }),
  .ZN({ S21020 })
);
OAI21_X1 #() 
OAI21_X1_1813_ (
  .A({ S25957[1157] }),
  .B1({ S21020 }),
  .B2({ S21018 }),
  .ZN({ S21021 })
);
NAND2_X1 #() 
NAND2_X1_3496_ (
  .A1({ S20817 }),
  .A2({ S20763 }),
  .ZN({ S21022 })
);
NAND2_X1 #() 
NAND2_X1_3497_ (
  .A1({ S20998 }),
  .A2({ S68 }),
  .ZN({ S21023 })
);
NAND3_X1 #() 
NAND3_X1_3696_ (
  .A1({ S21023 }),
  .A2({ S25957[1156] }),
  .A3({ S21022 }),
  .ZN({ S21024 })
);
NAND2_X1 #() 
NAND2_X1_3498_ (
  .A1({ S20828 }),
  .A2({ S20776 }),
  .ZN({ S21025 })
);
NAND3_X1 #() 
NAND3_X1_3697_ (
  .A1({ S20780 }),
  .A2({ S68 }),
  .A3({ S20762 }),
  .ZN({ S21026 })
);
NAND3_X1 #() 
NAND3_X1_3698_ (
  .A1({ S21025 }),
  .A2({ S21026 }),
  .A3({ S20774 }),
  .ZN({ S21027 })
);
AND2_X1 #() 
AND2_X1_218_ (
  .A1({ S21027 }),
  .A2({ S21024 }),
  .ZN({ S21028 })
);
OAI21_X1 #() 
OAI21_X1_1814_ (
  .A({ S21021 }),
  .B1({ S21028 }),
  .B2({ S25957[1157] }),
  .ZN({ S21029 })
);
NAND2_X1 #() 
NAND2_X1_3499_ (
  .A1({ S21029 }),
  .A2({ S25957[1158] }),
  .ZN({ S21030 })
);
NAND3_X1 #() 
NAND3_X1_3699_ (
  .A1({ S20819 }),
  .A2({ S25957[1153] }),
  .A3({ S25957[1154] }),
  .ZN({ S21031 })
);
INV_X1 #() 
INV_X1_1173_ (
  .A({ S20838 }),
  .ZN({ S21032 })
);
NAND2_X1 #() 
NAND2_X1_3500_ (
  .A1({ S21032 }),
  .A2({ S21031 }),
  .ZN({ S21033 })
);
OAI21_X1 #() 
OAI21_X1_1815_ (
  .A({ S21033 }),
  .B1({ S20786 }),
  .B2({ S20815 }),
  .ZN({ S21034 })
);
NOR2_X1 #() 
NOR2_X1_891_ (
  .A1({ S21034 }),
  .A2({ S20774 }),
  .ZN({ S21035 })
);
NAND2_X1 #() 
NAND2_X1_3501_ (
  .A1({ S20794 }),
  .A2({ S20840 }),
  .ZN({ S21036 })
);
NAND2_X1 #() 
NAND2_X1_3502_ (
  .A1({ S25957[1156] }),
  .A2({ S25957[1155] }),
  .ZN({ S21037 })
);
NAND3_X1 #() 
NAND3_X1_3700_ (
  .A1({ S20802 }),
  .A2({ S20975 }),
  .A3({ S25957[1156] }),
  .ZN({ S21038 })
);
AOI22_X1 #() 
AOI22_X1_401_ (
  .A1({ S25957[1155] }),
  .A2({ S21036 }),
  .B1({ S21038 }),
  .B2({ S21037 }),
  .ZN({ S21039 })
);
NAND2_X1 #() 
NAND2_X1_3503_ (
  .A1({ S20817 }),
  .A2({ S20787 }),
  .ZN({ S21040 })
);
OAI21_X1 #() 
OAI21_X1_1816_ (
  .A({ S21040 }),
  .B1({ S20963 }),
  .B2({ S20983 }),
  .ZN({ S21041 })
);
OAI21_X1 #() 
OAI21_X1_1817_ (
  .A({ S20784 }),
  .B1({ S21041 }),
  .B2({ S25957[1156] }),
  .ZN({ S21042 })
);
AOI21_X1 #() 
AOI21_X1_1891_ (
  .A({ S25957[1155] }),
  .B1({ S20794 }),
  .B2({ S20792 }),
  .ZN({ S21043 })
);
NAND2_X1 #() 
NAND2_X1_3504_ (
  .A1({ S20979 }),
  .A2({ S25957[1155] }),
  .ZN({ S21044 })
);
NAND2_X1 #() 
NAND2_X1_3505_ (
  .A1({ S21044 }),
  .A2({ S20774 }),
  .ZN({ S21045 })
);
OAI21_X1 #() 
OAI21_X1_1818_ (
  .A({ S25957[1157] }),
  .B1({ S21045 }),
  .B2({ S21043 }),
  .ZN({ S21046 })
);
OAI221_X1 #() 
OAI221_X1_106_ (
  .A({ S19194 }),
  .B1({ S21046 }),
  .B2({ S21039 }),
  .C1({ S21035 }),
  .C2({ S21042 }),
  .ZN({ S21047 })
);
NAND3_X1 #() 
NAND3_X1_3701_ (
  .A1({ S21030 }),
  .A2({ S21047 }),
  .A3({ S25957[1159] }),
  .ZN({ S21048 })
);
NAND2_X1 #() 
NAND2_X1_3506_ (
  .A1({ S20762 }),
  .A2({ S68 }),
  .ZN({ S21049 })
);
INV_X1 #() 
INV_X1_1174_ (
  .A({ S21049 }),
  .ZN({ S21050 })
);
AOI211_X1 #() 
AOI211_X1_56_ (
  .A({ S20774 }),
  .B({ S20861 }),
  .C1({ S20818 }),
  .C2({ S21050 }),
  .ZN({ S21051 })
);
AOI21_X1 #() 
AOI21_X1_1892_ (
  .A({ S20774 }),
  .B1({ S121 }),
  .B2({ S20775 }),
  .ZN({ S21052 })
);
NOR2_X1 #() 
NOR2_X1_892_ (
  .A1({ S20785 }),
  .A2({ S20819 }),
  .ZN({ S21053 })
);
OAI211_X1 #() 
OAI211_X1_1203_ (
  .A({ S21000 }),
  .B({ S20774 }),
  .C1({ S20847 }),
  .C2({ S21053 }),
  .ZN({ S21054 })
);
NAND2_X1 #() 
NAND2_X1_3507_ (
  .A1({ S21054 }),
  .A2({ S20784 }),
  .ZN({ S21055 })
);
NAND2_X1 #() 
NAND2_X1_3508_ (
  .A1({ S20793 }),
  .A2({ S25957[1154] }),
  .ZN({ S21056 })
);
NAND3_X1 #() 
NAND3_X1_3702_ (
  .A1({ S20758 }),
  .A2({ S76 }),
  .A3({ S20775 }),
  .ZN({ S21057 })
);
AOI21_X1 #() 
AOI21_X1_1893_ (
  .A({ S25957[1155] }),
  .B1({ S21057 }),
  .B2({ S21056 }),
  .ZN({ S21058 })
);
NAND2_X1 #() 
NAND2_X1_3509_ (
  .A1({ S20953 }),
  .A2({ S20774 }),
  .ZN({ S21059 })
);
OAI21_X1 #() 
OAI21_X1_1819_ (
  .A({ S25957[1157] }),
  .B1({ S21058 }),
  .B2({ S21059 }),
  .ZN({ S21060 })
);
OAI22_X1 #() 
OAI22_X1_97_ (
  .A1({ S21051 }),
  .A2({ S21055 }),
  .B1({ S21052 }),
  .B2({ S21060 }),
  .ZN({ S21061 })
);
AND2_X1 #() 
AND2_X1_219_ (
  .A1({ S20779 }),
  .A2({ S20984 }),
  .ZN({ S21062 })
);
OAI211_X1 #() 
OAI211_X1_1204_ (
  .A({ S20993 }),
  .B({ S20774 }),
  .C1({ S25957[1155] }),
  .C2({ S20758 }),
  .ZN({ S21063 })
);
OAI211_X1 #() 
OAI211_X1_1205_ (
  .A({ S25957[1157] }),
  .B({ S21063 }),
  .C1({ S21062 }),
  .C2({ S20774 }),
  .ZN({ S21064 })
);
NAND2_X1 #() 
NAND2_X1_3510_ (
  .A1({ S20821 }),
  .A2({ S68 }),
  .ZN({ S21065 })
);
AOI21_X1 #() 
AOI21_X1_1894_ (
  .A({ S25957[1156] }),
  .B1({ S21065 }),
  .B2({ S20904 }),
  .ZN({ S21066 })
);
NAND2_X1 #() 
NAND2_X1_3511_ (
  .A1({ S20833 }),
  .A2({ S20777 }),
  .ZN({ S21067 })
);
AND3_X1 #() 
AND3_X1_137_ (
  .A1({ S21067 }),
  .A2({ S21023 }),
  .A3({ S25957[1156] }),
  .ZN({ S21068 })
);
OAI21_X1 #() 
OAI21_X1_1820_ (
  .A({ S20784 }),
  .B1({ S21066 }),
  .B2({ S21068 }),
  .ZN({ S21069 })
);
NAND3_X1 #() 
NAND3_X1_3703_ (
  .A1({ S21064 }),
  .A2({ S21069 }),
  .A3({ S19194 }),
  .ZN({ S21070 })
);
OAI211_X1 #() 
OAI211_X1_1206_ (
  .A({ S21070 }),
  .B({ S19126 }),
  .C1({ S19194 }),
  .C2({ S21061 }),
  .ZN({ S21071 })
);
NAND3_X1 #() 
NAND3_X1_3704_ (
  .A1({ S21048 }),
  .A2({ S21071 }),
  .A3({ S25957[1260] }),
  .ZN({ S21072 })
);
INV_X1 #() 
INV_X1_1175_ (
  .A({ S25957[1260] }),
  .ZN({ S21073 })
);
AND2_X1 #() 
AND2_X1_220_ (
  .A1({ S21064 }),
  .A2({ S21069 }),
  .ZN({ S21074 })
);
NAND2_X1 #() 
NAND2_X1_3512_ (
  .A1({ S21061 }),
  .A2({ S25957[1158] }),
  .ZN({ S21075 })
);
OAI211_X1 #() 
OAI211_X1_1207_ (
  .A({ S19126 }),
  .B({ S21075 }),
  .C1({ S21074 }),
  .C2({ S25957[1158] }),
  .ZN({ S21076 })
);
OAI211_X1 #() 
OAI211_X1_1208_ (
  .A({ S21021 }),
  .B({ S25957[1158] }),
  .C1({ S21028 }),
  .C2({ S25957[1157] }),
  .ZN({ S21077 })
);
NAND2_X1 #() 
NAND2_X1_3513_ (
  .A1({ S21034 }),
  .A2({ S25957[1156] }),
  .ZN({ S21078 })
);
NAND2_X1 #() 
NAND2_X1_3514_ (
  .A1({ S21041 }),
  .A2({ S20774 }),
  .ZN({ S21079 })
);
AOI21_X1 #() 
AOI21_X1_1895_ (
  .A({ S25957[1157] }),
  .B1({ S21078 }),
  .B2({ S21079 }),
  .ZN({ S21080 })
);
NOR2_X1 #() 
NOR2_X1_893_ (
  .A1({ S21046 }),
  .A2({ S21039 }),
  .ZN({ S21081 })
);
OAI21_X1 #() 
OAI21_X1_1821_ (
  .A({ S19194 }),
  .B1({ S21080 }),
  .B2({ S21081 }),
  .ZN({ S21082 })
);
NAND3_X1 #() 
NAND3_X1_3705_ (
  .A1({ S21082 }),
  .A2({ S25957[1159] }),
  .A3({ S21077 }),
  .ZN({ S21083 })
);
NAND3_X1 #() 
NAND3_X1_3706_ (
  .A1({ S21083 }),
  .A2({ S21076 }),
  .A3({ S21073 }),
  .ZN({ S21084 })
);
NAND3_X1 #() 
NAND3_X1_3707_ (
  .A1({ S21084 }),
  .A2({ S25957[1228] }),
  .A3({ S21072 }),
  .ZN({ S21085 })
);
INV_X1 #() 
INV_X1_1176_ (
  .A({ S25957[1228] }),
  .ZN({ S21086 })
);
NAND3_X1 #() 
NAND3_X1_3708_ (
  .A1({ S21048 }),
  .A2({ S21071 }),
  .A3({ S21073 }),
  .ZN({ S21087 })
);
NAND3_X1 #() 
NAND3_X1_3709_ (
  .A1({ S21083 }),
  .A2({ S21076 }),
  .A3({ S25957[1260] }),
  .ZN({ S21088 })
);
NAND3_X1 #() 
NAND3_X1_3710_ (
  .A1({ S21088 }),
  .A2({ S21086 }),
  .A3({ S21087 }),
  .ZN({ S21089 })
);
NAND3_X1 #() 
NAND3_X1_3711_ (
  .A1({ S21085 }),
  .A2({ S21089 }),
  .A3({ S25956[12] }),
  .ZN({ S21090 })
);
NAND3_X1 #() 
NAND3_X1_3712_ (
  .A1({ S21084 }),
  .A2({ S21086 }),
  .A3({ S21072 }),
  .ZN({ S21091 })
);
NAND3_X1 #() 
NAND3_X1_3713_ (
  .A1({ S21088 }),
  .A2({ S25957[1228] }),
  .A3({ S21087 }),
  .ZN({ S21092 })
);
NAND3_X1 #() 
NAND3_X1_3714_ (
  .A1({ S21091 }),
  .A2({ S21092 }),
  .A3({ S5708 }),
  .ZN({ S21093 })
);
AND2_X1 #() 
AND2_X1_221_ (
  .A1({ S21093 }),
  .A2({ S21090 }),
  .ZN({ S25957[1036] })
);
NOR2_X1 #() 
NOR2_X1_894_ (
  .A1({ S16000 }),
  .A2({ S16042 }),
  .ZN({ S25957[1195] })
);
INV_X1 #() 
INV_X1_1177_ (
  .A({ S25957[1195] }),
  .ZN({ S21094 })
);
NAND2_X1 #() 
NAND2_X1_3515_ (
  .A1({ S16020 }),
  .A2({ S16031 }),
  .ZN({ S25957[1227] })
);
NAND2_X1 #() 
NAND2_X1_3516_ (
  .A1({ S15915 }),
  .A2({ S15948 }),
  .ZN({ S25957[1259] })
);
NAND3_X1 #() 
NAND3_X1_3715_ (
  .A1({ S20919 }),
  .A2({ S68 }),
  .A3({ S20776 }),
  .ZN({ S21095 })
);
NAND3_X1 #() 
NAND3_X1_3716_ (
  .A1({ S20802 }),
  .A2({ S20975 }),
  .A3({ S25957[1155] }),
  .ZN({ S21096 })
);
AOI21_X1 #() 
AOI21_X1_1896_ (
  .A({ S25957[1156] }),
  .B1({ S21096 }),
  .B2({ S21095 }),
  .ZN({ S21097 })
);
NAND3_X1 #() 
NAND3_X1_3717_ (
  .A1({ S21031 }),
  .A2({ S68 }),
  .A3({ S20776 }),
  .ZN({ S21098 })
);
NAND2_X1 #() 
NAND2_X1_3517_ (
  .A1({ S20793 }),
  .A2({ S20763 }),
  .ZN({ S21099 })
);
AOI21_X1 #() 
AOI21_X1_1897_ (
  .A({ S20774 }),
  .B1({ S21099 }),
  .B2({ S25957[1155] }),
  .ZN({ S21100 })
);
AND2_X1 #() 
AND2_X1_222_ (
  .A1({ S21100 }),
  .A2({ S21098 }),
  .ZN({ S21101 })
);
OAI21_X1 #() 
OAI21_X1_1822_ (
  .A({ S25957[1157] }),
  .B1({ S21101 }),
  .B2({ S21097 }),
  .ZN({ S21102 })
);
NAND2_X1 #() 
NAND2_X1_3518_ (
  .A1({ S20967 }),
  .A2({ S68 }),
  .ZN({ S21103 })
);
OAI21_X1 #() 
OAI21_X1_1823_ (
  .A({ S20977 }),
  .B1({ S21103 }),
  .B2({ S20809 }),
  .ZN({ S21104 })
);
NOR3_X1 #() 
NOR3_X1_122_ (
  .A1({ S20764 }),
  .A2({ S20842 }),
  .A3({ S25957[1156] }),
  .ZN({ S21105 })
);
AOI21_X1 #() 
AOI21_X1_1898_ (
  .A({ S21105 }),
  .B1({ S21104 }),
  .B2({ S25957[1156] }),
  .ZN({ S21106 })
);
OAI211_X1 #() 
OAI211_X1_1209_ (
  .A({ S21102 }),
  .B({ S25957[1158] }),
  .C1({ S21106 }),
  .C2({ S25957[1157] }),
  .ZN({ S21107 })
);
NAND2_X1 #() 
NAND2_X1_3519_ (
  .A1({ S20881 }),
  .A2({ S68 }),
  .ZN({ S21108 })
);
OAI211_X1 #() 
OAI211_X1_1210_ (
  .A({ S21108 }),
  .B({ S25957[1156] }),
  .C1({ S20992 }),
  .C2({ S20929 }),
  .ZN({ S21109 })
);
NAND2_X1 #() 
NAND2_X1_3520_ (
  .A1({ S20796 }),
  .A2({ S21050 }),
  .ZN({ S21110 })
);
AOI21_X1 #() 
AOI21_X1_1899_ (
  .A({ S68 }),
  .B1({ S20819 }),
  .B2({ S25957[1154] }),
  .ZN({ S21111 })
);
AOI21_X1 #() 
AOI21_X1_1900_ (
  .A({ S25957[1156] }),
  .B1({ S20914 }),
  .B2({ S21111 }),
  .ZN({ S21112 })
);
NAND2_X1 #() 
NAND2_X1_3521_ (
  .A1({ S21112 }),
  .A2({ S21110 }),
  .ZN({ S21113 })
);
AND2_X1 #() 
AND2_X1_223_ (
  .A1({ S21109 }),
  .A2({ S21113 }),
  .ZN({ S21114 })
);
NAND2_X1 #() 
NAND2_X1_3522_ (
  .A1({ S20780 }),
  .A2({ S20762 }),
  .ZN({ S21115 })
);
NAND2_X1 #() 
NAND2_X1_3523_ (
  .A1({ S21115 }),
  .A2({ S68 }),
  .ZN({ S21116 })
);
OAI211_X1 #() 
OAI211_X1_1211_ (
  .A({ S21116 }),
  .B({ S25957[1156] }),
  .C1({ S68 }),
  .C2({ S20794 }),
  .ZN({ S21117 })
);
NAND2_X1 #() 
NAND2_X1_3524_ (
  .A1({ S20793 }),
  .A2({ S20787 }),
  .ZN({ S21118 })
);
AOI22_X1 #() 
AOI22_X1_402_ (
  .A1({ S20828 }),
  .A2({ S20796 }),
  .B1({ S21118 }),
  .B2({ S68 }),
  .ZN({ S21119 })
);
NAND2_X1 #() 
NAND2_X1_3525_ (
  .A1({ S21119 }),
  .A2({ S20774 }),
  .ZN({ S21120 })
);
NAND3_X1 #() 
NAND3_X1_3718_ (
  .A1({ S21120 }),
  .A2({ S21117 }),
  .A3({ S20784 }),
  .ZN({ S21121 })
);
OAI211_X1 #() 
OAI211_X1_1212_ (
  .A({ S21121 }),
  .B({ S19194 }),
  .C1({ S21114 }),
  .C2({ S20784 }),
  .ZN({ S21122 })
);
NAND3_X1 #() 
NAND3_X1_3719_ (
  .A1({ S21122 }),
  .A2({ S21107 }),
  .A3({ S25957[1159] }),
  .ZN({ S21123 })
);
NAND3_X1 #() 
NAND3_X1_3720_ (
  .A1({ S20776 }),
  .A2({ S68 }),
  .A3({ S20785 }),
  .ZN({ S21124 })
);
NAND2_X1 #() 
NAND2_X1_3526_ (
  .A1({ S20948 }),
  .A2({ S20770 }),
  .ZN({ S21125 })
);
NAND3_X1 #() 
NAND3_X1_3721_ (
  .A1({ S21125 }),
  .A2({ S20774 }),
  .A3({ S21124 }),
  .ZN({ S21126 })
);
OAI211_X1 #() 
OAI211_X1_1213_ (
  .A({ S25957[1157] }),
  .B({ S21126 }),
  .C1({ S20839 }),
  .C2({ S20883 }),
  .ZN({ S21127 })
);
NAND3_X1 #() 
NAND3_X1_3722_ (
  .A1({ S20758 }),
  .A2({ S20787 }),
  .A3({ S68 }),
  .ZN({ S21128 })
);
INV_X1 #() 
INV_X1_1178_ (
  .A({ S21128 }),
  .ZN({ S21129 })
);
AOI22_X1 #() 
AOI22_X1_403_ (
  .A1({ S20790 }),
  .A2({ S21067 }),
  .B1({ S25957[1156] }),
  .B2({ S21129 }),
  .ZN({ S21130 })
);
OAI211_X1 #() 
OAI211_X1_1214_ (
  .A({ S21127 }),
  .B({ S25957[1158] }),
  .C1({ S21130 }),
  .C2({ S25957[1157] }),
  .ZN({ S21131 })
);
NAND4_X1 #() 
NAND4_X1_405_ (
  .A1({ S20932 }),
  .A2({ S20774 }),
  .A3({ S20785 }),
  .A4({ S25957[1152] }),
  .ZN({ S21132 })
);
NAND3_X1 #() 
NAND3_X1_3723_ (
  .A1({ S21103 }),
  .A2({ S25957[1156] }),
  .A3({ S20929 }),
  .ZN({ S21133 })
);
NAND2_X1 #() 
NAND2_X1_3527_ (
  .A1({ S21133 }),
  .A2({ S21132 }),
  .ZN({ S21134 })
);
OAI211_X1 #() 
OAI211_X1_1215_ (
  .A({ S25957[1155] }),
  .B({ S76 }),
  .C1({ S20758 }),
  .C2({ S25957[1154] }),
  .ZN({ S21135 })
);
NAND3_X1 #() 
NAND3_X1_3724_ (
  .A1({ S21135 }),
  .A2({ S20945 }),
  .A3({ S25957[1156] }),
  .ZN({ S21136 })
);
OAI211_X1 #() 
OAI211_X1_1216_ (
  .A({ S20780 }),
  .B({ S25957[1155] }),
  .C1({ S20819 }),
  .C2({ S20785 }),
  .ZN({ S21137 })
);
OAI211_X1 #() 
OAI211_X1_1217_ (
  .A({ S21137 }),
  .B({ S20774 }),
  .C1({ S20806 }),
  .C2({ S20855 }),
  .ZN({ S21138 })
);
NAND3_X1 #() 
NAND3_X1_3725_ (
  .A1({ S21138 }),
  .A2({ S20784 }),
  .A3({ S21136 }),
  .ZN({ S21139 })
);
OAI211_X1 #() 
OAI211_X1_1218_ (
  .A({ S19194 }),
  .B({ S21139 }),
  .C1({ S21134 }),
  .C2({ S20784 }),
  .ZN({ S21140 })
);
NAND3_X1 #() 
NAND3_X1_3726_ (
  .A1({ S21131 }),
  .A2({ S21140 }),
  .A3({ S19126 }),
  .ZN({ S21141 })
);
NAND3_X1 #() 
NAND3_X1_3727_ (
  .A1({ S21123 }),
  .A2({ S25957[1259] }),
  .A3({ S21141 }),
  .ZN({ S21142 })
);
INV_X1 #() 
INV_X1_1179_ (
  .A({ S25957[1259] }),
  .ZN({ S21143 })
);
INV_X1 #() 
INV_X1_1180_ (
  .A({ S21026 }),
  .ZN({ S21144 })
);
OAI211_X1 #() 
OAI211_X1_1219_ (
  .A({ S20985 }),
  .B({ S25957[1156] }),
  .C1({ S68 }),
  .C2({ S20776 }),
  .ZN({ S21145 })
);
OAI221_X1 #() 
OAI221_X1_107_ (
  .A({ S19194 }),
  .B1({ S21145 }),
  .B2({ S21144 }),
  .C1({ S21119 }),
  .C2({ S25957[1156] }),
  .ZN({ S21146 })
);
NAND2_X1 #() 
NAND2_X1_3528_ (
  .A1({ S21104 }),
  .A2({ S25957[1156] }),
  .ZN({ S21147 })
);
NOR2_X1 #() 
NOR2_X1_895_ (
  .A1({ S21105 }),
  .A2({ S19194 }),
  .ZN({ S21148 })
);
NAND2_X1 #() 
NAND2_X1_3529_ (
  .A1({ S21147 }),
  .A2({ S21148 }),
  .ZN({ S21149 })
);
AOI21_X1 #() 
AOI21_X1_1901_ (
  .A({ S19126 }),
  .B1({ S21149 }),
  .B2({ S21146 }),
  .ZN({ S21150 })
);
NAND2_X1 #() 
NAND2_X1_3530_ (
  .A1({ S21138 }),
  .A2({ S21136 }),
  .ZN({ S21151 })
);
NAND2_X1 #() 
NAND2_X1_3531_ (
  .A1({ S21151 }),
  .A2({ S19194 }),
  .ZN({ S21152 })
);
NAND2_X1 #() 
NAND2_X1_3532_ (
  .A1({ S20790 }),
  .A2({ S21067 }),
  .ZN({ S21153 })
);
NAND4_X1 #() 
NAND4_X1_406_ (
  .A1({ S25957[1156] }),
  .A2({ S20758 }),
  .A3({ S20787 }),
  .A4({ S68 }),
  .ZN({ S21154 })
);
NAND3_X1 #() 
NAND3_X1_3728_ (
  .A1({ S21153 }),
  .A2({ S25957[1158] }),
  .A3({ S21154 }),
  .ZN({ S21155 })
);
AOI21_X1 #() 
AOI21_X1_1902_ (
  .A({ S25957[1159] }),
  .B1({ S21155 }),
  .B2({ S21152 }),
  .ZN({ S21156 })
);
OAI21_X1 #() 
OAI21_X1_1824_ (
  .A({ S20784 }),
  .B1({ S21150 }),
  .B2({ S21156 }),
  .ZN({ S21157 })
);
NAND2_X1 #() 
NAND2_X1_3533_ (
  .A1({ S21134 }),
  .A2({ S19194 }),
  .ZN({ S21158 })
);
AOI22_X1 #() 
AOI22_X1_404_ (
  .A1({ S21032 }),
  .A2({ S20796 }),
  .B1({ S20881 }),
  .B2({ S25957[1155] }),
  .ZN({ S21159 })
);
NAND2_X1 #() 
NAND2_X1_3534_ (
  .A1({ S21125 }),
  .A2({ S21124 }),
  .ZN({ S21160 })
);
NAND2_X1 #() 
NAND2_X1_3535_ (
  .A1({ S21160 }),
  .A2({ S20774 }),
  .ZN({ S21161 })
);
OAI211_X1 #() 
OAI211_X1_1220_ (
  .A({ S21161 }),
  .B({ S25957[1158] }),
  .C1({ S21159 }),
  .C2({ S20774 }),
  .ZN({ S21162 })
);
AOI21_X1 #() 
AOI21_X1_1903_ (
  .A({ S25957[1159] }),
  .B1({ S21158 }),
  .B2({ S21162 }),
  .ZN({ S21163 })
);
NAND3_X1 #() 
NAND3_X1_3729_ (
  .A1({ S21109 }),
  .A2({ S19194 }),
  .A3({ S21113 }),
  .ZN({ S21164 })
);
NAND2_X1 #() 
NAND2_X1_3536_ (
  .A1({ S21096 }),
  .A2({ S21095 }),
  .ZN({ S21165 })
);
NAND2_X1 #() 
NAND2_X1_3537_ (
  .A1({ S21165 }),
  .A2({ S20774 }),
  .ZN({ S21166 })
);
AOI21_X1 #() 
AOI21_X1_1904_ (
  .A({ S19194 }),
  .B1({ S21100 }),
  .B2({ S21098 }),
  .ZN({ S21167 })
);
NAND2_X1 #() 
NAND2_X1_3538_ (
  .A1({ S21166 }),
  .A2({ S21167 }),
  .ZN({ S21168 })
);
AOI21_X1 #() 
AOI21_X1_1905_ (
  .A({ S19126 }),
  .B1({ S21168 }),
  .B2({ S21164 }),
  .ZN({ S21169 })
);
OAI21_X1 #() 
OAI21_X1_1825_ (
  .A({ S25957[1157] }),
  .B1({ S21163 }),
  .B2({ S21169 }),
  .ZN({ S21170 })
);
NAND3_X1 #() 
NAND3_X1_3730_ (
  .A1({ S21157 }),
  .A2({ S21170 }),
  .A3({ S21143 }),
  .ZN({ S21171 })
);
NAND3_X1 #() 
NAND3_X1_3731_ (
  .A1({ S21171 }),
  .A2({ S21142 }),
  .A3({ S25957[1227] }),
  .ZN({ S21172 })
);
INV_X1 #() 
INV_X1_1181_ (
  .A({ S25957[1227] }),
  .ZN({ S21173 })
);
NAND3_X1 #() 
NAND3_X1_3732_ (
  .A1({ S21123 }),
  .A2({ S21143 }),
  .A3({ S21141 }),
  .ZN({ S21174 })
);
NAND3_X1 #() 
NAND3_X1_3733_ (
  .A1({ S21157 }),
  .A2({ S21170 }),
  .A3({ S25957[1259] }),
  .ZN({ S21175 })
);
NAND3_X1 #() 
NAND3_X1_3734_ (
  .A1({ S21175 }),
  .A2({ S21174 }),
  .A3({ S21173 }),
  .ZN({ S21176 })
);
NAND3_X1 #() 
NAND3_X1_3735_ (
  .A1({ S21172 }),
  .A2({ S21176 }),
  .A3({ S21094 }),
  .ZN({ S21177 })
);
NAND3_X1 #() 
NAND3_X1_3736_ (
  .A1({ S21171 }),
  .A2({ S21142 }),
  .A3({ S21173 }),
  .ZN({ S21178 })
);
NAND3_X1 #() 
NAND3_X1_3737_ (
  .A1({ S21175 }),
  .A2({ S21174 }),
  .A3({ S25957[1227] }),
  .ZN({ S21179 })
);
NAND3_X1 #() 
NAND3_X1_3738_ (
  .A1({ S21178 }),
  .A2({ S21179 }),
  .A3({ S25957[1195] }),
  .ZN({ S21180 })
);
NAND3_X1 #() 
NAND3_X1_3739_ (
  .A1({ S21177 }),
  .A2({ S21180 }),
  .A3({ S65 }),
  .ZN({ S21181 })
);
NAND3_X1 #() 
NAND3_X1_3740_ (
  .A1({ S21172 }),
  .A2({ S21176 }),
  .A3({ S25957[1195] }),
  .ZN({ S21182 })
);
NAND3_X1 #() 
NAND3_X1_3741_ (
  .A1({ S21178 }),
  .A2({ S21179 }),
  .A3({ S21094 }),
  .ZN({ S21183 })
);
NAND3_X1 #() 
NAND3_X1_3742_ (
  .A1({ S21182 }),
  .A2({ S21183 }),
  .A3({ S25957[1163] }),
  .ZN({ S21184 })
);
NAND2_X1 #() 
NAND2_X1_3539_ (
  .A1({ S21181 }),
  .A2({ S21184 }),
  .ZN({ S77 })
);
NAND3_X1 #() 
NAND3_X1_3743_ (
  .A1({ S21182 }),
  .A2({ S21183 }),
  .A3({ S65 }),
  .ZN({ S21185 })
);
NAND3_X1 #() 
NAND3_X1_3744_ (
  .A1({ S21177 }),
  .A2({ S21180 }),
  .A3({ S25957[1163] }),
  .ZN({ S21186 })
);
NAND2_X1 #() 
NAND2_X1_3540_ (
  .A1({ S21185 }),
  .A2({ S21186 }),
  .ZN({ S25957[1035] })
);
NAND2_X1 #() 
NAND2_X1_3541_ (
  .A1({ S16538 }),
  .A2({ S16549 }),
  .ZN({ S25957[1224] })
);
INV_X1 #() 
INV_X1_1182_ (
  .A({ S25957[1224] }),
  .ZN({ S21187 })
);
NAND2_X1 #() 
NAND2_X1_3542_ (
  .A1({ S16462 }),
  .A2({ S16440 }),
  .ZN({ S25957[1256] })
);
NAND2_X1 #() 
NAND2_X1_3543_ (
  .A1({ S20926 }),
  .A2({ S25957[1155] }),
  .ZN({ S21188 })
);
NAND4_X1 #() 
NAND4_X1_407_ (
  .A1({ S20975 }),
  .A2({ S20895 }),
  .A3({ S20766 }),
  .A4({ S25957[1155] }),
  .ZN({ S21189 })
);
AOI21_X1 #() 
AOI21_X1_1906_ (
  .A({ S20774 }),
  .B1({ S20919 }),
  .B2({ S68 }),
  .ZN({ S21190 })
);
AOI22_X1 #() 
AOI22_X1_405_ (
  .A1({ S20863 }),
  .A2({ S21188 }),
  .B1({ S21190 }),
  .B2({ S21189 }),
  .ZN({ S21191 })
);
NAND3_X1 #() 
NAND3_X1_3745_ (
  .A1({ S20976 }),
  .A2({ S20774 }),
  .A3({ S20953 }),
  .ZN({ S21192 })
);
NAND4_X1 #() 
NAND4_X1_408_ (
  .A1({ S20949 }),
  .A2({ S20891 }),
  .A3({ S20778 }),
  .A4({ S25957[1156] }),
  .ZN({ S21193 })
);
NAND3_X1 #() 
NAND3_X1_3746_ (
  .A1({ S21192 }),
  .A2({ S20784 }),
  .A3({ S21193 }),
  .ZN({ S21194 })
);
OAI211_X1 #() 
OAI211_X1_1221_ (
  .A({ S25957[1158] }),
  .B({ S21194 }),
  .C1({ S21191 }),
  .C2({ S20784 }),
  .ZN({ S21195 })
);
AOI21_X1 #() 
AOI21_X1_1907_ (
  .A({ S25957[1155] }),
  .B1({ S20975 }),
  .B2({ S20895 }),
  .ZN({ S21196 })
);
NOR2_X1 #() 
NOR2_X1_896_ (
  .A1({ S21145 }),
  .A2({ S21196 }),
  .ZN({ S21197 })
);
NAND3_X1 #() 
NAND3_X1_3747_ (
  .A1({ S20904 }),
  .A2({ S20950 }),
  .A3({ S25957[1156] }),
  .ZN({ S21198 })
);
NAND3_X1 #() 
NAND3_X1_3748_ (
  .A1({ S20969 }),
  .A2({ S20878 }),
  .A3({ S20774 }),
  .ZN({ S21199 })
);
NAND3_X1 #() 
NAND3_X1_3749_ (
  .A1({ S21199 }),
  .A2({ S21198 }),
  .A3({ S25957[1157] }),
  .ZN({ S21200 })
);
AOI21_X1 #() 
AOI21_X1_1908_ (
  .A({ S68 }),
  .B1({ S20895 }),
  .B2({ S76 }),
  .ZN({ S21201 })
);
NAND2_X1 #() 
NAND2_X1_3544_ (
  .A1({ S20766 }),
  .A2({ S20785 }),
  .ZN({ S21202 })
);
NAND3_X1 #() 
NAND3_X1_3750_ (
  .A1({ S20787 }),
  .A2({ S68 }),
  .A3({ S20770 }),
  .ZN({ S21203 })
);
OAI21_X1 #() 
OAI21_X1_1826_ (
  .A({ S20774 }),
  .B1({ S21203 }),
  .B2({ S21202 }),
  .ZN({ S21204 })
);
OAI21_X1 #() 
OAI21_X1_1827_ (
  .A({ S20784 }),
  .B1({ S21204 }),
  .B2({ S21201 }),
  .ZN({ S21205 })
);
OAI211_X1 #() 
OAI211_X1_1222_ (
  .A({ S21200 }),
  .B({ S19194 }),
  .C1({ S21205 }),
  .C2({ S21197 }),
  .ZN({ S21206 })
);
NAND3_X1 #() 
NAND3_X1_3751_ (
  .A1({ S21195 }),
  .A2({ S21206 }),
  .A3({ S19126 }),
  .ZN({ S21207 })
);
OAI21_X1 #() 
OAI21_X1_1828_ (
  .A({ S25957[1155] }),
  .B1({ S21202 }),
  .B2({ S20803 }),
  .ZN({ S21208 })
);
NAND2_X1 #() 
NAND2_X1_3545_ (
  .A1({ S20830 }),
  .A2({ S21057 }),
  .ZN({ S21209 })
);
NAND3_X1 #() 
NAND3_X1_3752_ (
  .A1({ S21209 }),
  .A2({ S21208 }),
  .A3({ S20774 }),
  .ZN({ S21210 })
);
AOI21_X1 #() 
AOI21_X1_1909_ (
  .A({ S25957[1155] }),
  .B1({ S20818 }),
  .B2({ S20820 }),
  .ZN({ S21211 })
);
NOR2_X1 #() 
NOR2_X1_897_ (
  .A1({ S21056 }),
  .A2({ S68 }),
  .ZN({ S21212 })
);
OAI21_X1 #() 
OAI21_X1_1829_ (
  .A({ S25957[1156] }),
  .B1({ S21211 }),
  .B2({ S21212 }),
  .ZN({ S21213 })
);
AOI21_X1 #() 
AOI21_X1_1910_ (
  .A({ S20784 }),
  .B1({ S21213 }),
  .B2({ S21210 }),
  .ZN({ S21214 })
);
NOR2_X1 #() 
NOR2_X1_898_ (
  .A1({ S20967 }),
  .A2({ S68 }),
  .ZN({ S21215 })
);
AOI21_X1 #() 
AOI21_X1_1911_ (
  .A({ S21215 }),
  .B1({ S21038 }),
  .B2({ S21037 }),
  .ZN({ S21216 })
);
OAI21_X1 #() 
OAI21_X1_1830_ (
  .A({ S20784 }),
  .B1({ S21059 }),
  .B2({ S20964 }),
  .ZN({ S21217 })
);
OAI21_X1 #() 
OAI21_X1_1831_ (
  .A({ S25957[1158] }),
  .B1({ S21216 }),
  .B2({ S21217 }),
  .ZN({ S21218 })
);
NAND3_X1 #() 
NAND3_X1_3753_ (
  .A1({ S21044 }),
  .A2({ S20774 }),
  .A3({ S21016 }),
  .ZN({ S21219 })
);
NAND3_X1 #() 
NAND3_X1_3754_ (
  .A1({ S20770 }),
  .A2({ S20819 }),
  .A3({ S68 }),
  .ZN({ S21220 })
);
OR2_X1 #() 
OR2_X1_47_ (
  .A1({ S21220 }),
  .A2({ S20774 }),
  .ZN({ S21221 })
);
NAND3_X1 #() 
NAND3_X1_3755_ (
  .A1({ S20929 }),
  .A2({ S21128 }),
  .A3({ S25957[1156] }),
  .ZN({ S21222 })
);
NAND4_X1 #() 
NAND4_X1_409_ (
  .A1({ S21219 }),
  .A2({ S21221 }),
  .A3({ S25957[1157] }),
  .A4({ S21222 }),
  .ZN({ S21223 })
);
NAND2_X1 #() 
NAND2_X1_3546_ (
  .A1({ S25957[1155] }),
  .A2({ S20770 }),
  .ZN({ S21224 })
);
OAI211_X1 #() 
OAI211_X1_1223_ (
  .A({ S25957[1156] }),
  .B({ S21224 }),
  .C1({ S20992 }),
  .C2({ S25957[1155] }),
  .ZN({ S21225 })
);
NAND4_X1 #() 
NAND4_X1_410_ (
  .A1({ S20766 }),
  .A2({ S76 }),
  .A3({ S20787 }),
  .A4({ S68 }),
  .ZN({ S21226 })
);
NAND3_X1 #() 
NAND3_X1_3756_ (
  .A1({ S21226 }),
  .A2({ S21125 }),
  .A3({ S20774 }),
  .ZN({ S21227 })
);
NAND3_X1 #() 
NAND3_X1_3757_ (
  .A1({ S21225 }),
  .A2({ S20784 }),
  .A3({ S21227 }),
  .ZN({ S21228 })
);
NAND3_X1 #() 
NAND3_X1_3758_ (
  .A1({ S21223 }),
  .A2({ S19194 }),
  .A3({ S21228 }),
  .ZN({ S21229 })
);
OAI211_X1 #() 
OAI211_X1_1224_ (
  .A({ S21229 }),
  .B({ S25957[1159] }),
  .C1({ S21214 }),
  .C2({ S21218 }),
  .ZN({ S21230 })
);
NAND3_X1 #() 
NAND3_X1_3759_ (
  .A1({ S21230 }),
  .A2({ S25957[1256] }),
  .A3({ S21207 }),
  .ZN({ S21231 })
);
INV_X1 #() 
INV_X1_1183_ (
  .A({ S25957[1256] }),
  .ZN({ S21232 })
);
AOI21_X1 #() 
AOI21_X1_1912_ (
  .A({ S25957[1155] }),
  .B1({ S20802 }),
  .B2({ S20975 }),
  .ZN({ S21233 })
);
OAI21_X1 #() 
OAI21_X1_1832_ (
  .A({ S25957[1156] }),
  .B1({ S21215 }),
  .B2({ S21233 }),
  .ZN({ S21234 })
);
NAND2_X1 #() 
NAND2_X1_3547_ (
  .A1({ S20953 }),
  .A2({ S20963 }),
  .ZN({ S21235 })
);
NAND2_X1 #() 
NAND2_X1_3548_ (
  .A1({ S21235 }),
  .A2({ S20774 }),
  .ZN({ S21236 })
);
NAND3_X1 #() 
NAND3_X1_3760_ (
  .A1({ S21234 }),
  .A2({ S20784 }),
  .A3({ S21236 }),
  .ZN({ S21237 })
);
NAND3_X1 #() 
NAND3_X1_3761_ (
  .A1({ S21213 }),
  .A2({ S21210 }),
  .A3({ S25957[1157] }),
  .ZN({ S21238 })
);
NAND3_X1 #() 
NAND3_X1_3762_ (
  .A1({ S21237 }),
  .A2({ S21238 }),
  .A3({ S25957[1158] }),
  .ZN({ S21239 })
);
NAND2_X1 #() 
NAND2_X1_3549_ (
  .A1({ S21225 }),
  .A2({ S21227 }),
  .ZN({ S21240 })
);
NAND2_X1 #() 
NAND2_X1_3550_ (
  .A1({ S21240 }),
  .A2({ S20784 }),
  .ZN({ S21241 })
);
OAI211_X1 #() 
OAI211_X1_1225_ (
  .A({ S25957[1156] }),
  .B({ S21220 }),
  .C1({ S20886 }),
  .C2({ S21129 }),
  .ZN({ S21242 })
);
AOI21_X1 #() 
AOI21_X1_1913_ (
  .A({ S68 }),
  .B1({ S20777 }),
  .B2({ S21031 }),
  .ZN({ S21243 })
);
OAI21_X1 #() 
OAI21_X1_1833_ (
  .A({ S20774 }),
  .B1({ S21243 }),
  .B2({ S21017 }),
  .ZN({ S21244 })
);
NAND3_X1 #() 
NAND3_X1_3763_ (
  .A1({ S21244 }),
  .A2({ S21242 }),
  .A3({ S25957[1157] }),
  .ZN({ S21245 })
);
NAND3_X1 #() 
NAND3_X1_3764_ (
  .A1({ S21245 }),
  .A2({ S21241 }),
  .A3({ S19194 }),
  .ZN({ S21246 })
);
NAND3_X1 #() 
NAND3_X1_3765_ (
  .A1({ S21239 }),
  .A2({ S21246 }),
  .A3({ S25957[1159] }),
  .ZN({ S21247 })
);
NAND2_X1 #() 
NAND2_X1_3551_ (
  .A1({ S21192 }),
  .A2({ S21193 }),
  .ZN({ S21248 })
);
NAND2_X1 #() 
NAND2_X1_3552_ (
  .A1({ S21248 }),
  .A2({ S20784 }),
  .ZN({ S21249 })
);
NAND2_X1 #() 
NAND2_X1_3553_ (
  .A1({ S21190 }),
  .A2({ S21189 }),
  .ZN({ S21250 })
);
NAND2_X1 #() 
NAND2_X1_3554_ (
  .A1({ S21188 }),
  .A2({ S20863 }),
  .ZN({ S21251 })
);
NAND3_X1 #() 
NAND3_X1_3766_ (
  .A1({ S21251 }),
  .A2({ S21250 }),
  .A3({ S25957[1157] }),
  .ZN({ S21252 })
);
NAND3_X1 #() 
NAND3_X1_3767_ (
  .A1({ S21249 }),
  .A2({ S21252 }),
  .A3({ S25957[1158] }),
  .ZN({ S21253 })
);
OAI21_X1 #() 
OAI21_X1_1834_ (
  .A({ S21200 }),
  .B1({ S21205 }),
  .B2({ S21197 }),
  .ZN({ S21254 })
);
NAND2_X1 #() 
NAND2_X1_3555_ (
  .A1({ S21254 }),
  .A2({ S19194 }),
  .ZN({ S21255 })
);
NAND3_X1 #() 
NAND3_X1_3768_ (
  .A1({ S21255 }),
  .A2({ S19126 }),
  .A3({ S21253 }),
  .ZN({ S21256 })
);
NAND3_X1 #() 
NAND3_X1_3769_ (
  .A1({ S21247 }),
  .A2({ S21256 }),
  .A3({ S21232 }),
  .ZN({ S21257 })
);
NAND3_X1 #() 
NAND3_X1_3770_ (
  .A1({ S21257 }),
  .A2({ S21231 }),
  .A3({ S21187 }),
  .ZN({ S21258 })
);
NAND3_X1 #() 
NAND3_X1_3771_ (
  .A1({ S21230 }),
  .A2({ S21232 }),
  .A3({ S21207 }),
  .ZN({ S21259 })
);
NAND3_X1 #() 
NAND3_X1_3772_ (
  .A1({ S21247 }),
  .A2({ S21256 }),
  .A3({ S25957[1256] }),
  .ZN({ S21260 })
);
NAND3_X1 #() 
NAND3_X1_3773_ (
  .A1({ S21260 }),
  .A2({ S21259 }),
  .A3({ S25957[1224] }),
  .ZN({ S21261 })
);
AOI21_X1 #() 
AOI21_X1_1914_ (
  .A({ S5639 }),
  .B1({ S21258 }),
  .B2({ S21261 }),
  .ZN({ S21262 })
);
NAND3_X1 #() 
NAND3_X1_3774_ (
  .A1({ S21257 }),
  .A2({ S21231 }),
  .A3({ S25957[1224] }),
  .ZN({ S21263 })
);
NAND3_X1 #() 
NAND3_X1_3775_ (
  .A1({ S21260 }),
  .A2({ S21259 }),
  .A3({ S21187 }),
  .ZN({ S21264 })
);
AOI21_X1 #() 
AOI21_X1_1915_ (
  .A({ S25956[8] }),
  .B1({ S21263 }),
  .B2({ S21264 }),
  .ZN({ S21265 })
);
NOR2_X1 #() 
NOR2_X1_899_ (
  .A1({ S21262 }),
  .A2({ S21265 }),
  .ZN({ S25957[1032] })
);
NAND2_X1 #() 
NAND2_X1_3556_ (
  .A1({ S17262 }),
  .A2({ S17273 }),
  .ZN({ S25957[1225] })
);
INV_X1 #() 
INV_X1_1184_ (
  .A({ S25957[1225] }),
  .ZN({ S21266 })
);
NAND2_X1 #() 
NAND2_X1_3557_ (
  .A1({ S17186 }),
  .A2({ S17078 }),
  .ZN({ S25957[1257] })
);
OAI211_X1 #() 
OAI211_X1_1226_ (
  .A({ S25957[1156] }),
  .B({ S21220 }),
  .C1({ S20946 }),
  .C2({ S20944 }),
  .ZN({ S21267 })
);
NAND2_X1 #() 
NAND2_X1_3558_ (
  .A1({ S20820 }),
  .A2({ S68 }),
  .ZN({ S21268 })
);
NAND2_X1 #() 
NAND2_X1_3559_ (
  .A1({ S20758 }),
  .A2({ S20787 }),
  .ZN({ S21269 })
);
NAND3_X1 #() 
NAND3_X1_3776_ (
  .A1({ S20758 }),
  .A2({ S20780 }),
  .A3({ S25957[1155] }),
  .ZN({ S21270 })
);
OAI211_X1 #() 
OAI211_X1_1227_ (
  .A({ S20774 }),
  .B({ S21270 }),
  .C1({ S21268 }),
  .C2({ S21269 }),
  .ZN({ S21271 })
);
NAND3_X1 #() 
NAND3_X1_3777_ (
  .A1({ S21267 }),
  .A2({ S21271 }),
  .A3({ S20784 }),
  .ZN({ S21272 })
);
AOI21_X1 #() 
AOI21_X1_1916_ (
  .A({ S68 }),
  .B1({ S20796 }),
  .B2({ S20956 }),
  .ZN({ S21273 })
);
NAND3_X1 #() 
NAND3_X1_3778_ (
  .A1({ S20781 }),
  .A2({ S20977 }),
  .A3({ S25957[1156] }),
  .ZN({ S21274 })
);
NAND2_X1 #() 
NAND2_X1_3560_ (
  .A1({ S20771 }),
  .A2({ S20774 }),
  .ZN({ S21275 })
);
OAI211_X1 #() 
OAI211_X1_1228_ (
  .A({ S25957[1157] }),
  .B({ S21274 }),
  .C1({ S21273 }),
  .C2({ S21275 }),
  .ZN({ S21276 })
);
NAND3_X1 #() 
NAND3_X1_3779_ (
  .A1({ S21272 }),
  .A2({ S21276 }),
  .A3({ S25957[1158] }),
  .ZN({ S21277 })
);
NAND3_X1 #() 
NAND3_X1_3780_ (
  .A1({ S21124 }),
  .A2({ S20985 }),
  .A3({ S20774 }),
  .ZN({ S21278 })
);
AOI21_X1 #() 
AOI21_X1_1917_ (
  .A({ S68 }),
  .B1({ S20967 }),
  .B2({ S20766 }),
  .ZN({ S21279 })
);
OAI211_X1 #() 
OAI211_X1_1229_ (
  .A({ S25957[1157] }),
  .B({ S21278 }),
  .C1({ S21279 }),
  .C2({ S20772 }),
  .ZN({ S21280 })
);
OAI21_X1 #() 
OAI21_X1_1835_ (
  .A({ S20774 }),
  .B1({ S20963 }),
  .B2({ S20983 }),
  .ZN({ S21281 })
);
NAND2_X1 #() 
NAND2_X1_3561_ (
  .A1({ S20786 }),
  .A2({ S25957[1155] }),
  .ZN({ S21282 })
);
OAI211_X1 #() 
OAI211_X1_1230_ (
  .A({ S25957[1156] }),
  .B({ S21282 }),
  .C1({ S20892 }),
  .C2({ S25957[1155] }),
  .ZN({ S21283 })
);
OAI211_X1 #() 
OAI211_X1_1231_ (
  .A({ S21283 }),
  .B({ S20784 }),
  .C1({ S21281 }),
  .C2({ S20795 }),
  .ZN({ S21284 })
);
NAND3_X1 #() 
NAND3_X1_3781_ (
  .A1({ S21284 }),
  .A2({ S21280 }),
  .A3({ S19194 }),
  .ZN({ S21285 })
);
NAND3_X1 #() 
NAND3_X1_3782_ (
  .A1({ S21285 }),
  .A2({ S21277 }),
  .A3({ S25957[1159] }),
  .ZN({ S21286 })
);
AOI21_X1 #() 
AOI21_X1_1918_ (
  .A({ S20788 }),
  .B1({ S76 }),
  .B2({ S20849 }),
  .ZN({ S21287 })
);
NOR2_X1 #() 
NOR2_X1_900_ (
  .A1({ S20778 }),
  .A2({ S25957[1152] }),
  .ZN({ S21288 })
);
OAI21_X1 #() 
OAI21_X1_1836_ (
  .A({ S25957[1156] }),
  .B1({ S21288 }),
  .B2({ S20855 }),
  .ZN({ S21289 })
);
AOI21_X1 #() 
AOI21_X1_1919_ (
  .A({ S20817 }),
  .B1({ S20919 }),
  .B2({ S20763 }),
  .ZN({ S21290 })
);
AOI21_X1 #() 
AOI21_X1_1920_ (
  .A({ S20784 }),
  .B1({ S21290 }),
  .B2({ S20774 }),
  .ZN({ S21291 })
);
OAI21_X1 #() 
OAI21_X1_1837_ (
  .A({ S21291 }),
  .B1({ S21287 }),
  .B2({ S21289 }),
  .ZN({ S21292 })
);
OAI21_X1 #() 
OAI21_X1_1838_ (
  .A({ S25957[1156] }),
  .B1({ S21268 }),
  .B2({ S20896 }),
  .ZN({ S21293 })
);
OAI211_X1 #() 
OAI211_X1_1232_ (
  .A({ S20912 }),
  .B({ S20774 }),
  .C1({ S20967 }),
  .C2({ S68 }),
  .ZN({ S21294 })
);
OAI211_X1 #() 
OAI211_X1_1233_ (
  .A({ S21294 }),
  .B({ S20784 }),
  .C1({ S21293 }),
  .C2({ S21273 }),
  .ZN({ S21295 })
);
NAND3_X1 #() 
NAND3_X1_3783_ (
  .A1({ S21295 }),
  .A2({ S21292 }),
  .A3({ S25957[1158] }),
  .ZN({ S21296 })
);
NAND2_X1 #() 
NAND2_X1_3562_ (
  .A1({ S20914 }),
  .A2({ S21111 }),
  .ZN({ S21297 })
);
AOI21_X1 #() 
AOI21_X1_1921_ (
  .A({ S20774 }),
  .B1({ S21297 }),
  .B2({ S21019 }),
  .ZN({ S21298 })
);
OAI21_X1 #() 
OAI21_X1_1839_ (
  .A({ S25957[1157] }),
  .B1({ S21298 }),
  .B2({ S20790 }),
  .ZN({ S21299 })
);
NAND4_X1 #() 
NAND4_X1_411_ (
  .A1({ S21026 }),
  .A2({ S20804 }),
  .A3({ S20860 }),
  .A4({ S25957[1156] }),
  .ZN({ S21300 })
);
OAI211_X1 #() 
OAI211_X1_1234_ (
  .A({ S20852 }),
  .B({ S20774 }),
  .C1({ S20781 }),
  .C2({ S21202 }),
  .ZN({ S21301 })
);
NAND3_X1 #() 
NAND3_X1_3784_ (
  .A1({ S21301 }),
  .A2({ S21300 }),
  .A3({ S20784 }),
  .ZN({ S21302 })
);
NAND3_X1 #() 
NAND3_X1_3785_ (
  .A1({ S21299 }),
  .A2({ S21302 }),
  .A3({ S19194 }),
  .ZN({ S21303 })
);
NAND3_X1 #() 
NAND3_X1_3786_ (
  .A1({ S21296 }),
  .A2({ S21303 }),
  .A3({ S19126 }),
  .ZN({ S21304 })
);
NAND3_X1 #() 
NAND3_X1_3787_ (
  .A1({ S21304 }),
  .A2({ S21286 }),
  .A3({ S25957[1257] }),
  .ZN({ S21305 })
);
INV_X1 #() 
INV_X1_1185_ (
  .A({ S25957[1257] }),
  .ZN({ S21306 })
);
NAND2_X1 #() 
NAND2_X1_3563_ (
  .A1({ S21304 }),
  .A2({ S21286 }),
  .ZN({ S21307 })
);
NAND2_X1 #() 
NAND2_X1_3564_ (
  .A1({ S21307 }),
  .A2({ S21306 }),
  .ZN({ S21308 })
);
NAND3_X1 #() 
NAND3_X1_3788_ (
  .A1({ S21308 }),
  .A2({ S21266 }),
  .A3({ S21305 }),
  .ZN({ S21309 })
);
NAND3_X1 #() 
NAND3_X1_3789_ (
  .A1({ S21304 }),
  .A2({ S21286 }),
  .A3({ S21306 }),
  .ZN({ S21310 })
);
NAND2_X1 #() 
NAND2_X1_3565_ (
  .A1({ S21307 }),
  .A2({ S25957[1257] }),
  .ZN({ S21311 })
);
NAND3_X1 #() 
NAND3_X1_3790_ (
  .A1({ S21311 }),
  .A2({ S25957[1225] }),
  .A3({ S21310 }),
  .ZN({ S21312 })
);
AOI21_X1 #() 
AOI21_X1_1922_ (
  .A({ S5628 }),
  .B1({ S21309 }),
  .B2({ S21312 }),
  .ZN({ S21313 })
);
NAND3_X1 #() 
NAND3_X1_3791_ (
  .A1({ S21308 }),
  .A2({ S25957[1225] }),
  .A3({ S21305 }),
  .ZN({ S21314 })
);
NAND3_X1 #() 
NAND3_X1_3792_ (
  .A1({ S21311 }),
  .A2({ S21266 }),
  .A3({ S21310 }),
  .ZN({ S21315 })
);
AOI21_X1 #() 
AOI21_X1_1923_ (
  .A({ S25956[9] }),
  .B1({ S21314 }),
  .B2({ S21315 }),
  .ZN({ S21316 })
);
NOR2_X1 #() 
NOR2_X1_901_ (
  .A1({ S21313 }),
  .A2({ S21316 }),
  .ZN({ S25957[1033] })
);
NAND2_X1 #() 
NAND2_X1_3566_ (
  .A1({ S17911 }),
  .A2({ S17922 }),
  .ZN({ S21317 })
);
INV_X1 #() 
INV_X1_1186_ (
  .A({ S21317 }),
  .ZN({ S25957[1258] })
);
NAND3_X1 #() 
NAND3_X1_3793_ (
  .A1({ S21057 }),
  .A2({ S25957[1155] }),
  .A3({ S21056 }),
  .ZN({ S21318 })
);
NAND3_X1 #() 
NAND3_X1_3794_ (
  .A1({ S21318 }),
  .A2({ S20774 }),
  .A3({ S20931 }),
  .ZN({ S21319 })
);
NAND3_X1 #() 
NAND3_X1_3795_ (
  .A1({ S20849 }),
  .A2({ S68 }),
  .A3({ S76 }),
  .ZN({ S21320 })
);
AOI21_X1 #() 
AOI21_X1_1924_ (
  .A({ S20774 }),
  .B1({ S21115 }),
  .B2({ S25957[1155] }),
  .ZN({ S21321 })
);
AOI21_X1 #() 
AOI21_X1_1925_ (
  .A({ S20784 }),
  .B1({ S21321 }),
  .B2({ S21320 }),
  .ZN({ S21322 })
);
NAND2_X1 #() 
NAND2_X1_3567_ (
  .A1({ S21322 }),
  .A2({ S21319 }),
  .ZN({ S21323 })
);
NAND2_X1 #() 
NAND2_X1_3568_ (
  .A1({ S20807 }),
  .A2({ S68 }),
  .ZN({ S21324 })
);
NAND3_X1 #() 
NAND3_X1_3796_ (
  .A1({ S21025 }),
  .A2({ S21324 }),
  .A3({ S20774 }),
  .ZN({ S21325 })
);
NAND2_X1 #() 
NAND2_X1_3569_ (
  .A1({ S20850 }),
  .A2({ S21111 }),
  .ZN({ S21326 })
);
NAND2_X1 #() 
NAND2_X1_3570_ (
  .A1({ S21326 }),
  .A2({ S20995 }),
  .ZN({ S21327 })
);
NAND3_X1 #() 
NAND3_X1_3797_ (
  .A1({ S21327 }),
  .A2({ S21325 }),
  .A3({ S20784 }),
  .ZN({ S21328 })
);
NAND3_X1 #() 
NAND3_X1_3798_ (
  .A1({ S21328 }),
  .A2({ S21323 }),
  .A3({ S25957[1158] }),
  .ZN({ S21329 })
);
NAND3_X1 #() 
NAND3_X1_3799_ (
  .A1({ S25957[1155] }),
  .A2({ S20762 }),
  .A3({ S25957[1152] }),
  .ZN({ S21330 })
);
OAI211_X1 #() 
OAI211_X1_1235_ (
  .A({ S25957[1156] }),
  .B({ S21330 }),
  .C1({ S20781 }),
  .C2({ S21202 }),
  .ZN({ S21331 })
);
NAND3_X1 #() 
NAND3_X1_3800_ (
  .A1({ S25957[1155] }),
  .A2({ S25957[1152] }),
  .A3({ S25957[1153] }),
  .ZN({ S21332 })
);
NAND4_X1 #() 
NAND4_X1_412_ (
  .A1({ S21040 }),
  .A2({ S21203 }),
  .A3({ S21332 }),
  .A4({ S20774 }),
  .ZN({ S21333 })
);
NAND3_X1 #() 
NAND3_X1_3801_ (
  .A1({ S21331 }),
  .A2({ S21333 }),
  .A3({ S25957[1157] }),
  .ZN({ S21334 })
);
OAI211_X1 #() 
OAI211_X1_1236_ (
  .A({ S20899 }),
  .B({ S20774 }),
  .C1({ S20891 }),
  .C2({ S25957[1155] }),
  .ZN({ S21335 })
);
NAND2_X1 #() 
NAND2_X1_3571_ (
  .A1({ S20785 }),
  .A2({ S68 }),
  .ZN({ S21336 })
);
NAND3_X1 #() 
NAND3_X1_3802_ (
  .A1({ S20763 }),
  .A2({ S25957[1155] }),
  .A3({ S25957[1153] }),
  .ZN({ S21337 })
);
NAND3_X1 #() 
NAND3_X1_3803_ (
  .A1({ S21337 }),
  .A2({ S25957[1156] }),
  .A3({ S21336 }),
  .ZN({ S21338 })
);
NAND3_X1 #() 
NAND3_X1_3804_ (
  .A1({ S21335 }),
  .A2({ S21338 }),
  .A3({ S20784 }),
  .ZN({ S21339 })
);
NAND3_X1 #() 
NAND3_X1_3805_ (
  .A1({ S21334 }),
  .A2({ S21339 }),
  .A3({ S19194 }),
  .ZN({ S21340 })
);
NAND3_X1 #() 
NAND3_X1_3806_ (
  .A1({ S21329 }),
  .A2({ S25957[1159] }),
  .A3({ S21340 }),
  .ZN({ S21341 })
);
NAND3_X1 #() 
NAND3_X1_3807_ (
  .A1({ S20831 }),
  .A2({ S25957[1155] }),
  .A3({ S20895 }),
  .ZN({ S21342 })
);
NAND3_X1 #() 
NAND3_X1_3808_ (
  .A1({ S21342 }),
  .A2({ S20774 }),
  .A3({ S20900 }),
  .ZN({ S21343 })
);
OAI211_X1 #() 
OAI211_X1_1237_ (
  .A({ S20787 }),
  .B({ S25957[1155] }),
  .C1({ S20762 }),
  .C2({ S25957[1152] }),
  .ZN({ S21344 })
);
OAI211_X1 #() 
OAI211_X1_1238_ (
  .A({ S25957[1156] }),
  .B({ S21344 }),
  .C1({ S20806 }),
  .C2({ S21049 }),
  .ZN({ S21345 })
);
NAND3_X1 #() 
NAND3_X1_3809_ (
  .A1({ S21343 }),
  .A2({ S21345 }),
  .A3({ S25957[1157] }),
  .ZN({ S21346 })
);
OAI211_X1 #() 
OAI211_X1_1239_ (
  .A({ S21337 }),
  .B({ S25957[1156] }),
  .C1({ S20771 }),
  .C2({ S21053 }),
  .ZN({ S21347 })
);
NAND3_X1 #() 
NAND3_X1_3810_ (
  .A1({ S21188 }),
  .A2({ S21209 }),
  .A3({ S20774 }),
  .ZN({ S21348 })
);
NAND3_X1 #() 
NAND3_X1_3811_ (
  .A1({ S21348 }),
  .A2({ S20784 }),
  .A3({ S21347 }),
  .ZN({ S21349 })
);
NAND3_X1 #() 
NAND3_X1_3812_ (
  .A1({ S21349 }),
  .A2({ S19194 }),
  .A3({ S21346 }),
  .ZN({ S21350 })
);
NAND3_X1 #() 
NAND3_X1_3813_ (
  .A1({ S20802 }),
  .A2({ S20975 }),
  .A3({ S68 }),
  .ZN({ S21351 })
);
AND3_X1 #() 
AND3_X1_138_ (
  .A1({ S21351 }),
  .A2({ S21337 }),
  .A3({ S20774 }),
  .ZN({ S21352 })
);
NAND3_X1 #() 
NAND3_X1_3814_ (
  .A1({ S20849 }),
  .A2({ S25957[1156] }),
  .A3({ S68 }),
  .ZN({ S21353 })
);
NAND2_X1 #() 
NAND2_X1_3572_ (
  .A1({ S25957[1156] }),
  .A2({ S20787 }),
  .ZN({ S21354 })
);
OAI211_X1 #() 
OAI211_X1_1240_ (
  .A({ S21353 }),
  .B({ S20784 }),
  .C1({ S20946 }),
  .C2({ S21354 }),
  .ZN({ S21355 })
);
NOR2_X1 #() 
NOR2_X1_902_ (
  .A1({ S21352 }),
  .A2({ S21355 }),
  .ZN({ S21356 })
);
NAND3_X1 #() 
NAND3_X1_3815_ (
  .A1({ S20967 }),
  .A2({ S21057 }),
  .A3({ S25957[1155] }),
  .ZN({ S21357 })
);
OAI21_X1 #() 
OAI21_X1_1840_ (
  .A({ S20774 }),
  .B1({ S21336 }),
  .B2({ S20819 }),
  .ZN({ S21358 })
);
INV_X1 #() 
INV_X1_1187_ (
  .A({ S21358 }),
  .ZN({ S21359 })
);
NAND4_X1 #() 
NAND4_X1_413_ (
  .A1({ S20776 }),
  .A2({ S25957[1156] }),
  .A3({ S20762 }),
  .A4({ S25957[1155] }),
  .ZN({ S21360 })
);
NAND3_X1 #() 
NAND3_X1_3816_ (
  .A1({ S25957[1157] }),
  .A2({ S21154 }),
  .A3({ S21360 }),
  .ZN({ S21361 })
);
AOI21_X1 #() 
AOI21_X1_1926_ (
  .A({ S21361 }),
  .B1({ S21359 }),
  .B2({ S21357 }),
  .ZN({ S21362 })
);
OAI21_X1 #() 
OAI21_X1_1841_ (
  .A({ S25957[1158] }),
  .B1({ S21356 }),
  .B2({ S21362 }),
  .ZN({ S21363 })
);
NAND3_X1 #() 
NAND3_X1_3817_ (
  .A1({ S21363 }),
  .A2({ S21350 }),
  .A3({ S19126 }),
  .ZN({ S21364 })
);
NAND3_X1 #() 
NAND3_X1_3818_ (
  .A1({ S21364 }),
  .A2({ S25957[1258] }),
  .A3({ S21341 }),
  .ZN({ S21365 })
);
AOI21_X1 #() 
AOI21_X1_1927_ (
  .A({ S25957[1157] }),
  .B1({ S21326 }),
  .B2({ S20995 }),
  .ZN({ S21366 })
);
AOI22_X1 #() 
AOI22_X1_406_ (
  .A1({ S21366 }),
  .A2({ S21325 }),
  .B1({ S21322 }),
  .B2({ S21319 }),
  .ZN({ S21367 })
);
NAND2_X1 #() 
NAND2_X1_3573_ (
  .A1({ S21334 }),
  .A2({ S21339 }),
  .ZN({ S21368 })
);
NAND2_X1 #() 
NAND2_X1_3574_ (
  .A1({ S21368 }),
  .A2({ S19194 }),
  .ZN({ S21369 })
);
OAI211_X1 #() 
OAI211_X1_1241_ (
  .A({ S21369 }),
  .B({ S25957[1159] }),
  .C1({ S21367 }),
  .C2({ S19194 }),
  .ZN({ S21370 })
);
NAND3_X1 #() 
NAND3_X1_3819_ (
  .A1({ S20830 }),
  .A2({ S21057 }),
  .A3({ S20774 }),
  .ZN({ S21371 })
);
OAI21_X1 #() 
OAI21_X1_1842_ (
  .A({ S21337 }),
  .B1({ S20771 }),
  .B2({ S21053 }),
  .ZN({ S21372 })
);
NAND2_X1 #() 
NAND2_X1_3575_ (
  .A1({ S21372 }),
  .A2({ S25957[1156] }),
  .ZN({ S21373 })
);
NAND4_X1 #() 
NAND4_X1_414_ (
  .A1({ S21373 }),
  .A2({ S21371 }),
  .A3({ S20927 }),
  .A4({ S20784 }),
  .ZN({ S21374 })
);
NAND2_X1 #() 
NAND2_X1_3576_ (
  .A1({ S21343 }),
  .A2({ S21345 }),
  .ZN({ S21375 })
);
NAND2_X1 #() 
NAND2_X1_3577_ (
  .A1({ S21375 }),
  .A2({ S25957[1157] }),
  .ZN({ S21376 })
);
NAND3_X1 #() 
NAND3_X1_3820_ (
  .A1({ S21376 }),
  .A2({ S19194 }),
  .A3({ S21374 }),
  .ZN({ S21377 })
);
NOR2_X1 #() 
NOR2_X1_903_ (
  .A1({ S20854 }),
  .A2({ S21358 }),
  .ZN({ S21378 })
);
OAI221_X1 #() 
OAI221_X1_108_ (
  .A({ S25957[1158] }),
  .B1({ S21352 }),
  .B2({ S21355 }),
  .C1({ S21378 }),
  .C2({ S21361 }),
  .ZN({ S21379 })
);
NAND3_X1 #() 
NAND3_X1_3821_ (
  .A1({ S21379 }),
  .A2({ S21377 }),
  .A3({ S19126 }),
  .ZN({ S21380 })
);
NAND3_X1 #() 
NAND3_X1_3822_ (
  .A1({ S21380 }),
  .A2({ S21370 }),
  .A3({ S21317 }),
  .ZN({ S21381 })
);
AOI21_X1 #() 
AOI21_X1_1928_ (
  .A({ S25956[42] }),
  .B1({ S21381 }),
  .B2({ S21365 }),
  .ZN({ S21382 })
);
NAND3_X1 #() 
NAND3_X1_3823_ (
  .A1({ S21364 }),
  .A2({ S21317 }),
  .A3({ S21341 }),
  .ZN({ S21383 })
);
NAND3_X1 #() 
NAND3_X1_3824_ (
  .A1({ S21380 }),
  .A2({ S21370 }),
  .A3({ S25957[1258] }),
  .ZN({ S21384 })
);
AOI21_X1 #() 
AOI21_X1_1929_ (
  .A({ S17348 }),
  .B1({ S21384 }),
  .B2({ S21383 }),
  .ZN({ S21385 })
);
OAI21_X1 #() 
OAI21_X1_1843_ (
  .A({ S25957[1162] }),
  .B1({ S21382 }),
  .B2({ S21385 }),
  .ZN({ S21386 })
);
NAND3_X1 #() 
NAND3_X1_3825_ (
  .A1({ S21384 }),
  .A2({ S21383 }),
  .A3({ S17348 }),
  .ZN({ S21387 })
);
NAND3_X1 #() 
NAND3_X1_3826_ (
  .A1({ S21381 }),
  .A2({ S21365 }),
  .A3({ S25956[42] }),
  .ZN({ S21388 })
);
NAND3_X1 #() 
NAND3_X1_3827_ (
  .A1({ S21387 }),
  .A2({ S21388 }),
  .A3({ S20138 }),
  .ZN({ S21389 })
);
NAND2_X1 #() 
NAND2_X1_3578_ (
  .A1({ S21386 }),
  .A2({ S21389 }),
  .ZN({ S25957[1034] })
);
NAND3_X1 #() 
NAND3_X1_3828_ (
  .A1({ S20021 }),
  .A2({ S25956[24] }),
  .A3({ S20022 }),
  .ZN({ S21390 })
);
NAND3_X1 #() 
NAND3_X1_3829_ (
  .A1({ S20015 }),
  .A2({ S18242 }),
  .A3({ S20019 }),
  .ZN({ S21391 })
);
OAI21_X1 #() 
OAI21_X1_1844_ (
  .A({ S18383 }),
  .B1({ S20066 }),
  .B2({ S20067 }),
  .ZN({ S21392 })
);
NAND3_X1 #() 
NAND3_X1_3830_ (
  .A1({ S20070 }),
  .A2({ S25956[25] }),
  .A3({ S20069 }),
  .ZN({ S21393 })
);
NAND4_X1 #() 
NAND4_X1_415_ (
  .A1({ S21390 }),
  .A2({ S21391 }),
  .A3({ S21392 }),
  .A4({ S21393 }),
  .ZN({ S21394 })
);
INV_X1 #() 
INV_X1_1188_ (
  .A({ S21394 }),
  .ZN({ S78 })
);
NAND4_X1 #() 
NAND4_X1_416_ (
  .A1({ S20020 }),
  .A2({ S20023 }),
  .A3({ S20068 }),
  .A4({ S20071 }),
  .ZN({ S79 })
);
INV_X1 #() 
INV_X1_1189_ (
  .A({ S19125 }),
  .ZN({ S25957[1223] })
);
INV_X1 #() 
INV_X1_1190_ (
  .A({ S25957[1183] }),
  .ZN({ S21395 })
);
OAI21_X1 #() 
OAI21_X1_1845_ (
  .A({ S18113 }),
  .B1({ S19876 }),
  .B2({ S19880 }),
  .ZN({ S21396 })
);
NAND3_X1 #() 
NAND3_X1_3831_ (
  .A1({ S19882 }),
  .A2({ S19883 }),
  .A3({ S25956[28] }),
  .ZN({ S21397 })
);
NAND2_X1 #() 
NAND2_X1_3579_ (
  .A1({ S21396 }),
  .A2({ S21397 }),
  .ZN({ S21398 })
);
NAND2_X1 #() 
NAND2_X1_3580_ (
  .A1({ S21392 }),
  .A2({ S21393 }),
  .ZN({ S21399 })
);
NAND3_X1 #() 
NAND3_X1_3832_ (
  .A1({ S21399 }),
  .A2({ S20121 }),
  .A3({ S20124 }),
  .ZN({ S21400 })
);
NAND4_X1 #() 
NAND4_X1_417_ (
  .A1({ S20020 }),
  .A2({ S20023 }),
  .A3({ S21392 }),
  .A4({ S21393 }),
  .ZN({ S21401 })
);
NAND2_X1 #() 
NAND2_X1_3581_ (
  .A1({ S21400 }),
  .A2({ S21401 }),
  .ZN({ S21402 })
);
NAND2_X1 #() 
NAND2_X1_3582_ (
  .A1({ S21402 }),
  .A2({ S25957[1179] }),
  .ZN({ S21403 })
);
NAND2_X1 #() 
NAND2_X1_3583_ (
  .A1({ S21401 }),
  .A2({ S71 }),
  .ZN({ S21404 })
);
AOI21_X1 #() 
AOI21_X1_1930_ (
  .A({ S21398 }),
  .B1({ S21403 }),
  .B2({ S21404 }),
  .ZN({ S21405 })
);
NOR2_X1 #() 
NOR2_X1_904_ (
  .A1({ S71 }),
  .A2({ S25957[1177] }),
  .ZN({ S21406 })
);
NAND2_X1 #() 
NAND2_X1_3584_ (
  .A1({ S79 }),
  .A2({ S25957[1178] }),
  .ZN({ S21407 })
);
NAND2_X1 #() 
NAND2_X1_3585_ (
  .A1({ S21390 }),
  .A2({ S21391 }),
  .ZN({ S21408 })
);
OAI21_X1 #() 
OAI21_X1_1846_ (
  .A({ S18198 }),
  .B1({ S20116 }),
  .B2({ S20120 }),
  .ZN({ S21409 })
);
NAND3_X1 #() 
NAND3_X1_3833_ (
  .A1({ S20122 }),
  .A2({ S20123 }),
  .A3({ S25956[26] }),
  .ZN({ S21410 })
);
NAND2_X1 #() 
NAND2_X1_3586_ (
  .A1({ S21409 }),
  .A2({ S21410 }),
  .ZN({ S21411 })
);
NAND3_X1 #() 
NAND3_X1_3834_ (
  .A1({ S21411 }),
  .A2({ S21408 }),
  .A3({ S21399 }),
  .ZN({ S21412 })
);
NAND2_X1 #() 
NAND2_X1_3587_ (
  .A1({ S21412 }),
  .A2({ S21407 }),
  .ZN({ S21413 })
);
AOI211_X1 #() 
AOI211_X1_57_ (
  .A({ S25957[1180] }),
  .B({ S21413 }),
  .C1({ S25957[1176] }),
  .C2({ S21406 }),
  .ZN({ S21414 })
);
OR3_X1 #() 
OR3_X1_21_ (
  .A1({ S21414 }),
  .A2({ S21405 }),
  .A3({ S25957[1181] }),
  .ZN({ S21415 })
);
NAND4_X1 #() 
NAND4_X1_418_ (
  .A1({ S21390 }),
  .A2({ S21391 }),
  .A3({ S20068 }),
  .A4({ S20071 }),
  .ZN({ S21416 })
);
INV_X1 #() 
INV_X1_1191_ (
  .A({ S21416 }),
  .ZN({ S21417 })
);
NOR2_X1 #() 
NOR2_X1_905_ (
  .A1({ S21401 }),
  .A2({ S21411 }),
  .ZN({ S21418 })
);
NOR2_X1 #() 
NOR2_X1_906_ (
  .A1({ S21418 }),
  .A2({ S21417 }),
  .ZN({ S21419 })
);
NOR2_X1 #() 
NOR2_X1_907_ (
  .A1({ S25957[1178] }),
  .A2({ S25957[1177] }),
  .ZN({ S21420 })
);
NAND2_X1 #() 
NAND2_X1_3588_ (
  .A1({ S21420 }),
  .A2({ S71 }),
  .ZN({ S21421 })
);
NAND2_X1 #() 
NAND2_X1_3589_ (
  .A1({ S21421 }),
  .A2({ S21398 }),
  .ZN({ S21422 })
);
NAND4_X1 #() 
NAND4_X1_419_ (
  .A1({ S21409 }),
  .A2({ S21410 }),
  .A3({ S21390 }),
  .A4({ S21391 }),
  .ZN({ S21423 })
);
AOI21_X1 #() 
AOI21_X1_1931_ (
  .A({ S25957[1179] }),
  .B1({ S21423 }),
  .B2({ S21401 }),
  .ZN({ S21424 })
);
AOI211_X1 #() 
AOI211_X1_58_ (
  .A({ S21424 }),
  .B({ S21422 }),
  .C1({ S21419 }),
  .C2({ S25957[1179] }),
  .ZN({ S21425 })
);
NAND3_X1 #() 
NAND3_X1_3835_ (
  .A1({ S21411 }),
  .A2({ S25957[1176] }),
  .A3({ S21399 }),
  .ZN({ S21426 })
);
AOI21_X1 #() 
AOI21_X1_1932_ (
  .A({ S71 }),
  .B1({ S25957[1178] }),
  .B2({ S21408 }),
  .ZN({ S21427 })
);
NAND4_X1 #() 
NAND4_X1_420_ (
  .A1({ S20121 }),
  .A2({ S20124 }),
  .A3({ S20020 }),
  .A4({ S20023 }),
  .ZN({ S21428 })
);
NOR2_X1 #() 
NOR2_X1_908_ (
  .A1({ S25957[1179] }),
  .A2({ S21399 }),
  .ZN({ S21429 })
);
AOI22_X1 #() 
AOI22_X1_407_ (
  .A1({ S21427 }),
  .A2({ S21426 }),
  .B1({ S21429 }),
  .B2({ S21428 }),
  .ZN({ S21430 })
);
OAI21_X1 #() 
OAI21_X1_1847_ (
  .A({ S25957[1181] }),
  .B1({ S21430 }),
  .B2({ S21398 }),
  .ZN({ S21431 })
);
OAI211_X1 #() 
OAI211_X1_1242_ (
  .A({ S21415 }),
  .B({ S25957[1182] }),
  .C1({ S21425 }),
  .C2({ S21431 }),
  .ZN({ S21432 })
);
INV_X1 #() 
INV_X1_1192_ (
  .A({ S25957[1182] }),
  .ZN({ S21433 })
);
NAND3_X1 #() 
NAND3_X1_3836_ (
  .A1({ S21394 }),
  .A2({ S79 }),
  .A3({ S25957[1178] }),
  .ZN({ S21434 })
);
NAND3_X1 #() 
NAND3_X1_3837_ (
  .A1({ S21401 }),
  .A2({ S21416 }),
  .A3({ S21411 }),
  .ZN({ S21435 })
);
AOI21_X1 #() 
AOI21_X1_1933_ (
  .A({ S71 }),
  .B1({ S21434 }),
  .B2({ S21435 }),
  .ZN({ S21436 })
);
INV_X1 #() 
INV_X1_1193_ (
  .A({ S21436 }),
  .ZN({ S21437 })
);
NAND2_X1 #() 
NAND2_X1_3590_ (
  .A1({ S25957[1178] }),
  .A2({ S25957[1177] }),
  .ZN({ S21438 })
);
NAND4_X1 #() 
NAND4_X1_421_ (
  .A1({ S20121 }),
  .A2({ S20124 }),
  .A3({ S21390 }),
  .A4({ S21391 }),
  .ZN({ S21439 })
);
NAND3_X1 #() 
NAND3_X1_3838_ (
  .A1({ S21438 }),
  .A2({ S71 }),
  .A3({ S21439 }),
  .ZN({ S21440 })
);
AOI21_X1 #() 
AOI21_X1_1934_ (
  .A({ S21398 }),
  .B1({ S21437 }),
  .B2({ S21440 }),
  .ZN({ S21441 })
);
NAND3_X1 #() 
NAND3_X1_3839_ (
  .A1({ S19808 }),
  .A2({ S19811 }),
  .A3({ S18103 }),
  .ZN({ S21442 })
);
NAND2_X1 #() 
NAND2_X1_3591_ (
  .A1({ S25957[1213] }),
  .A2({ S25956[29] }),
  .ZN({ S21443 })
);
NAND2_X1 #() 
NAND2_X1_3592_ (
  .A1({ S21443 }),
  .A2({ S21442 }),
  .ZN({ S21444 })
);
NAND2_X1 #() 
NAND2_X1_3593_ (
  .A1({ S21416 }),
  .A2({ S25957[1178] }),
  .ZN({ S21445 })
);
NAND3_X1 #() 
NAND3_X1_3840_ (
  .A1({ S21394 }),
  .A2({ S79 }),
  .A3({ S21411 }),
  .ZN({ S21446 })
);
NAND2_X1 #() 
NAND2_X1_3594_ (
  .A1({ S21446 }),
  .A2({ S21445 }),
  .ZN({ S21447 })
);
OAI21_X1 #() 
OAI21_X1_1848_ (
  .A({ S21398 }),
  .B1({ S21400 }),
  .B2({ S71 }),
  .ZN({ S21448 })
);
INV_X1 #() 
INV_X1_1194_ (
  .A({ S21448 }),
  .ZN({ S21449 })
);
OAI21_X1 #() 
OAI21_X1_1849_ (
  .A({ S21449 }),
  .B1({ S21447 }),
  .B2({ S25957[1179] }),
  .ZN({ S21450 })
);
NAND2_X1 #() 
NAND2_X1_3595_ (
  .A1({ S21450 }),
  .A2({ S21444 }),
  .ZN({ S21451 })
);
INV_X1 #() 
INV_X1_1195_ (
  .A({ S21423 }),
  .ZN({ S21452 })
);
NAND3_X1 #() 
NAND3_X1_3841_ (
  .A1({ S25957[1177] }),
  .A2({ S19959 }),
  .A3({ S19960 }),
  .ZN({ S21453 })
);
NOR2_X1 #() 
NOR2_X1_909_ (
  .A1({ S21452 }),
  .A2({ S21453 }),
  .ZN({ S21454 })
);
NAND2_X1 #() 
NAND2_X1_3596_ (
  .A1({ S25957[1179] }),
  .A2({ S21399 }),
  .ZN({ S21455 })
);
NAND2_X1 #() 
NAND2_X1_3597_ (
  .A1({ S21452 }),
  .A2({ S25957[1179] }),
  .ZN({ S21456 })
);
NAND2_X1 #() 
NAND2_X1_3598_ (
  .A1({ S21456 }),
  .A2({ S21455 }),
  .ZN({ S21457 })
);
OAI21_X1 #() 
OAI21_X1_1850_ (
  .A({ S25957[1180] }),
  .B1({ S21457 }),
  .B2({ S21454 }),
  .ZN({ S21458 })
);
NOR2_X1 #() 
NOR2_X1_910_ (
  .A1({ S71 }),
  .A2({ S25957[1176] }),
  .ZN({ S21459 })
);
INV_X1 #() 
INV_X1_1196_ (
  .A({ S21459 }),
  .ZN({ S21460 })
);
NAND4_X1 #() 
NAND4_X1_422_ (
  .A1({ S21460 }),
  .A2({ S21412 }),
  .A3({ S21398 }),
  .A4({ S21455 }),
  .ZN({ S21461 })
);
NAND3_X1 #() 
NAND3_X1_3842_ (
  .A1({ S21458 }),
  .A2({ S25957[1181] }),
  .A3({ S21461 }),
  .ZN({ S21462 })
);
OAI211_X1 #() 
OAI211_X1_1243_ (
  .A({ S21462 }),
  .B({ S21433 }),
  .C1({ S21441 }),
  .C2({ S21451 }),
  .ZN({ S21463 })
);
AOI21_X1 #() 
AOI21_X1_1935_ (
  .A({ S21395 }),
  .B1({ S21432 }),
  .B2({ S21463 }),
  .ZN({ S21464 })
);
NAND3_X1 #() 
NAND3_X1_3843_ (
  .A1({ S21411 }),
  .A2({ S25957[1176] }),
  .A3({ S25957[1177] }),
  .ZN({ S21465 })
);
OAI21_X1 #() 
OAI21_X1_1851_ (
  .A({ S25957[1179] }),
  .B1({ S79 }),
  .B2({ S21411 }),
  .ZN({ S21466 })
);
INV_X1 #() 
INV_X1_1197_ (
  .A({ S21466 }),
  .ZN({ S21467 })
);
OAI21_X1 #() 
OAI21_X1_1852_ (
  .A({ S21408 }),
  .B1({ S21411 }),
  .B2({ S25957[1177] }),
  .ZN({ S21468 })
);
AOI21_X1 #() 
AOI21_X1_1936_ (
  .A({ S21398 }),
  .B1({ S21468 }),
  .B2({ S71 }),
  .ZN({ S21469 })
);
INV_X1 #() 
INV_X1_1198_ (
  .A({ S21469 }),
  .ZN({ S21470 })
);
AOI21_X1 #() 
AOI21_X1_1937_ (
  .A({ S21470 }),
  .B1({ S21467 }),
  .B2({ S21465 }),
  .ZN({ S21471 })
);
NAND2_X1 #() 
NAND2_X1_3599_ (
  .A1({ S25957[1178] }),
  .A2({ S21399 }),
  .ZN({ S21472 })
);
NAND2_X1 #() 
NAND2_X1_3600_ (
  .A1({ S21416 }),
  .A2({ S21411 }),
  .ZN({ S21473 })
);
NAND3_X1 #() 
NAND3_X1_3844_ (
  .A1({ S21473 }),
  .A2({ S25957[1179] }),
  .A3({ S21472 }),
  .ZN({ S21474 })
);
INV_X1 #() 
INV_X1_1199_ (
  .A({ S21474 }),
  .ZN({ S21475 })
);
AOI21_X1 #() 
AOI21_X1_1938_ (
  .A({ S25957[1179] }),
  .B1({ S21394 }),
  .B2({ S25957[1178] }),
  .ZN({ S21476 })
);
NOR3_X1 #() 
NOR3_X1_123_ (
  .A1({ S21475 }),
  .A2({ S21476 }),
  .A3({ S25957[1180] }),
  .ZN({ S21477 })
);
OR3_X1 #() 
OR3_X1_22_ (
  .A1({ S21471 }),
  .A2({ S21477 }),
  .A3({ S21444 }),
  .ZN({ S21478 })
);
OAI211_X1 #() 
OAI211_X1_1244_ (
  .A({ S21423 }),
  .B({ S25957[1179] }),
  .C1({ S21399 }),
  .C2({ S25957[1178] }),
  .ZN({ S21479 })
);
NAND2_X1 #() 
NAND2_X1_3601_ (
  .A1({ S21394 }),
  .A2({ S25957[1178] }),
  .ZN({ S21480 })
);
NAND2_X1 #() 
NAND2_X1_3602_ (
  .A1({ S21480 }),
  .A2({ S21473 }),
  .ZN({ S21481 })
);
AOI21_X1 #() 
AOI21_X1_1939_ (
  .A({ S25957[1180] }),
  .B1({ S21481 }),
  .B2({ S71 }),
  .ZN({ S21482 })
);
NAND3_X1 #() 
NAND3_X1_3845_ (
  .A1({ S21401 }),
  .A2({ S21416 }),
  .A3({ S25957[1178] }),
  .ZN({ S21483 })
);
AOI21_X1 #() 
AOI21_X1_1940_ (
  .A({ S25957[1179] }),
  .B1({ S21483 }),
  .B2({ S21428 }),
  .ZN({ S21484 })
);
AOI21_X1 #() 
AOI21_X1_1941_ (
  .A({ S71 }),
  .B1({ S21435 }),
  .B2({ S21480 }),
  .ZN({ S21485 })
);
NOR3_X1 #() 
NOR3_X1_124_ (
  .A1({ S21485 }),
  .A2({ S21484 }),
  .A3({ S21398 }),
  .ZN({ S21486 })
);
AOI21_X1 #() 
AOI21_X1_1942_ (
  .A({ S21486 }),
  .B1({ S21482 }),
  .B2({ S21479 }),
  .ZN({ S21487 })
);
OAI211_X1 #() 
OAI211_X1_1245_ (
  .A({ S21478 }),
  .B({ S25957[1182] }),
  .C1({ S25957[1181] }),
  .C2({ S21487 }),
  .ZN({ S21488 })
);
AOI21_X1 #() 
AOI21_X1_1943_ (
  .A({ S25957[1179] }),
  .B1({ S25957[1178] }),
  .B2({ S25957[1177] }),
  .ZN({ S21489 })
);
NAND2_X1 #() 
NAND2_X1_3603_ (
  .A1({ S21394 }),
  .A2({ S21411 }),
  .ZN({ S21490 })
);
AOI21_X1 #() 
AOI21_X1_1944_ (
  .A({ S71 }),
  .B1({ S21438 }),
  .B2({ S79 }),
  .ZN({ S21491 })
);
AOI21_X1 #() 
AOI21_X1_1945_ (
  .A({ S21491 }),
  .B1({ S21490 }),
  .B2({ S21489 }),
  .ZN({ S21492 })
);
NAND4_X1 #() 
NAND4_X1_423_ (
  .A1({ S19959 }),
  .A2({ S21390 }),
  .A3({ S21391 }),
  .A4({ S19960 }),
  .ZN({ S21493 })
);
NAND2_X1 #() 
NAND2_X1_3604_ (
  .A1({ S21423 }),
  .A2({ S25957[1179] }),
  .ZN({ S21494 })
);
OAI21_X1 #() 
OAI21_X1_1853_ (
  .A({ S21493 }),
  .B1({ S21494 }),
  .B2({ S21420 }),
  .ZN({ S21495 })
);
OR2_X1 #() 
OR2_X1_48_ (
  .A1({ S21495 }),
  .A2({ S21398 }),
  .ZN({ S21496 })
);
OAI211_X1 #() 
OAI211_X1_1246_ (
  .A({ S21496 }),
  .B({ S25957[1181] }),
  .C1({ S25957[1180] }),
  .C2({ S21492 }),
  .ZN({ S21497 })
);
NAND3_X1 #() 
NAND3_X1_3846_ (
  .A1({ S21434 }),
  .A2({ S71 }),
  .A3({ S21465 }),
  .ZN({ S21498 })
);
OAI21_X1 #() 
OAI21_X1_1854_ (
  .A({ S21498 }),
  .B1({ S71 }),
  .B2({ S21418 }),
  .ZN({ S21499 })
);
NOR2_X1 #() 
NOR2_X1_911_ (
  .A1({ S21404 }),
  .A2({ S21445 }),
  .ZN({ S21500 })
);
OAI21_X1 #() 
OAI21_X1_1855_ (
  .A({ S21398 }),
  .B1({ S21480 }),
  .B2({ S71 }),
  .ZN({ S21501 })
);
OAI22_X1 #() 
OAI22_X1_98_ (
  .A1({ S21499 }),
  .A2({ S21398 }),
  .B1({ S21500 }),
  .B2({ S21501 }),
  .ZN({ S21502 })
);
OAI211_X1 #() 
OAI211_X1_1247_ (
  .A({ S21497 }),
  .B({ S21433 }),
  .C1({ S25957[1181] }),
  .C2({ S21502 }),
  .ZN({ S21503 })
);
AOI21_X1 #() 
AOI21_X1_1946_ (
  .A({ S25957[1183] }),
  .B1({ S21488 }),
  .B2({ S21503 }),
  .ZN({ S21504 })
);
NOR2_X1 #() 
NOR2_X1_912_ (
  .A1({ S21504 }),
  .A2({ S21464 }),
  .ZN({ S21505 })
);
NAND2_X1 #() 
NAND2_X1_3605_ (
  .A1({ S21505 }),
  .A2({ S19124 }),
  .ZN({ S21506 })
);
INV_X1 #() 
INV_X1_1200_ (
  .A({ S19124 }),
  .ZN({ S25957[1255] })
);
OAI21_X1 #() 
OAI21_X1_1856_ (
  .A({ S25957[1255] }),
  .B1({ S21504 }),
  .B2({ S21464 }),
  .ZN({ S21507 })
);
NAND3_X1 #() 
NAND3_X1_3847_ (
  .A1({ S21506 }),
  .A2({ S25957[1223] }),
  .A3({ S21507 }),
  .ZN({ S21508 })
);
NAND2_X1 #() 
NAND2_X1_3606_ (
  .A1({ S21506 }),
  .A2({ S21507 }),
  .ZN({ S25957[1127] })
);
NAND2_X1 #() 
NAND2_X1_3607_ (
  .A1({ S25957[1127] }),
  .A2({ S19125 }),
  .ZN({ S21509 })
);
NAND2_X1 #() 
NAND2_X1_3608_ (
  .A1({ S21509 }),
  .A2({ S21508 }),
  .ZN({ S25957[1095] })
);
NAND2_X1 #() 
NAND2_X1_3609_ (
  .A1({ S25957[1095] }),
  .A2({ S25956[7] }),
  .ZN({ S21510 })
);
NAND3_X1 #() 
NAND3_X1_3848_ (
  .A1({ S21509 }),
  .A2({ S11609 }),
  .A3({ S21508 }),
  .ZN({ S21511 })
);
NAND2_X1 #() 
NAND2_X1_3610_ (
  .A1({ S21510 }),
  .A2({ S21511 }),
  .ZN({ S21512 })
);
INV_X1 #() 
INV_X1_1201_ (
  .A({ S21512 }),
  .ZN({ S25957[1031] })
);
INV_X1 #() 
INV_X1_1202_ (
  .A({ S25957[1222] }),
  .ZN({ S21513 })
);
INV_X1 #() 
INV_X1_1203_ (
  .A({ S25957[1254] }),
  .ZN({ S21514 })
);
AOI21_X1 #() 
AOI21_X1_1947_ (
  .A({ S25957[1179] }),
  .B1({ S21446 }),
  .B2({ S21423 }),
  .ZN({ S21515 })
);
AOI21_X1 #() 
AOI21_X1_1948_ (
  .A({ S71 }),
  .B1({ S21445 }),
  .B2({ S21439 }),
  .ZN({ S21516 })
);
NOR3_X1 #() 
NOR3_X1_125_ (
  .A1({ S21515 }),
  .A2({ S21516 }),
  .A3({ S21398 }),
  .ZN({ S21517 })
);
INV_X1 #() 
INV_X1_1204_ (
  .A({ S21482 }),
  .ZN({ S21518 })
);
AOI21_X1 #() 
AOI21_X1_1949_ (
  .A({ S71 }),
  .B1({ S21465 }),
  .B2({ S21407 }),
  .ZN({ S21519 })
);
NOR2_X1 #() 
NOR2_X1_913_ (
  .A1({ S21518 }),
  .A2({ S21519 }),
  .ZN({ S21520 })
);
OAI21_X1 #() 
OAI21_X1_1857_ (
  .A({ S25957[1182] }),
  .B1({ S21520 }),
  .B2({ S21517 }),
  .ZN({ S21521 })
);
NAND3_X1 #() 
NAND3_X1_3849_ (
  .A1({ S25957[1178] }),
  .A2({ S21408 }),
  .A3({ S25957[1177] }),
  .ZN({ S21522 })
);
AOI21_X1 #() 
AOI21_X1_1950_ (
  .A({ S71 }),
  .B1({ S21522 }),
  .B2({ S21439 }),
  .ZN({ S21523 })
);
OAI21_X1 #() 
OAI21_X1_1858_ (
  .A({ S21398 }),
  .B1({ S21515 }),
  .B2({ S21523 }),
  .ZN({ S21524 })
);
NOR2_X1 #() 
NOR2_X1_914_ (
  .A1({ S21473 }),
  .A2({ S25957[1179] }),
  .ZN({ S21525 })
);
OAI211_X1 #() 
OAI211_X1_1248_ (
  .A({ S21455 }),
  .B({ S25957[1180] }),
  .C1({ S71 }),
  .C2({ S21423 }),
  .ZN({ S21526 })
);
OAI211_X1 #() 
OAI211_X1_1249_ (
  .A({ S21524 }),
  .B({ S21433 }),
  .C1({ S21525 }),
  .C2({ S21526 }),
  .ZN({ S21527 })
);
AOI21_X1 #() 
AOI21_X1_1951_ (
  .A({ S25957[1181] }),
  .B1({ S21521 }),
  .B2({ S21527 }),
  .ZN({ S21528 })
);
NAND2_X1 #() 
NAND2_X1_3611_ (
  .A1({ S79 }),
  .A2({ S21411 }),
  .ZN({ S21529 })
);
NAND2_X1 #() 
NAND2_X1_3612_ (
  .A1({ S21434 }),
  .A2({ S21529 }),
  .ZN({ S21530 })
);
NAND2_X1 #() 
NAND2_X1_3613_ (
  .A1({ S21401 }),
  .A2({ S21411 }),
  .ZN({ S21531 })
);
NAND2_X1 #() 
NAND2_X1_3614_ (
  .A1({ S21531 }),
  .A2({ S21438 }),
  .ZN({ S21532 })
);
NAND2_X1 #() 
NAND2_X1_3615_ (
  .A1({ S21532 }),
  .A2({ S25957[1179] }),
  .ZN({ S21533 })
);
OAI211_X1 #() 
OAI211_X1_1250_ (
  .A({ S21533 }),
  .B({ S21398 }),
  .C1({ S25957[1179] }),
  .C2({ S21530 }),
  .ZN({ S21534 })
);
NAND4_X1 #() 
NAND4_X1_424_ (
  .A1({ S19959 }),
  .A2({ S20121 }),
  .A3({ S19960 }),
  .A4({ S20124 }),
  .ZN({ S21535 })
);
OAI22_X1 #() 
OAI22_X1_99_ (
  .A1({ S21438 }),
  .A2({ S71 }),
  .B1({ S21535 }),
  .B2({ S21401 }),
  .ZN({ S21536 })
);
OAI21_X1 #() 
OAI21_X1_1859_ (
  .A({ S25957[1180] }),
  .B1({ S21500 }),
  .B2({ S21536 }),
  .ZN({ S21537 })
);
NAND3_X1 #() 
NAND3_X1_3850_ (
  .A1({ S21534 }),
  .A2({ S21433 }),
  .A3({ S21537 }),
  .ZN({ S21538 })
);
AOI21_X1 #() 
AOI21_X1_1952_ (
  .A({ S21429 }),
  .B1({ S21402 }),
  .B2({ S25957[1179] }),
  .ZN({ S21539 })
);
NAND4_X1 #() 
NAND4_X1_425_ (
  .A1({ S21409 }),
  .A2({ S21410 }),
  .A3({ S20020 }),
  .A4({ S20023 }),
  .ZN({ S21540 })
);
NAND3_X1 #() 
NAND3_X1_3851_ (
  .A1({ S21406 }),
  .A2({ S21540 }),
  .A3({ S21439 }),
  .ZN({ S21541 })
);
OAI211_X1 #() 
OAI211_X1_1251_ (
  .A({ S21541 }),
  .B({ S25957[1180] }),
  .C1({ S25957[1179] }),
  .C2({ S21407 }),
  .ZN({ S21542 })
);
OAI211_X1 #() 
OAI211_X1_1252_ (
  .A({ S25957[1182] }),
  .B({ S21542 }),
  .C1({ S21539 }),
  .C2({ S25957[1180] }),
  .ZN({ S21543 })
);
AOI21_X1 #() 
AOI21_X1_1953_ (
  .A({ S21444 }),
  .B1({ S21538 }),
  .B2({ S21543 }),
  .ZN({ S21544 })
);
OR3_X1 #() 
OR3_X1_23_ (
  .A1({ S21528 }),
  .A2({ S21544 }),
  .A3({ S21395 }),
  .ZN({ S21545 })
);
NAND3_X1 #() 
NAND3_X1_3852_ (
  .A1({ S21400 }),
  .A2({ S71 }),
  .A3({ S21408 }),
  .ZN({ S21546 })
);
NOR2_X1 #() 
NOR2_X1_915_ (
  .A1({ S25957[1178] }),
  .A2({ S21399 }),
  .ZN({ S21547 })
);
AOI21_X1 #() 
AOI21_X1_1954_ (
  .A({ S21398 }),
  .B1({ S21547 }),
  .B2({ S25957[1179] }),
  .ZN({ S21548 })
);
AOI21_X1 #() 
AOI21_X1_1955_ (
  .A({ S21516 }),
  .B1({ S21434 }),
  .B2({ S71 }),
  .ZN({ S21549 })
);
AOI22_X1 #() 
AOI22_X1_408_ (
  .A1({ S21549 }),
  .A2({ S21398 }),
  .B1({ S21546 }),
  .B2({ S21548 }),
  .ZN({ S21550 })
);
NOR2_X1 #() 
NOR2_X1_916_ (
  .A1({ S21550 }),
  .A2({ S21433 }),
  .ZN({ S21551 })
);
AOI21_X1 #() 
AOI21_X1_1956_ (
  .A({ S21398 }),
  .B1({ S21426 }),
  .B2({ S71 }),
  .ZN({ S21552 })
);
NAND2_X1 #() 
NAND2_X1_3616_ (
  .A1({ S21522 }),
  .A2({ S21531 }),
  .ZN({ S21553 })
);
NAND2_X1 #() 
NAND2_X1_3617_ (
  .A1({ S21553 }),
  .A2({ S25957[1179] }),
  .ZN({ S21554 })
);
NOR2_X1 #() 
NOR2_X1_917_ (
  .A1({ S21554 }),
  .A2({ S25957[1180] }),
  .ZN({ S21555 })
);
AOI211_X1 #() 
AOI211_X1_59_ (
  .A({ S25957[1182] }),
  .B({ S21555 }),
  .C1({ S21474 }),
  .C2({ S21552 }),
  .ZN({ S21556 })
);
OAI21_X1 #() 
OAI21_X1_1860_ (
  .A({ S21444 }),
  .B1({ S21556 }),
  .B2({ S21551 }),
  .ZN({ S21557 })
);
NAND2_X1 #() 
NAND2_X1_3618_ (
  .A1({ S21489 }),
  .A2({ S21426 }),
  .ZN({ S21558 })
);
NAND2_X1 #() 
NAND2_X1_3619_ (
  .A1({ S21472 }),
  .A2({ S25957[1179] }),
  .ZN({ S21559 })
);
OR2_X1 #() 
OR2_X1_49_ (
  .A1({ S21559 }),
  .A2({ S21547 }),
  .ZN({ S21560 })
);
AOI21_X1 #() 
AOI21_X1_1957_ (
  .A({ S25957[1180] }),
  .B1({ S21560 }),
  .B2({ S21558 }),
  .ZN({ S21561 })
);
NAND2_X1 #() 
NAND2_X1_3620_ (
  .A1({ S21439 }),
  .A2({ S71 }),
  .ZN({ S21562 })
);
NAND2_X1 #() 
NAND2_X1_3621_ (
  .A1({ S21467 }),
  .A2({ S21394 }),
  .ZN({ S21563 })
);
AOI21_X1 #() 
AOI21_X1_1958_ (
  .A({ S21398 }),
  .B1({ S21563 }),
  .B2({ S21562 }),
  .ZN({ S21564 })
);
NOR3_X1 #() 
NOR3_X1_126_ (
  .A1({ S21561 }),
  .A2({ S21564 }),
  .A3({ S25957[1182] }),
  .ZN({ S21565 })
);
NAND3_X1 #() 
NAND3_X1_3853_ (
  .A1({ S21480 }),
  .A2({ S71 }),
  .A3({ S21439 }),
  .ZN({ S21566 })
);
NAND2_X1 #() 
NAND2_X1_3622_ (
  .A1({ S21423 }),
  .A2({ S21401 }),
  .ZN({ S21567 })
);
AOI21_X1 #() 
AOI21_X1_1959_ (
  .A({ S21398 }),
  .B1({ S21567 }),
  .B2({ S25957[1179] }),
  .ZN({ S21568 })
);
NAND2_X1 #() 
NAND2_X1_3623_ (
  .A1({ S21439 }),
  .A2({ S25957[1177] }),
  .ZN({ S21569 })
);
AOI21_X1 #() 
AOI21_X1_1960_ (
  .A({ S25957[1180] }),
  .B1({ S21456 }),
  .B2({ S21569 }),
  .ZN({ S21570 })
);
AOI211_X1 #() 
AOI211_X1_60_ (
  .A({ S21570 }),
  .B({ S21433 }),
  .C1({ S21568 }),
  .C2({ S21566 }),
  .ZN({ S21571 })
);
OAI21_X1 #() 
OAI21_X1_1861_ (
  .A({ S25957[1181] }),
  .B1({ S21571 }),
  .B2({ S21565 }),
  .ZN({ S21572 })
);
NAND3_X1 #() 
NAND3_X1_3854_ (
  .A1({ S21557 }),
  .A2({ S21572 }),
  .A3({ S21395 }),
  .ZN({ S21573 })
);
NAND3_X1 #() 
NAND3_X1_3855_ (
  .A1({ S21545 }),
  .A2({ S21514 }),
  .A3({ S21573 }),
  .ZN({ S21574 })
);
NAND2_X1 #() 
NAND2_X1_3624_ (
  .A1({ S21545 }),
  .A2({ S21573 }),
  .ZN({ S21575 })
);
NAND2_X1 #() 
NAND2_X1_3625_ (
  .A1({ S21575 }),
  .A2({ S25957[1254] }),
  .ZN({ S21576 })
);
NAND2_X1 #() 
NAND2_X1_3626_ (
  .A1({ S21576 }),
  .A2({ S21574 }),
  .ZN({ S25957[1126] })
);
NAND2_X1 #() 
NAND2_X1_3627_ (
  .A1({ S25957[1126] }),
  .A2({ S21513 }),
  .ZN({ S21577 })
);
NAND3_X1 #() 
NAND3_X1_3856_ (
  .A1({ S21576 }),
  .A2({ S21574 }),
  .A3({ S25957[1222] }),
  .ZN({ S21578 })
);
NAND2_X1 #() 
NAND2_X1_3628_ (
  .A1({ S21577 }),
  .A2({ S21578 }),
  .ZN({ S25957[1094] })
);
NAND2_X1 #() 
NAND2_X1_3629_ (
  .A1({ S25957[1094] }),
  .A2({ S25956[6] }),
  .ZN({ S21579 })
);
NAND3_X1 #() 
NAND3_X1_3857_ (
  .A1({ S21577 }),
  .A2({ S21578 }),
  .A3({ S11620 }),
  .ZN({ S21580 })
);
NAND2_X1 #() 
NAND2_X1_3630_ (
  .A1({ S21579 }),
  .A2({ S21580 }),
  .ZN({ S21581 })
);
INV_X1 #() 
INV_X1_1205_ (
  .A({ S21581 }),
  .ZN({ S25957[1030] })
);
INV_X1 #() 
INV_X1_1206_ (
  .A({ S25957[1253] }),
  .ZN({ S21582 })
);
NAND3_X1 #() 
NAND3_X1_3858_ (
  .A1({ S21428 }),
  .A2({ S71 }),
  .A3({ S21394 }),
  .ZN({ S21583 })
);
OAI21_X1 #() 
OAI21_X1_1862_ (
  .A({ S21583 }),
  .B1({ S21481 }),
  .B2({ S71 }),
  .ZN({ S21584 })
);
AOI21_X1 #() 
AOI21_X1_1961_ (
  .A({ S25957[1179] }),
  .B1({ S21408 }),
  .B2({ S25957[1177] }),
  .ZN({ S21585 })
);
NAND2_X1 #() 
NAND2_X1_3631_ (
  .A1({ S21585 }),
  .A2({ S21400 }),
  .ZN({ S21586 })
);
NOR2_X1 #() 
NOR2_X1_918_ (
  .A1({ S21406 }),
  .A2({ S25957[1180] }),
  .ZN({ S21587 })
);
AOI21_X1 #() 
AOI21_X1_1962_ (
  .A({ S21444 }),
  .B1({ S21586 }),
  .B2({ S21587 }),
  .ZN({ S21588 })
);
OAI21_X1 #() 
OAI21_X1_1863_ (
  .A({ S21588 }),
  .B1({ S21584 }),
  .B2({ S21398 }),
  .ZN({ S21589 })
);
AOI21_X1 #() 
AOI21_X1_1963_ (
  .A({ S71 }),
  .B1({ S21434 }),
  .B2({ S21412 }),
  .ZN({ S21590 })
);
AOI211_X1 #() 
AOI211_X1_61_ (
  .A({ S25957[1180] }),
  .B({ S21590 }),
  .C1({ S71 }),
  .C2({ S21465 }),
  .ZN({ S21591 })
);
AOI21_X1 #() 
AOI21_X1_1964_ (
  .A({ S25957[1178] }),
  .B1({ S21401 }),
  .B2({ S21416 }),
  .ZN({ S21592 })
);
NAND2_X1 #() 
NAND2_X1_3632_ (
  .A1({ S21592 }),
  .A2({ S25957[1179] }),
  .ZN({ S21593 })
);
NAND3_X1 #() 
NAND3_X1_3859_ (
  .A1({ S21439 }),
  .A2({ S71 }),
  .A3({ S21399 }),
  .ZN({ S21594 })
);
AOI21_X1 #() 
AOI21_X1_1965_ (
  .A({ S21398 }),
  .B1({ S21593 }),
  .B2({ S21594 }),
  .ZN({ S21595 })
);
OR2_X1 #() 
OR2_X1_50_ (
  .A1({ S21595 }),
  .A2({ S25957[1181] }),
  .ZN({ S21596 })
);
OAI211_X1 #() 
OAI211_X1_1253_ (
  .A({ S21433 }),
  .B({ S21589 }),
  .C1({ S21596 }),
  .C2({ S21591 }),
  .ZN({ S21597 })
);
NAND2_X1 #() 
NAND2_X1_3633_ (
  .A1({ S21585 }),
  .A2({ S21473 }),
  .ZN({ S21598 })
);
AOI21_X1 #() 
AOI21_X1_1966_ (
  .A({ S21398 }),
  .B1({ S21459 }),
  .B2({ S21400 }),
  .ZN({ S21599 })
);
NAND2_X1 #() 
NAND2_X1_3634_ (
  .A1({ S21423 }),
  .A2({ S21399 }),
  .ZN({ S21600 })
);
NAND2_X1 #() 
NAND2_X1_3635_ (
  .A1({ S21600 }),
  .A2({ S71 }),
  .ZN({ S21601 })
);
AOI22_X1 #() 
AOI22_X1_409_ (
  .A1({ S21409 }),
  .A2({ S21410 }),
  .B1({ S21391 }),
  .B2({ S21390 }),
  .ZN({ S21602 })
);
OAI21_X1 #() 
OAI21_X1_1864_ (
  .A({ S25957[1179] }),
  .B1({ S21602 }),
  .B2({ S21399 }),
  .ZN({ S21603 })
);
NAND3_X1 #() 
NAND3_X1_3860_ (
  .A1({ S21601 }),
  .A2({ S21456 }),
  .A3({ S21603 }),
  .ZN({ S21604 })
);
AOI22_X1 #() 
AOI22_X1_410_ (
  .A1({ S21604 }),
  .A2({ S21398 }),
  .B1({ S21598 }),
  .B2({ S21599 }),
  .ZN({ S21605 })
);
INV_X1 #() 
INV_X1_1207_ (
  .A({ S21516 }),
  .ZN({ S21606 })
);
NAND3_X1 #() 
NAND3_X1_3861_ (
  .A1({ S21606 }),
  .A2({ S21398 }),
  .A3({ S21483 }),
  .ZN({ S21607 })
);
NAND2_X1 #() 
NAND2_X1_3636_ (
  .A1({ S21585 }),
  .A2({ S25957[1178] }),
  .ZN({ S21608 })
);
NAND2_X1 #() 
NAND2_X1_3637_ (
  .A1({ S21531 }),
  .A2({ S25957[1179] }),
  .ZN({ S21609 })
);
NAND3_X1 #() 
NAND3_X1_3862_ (
  .A1({ S21608 }),
  .A2({ S25957[1180] }),
  .A3({ S21609 }),
  .ZN({ S21610 })
);
NAND3_X1 #() 
NAND3_X1_3863_ (
  .A1({ S21607 }),
  .A2({ S21444 }),
  .A3({ S21610 }),
  .ZN({ S21611 })
);
OAI211_X1 #() 
OAI211_X1_1254_ (
  .A({ S21611 }),
  .B({ S25957[1182] }),
  .C1({ S21444 }),
  .C2({ S21605 }),
  .ZN({ S21612 })
);
NAND3_X1 #() 
NAND3_X1_3864_ (
  .A1({ S21597 }),
  .A2({ S25957[1183] }),
  .A3({ S21612 }),
  .ZN({ S21613 })
);
NAND3_X1 #() 
NAND3_X1_3865_ (
  .A1({ S21473 }),
  .A2({ S71 }),
  .A3({ S21472 }),
  .ZN({ S21614 })
);
NOR2_X1 #() 
NOR2_X1_919_ (
  .A1({ S21401 }),
  .A2({ S25957[1178] }),
  .ZN({ S21615 })
);
INV_X1 #() 
INV_X1_1208_ (
  .A({ S21615 }),
  .ZN({ S21616 })
);
NAND3_X1 #() 
NAND3_X1_3866_ (
  .A1({ S21616 }),
  .A2({ S25957[1179] }),
  .A3({ S21483 }),
  .ZN({ S21617 })
);
AOI21_X1 #() 
AOI21_X1_1967_ (
  .A({ S21398 }),
  .B1({ S21617 }),
  .B2({ S21614 }),
  .ZN({ S21618 })
);
OAI21_X1 #() 
OAI21_X1_1865_ (
  .A({ S71 }),
  .B1({ S21401 }),
  .B2({ S25957[1178] }),
  .ZN({ S21619 })
);
NAND3_X1 #() 
NAND3_X1_3867_ (
  .A1({ S21480 }),
  .A2({ S25957[1179] }),
  .A3({ S21439 }),
  .ZN({ S21620 })
);
OAI21_X1 #() 
OAI21_X1_1866_ (
  .A({ S21620 }),
  .B1({ S21452 }),
  .B2({ S21619 }),
  .ZN({ S21621 })
);
NAND3_X1 #() 
NAND3_X1_3868_ (
  .A1({ S25957[1178] }),
  .A2({ S25957[1176] }),
  .A3({ S25957[1177] }),
  .ZN({ S21622 })
);
NAND3_X1 #() 
NAND3_X1_3869_ (
  .A1({ S21622 }),
  .A2({ S21490 }),
  .A3({ S71 }),
  .ZN({ S21623 })
);
NAND3_X1 #() 
NAND3_X1_3870_ (
  .A1({ S21416 }),
  .A2({ S25957[1179] }),
  .A3({ S21411 }),
  .ZN({ S21624 })
);
AND2_X1 #() 
AND2_X1_224_ (
  .A1({ S21624 }),
  .A2({ S25957[1180] }),
  .ZN({ S21625 })
);
AOI22_X1 #() 
AOI22_X1_411_ (
  .A1({ S21621 }),
  .A2({ S21398 }),
  .B1({ S21625 }),
  .B2({ S21623 }),
  .ZN({ S21626 })
);
NAND2_X1 #() 
NAND2_X1_3638_ (
  .A1({ S21585 }),
  .A2({ S21439 }),
  .ZN({ S21627 })
);
NAND3_X1 #() 
NAND3_X1_3871_ (
  .A1({ S21627 }),
  .A2({ S21398 }),
  .A3({ S21460 }),
  .ZN({ S21628 })
);
NAND2_X1 #() 
NAND2_X1_3639_ (
  .A1({ S21628 }),
  .A2({ S25957[1181] }),
  .ZN({ S21629 })
);
OAI22_X1 #() 
OAI22_X1_100_ (
  .A1({ S21626 }),
  .A2({ S25957[1181] }),
  .B1({ S21629 }),
  .B2({ S21618 }),
  .ZN({ S21630 })
);
NOR2_X1 #() 
NOR2_X1_920_ (
  .A1({ S21394 }),
  .A2({ S25957[1179] }),
  .ZN({ S21631 })
);
AOI22_X1 #() 
AOI22_X1_412_ (
  .A1({ S21631 }),
  .A2({ S25957[1178] }),
  .B1({ S21417 }),
  .B2({ S25957[1179] }),
  .ZN({ S21632 })
);
INV_X1 #() 
INV_X1_1209_ (
  .A({ S21426 }),
  .ZN({ S21633 })
);
NAND2_X1 #() 
NAND2_X1_3640_ (
  .A1({ S21483 }),
  .A2({ S25957[1179] }),
  .ZN({ S21634 })
);
NAND4_X1 #() 
NAND4_X1_426_ (
  .A1({ S21428 }),
  .A2({ S21416 }),
  .A3({ S21401 }),
  .A4({ S71 }),
  .ZN({ S21635 })
);
OAI211_X1 #() 
OAI211_X1_1255_ (
  .A({ S25957[1180] }),
  .B({ S21635 }),
  .C1({ S21634 }),
  .C2({ S21633 }),
  .ZN({ S21636 })
);
OAI211_X1 #() 
OAI211_X1_1256_ (
  .A({ S21636 }),
  .B({ S21444 }),
  .C1({ S25957[1180] }),
  .C2({ S21632 }),
  .ZN({ S21637 })
);
OAI21_X1 #() 
OAI21_X1_1867_ (
  .A({ S21619 }),
  .B1({ S71 }),
  .B2({ S21490 }),
  .ZN({ S21638 })
);
INV_X1 #() 
INV_X1_1210_ (
  .A({ S21540 }),
  .ZN({ S21639 })
);
OAI21_X1 #() 
OAI21_X1_1868_ (
  .A({ S71 }),
  .B1({ S21569 }),
  .B2({ S21639 }),
  .ZN({ S21640 })
);
AOI21_X1 #() 
AOI21_X1_1968_ (
  .A({ S25957[1180] }),
  .B1({ S25957[1179] }),
  .B2({ S21423 }),
  .ZN({ S21641 })
);
AOI22_X1 #() 
AOI22_X1_413_ (
  .A1({ S21638 }),
  .A2({ S25957[1180] }),
  .B1({ S21640 }),
  .B2({ S21641 }),
  .ZN({ S21642 })
);
AOI21_X1 #() 
AOI21_X1_1969_ (
  .A({ S25957[1182] }),
  .B1({ S21642 }),
  .B2({ S25957[1181] }),
  .ZN({ S21643 })
);
AOI22_X1 #() 
AOI22_X1_414_ (
  .A1({ S21630 }),
  .A2({ S25957[1182] }),
  .B1({ S21637 }),
  .B2({ S21643 }),
  .ZN({ S21644 })
);
OAI21_X1 #() 
OAI21_X1_1869_ (
  .A({ S21613 }),
  .B1({ S21644 }),
  .B2({ S25957[1183] }),
  .ZN({ S21645 })
);
NAND2_X1 #() 
NAND2_X1_3641_ (
  .A1({ S21645 }),
  .A2({ S21582 }),
  .ZN({ S21646 })
);
OAI211_X1 #() 
OAI211_X1_1257_ (
  .A({ S21613 }),
  .B({ S25957[1253] }),
  .C1({ S21644 }),
  .C2({ S25957[1183] }),
  .ZN({ S21647 })
);
AOI21_X1 #() 
AOI21_X1_1970_ (
  .A({ S25957[1221] }),
  .B1({ S21646 }),
  .B2({ S21647 }),
  .ZN({ S21648 })
);
INV_X1 #() 
INV_X1_1211_ (
  .A({ S25957[1221] }),
  .ZN({ S21649 })
);
OAI211_X1 #() 
OAI211_X1_1258_ (
  .A({ S21613 }),
  .B({ S21582 }),
  .C1({ S21644 }),
  .C2({ S25957[1183] }),
  .ZN({ S21650 })
);
NAND2_X1 #() 
NAND2_X1_3642_ (
  .A1({ S21645 }),
  .A2({ S25957[1253] }),
  .ZN({ S21651 })
);
AOI21_X1 #() 
AOI21_X1_1971_ (
  .A({ S21649 }),
  .B1({ S21651 }),
  .B2({ S21650 }),
  .ZN({ S21652 })
);
OAI21_X1 #() 
OAI21_X1_1870_ (
  .A({ S25956[5] }),
  .B1({ S21648 }),
  .B2({ S21652 }),
  .ZN({ S21653 })
);
NAND3_X1 #() 
NAND3_X1_3872_ (
  .A1({ S21651 }),
  .A2({ S21649 }),
  .A3({ S21650 }),
  .ZN({ S21654 })
);
NAND2_X1 #() 
NAND2_X1_3643_ (
  .A1({ S21651 }),
  .A2({ S21650 }),
  .ZN({ S25957[1125] })
);
NAND2_X1 #() 
NAND2_X1_3644_ (
  .A1({ S25957[1125] }),
  .A2({ S25957[1221] }),
  .ZN({ S21655 })
);
NAND3_X1 #() 
NAND3_X1_3873_ (
  .A1({ S21655 }),
  .A2({ S11631 }),
  .A3({ S21654 }),
  .ZN({ S21656 })
);
NAND2_X1 #() 
NAND2_X1_3645_ (
  .A1({ S21656 }),
  .A2({ S21653 }),
  .ZN({ S25957[1029] })
);
NOR2_X1 #() 
NOR2_X1_921_ (
  .A1({ S19308 }),
  .A2({ S19306 }),
  .ZN({ S25957[1188] })
);
INV_X1 #() 
INV_X1_1212_ (
  .A({ S25957[1188] }),
  .ZN({ S21657 })
);
NAND3_X1 #() 
NAND3_X1_3874_ (
  .A1({ S25957[1178] }),
  .A2({ S21408 }),
  .A3({ S21399 }),
  .ZN({ S21658 })
);
NAND2_X1 #() 
NAND2_X1_3646_ (
  .A1({ S21658 }),
  .A2({ S71 }),
  .ZN({ S21659 })
);
NAND2_X1 #() 
NAND2_X1_3647_ (
  .A1({ S21625 }),
  .A2({ S21659 }),
  .ZN({ S21660 })
);
OAI211_X1 #() 
OAI211_X1_1259_ (
  .A({ S71 }),
  .B({ S21408 }),
  .C1({ S25957[1178] }),
  .C2({ S21399 }),
  .ZN({ S21661 })
);
OAI211_X1 #() 
OAI211_X1_1260_ (
  .A({ S21661 }),
  .B({ S21398 }),
  .C1({ S21494 }),
  .C2({ S21420 }),
  .ZN({ S21662 })
);
NAND3_X1 #() 
NAND3_X1_3875_ (
  .A1({ S21660 }),
  .A2({ S21662 }),
  .A3({ S25957[1181] }),
  .ZN({ S21663 })
);
INV_X1 #() 
INV_X1_1213_ (
  .A({ S21439 }),
  .ZN({ S21664 })
);
NOR2_X1 #() 
NOR2_X1_922_ (
  .A1({ S21664 }),
  .A2({ S21455 }),
  .ZN({ S21665 })
);
NOR2_X1 #() 
NOR2_X1_923_ (
  .A1({ S21420 }),
  .A2({ S21404 }),
  .ZN({ S21666 })
);
OAI21_X1 #() 
OAI21_X1_1871_ (
  .A({ S25957[1180] }),
  .B1({ S21666 }),
  .B2({ S21665 }),
  .ZN({ S21667 })
);
AOI22_X1 #() 
AOI22_X1_415_ (
  .A1({ S21535 }),
  .A2({ S21493 }),
  .B1({ S21411 }),
  .B2({ S21399 }),
  .ZN({ S21668 })
);
OAI21_X1 #() 
OAI21_X1_1872_ (
  .A({ S21398 }),
  .B1({ S21491 }),
  .B2({ S21668 }),
  .ZN({ S21669 })
);
NAND2_X1 #() 
NAND2_X1_3648_ (
  .A1({ S21667 }),
  .A2({ S21669 }),
  .ZN({ S21670 })
);
NAND2_X1 #() 
NAND2_X1_3649_ (
  .A1({ S21670 }),
  .A2({ S21444 }),
  .ZN({ S21671 })
);
NAND3_X1 #() 
NAND3_X1_3876_ (
  .A1({ S21671 }),
  .A2({ S25957[1182] }),
  .A3({ S21663 }),
  .ZN({ S21672 })
);
AOI21_X1 #() 
AOI21_X1_1972_ (
  .A({ S25957[1179] }),
  .B1({ S21435 }),
  .B2({ S21480 }),
  .ZN({ S21673 })
);
NAND3_X1 #() 
NAND3_X1_3877_ (
  .A1({ S25957[1179] }),
  .A2({ S21408 }),
  .A3({ S25957[1177] }),
  .ZN({ S21674 })
);
NAND2_X1 #() 
NAND2_X1_3650_ (
  .A1({ S21624 }),
  .A2({ S21674 }),
  .ZN({ S21675 })
);
OR2_X1 #() 
OR2_X1_51_ (
  .A1({ S21673 }),
  .A2({ S21675 }),
  .ZN({ S21676 })
);
NAND2_X1 #() 
NAND2_X1_3651_ (
  .A1({ S21417 }),
  .A2({ S21535 }),
  .ZN({ S21677 })
);
NAND2_X1 #() 
NAND2_X1_3652_ (
  .A1({ S21616 }),
  .A2({ S21677 }),
  .ZN({ S21678 })
);
AOI21_X1 #() 
AOI21_X1_1973_ (
  .A({ S21444 }),
  .B1({ S21678 }),
  .B2({ S25957[1180] }),
  .ZN({ S21679 })
);
OAI21_X1 #() 
OAI21_X1_1873_ (
  .A({ S21679 }),
  .B1({ S21676 }),
  .B2({ S25957[1180] }),
  .ZN({ S21680 })
);
NAND3_X1 #() 
NAND3_X1_3878_ (
  .A1({ S21522 }),
  .A2({ S21465 }),
  .A3({ S71 }),
  .ZN({ S21681 })
);
OAI211_X1 #() 
OAI211_X1_1261_ (
  .A({ S25957[1180] }),
  .B({ S21681 }),
  .C1({ S21403 }),
  .C2({ S21547 }),
  .ZN({ S21682 })
);
NOR2_X1 #() 
NOR2_X1_924_ (
  .A1({ S21452 }),
  .A2({ S21455 }),
  .ZN({ S21683 })
);
AOI21_X1 #() 
AOI21_X1_1974_ (
  .A({ S25957[1179] }),
  .B1({ S21522 }),
  .B2({ S21531 }),
  .ZN({ S21684 })
);
INV_X1 #() 
INV_X1_1214_ (
  .A({ S21684 }),
  .ZN({ S21685 })
);
NAND2_X1 #() 
NAND2_X1_3653_ (
  .A1({ S21685 }),
  .A2({ S21398 }),
  .ZN({ S21686 })
);
OAI211_X1 #() 
OAI211_X1_1262_ (
  .A({ S21682 }),
  .B({ S21444 }),
  .C1({ S21686 }),
  .C2({ S21683 }),
  .ZN({ S21687 })
);
NAND3_X1 #() 
NAND3_X1_3879_ (
  .A1({ S21687 }),
  .A2({ S21680 }),
  .A3({ S21433 }),
  .ZN({ S21688 })
);
NAND3_X1 #() 
NAND3_X1_3880_ (
  .A1({ S21688 }),
  .A2({ S25957[1183] }),
  .A3({ S21672 }),
  .ZN({ S21689 })
);
NAND2_X1 #() 
NAND2_X1_3654_ (
  .A1({ S21407 }),
  .A2({ S71 }),
  .ZN({ S21690 })
);
NOR2_X1 #() 
NOR2_X1_925_ (
  .A1({ S21690 }),
  .A2({ S21420 }),
  .ZN({ S21691 })
);
NAND3_X1 #() 
NAND3_X1_3881_ (
  .A1({ S21465 }),
  .A2({ S71 }),
  .A3({ S21540 }),
  .ZN({ S21692 })
);
AOI21_X1 #() 
AOI21_X1_1975_ (
  .A({ S25957[1180] }),
  .B1({ S25957[1179] }),
  .B2({ S25957[1178] }),
  .ZN({ S21693 })
);
NAND2_X1 #() 
NAND2_X1_3655_ (
  .A1({ S21692 }),
  .A2({ S21693 }),
  .ZN({ S21694 })
);
OAI21_X1 #() 
OAI21_X1_1874_ (
  .A({ S21694 }),
  .B1({ S21691 }),
  .B2({ S21526 }),
  .ZN({ S21695 })
);
INV_X1 #() 
INV_X1_1215_ (
  .A({ S122 }),
  .ZN({ S21696 })
);
OAI21_X1 #() 
OAI21_X1_1875_ (
  .A({ S25957[1180] }),
  .B1({ S21696 }),
  .B2({ S25957[1178] }),
  .ZN({ S21697 })
);
NAND4_X1 #() 
NAND4_X1_427_ (
  .A1({ S21394 }),
  .A2({ S79 }),
  .A3({ S71 }),
  .A4({ S21411 }),
  .ZN({ S21698 })
);
NAND4_X1 #() 
NAND4_X1_428_ (
  .A1({ S21608 }),
  .A2({ S21620 }),
  .A3({ S21398 }),
  .A4({ S21698 }),
  .ZN({ S21699 })
);
NAND3_X1 #() 
NAND3_X1_3882_ (
  .A1({ S21699 }),
  .A2({ S25957[1181] }),
  .A3({ S21697 }),
  .ZN({ S21700 })
);
OAI211_X1 #() 
OAI211_X1_1263_ (
  .A({ S21700 }),
  .B({ S25957[1182] }),
  .C1({ S21695 }),
  .C2({ S25957[1181] }),
  .ZN({ S21701 })
);
AOI21_X1 #() 
AOI21_X1_1976_ (
  .A({ S21631 }),
  .B1({ S21592 }),
  .B2({ S25957[1179] }),
  .ZN({ S21702 })
);
NAND3_X1 #() 
NAND3_X1_3883_ (
  .A1({ S21608 }),
  .A2({ S21474 }),
  .A3({ S25957[1180] }),
  .ZN({ S21703 })
);
OAI21_X1 #() 
OAI21_X1_1876_ (
  .A({ S21703 }),
  .B1({ S25957[1180] }),
  .B2({ S21702 }),
  .ZN({ S21704 })
);
NAND2_X1 #() 
NAND2_X1_3656_ (
  .A1({ S21704 }),
  .A2({ S25957[1181] }),
  .ZN({ S21705 })
);
NAND2_X1 #() 
NAND2_X1_3657_ (
  .A1({ S21439 }),
  .A2({ S21401 }),
  .ZN({ S21706 })
);
NAND2_X1 #() 
NAND2_X1_3658_ (
  .A1({ S21706 }),
  .A2({ S25957[1179] }),
  .ZN({ S21707 })
);
NAND3_X1 #() 
NAND3_X1_3884_ (
  .A1({ S21658 }),
  .A2({ S21529 }),
  .A3({ S71 }),
  .ZN({ S21708 })
);
AOI21_X1 #() 
AOI21_X1_1977_ (
  .A({ S25957[1180] }),
  .B1({ S21708 }),
  .B2({ S21707 }),
  .ZN({ S21709 })
);
NAND3_X1 #() 
NAND3_X1_3885_ (
  .A1({ S21473 }),
  .A2({ S25957[1179] }),
  .A3({ S21423 }),
  .ZN({ S21710 })
);
AND3_X1 #() 
AND3_X1_139_ (
  .A1({ S21586 }),
  .A2({ S25957[1180] }),
  .A3({ S21710 }),
  .ZN({ S21711 })
);
OAI21_X1 #() 
OAI21_X1_1877_ (
  .A({ S21444 }),
  .B1({ S21711 }),
  .B2({ S21709 }),
  .ZN({ S21712 })
);
NAND3_X1 #() 
NAND3_X1_3886_ (
  .A1({ S21705 }),
  .A2({ S21712 }),
  .A3({ S21433 }),
  .ZN({ S21713 })
);
NAND3_X1 #() 
NAND3_X1_3887_ (
  .A1({ S21713 }),
  .A2({ S21701 }),
  .A3({ S21395 }),
  .ZN({ S21714 })
);
NAND3_X1 #() 
NAND3_X1_3888_ (
  .A1({ S21689 }),
  .A2({ S21714 }),
  .A3({ S25957[1252] }),
  .ZN({ S21715 })
);
NAND2_X1 #() 
NAND2_X1_3659_ (
  .A1({ S21660 }),
  .A2({ S21662 }),
  .ZN({ S21716 })
);
NAND2_X1 #() 
NAND2_X1_3660_ (
  .A1({ S21716 }),
  .A2({ S25957[1181] }),
  .ZN({ S21717 })
);
OAI211_X1 #() 
OAI211_X1_1264_ (
  .A({ S21717 }),
  .B({ S25957[1182] }),
  .C1({ S25957[1181] }),
  .C2({ S21670 }),
  .ZN({ S21718 })
);
OAI21_X1 #() 
OAI21_X1_1878_ (
  .A({ S21398 }),
  .B1({ S21673 }),
  .B2({ S21675 }),
  .ZN({ S21719 })
);
OAI211_X1 #() 
OAI211_X1_1265_ (
  .A({ S21719 }),
  .B({ S25957[1181] }),
  .C1({ S21398 }),
  .C2({ S21678 }),
  .ZN({ S21720 })
);
OAI21_X1 #() 
OAI21_X1_1879_ (
  .A({ S21681 }),
  .B1({ S21403 }),
  .B2({ S21547 }),
  .ZN({ S21721 })
);
NAND2_X1 #() 
NAND2_X1_3661_ (
  .A1({ S21721 }),
  .A2({ S25957[1180] }),
  .ZN({ S21722 })
);
OAI21_X1 #() 
OAI21_X1_1880_ (
  .A({ S21398 }),
  .B1({ S21684 }),
  .B2({ S21683 }),
  .ZN({ S21723 })
);
NAND3_X1 #() 
NAND3_X1_3889_ (
  .A1({ S21722 }),
  .A2({ S21444 }),
  .A3({ S21723 }),
  .ZN({ S21724 })
);
NAND3_X1 #() 
NAND3_X1_3890_ (
  .A1({ S21724 }),
  .A2({ S21720 }),
  .A3({ S21433 }),
  .ZN({ S21725 })
);
NAND3_X1 #() 
NAND3_X1_3891_ (
  .A1({ S21725 }),
  .A2({ S21718 }),
  .A3({ S25957[1183] }),
  .ZN({ S21726 })
);
OAI21_X1 #() 
OAI21_X1_1881_ (
  .A({ S21700 }),
  .B1({ S21695 }),
  .B2({ S25957[1181] }),
  .ZN({ S21727 })
);
NAND2_X1 #() 
NAND2_X1_3662_ (
  .A1({ S21727 }),
  .A2({ S25957[1182] }),
  .ZN({ S21728 })
);
OAI211_X1 #() 
OAI211_X1_1266_ (
  .A({ S21703 }),
  .B({ S25957[1181] }),
  .C1({ S25957[1180] }),
  .C2({ S21702 }),
  .ZN({ S21729 })
);
NAND3_X1 #() 
NAND3_X1_3892_ (
  .A1({ S21586 }),
  .A2({ S21710 }),
  .A3({ S25957[1180] }),
  .ZN({ S21730 })
);
NAND2_X1 #() 
NAND2_X1_3663_ (
  .A1({ S21730 }),
  .A2({ S21444 }),
  .ZN({ S21731 })
);
OAI211_X1 #() 
OAI211_X1_1267_ (
  .A({ S21729 }),
  .B({ S21433 }),
  .C1({ S21709 }),
  .C2({ S21731 }),
  .ZN({ S21732 })
);
NAND3_X1 #() 
NAND3_X1_3893_ (
  .A1({ S21728 }),
  .A2({ S21395 }),
  .A3({ S21732 }),
  .ZN({ S21733 })
);
NAND3_X1 #() 
NAND3_X1_3894_ (
  .A1({ S21733 }),
  .A2({ S21726 }),
  .A3({ S19304 }),
  .ZN({ S21734 })
);
NAND3_X1 #() 
NAND3_X1_3895_ (
  .A1({ S21734 }),
  .A2({ S21715 }),
  .A3({ S19311 }),
  .ZN({ S21735 })
);
NAND3_X1 #() 
NAND3_X1_3896_ (
  .A1({ S21733 }),
  .A2({ S21726 }),
  .A3({ S25957[1252] }),
  .ZN({ S21736 })
);
NAND3_X1 #() 
NAND3_X1_3897_ (
  .A1({ S21689 }),
  .A2({ S21714 }),
  .A3({ S19304 }),
  .ZN({ S21737 })
);
NAND3_X1 #() 
NAND3_X1_3898_ (
  .A1({ S21736 }),
  .A2({ S21737 }),
  .A3({ S25957[1220] }),
  .ZN({ S21738 })
);
NAND3_X1 #() 
NAND3_X1_3899_ (
  .A1({ S21735 }),
  .A2({ S21738 }),
  .A3({ S21657 }),
  .ZN({ S21739 })
);
NAND3_X1 #() 
NAND3_X1_3900_ (
  .A1({ S21734 }),
  .A2({ S21715 }),
  .A3({ S25957[1220] }),
  .ZN({ S21740 })
);
NAND3_X1 #() 
NAND3_X1_3901_ (
  .A1({ S21736 }),
  .A2({ S21737 }),
  .A3({ S19311 }),
  .ZN({ S21741 })
);
NAND3_X1 #() 
NAND3_X1_3902_ (
  .A1({ S21740 }),
  .A2({ S21741 }),
  .A3({ S25957[1188] }),
  .ZN({ S21742 })
);
NAND3_X1 #() 
NAND3_X1_3903_ (
  .A1({ S21739 }),
  .A2({ S21742 }),
  .A3({ S20774 }),
  .ZN({ S21743 })
);
NAND3_X1 #() 
NAND3_X1_3904_ (
  .A1({ S21740 }),
  .A2({ S21741 }),
  .A3({ S21657 }),
  .ZN({ S21744 })
);
NAND3_X1 #() 
NAND3_X1_3905_ (
  .A1({ S21735 }),
  .A2({ S21738 }),
  .A3({ S25957[1188] }),
  .ZN({ S21745 })
);
NAND3_X1 #() 
NAND3_X1_3906_ (
  .A1({ S21744 }),
  .A2({ S21745 }),
  .A3({ S25957[1156] }),
  .ZN({ S21746 })
);
NAND2_X1 #() 
NAND2_X1_3664_ (
  .A1({ S21743 }),
  .A2({ S21746 }),
  .ZN({ S25957[1028] })
);
NAND2_X1 #() 
NAND2_X1_3665_ (
  .A1({ S19369 }),
  .A2({ S19367 }),
  .ZN({ S25957[1219] })
);
NAND4_X1 #() 
NAND4_X1_429_ (
  .A1({ S21540 }),
  .A2({ S21416 }),
  .A3({ S21401 }),
  .A4({ S71 }),
  .ZN({ S21747 })
);
NAND3_X1 #() 
NAND3_X1_3907_ (
  .A1({ S21445 }),
  .A2({ S21531 }),
  .A3({ S25957[1179] }),
  .ZN({ S21748 })
);
AOI21_X1 #() 
AOI21_X1_1978_ (
  .A({ S25957[1180] }),
  .B1({ S21748 }),
  .B2({ S21747 }),
  .ZN({ S21749 })
);
NAND3_X1 #() 
NAND3_X1_3908_ (
  .A1({ S21522 }),
  .A2({ S71 }),
  .A3({ S21416 }),
  .ZN({ S21750 })
);
AOI21_X1 #() 
AOI21_X1_1979_ (
  .A({ S21398 }),
  .B1({ S21706 }),
  .B2({ S25957[1179] }),
  .ZN({ S21751 })
);
NAND2_X1 #() 
NAND2_X1_3666_ (
  .A1({ S21751 }),
  .A2({ S21750 }),
  .ZN({ S21752 })
);
NAND2_X1 #() 
NAND2_X1_3667_ (
  .A1({ S21752 }),
  .A2({ S25957[1181] }),
  .ZN({ S21753 })
);
NOR2_X1 #() 
NOR2_X1_926_ (
  .A1({ S21753 }),
  .A2({ S21749 }),
  .ZN({ S21754 })
);
NAND2_X1 #() 
NAND2_X1_3668_ (
  .A1({ S21483 }),
  .A2({ S71 }),
  .ZN({ S21755 })
);
OAI21_X1 #() 
OAI21_X1_1882_ (
  .A({ S21603 }),
  .B1({ S21755 }),
  .B2({ S21633 }),
  .ZN({ S21756 })
);
OAI211_X1 #() 
OAI211_X1_1268_ (
  .A({ S21567 }),
  .B({ S21398 }),
  .C1({ S71 }),
  .C2({ S21411 }),
  .ZN({ S21757 })
);
NAND2_X1 #() 
NAND2_X1_3669_ (
  .A1({ S21757 }),
  .A2({ S21444 }),
  .ZN({ S21758 })
);
AOI21_X1 #() 
AOI21_X1_1980_ (
  .A({ S21758 }),
  .B1({ S21756 }),
  .B2({ S25957[1180] }),
  .ZN({ S21759 })
);
OAI21_X1 #() 
OAI21_X1_1883_ (
  .A({ S25957[1182] }),
  .B1({ S21754 }),
  .B2({ S21759 }),
  .ZN({ S21760 })
);
NAND3_X1 #() 
NAND3_X1_3909_ (
  .A1({ S21434 }),
  .A2({ S71 }),
  .A3({ S21400 }),
  .ZN({ S21761 })
);
NAND4_X1 #() 
NAND4_X1_430_ (
  .A1({ S21540 }),
  .A2({ S21439 }),
  .A3({ S25957[1179] }),
  .A4({ S25957[1177] }),
  .ZN({ S21762 })
);
AND2_X1 #() 
AND2_X1_225_ (
  .A1({ S21762 }),
  .A2({ S21398 }),
  .ZN({ S21763 })
);
NAND2_X1 #() 
NAND2_X1_3670_ (
  .A1({ S21445 }),
  .A2({ S21439 }),
  .ZN({ S21764 })
);
NAND2_X1 #() 
NAND2_X1_3671_ (
  .A1({ S21764 }),
  .A2({ S71 }),
  .ZN({ S21765 })
);
AOI21_X1 #() 
AOI21_X1_1981_ (
  .A({ S21398 }),
  .B1({ S21467 }),
  .B2({ S21446 }),
  .ZN({ S21766 })
);
AOI22_X1 #() 
AOI22_X1_416_ (
  .A1({ S21766 }),
  .A2({ S21765 }),
  .B1({ S21763 }),
  .B2({ S21761 }),
  .ZN({ S21767 })
);
NAND2_X1 #() 
NAND2_X1_3672_ (
  .A1({ S21417 }),
  .A2({ S25957[1179] }),
  .ZN({ S21768 })
);
NAND2_X1 #() 
NAND2_X1_3673_ (
  .A1({ S21609 }),
  .A2({ S21768 }),
  .ZN({ S21769 })
);
OAI21_X1 #() 
OAI21_X1_1884_ (
  .A({ S25957[1180] }),
  .B1({ S21769 }),
  .B2({ S21668 }),
  .ZN({ S21770 })
);
NAND2_X1 #() 
NAND2_X1_3674_ (
  .A1({ S21600 }),
  .A2({ S21622 }),
  .ZN({ S21771 })
);
AOI21_X1 #() 
AOI21_X1_1982_ (
  .A({ S21424 }),
  .B1({ S21771 }),
  .B2({ S25957[1179] }),
  .ZN({ S21772 })
);
NAND2_X1 #() 
NAND2_X1_3675_ (
  .A1({ S21772 }),
  .A2({ S21398 }),
  .ZN({ S21773 })
);
NAND3_X1 #() 
NAND3_X1_3910_ (
  .A1({ S21773 }),
  .A2({ S21444 }),
  .A3({ S21770 }),
  .ZN({ S21774 })
);
OAI211_X1 #() 
OAI211_X1_1269_ (
  .A({ S21774 }),
  .B({ S21433 }),
  .C1({ S21767 }),
  .C2({ S21444 }),
  .ZN({ S21775 })
);
NAND3_X1 #() 
NAND3_X1_3911_ (
  .A1({ S21775 }),
  .A2({ S21760 }),
  .A3({ S25957[1183] }),
  .ZN({ S21776 })
);
OAI21_X1 #() 
OAI21_X1_1885_ (
  .A({ S79 }),
  .B1({ S21394 }),
  .B2({ S25957[1178] }),
  .ZN({ S21777 })
);
OAI21_X1 #() 
OAI21_X1_1886_ (
  .A({ S21614 }),
  .B1({ S71 }),
  .B2({ S21777 }),
  .ZN({ S21778 })
);
NOR2_X1 #() 
NOR2_X1_927_ (
  .A1({ S21778 }),
  .A2({ S21398 }),
  .ZN({ S21779 })
);
AND2_X1 #() 
AND2_X1_226_ (
  .A1({ S21483 }),
  .A2({ S21428 }),
  .ZN({ S21780 })
);
NAND2_X1 #() 
NAND2_X1_3676_ (
  .A1({ S21427 }),
  .A2({ S21465 }),
  .ZN({ S21781 })
);
OAI211_X1 #() 
OAI211_X1_1270_ (
  .A({ S21398 }),
  .B({ S21781 }),
  .C1({ S21780 }),
  .C2({ S25957[1179] }),
  .ZN({ S21782 })
);
NAND2_X1 #() 
NAND2_X1_3677_ (
  .A1({ S21782 }),
  .A2({ S21444 }),
  .ZN({ S21783 })
);
NAND3_X1 #() 
NAND3_X1_3912_ (
  .A1({ S21755 }),
  .A2({ S25957[1180] }),
  .A3({ S21466 }),
  .ZN({ S21784 })
);
NAND4_X1 #() 
NAND4_X1_431_ (
  .A1({ S21559 }),
  .A2({ S21398 }),
  .A3({ S21540 }),
  .A4({ S21473 }),
  .ZN({ S21785 })
);
NAND3_X1 #() 
NAND3_X1_3913_ (
  .A1({ S21784 }),
  .A2({ S21785 }),
  .A3({ S25957[1181] }),
  .ZN({ S21786 })
);
OAI211_X1 #() 
OAI211_X1_1271_ (
  .A({ S21433 }),
  .B({ S21786 }),
  .C1({ S21783 }),
  .C2({ S21779 }),
  .ZN({ S21787 })
);
NAND3_X1 #() 
NAND3_X1_3914_ (
  .A1({ S21606 }),
  .A2({ S21498 }),
  .A3({ S25957[1180] }),
  .ZN({ S21788 })
);
INV_X1 #() 
INV_X1_1216_ (
  .A({ S79 }),
  .ZN({ S21789 })
);
NOR2_X1 #() 
NOR2_X1_928_ (
  .A1({ S21411 }),
  .A2({ S21399 }),
  .ZN({ S21790 })
);
OAI21_X1 #() 
OAI21_X1_1887_ (
  .A({ S71 }),
  .B1({ S21790 }),
  .B2({ S21789 }),
  .ZN({ S21791 })
);
AOI21_X1 #() 
AOI21_X1_1983_ (
  .A({ S25957[1180] }),
  .B1({ S21459 }),
  .B2({ S21438 }),
  .ZN({ S21792 })
);
AOI21_X1 #() 
AOI21_X1_1984_ (
  .A({ S21444 }),
  .B1({ S21792 }),
  .B2({ S21791 }),
  .ZN({ S21793 })
);
NAND2_X1 #() 
NAND2_X1_3678_ (
  .A1({ S21788 }),
  .A2({ S21793 }),
  .ZN({ S21794 })
);
NAND3_X1 #() 
NAND3_X1_3915_ (
  .A1({ S21423 }),
  .A2({ S21394 }),
  .A3({ S71 }),
  .ZN({ S21795 })
);
NOR2_X1 #() 
NOR2_X1_929_ (
  .A1({ S21795 }),
  .A2({ S21398 }),
  .ZN({ S21796 })
);
AOI21_X1 #() 
AOI21_X1_1985_ (
  .A({ S21796 }),
  .B1({ S21482 }),
  .B2({ S21710 }),
  .ZN({ S21797 })
);
OAI211_X1 #() 
OAI211_X1_1272_ (
  .A({ S21794 }),
  .B({ S25957[1182] }),
  .C1({ S21797 }),
  .C2({ S25957[1181] }),
  .ZN({ S21798 })
);
NAND3_X1 #() 
NAND3_X1_3916_ (
  .A1({ S21787 }),
  .A2({ S21395 }),
  .A3({ S21798 }),
  .ZN({ S21799 })
);
NAND3_X1 #() 
NAND3_X1_3917_ (
  .A1({ S21776 }),
  .A2({ S21799 }),
  .A3({ S25957[1251] }),
  .ZN({ S21800 })
);
INV_X1 #() 
INV_X1_1217_ (
  .A({ S21749 }),
  .ZN({ S21801 })
);
NAND3_X1 #() 
NAND3_X1_3918_ (
  .A1({ S21801 }),
  .A2({ S25957[1181] }),
  .A3({ S21752 }),
  .ZN({ S21802 })
);
AND2_X1 #() 
AND2_X1_227_ (
  .A1({ S21756 }),
  .A2({ S25957[1180] }),
  .ZN({ S21803 })
);
OAI211_X1 #() 
OAI211_X1_1273_ (
  .A({ S21802 }),
  .B({ S25957[1182] }),
  .C1({ S21803 }),
  .C2({ S21758 }),
  .ZN({ S21804 })
);
NAND3_X1 #() 
NAND3_X1_3919_ (
  .A1({ S21400 }),
  .A2({ S71 }),
  .A3({ S21540 }),
  .ZN({ S21805 })
);
NAND2_X1 #() 
NAND2_X1_3679_ (
  .A1({ S21805 }),
  .A2({ S25957[1180] }),
  .ZN({ S21806 })
);
OAI221_X1 #() 
OAI221_X1_109_ (
  .A({ S21444 }),
  .B1({ S21769 }),
  .B2({ S21806 }),
  .C1({ S21772 }),
  .C2({ S25957[1180] }),
  .ZN({ S21807 })
);
NAND2_X1 #() 
NAND2_X1_3680_ (
  .A1({ S21763 }),
  .A2({ S21761 }),
  .ZN({ S21808 })
);
NAND2_X1 #() 
NAND2_X1_3681_ (
  .A1({ S21766 }),
  .A2({ S21765 }),
  .ZN({ S21809 })
);
NAND3_X1 #() 
NAND3_X1_3920_ (
  .A1({ S21809 }),
  .A2({ S21808 }),
  .A3({ S25957[1181] }),
  .ZN({ S21810 })
);
NAND3_X1 #() 
NAND3_X1_3921_ (
  .A1({ S21807 }),
  .A2({ S21810 }),
  .A3({ S21433 }),
  .ZN({ S21811 })
);
NAND3_X1 #() 
NAND3_X1_3922_ (
  .A1({ S21804 }),
  .A2({ S21811 }),
  .A3({ S25957[1183] }),
  .ZN({ S21812 })
);
NAND2_X1 #() 
NAND2_X1_3682_ (
  .A1({ S21482 }),
  .A2({ S21710 }),
  .ZN({ S21813 })
);
NOR2_X1 #() 
NOR2_X1_930_ (
  .A1({ S21796 }),
  .A2({ S25957[1181] }),
  .ZN({ S21814 })
);
NAND2_X1 #() 
NAND2_X1_3683_ (
  .A1({ S21813 }),
  .A2({ S21814 }),
  .ZN({ S21815 })
);
NOR2_X1 #() 
NOR2_X1_931_ (
  .A1({ S21516 }),
  .A2({ S21398 }),
  .ZN({ S21816 })
);
AOI22_X1 #() 
AOI22_X1_417_ (
  .A1({ S21816 }),
  .A2({ S21498 }),
  .B1({ S21791 }),
  .B2({ S21792 }),
  .ZN({ S21817 })
);
OAI211_X1 #() 
OAI211_X1_1274_ (
  .A({ S21815 }),
  .B({ S25957[1182] }),
  .C1({ S21817 }),
  .C2({ S21444 }),
  .ZN({ S21818 })
);
INV_X1 #() 
INV_X1_1218_ (
  .A({ S21781 }),
  .ZN({ S21819 })
);
OAI21_X1 #() 
OAI21_X1_1888_ (
  .A({ S21398 }),
  .B1({ S21819 }),
  .B2({ S21484 }),
  .ZN({ S21820 })
);
AOI21_X1 #() 
AOI21_X1_1986_ (
  .A({ S25957[1181] }),
  .B1({ S21778 }),
  .B2({ S25957[1180] }),
  .ZN({ S21821 })
);
NAND2_X1 #() 
NAND2_X1_3684_ (
  .A1({ S21821 }),
  .A2({ S21820 }),
  .ZN({ S21822 })
);
NAND2_X1 #() 
NAND2_X1_3685_ (
  .A1({ S21784 }),
  .A2({ S21785 }),
  .ZN({ S21823 })
);
NAND2_X1 #() 
NAND2_X1_3686_ (
  .A1({ S21823 }),
  .A2({ S25957[1181] }),
  .ZN({ S21824 })
);
NAND3_X1 #() 
NAND3_X1_3923_ (
  .A1({ S21822 }),
  .A2({ S21824 }),
  .A3({ S21433 }),
  .ZN({ S21825 })
);
NAND3_X1 #() 
NAND3_X1_3924_ (
  .A1({ S21825 }),
  .A2({ S21818 }),
  .A3({ S21395 }),
  .ZN({ S21826 })
);
NAND3_X1 #() 
NAND3_X1_3925_ (
  .A1({ S21812 }),
  .A2({ S21826 }),
  .A3({ S19368 }),
  .ZN({ S21827 })
);
NAND3_X1 #() 
NAND3_X1_3926_ (
  .A1({ S21800 }),
  .A2({ S21827 }),
  .A3({ S25957[1219] }),
  .ZN({ S21828 })
);
INV_X1 #() 
INV_X1_1219_ (
  .A({ S25957[1219] }),
  .ZN({ S21829 })
);
NAND3_X1 #() 
NAND3_X1_3927_ (
  .A1({ S21776 }),
  .A2({ S21799 }),
  .A3({ S19368 }),
  .ZN({ S21830 })
);
NAND3_X1 #() 
NAND3_X1_3928_ (
  .A1({ S21812 }),
  .A2({ S21826 }),
  .A3({ S25957[1251] }),
  .ZN({ S21831 })
);
NAND3_X1 #() 
NAND3_X1_3929_ (
  .A1({ S21830 }),
  .A2({ S21831 }),
  .A3({ S21829 }),
  .ZN({ S21832 })
);
NAND3_X1 #() 
NAND3_X1_3930_ (
  .A1({ S21828 }),
  .A2({ S21832 }),
  .A3({ S25956[3] }),
  .ZN({ S21833 })
);
NAND3_X1 #() 
NAND3_X1_3931_ (
  .A1({ S21800 }),
  .A2({ S21827 }),
  .A3({ S21829 }),
  .ZN({ S21834 })
);
NAND3_X1 #() 
NAND3_X1_3932_ (
  .A1({ S21830 }),
  .A2({ S21831 }),
  .A3({ S25957[1219] }),
  .ZN({ S21835 })
);
NAND3_X1 #() 
NAND3_X1_3933_ (
  .A1({ S21834 }),
  .A2({ S21835 }),
  .A3({ S11664 }),
  .ZN({ S21836 })
);
NAND2_X1 #() 
NAND2_X1_3687_ (
  .A1({ S21833 }),
  .A2({ S21836 }),
  .ZN({ S80 })
);
AND2_X1 #() 
AND2_X1_228_ (
  .A1({ S21836 }),
  .A2({ S21833 }),
  .ZN({ S25957[1027] })
);
NAND2_X1 #() 
NAND2_X1_3688_ (
  .A1({ S19425 }),
  .A2({ S19426 }),
  .ZN({ S25957[1216] })
);
INV_X1 #() 
INV_X1_1220_ (
  .A({ S25957[1216] }),
  .ZN({ S21837 })
);
INV_X1 #() 
INV_X1_1221_ (
  .A({ S25957[1248] }),
  .ZN({ S21838 })
);
NAND3_X1 #() 
NAND3_X1_3934_ (
  .A1({ S21445 }),
  .A2({ S21531 }),
  .A3({ S71 }),
  .ZN({ S21839 })
);
AOI21_X1 #() 
AOI21_X1_1987_ (
  .A({ S21398 }),
  .B1({ S21634 }),
  .B2({ S21839 }),
  .ZN({ S21840 })
);
NAND3_X1 #() 
NAND3_X1_3935_ (
  .A1({ S21620 }),
  .A2({ S21398 }),
  .A3({ S21619 }),
  .ZN({ S21841 })
);
INV_X1 #() 
INV_X1_1222_ (
  .A({ S21841 }),
  .ZN({ S21842 })
);
OAI21_X1 #() 
OAI21_X1_1889_ (
  .A({ S21444 }),
  .B1({ S21842 }),
  .B2({ S21840 }),
  .ZN({ S21843 })
);
OAI211_X1 #() 
OAI211_X1_1275_ (
  .A({ S21540 }),
  .B({ S25957[1179] }),
  .C1({ S21416 }),
  .C2({ S25957[1178] }),
  .ZN({ S21844 })
);
NAND2_X1 #() 
NAND2_X1_3689_ (
  .A1({ S21438 }),
  .A2({ S71 }),
  .ZN({ S21845 })
);
OAI211_X1 #() 
OAI211_X1_1276_ (
  .A({ S21844 }),
  .B({ S21398 }),
  .C1({ S21845 }),
  .C2({ S21592 }),
  .ZN({ S21846 })
);
NOR2_X1 #() 
NOR2_X1_932_ (
  .A1({ S71 }),
  .A2({ S21411 }),
  .ZN({ S21847 })
);
AOI22_X1 #() 
AOI22_X1_418_ (
  .A1({ S21413 }),
  .A2({ S71 }),
  .B1({ S21847 }),
  .B2({ S21401 }),
  .ZN({ S21848 })
);
OAI211_X1 #() 
OAI211_X1_1277_ (
  .A({ S25957[1181] }),
  .B({ S21846 }),
  .C1({ S21848 }),
  .C2({ S21398 }),
  .ZN({ S21849 })
);
AOI21_X1 #() 
AOI21_X1_1988_ (
  .A({ S21433 }),
  .B1({ S21843 }),
  .B2({ S21849 }),
  .ZN({ S21850 })
);
AOI22_X1 #() 
AOI22_X1_419_ (
  .A1({ S21466 }),
  .A2({ S21795 }),
  .B1({ S21489 }),
  .B2({ S21408 }),
  .ZN({ S21851 })
);
NAND4_X1 #() 
NAND4_X1_432_ (
  .A1({ S21659 }),
  .A2({ S21624 }),
  .A3({ S21398 }),
  .A4({ S21674 }),
  .ZN({ S21852 })
);
OAI211_X1 #() 
OAI211_X1_1278_ (
  .A({ S25957[1181] }),
  .B({ S21852 }),
  .C1({ S21851 }),
  .C2({ S21398 }),
  .ZN({ S21853 })
);
NAND2_X1 #() 
NAND2_X1_3690_ (
  .A1({ S21438 }),
  .A2({ S25957[1179] }),
  .ZN({ S21854 })
);
OAI211_X1 #() 
OAI211_X1_1279_ (
  .A({ S21854 }),
  .B({ S25957[1180] }),
  .C1({ S21592 }),
  .C2({ S25957[1179] }),
  .ZN({ S21855 })
);
NAND4_X1 #() 
NAND4_X1_433_ (
  .A1({ S21423 }),
  .A2({ S21428 }),
  .A3({ S71 }),
  .A4({ S79 }),
  .ZN({ S21856 })
);
AOI21_X1 #() 
AOI21_X1_1989_ (
  .A({ S25957[1181] }),
  .B1({ S21792 }),
  .B2({ S21856 }),
  .ZN({ S21857 })
);
AOI21_X1 #() 
AOI21_X1_1990_ (
  .A({ S25957[1182] }),
  .B1({ S21857 }),
  .B2({ S21855 }),
  .ZN({ S21858 })
);
NAND2_X1 #() 
NAND2_X1_3691_ (
  .A1({ S21858 }),
  .A2({ S21853 }),
  .ZN({ S21859 })
);
NAND2_X1 #() 
NAND2_X1_3692_ (
  .A1({ S21859 }),
  .A2({ S25957[1183] }),
  .ZN({ S21860 })
);
NOR2_X1 #() 
NOR2_X1_933_ (
  .A1({ S21860 }),
  .A2({ S21850 }),
  .ZN({ S21861 })
);
NAND2_X1 #() 
NAND2_X1_3693_ (
  .A1({ S21622 }),
  .A2({ S21428 }),
  .ZN({ S21862 })
);
NAND3_X1 #() 
NAND3_X1_3936_ (
  .A1({ S21540 }),
  .A2({ S71 }),
  .A3({ S21401 }),
  .ZN({ S21863 })
);
NAND3_X1 #() 
NAND3_X1_3937_ (
  .A1({ S21400 }),
  .A2({ S25957[1179] }),
  .A3({ S79 }),
  .ZN({ S21864 })
);
OAI211_X1 #() 
OAI211_X1_1280_ (
  .A({ S25957[1180] }),
  .B({ S21863 }),
  .C1({ S21862 }),
  .C2({ S21864 }),
  .ZN({ S21865 })
);
NOR2_X1 #() 
NOR2_X1_934_ (
  .A1({ S21602 }),
  .A2({ S25957[1179] }),
  .ZN({ S21866 })
);
NOR2_X1 #() 
NOR2_X1_935_ (
  .A1({ S21866 }),
  .A2({ S25957[1180] }),
  .ZN({ S21867 })
);
NAND2_X1 #() 
NAND2_X1_3694_ (
  .A1({ S21554 }),
  .A2({ S21867 }),
  .ZN({ S21868 })
);
AOI21_X1 #() 
AOI21_X1_1991_ (
  .A({ S21444 }),
  .B1({ S21868 }),
  .B2({ S21865 }),
  .ZN({ S21869 })
);
NAND3_X1 #() 
NAND3_X1_3938_ (
  .A1({ S21601 }),
  .A2({ S21620 }),
  .A3({ S21398 }),
  .ZN({ S21870 })
);
NAND3_X1 #() 
NAND3_X1_3939_ (
  .A1({ S21532 }),
  .A2({ S21460 }),
  .A3({ S25957[1180] }),
  .ZN({ S21871 })
);
AND3_X1 #() 
AND3_X1_140_ (
  .A1({ S21870 }),
  .A2({ S21444 }),
  .A3({ S21871 }),
  .ZN({ S21872 })
);
OAI21_X1 #() 
OAI21_X1_1890_ (
  .A({ S25957[1182] }),
  .B1({ S21869 }),
  .B2({ S21872 }),
  .ZN({ S21873 })
);
AOI21_X1 #() 
AOI21_X1_1992_ (
  .A({ S25957[1179] }),
  .B1({ S21600 }),
  .B2({ S21622 }),
  .ZN({ S21874 })
);
OAI21_X1 #() 
OAI21_X1_1891_ (
  .A({ S25957[1180] }),
  .B1({ S21769 }),
  .B2({ S21874 }),
  .ZN({ S21875 })
);
NAND3_X1 #() 
NAND3_X1_3940_ (
  .A1({ S21622 }),
  .A2({ S25957[1179] }),
  .A3({ S79 }),
  .ZN({ S21876 })
);
OAI211_X1 #() 
OAI211_X1_1281_ (
  .A({ S21876 }),
  .B({ S21398 }),
  .C1({ S21659 }),
  .C2({ S21633 }),
  .ZN({ S21877 })
);
NAND3_X1 #() 
NAND3_X1_3941_ (
  .A1({ S21875 }),
  .A2({ S21877 }),
  .A3({ S21444 }),
  .ZN({ S21878 })
);
NAND3_X1 #() 
NAND3_X1_3942_ (
  .A1({ S21541 }),
  .A2({ S21635 }),
  .A3({ S21398 }),
  .ZN({ S21879 })
);
NAND2_X1 #() 
NAND2_X1_3695_ (
  .A1({ S21751 }),
  .A2({ S21627 }),
  .ZN({ S21880 })
);
NAND2_X1 #() 
NAND2_X1_3696_ (
  .A1({ S21880 }),
  .A2({ S21879 }),
  .ZN({ S21881 })
);
AOI21_X1 #() 
AOI21_X1_1993_ (
  .A({ S25957[1182] }),
  .B1({ S21881 }),
  .B2({ S25957[1181] }),
  .ZN({ S21882 })
);
NAND2_X1 #() 
NAND2_X1_3697_ (
  .A1({ S21882 }),
  .A2({ S21878 }),
  .ZN({ S21883 })
);
AOI21_X1 #() 
AOI21_X1_1994_ (
  .A({ S25957[1183] }),
  .B1({ S21883 }),
  .B2({ S21873 }),
  .ZN({ S21884 })
);
OAI21_X1 #() 
OAI21_X1_1892_ (
  .A({ S21838 }),
  .B1({ S21884 }),
  .B2({ S21861 }),
  .ZN({ S21885 })
);
NAND2_X1 #() 
NAND2_X1_3698_ (
  .A1({ S21401 }),
  .A2({ S25957[1178] }),
  .ZN({ S21886 })
);
OAI21_X1 #() 
OAI21_X1_1893_ (
  .A({ S21708 }),
  .B1({ S71 }),
  .B2({ S21886 }),
  .ZN({ S21887 })
);
NAND2_X1 #() 
NAND2_X1_3699_ (
  .A1({ S21887 }),
  .A2({ S25957[1180] }),
  .ZN({ S21888 })
);
AOI21_X1 #() 
AOI21_X1_1995_ (
  .A({ S21444 }),
  .B1({ S21888 }),
  .B2({ S21846 }),
  .ZN({ S21889 })
);
NAND2_X1 #() 
NAND2_X1_3700_ (
  .A1({ S21841 }),
  .A2({ S21444 }),
  .ZN({ S21890 })
);
OAI21_X1 #() 
OAI21_X1_1894_ (
  .A({ S25957[1182] }),
  .B1({ S21890 }),
  .B2({ S21840 }),
  .ZN({ S21891 })
);
OAI211_X1 #() 
OAI211_X1_1282_ (
  .A({ S21859 }),
  .B({ S25957[1183] }),
  .C1({ S21889 }),
  .C2({ S21891 }),
  .ZN({ S21892 })
);
NAND3_X1 #() 
NAND3_X1_3943_ (
  .A1({ S21434 }),
  .A2({ S25957[1179] }),
  .A3({ S21465 }),
  .ZN({ S21893 })
);
NAND3_X1 #() 
NAND3_X1_3944_ (
  .A1({ S21893 }),
  .A2({ S25957[1180] }),
  .A3({ S21546 }),
  .ZN({ S21894 })
);
AOI21_X1 #() 
AOI21_X1_1996_ (
  .A({ S71 }),
  .B1({ S21522 }),
  .B2({ S21531 }),
  .ZN({ S21895 })
);
OAI21_X1 #() 
OAI21_X1_1895_ (
  .A({ S21398 }),
  .B1({ S21895 }),
  .B2({ S21866 }),
  .ZN({ S21896 })
);
NAND3_X1 #() 
NAND3_X1_3945_ (
  .A1({ S21896 }),
  .A2({ S25957[1181] }),
  .A3({ S21894 }),
  .ZN({ S21897 })
);
NAND3_X1 #() 
NAND3_X1_3946_ (
  .A1({ S21870 }),
  .A2({ S21444 }),
  .A3({ S21871 }),
  .ZN({ S21898 })
);
NAND2_X1 #() 
NAND2_X1_3701_ (
  .A1({ S21897 }),
  .A2({ S21898 }),
  .ZN({ S21899 })
);
AOI22_X1 #() 
AOI22_X1_420_ (
  .A1({ S21899 }),
  .A2({ S25957[1182] }),
  .B1({ S21882 }),
  .B2({ S21878 }),
  .ZN({ S21900 })
);
OAI211_X1 #() 
OAI211_X1_1283_ (
  .A({ S25957[1248] }),
  .B({ S21892 }),
  .C1({ S21900 }),
  .C2({ S25957[1183] }),
  .ZN({ S21901 })
);
NAND3_X1 #() 
NAND3_X1_3947_ (
  .A1({ S21885 }),
  .A2({ S21837 }),
  .A3({ S21901 }),
  .ZN({ S21902 })
);
OAI211_X1 #() 
OAI211_X1_1284_ (
  .A({ S21838 }),
  .B({ S21892 }),
  .C1({ S21900 }),
  .C2({ S25957[1183] }),
  .ZN({ S21903 })
);
OAI21_X1 #() 
OAI21_X1_1896_ (
  .A({ S25957[1248] }),
  .B1({ S21884 }),
  .B2({ S21861 }),
  .ZN({ S21904 })
);
NAND3_X1 #() 
NAND3_X1_3948_ (
  .A1({ S21904 }),
  .A2({ S25957[1216] }),
  .A3({ S21903 }),
  .ZN({ S21905 })
);
AOI21_X1 #() 
AOI21_X1_1997_ (
  .A({ S11550 }),
  .B1({ S21902 }),
  .B2({ S21905 }),
  .ZN({ S21906 })
);
NAND3_X1 #() 
NAND3_X1_3949_ (
  .A1({ S21885 }),
  .A2({ S25957[1216] }),
  .A3({ S21901 }),
  .ZN({ S21907 })
);
NAND3_X1 #() 
NAND3_X1_3950_ (
  .A1({ S21904 }),
  .A2({ S21837 }),
  .A3({ S21903 }),
  .ZN({ S21908 })
);
AOI21_X1 #() 
AOI21_X1_1998_ (
  .A({ S25956[0] }),
  .B1({ S21907 }),
  .B2({ S21908 }),
  .ZN({ S21909 })
);
NOR2_X1 #() 
NOR2_X1_936_ (
  .A1({ S21906 }),
  .A2({ S21909 }),
  .ZN({ S25957[1024] })
);
NAND2_X1 #() 
NAND2_X1_3702_ (
  .A1({ S19480 }),
  .A2({ S19481 }),
  .ZN({ S25957[1217] })
);
INV_X1 #() 
INV_X1_1223_ (
  .A({ S25957[1217] }),
  .ZN({ S21910 })
);
NAND2_X1 #() 
NAND2_X1_3703_ (
  .A1({ S19473 }),
  .A2({ S19470 }),
  .ZN({ S25957[1249] })
);
INV_X1 #() 
INV_X1_1224_ (
  .A({ S25957[1249] }),
  .ZN({ S21911 })
);
NOR2_X1 #() 
NOR2_X1_937_ (
  .A1({ S21634 }),
  .A2({ S21615 }),
  .ZN({ S21912 })
);
OAI21_X1 #() 
OAI21_X1_1897_ (
  .A({ S25957[1180] }),
  .B1({ S21845 }),
  .B2({ S25957[1176] }),
  .ZN({ S21913 })
);
INV_X1 #() 
INV_X1_1225_ (
  .A({ S21412 }),
  .ZN({ S21914 })
);
NAND3_X1 #() 
NAND3_X1_3951_ (
  .A1({ S21540 }),
  .A2({ S25957[1179] }),
  .A3({ S21394 }),
  .ZN({ S21915 })
);
OAI211_X1 #() 
OAI211_X1_1285_ (
  .A({ S21398 }),
  .B({ S21915 }),
  .C1({ S21914 }),
  .C2({ S21795 }),
  .ZN({ S21916 })
);
OAI211_X1 #() 
OAI211_X1_1286_ (
  .A({ S21444 }),
  .B({ S21916 }),
  .C1({ S21912 }),
  .C2({ S21913 }),
  .ZN({ S21917 })
);
NOR2_X1 #() 
NOR2_X1_938_ (
  .A1({ S21862 }),
  .A2({ S21864 }),
  .ZN({ S21918 })
);
NAND2_X1 #() 
NAND2_X1_3704_ (
  .A1({ S21480 }),
  .A2({ S71 }),
  .ZN({ S21919 })
);
NAND3_X1 #() 
NAND3_X1_3952_ (
  .A1({ S21919 }),
  .A2({ S21603 }),
  .A3({ S25957[1180] }),
  .ZN({ S21920 })
);
NAND2_X1 #() 
NAND2_X1_3705_ (
  .A1({ S21522 }),
  .A2({ S71 }),
  .ZN({ S21921 })
);
NAND2_X1 #() 
NAND2_X1_3706_ (
  .A1({ S21921 }),
  .A2({ S21398 }),
  .ZN({ S21922 })
);
OAI211_X1 #() 
OAI211_X1_1287_ (
  .A({ S21920 }),
  .B({ S25957[1181] }),
  .C1({ S21918 }),
  .C2({ S21922 }),
  .ZN({ S21923 })
);
AOI21_X1 #() 
AOI21_X1_1999_ (
  .A({ S21433 }),
  .B1({ S21917 }),
  .B2({ S21923 }),
  .ZN({ S21924 })
);
OAI21_X1 #() 
OAI21_X1_1898_ (
  .A({ S21469 }),
  .B1({ S21780 }),
  .B2({ S71 }),
  .ZN({ S21925 })
);
AOI21_X1 #() 
AOI21_X1_2000_ (
  .A({ S25957[1180] }),
  .B1({ S21531 }),
  .B2({ S25957[1179] }),
  .ZN({ S21926 })
);
AOI21_X1 #() 
AOI21_X1_2001_ (
  .A({ S21444 }),
  .B1({ S21791 }),
  .B2({ S21926 }),
  .ZN({ S21927 })
);
INV_X1 #() 
INV_X1_1226_ (
  .A({ S21485 }),
  .ZN({ S21928 })
);
NAND3_X1 #() 
NAND3_X1_3953_ (
  .A1({ S21928 }),
  .A2({ S21398 }),
  .A3({ S21685 }),
  .ZN({ S21929 })
);
OAI211_X1 #() 
OAI211_X1_1288_ (
  .A({ S21472 }),
  .B({ S71 }),
  .C1({ S25957[1178] }),
  .C2({ S21401 }),
  .ZN({ S21930 })
);
AOI21_X1 #() 
AOI21_X1_2002_ (
  .A({ S25957[1181] }),
  .B1({ S21548 }),
  .B2({ S21930 }),
  .ZN({ S21931 })
);
AOI22_X1 #() 
AOI22_X1_421_ (
  .A1({ S21929 }),
  .A2({ S21931 }),
  .B1({ S21925 }),
  .B2({ S21927 }),
  .ZN({ S21932 })
);
OAI21_X1 #() 
OAI21_X1_1899_ (
  .A({ S25957[1183] }),
  .B1({ S21932 }),
  .B2({ S25957[1182] }),
  .ZN({ S21933 })
);
NAND3_X1 #() 
NAND3_X1_3954_ (
  .A1({ S21453 }),
  .A2({ S21535 }),
  .A3({ S21493 }),
  .ZN({ S21934 })
);
AOI22_X1 #() 
AOI22_X1_422_ (
  .A1({ S21934 }),
  .A2({ S21439 }),
  .B1({ S21777 }),
  .B2({ S25957[1179] }),
  .ZN({ S21935 })
);
NAND3_X1 #() 
NAND3_X1_3955_ (
  .A1({ S21412 }),
  .A2({ S21455 }),
  .A3({ S21423 }),
  .ZN({ S21936 })
);
NAND2_X1 #() 
NAND2_X1_3707_ (
  .A1({ S21936 }),
  .A2({ S21398 }),
  .ZN({ S21937 })
);
OAI211_X1 #() 
OAI211_X1_1289_ (
  .A({ S21937 }),
  .B({ S25957[1181] }),
  .C1({ S21935 }),
  .C2({ S21398 }),
  .ZN({ S21938 })
);
NAND4_X1 #() 
NAND4_X1_434_ (
  .A1({ S21401 }),
  .A2({ S21416 }),
  .A3({ S25957[1179] }),
  .A4({ S25957[1178] }),
  .ZN({ S21939 })
);
AOI21_X1 #() 
AOI21_X1_2003_ (
  .A({ S25957[1180] }),
  .B1({ S21566 }),
  .B2({ S21939 }),
  .ZN({ S21940 })
);
AOI21_X1 #() 
AOI21_X1_2004_ (
  .A({ S21602 }),
  .B1({ S21406 }),
  .B2({ S21423 }),
  .ZN({ S21941 })
);
NOR2_X1 #() 
NOR2_X1_939_ (
  .A1({ S21941 }),
  .A2({ S21429 }),
  .ZN({ S21942 })
);
NAND2_X1 #() 
NAND2_X1_3708_ (
  .A1({ S21622 }),
  .A2({ S25957[1180] }),
  .ZN({ S21943 })
);
OAI21_X1 #() 
OAI21_X1_1900_ (
  .A({ S21444 }),
  .B1({ S21942 }),
  .B2({ S21943 }),
  .ZN({ S21944 })
);
OAI211_X1 #() 
OAI211_X1_1290_ (
  .A({ S21938 }),
  .B({ S25957[1182] }),
  .C1({ S21944 }),
  .C2({ S21940 }),
  .ZN({ S21945 })
);
NOR2_X1 #() 
NOR2_X1_940_ (
  .A1({ S21526 }),
  .A2({ S21668 }),
  .ZN({ S21946 })
);
AOI21_X1 #() 
AOI21_X1_2005_ (
  .A({ S21448 }),
  .B1({ S21476 }),
  .B2({ S21473 }),
  .ZN({ S21947 })
);
OAI21_X1 #() 
OAI21_X1_1901_ (
  .A({ S21444 }),
  .B1({ S21947 }),
  .B2({ S21946 }),
  .ZN({ S21948 })
);
AOI21_X1 #() 
AOI21_X1_2006_ (
  .A({ S21398 }),
  .B1({ S21762 }),
  .B2({ S21661 }),
  .ZN({ S21949 })
);
INV_X1 #() 
INV_X1_1227_ (
  .A({ S21949 }),
  .ZN({ S21950 })
);
NAND3_X1 #() 
NAND3_X1_3956_ (
  .A1({ S21518 }),
  .A2({ S21950 }),
  .A3({ S25957[1181] }),
  .ZN({ S21951 })
);
NAND3_X1 #() 
NAND3_X1_3957_ (
  .A1({ S21951 }),
  .A2({ S21948 }),
  .A3({ S21433 }),
  .ZN({ S21952 })
);
NAND3_X1 #() 
NAND3_X1_3958_ (
  .A1({ S21945 }),
  .A2({ S21952 }),
  .A3({ S21395 }),
  .ZN({ S21953 })
);
OAI211_X1 #() 
OAI211_X1_1291_ (
  .A({ S21953 }),
  .B({ S21911 }),
  .C1({ S21933 }),
  .C2({ S21924 }),
  .ZN({ S21954 })
);
NAND2_X1 #() 
NAND2_X1_3709_ (
  .A1({ S21925 }),
  .A2({ S21927 }),
  .ZN({ S21955 })
);
NAND2_X1 #() 
NAND2_X1_3710_ (
  .A1({ S21929 }),
  .A2({ S21931 }),
  .ZN({ S21956 })
);
AOI21_X1 #() 
AOI21_X1_2007_ (
  .A({ S25957[1182] }),
  .B1({ S21956 }),
  .B2({ S21955 }),
  .ZN({ S21957 })
);
OAI21_X1 #() 
OAI21_X1_1902_ (
  .A({ S25957[1183] }),
  .B1({ S21957 }),
  .B2({ S21924 }),
  .ZN({ S21958 })
);
AND2_X1 #() 
AND2_X1_229_ (
  .A1({ S21777 }),
  .A2({ S25957[1179] }),
  .ZN({ S21959 })
);
NAND3_X1 #() 
NAND3_X1_3959_ (
  .A1({ S21587 }),
  .A2({ S21423 }),
  .A3({ S21412 }),
  .ZN({ S21960 })
);
OAI21_X1 #() 
OAI21_X1_1903_ (
  .A({ S25957[1180] }),
  .B1({ S21659 }),
  .B2({ S21664 }),
  .ZN({ S21961 })
);
OAI211_X1 #() 
OAI211_X1_1292_ (
  .A({ S25957[1181] }),
  .B({ S21960 }),
  .C1({ S21961 }),
  .C2({ S21959 }),
  .ZN({ S21962 })
);
OAI21_X1 #() 
OAI21_X1_1904_ (
  .A({ S21428 }),
  .B1({ S21452 }),
  .B2({ S21455 }),
  .ZN({ S21963 })
);
AOI21_X1 #() 
AOI21_X1_2008_ (
  .A({ S21943 }),
  .B1({ S21963 }),
  .B2({ S21453 }),
  .ZN({ S21964 })
);
OAI21_X1 #() 
OAI21_X1_1905_ (
  .A({ S21444 }),
  .B1({ S21964 }),
  .B2({ S21940 }),
  .ZN({ S21965 })
);
AOI21_X1 #() 
AOI21_X1_2009_ (
  .A({ S21433 }),
  .B1({ S21965 }),
  .B2({ S21962 }),
  .ZN({ S21966 })
);
OAI21_X1 #() 
OAI21_X1_1906_ (
  .A({ S25957[1181] }),
  .B1({ S21482 }),
  .B2({ S21949 }),
  .ZN({ S21967 })
);
NAND4_X1 #() 
NAND4_X1_435_ (
  .A1({ S21456 }),
  .A2({ S21805 }),
  .A3({ S25957[1180] }),
  .A4({ S21455 }),
  .ZN({ S21968 })
);
OAI21_X1 #() 
OAI21_X1_1907_ (
  .A({ S21449 }),
  .B1({ S21481 }),
  .B2({ S25957[1179] }),
  .ZN({ S21969 })
);
NAND3_X1 #() 
NAND3_X1_3960_ (
  .A1({ S21969 }),
  .A2({ S21444 }),
  .A3({ S21968 }),
  .ZN({ S21970 })
);
AOI21_X1 #() 
AOI21_X1_2010_ (
  .A({ S25957[1182] }),
  .B1({ S21970 }),
  .B2({ S21967 }),
  .ZN({ S21971 })
);
OAI21_X1 #() 
OAI21_X1_1908_ (
  .A({ S21395 }),
  .B1({ S21966 }),
  .B2({ S21971 }),
  .ZN({ S21972 })
);
NAND3_X1 #() 
NAND3_X1_3961_ (
  .A1({ S21958 }),
  .A2({ S21972 }),
  .A3({ S25957[1249] }),
  .ZN({ S21973 })
);
NAND3_X1 #() 
NAND3_X1_3962_ (
  .A1({ S21973 }),
  .A2({ S21954 }),
  .A3({ S21910 }),
  .ZN({ S21974 })
);
OAI211_X1 #() 
OAI211_X1_1293_ (
  .A({ S21953 }),
  .B({ S25957[1249] }),
  .C1({ S21933 }),
  .C2({ S21924 }),
  .ZN({ S21975 })
);
NAND3_X1 #() 
NAND3_X1_3963_ (
  .A1({ S21958 }),
  .A2({ S21972 }),
  .A3({ S21911 }),
  .ZN({ S21976 })
);
NAND3_X1 #() 
NAND3_X1_3964_ (
  .A1({ S21976 }),
  .A2({ S21975 }),
  .A3({ S25957[1217] }),
  .ZN({ S21977 })
);
AOI21_X1 #() 
AOI21_X1_2011_ (
  .A({ S11539 }),
  .B1({ S21974 }),
  .B2({ S21977 }),
  .ZN({ S21978 })
);
NAND3_X1 #() 
NAND3_X1_3965_ (
  .A1({ S21973 }),
  .A2({ S21954 }),
  .A3({ S25957[1217] }),
  .ZN({ S21979 })
);
NAND3_X1 #() 
NAND3_X1_3966_ (
  .A1({ S21976 }),
  .A2({ S21975 }),
  .A3({ S21910 }),
  .ZN({ S21980 })
);
AOI21_X1 #() 
AOI21_X1_2012_ (
  .A({ S25956[1] }),
  .B1({ S21979 }),
  .B2({ S21980 }),
  .ZN({ S21981 })
);
NOR2_X1 #() 
NOR2_X1_941_ (
  .A1({ S21978 }),
  .A2({ S21981 }),
  .ZN({ S25957[1025] })
);
INV_X1 #() 
INV_X1_1228_ (
  .A({ S19534 }),
  .ZN({ S25957[1218] })
);
INV_X1 #() 
INV_X1_1229_ (
  .A({ S19530 }),
  .ZN({ S25957[1250] })
);
OAI21_X1 #() 
OAI21_X1_1909_ (
  .A({ S71 }),
  .B1({ S25957[1178] }),
  .B2({ S21399 }),
  .ZN({ S21982 })
);
OAI21_X1 #() 
OAI21_X1_1910_ (
  .A({ S21398 }),
  .B1({ S21982 }),
  .B2({ S21408 }),
  .ZN({ S21983 })
);
NAND4_X1 #() 
NAND4_X1_436_ (
  .A1({ S25957[1180] }),
  .A2({ S21400 }),
  .A3({ S25957[1179] }),
  .A4({ S21416 }),
  .ZN({ S21984 })
);
OAI21_X1 #() 
OAI21_X1_1911_ (
  .A({ S21984 }),
  .B1({ S21436 }),
  .B2({ S21983 }),
  .ZN({ S21985 })
);
NAND2_X1 #() 
NAND2_X1_3711_ (
  .A1({ S21985 }),
  .A2({ S25957[1181] }),
  .ZN({ S21986 })
);
NAND3_X1 #() 
NAND3_X1_3967_ (
  .A1({ S21439 }),
  .A2({ S25957[1179] }),
  .A3({ S25957[1177] }),
  .ZN({ S21987 })
);
AND3_X1 #() 
AND3_X1_141_ (
  .A1({ S21839 }),
  .A2({ S21987 }),
  .A3({ S21398 }),
  .ZN({ S21988 })
);
NAND2_X1 #() 
NAND2_X1_3712_ (
  .A1({ S21790 }),
  .A2({ S71 }),
  .ZN({ S21989 })
);
OAI211_X1 #() 
OAI211_X1_1294_ (
  .A({ S21423 }),
  .B({ S25957[1179] }),
  .C1({ S21401 }),
  .C2({ S25957[1178] }),
  .ZN({ S21990 })
);
AOI21_X1 #() 
AOI21_X1_2013_ (
  .A({ S21398 }),
  .B1({ S21989 }),
  .B2({ S21990 }),
  .ZN({ S21991 })
);
OAI21_X1 #() 
OAI21_X1_1912_ (
  .A({ S21444 }),
  .B1({ S21988 }),
  .B2({ S21991 }),
  .ZN({ S21992 })
);
NOR2_X1 #() 
NOR2_X1_942_ (
  .A1({ S21433 }),
  .A2({ S21796 }),
  .ZN({ S21993 })
);
NAND3_X1 #() 
NAND3_X1_3968_ (
  .A1({ S21992 }),
  .A2({ S21986 }),
  .A3({ S21993 }),
  .ZN({ S21994 })
);
OAI21_X1 #() 
OAI21_X1_1913_ (
  .A({ S21398 }),
  .B1({ S21845 }),
  .B2({ S21592 }),
  .ZN({ S21995 })
);
NAND3_X1 #() 
NAND3_X1_3969_ (
  .A1({ S21681 }),
  .A2({ S25957[1180] }),
  .A3({ S21987 }),
  .ZN({ S21996 })
);
OAI211_X1 #() 
OAI211_X1_1295_ (
  .A({ S21996 }),
  .B({ S21444 }),
  .C1({ S21995 }),
  .C2({ S21895 }),
  .ZN({ S21997 })
);
NAND3_X1 #() 
NAND3_X1_3970_ (
  .A1({ S21412 }),
  .A2({ S25957[1179] }),
  .A3({ S21423 }),
  .ZN({ S21998 })
);
NAND3_X1 #() 
NAND3_X1_3971_ (
  .A1({ S21761 }),
  .A2({ S21998 }),
  .A3({ S25957[1180] }),
  .ZN({ S21999 })
);
NAND3_X1 #() 
NAND3_X1_3972_ (
  .A1({ S21622 }),
  .A2({ S21490 }),
  .A3({ S25957[1179] }),
  .ZN({ S22000 })
);
AOI21_X1 #() 
AOI21_X1_2014_ (
  .A({ S25957[1180] }),
  .B1({ S21429 }),
  .B2({ S21602 }),
  .ZN({ S22001 })
);
AOI21_X1 #() 
AOI21_X1_2015_ (
  .A({ S21444 }),
  .B1({ S22001 }),
  .B2({ S22000 }),
  .ZN({ S22002 })
);
AOI21_X1 #() 
AOI21_X1_2016_ (
  .A({ S25957[1182] }),
  .B1({ S22002 }),
  .B2({ S21999 }),
  .ZN({ S22003 })
);
AOI21_X1 #() 
AOI21_X1_2017_ (
  .A({ S25957[1183] }),
  .B1({ S22003 }),
  .B2({ S21997 }),
  .ZN({ S22004 })
);
NAND2_X1 #() 
NAND2_X1_3713_ (
  .A1({ S22004 }),
  .A2({ S21994 }),
  .ZN({ S22005 })
);
NOR2_X1 #() 
NOR2_X1_943_ (
  .A1({ S21422 }),
  .A2({ S21491 }),
  .ZN({ S22006 })
);
NAND4_X1 #() 
NAND4_X1_437_ (
  .A1({ S21989 }),
  .A2({ S21479 }),
  .A3({ S25957[1180] }),
  .A4({ S21698 }),
  .ZN({ S22007 })
);
NAND3_X1 #() 
NAND3_X1_3973_ (
  .A1({ S21446 }),
  .A2({ S25957[1179] }),
  .A3({ S21886 }),
  .ZN({ S22008 })
);
NAND3_X1 #() 
NAND3_X1_3974_ (
  .A1({ S22008 }),
  .A2({ S21398 }),
  .A3({ S21845 }),
  .ZN({ S22009 })
);
NAND3_X1 #() 
NAND3_X1_3975_ (
  .A1({ S22009 }),
  .A2({ S22007 }),
  .A3({ S25957[1181] }),
  .ZN({ S22010 })
);
NAND2_X1 #() 
NAND2_X1_3714_ (
  .A1({ S21594 }),
  .A2({ S25957[1180] }),
  .ZN({ S22011 })
);
NOR2_X1 #() 
NOR2_X1_944_ (
  .A1({ S21447 }),
  .A2({ S71 }),
  .ZN({ S22012 })
);
OAI21_X1 #() 
OAI21_X1_1914_ (
  .A({ S21444 }),
  .B1({ S22012 }),
  .B2({ S22011 }),
  .ZN({ S22013 })
);
OAI211_X1 #() 
OAI211_X1_1296_ (
  .A({ S25957[1182] }),
  .B({ S22010 }),
  .C1({ S22013 }),
  .C2({ S22006 }),
  .ZN({ S22014 })
);
NAND3_X1 #() 
NAND3_X1_3976_ (
  .A1({ S21400 }),
  .A2({ S25957[1179] }),
  .A3({ S25957[1176] }),
  .ZN({ S22015 })
);
OAI211_X1 #() 
OAI211_X1_1297_ (
  .A({ S25957[1180] }),
  .B({ S22015 }),
  .C1({ S21481 }),
  .C2({ S25957[1179] }),
  .ZN({ S22016 })
);
OAI211_X1 #() 
OAI211_X1_1298_ (
  .A({ S25957[1179] }),
  .B({ S21401 }),
  .C1({ S21416 }),
  .C2({ S21411 }),
  .ZN({ S22017 })
);
NAND3_X1 #() 
NAND3_X1_3977_ (
  .A1({ S21690 }),
  .A2({ S22017 }),
  .A3({ S21398 }),
  .ZN({ S22018 })
);
NAND3_X1 #() 
NAND3_X1_3978_ (
  .A1({ S22016 }),
  .A2({ S25957[1181] }),
  .A3({ S22018 }),
  .ZN({ S22019 })
);
NAND3_X1 #() 
NAND3_X1_3979_ (
  .A1({ S21987 }),
  .A2({ S25957[1180] }),
  .A3({ S21982 }),
  .ZN({ S22020 })
);
OAI211_X1 #() 
OAI211_X1_1299_ (
  .A({ S22020 }),
  .B({ S21444 }),
  .C1({ S25957[1180] }),
  .C2({ S21536 }),
  .ZN({ S22021 })
);
NAND3_X1 #() 
NAND3_X1_3980_ (
  .A1({ S22019 }),
  .A2({ S21433 }),
  .A3({ S22021 }),
  .ZN({ S22022 })
);
NAND3_X1 #() 
NAND3_X1_3981_ (
  .A1({ S22014 }),
  .A2({ S25957[1183] }),
  .A3({ S22022 }),
  .ZN({ S22023 })
);
NAND3_X1 #() 
NAND3_X1_3982_ (
  .A1({ S22023 }),
  .A2({ S22005 }),
  .A3({ S25957[1250] }),
  .ZN({ S22024 })
);
NAND2_X1 #() 
NAND2_X1_3715_ (
  .A1({ S22023 }),
  .A2({ S22005 }),
  .ZN({ S22025 })
);
NAND2_X1 #() 
NAND2_X1_3716_ (
  .A1({ S22025 }),
  .A2({ S19530 }),
  .ZN({ S22026 })
);
NAND3_X1 #() 
NAND3_X1_3983_ (
  .A1({ S22026 }),
  .A2({ S25957[1218] }),
  .A3({ S22024 }),
  .ZN({ S22027 })
);
NAND3_X1 #() 
NAND3_X1_3984_ (
  .A1({ S22023 }),
  .A2({ S22005 }),
  .A3({ S19530 }),
  .ZN({ S22028 })
);
NAND2_X1 #() 
NAND2_X1_3717_ (
  .A1({ S22025 }),
  .A2({ S25957[1250] }),
  .ZN({ S22029 })
);
NAND3_X1 #() 
NAND3_X1_3985_ (
  .A1({ S22029 }),
  .A2({ S19534 }),
  .A3({ S22028 }),
  .ZN({ S22030 })
);
NAND3_X1 #() 
NAND3_X1_3986_ (
  .A1({ S22027 }),
  .A2({ S22030 }),
  .A3({ S11642 }),
  .ZN({ S22031 })
);
NAND3_X1 #() 
NAND3_X1_3987_ (
  .A1({ S22029 }),
  .A2({ S25957[1218] }),
  .A3({ S22028 }),
  .ZN({ S22032 })
);
NAND3_X1 #() 
NAND3_X1_3988_ (
  .A1({ S22026 }),
  .A2({ S19534 }),
  .A3({ S22024 }),
  .ZN({ S22033 })
);
NAND3_X1 #() 
NAND3_X1_3989_ (
  .A1({ S22032 }),
  .A2({ S22033 }),
  .A3({ S25956[2] }),
  .ZN({ S22034 })
);
NAND2_X1 #() 
NAND2_X1_3718_ (
  .A1({ S22031 }),
  .A2({ S22034 }),
  .ZN({ S25957[1026] })
);
NAND2_X1 #() 
NAND2_X1_3719_ (
  .A1({ S25957[1168] }),
  .A2({ S25957[1169] }),
  .ZN({ S22035 })
);
INV_X1 #() 
INV_X1_1230_ (
  .A({ S22035 }),
  .ZN({ S81 })
);
NAND4_X1 #() 
NAND4_X1_438_ (
  .A1({ S10379 }),
  .A2({ S10417 }),
  .A3({ S10915 }),
  .A4({ S10948 }),
  .ZN({ S82 })
);
NAND2_X1 #() 
NAND2_X1_3720_ (
  .A1({ S25957[1170] }),
  .A2({ S20616 }),
  .ZN({ S22036 })
);
NAND4_X1 #() 
NAND4_X1_439_ (
  .A1({ S20614 }),
  .A2({ S20615 }),
  .A3({ S10915 }),
  .A4({ S10948 }),
  .ZN({ S22037 })
);
OAI211_X1 #() 
OAI211_X1_1300_ (
  .A({ S22036 }),
  .B({ S25957[1171] }),
  .C1({ S22037 }),
  .C2({ S25957[1170] }),
  .ZN({ S22038 })
);
INV_X1 #() 
INV_X1_1231_ (
  .A({ S22038 }),
  .ZN({ S22039 })
);
NOR2_X1 #() 
NOR2_X1_945_ (
  .A1({ S25957[1170] }),
  .A2({ S25957[1168] }),
  .ZN({ S22040 })
);
NOR2_X1 #() 
NOR2_X1_946_ (
  .A1({ S22040 }),
  .A2({ S25957[1171] }),
  .ZN({ S22041 })
);
AOI21_X1 #() 
AOI21_X1_2018_ (
  .A({ S22039 }),
  .B1({ S25957[1169] }),
  .B2({ S22041 }),
  .ZN({ S22042 })
);
NOR2_X1 #() 
NOR2_X1_947_ (
  .A1({ S22035 }),
  .A2({ S25957[1170] }),
  .ZN({ S22043 })
);
NAND3_X1 #() 
NAND3_X1_3990_ (
  .A1({ S20676 }),
  .A2({ S25957[1170] }),
  .A3({ S20616 }),
  .ZN({ S22044 })
);
NAND2_X1 #() 
NAND2_X1_3721_ (
  .A1({ S22044 }),
  .A2({ S50 }),
  .ZN({ S22045 })
);
AOI22_X1 #() 
AOI22_X1_423_ (
  .A1({ S20614 }),
  .A2({ S20615 }),
  .B1({ S10915 }),
  .B2({ S10948 }),
  .ZN({ S22046 })
);
NAND2_X1 #() 
NAND2_X1_3722_ (
  .A1({ S22046 }),
  .A2({ S25957[1170] }),
  .ZN({ S22047 })
);
NAND2_X1 #() 
NAND2_X1_3723_ (
  .A1({ S22047 }),
  .A2({ S22037 }),
  .ZN({ S22048 })
);
OAI221_X1 #() 
OAI221_X1_110_ (
  .A({ S9119 }),
  .B1({ S22045 }),
  .B2({ S22043 }),
  .C1({ S50 }),
  .C2({ S22048 }),
  .ZN({ S22049 })
);
OAI211_X1 #() 
OAI211_X1_1301_ (
  .A({ S22049 }),
  .B({ S25957[1173] }),
  .C1({ S22042 }),
  .C2({ S9119 }),
  .ZN({ S22050 })
);
INV_X1 #() 
INV_X1_1232_ (
  .A({ S25957[1173] }),
  .ZN({ S22051 })
);
NAND2_X1 #() 
NAND2_X1_3724_ (
  .A1({ S20616 }),
  .A2({ S25957[1169] }),
  .ZN({ S22052 })
);
NAND2_X1 #() 
NAND2_X1_3725_ (
  .A1({ S22052 }),
  .A2({ S50 }),
  .ZN({ S22053 })
);
INV_X1 #() 
INV_X1_1233_ (
  .A({ S22053 }),
  .ZN({ S22054 })
);
NAND4_X1 #() 
NAND4_X1_440_ (
  .A1({ S11476 }),
  .A2({ S11518 }),
  .A3({ S10915 }),
  .A4({ S10948 }),
  .ZN({ S22055 })
);
AOI21_X1 #() 
AOI21_X1_2019_ (
  .A({ S50 }),
  .B1({ S22052 }),
  .B2({ S22055 }),
  .ZN({ S22056 })
);
OAI21_X1 #() 
OAI21_X1_1915_ (
  .A({ S25957[1172] }),
  .B1({ S22054 }),
  .B2({ S22056 }),
  .ZN({ S22057 })
);
NAND2_X1 #() 
NAND2_X1_3726_ (
  .A1({ S82 }),
  .A2({ S20682 }),
  .ZN({ S22058 })
);
NAND2_X1 #() 
NAND2_X1_3727_ (
  .A1({ S22044 }),
  .A2({ S22058 }),
  .ZN({ S22059 })
);
INV_X1 #() 
INV_X1_1234_ (
  .A({ S22037 }),
  .ZN({ S22060 })
);
NAND2_X1 #() 
NAND2_X1_3728_ (
  .A1({ S22060 }),
  .A2({ S25957[1171] }),
  .ZN({ S22061 })
);
NAND3_X1 #() 
NAND3_X1_3991_ (
  .A1({ S22059 }),
  .A2({ S9119 }),
  .A3({ S22061 }),
  .ZN({ S22062 })
);
NAND3_X1 #() 
NAND3_X1_3992_ (
  .A1({ S22057 }),
  .A2({ S22062 }),
  .A3({ S22051 }),
  .ZN({ S22063 })
);
AND3_X1 #() 
AND3_X1_142_ (
  .A1({ S22050 }),
  .A2({ S25957[1174] }),
  .A3({ S22063 }),
  .ZN({ S22064 })
);
NAND2_X1 #() 
NAND2_X1_3729_ (
  .A1({ S25957[1170] }),
  .A2({ S25957[1168] }),
  .ZN({ S22065 })
);
NOR2_X1 #() 
NOR2_X1_948_ (
  .A1({ S20676 }),
  .A2({ S25957[1171] }),
  .ZN({ S22066 })
);
NAND2_X1 #() 
NAND2_X1_3730_ (
  .A1({ S22066 }),
  .A2({ S22065 }),
  .ZN({ S22067 })
);
NOR2_X1 #() 
NOR2_X1_949_ (
  .A1({ S20682 }),
  .A2({ S20616 }),
  .ZN({ S22068 })
);
OAI21_X1 #() 
OAI21_X1_1916_ (
  .A({ S25957[1171] }),
  .B1({ S22068 }),
  .B2({ S20676 }),
  .ZN({ S22069 })
);
AOI21_X1 #() 
AOI21_X1_2020_ (
  .A({ S9119 }),
  .B1({ S22069 }),
  .B2({ S22067 }),
  .ZN({ S22070 })
);
OAI21_X1 #() 
OAI21_X1_1917_ (
  .A({ S50 }),
  .B1({ S82 }),
  .B2({ S25957[1170] }),
  .ZN({ S22071 })
);
AOI21_X1 #() 
AOI21_X1_2021_ (
  .A({ S25957[1172] }),
  .B1({ S22071 }),
  .B2({ S22035 }),
  .ZN({ S22072 })
);
NOR3_X1 #() 
NOR3_X1_127_ (
  .A1({ S22070 }),
  .A2({ S22072 }),
  .A3({ S22051 }),
  .ZN({ S22073 })
);
NAND2_X1 #() 
NAND2_X1_3731_ (
  .A1({ S22036 }),
  .A2({ S50 }),
  .ZN({ S22074 })
);
INV_X1 #() 
INV_X1_1235_ (
  .A({ S22074 }),
  .ZN({ S22075 })
);
NAND2_X1 #() 
NAND2_X1_3732_ (
  .A1({ S25957[1170] }),
  .A2({ S25957[1169] }),
  .ZN({ S22076 })
);
NAND3_X1 #() 
NAND3_X1_3993_ (
  .A1({ S22076 }),
  .A2({ S25957[1168] }),
  .A3({ S22055 }),
  .ZN({ S22077 })
);
NAND2_X1 #() 
NAND2_X1_3733_ (
  .A1({ S22077 }),
  .A2({ S82 }),
  .ZN({ S22078 })
);
NAND2_X1 #() 
NAND2_X1_3734_ (
  .A1({ S22078 }),
  .A2({ S22075 }),
  .ZN({ S22079 })
);
INV_X1 #() 
INV_X1_1236_ (
  .A({ S22055 }),
  .ZN({ S22080 })
);
AOI21_X1 #() 
AOI21_X1_2022_ (
  .A({ S25957[1172] }),
  .B1({ S22080 }),
  .B2({ S25957[1171] }),
  .ZN({ S22081 })
);
AOI21_X1 #() 
AOI21_X1_2023_ (
  .A({ S20682 }),
  .B1({ S22052 }),
  .B2({ S22037 }),
  .ZN({ S22082 })
);
NAND2_X1 #() 
NAND2_X1_3735_ (
  .A1({ S22037 }),
  .A2({ S20682 }),
  .ZN({ S22083 })
);
NOR2_X1 #() 
NOR2_X1_950_ (
  .A1({ S22083 }),
  .A2({ S22046 }),
  .ZN({ S22084 })
);
OAI21_X1 #() 
OAI21_X1_1918_ (
  .A({ S25957[1171] }),
  .B1({ S22084 }),
  .B2({ S22082 }),
  .ZN({ S22085 })
);
NAND2_X1 #() 
NAND2_X1_3736_ (
  .A1({ S20682 }),
  .A2({ S25957[1168] }),
  .ZN({ S22086 })
);
NAND2_X1 #() 
NAND2_X1_3737_ (
  .A1({ S22086 }),
  .A2({ S50 }),
  .ZN({ S22087 })
);
INV_X1 #() 
INV_X1_1237_ (
  .A({ S22087 }),
  .ZN({ S22088 })
);
NAND2_X1 #() 
NAND2_X1_3738_ (
  .A1({ S22088 }),
  .A2({ S22076 }),
  .ZN({ S22089 })
);
AOI21_X1 #() 
AOI21_X1_2024_ (
  .A({ S9119 }),
  .B1({ S22085 }),
  .B2({ S22089 }),
  .ZN({ S22090 })
);
AOI21_X1 #() 
AOI21_X1_2025_ (
  .A({ S22090 }),
  .B1({ S22081 }),
  .B2({ S22079 }),
  .ZN({ S22091 })
);
AOI211_X1 #() 
AOI211_X1_62_ (
  .A({ S22073 }),
  .B({ S25957[1174] }),
  .C1({ S22091 }),
  .C2({ S22051 }),
  .ZN({ S22092 })
);
OAI21_X1 #() 
OAI21_X1_1919_ (
  .A({ S25957[1175] }),
  .B1({ S22092 }),
  .B2({ S22064 }),
  .ZN({ S22093 })
);
INV_X1 #() 
INV_X1_1238_ (
  .A({ S25957[1175] }),
  .ZN({ S22094 })
);
NAND2_X1 #() 
NAND2_X1_3739_ (
  .A1({ S20682 }),
  .A2({ S25957[1169] }),
  .ZN({ S22095 })
);
NAND2_X1 #() 
NAND2_X1_3740_ (
  .A1({ S22065 }),
  .A2({ S25957[1171] }),
  .ZN({ S22096 })
);
INV_X1 #() 
INV_X1_1239_ (
  .A({ S22096 }),
  .ZN({ S22097 })
);
NAND2_X1 #() 
NAND2_X1_3741_ (
  .A1({ S22097 }),
  .A2({ S22095 }),
  .ZN({ S22098 })
);
NAND2_X1 #() 
NAND2_X1_3742_ (
  .A1({ S22035 }),
  .A2({ S25957[1170] }),
  .ZN({ S22099 })
);
NAND2_X1 #() 
NAND2_X1_3743_ (
  .A1({ S22099 }),
  .A2({ S22083 }),
  .ZN({ S22100 })
);
AOI21_X1 #() 
AOI21_X1_2026_ (
  .A({ S25957[1172] }),
  .B1({ S22100 }),
  .B2({ S50 }),
  .ZN({ S22101 })
);
NOR2_X1 #() 
NOR2_X1_951_ (
  .A1({ S22046 }),
  .A2({ S25957[1170] }),
  .ZN({ S22102 })
);
NAND2_X1 #() 
NAND2_X1_3744_ (
  .A1({ S22102 }),
  .A2({ S22037 }),
  .ZN({ S22103 })
);
AOI21_X1 #() 
AOI21_X1_2027_ (
  .A({ S50 }),
  .B1({ S22103 }),
  .B2({ S22099 }),
  .ZN({ S22104 })
);
OAI21_X1 #() 
OAI21_X1_1920_ (
  .A({ S25957[1172] }),
  .B1({ S22082 }),
  .B2({ S22087 }),
  .ZN({ S22105 })
);
OAI21_X1 #() 
OAI21_X1_1921_ (
  .A({ S22051 }),
  .B1({ S22104 }),
  .B2({ S22105 }),
  .ZN({ S22106 })
);
AOI21_X1 #() 
AOI21_X1_2028_ (
  .A({ S22106 }),
  .B1({ S22101 }),
  .B2({ S22098 }),
  .ZN({ S22107 })
);
NOR2_X1 #() 
NOR2_X1_952_ (
  .A1({ S82 }),
  .A2({ S20682 }),
  .ZN({ S22108 })
);
NOR3_X1 #() 
NOR3_X1_128_ (
  .A1({ S22043 }),
  .A2({ S22108 }),
  .A3({ S50 }),
  .ZN({ S22109 })
);
NAND2_X1 #() 
NAND2_X1_3745_ (
  .A1({ S22047 }),
  .A2({ S50 }),
  .ZN({ S22110 })
);
OAI21_X1 #() 
OAI21_X1_1922_ (
  .A({ S25957[1172] }),
  .B1({ S22110 }),
  .B2({ S22040 }),
  .ZN({ S22111 })
);
AOI21_X1 #() 
AOI21_X1_2029_ (
  .A({ S50 }),
  .B1({ S20676 }),
  .B2({ S25957[1170] }),
  .ZN({ S22112 })
);
NAND2_X1 #() 
NAND2_X1_3746_ (
  .A1({ S22112 }),
  .A2({ S22083 }),
  .ZN({ S22113 })
);
NAND2_X1 #() 
NAND2_X1_3747_ (
  .A1({ S20676 }),
  .A2({ S25957[1170] }),
  .ZN({ S22114 })
);
NAND3_X1 #() 
NAND3_X1_3994_ (
  .A1({ S22114 }),
  .A2({ S22036 }),
  .A3({ S50 }),
  .ZN({ S22115 })
);
NAND3_X1 #() 
NAND3_X1_3995_ (
  .A1({ S22113 }),
  .A2({ S9119 }),
  .A3({ S22115 }),
  .ZN({ S22116 })
);
OAI21_X1 #() 
OAI21_X1_1923_ (
  .A({ S22116 }),
  .B1({ S22109 }),
  .B2({ S22111 }),
  .ZN({ S22117 })
);
AOI21_X1 #() 
AOI21_X1_2030_ (
  .A({ S22107 }),
  .B1({ S25957[1173] }),
  .B2({ S22117 }),
  .ZN({ S22118 })
);
NAND2_X1 #() 
NAND2_X1_3748_ (
  .A1({ S50 }),
  .A2({ S25957[1168] }),
  .ZN({ S22119 })
);
NAND2_X1 #() 
NAND2_X1_3749_ (
  .A1({ S22097 }),
  .A2({ S22055 }),
  .ZN({ S22120 })
);
AOI21_X1 #() 
AOI21_X1_2031_ (
  .A({ S9119 }),
  .B1({ S22120 }),
  .B2({ S22119 }),
  .ZN({ S22121 })
);
AOI21_X1 #() 
AOI21_X1_2032_ (
  .A({ S25957[1171] }),
  .B1({ S25957[1170] }),
  .B2({ S25957[1169] }),
  .ZN({ S22122 })
);
INV_X1 #() 
INV_X1_1240_ (
  .A({ S22122 }),
  .ZN({ S22123 })
);
NOR3_X1 #() 
NOR3_X1_129_ (
  .A1({ S22123 }),
  .A2({ S22040 }),
  .A3({ S22080 }),
  .ZN({ S22124 })
);
NAND3_X1 #() 
NAND3_X1_3996_ (
  .A1({ S22095 }),
  .A2({ S25957[1171] }),
  .A3({ S22037 }),
  .ZN({ S22125 })
);
NAND2_X1 #() 
NAND2_X1_3750_ (
  .A1({ S22125 }),
  .A2({ S9119 }),
  .ZN({ S22126 })
);
NOR2_X1 #() 
NOR2_X1_953_ (
  .A1({ S22124 }),
  .A2({ S22126 }),
  .ZN({ S22127 })
);
OAI21_X1 #() 
OAI21_X1_1924_ (
  .A({ S25957[1173] }),
  .B1({ S22121 }),
  .B2({ S22127 }),
  .ZN({ S22128 })
);
INV_X1 #() 
INV_X1_1241_ (
  .A({ S22082 }),
  .ZN({ S22129 })
);
NOR2_X1 #() 
NOR2_X1_954_ (
  .A1({ S22043 }),
  .A2({ S25957[1171] }),
  .ZN({ S22130 })
);
NAND2_X1 #() 
NAND2_X1_3751_ (
  .A1({ S22130 }),
  .A2({ S22129 }),
  .ZN({ S22131 })
);
NAND2_X1 #() 
NAND2_X1_3752_ (
  .A1({ S22131 }),
  .A2({ S25957[1172] }),
  .ZN({ S22132 })
);
AOI21_X1 #() 
AOI21_X1_2033_ (
  .A({ S22132 }),
  .B1({ S22047 }),
  .B2({ S25957[1171] }),
  .ZN({ S22133 })
);
NAND2_X1 #() 
NAND2_X1_3753_ (
  .A1({ S22037 }),
  .A2({ S25957[1170] }),
  .ZN({ S22134 })
);
OAI221_X1 #() 
OAI221_X1_111_ (
  .A({ S9119 }),
  .B1({ S22053 }),
  .B2({ S22134 }),
  .C1({ S22099 }),
  .C2({ S50 }),
  .ZN({ S22135 })
);
NAND2_X1 #() 
NAND2_X1_3754_ (
  .A1({ S22135 }),
  .A2({ S22051 }),
  .ZN({ S22136 })
);
OAI211_X1 #() 
OAI211_X1_1302_ (
  .A({ S22128 }),
  .B({ S7741 }),
  .C1({ S22133 }),
  .C2({ S22136 }),
  .ZN({ S22137 })
);
OAI21_X1 #() 
OAI21_X1_1925_ (
  .A({ S22137 }),
  .B1({ S22118 }),
  .B2({ S7741 }),
  .ZN({ S22138 })
);
NAND2_X1 #() 
NAND2_X1_3755_ (
  .A1({ S22138 }),
  .A2({ S22094 }),
  .ZN({ S22139 })
);
AND2_X1 #() 
AND2_X1_230_ (
  .A1({ S22139 }),
  .A2({ S22093 }),
  .ZN({ S22140 })
);
NAND2_X1 #() 
NAND2_X1_3756_ (
  .A1({ S22140 }),
  .A2({ S25957[1279] }),
  .ZN({ S22141 })
);
OR2_X1 #() 
OR2_X1_52_ (
  .A1({ S22140 }),
  .A2({ S25957[1279] }),
  .ZN({ S22142 })
);
NAND2_X1 #() 
NAND2_X1_3757_ (
  .A1({ S22142 }),
  .A2({ S22141 }),
  .ZN({ S22143 })
);
INV_X1 #() 
INV_X1_1242_ (
  .A({ S22143 }),
  .ZN({ S25957[1151] })
);
NAND2_X1 #() 
NAND2_X1_3758_ (
  .A1({ S25957[1151] }),
  .A2({ S25957[1247] }),
  .ZN({ S22144 })
);
INV_X1 #() 
INV_X1_1243_ (
  .A({ S25957[1247] }),
  .ZN({ S22145 })
);
NAND2_X1 #() 
NAND2_X1_3759_ (
  .A1({ S22143 }),
  .A2({ S22145 }),
  .ZN({ S22146 })
);
NAND3_X1 #() 
NAND3_X1_3997_ (
  .A1({ S22144 }),
  .A2({ S25956[31] }),
  .A3({ S22146 }),
  .ZN({ S22147 })
);
NAND2_X1 #() 
NAND2_X1_3760_ (
  .A1({ S22144 }),
  .A2({ S22146 }),
  .ZN({ S22148 })
);
NAND2_X1 #() 
NAND2_X1_3761_ (
  .A1({ S22148 }),
  .A2({ S18081 }),
  .ZN({ S22149 })
);
NAND2_X1 #() 
NAND2_X1_3762_ (
  .A1({ S22149 }),
  .A2({ S22147 }),
  .ZN({ S22150 })
);
INV_X1 #() 
INV_X1_1244_ (
  .A({ S22150 }),
  .ZN({ S25957[1055] })
);
NOR2_X1 #() 
NOR2_X1_955_ (
  .A1({ S19731 }),
  .A2({ S19732 }),
  .ZN({ S25957[1214] })
);
NAND2_X1 #() 
NAND2_X1_3763_ (
  .A1({ S19728 }),
  .A2({ S19729 }),
  .ZN({ S25957[1246] })
);
INV_X1 #() 
INV_X1_1245_ (
  .A({ S25957[1246] }),
  .ZN({ S22151 })
);
NAND2_X1 #() 
NAND2_X1_3764_ (
  .A1({ S20682 }),
  .A2({ S20616 }),
  .ZN({ S22152 })
);
NOR2_X1 #() 
NOR2_X1_956_ (
  .A1({ S22084 }),
  .A2({ S22074 }),
  .ZN({ S22153 })
);
NAND3_X1 #() 
NAND3_X1_3998_ (
  .A1({ S22065 }),
  .A2({ S25957[1171] }),
  .A3({ S82 }),
  .ZN({ S22154 })
);
INV_X1 #() 
INV_X1_1246_ (
  .A({ S22154 }),
  .ZN({ S22155 })
);
AOI21_X1 #() 
AOI21_X1_2034_ (
  .A({ S22153 }),
  .B1({ S22152 }),
  .B2({ S22155 }),
  .ZN({ S22156 })
);
OAI211_X1 #() 
OAI211_X1_1303_ (
  .A({ S22069 }),
  .B({ S25957[1172] }),
  .C1({ S25957[1171] }),
  .C2({ S22083 }),
  .ZN({ S22157 })
);
OAI211_X1 #() 
OAI211_X1_1304_ (
  .A({ S22051 }),
  .B({ S22157 }),
  .C1({ S22156 }),
  .C2({ S25957[1172] }),
  .ZN({ S22158 })
);
NOR2_X1 #() 
NOR2_X1_957_ (
  .A1({ S22134 }),
  .A2({ S22046 }),
  .ZN({ S22159 })
);
NOR2_X1 #() 
NOR2_X1_958_ (
  .A1({ S22052 }),
  .A2({ S25957[1170] }),
  .ZN({ S22160 })
);
OAI21_X1 #() 
OAI21_X1_1926_ (
  .A({ S50 }),
  .B1({ S22159 }),
  .B2({ S22160 }),
  .ZN({ S22161 })
);
NOR2_X1 #() 
NOR2_X1_959_ (
  .A1({ S50 }),
  .A2({ S20682 }),
  .ZN({ S22162 })
);
AOI21_X1 #() 
AOI21_X1_2035_ (
  .A({ S9119 }),
  .B1({ S22162 }),
  .B2({ S25957[1169] }),
  .ZN({ S22163 })
);
NAND2_X1 #() 
NAND2_X1_3765_ (
  .A1({ S22052 }),
  .A2({ S20682 }),
  .ZN({ S22164 })
);
NAND2_X1 #() 
NAND2_X1_3766_ (
  .A1({ S22164 }),
  .A2({ S22076 }),
  .ZN({ S22165 })
);
INV_X1 #() 
INV_X1_1247_ (
  .A({ S22165 }),
  .ZN({ S22166 })
);
INV_X1 #() 
INV_X1_1248_ (
  .A({ S82 }),
  .ZN({ S22167 })
);
NAND3_X1 #() 
NAND3_X1_3999_ (
  .A1({ S25957[1170] }),
  .A2({ S25957[1168] }),
  .A3({ S25957[1169] }),
  .ZN({ S22168 })
);
INV_X1 #() 
INV_X1_1249_ (
  .A({ S22168 }),
  .ZN({ S22169 })
);
OAI21_X1 #() 
OAI21_X1_1927_ (
  .A({ S50 }),
  .B1({ S22169 }),
  .B2({ S22167 }),
  .ZN({ S22170 })
);
OAI21_X1 #() 
OAI21_X1_1928_ (
  .A({ S22170 }),
  .B1({ S22166 }),
  .B2({ S50 }),
  .ZN({ S22171 })
);
AOI22_X1 #() 
AOI22_X1_424_ (
  .A1({ S22171 }),
  .A2({ S9119 }),
  .B1({ S22161 }),
  .B2({ S22163 }),
  .ZN({ S22172 })
);
OAI21_X1 #() 
OAI21_X1_1929_ (
  .A({ S22158 }),
  .B1({ S22051 }),
  .B2({ S22172 }),
  .ZN({ S22173 })
);
AOI21_X1 #() 
AOI21_X1_2036_ (
  .A({ S50 }),
  .B1({ S22134 }),
  .B2({ S22086 }),
  .ZN({ S22174 })
);
NOR3_X1 #() 
NOR3_X1_130_ (
  .A1({ S22153 }),
  .A2({ S22174 }),
  .A3({ S9119 }),
  .ZN({ S22175 })
);
OR2_X1 #() 
OR2_X1_53_ (
  .A1({ S22056 }),
  .A2({ S22066 }),
  .ZN({ S22176 })
);
NAND3_X1 #() 
NAND3_X1_4000_ (
  .A1({ S22134 }),
  .A2({ S22058 }),
  .A3({ S25957[1171] }),
  .ZN({ S22177 })
);
NAND2_X1 #() 
NAND2_X1_3767_ (
  .A1({ S22065 }),
  .A2({ S22076 }),
  .ZN({ S22178 })
);
AOI21_X1 #() 
AOI21_X1_2037_ (
  .A({ S9119 }),
  .B1({ S22178 }),
  .B2({ S50 }),
  .ZN({ S22179 })
);
AOI22_X1 #() 
AOI22_X1_425_ (
  .A1({ S22176 }),
  .A2({ S9119 }),
  .B1({ S22179 }),
  .B2({ S22177 }),
  .ZN({ S22180 })
);
NAND3_X1 #() 
NAND3_X1_4001_ (
  .A1({ S22152 }),
  .A2({ S25957[1171] }),
  .A3({ S22055 }),
  .ZN({ S22181 })
);
OAI21_X1 #() 
OAI21_X1_1930_ (
  .A({ S22101 }),
  .B1({ S22167 }),
  .B2({ S22181 }),
  .ZN({ S22182 })
);
NAND2_X1 #() 
NAND2_X1_3768_ (
  .A1({ S22182 }),
  .A2({ S22051 }),
  .ZN({ S22183 })
);
OAI22_X1 #() 
OAI22_X1_101_ (
  .A1({ S22183 }),
  .A2({ S22175 }),
  .B1({ S22180 }),
  .B2({ S22051 }),
  .ZN({ S22184 })
);
NAND2_X1 #() 
NAND2_X1_3769_ (
  .A1({ S22184 }),
  .A2({ S25957[1174] }),
  .ZN({ S22185 })
);
OAI211_X1 #() 
OAI211_X1_1305_ (
  .A({ S22185 }),
  .B({ S25957[1175] }),
  .C1({ S22173 }),
  .C2({ S25957[1174] }),
  .ZN({ S22186 })
);
NAND2_X1 #() 
NAND2_X1_3770_ (
  .A1({ S22044 }),
  .A2({ S25957[1171] }),
  .ZN({ S22187 })
);
INV_X1 #() 
INV_X1_1250_ (
  .A({ S22187 }),
  .ZN({ S22188 })
);
AOI211_X1 #() 
AOI211_X1_63_ (
  .A({ S9119 }),
  .B({ S22088 }),
  .C1({ S22188 }),
  .C2({ S22035 }),
  .ZN({ S22189 })
);
NOR2_X1 #() 
NOR2_X1_960_ (
  .A1({ S22037 }),
  .A2({ S25957[1170] }),
  .ZN({ S22190 })
);
INV_X1 #() 
INV_X1_1251_ (
  .A({ S22190 }),
  .ZN({ S22191 })
);
AOI22_X1 #() 
AOI22_X1_426_ (
  .A1({ S22191 }),
  .A2({ S22122 }),
  .B1({ S22112 }),
  .B2({ S22095 }),
  .ZN({ S22192 })
);
AOI21_X1 #() 
AOI21_X1_2038_ (
  .A({ S22189 }),
  .B1({ S9119 }),
  .B2({ S22192 }),
  .ZN({ S22193 })
);
OAI211_X1 #() 
OAI211_X1_1306_ (
  .A({ S22113 }),
  .B({ S25957[1172] }),
  .C1({ S25957[1171] }),
  .C2({ S22190 }),
  .ZN({ S22194 })
);
INV_X1 #() 
INV_X1_1252_ (
  .A({ S22047 }),
  .ZN({ S22195 })
);
OAI21_X1 #() 
OAI21_X1_1931_ (
  .A({ S25957[1171] }),
  .B1({ S22195 }),
  .B2({ S22102 }),
  .ZN({ S22196 })
);
OAI211_X1 #() 
OAI211_X1_1307_ (
  .A({ S22194 }),
  .B({ S22051 }),
  .C1({ S25957[1172] }),
  .C2({ S22196 }),
  .ZN({ S22197 })
);
OAI21_X1 #() 
OAI21_X1_1932_ (
  .A({ S22197 }),
  .B1({ S22193 }),
  .B2({ S22051 }),
  .ZN({ S22198 })
);
AOI211_X1 #() 
AOI211_X1_64_ (
  .A({ S25957[1172] }),
  .B({ S22174 }),
  .C1({ S50 }),
  .C2({ S22129 }),
  .ZN({ S22199 })
);
NAND2_X1 #() 
NAND2_X1_3771_ (
  .A1({ S22065 }),
  .A2({ S22052 }),
  .ZN({ S22200 })
);
NAND2_X1 #() 
NAND2_X1_3772_ (
  .A1({ S22200 }),
  .A2({ S25957[1171] }),
  .ZN({ S22201 })
);
AOI21_X1 #() 
AOI21_X1_2039_ (
  .A({ S9119 }),
  .B1({ S22088 }),
  .B2({ S22099 }),
  .ZN({ S22202 })
);
NAND2_X1 #() 
NAND2_X1_3773_ (
  .A1({ S20676 }),
  .A2({ S50 }),
  .ZN({ S22203 })
);
AND3_X1 #() 
AND3_X1_143_ (
  .A1({ S22200 }),
  .A2({ S9119 }),
  .A3({ S22203 }),
  .ZN({ S22204 })
);
AOI21_X1 #() 
AOI21_X1_2040_ (
  .A({ S22204 }),
  .B1({ S22202 }),
  .B2({ S22201 }),
  .ZN({ S22205 })
);
NAND3_X1 #() 
NAND3_X1_4002_ (
  .A1({ S22055 }),
  .A2({ S50 }),
  .A3({ S20616 }),
  .ZN({ S22206 })
);
OAI211_X1 #() 
OAI211_X1_1308_ (
  .A({ S22206 }),
  .B({ S25957[1172] }),
  .C1({ S50 }),
  .C2({ S22095 }),
  .ZN({ S22207 })
);
NAND2_X1 #() 
NAND2_X1_3774_ (
  .A1({ S22207 }),
  .A2({ S22051 }),
  .ZN({ S22208 })
);
OAI22_X1 #() 
OAI22_X1_102_ (
  .A1({ S22205 }),
  .A2({ S22051 }),
  .B1({ S22199 }),
  .B2({ S22208 }),
  .ZN({ S22209 })
);
NAND2_X1 #() 
NAND2_X1_3775_ (
  .A1({ S22209 }),
  .A2({ S25957[1174] }),
  .ZN({ S22210 })
);
OAI211_X1 #() 
OAI211_X1_1309_ (
  .A({ S22210 }),
  .B({ S22094 }),
  .C1({ S22198 }),
  .C2({ S25957[1174] }),
  .ZN({ S22211 })
);
NAND3_X1 #() 
NAND3_X1_4003_ (
  .A1({ S22186 }),
  .A2({ S25957[1278] }),
  .A3({ S22211 }),
  .ZN({ S22212 })
);
NAND2_X1 #() 
NAND2_X1_3776_ (
  .A1({ S22186 }),
  .A2({ S22211 }),
  .ZN({ S22213 })
);
NAND2_X1 #() 
NAND2_X1_3777_ (
  .A1({ S22213 }),
  .A2({ S19727 }),
  .ZN({ S22214 })
);
NAND2_X1 #() 
NAND2_X1_3778_ (
  .A1({ S22214 }),
  .A2({ S22212 }),
  .ZN({ S25957[1150] })
);
NAND2_X1 #() 
NAND2_X1_3779_ (
  .A1({ S25957[1150] }),
  .A2({ S22151 }),
  .ZN({ S22215 })
);
NAND3_X1 #() 
NAND3_X1_4004_ (
  .A1({ S22214 }),
  .A2({ S25957[1246] }),
  .A3({ S22212 }),
  .ZN({ S22216 })
);
NAND2_X1 #() 
NAND2_X1_3780_ (
  .A1({ S22215 }),
  .A2({ S22216 }),
  .ZN({ S25957[1118] })
);
NAND2_X1 #() 
NAND2_X1_3781_ (
  .A1({ S25957[1118] }),
  .A2({ S25956[30] }),
  .ZN({ S22217 })
);
NAND3_X1 #() 
NAND3_X1_4005_ (
  .A1({ S22215 }),
  .A2({ S22216 }),
  .A3({ S18092 }),
  .ZN({ S22218 })
);
NAND2_X1 #() 
NAND2_X1_3782_ (
  .A1({ S22217 }),
  .A2({ S22218 }),
  .ZN({ S22219 })
);
INV_X1 #() 
INV_X1_1253_ (
  .A({ S22219 }),
  .ZN({ S25957[1054] })
);
NOR2_X1 #() 
NOR2_X1_961_ (
  .A1({ S19806 }),
  .A2({ S19807 }),
  .ZN({ S25957[1245] })
);
NAND2_X1 #() 
NAND2_X1_3783_ (
  .A1({ S19804 }),
  .A2({ S19801 }),
  .ZN({ S25957[1277] })
);
INV_X1 #() 
INV_X1_1254_ (
  .A({ S25957[1277] }),
  .ZN({ S22220 })
);
NAND2_X1 #() 
NAND2_X1_3784_ (
  .A1({ S22054 }),
  .A2({ S25957[1170] }),
  .ZN({ S22221 })
);
NAND2_X1 #() 
NAND2_X1_3785_ (
  .A1({ S22164 }),
  .A2({ S25957[1171] }),
  .ZN({ S22222 })
);
NAND3_X1 #() 
NAND3_X1_4006_ (
  .A1({ S22221 }),
  .A2({ S25957[1172] }),
  .A3({ S22222 }),
  .ZN({ S22223 })
);
INV_X1 #() 
INV_X1_1255_ (
  .A({ S22159 }),
  .ZN({ S22224 })
);
NAND2_X1 #() 
NAND2_X1_3786_ (
  .A1({ S22224 }),
  .A2({ S9119 }),
  .ZN({ S22225 })
);
OAI21_X1 #() 
OAI21_X1_1933_ (
  .A({ S22223 }),
  .B1({ S22225 }),
  .B2({ S22174 }),
  .ZN({ S22226 })
);
NAND3_X1 #() 
NAND3_X1_4007_ (
  .A1({ S22076 }),
  .A2({ S22035 }),
  .A3({ S25957[1171] }),
  .ZN({ S22227 })
);
INV_X1 #() 
INV_X1_1256_ (
  .A({ S22227 }),
  .ZN({ S22228 })
);
OAI211_X1 #() 
OAI211_X1_1310_ (
  .A({ S22065 }),
  .B({ S9119 }),
  .C1({ S25957[1171] }),
  .C2({ S20676 }),
  .ZN({ S22229 })
);
NAND2_X1 #() 
NAND2_X1_3787_ (
  .A1({ S20616 }),
  .A2({ S25957[1171] }),
  .ZN({ S22230 })
);
INV_X1 #() 
INV_X1_1257_ (
  .A({ S22230 }),
  .ZN({ S22231 })
);
AOI22_X1 #() 
AOI22_X1_427_ (
  .A1({ S22054 }),
  .A2({ S22083 }),
  .B1({ S22231 }),
  .B2({ S22055 }),
  .ZN({ S22232 })
);
OAI221_X1 #() 
OAI221_X1_112_ (
  .A({ S25957[1173] }),
  .B1({ S22228 }),
  .B2({ S22229 }),
  .C1({ S22232 }),
  .C2({ S9119 }),
  .ZN({ S22233 })
);
OAI21_X1 #() 
OAI21_X1_1934_ (
  .A({ S22233 }),
  .B1({ S22226 }),
  .B2({ S25957[1173] }),
  .ZN({ S22234 })
);
NAND2_X1 #() 
NAND2_X1_3788_ (
  .A1({ S22234 }),
  .A2({ S25957[1174] }),
  .ZN({ S22235 })
);
AOI21_X1 #() 
AOI21_X1_2041_ (
  .A({ S9119 }),
  .B1({ S22041 }),
  .B2({ S22035 }),
  .ZN({ S22236 })
);
OAI21_X1 #() 
OAI21_X1_1935_ (
  .A({ S22236 }),
  .B1({ S50 }),
  .B2({ S22100 }),
  .ZN({ S22237 })
);
NAND2_X1 #() 
NAND2_X1_3789_ (
  .A1({ S22054 }),
  .A2({ S22055 }),
  .ZN({ S22238 })
);
NAND2_X1 #() 
NAND2_X1_3790_ (
  .A1({ S20676 }),
  .A2({ S25957[1171] }),
  .ZN({ S22239 })
);
AND2_X1 #() 
AND2_X1_231_ (
  .A1({ S22239 }),
  .A2({ S9119 }),
  .ZN({ S22240 })
);
AOI21_X1 #() 
AOI21_X1_2042_ (
  .A({ S22051 }),
  .B1({ S22238 }),
  .B2({ S22240 }),
  .ZN({ S22241 })
);
NOR2_X1 #() 
NOR2_X1_962_ (
  .A1({ S82 }),
  .A2({ S25957[1170] }),
  .ZN({ S22242 })
);
OR2_X1 #() 
OR2_X1_54_ (
  .A1({ S22082 }),
  .A2({ S22242 }),
  .ZN({ S22243 })
);
AOI21_X1 #() 
AOI21_X1_2043_ (
  .A({ S22130 }),
  .B1({ S22243 }),
  .B2({ S25957[1171] }),
  .ZN({ S22244 })
);
NAND3_X1 #() 
NAND3_X1_4008_ (
  .A1({ S22035 }),
  .A2({ S20682 }),
  .A3({ S82 }),
  .ZN({ S22245 })
);
NOR2_X1 #() 
NOR2_X1_963_ (
  .A1({ S22245 }),
  .A2({ S50 }),
  .ZN({ S22246 })
);
NOR2_X1 #() 
NOR2_X1_964_ (
  .A1({ S25957[1170] }),
  .A2({ S20616 }),
  .ZN({ S22247 })
);
OAI21_X1 #() 
OAI21_X1_1936_ (
  .A({ S25957[1172] }),
  .B1({ S22203 }),
  .B2({ S22247 }),
  .ZN({ S22248 })
);
OAI22_X1 #() 
OAI22_X1_103_ (
  .A1({ S22244 }),
  .A2({ S25957[1172] }),
  .B1({ S22246 }),
  .B2({ S22248 }),
  .ZN({ S22249 })
);
AOI22_X1 #() 
AOI22_X1_428_ (
  .A1({ S22249 }),
  .A2({ S22051 }),
  .B1({ S22237 }),
  .B2({ S22241 }),
  .ZN({ S22250 })
);
OAI21_X1 #() 
OAI21_X1_1937_ (
  .A({ S22235 }),
  .B1({ S22250 }),
  .B2({ S25957[1174] }),
  .ZN({ S22251 })
);
NAND2_X1 #() 
NAND2_X1_3791_ (
  .A1({ S22251 }),
  .A2({ S25957[1175] }),
  .ZN({ S22252 })
);
AOI21_X1 #() 
AOI21_X1_2044_ (
  .A({ S50 }),
  .B1({ S22168 }),
  .B2({ S22152 }),
  .ZN({ S22253 })
);
NAND2_X1 #() 
NAND2_X1_3792_ (
  .A1({ S22164 }),
  .A2({ S22036 }),
  .ZN({ S22254 })
);
AOI21_X1 #() 
AOI21_X1_2045_ (
  .A({ S22253 }),
  .B1({ S50 }),
  .B2({ S22254 }),
  .ZN({ S22255 })
);
NAND4_X1 #() 
NAND4_X1_441_ (
  .A1({ S22168 }),
  .A2({ S22152 }),
  .A3({ S22055 }),
  .A4({ S50 }),
  .ZN({ S22256 })
);
NAND3_X1 #() 
NAND3_X1_4009_ (
  .A1({ S22037 }),
  .A2({ S25957[1171] }),
  .A3({ S20682 }),
  .ZN({ S22257 })
);
AND2_X1 #() 
AND2_X1_232_ (
  .A1({ S22257 }),
  .A2({ S25957[1172] }),
  .ZN({ S22258 })
);
AOI21_X1 #() 
AOI21_X1_2046_ (
  .A({ S7741 }),
  .B1({ S22256 }),
  .B2({ S22258 }),
  .ZN({ S22259 })
);
OAI21_X1 #() 
OAI21_X1_1938_ (
  .A({ S22259 }),
  .B1({ S25957[1172] }),
  .B2({ S22255 }),
  .ZN({ S22260 })
);
NAND4_X1 #() 
NAND4_X1_442_ (
  .A1({ S22152 }),
  .A2({ S22052 }),
  .A3({ S50 }),
  .A4({ S22037 }),
  .ZN({ S22261 })
);
NAND3_X1 #() 
NAND3_X1_4010_ (
  .A1({ S22224 }),
  .A2({ S25957[1171] }),
  .A3({ S22191 }),
  .ZN({ S22262 })
);
NAND3_X1 #() 
NAND3_X1_4011_ (
  .A1({ S22262 }),
  .A2({ S25957[1172] }),
  .A3({ S22261 }),
  .ZN({ S22263 })
);
OAI21_X1 #() 
OAI21_X1_1939_ (
  .A({ S22061 }),
  .B1({ S25957[1171] }),
  .B2({ S22168 }),
  .ZN({ S22264 })
);
NAND2_X1 #() 
NAND2_X1_3793_ (
  .A1({ S22264 }),
  .A2({ S9119 }),
  .ZN({ S22265 })
);
NAND3_X1 #() 
NAND3_X1_4012_ (
  .A1({ S22263 }),
  .A2({ S7741 }),
  .A3({ S22265 }),
  .ZN({ S22266 })
);
AOI21_X1 #() 
AOI21_X1_2047_ (
  .A({ S25957[1173] }),
  .B1({ S22266 }),
  .B2({ S22260 }),
  .ZN({ S22267 })
);
AOI21_X1 #() 
AOI21_X1_2048_ (
  .A({ S50 }),
  .B1({ S22046 }),
  .B2({ S20682 }),
  .ZN({ S22268 })
);
INV_X1 #() 
INV_X1_1258_ (
  .A({ S22268 }),
  .ZN({ S22269 })
);
NAND3_X1 #() 
NAND3_X1_4013_ (
  .A1({ S22083 }),
  .A2({ S22114 }),
  .A3({ S50 }),
  .ZN({ S22270 })
);
OAI21_X1 #() 
OAI21_X1_1940_ (
  .A({ S22270 }),
  .B1({ S22269 }),
  .B2({ S22159 }),
  .ZN({ S22271 })
);
OAI21_X1 #() 
OAI21_X1_1941_ (
  .A({ S22230 }),
  .B1({ S22053 }),
  .B2({ S22247 }),
  .ZN({ S22272 })
);
AOI21_X1 #() 
AOI21_X1_2049_ (
  .A({ S7741 }),
  .B1({ S9119 }),
  .B2({ S22272 }),
  .ZN({ S22273 })
);
OAI21_X1 #() 
OAI21_X1_1942_ (
  .A({ S22273 }),
  .B1({ S9119 }),
  .B2({ S22271 }),
  .ZN({ S22274 })
);
NAND2_X1 #() 
NAND2_X1_3794_ (
  .A1({ S22066 }),
  .A2({ S22040 }),
  .ZN({ S22275 })
);
NAND3_X1 #() 
NAND3_X1_4014_ (
  .A1({ S22275 }),
  .A2({ S25957[1172] }),
  .A3({ S22181 }),
  .ZN({ S22276 })
);
NAND3_X1 #() 
NAND3_X1_4015_ (
  .A1({ S25957[1170] }),
  .A2({ S25957[1168] }),
  .A3({ S25957[1171] }),
  .ZN({ S22277 })
);
INV_X1 #() 
INV_X1_1259_ (
  .A({ S22277 }),
  .ZN({ S22278 })
);
OAI21_X1 #() 
OAI21_X1_1943_ (
  .A({ S22204 }),
  .B1({ S22278 }),
  .B2({ S22075 }),
  .ZN({ S22279 })
);
NAND3_X1 #() 
NAND3_X1_4016_ (
  .A1({ S22279 }),
  .A2({ S7741 }),
  .A3({ S22276 }),
  .ZN({ S22280 })
);
AOI21_X1 #() 
AOI21_X1_2050_ (
  .A({ S22051 }),
  .B1({ S22274 }),
  .B2({ S22280 }),
  .ZN({ S22281 })
);
OR3_X1 #() 
OR3_X1_24_ (
  .A1({ S22267 }),
  .A2({ S22281 }),
  .A3({ S25957[1175] }),
  .ZN({ S22282 })
);
NAND3_X1 #() 
NAND3_X1_4017_ (
  .A1({ S22252 }),
  .A2({ S22282 }),
  .A3({ S22220 }),
  .ZN({ S22283 })
);
OR2_X1 #() 
OR2_X1_55_ (
  .A1({ S22251 }),
  .A2({ S22094 }),
  .ZN({ S22284 })
);
OAI21_X1 #() 
OAI21_X1_1944_ (
  .A({ S22094 }),
  .B1({ S22267 }),
  .B2({ S22281 }),
  .ZN({ S22285 })
);
NAND3_X1 #() 
NAND3_X1_4018_ (
  .A1({ S22284 }),
  .A2({ S25957[1277] }),
  .A3({ S22285 }),
  .ZN({ S22286 })
);
NAND2_X1 #() 
NAND2_X1_3795_ (
  .A1({ S22286 }),
  .A2({ S22283 }),
  .ZN({ S25957[1149] })
);
NAND2_X1 #() 
NAND2_X1_3796_ (
  .A1({ S25957[1149] }),
  .A2({ S25957[1245] }),
  .ZN({ S22287 })
);
INV_X1 #() 
INV_X1_1260_ (
  .A({ S25957[1245] }),
  .ZN({ S22288 })
);
NAND3_X1 #() 
NAND3_X1_4019_ (
  .A1({ S22286 }),
  .A2({ S22288 }),
  .A3({ S22283 }),
  .ZN({ S22289 })
);
NAND3_X1 #() 
NAND3_X1_4020_ (
  .A1({ S22287 }),
  .A2({ S22289 }),
  .A3({ S18103 }),
  .ZN({ S22290 })
);
NAND2_X1 #() 
NAND2_X1_3797_ (
  .A1({ S25957[1149] }),
  .A2({ S22288 }),
  .ZN({ S22291 })
);
NAND3_X1 #() 
NAND3_X1_4021_ (
  .A1({ S22286 }),
  .A2({ S25957[1245] }),
  .A3({ S22283 }),
  .ZN({ S22292 })
);
NAND3_X1 #() 
NAND3_X1_4022_ (
  .A1({ S22291 }),
  .A2({ S22292 }),
  .A3({ S25956[29] }),
  .ZN({ S22293 })
);
AND2_X1 #() 
AND2_X1_233_ (
  .A1({ S22293 }),
  .A2({ S22290 }),
  .ZN({ S22294 })
);
INV_X1 #() 
INV_X1_1261_ (
  .A({ S22294 }),
  .ZN({ S25957[1053] })
);
NOR2_X1 #() 
NOR2_X1_965_ (
  .A1({ S19876 }),
  .A2({ S19880 }),
  .ZN({ S25957[1212] })
);
NAND2_X1 #() 
NAND2_X1_3798_ (
  .A1({ S19878 }),
  .A2({ S19879 }),
  .ZN({ S25957[1244] })
);
NAND2_X1 #() 
NAND2_X1_3799_ (
  .A1({ S19871 }),
  .A2({ S19867 }),
  .ZN({ S25957[1276] })
);
AOI21_X1 #() 
AOI21_X1_2051_ (
  .A({ S25957[1171] }),
  .B1({ S22164 }),
  .B2({ S22047 }),
  .ZN({ S22295 })
);
NAND2_X1 #() 
NAND2_X1_3800_ (
  .A1({ S22065 }),
  .A2({ S20676 }),
  .ZN({ S22296 })
);
NOR2_X1 #() 
NOR2_X1_966_ (
  .A1({ S22296 }),
  .A2({ S50 }),
  .ZN({ S22297 })
);
NOR3_X1 #() 
NOR3_X1_131_ (
  .A1({ S22295 }),
  .A2({ S22297 }),
  .A3({ S25957[1172] }),
  .ZN({ S22298 })
);
NAND2_X1 #() 
NAND2_X1_3801_ (
  .A1({ S22056 }),
  .A2({ S22095 }),
  .ZN({ S22299 })
);
AOI21_X1 #() 
AOI21_X1_2052_ (
  .A({ S9119 }),
  .B1({ S22130 }),
  .B2({ S22047 }),
  .ZN({ S22300 })
);
AOI21_X1 #() 
AOI21_X1_2053_ (
  .A({ S22298 }),
  .B1({ S22299 }),
  .B2({ S22300 }),
  .ZN({ S22301 })
);
NAND2_X1 #() 
NAND2_X1_3802_ (
  .A1({ S22164 }),
  .A2({ S22134 }),
  .ZN({ S22302 })
);
NAND2_X1 #() 
NAND2_X1_3803_ (
  .A1({ S22302 }),
  .A2({ S50 }),
  .ZN({ S22303 })
);
OAI211_X1 #() 
OAI211_X1_1311_ (
  .A({ S22303 }),
  .B({ S25957[1172] }),
  .C1({ S22060 }),
  .C2({ S22269 }),
  .ZN({ S22304 })
);
AOI21_X1 #() 
AOI21_X1_2054_ (
  .A({ S25957[1171] }),
  .B1({ S22103 }),
  .B2({ S22099 }),
  .ZN({ S22305 })
);
AOI21_X1 #() 
AOI21_X1_2055_ (
  .A({ S50 }),
  .B1({ S22047 }),
  .B2({ S22083 }),
  .ZN({ S22306 })
);
NOR3_X1 #() 
NOR3_X1_132_ (
  .A1({ S22305 }),
  .A2({ S22306 }),
  .A3({ S25957[1172] }),
  .ZN({ S22307 })
);
NOR2_X1 #() 
NOR2_X1_967_ (
  .A1({ S22307 }),
  .A2({ S22051 }),
  .ZN({ S22308 })
);
AOI22_X1 #() 
AOI22_X1_429_ (
  .A1({ S22304 }),
  .A2({ S22308 }),
  .B1({ S22301 }),
  .B2({ S22051 }),
  .ZN({ S22309 })
);
NAND2_X1 #() 
NAND2_X1_3804_ (
  .A1({ S22309 }),
  .A2({ S7741 }),
  .ZN({ S22310 })
);
NAND3_X1 #() 
NAND3_X1_4023_ (
  .A1({ S22036 }),
  .A2({ S50 }),
  .A3({ S22055 }),
  .ZN({ S22311 })
);
INV_X1 #() 
INV_X1_1262_ (
  .A({ S22311 }),
  .ZN({ S22312 })
);
OAI211_X1 #() 
OAI211_X1_1312_ (
  .A({ S22238 }),
  .B({ S25957[1172] }),
  .C1({ S22239 }),
  .C2({ S22247 }),
  .ZN({ S22313 })
);
OAI21_X1 #() 
OAI21_X1_1945_ (
  .A({ S22313 }),
  .B1({ S22126 }),
  .B2({ S22312 }),
  .ZN({ S22314 })
);
NAND2_X1 #() 
NAND2_X1_3805_ (
  .A1({ S22258 }),
  .A2({ S22045 }),
  .ZN({ S22315 })
);
NAND3_X1 #() 
NAND3_X1_4024_ (
  .A1({ S22095 }),
  .A2({ S50 }),
  .A3({ S20616 }),
  .ZN({ S22316 })
);
NAND3_X1 #() 
NAND3_X1_4025_ (
  .A1({ S22120 }),
  .A2({ S9119 }),
  .A3({ S22316 }),
  .ZN({ S22317 })
);
NAND3_X1 #() 
NAND3_X1_4026_ (
  .A1({ S22317 }),
  .A2({ S22315 }),
  .A3({ S25957[1173] }),
  .ZN({ S22318 })
);
OAI21_X1 #() 
OAI21_X1_1946_ (
  .A({ S22318 }),
  .B1({ S22314 }),
  .B2({ S25957[1173] }),
  .ZN({ S22319 })
);
OR2_X1 #() 
OR2_X1_56_ (
  .A1({ S22319 }),
  .A2({ S7741 }),
  .ZN({ S22320 })
);
NAND3_X1 #() 
NAND3_X1_4027_ (
  .A1({ S22310 }),
  .A2({ S22320 }),
  .A3({ S25957[1175] }),
  .ZN({ S22321 })
);
AOI21_X1 #() 
AOI21_X1_2056_ (
  .A({ S9119 }),
  .B1({ S123 }),
  .B2({ S20682 }),
  .ZN({ S22322 })
);
NOR2_X1 #() 
NOR2_X1_968_ (
  .A1({ S22162 }),
  .A2({ S25957[1172] }),
  .ZN({ S22323 })
);
OAI21_X1 #() 
OAI21_X1_1947_ (
  .A({ S22323 }),
  .B1({ S22074 }),
  .B2({ S22043 }),
  .ZN({ S22324 })
);
NAND2_X1 #() 
NAND2_X1_3806_ (
  .A1({ S22055 }),
  .A2({ S50 }),
  .ZN({ S22325 })
);
OAI211_X1 #() 
OAI211_X1_1313_ (
  .A({ S22069 }),
  .B({ S25957[1172] }),
  .C1({ S22178 }),
  .C2({ S22325 }),
  .ZN({ S22326 })
);
NAND3_X1 #() 
NAND3_X1_4028_ (
  .A1({ S22326 }),
  .A2({ S22051 }),
  .A3({ S22324 }),
  .ZN({ S22327 })
);
INV_X1 #() 
INV_X1_1263_ (
  .A({ S22253 }),
  .ZN({ S22328 })
);
AOI21_X1 #() 
AOI21_X1_2057_ (
  .A({ S25957[1170] }),
  .B1({ S22052 }),
  .B2({ S22037 }),
  .ZN({ S22329 })
);
NAND2_X1 #() 
NAND2_X1_3807_ (
  .A1({ S22329 }),
  .A2({ S50 }),
  .ZN({ S22330 })
);
NAND4_X1 #() 
NAND4_X1_443_ (
  .A1({ S22328 }),
  .A2({ S22330 }),
  .A3({ S9119 }),
  .A4({ S22221 }),
  .ZN({ S22331 })
);
NAND2_X1 #() 
NAND2_X1_3808_ (
  .A1({ S22331 }),
  .A2({ S25957[1173] }),
  .ZN({ S22332 })
);
OAI21_X1 #() 
OAI21_X1_1948_ (
  .A({ S22327 }),
  .B1({ S22332 }),
  .B2({ S22322 }),
  .ZN({ S22333 })
);
NAND2_X1 #() 
NAND2_X1_3809_ (
  .A1({ S22333 }),
  .A2({ S25957[1174] }),
  .ZN({ S22334 })
);
NAND3_X1 #() 
NAND3_X1_4029_ (
  .A1({ S22044 }),
  .A2({ S22058 }),
  .A3({ S50 }),
  .ZN({ S22335 })
);
AND2_X1 #() 
AND2_X1_234_ (
  .A1({ S22335 }),
  .A2({ S22154 }),
  .ZN({ S22336 })
);
NAND3_X1 #() 
NAND3_X1_4030_ (
  .A1({ S22083 }),
  .A2({ S25957[1171] }),
  .A3({ S22065 }),
  .ZN({ S22337 })
);
NAND3_X1 #() 
NAND3_X1_4031_ (
  .A1({ S22238 }),
  .A2({ S25957[1172] }),
  .A3({ S22337 }),
  .ZN({ S22338 })
);
OAI211_X1 #() 
OAI211_X1_1314_ (
  .A({ S22051 }),
  .B({ S22338 }),
  .C1({ S22336 }),
  .C2({ S25957[1172] }),
  .ZN({ S22339 })
);
NAND3_X1 #() 
NAND3_X1_4032_ (
  .A1({ S22221 }),
  .A2({ S25957[1172] }),
  .A3({ S22113 }),
  .ZN({ S22340 })
);
AOI21_X1 #() 
AOI21_X1_2058_ (
  .A({ S22246 }),
  .B1({ S81 }),
  .B2({ S50 }),
  .ZN({ S22341 })
);
OAI211_X1 #() 
OAI211_X1_1315_ (
  .A({ S25957[1173] }),
  .B({ S22340 }),
  .C1({ S22341 }),
  .C2({ S25957[1172] }),
  .ZN({ S22342 })
);
NAND3_X1 #() 
NAND3_X1_4033_ (
  .A1({ S22342 }),
  .A2({ S7741 }),
  .A3({ S22339 }),
  .ZN({ S22343 })
);
NAND2_X1 #() 
NAND2_X1_3810_ (
  .A1({ S22334 }),
  .A2({ S22343 }),
  .ZN({ S22344 })
);
NAND2_X1 #() 
NAND2_X1_3811_ (
  .A1({ S22344 }),
  .A2({ S22094 }),
  .ZN({ S22345 })
);
NAND3_X1 #() 
NAND3_X1_4034_ (
  .A1({ S22321 }),
  .A2({ S22345 }),
  .A3({ S25957[1276] }),
  .ZN({ S22346 })
);
INV_X1 #() 
INV_X1_1264_ (
  .A({ S25957[1276] }),
  .ZN({ S22347 })
);
NAND2_X1 #() 
NAND2_X1_3812_ (
  .A1({ S22319 }),
  .A2({ S25957[1174] }),
  .ZN({ S22348 })
);
OAI211_X1 #() 
OAI211_X1_1316_ (
  .A({ S22348 }),
  .B({ S25957[1175] }),
  .C1({ S22309 }),
  .C2({ S25957[1174] }),
  .ZN({ S22349 })
);
NAND3_X1 #() 
NAND3_X1_4035_ (
  .A1({ S22334 }),
  .A2({ S22343 }),
  .A3({ S22094 }),
  .ZN({ S22350 })
);
NAND3_X1 #() 
NAND3_X1_4036_ (
  .A1({ S22349 }),
  .A2({ S22350 }),
  .A3({ S22347 }),
  .ZN({ S22351 })
);
NAND3_X1 #() 
NAND3_X1_4037_ (
  .A1({ S22346 }),
  .A2({ S25957[1244] }),
  .A3({ S22351 }),
  .ZN({ S22352 })
);
INV_X1 #() 
INV_X1_1265_ (
  .A({ S25957[1244] }),
  .ZN({ S22353 })
);
NAND3_X1 #() 
NAND3_X1_4038_ (
  .A1({ S22321 }),
  .A2({ S22345 }),
  .A3({ S22347 }),
  .ZN({ S22354 })
);
NAND3_X1 #() 
NAND3_X1_4039_ (
  .A1({ S22349 }),
  .A2({ S22350 }),
  .A3({ S25957[1276] }),
  .ZN({ S22355 })
);
NAND3_X1 #() 
NAND3_X1_4040_ (
  .A1({ S22354 }),
  .A2({ S22353 }),
  .A3({ S22355 }),
  .ZN({ S22356 })
);
NAND3_X1 #() 
NAND3_X1_4041_ (
  .A1({ S22352 }),
  .A2({ S22356 }),
  .A3({ S25956[28] }),
  .ZN({ S22357 })
);
NAND3_X1 #() 
NAND3_X1_4042_ (
  .A1({ S22346 }),
  .A2({ S22353 }),
  .A3({ S22351 }),
  .ZN({ S22358 })
);
NAND3_X1 #() 
NAND3_X1_4043_ (
  .A1({ S22354 }),
  .A2({ S25957[1244] }),
  .A3({ S22355 }),
  .ZN({ S22359 })
);
NAND3_X1 #() 
NAND3_X1_4044_ (
  .A1({ S22358 }),
  .A2({ S22359 }),
  .A3({ S18113 }),
  .ZN({ S22360 })
);
AND2_X1 #() 
AND2_X1_235_ (
  .A1({ S22360 }),
  .A2({ S22357 }),
  .ZN({ S25957[1052] })
);
NAND2_X1 #() 
NAND2_X1_3813_ (
  .A1({ S19952 }),
  .A2({ S19953 }),
  .ZN({ S25957[1243] })
);
NAND2_X1 #() 
NAND2_X1_3814_ (
  .A1({ S19945 }),
  .A2({ S19937 }),
  .ZN({ S25957[1275] })
);
INV_X1 #() 
INV_X1_1266_ (
  .A({ S25957[1275] }),
  .ZN({ S22361 })
);
NOR2_X1 #() 
NOR2_X1_969_ (
  .A1({ S22159 }),
  .A2({ S25957[1171] }),
  .ZN({ S22362 })
);
AOI21_X1 #() 
AOI21_X1_2059_ (
  .A({ S22228 }),
  .B1({ S22362 }),
  .B2({ S22191 }),
  .ZN({ S22363 })
);
NAND2_X1 #() 
NAND2_X1_3815_ (
  .A1({ S22323 }),
  .A2({ S22200 }),
  .ZN({ S22364 })
);
NAND2_X1 #() 
NAND2_X1_3816_ (
  .A1({ S22364 }),
  .A2({ S22051 }),
  .ZN({ S22365 })
);
INV_X1 #() 
INV_X1_1267_ (
  .A({ S22365 }),
  .ZN({ S22366 })
);
OAI21_X1 #() 
OAI21_X1_1949_ (
  .A({ S22366 }),
  .B1({ S22363 }),
  .B2({ S9119 }),
  .ZN({ S22367 })
);
OAI21_X1 #() 
OAI21_X1_1950_ (
  .A({ S22154 }),
  .B1({ S22048 }),
  .B2({ S25957[1171] }),
  .ZN({ S22368 })
);
NAND2_X1 #() 
NAND2_X1_3817_ (
  .A1({ S22368 }),
  .A2({ S25957[1172] }),
  .ZN({ S22369 })
);
AOI21_X1 #() 
AOI21_X1_2060_ (
  .A({ S25957[1171] }),
  .B1({ S22055 }),
  .B2({ S20616 }),
  .ZN({ S22370 })
);
AOI21_X1 #() 
AOI21_X1_2061_ (
  .A({ S25957[1172] }),
  .B1({ S22370 }),
  .B2({ S22037 }),
  .ZN({ S22371 })
);
OAI21_X1 #() 
OAI21_X1_1951_ (
  .A({ S22371 }),
  .B1({ S50 }),
  .B2({ S22302 }),
  .ZN({ S22372 })
);
NAND2_X1 #() 
NAND2_X1_3818_ (
  .A1({ S22369 }),
  .A2({ S22372 }),
  .ZN({ S22373 })
);
NAND2_X1 #() 
NAND2_X1_3819_ (
  .A1({ S22373 }),
  .A2({ S25957[1173] }),
  .ZN({ S22374 })
);
AOI21_X1 #() 
AOI21_X1_2062_ (
  .A({ S22094 }),
  .B1({ S22374 }),
  .B2({ S22367 }),
  .ZN({ S22375 })
);
NAND2_X1 #() 
NAND2_X1_3820_ (
  .A1({ S22101 }),
  .A2({ S22337 }),
  .ZN({ S22376 })
);
NAND3_X1 #() 
NAND3_X1_4045_ (
  .A1({ S22065 }),
  .A2({ S22035 }),
  .A3({ S50 }),
  .ZN({ S22377 })
);
NOR2_X1 #() 
NOR2_X1_970_ (
  .A1({ S22377 }),
  .A2({ S9119 }),
  .ZN({ S22378 })
);
NOR2_X1 #() 
NOR2_X1_971_ (
  .A1({ S22378 }),
  .A2({ S25957[1173] }),
  .ZN({ S22379 })
);
NAND2_X1 #() 
NAND2_X1_3821_ (
  .A1({ S22376 }),
  .A2({ S22379 }),
  .ZN({ S22380 })
);
AOI21_X1 #() 
AOI21_X1_2063_ (
  .A({ S22174 }),
  .B1({ S22130 }),
  .B2({ S22129 }),
  .ZN({ S22381 })
);
NAND3_X1 #() 
NAND3_X1_4046_ (
  .A1({ S22095 }),
  .A2({ S50 }),
  .A3({ S22037 }),
  .ZN({ S22382 })
);
NAND2_X1 #() 
NAND2_X1_3822_ (
  .A1({ S22231 }),
  .A2({ S22076 }),
  .ZN({ S22383 })
);
NAND2_X1 #() 
NAND2_X1_3823_ (
  .A1({ S22383 }),
  .A2({ S22382 }),
  .ZN({ S22384 })
);
NAND2_X1 #() 
NAND2_X1_3824_ (
  .A1({ S22384 }),
  .A2({ S9119 }),
  .ZN({ S22385 })
);
OAI211_X1 #() 
OAI211_X1_1317_ (
  .A({ S25957[1173] }),
  .B({ S22385 }),
  .C1({ S22381 }),
  .C2({ S9119 }),
  .ZN({ S22386 })
);
AOI21_X1 #() 
AOI21_X1_2064_ (
  .A({ S25957[1175] }),
  .B1({ S22386 }),
  .B2({ S22380 }),
  .ZN({ S22387 })
);
OAI21_X1 #() 
OAI21_X1_1952_ (
  .A({ S25957[1174] }),
  .B1({ S22375 }),
  .B2({ S22387 }),
  .ZN({ S22388 })
);
NAND2_X1 #() 
NAND2_X1_3825_ (
  .A1({ S22296 }),
  .A2({ S22168 }),
  .ZN({ S22389 })
);
AOI22_X1 #() 
AOI22_X1_430_ (
  .A1({ S22389 }),
  .A2({ S25957[1171] }),
  .B1({ S22088 }),
  .B2({ S82 }),
  .ZN({ S22390 })
);
OAI211_X1 #() 
OAI211_X1_1318_ (
  .A({ S25957[1172] }),
  .B({ S22311 }),
  .C1({ S22084 }),
  .C2({ S50 }),
  .ZN({ S22391 })
);
OAI211_X1 #() 
OAI211_X1_1319_ (
  .A({ S22391 }),
  .B({ S22051 }),
  .C1({ S22390 }),
  .C2({ S25957[1172] }),
  .ZN({ S22392 })
);
NAND2_X1 #() 
NAND2_X1_3826_ (
  .A1({ S22134 }),
  .A2({ S22086 }),
  .ZN({ S22393 })
);
NAND2_X1 #() 
NAND2_X1_3827_ (
  .A1({ S22393 }),
  .A2({ S50 }),
  .ZN({ S22394 })
);
OAI211_X1 #() 
OAI211_X1_1320_ (
  .A({ S22394 }),
  .B({ S25957[1172] }),
  .C1({ S22329 }),
  .C2({ S22187 }),
  .ZN({ S22395 })
);
OR2_X1 #() 
OR2_X1_57_ (
  .A1({ S22082 }),
  .A2({ S22325 }),
  .ZN({ S22396 })
);
NAND2_X1 #() 
NAND2_X1_3828_ (
  .A1({ S25957[1169] }),
  .A2({ S25957[1171] }),
  .ZN({ S22397 })
);
INV_X1 #() 
INV_X1_1268_ (
  .A({ S22397 }),
  .ZN({ S22398 })
);
NAND3_X1 #() 
NAND3_X1_4047_ (
  .A1({ S22398 }),
  .A2({ S22036 }),
  .A3({ S22086 }),
  .ZN({ S22399 })
);
AND2_X1 #() 
AND2_X1_236_ (
  .A1({ S22399 }),
  .A2({ S9119 }),
  .ZN({ S22400 })
);
NAND2_X1 #() 
NAND2_X1_3829_ (
  .A1({ S22400 }),
  .A2({ S22396 }),
  .ZN({ S22401 })
);
NAND3_X1 #() 
NAND3_X1_4048_ (
  .A1({ S22401 }),
  .A2({ S22395 }),
  .A3({ S25957[1173] }),
  .ZN({ S22402 })
);
AOI21_X1 #() 
AOI21_X1_2065_ (
  .A({ S22094 }),
  .B1({ S22392 }),
  .B2({ S22402 }),
  .ZN({ S22403 })
);
OAI211_X1 #() 
OAI211_X1_1321_ (
  .A({ S25957[1171] }),
  .B({ S82 }),
  .C1({ S22035 }),
  .C2({ S25957[1170] }),
  .ZN({ S22404 })
);
NAND3_X1 #() 
NAND3_X1_4049_ (
  .A1({ S22270 }),
  .A2({ S22404 }),
  .A3({ S25957[1172] }),
  .ZN({ S22405 })
);
OAI211_X1 #() 
OAI211_X1_1322_ (
  .A({ S22036 }),
  .B({ S25957[1171] }),
  .C1({ S22035 }),
  .C2({ S25957[1170] }),
  .ZN({ S22406 })
);
OAI211_X1 #() 
OAI211_X1_1323_ (
  .A({ S22406 }),
  .B({ S9119 }),
  .C1({ S22082 }),
  .C2({ S22087 }),
  .ZN({ S22407 })
);
NAND3_X1 #() 
NAND3_X1_4050_ (
  .A1({ S22407 }),
  .A2({ S22405 }),
  .A3({ S22051 }),
  .ZN({ S22408 })
);
NAND2_X1 #() 
NAND2_X1_3830_ (
  .A1({ S22397 }),
  .A2({ S25957[1170] }),
  .ZN({ S22409 })
);
NAND2_X1 #() 
NAND2_X1_3831_ (
  .A1({ S22409 }),
  .A2({ S22203 }),
  .ZN({ S22410 })
);
NAND3_X1 #() 
NAND3_X1_4051_ (
  .A1({ S22410 }),
  .A2({ S9119 }),
  .A3({ S25957[1168] }),
  .ZN({ S22411 })
);
NAND2_X1 #() 
NAND2_X1_3832_ (
  .A1({ S22187 }),
  .A2({ S25957[1172] }),
  .ZN({ S22412 })
);
OAI211_X1 #() 
OAI211_X1_1324_ (
  .A({ S22411 }),
  .B({ S25957[1173] }),
  .C1({ S22412 }),
  .C2({ S22362 }),
  .ZN({ S22413 })
);
AND3_X1 #() 
AND3_X1_144_ (
  .A1({ S22413 }),
  .A2({ S22408 }),
  .A3({ S22094 }),
  .ZN({ S22414 })
);
OAI21_X1 #() 
OAI21_X1_1953_ (
  .A({ S7741 }),
  .B1({ S22403 }),
  .B2({ S22414 }),
  .ZN({ S22415 })
);
NAND3_X1 #() 
NAND3_X1_4052_ (
  .A1({ S22388 }),
  .A2({ S22415 }),
  .A3({ S22361 }),
  .ZN({ S22416 })
);
NAND3_X1 #() 
NAND3_X1_4053_ (
  .A1({ S22224 }),
  .A2({ S50 }),
  .A3({ S22191 }),
  .ZN({ S22417 })
);
NAND2_X1 #() 
NAND2_X1_3833_ (
  .A1({ S22417 }),
  .A2({ S22227 }),
  .ZN({ S22418 })
);
AOI21_X1 #() 
AOI21_X1_2066_ (
  .A({ S22365 }),
  .B1({ S22418 }),
  .B2({ S25957[1172] }),
  .ZN({ S22419 })
);
AOI21_X1 #() 
AOI21_X1_2067_ (
  .A({ S22051 }),
  .B1({ S22369 }),
  .B2({ S22372 }),
  .ZN({ S22420 })
);
OAI21_X1 #() 
OAI21_X1_1954_ (
  .A({ S25957[1174] }),
  .B1({ S22419 }),
  .B2({ S22420 }),
  .ZN({ S22421 })
);
NAND2_X1 #() 
NAND2_X1_3834_ (
  .A1({ S22392 }),
  .A2({ S22402 }),
  .ZN({ S22422 })
);
NAND2_X1 #() 
NAND2_X1_3835_ (
  .A1({ S22422 }),
  .A2({ S7741 }),
  .ZN({ S22423 })
);
NAND3_X1 #() 
NAND3_X1_4054_ (
  .A1({ S22423 }),
  .A2({ S22421 }),
  .A3({ S25957[1175] }),
  .ZN({ S22424 })
);
AND2_X1 #() 
AND2_X1_237_ (
  .A1({ S22386 }),
  .A2({ S22380 }),
  .ZN({ S22425 })
);
NAND3_X1 #() 
NAND3_X1_4055_ (
  .A1({ S22413 }),
  .A2({ S22408 }),
  .A3({ S7741 }),
  .ZN({ S22426 })
);
OAI211_X1 #() 
OAI211_X1_1325_ (
  .A({ S22094 }),
  .B({ S22426 }),
  .C1({ S22425 }),
  .C2({ S7741 }),
  .ZN({ S22427 })
);
NAND3_X1 #() 
NAND3_X1_4056_ (
  .A1({ S22424 }),
  .A2({ S22427 }),
  .A3({ S25957[1275] }),
  .ZN({ S22428 })
);
NAND3_X1 #() 
NAND3_X1_4057_ (
  .A1({ S22416 }),
  .A2({ S22428 }),
  .A3({ S25957[1243] }),
  .ZN({ S22429 })
);
INV_X1 #() 
INV_X1_1269_ (
  .A({ S25957[1243] }),
  .ZN({ S22430 })
);
NAND3_X1 #() 
NAND3_X1_4058_ (
  .A1({ S22424 }),
  .A2({ S22427 }),
  .A3({ S22361 }),
  .ZN({ S22431 })
);
NAND3_X1 #() 
NAND3_X1_4059_ (
  .A1({ S22388 }),
  .A2({ S22415 }),
  .A3({ S25957[1275] }),
  .ZN({ S22432 })
);
NAND3_X1 #() 
NAND3_X1_4060_ (
  .A1({ S22432 }),
  .A2({ S22431 }),
  .A3({ S22430 }),
  .ZN({ S22433 })
);
NAND3_X1 #() 
NAND3_X1_4061_ (
  .A1({ S22429 }),
  .A2({ S22433 }),
  .A3({ S25956[27] }),
  .ZN({ S22434 })
);
NAND3_X1 #() 
NAND3_X1_4062_ (
  .A1({ S22416 }),
  .A2({ S22428 }),
  .A3({ S22430 }),
  .ZN({ S22435 })
);
NAND3_X1 #() 
NAND3_X1_4063_ (
  .A1({ S22432 }),
  .A2({ S22431 }),
  .A3({ S25957[1243] }),
  .ZN({ S22436 })
);
NAND3_X1 #() 
NAND3_X1_4064_ (
  .A1({ S22435 }),
  .A2({ S22436 }),
  .A3({ S18124 }),
  .ZN({ S22437 })
);
NAND2_X1 #() 
NAND2_X1_3836_ (
  .A1({ S22434 }),
  .A2({ S22437 }),
  .ZN({ S83 })
);
AND2_X1 #() 
AND2_X1_238_ (
  .A1({ S22437 }),
  .A2({ S22434 }),
  .ZN({ S25957[1051] })
);
NOR2_X1 #() 
NOR2_X1_972_ (
  .A1({ S20010 }),
  .A2({ S20014 }),
  .ZN({ S25957[1240] })
);
NAND2_X1 #() 
NAND2_X1_3837_ (
  .A1({ S20013 }),
  .A2({ S20012 }),
  .ZN({ S25957[1272] })
);
INV_X1 #() 
INV_X1_1270_ (
  .A({ S25957[1272] }),
  .ZN({ S22438 })
);
AOI21_X1 #() 
AOI21_X1_2068_ (
  .A({ S25957[1171] }),
  .B1({ S22164 }),
  .B2({ S22134 }),
  .ZN({ S22439 })
);
NAND3_X1 #() 
NAND3_X1_4065_ (
  .A1({ S22162 }),
  .A2({ S22052 }),
  .A3({ S22037 }),
  .ZN({ S22440 })
);
INV_X1 #() 
INV_X1_1271_ (
  .A({ S22440 }),
  .ZN({ S22441 })
);
OAI21_X1 #() 
OAI21_X1_1955_ (
  .A({ S25957[1172] }),
  .B1({ S22441 }),
  .B2({ S22439 }),
  .ZN({ S22442 })
);
NAND2_X1 #() 
NAND2_X1_3838_ (
  .A1({ S22095 }),
  .A2({ S50 }),
  .ZN({ S22443 })
);
NAND2_X1 #() 
NAND2_X1_3839_ (
  .A1({ S22443 }),
  .A2({ S22119 }),
  .ZN({ S22444 })
);
OAI21_X1 #() 
OAI21_X1_1956_ (
  .A({ S9119 }),
  .B1({ S22444 }),
  .B2({ S22253 }),
  .ZN({ S22445 })
);
NAND3_X1 #() 
NAND3_X1_4066_ (
  .A1({ S22442 }),
  .A2({ S22051 }),
  .A3({ S22445 }),
  .ZN({ S22446 })
);
NAND2_X1 #() 
NAND2_X1_3840_ (
  .A1({ S22245 }),
  .A2({ S22122 }),
  .ZN({ S22447 })
);
NAND3_X1 #() 
NAND3_X1_4067_ (
  .A1({ S22447 }),
  .A2({ S9119 }),
  .A3({ S22038 }),
  .ZN({ S22448 })
);
NAND2_X1 #() 
NAND2_X1_3841_ (
  .A1({ S22162 }),
  .A2({ S22052 }),
  .ZN({ S22449 })
);
AOI21_X1 #() 
AOI21_X1_2069_ (
  .A({ S9119 }),
  .B1({ S22335 }),
  .B2({ S22449 }),
  .ZN({ S22450 })
);
NOR2_X1 #() 
NOR2_X1_973_ (
  .A1({ S22450 }),
  .A2({ S22051 }),
  .ZN({ S22451 })
);
NAND2_X1 #() 
NAND2_X1_3842_ (
  .A1({ S22451 }),
  .A2({ S22448 }),
  .ZN({ S22452 })
);
NAND3_X1 #() 
NAND3_X1_4068_ (
  .A1({ S22452 }),
  .A2({ S22446 }),
  .A3({ S25957[1174] }),
  .ZN({ S22453 })
);
AOI22_X1 #() 
AOI22_X1_431_ (
  .A1({ S22187 }),
  .A2({ S22377 }),
  .B1({ S22122 }),
  .B2({ S20616 }),
  .ZN({ S22454 })
);
AOI21_X1 #() 
AOI21_X1_2070_ (
  .A({ S25957[1172] }),
  .B1({ S25957[1171] }),
  .B2({ S22046 }),
  .ZN({ S22455 })
);
NAND3_X1 #() 
NAND3_X1_4069_ (
  .A1({ S22455 }),
  .A2({ S22045 }),
  .A3({ S22257 }),
  .ZN({ S22456 })
);
OAI21_X1 #() 
OAI21_X1_1957_ (
  .A({ S22456 }),
  .B1({ S22454 }),
  .B2({ S9119 }),
  .ZN({ S22457 })
);
NAND2_X1 #() 
NAND2_X1_3843_ (
  .A1({ S22457 }),
  .A2({ S25957[1173] }),
  .ZN({ S22458 })
);
NAND4_X1 #() 
NAND4_X1_444_ (
  .A1({ S22065 }),
  .A2({ S22152 }),
  .A3({ S50 }),
  .A4({ S82 }),
  .ZN({ S22459 })
);
AOI21_X1 #() 
AOI21_X1_2071_ (
  .A({ S25957[1172] }),
  .B1({ S22459 }),
  .B2({ S22383 }),
  .ZN({ S22460 })
);
INV_X1 #() 
INV_X1_1272_ (
  .A({ S22460 }),
  .ZN({ S22461 })
);
AOI21_X1 #() 
AOI21_X1_2072_ (
  .A({ S25957[1173] }),
  .B1({ S22330 }),
  .B2({ S22163 }),
  .ZN({ S22462 })
);
AOI21_X1 #() 
AOI21_X1_2073_ (
  .A({ S25957[1174] }),
  .B1({ S22461 }),
  .B2({ S22462 }),
  .ZN({ S22463 })
);
NAND2_X1 #() 
NAND2_X1_3844_ (
  .A1({ S22458 }),
  .A2({ S22463 }),
  .ZN({ S22464 })
);
NAND3_X1 #() 
NAND3_X1_4070_ (
  .A1({ S22453 }),
  .A2({ S22464 }),
  .A3({ S25957[1175] }),
  .ZN({ S22465 })
);
NAND2_X1 #() 
NAND2_X1_3845_ (
  .A1({ S22114 }),
  .A2({ S22230 }),
  .ZN({ S22466 })
);
OAI21_X1 #() 
OAI21_X1_1958_ (
  .A({ S25957[1172] }),
  .B1({ S22466 }),
  .B2({ S22160 }),
  .ZN({ S22467 })
);
NOR2_X1 #() 
NOR2_X1_974_ (
  .A1({ S22325 }),
  .A2({ S22167 }),
  .ZN({ S22468 })
);
OAI21_X1 #() 
OAI21_X1_1959_ (
  .A({ S9119 }),
  .B1({ S22253 }),
  .B2({ S22468 }),
  .ZN({ S22469 })
);
NAND3_X1 #() 
NAND3_X1_4071_ (
  .A1({ S22469 }),
  .A2({ S22051 }),
  .A3({ S22467 }),
  .ZN({ S22470 })
);
OAI21_X1 #() 
OAI21_X1_1960_ (
  .A({ S25957[1171] }),
  .B1({ S22082 }),
  .B2({ S22043 }),
  .ZN({ S22471 })
);
NOR2_X1 #() 
NOR2_X1_975_ (
  .A1({ S22370 }),
  .A2({ S9119 }),
  .ZN({ S22472 })
);
NAND2_X1 #() 
NAND2_X1_3846_ (
  .A1({ S22471 }),
  .A2({ S22472 }),
  .ZN({ S22473 })
);
NOR2_X1 #() 
NOR2_X1_976_ (
  .A1({ S22041 }),
  .A2({ S25957[1172] }),
  .ZN({ S22474 })
);
NAND2_X1 #() 
NAND2_X1_3847_ (
  .A1({ S22196 }),
  .A2({ S22474 }),
  .ZN({ S22475 })
);
NAND3_X1 #() 
NAND3_X1_4072_ (
  .A1({ S22475 }),
  .A2({ S22473 }),
  .A3({ S25957[1173] }),
  .ZN({ S22476 })
);
NAND3_X1 #() 
NAND3_X1_4073_ (
  .A1({ S22476 }),
  .A2({ S22470 }),
  .A3({ S25957[1174] }),
  .ZN({ S22477 })
);
NOR2_X1 #() 
NOR2_X1_977_ (
  .A1({ S22084 }),
  .A2({ S50 }),
  .ZN({ S22478 })
);
AOI21_X1 #() 
AOI21_X1_2074_ (
  .A({ S25957[1171] }),
  .B1({ S22296 }),
  .B2({ S22168 }),
  .ZN({ S22479 })
);
OAI21_X1 #() 
OAI21_X1_1961_ (
  .A({ S22051 }),
  .B1({ S22478 }),
  .B2({ S22479 }),
  .ZN({ S22480 })
);
OAI21_X1 #() 
OAI21_X1_1962_ (
  .A({ S22154 }),
  .B1({ S22053 }),
  .B2({ S22247 }),
  .ZN({ S22481 })
);
AOI21_X1 #() 
AOI21_X1_2075_ (
  .A({ S9119 }),
  .B1({ S22481 }),
  .B2({ S25957[1173] }),
  .ZN({ S22482 })
);
NAND2_X1 #() 
NAND2_X1_3848_ (
  .A1({ S22480 }),
  .A2({ S22482 }),
  .ZN({ S22483 })
);
NAND2_X1 #() 
NAND2_X1_3849_ (
  .A1({ S22177 }),
  .A2({ S22261 }),
  .ZN({ S22484 })
);
NAND2_X1 #() 
NAND2_X1_3850_ (
  .A1({ S22484 }),
  .A2({ S25957[1173] }),
  .ZN({ S22485 })
);
NAND3_X1 #() 
NAND3_X1_4074_ (
  .A1({ S22168 }),
  .A2({ S25957[1171] }),
  .A3({ S82 }),
  .ZN({ S22486 })
);
OAI211_X1 #() 
OAI211_X1_1326_ (
  .A({ S22051 }),
  .B({ S22486 }),
  .C1({ S22045 }),
  .C2({ S22190 }),
  .ZN({ S22487 })
);
NAND3_X1 #() 
NAND3_X1_4075_ (
  .A1({ S22485 }),
  .A2({ S9119 }),
  .A3({ S22487 }),
  .ZN({ S22488 })
);
NAND3_X1 #() 
NAND3_X1_4076_ (
  .A1({ S22483 }),
  .A2({ S7741 }),
  .A3({ S22488 }),
  .ZN({ S22489 })
);
NAND3_X1 #() 
NAND3_X1_4077_ (
  .A1({ S22489 }),
  .A2({ S22477 }),
  .A3({ S22094 }),
  .ZN({ S22490 })
);
NAND3_X1 #() 
NAND3_X1_4078_ (
  .A1({ S22465 }),
  .A2({ S22490 }),
  .A3({ S22438 }),
  .ZN({ S22491 })
);
OAI211_X1 #() 
OAI211_X1_1327_ (
  .A({ S22456 }),
  .B({ S25957[1173] }),
  .C1({ S22454 }),
  .C2({ S9119 }),
  .ZN({ S22492 })
);
AND2_X1 #() 
AND2_X1_239_ (
  .A1({ S22330 }),
  .A2({ S22163 }),
  .ZN({ S22493 })
);
OAI21_X1 #() 
OAI21_X1_1963_ (
  .A({ S22051 }),
  .B1({ S22493 }),
  .B2({ S22460 }),
  .ZN({ S22494 })
);
NAND3_X1 #() 
NAND3_X1_4079_ (
  .A1({ S22494 }),
  .A2({ S7741 }),
  .A3({ S22492 }),
  .ZN({ S22495 })
);
INV_X1 #() 
INV_X1_1273_ (
  .A({ S22448 }),
  .ZN({ S22496 })
);
OAI21_X1 #() 
OAI21_X1_1964_ (
  .A({ S25957[1173] }),
  .B1({ S22496 }),
  .B2({ S22450 }),
  .ZN({ S22497 })
);
NAND3_X1 #() 
NAND3_X1_4080_ (
  .A1({ S22303 }),
  .A2({ S25957[1172] }),
  .A3({ S22440 }),
  .ZN({ S22498 })
);
NAND4_X1 #() 
NAND4_X1_445_ (
  .A1({ S22328 }),
  .A2({ S22443 }),
  .A3({ S9119 }),
  .A4({ S22119 }),
  .ZN({ S22499 })
);
NAND3_X1 #() 
NAND3_X1_4081_ (
  .A1({ S22498 }),
  .A2({ S22499 }),
  .A3({ S22051 }),
  .ZN({ S22500 })
);
NAND3_X1 #() 
NAND3_X1_4082_ (
  .A1({ S22497 }),
  .A2({ S22500 }),
  .A3({ S25957[1174] }),
  .ZN({ S22501 })
);
NAND3_X1 #() 
NAND3_X1_4083_ (
  .A1({ S22501 }),
  .A2({ S22495 }),
  .A3({ S25957[1175] }),
  .ZN({ S22502 })
);
AND2_X1 #() 
AND2_X1_240_ (
  .A1({ S22487 }),
  .A2({ S9119 }),
  .ZN({ S22503 })
);
AOI22_X1 #() 
AOI22_X1_432_ (
  .A1({ S22503 }),
  .A2({ S22485 }),
  .B1({ S22480 }),
  .B2({ S22482 }),
  .ZN({ S22504 })
);
AOI22_X1 #() 
AOI22_X1_433_ (
  .A1({ S22196 }),
  .A2({ S22474 }),
  .B1({ S22471 }),
  .B2({ S22472 }),
  .ZN({ S22505 })
);
INV_X1 #() 
INV_X1_1274_ (
  .A({ S22468 }),
  .ZN({ S22506 })
);
NAND3_X1 #() 
NAND3_X1_4084_ (
  .A1({ S22328 }),
  .A2({ S22506 }),
  .A3({ S9119 }),
  .ZN({ S22507 })
);
NAND3_X1 #() 
NAND3_X1_4085_ (
  .A1({ S22165 }),
  .A2({ S25957[1172] }),
  .A3({ S22230 }),
  .ZN({ S22508 })
);
NAND3_X1 #() 
NAND3_X1_4086_ (
  .A1({ S22507 }),
  .A2({ S22051 }),
  .A3({ S22508 }),
  .ZN({ S22509 })
);
OAI211_X1 #() 
OAI211_X1_1328_ (
  .A({ S22509 }),
  .B({ S25957[1174] }),
  .C1({ S22505 }),
  .C2({ S22051 }),
  .ZN({ S22510 })
);
OAI211_X1 #() 
OAI211_X1_1329_ (
  .A({ S22510 }),
  .B({ S22094 }),
  .C1({ S22504 }),
  .C2({ S25957[1174] }),
  .ZN({ S22511 })
);
NAND3_X1 #() 
NAND3_X1_4087_ (
  .A1({ S22511 }),
  .A2({ S22502 }),
  .A3({ S25957[1272] }),
  .ZN({ S22512 })
);
NAND3_X1 #() 
NAND3_X1_4088_ (
  .A1({ S22512 }),
  .A2({ S22491 }),
  .A3({ S25957[1240] }),
  .ZN({ S22513 })
);
INV_X1 #() 
INV_X1_1275_ (
  .A({ S25957[1240] }),
  .ZN({ S22514 })
);
NAND3_X1 #() 
NAND3_X1_4089_ (
  .A1({ S22511 }),
  .A2({ S22502 }),
  .A3({ S22438 }),
  .ZN({ S22515 })
);
NAND3_X1 #() 
NAND3_X1_4090_ (
  .A1({ S22465 }),
  .A2({ S22490 }),
  .A3({ S25957[1272] }),
  .ZN({ S22516 })
);
NAND3_X1 #() 
NAND3_X1_4091_ (
  .A1({ S22515 }),
  .A2({ S22516 }),
  .A3({ S22514 }),
  .ZN({ S22517 })
);
NAND3_X1 #() 
NAND3_X1_4092_ (
  .A1({ S22513 }),
  .A2({ S22517 }),
  .A3({ S25956[24] }),
  .ZN({ S22518 })
);
NAND3_X1 #() 
NAND3_X1_4093_ (
  .A1({ S22512 }),
  .A2({ S22491 }),
  .A3({ S22514 }),
  .ZN({ S22519 })
);
NAND3_X1 #() 
NAND3_X1_4094_ (
  .A1({ S22515 }),
  .A2({ S22516 }),
  .A3({ S25957[1240] }),
  .ZN({ S22520 })
);
NAND3_X1 #() 
NAND3_X1_4095_ (
  .A1({ S22519 }),
  .A2({ S22520 }),
  .A3({ S18242 }),
  .ZN({ S22521 })
);
AND2_X1 #() 
AND2_X1_241_ (
  .A1({ S22521 }),
  .A2({ S22518 }),
  .ZN({ S25957[1048] })
);
NAND2_X1 #() 
NAND2_X1_3851_ (
  .A1({ S20064 }),
  .A2({ S20063 }),
  .ZN({ S25957[1273] })
);
INV_X1 #() 
INV_X1_1276_ (
  .A({ S25957[1273] }),
  .ZN({ S22522 })
);
AOI21_X1 #() 
AOI21_X1_2076_ (
  .A({ S9119 }),
  .B1({ S22399 }),
  .B2({ S22316 }),
  .ZN({ S22523 })
);
OAI21_X1 #() 
OAI21_X1_1965_ (
  .A({ S25957[1173] }),
  .B1({ S22101 }),
  .B2({ S22523 }),
  .ZN({ S22524 })
);
NAND3_X1 #() 
NAND3_X1_4096_ (
  .A1({ S22069 }),
  .A2({ S25957[1172] }),
  .A3({ S22311 }),
  .ZN({ S22525 })
);
INV_X1 #() 
INV_X1_1277_ (
  .A({ S22083 }),
  .ZN({ S22526 })
);
OAI21_X1 #() 
OAI21_X1_1966_ (
  .A({ S22081 }),
  .B1({ S22115 }),
  .B2({ S22526 }),
  .ZN({ S22527 })
);
NAND3_X1 #() 
NAND3_X1_4097_ (
  .A1({ S22527 }),
  .A2({ S22525 }),
  .A3({ S22051 }),
  .ZN({ S22528 })
);
NAND3_X1 #() 
NAND3_X1_4098_ (
  .A1({ S22524 }),
  .A2({ S7741 }),
  .A3({ S22528 }),
  .ZN({ S22529 })
);
AOI21_X1 #() 
AOI21_X1_2077_ (
  .A({ S22096 }),
  .B1({ S22077 }),
  .B2({ S82 }),
  .ZN({ S22530 })
);
OAI21_X1 #() 
OAI21_X1_1967_ (
  .A({ S25957[1172] }),
  .B1({ S22087 }),
  .B2({ S22108 }),
  .ZN({ S22531 })
);
NOR2_X1 #() 
NOR2_X1_978_ (
  .A1({ S22242 }),
  .A2({ S22068 }),
  .ZN({ S22532 })
);
AOI21_X1 #() 
AOI21_X1_2078_ (
  .A({ S22051 }),
  .B1({ S22240 }),
  .B2({ S22532 }),
  .ZN({ S22533 })
);
OAI21_X1 #() 
OAI21_X1_1968_ (
  .A({ S22533 }),
  .B1({ S22530 }),
  .B2({ S22531 }),
  .ZN({ S22534 })
);
AOI22_X1 #() 
AOI22_X1_434_ (
  .A1({ S22099 }),
  .A2({ S22086 }),
  .B1({ S22277 }),
  .B2({ S22397 }),
  .ZN({ S22535 })
);
OAI21_X1 #() 
OAI21_X1_1969_ (
  .A({ S25957[1172] }),
  .B1({ S22169 }),
  .B2({ S22071 }),
  .ZN({ S22536 })
);
INV_X1 #() 
INV_X1_1278_ (
  .A({ S22099 }),
  .ZN({ S22537 })
);
OAI211_X1 #() 
OAI211_X1_1330_ (
  .A({ S22440 }),
  .B({ S9119 }),
  .C1({ S22537 }),
  .C2({ S22087 }),
  .ZN({ S22538 })
);
OAI211_X1 #() 
OAI211_X1_1331_ (
  .A({ S22538 }),
  .B({ S22051 }),
  .C1({ S22535 }),
  .C2({ S22536 }),
  .ZN({ S22539 })
);
NAND3_X1 #() 
NAND3_X1_4099_ (
  .A1({ S22539 }),
  .A2({ S22534 }),
  .A3({ S25957[1174] }),
  .ZN({ S22540 })
);
NAND3_X1 #() 
NAND3_X1_4100_ (
  .A1({ S22540 }),
  .A2({ S22529 }),
  .A3({ S22094 }),
  .ZN({ S22541 })
);
NOR3_X1 #() 
NOR3_X1_133_ (
  .A1({ S22104 }),
  .A2({ S22295 }),
  .A3({ S25957[1172] }),
  .ZN({ S22542 })
);
NAND2_X1 #() 
NAND2_X1_3852_ (
  .A1({ S25957[1172] }),
  .A2({ S50 }),
  .ZN({ S22543 })
);
NAND3_X1 #() 
NAND3_X1_4101_ (
  .A1({ S25957[1172] }),
  .A2({ S25957[1171] }),
  .A3({ S22095 }),
  .ZN({ S22544 })
);
OAI211_X1 #() 
OAI211_X1_1332_ (
  .A({ S22051 }),
  .B({ S22544 }),
  .C1({ S22165 }),
  .C2({ S22543 }),
  .ZN({ S22545 })
);
NOR3_X1 #() 
NOR3_X1_134_ (
  .A1({ S22082 }),
  .A2({ S22247 }),
  .A3({ S50 }),
  .ZN({ S22546 })
);
NAND3_X1 #() 
NAND3_X1_4102_ (
  .A1({ S22222 }),
  .A2({ S22382 }),
  .A3({ S9119 }),
  .ZN({ S22547 })
);
OAI211_X1 #() 
OAI211_X1_1333_ (
  .A({ S25957[1173] }),
  .B({ S22547 }),
  .C1({ S22111 }),
  .C2({ S22546 }),
  .ZN({ S22548 })
);
OAI211_X1 #() 
OAI211_X1_1334_ (
  .A({ S22548 }),
  .B({ S7741 }),
  .C1({ S22542 }),
  .C2({ S22545 }),
  .ZN({ S22549 })
);
NAND2_X1 #() 
NAND2_X1_3853_ (
  .A1({ S22122 }),
  .A2({ S20616 }),
  .ZN({ S22550 })
);
OAI211_X1 #() 
OAI211_X1_1335_ (
  .A({ S25957[1172] }),
  .B({ S22550 }),
  .C1({ S22269 }),
  .C2({ S22159 }),
  .ZN({ S22551 })
);
NAND3_X1 #() 
NAND3_X1_4103_ (
  .A1({ S22036 }),
  .A2({ S22035 }),
  .A3({ S25957[1171] }),
  .ZN({ S22552 })
);
OAI211_X1 #() 
OAI211_X1_1336_ (
  .A({ S22552 }),
  .B({ S9119 }),
  .C1({ S22377 }),
  .C2({ S22242 }),
  .ZN({ S22553 })
);
NAND3_X1 #() 
NAND3_X1_4104_ (
  .A1({ S22551 }),
  .A2({ S22051 }),
  .A3({ S22553 }),
  .ZN({ S22554 })
);
NAND3_X1 #() 
NAND3_X1_4105_ (
  .A1({ S22115 }),
  .A2({ S22227 }),
  .A3({ S25957[1172] }),
  .ZN({ S22555 })
);
NAND2_X1 #() 
NAND2_X1_3854_ (
  .A1({ S22110 }),
  .A2({ S9119 }),
  .ZN({ S22556 })
);
OAI211_X1 #() 
OAI211_X1_1337_ (
  .A({ S25957[1173] }),
  .B({ S22555 }),
  .C1({ S22556 }),
  .C2({ S22535 }),
  .ZN({ S22557 })
);
NAND3_X1 #() 
NAND3_X1_4106_ (
  .A1({ S22554 }),
  .A2({ S25957[1174] }),
  .A3({ S22557 }),
  .ZN({ S22558 })
);
NAND3_X1 #() 
NAND3_X1_4107_ (
  .A1({ S22549 }),
  .A2({ S25957[1175] }),
  .A3({ S22558 }),
  .ZN({ S22559 })
);
NAND3_X1 #() 
NAND3_X1_4108_ (
  .A1({ S22559 }),
  .A2({ S22541 }),
  .A3({ S22522 }),
  .ZN({ S22560 })
);
NAND2_X1 #() 
NAND2_X1_3855_ (
  .A1({ S22559 }),
  .A2({ S22541 }),
  .ZN({ S22561 })
);
NAND2_X1 #() 
NAND2_X1_3856_ (
  .A1({ S22561 }),
  .A2({ S25957[1273] }),
  .ZN({ S22562 })
);
AOI21_X1 #() 
AOI21_X1_2079_ (
  .A({ S25956[57] }),
  .B1({ S22562 }),
  .B2({ S22560 }),
  .ZN({ S22563 })
);
NAND3_X1 #() 
NAND3_X1_4109_ (
  .A1({ S22559 }),
  .A2({ S22541 }),
  .A3({ S25957[1273] }),
  .ZN({ S22564 })
);
NAND2_X1 #() 
NAND2_X1_3857_ (
  .A1({ S22561 }),
  .A2({ S22522 }),
  .ZN({ S22565 })
);
AOI21_X1 #() 
AOI21_X1_2080_ (
  .A({ S20024 }),
  .B1({ S22565 }),
  .B2({ S22564 }),
  .ZN({ S22566 })
);
OAI21_X1 #() 
OAI21_X1_1970_ (
  .A({ S25957[1177] }),
  .B1({ S22563 }),
  .B2({ S22566 }),
  .ZN({ S22567 })
);
NAND3_X1 #() 
NAND3_X1_4110_ (
  .A1({ S22565 }),
  .A2({ S20024 }),
  .A3({ S22564 }),
  .ZN({ S22568 })
);
NAND3_X1 #() 
NAND3_X1_4111_ (
  .A1({ S22562 }),
  .A2({ S25956[57] }),
  .A3({ S22560 }),
  .ZN({ S22569 })
);
NAND3_X1 #() 
NAND3_X1_4112_ (
  .A1({ S22568 }),
  .A2({ S22569 }),
  .A3({ S21399 }),
  .ZN({ S22570 })
);
NAND2_X1 #() 
NAND2_X1_3858_ (
  .A1({ S22567 }),
  .A2({ S22570 }),
  .ZN({ S25957[1049] })
);
NOR2_X1 #() 
NOR2_X1_979_ (
  .A1({ S20116 }),
  .A2({ S20120 }),
  .ZN({ S25957[1210] })
);
NAND2_X1 #() 
NAND2_X1_3859_ (
  .A1({ S20118 }),
  .A2({ S20119 }),
  .ZN({ S25957[1242] })
);
INV_X1 #() 
INV_X1_1279_ (
  .A({ S25957[1242] }),
  .ZN({ S22571 })
);
NAND2_X1 #() 
NAND2_X1_3860_ (
  .A1({ S20111 }),
  .A2({ S20109 }),
  .ZN({ S25957[1274] })
);
INV_X1 #() 
INV_X1_1280_ (
  .A({ S25957[1274] }),
  .ZN({ S22572 })
);
NOR2_X1 #() 
NOR2_X1_980_ (
  .A1({ S22443 }),
  .A2({ S20616 }),
  .ZN({ S22573 })
);
NOR2_X1 #() 
NOR2_X1_981_ (
  .A1({ S22573 }),
  .A2({ S25957[1172] }),
  .ZN({ S22574 })
);
NAND4_X1 #() 
NAND4_X1_446_ (
  .A1({ S25957[1172] }),
  .A2({ S25957[1171] }),
  .A3({ S22055 }),
  .A4({ S22037 }),
  .ZN({ S22575 })
);
OAI211_X1 #() 
OAI211_X1_1338_ (
  .A({ S22575 }),
  .B({ S25957[1173] }),
  .C1({ S9119 }),
  .C2({ S22377 }),
  .ZN({ S22576 })
);
AOI21_X1 #() 
AOI21_X1_2081_ (
  .A({ S22576 }),
  .B1({ S22574 }),
  .B2({ S22085 }),
  .ZN({ S22577 })
);
NAND3_X1 #() 
NAND3_X1_4113_ (
  .A1({ S22077 }),
  .A2({ S25957[1172] }),
  .A3({ S50 }),
  .ZN({ S22578 })
);
AOI21_X1 #() 
AOI21_X1_2082_ (
  .A({ S25957[1172] }),
  .B1({ S22398 }),
  .B2({ S22086 }),
  .ZN({ S22579 })
);
OAI21_X1 #() 
OAI21_X1_1971_ (
  .A({ S22579 }),
  .B1({ S22302 }),
  .B2({ S25957[1171] }),
  .ZN({ S22580 })
);
NOR2_X1 #() 
NOR2_X1_982_ (
  .A1({ S22068 }),
  .A2({ S9119 }),
  .ZN({ S22581 })
);
AOI21_X1 #() 
AOI21_X1_2083_ (
  .A({ S25957[1173] }),
  .B1({ S22581 }),
  .B2({ S22268 }),
  .ZN({ S22582 })
);
AND3_X1 #() 
AND3_X1_145_ (
  .A1({ S22580 }),
  .A2({ S22578 }),
  .A3({ S22582 }),
  .ZN({ S22583 })
);
OAI21_X1 #() 
OAI21_X1_1972_ (
  .A({ S25957[1174] }),
  .B1({ S22583 }),
  .B2({ S22577 }),
  .ZN({ S22584 })
);
OAI221_X1 #() 
OAI221_X1_113_ (
  .A({ S25957[1172] }),
  .B1({ S22096 }),
  .B2({ S22242 }),
  .C1({ S22082 }),
  .C2({ S22325 }),
  .ZN({ S22585 })
);
OAI211_X1 #() 
OAI211_X1_1339_ (
  .A({ S22275 }),
  .B({ S9119 }),
  .C1({ S22181 }),
  .C2({ S22169 }),
  .ZN({ S22586 })
);
NAND3_X1 #() 
NAND3_X1_4114_ (
  .A1({ S22585 }),
  .A2({ S22586 }),
  .A3({ S25957[1173] }),
  .ZN({ S22587 })
);
NAND2_X1 #() 
NAND2_X1_3861_ (
  .A1({ S22398 }),
  .A2({ S22086 }),
  .ZN({ S22588 })
);
OAI211_X1 #() 
OAI211_X1_1340_ (
  .A({ S25957[1172] }),
  .B({ S22588 }),
  .C1({ S22110 }),
  .C2({ S22043 }),
  .ZN({ S22589 })
);
NAND3_X1 #() 
NAND3_X1_4115_ (
  .A1({ S22196 }),
  .A2({ S9119 }),
  .A3({ S22447 }),
  .ZN({ S22590 })
);
NAND3_X1 #() 
NAND3_X1_4116_ (
  .A1({ S22590 }),
  .A2({ S22051 }),
  .A3({ S22589 }),
  .ZN({ S22591 })
);
NAND3_X1 #() 
NAND3_X1_4117_ (
  .A1({ S22591 }),
  .A2({ S7741 }),
  .A3({ S22587 }),
  .ZN({ S22592 })
);
NAND3_X1 #() 
NAND3_X1_4118_ (
  .A1({ S22584 }),
  .A2({ S22592 }),
  .A3({ S22094 }),
  .ZN({ S22593 })
);
OAI211_X1 #() 
OAI211_X1_1341_ (
  .A({ S22098 }),
  .B({ S25957[1172] }),
  .C1({ S25957[1171] }),
  .C2({ S22078 }),
  .ZN({ S22594 })
);
NAND4_X1 #() 
NAND4_X1_447_ (
  .A1({ S22245 }),
  .A2({ S22114 }),
  .A3({ S22065 }),
  .A4({ S25957[1171] }),
  .ZN({ S22595 })
);
NAND3_X1 #() 
NAND3_X1_4119_ (
  .A1({ S22595 }),
  .A2({ S9119 }),
  .A3({ S22123 }),
  .ZN({ S22596 })
);
NAND3_X1 #() 
NAND3_X1_4120_ (
  .A1({ S22594 }),
  .A2({ S25957[1173] }),
  .A3({ S22596 }),
  .ZN({ S22597 })
);
AND3_X1 #() 
AND3_X1_146_ (
  .A1({ S22245 }),
  .A2({ S22134 }),
  .A3({ S25957[1171] }),
  .ZN({ S22598 })
);
NOR2_X1 #() 
NOR2_X1_983_ (
  .A1({ S22055 }),
  .A2({ S25957[1171] }),
  .ZN({ S22599 })
);
OAI221_X1 #() 
OAI221_X1_114_ (
  .A({ S22051 }),
  .B1({ S22126 }),
  .B2({ S22599 }),
  .C1({ S22598 }),
  .C2({ S22248 }),
  .ZN({ S22600 })
);
NAND3_X1 #() 
NAND3_X1_4121_ (
  .A1({ S22597 }),
  .A2({ S25957[1174] }),
  .A3({ S22600 }),
  .ZN({ S22601 })
);
OAI211_X1 #() 
OAI211_X1_1342_ (
  .A({ S22275 }),
  .B({ S9119 }),
  .C1({ S50 }),
  .C2({ S22076 }),
  .ZN({ S22602 })
);
AOI21_X1 #() 
AOI21_X1_2084_ (
  .A({ S9119 }),
  .B1({ S22095 }),
  .B2({ S50 }),
  .ZN({ S22603 })
);
AOI21_X1 #() 
AOI21_X1_2085_ (
  .A({ S25957[1173] }),
  .B1({ S22603 }),
  .B2({ S22588 }),
  .ZN({ S22604 })
);
NAND3_X1 #() 
NAND3_X1_4122_ (
  .A1({ S22055 }),
  .A2({ S25957[1171] }),
  .A3({ S25957[1168] }),
  .ZN({ S22605 })
);
OAI211_X1 #() 
OAI211_X1_1343_ (
  .A({ S25957[1172] }),
  .B({ S22605 }),
  .C1({ S22115 }),
  .C2({ S22526 }),
  .ZN({ S22606 })
);
AOI21_X1 #() 
AOI21_X1_2086_ (
  .A({ S22167 }),
  .B1({ S22409 }),
  .B2({ S22230 }),
  .ZN({ S22607 })
);
AOI21_X1 #() 
AOI21_X1_2087_ (
  .A({ S22051 }),
  .B1({ S22607 }),
  .B2({ S9119 }),
  .ZN({ S22608 })
);
AOI22_X1 #() 
AOI22_X1_435_ (
  .A1({ S22608 }),
  .A2({ S22606 }),
  .B1({ S22602 }),
  .B2({ S22604 }),
  .ZN({ S22609 })
);
AOI21_X1 #() 
AOI21_X1_2088_ (
  .A({ S22094 }),
  .B1({ S22609 }),
  .B2({ S7741 }),
  .ZN({ S22610 })
);
NAND2_X1 #() 
NAND2_X1_3862_ (
  .A1({ S22601 }),
  .A2({ S22610 }),
  .ZN({ S22611 })
);
NAND3_X1 #() 
NAND3_X1_4123_ (
  .A1({ S22593 }),
  .A2({ S22611 }),
  .A3({ S22572 }),
  .ZN({ S22612 })
);
NAND2_X1 #() 
NAND2_X1_3863_ (
  .A1({ S22593 }),
  .A2({ S22611 }),
  .ZN({ S22613 })
);
NAND2_X1 #() 
NAND2_X1_3864_ (
  .A1({ S22613 }),
  .A2({ S25957[1274] }),
  .ZN({ S22614 })
);
NAND3_X1 #() 
NAND3_X1_4124_ (
  .A1({ S22614 }),
  .A2({ S22571 }),
  .A3({ S22612 }),
  .ZN({ S22615 })
);
NAND2_X1 #() 
NAND2_X1_3865_ (
  .A1({ S22613 }),
  .A2({ S22572 }),
  .ZN({ S22616 })
);
NAND3_X1 #() 
NAND3_X1_4125_ (
  .A1({ S22593 }),
  .A2({ S22611 }),
  .A3({ S25957[1274] }),
  .ZN({ S22617 })
);
NAND3_X1 #() 
NAND3_X1_4126_ (
  .A1({ S22616 }),
  .A2({ S25957[1242] }),
  .A3({ S22617 }),
  .ZN({ S22618 })
);
AOI21_X1 #() 
AOI21_X1_2089_ (
  .A({ S25957[1210] }),
  .B1({ S22615 }),
  .B2({ S22618 }),
  .ZN({ S22619 })
);
AND3_X1 #() 
AND3_X1_147_ (
  .A1({ S22618 }),
  .A2({ S22615 }),
  .A3({ S25957[1210] }),
  .ZN({ S22620 })
);
OAI21_X1 #() 
OAI21_X1_1973_ (
  .A({ S25957[1178] }),
  .B1({ S22620 }),
  .B2({ S22619 }),
  .ZN({ S22621 })
);
INV_X1 #() 
INV_X1_1281_ (
  .A({ S25957[1210] }),
  .ZN({ S22622 })
);
AOI21_X1 #() 
AOI21_X1_2090_ (
  .A({ S25957[1242] }),
  .B1({ S22616 }),
  .B2({ S22617 }),
  .ZN({ S22623 })
);
AOI21_X1 #() 
AOI21_X1_2091_ (
  .A({ S22571 }),
  .B1({ S22614 }),
  .B2({ S22612 }),
  .ZN({ S22624 })
);
OAI21_X1 #() 
OAI21_X1_1974_ (
  .A({ S22622 }),
  .B1({ S22623 }),
  .B2({ S22624 }),
  .ZN({ S22625 })
);
NAND3_X1 #() 
NAND3_X1_4127_ (
  .A1({ S22615 }),
  .A2({ S22618 }),
  .A3({ S25957[1210] }),
  .ZN({ S22626 })
);
NAND3_X1 #() 
NAND3_X1_4128_ (
  .A1({ S22625 }),
  .A2({ S21411 }),
  .A3({ S22626 }),
  .ZN({ S22627 })
);
NAND2_X1 #() 
NAND2_X1_3866_ (
  .A1({ S22621 }),
  .A2({ S22627 }),
  .ZN({ S25957[1050] })
);
NAND3_X1 #() 
NAND3_X1_4129_ (
  .A1({ S21263 }),
  .A2({ S21264 }),
  .A3({ S25956[8] }),
  .ZN({ S22628 })
);
NAND3_X1 #() 
NAND3_X1_4130_ (
  .A1({ S21258 }),
  .A2({ S21261 }),
  .A3({ S5639 }),
  .ZN({ S22629 })
);
NAND3_X1 #() 
NAND3_X1_4131_ (
  .A1({ S21314 }),
  .A2({ S21315 }),
  .A3({ S25956[9] }),
  .ZN({ S22630 })
);
NAND3_X1 #() 
NAND3_X1_4132_ (
  .A1({ S21309 }),
  .A2({ S21312 }),
  .A3({ S5628 }),
  .ZN({ S22631 })
);
NAND4_X1 #() 
NAND4_X1_448_ (
  .A1({ S22630 }),
  .A2({ S22631 }),
  .A3({ S22628 }),
  .A4({ S22629 }),
  .ZN({ S22632 })
);
INV_X1 #() 
INV_X1_1282_ (
  .A({ S22632 }),
  .ZN({ S84 })
);
NAND2_X1 #() 
NAND2_X1_3867_ (
  .A1({ S22628 }),
  .A2({ S22629 }),
  .ZN({ S22633 })
);
NAND2_X1 #() 
NAND2_X1_3868_ (
  .A1({ S22630 }),
  .A2({ S22631 }),
  .ZN({ S22634 })
);
NAND2_X1 #() 
NAND2_X1_3869_ (
  .A1({ S22634 }),
  .A2({ S22633 }),
  .ZN({ S85 })
);
XOR2_X1 #() 
XOR2_X1_71_ (
  .A({ S25957[1143] }),
  .B({ S25956[55] }),
  .Z({ S25957[1079] })
);
NAND2_X1 #() 
NAND2_X1_3870_ (
  .A1({ S20941 }),
  .A2({ S20942 }),
  .ZN({ S22635 })
);
NAND2_X1 #() 
NAND2_X1_3871_ (
  .A1({ S21090 }),
  .A2({ S21093 }),
  .ZN({ S22636 })
);
NAND2_X1 #() 
NAND2_X1_3872_ (
  .A1({ S17900 }),
  .A2({ S17933 }),
  .ZN({ S22637 })
);
INV_X1 #() 
INV_X1_1283_ (
  .A({ S22637 }),
  .ZN({ S25957[1226] })
);
NAND3_X1 #() 
NAND3_X1_4133_ (
  .A1({ S21384 }),
  .A2({ S21383 }),
  .A3({ S25957[1226] }),
  .ZN({ S22638 })
);
NAND3_X1 #() 
NAND3_X1_4134_ (
  .A1({ S21381 }),
  .A2({ S21365 }),
  .A3({ S22637 }),
  .ZN({ S22639 })
);
NAND3_X1 #() 
NAND3_X1_4135_ (
  .A1({ S22638 }),
  .A2({ S22639 }),
  .A3({ S5730 }),
  .ZN({ S22640 })
);
NAND3_X1 #() 
NAND3_X1_4136_ (
  .A1({ S21381 }),
  .A2({ S21365 }),
  .A3({ S25957[1226] }),
  .ZN({ S22641 })
);
NAND3_X1 #() 
NAND3_X1_4137_ (
  .A1({ S21384 }),
  .A2({ S21383 }),
  .A3({ S22637 }),
  .ZN({ S22642 })
);
NAND3_X1 #() 
NAND3_X1_4138_ (
  .A1({ S22641 }),
  .A2({ S22642 }),
  .A3({ S25956[10] }),
  .ZN({ S22643 })
);
NAND2_X1 #() 
NAND2_X1_3873_ (
  .A1({ S22640 }),
  .A2({ S22643 }),
  .ZN({ S22644 })
);
NAND2_X1 #() 
NAND2_X1_3874_ (
  .A1({ S22644 }),
  .A2({ S22633 }),
  .ZN({ S22645 })
);
NAND2_X1 #() 
NAND2_X1_3875_ (
  .A1({ S22645 }),
  .A2({ S25957[1033] }),
  .ZN({ S22646 })
);
NAND4_X1 #() 
NAND4_X1_449_ (
  .A1({ S21386 }),
  .A2({ S21389 }),
  .A3({ S22630 }),
  .A4({ S22631 }),
  .ZN({ S22647 })
);
NAND4_X1 #() 
NAND4_X1_450_ (
  .A1({ S22640 }),
  .A2({ S22643 }),
  .A3({ S22628 }),
  .A4({ S22629 }),
  .ZN({ S22648 })
);
NAND3_X1 #() 
NAND3_X1_4139_ (
  .A1({ S22645 }),
  .A2({ S22647 }),
  .A3({ S22648 }),
  .ZN({ S22649 })
);
NAND2_X1 #() 
NAND2_X1_3876_ (
  .A1({ S22649 }),
  .A2({ S25957[1035] }),
  .ZN({ S22650 })
);
OAI21_X1 #() 
OAI21_X1_1975_ (
  .A({ S22650 }),
  .B1({ S25957[1035] }),
  .B2({ S22646 }),
  .ZN({ S22651 })
);
NOR2_X1 #() 
NOR2_X1_984_ (
  .A1({ S22651 }),
  .A2({ S22636 }),
  .ZN({ S22652 })
);
NAND3_X1 #() 
NAND3_X1_4140_ (
  .A1({ S25957[1034] }),
  .A2({ S22633 }),
  .A3({ S22634 }),
  .ZN({ S22653 })
);
NAND2_X1 #() 
NAND2_X1_3877_ (
  .A1({ S85 }),
  .A2({ S22644 }),
  .ZN({ S22654 })
);
NAND2_X1 #() 
NAND2_X1_3878_ (
  .A1({ S22654 }),
  .A2({ S22653 }),
  .ZN({ S22655 })
);
OAI211_X1 #() 
OAI211_X1_1344_ (
  .A({ S22628 }),
  .B({ S22629 }),
  .C1({ S21316 }),
  .C2({ S21313 }),
  .ZN({ S22656 })
);
INV_X1 #() 
INV_X1_1284_ (
  .A({ S22656 }),
  .ZN({ S22657 })
);
NAND2_X1 #() 
NAND2_X1_3879_ (
  .A1({ S22657 }),
  .A2({ S25957[1035] }),
  .ZN({ S22658 })
);
AOI21_X1 #() 
AOI21_X1_2092_ (
  .A({ S25957[1036] }),
  .B1({ S22655 }),
  .B2({ S22658 }),
  .ZN({ S22659 })
);
NAND3_X1 #() 
NAND3_X1_4141_ (
  .A1({ S22633 }),
  .A2({ S22640 }),
  .A3({ S22643 }),
  .ZN({ S22660 })
);
NAND2_X1 #() 
NAND2_X1_3880_ (
  .A1({ S22660 }),
  .A2({ S22632 }),
  .ZN({ S22661 })
);
INV_X1 #() 
INV_X1_1285_ (
  .A({ S22661 }),
  .ZN({ S22662 })
);
NAND4_X1 #() 
NAND4_X1_451_ (
  .A1({ S22630 }),
  .A2({ S22631 }),
  .A3({ S22640 }),
  .A4({ S22643 }),
  .ZN({ S22663 })
);
NAND2_X1 #() 
NAND2_X1_3881_ (
  .A1({ S77 }),
  .A2({ S22663 }),
  .ZN({ S22664 })
);
NAND3_X1 #() 
NAND3_X1_4142_ (
  .A1({ S22633 }),
  .A2({ S22630 }),
  .A3({ S22631 }),
  .ZN({ S22665 })
);
NAND2_X1 #() 
NAND2_X1_3882_ (
  .A1({ S22656 }),
  .A2({ S22665 }),
  .ZN({ S22666 })
);
NAND3_X1 #() 
NAND3_X1_4143_ (
  .A1({ S22666 }),
  .A2({ S25957[1035] }),
  .A3({ S22647 }),
  .ZN({ S22667 })
);
OAI21_X1 #() 
OAI21_X1_1976_ (
  .A({ S22667 }),
  .B1({ S22662 }),
  .B2({ S22664 }),
  .ZN({ S22668 })
);
OAI21_X1 #() 
OAI21_X1_1977_ (
  .A({ S25957[1037] }),
  .B1({ S22668 }),
  .B2({ S25957[1036] }),
  .ZN({ S22669 })
);
NOR2_X1 #() 
NOR2_X1_985_ (
  .A1({ S25957[1032] }),
  .A2({ S22634 }),
  .ZN({ S22670 })
);
AOI22_X1 #() 
AOI22_X1_436_ (
  .A1({ S21185 }),
  .A2({ S21186 }),
  .B1({ S25957[1034] }),
  .B2({ S22634 }),
  .ZN({ S22671 })
);
NAND2_X1 #() 
NAND2_X1_3883_ (
  .A1({ S22671 }),
  .A2({ S22632 }),
  .ZN({ S22672 })
);
OAI21_X1 #() 
OAI21_X1_1978_ (
  .A({ S22672 }),
  .B1({ S25957[1035] }),
  .B2({ S22670 }),
  .ZN({ S22673 })
);
OAI21_X1 #() 
OAI21_X1_1979_ (
  .A({ S21015 }),
  .B1({ S22673 }),
  .B2({ S22636 }),
  .ZN({ S22674 })
);
OAI22_X1 #() 
OAI22_X1_104_ (
  .A1({ S22674 }),
  .A2({ S22659 }),
  .B1({ S22669 }),
  .B2({ S22652 }),
  .ZN({ S22675 })
);
INV_X1 #() 
INV_X1_1286_ (
  .A({ S22648 }),
  .ZN({ S22676 })
);
NAND2_X1 #() 
NAND2_X1_3884_ (
  .A1({ S77 }),
  .A2({ S25957[1033] }),
  .ZN({ S22677 })
);
OAI21_X1 #() 
OAI21_X1_1980_ (
  .A({ S25957[1035] }),
  .B1({ S22634 }),
  .B2({ S22676 }),
  .ZN({ S22678 })
);
OAI21_X1 #() 
OAI21_X1_1981_ (
  .A({ S22678 }),
  .B1({ S22677 }),
  .B2({ S22676 }),
  .ZN({ S22679 })
);
NOR2_X1 #() 
NOR2_X1_986_ (
  .A1({ S22679 }),
  .A2({ S22636 }),
  .ZN({ S22680 })
);
NAND3_X1 #() 
NAND3_X1_4144_ (
  .A1({ S22660 }),
  .A2({ S21185 }),
  .A3({ S21186 }),
  .ZN({ S22681 })
);
NAND3_X1 #() 
NAND3_X1_4145_ (
  .A1({ S25957[1032] }),
  .A2({ S22634 }),
  .A3({ S22644 }),
  .ZN({ S22682 })
);
NAND4_X1 #() 
NAND4_X1_452_ (
  .A1({ S21386 }),
  .A2({ S21389 }),
  .A3({ S22628 }),
  .A4({ S22629 }),
  .ZN({ S22683 })
);
NAND2_X1 #() 
NAND2_X1_3885_ (
  .A1({ S22683 }),
  .A2({ S25957[1033] }),
  .ZN({ S22684 })
);
AOI21_X1 #() 
AOI21_X1_2093_ (
  .A({ S25957[1035] }),
  .B1({ S22682 }),
  .B2({ S22684 }),
  .ZN({ S22685 })
);
NAND2_X1 #() 
NAND2_X1_3886_ (
  .A1({ S22634 }),
  .A2({ S22644 }),
  .ZN({ S22686 })
);
INV_X1 #() 
INV_X1_1287_ (
  .A({ S22686 }),
  .ZN({ S22687 })
);
NAND2_X1 #() 
NAND2_X1_3887_ (
  .A1({ S25957[1035] }),
  .A2({ S22687 }),
  .ZN({ S22688 })
);
AOI211_X1 #() 
AOI211_X1_65_ (
  .A({ S25957[1036] }),
  .B({ S22685 }),
  .C1({ S22681 }),
  .C2({ S22688 }),
  .ZN({ S22689 })
);
NOR2_X1 #() 
NOR2_X1_987_ (
  .A1({ S22645 }),
  .A2({ S25957[1033] }),
  .ZN({ S22690 })
);
OAI21_X1 #() 
OAI21_X1_1982_ (
  .A({ S22632 }),
  .B1({ S22690 }),
  .B2({ S25957[1035] }),
  .ZN({ S22691 })
);
OAI21_X1 #() 
OAI21_X1_1983_ (
  .A({ S25957[1037] }),
  .B1({ S22691 }),
  .B2({ S25957[1036] }),
  .ZN({ S22692 })
);
NAND3_X1 #() 
NAND3_X1_4146_ (
  .A1({ S22656 }),
  .A2({ S22665 }),
  .A3({ S22644 }),
  .ZN({ S22693 })
);
NAND3_X1 #() 
NAND3_X1_4147_ (
  .A1({ S85 }),
  .A2({ S25957[1034] }),
  .A3({ S22632 }),
  .ZN({ S22694 })
);
AOI21_X1 #() 
AOI21_X1_2094_ (
  .A({ S77 }),
  .B1({ S22693 }),
  .B2({ S22694 }),
  .ZN({ S22695 })
);
INV_X1 #() 
INV_X1_1288_ (
  .A({ S22663 }),
  .ZN({ S22696 })
);
NAND3_X1 #() 
NAND3_X1_4148_ (
  .A1({ S21186 }),
  .A2({ S22683 }),
  .A3({ S21185 }),
  .ZN({ S22697 })
);
OAI21_X1 #() 
OAI21_X1_1984_ (
  .A({ S25957[1036] }),
  .B1({ S22697 }),
  .B2({ S22696 }),
  .ZN({ S22698 })
);
OAI21_X1 #() 
OAI21_X1_1985_ (
  .A({ S21015 }),
  .B1({ S22695 }),
  .B2({ S22698 }),
  .ZN({ S22699 })
);
OAI221_X1 #() 
OAI221_X1_115_ (
  .A({ S22635 }),
  .B1({ S22680 }),
  .B2({ S22692 }),
  .C1({ S22689 }),
  .C2({ S22699 }),
  .ZN({ S22700 })
);
OAI211_X1 #() 
OAI211_X1_1345_ (
  .A({ S22700 }),
  .B({ S25957[1039] }),
  .C1({ S22635 }),
  .C2({ S22675 }),
  .ZN({ S22701 })
);
NAND3_X1 #() 
NAND3_X1_4149_ (
  .A1({ S22656 }),
  .A2({ S22665 }),
  .A3({ S25957[1034] }),
  .ZN({ S22702 })
);
AOI21_X1 #() 
AOI21_X1_2095_ (
  .A({ S25957[1035] }),
  .B1({ S22702 }),
  .B2({ S22645 }),
  .ZN({ S22703 })
);
NAND2_X1 #() 
NAND2_X1_3888_ (
  .A1({ S22632 }),
  .A2({ S25957[1034] }),
  .ZN({ S22704 })
);
AOI21_X1 #() 
AOI21_X1_2096_ (
  .A({ S77 }),
  .B1({ S22693 }),
  .B2({ S22704 }),
  .ZN({ S22705 })
);
NOR3_X1 #() 
NOR3_X1_135_ (
  .A1({ S22705 }),
  .A2({ S22703 }),
  .A3({ S22636 }),
  .ZN({ S22706 })
);
NAND3_X1 #() 
NAND3_X1_4150_ (
  .A1({ S22661 }),
  .A2({ S25957[1035] }),
  .A3({ S22663 }),
  .ZN({ S22707 })
);
AOI21_X1 #() 
AOI21_X1_2097_ (
  .A({ S25957[1032] }),
  .B1({ S22634 }),
  .B2({ S25957[1034] }),
  .ZN({ S22708 })
);
NAND2_X1 #() 
NAND2_X1_3889_ (
  .A1({ S22708 }),
  .A2({ S77 }),
  .ZN({ S22709 })
);
AOI21_X1 #() 
AOI21_X1_2098_ (
  .A({ S22636 }),
  .B1({ S22707 }),
  .B2({ S22709 }),
  .ZN({ S22710 })
);
NAND2_X1 #() 
NAND2_X1_3890_ (
  .A1({ S22656 }),
  .A2({ S22644 }),
  .ZN({ S22711 })
);
NAND2_X1 #() 
NAND2_X1_3891_ (
  .A1({ S22671 }),
  .A2({ S22711 }),
  .ZN({ S22712 })
);
NAND3_X1 #() 
NAND3_X1_4151_ (
  .A1({ S22704 }),
  .A2({ S21185 }),
  .A3({ S21186 }),
  .ZN({ S22713 })
);
NAND3_X1 #() 
NAND3_X1_4152_ (
  .A1({ S22712 }),
  .A2({ S22636 }),
  .A3({ S22713 }),
  .ZN({ S22714 })
);
INV_X1 #() 
INV_X1_1289_ (
  .A({ S22714 }),
  .ZN({ S22715 })
);
OAI21_X1 #() 
OAI21_X1_1986_ (
  .A({ S25957[1037] }),
  .B1({ S22715 }),
  .B2({ S22710 }),
  .ZN({ S22716 })
);
INV_X1 #() 
INV_X1_1290_ (
  .A({ S22647 }),
  .ZN({ S22717 })
);
NAND3_X1 #() 
NAND3_X1_4153_ (
  .A1({ S21181 }),
  .A2({ S21184 }),
  .A3({ S22648 }),
  .ZN({ S22718 })
);
NOR2_X1 #() 
NOR2_X1_988_ (
  .A1({ S22718 }),
  .A2({ S22717 }),
  .ZN({ S22719 })
);
NAND2_X1 #() 
NAND2_X1_3892_ (
  .A1({ S22711 }),
  .A2({ S22704 }),
  .ZN({ S22720 })
);
AOI21_X1 #() 
AOI21_X1_2099_ (
  .A({ S25957[1036] }),
  .B1({ S22720 }),
  .B2({ S77 }),
  .ZN({ S22721 })
);
INV_X1 #() 
INV_X1_1291_ (
  .A({ S22721 }),
  .ZN({ S22722 })
);
OAI21_X1 #() 
OAI21_X1_1987_ (
  .A({ S21015 }),
  .B1({ S22722 }),
  .B2({ S22719 }),
  .ZN({ S22723 })
);
OAI211_X1 #() 
OAI211_X1_1346_ (
  .A({ S22716 }),
  .B({ S25957[1038] }),
  .C1({ S22706 }),
  .C2({ S22723 }),
  .ZN({ S22724 })
);
INV_X1 #() 
INV_X1_1292_ (
  .A({ S22724 }),
  .ZN({ S22725 })
);
NAND2_X1 #() 
NAND2_X1_3893_ (
  .A1({ S20874 }),
  .A2({ S20875 }),
  .ZN({ S22726 })
);
NAND2_X1 #() 
NAND2_X1_3894_ (
  .A1({ S77 }),
  .A2({ S25957[1032] }),
  .ZN({ S22727 })
);
INV_X1 #() 
INV_X1_1293_ (
  .A({ S22718 }),
  .ZN({ S22728 })
);
NAND2_X1 #() 
NAND2_X1_3895_ (
  .A1({ S22728 }),
  .A2({ S22686 }),
  .ZN({ S22729 })
);
AND2_X1 #() 
AND2_X1_242_ (
  .A1({ S22729 }),
  .A2({ S22727 }),
  .ZN({ S22730 })
);
NAND2_X1 #() 
NAND2_X1_3896_ (
  .A1({ S22686 }),
  .A2({ S22645 }),
  .ZN({ S22731 })
);
NAND2_X1 #() 
NAND2_X1_3897_ (
  .A1({ S85 }),
  .A2({ S22663 }),
  .ZN({ S22732 })
);
NAND2_X1 #() 
NAND2_X1_3898_ (
  .A1({ S22732 }),
  .A2({ S25957[1035] }),
  .ZN({ S22733 })
);
OAI211_X1 #() 
OAI211_X1_1347_ (
  .A({ S22733 }),
  .B({ S22636 }),
  .C1({ S22664 }),
  .C2({ S22731 }),
  .ZN({ S22734 })
);
OAI211_X1 #() 
OAI211_X1_1348_ (
  .A({ S25957[1037] }),
  .B({ S22734 }),
  .C1({ S22730 }),
  .C2({ S22636 }),
  .ZN({ S22735 })
);
OAI211_X1 #() 
OAI211_X1_1349_ (
  .A({ S21185 }),
  .B({ S21186 }),
  .C1({ S22632 }),
  .C2({ S25957[1034] }),
  .ZN({ S22736 })
);
INV_X1 #() 
INV_X1_1294_ (
  .A({ S22736 }),
  .ZN({ S22737 })
);
NAND2_X1 #() 
NAND2_X1_3899_ (
  .A1({ S22737 }),
  .A2({ S22694 }),
  .ZN({ S22738 })
);
NAND3_X1 #() 
NAND3_X1_4154_ (
  .A1({ S25957[1033] }),
  .A2({ S25957[1034] }),
  .A3({ S22633 }),
  .ZN({ S22739 })
);
AOI21_X1 #() 
AOI21_X1_2100_ (
  .A({ S22636 }),
  .B1({ S25957[1035] }),
  .B2({ S22739 }),
  .ZN({ S22740 })
);
INV_X1 #() 
INV_X1_1295_ (
  .A({ S22704 }),
  .ZN({ S22741 })
);
NAND2_X1 #() 
NAND2_X1_3900_ (
  .A1({ S22741 }),
  .A2({ S25957[1035] }),
  .ZN({ S22742 })
);
NOR2_X1 #() 
NOR2_X1_989_ (
  .A1({ S22702 }),
  .A2({ S25957[1035] }),
  .ZN({ S22743 })
);
NOR2_X1 #() 
NOR2_X1_990_ (
  .A1({ S22743 }),
  .A2({ S25957[1036] }),
  .ZN({ S22744 })
);
AOI22_X1 #() 
AOI22_X1_437_ (
  .A1({ S22744 }),
  .A2({ S22742 }),
  .B1({ S22740 }),
  .B2({ S22738 }),
  .ZN({ S22745 })
);
OAI21_X1 #() 
OAI21_X1_1988_ (
  .A({ S22735 }),
  .B1({ S22745 }),
  .B2({ S25957[1037] }),
  .ZN({ S22746 })
);
OAI21_X1 #() 
OAI21_X1_1989_ (
  .A({ S22726 }),
  .B1({ S22746 }),
  .B2({ S25957[1038] }),
  .ZN({ S22747 })
);
OR2_X1 #() 
OR2_X1_58_ (
  .A1({ S22747 }),
  .A2({ S22725 }),
  .ZN({ S22748 })
);
NAND2_X1 #() 
NAND2_X1_3901_ (
  .A1({ S22748 }),
  .A2({ S22701 }),
  .ZN({ S22749 })
);
NOR2_X1 #() 
NOR2_X1_991_ (
  .A1({ S22749 }),
  .A2({ S6989 }),
  .ZN({ S22750 })
);
NAND2_X1 #() 
NAND2_X1_3902_ (
  .A1({ S22749 }),
  .A2({ S6989 }),
  .ZN({ S22751 })
);
INV_X1 #() 
INV_X1_1296_ (
  .A({ S22751 }),
  .ZN({ S22752 })
);
OAI21_X1 #() 
OAI21_X1_1990_ (
  .A({ S25957[1079] }),
  .B1({ S22752 }),
  .B2({ S22750 }),
  .ZN({ S22753 })
);
OR3_X1 #() 
OR3_X1_25_ (
  .A1({ S22752 }),
  .A2({ S22750 }),
  .A3({ S25957[1079] }),
  .ZN({ S22754 })
);
NAND3_X1 #() 
NAND3_X1_4155_ (
  .A1({ S22754 }),
  .A2({ S20242 }),
  .A3({ S22753 }),
  .ZN({ S22755 })
);
NAND2_X1 #() 
NAND2_X1_3903_ (
  .A1({ S22754 }),
  .A2({ S22753 }),
  .ZN({ S25957[951] })
);
NAND2_X1 #() 
NAND2_X1_3904_ (
  .A1({ S25957[951] }),
  .A2({ S25957[1047] }),
  .ZN({ S22756 })
);
AND2_X1 #() 
AND2_X1_243_ (
  .A1({ S22756 }),
  .A2({ S22755 }),
  .ZN({ S25957[919] })
);
XOR2_X1 #() 
XOR2_X1_72_ (
  .A({ S25957[1110] }),
  .B({ S25957[1206] }),
  .Z({ S25957[1078] })
);
INV_X1 #() 
INV_X1_1297_ (
  .A({ S25957[1078] }),
  .ZN({ S22757 })
);
AOI21_X1 #() 
AOI21_X1_2101_ (
  .A({ S25957[1036] }),
  .B1({ S22672 }),
  .B2({ S22677 }),
  .ZN({ S22758 })
);
INV_X1 #() 
INV_X1_1298_ (
  .A({ S22683 }),
  .ZN({ S22759 })
);
NAND3_X1 #() 
NAND3_X1_4156_ (
  .A1({ S21181 }),
  .A2({ S21184 }),
  .A3({ S22634 }),
  .ZN({ S22760 })
);
NOR2_X1 #() 
NOR2_X1_992_ (
  .A1({ S22760 }),
  .A2({ S22759 }),
  .ZN({ S22761 })
);
NAND2_X1 #() 
NAND2_X1_3905_ (
  .A1({ S85 }),
  .A2({ S25957[1034] }),
  .ZN({ S22762 })
);
OAI21_X1 #() 
OAI21_X1_1991_ (
  .A({ S25957[1036] }),
  .B1({ S22762 }),
  .B2({ S25957[1035] }),
  .ZN({ S22763 })
);
AOI21_X1 #() 
AOI21_X1_2102_ (
  .A({ S22763 }),
  .B1({ S22761 }),
  .B2({ S22660 }),
  .ZN({ S22764 })
);
OAI21_X1 #() 
OAI21_X1_1992_ (
  .A({ S25957[1037] }),
  .B1({ S22764 }),
  .B2({ S22758 }),
  .ZN({ S22765 })
);
NAND2_X1 #() 
NAND2_X1_3906_ (
  .A1({ S22720 }),
  .A2({ S77 }),
  .ZN({ S22766 })
);
NAND2_X1 #() 
NAND2_X1_3907_ (
  .A1({ S22632 }),
  .A2({ S22644 }),
  .ZN({ S22767 })
);
NOR2_X1 #() 
NOR2_X1_993_ (
  .A1({ S77 }),
  .A2({ S22767 }),
  .ZN({ S22768 })
);
NAND2_X1 #() 
NAND2_X1_3908_ (
  .A1({ S25957[1035] }),
  .A2({ S22653 }),
  .ZN({ S22769 })
);
AOI21_X1 #() 
AOI21_X1_2103_ (
  .A({ S22768 }),
  .B1({ S22766 }),
  .B2({ S22769 }),
  .ZN({ S22770 })
);
INV_X1 #() 
INV_X1_1299_ (
  .A({ S22681 }),
  .ZN({ S22771 })
);
NAND2_X1 #() 
NAND2_X1_3909_ (
  .A1({ S22771 }),
  .A2({ S22693 }),
  .ZN({ S22772 })
);
NAND3_X1 #() 
NAND3_X1_4157_ (
  .A1({ S22660 }),
  .A2({ S22632 }),
  .A3({ S22683 }),
  .ZN({ S22773 })
);
AOI21_X1 #() 
AOI21_X1_2104_ (
  .A({ S22636 }),
  .B1({ S22773 }),
  .B2({ S25957[1035] }),
  .ZN({ S22774 })
);
AOI21_X1 #() 
AOI21_X1_2105_ (
  .A({ S25957[1037] }),
  .B1({ S22772 }),
  .B2({ S22774 }),
  .ZN({ S22775 })
);
OAI21_X1 #() 
OAI21_X1_1993_ (
  .A({ S22775 }),
  .B1({ S22770 }),
  .B2({ S25957[1036] }),
  .ZN({ S22776 })
);
NAND3_X1 #() 
NAND3_X1_4158_ (
  .A1({ S22776 }),
  .A2({ S25957[1038] }),
  .A3({ S22765 }),
  .ZN({ S22777 })
);
NAND2_X1 #() 
NAND2_X1_3910_ (
  .A1({ S77 }),
  .A2({ S22647 }),
  .ZN({ S22778 })
);
OAI211_X1 #() 
OAI211_X1_1350_ (
  .A({ S22640 }),
  .B({ S22643 }),
  .C1({ S21316 }),
  .C2({ S21313 }),
  .ZN({ S22779 })
);
OAI21_X1 #() 
OAI21_X1_1994_ (
  .A({ S22779 }),
  .B1({ S22647 }),
  .B2({ S25957[1032] }),
  .ZN({ S22780 })
);
OAI22_X1 #() 
OAI22_X1_105_ (
  .A1({ S22778 }),
  .A2({ S22666 }),
  .B1({ S22780 }),
  .B2({ S77 }),
  .ZN({ S22781 })
);
NAND2_X1 #() 
NAND2_X1_3911_ (
  .A1({ S25957[1035] }),
  .A2({ S22696 }),
  .ZN({ S22782 })
);
NAND3_X1 #() 
NAND3_X1_4159_ (
  .A1({ S25957[1033] }),
  .A2({ S22633 }),
  .A3({ S22644 }),
  .ZN({ S22783 })
);
OAI21_X1 #() 
OAI21_X1_1995_ (
  .A({ S22782 }),
  .B1({ S25957[1035] }),
  .B2({ S22783 }),
  .ZN({ S22784 })
);
OAI21_X1 #() 
OAI21_X1_1996_ (
  .A({ S25957[1036] }),
  .B1({ S22784 }),
  .B2({ S22743 }),
  .ZN({ S22785 })
);
OAI21_X1 #() 
OAI21_X1_1997_ (
  .A({ S22785 }),
  .B1({ S25957[1036] }),
  .B2({ S22781 }),
  .ZN({ S22786 })
);
NAND2_X1 #() 
NAND2_X1_3912_ (
  .A1({ S22786 }),
  .A2({ S25957[1037] }),
  .ZN({ S22787 })
);
NAND2_X1 #() 
NAND2_X1_3913_ (
  .A1({ S22645 }),
  .A2({ S22647 }),
  .ZN({ S22788 })
);
OAI21_X1 #() 
OAI21_X1_1998_ (
  .A({ S22760 }),
  .B1({ S77 }),
  .B2({ S22648 }),
  .ZN({ S22789 })
);
AOI21_X1 #() 
AOI21_X1_2106_ (
  .A({ S22789 }),
  .B1({ S22788 }),
  .B2({ S77 }),
  .ZN({ S22790 })
);
OAI21_X1 #() 
OAI21_X1_1999_ (
  .A({ S22683 }),
  .B1({ S22663 }),
  .B2({ S25957[1032] }),
  .ZN({ S22791 })
);
NAND2_X1 #() 
NAND2_X1_3914_ (
  .A1({ S22791 }),
  .A2({ S25957[1035] }),
  .ZN({ S22792 })
);
NAND3_X1 #() 
NAND3_X1_4160_ (
  .A1({ S22772 }),
  .A2({ S22636 }),
  .A3({ S22792 }),
  .ZN({ S22793 })
);
OAI211_X1 #() 
OAI211_X1_1351_ (
  .A({ S22793 }),
  .B({ S21015 }),
  .C1({ S22790 }),
  .C2({ S22636 }),
  .ZN({ S22794 })
);
NAND3_X1 #() 
NAND3_X1_4161_ (
  .A1({ S22787 }),
  .A2({ S22794 }),
  .A3({ S22635 }),
  .ZN({ S22795 })
);
NAND3_X1 #() 
NAND3_X1_4162_ (
  .A1({ S22795 }),
  .A2({ S25957[1039] }),
  .A3({ S22777 }),
  .ZN({ S22796 })
);
NAND2_X1 #() 
NAND2_X1_3915_ (
  .A1({ S22686 }),
  .A2({ S22633 }),
  .ZN({ S22797 })
);
NAND4_X1 #() 
NAND4_X1_453_ (
  .A1({ S21181 }),
  .A2({ S21184 }),
  .A3({ S25957[1033] }),
  .A4({ S22644 }),
  .ZN({ S22798 })
);
OAI21_X1 #() 
OAI21_X1_2000_ (
  .A({ S22798 }),
  .B1({ S25957[1035] }),
  .B2({ S22797 }),
  .ZN({ S22799 })
);
NAND2_X1 #() 
NAND2_X1_3916_ (
  .A1({ S22694 }),
  .A2({ S77 }),
  .ZN({ S22800 })
);
NAND2_X1 #() 
NAND2_X1_3917_ (
  .A1({ S22773 }),
  .A2({ S25957[1035] }),
  .ZN({ S22801 })
);
AOI21_X1 #() 
AOI21_X1_2107_ (
  .A({ S25957[1036] }),
  .B1({ S22801 }),
  .B2({ S22800 }),
  .ZN({ S22802 })
);
AOI211_X1 #() 
AOI211_X1_66_ (
  .A({ S25957[1037] }),
  .B({ S22802 }),
  .C1({ S25957[1036] }),
  .C2({ S22799 }),
  .ZN({ S22803 })
);
OAI21_X1 #() 
OAI21_X1_2001_ (
  .A({ S22645 }),
  .B1({ S22634 }),
  .B2({ S22648 }),
  .ZN({ S22804 })
);
NAND2_X1 #() 
NAND2_X1_3918_ (
  .A1({ S22804 }),
  .A2({ S77 }),
  .ZN({ S22805 })
);
NAND2_X1 #() 
NAND2_X1_3919_ (
  .A1({ S85 }),
  .A2({ S22683 }),
  .ZN({ S22806 })
);
OAI211_X1 #() 
OAI211_X1_1352_ (
  .A({ S22805 }),
  .B({ S25957[1036] }),
  .C1({ S77 }),
  .C2({ S22806 }),
  .ZN({ S22807 })
);
NAND2_X1 #() 
NAND2_X1_3920_ (
  .A1({ S25957[1035] }),
  .A2({ S22676 }),
  .ZN({ S22808 })
);
INV_X1 #() 
INV_X1_1300_ (
  .A({ S22808 }),
  .ZN({ S22809 })
);
NAND2_X1 #() 
NAND2_X1_3921_ (
  .A1({ S22665 }),
  .A2({ S22663 }),
  .ZN({ S22810 })
);
OAI21_X1 #() 
OAI21_X1_2002_ (
  .A({ S22636 }),
  .B1({ S22809 }),
  .B2({ S22810 }),
  .ZN({ S22811 })
);
AND3_X1 #() 
AND3_X1_148_ (
  .A1({ S22811 }),
  .A2({ S22807 }),
  .A3({ S25957[1037] }),
  .ZN({ S22812 })
);
OAI21_X1 #() 
OAI21_X1_2003_ (
  .A({ S25957[1038] }),
  .B1({ S22803 }),
  .B2({ S22812 }),
  .ZN({ S22813 })
);
AOI21_X1 #() 
AOI21_X1_2108_ (
  .A({ S25957[1036] }),
  .B1({ S25957[1035] }),
  .B2({ S22687 }),
  .ZN({ S22814 })
);
NAND2_X1 #() 
NAND2_X1_3922_ (
  .A1({ S22814 }),
  .A2({ S22792 }),
  .ZN({ S22815 })
);
AOI22_X1 #() 
AOI22_X1_438_ (
  .A1({ S22671 }),
  .A2({ S22711 }),
  .B1({ S77 }),
  .B2({ S22682 }),
  .ZN({ S22816 })
);
OAI21_X1 #() 
OAI21_X1_2004_ (
  .A({ S22815 }),
  .B1({ S22816 }),
  .B2({ S22636 }),
  .ZN({ S22817 })
);
NAND3_X1 #() 
NAND3_X1_4163_ (
  .A1({ S22779 }),
  .A2({ S21181 }),
  .A3({ S21184 }),
  .ZN({ S22818 })
);
NAND3_X1 #() 
NAND3_X1_4164_ (
  .A1({ S22779 }),
  .A2({ S22645 }),
  .A3({ S22647 }),
  .ZN({ S22819 })
);
NAND2_X1 #() 
NAND2_X1_3923_ (
  .A1({ S22819 }),
  .A2({ S77 }),
  .ZN({ S22820 })
);
OAI21_X1 #() 
OAI21_X1_2005_ (
  .A({ S22820 }),
  .B1({ S22717 }),
  .B2({ S22818 }),
  .ZN({ S22821 })
);
OAI211_X1 #() 
OAI211_X1_1353_ (
  .A({ S25957[1036] }),
  .B({ S22697 }),
  .C1({ S22769 }),
  .C2({ S84 }),
  .ZN({ S22822 })
);
OAI211_X1 #() 
OAI211_X1_1354_ (
  .A({ S25957[1037] }),
  .B({ S22822 }),
  .C1({ S22821 }),
  .C2({ S25957[1036] }),
  .ZN({ S22823 })
);
OAI211_X1 #() 
OAI211_X1_1355_ (
  .A({ S22823 }),
  .B({ S22635 }),
  .C1({ S25957[1037] }),
  .C2({ S22817 }),
  .ZN({ S22824 })
);
NAND3_X1 #() 
NAND3_X1_4165_ (
  .A1({ S22813 }),
  .A2({ S22726 }),
  .A3({ S22824 }),
  .ZN({ S22825 })
);
NAND3_X1 #() 
NAND3_X1_4166_ (
  .A1({ S22825 }),
  .A2({ S22796 }),
  .A3({ S25957[1238] }),
  .ZN({ S22826 })
);
INV_X1 #() 
INV_X1_1301_ (
  .A({ S22826 }),
  .ZN({ S22827 })
);
AOI21_X1 #() 
AOI21_X1_2109_ (
  .A({ S25957[1238] }),
  .B1({ S22825 }),
  .B2({ S22796 }),
  .ZN({ S22828 })
);
OAI21_X1 #() 
OAI21_X1_2006_ (
  .A({ S22757 }),
  .B1({ S22827 }),
  .B2({ S22828 }),
  .ZN({ S22829 })
);
NOR2_X1 #() 
NOR2_X1_994_ (
  .A1({ S22827 }),
  .A2({ S22828 }),
  .ZN({ S25957[982] })
);
NAND2_X1 #() 
NAND2_X1_3924_ (
  .A1({ S25957[982] }),
  .A2({ S25957[1078] }),
  .ZN({ S22830 })
);
NAND3_X1 #() 
NAND3_X1_4167_ (
  .A1({ S22830 }),
  .A2({ S25957[1046] }),
  .A3({ S22829 }),
  .ZN({ S22831 })
);
AND2_X1 #() 
AND2_X1_244_ (
  .A1({ S20317 }),
  .A2({ S20316 }),
  .ZN({ S22832 })
);
OAI21_X1 #() 
OAI21_X1_2007_ (
  .A({ S25957[1078] }),
  .B1({ S22827 }),
  .B2({ S22828 }),
  .ZN({ S22833 })
);
NAND2_X1 #() 
NAND2_X1_3925_ (
  .A1({ S25957[982] }),
  .A2({ S22757 }),
  .ZN({ S22834 })
);
NAND3_X1 #() 
NAND3_X1_4168_ (
  .A1({ S22834 }),
  .A2({ S22832 }),
  .A3({ S22833 }),
  .ZN({ S22835 })
);
NAND2_X1 #() 
NAND2_X1_3926_ (
  .A1({ S22831 }),
  .A2({ S22835 }),
  .ZN({ S22836 })
);
INV_X1 #() 
INV_X1_1302_ (
  .A({ S22836 }),
  .ZN({ S25957[918] })
);
NAND2_X1 #() 
NAND2_X1_3927_ (
  .A1({ S20385 }),
  .A2({ S20389 }),
  .ZN({ S22837 })
);
XNOR2_X1 #() 
XNOR2_X1_169_ (
  .A({ S22837 }),
  .B({ S25957[1205] }),
  .ZN({ S25957[1077] })
);
INV_X1 #() 
INV_X1_1303_ (
  .A({ S25957[1077] }),
  .ZN({ S22838 })
);
AOI22_X1 #() 
AOI22_X1_439_ (
  .A1({ S22630 }),
  .A2({ S22631 }),
  .B1({ S22629 }),
  .B2({ S22628 }),
  .ZN({ S22839 })
);
NAND2_X1 #() 
NAND2_X1_3928_ (
  .A1({ S22839 }),
  .A2({ S22644 }),
  .ZN({ S22840 })
);
AOI21_X1 #() 
AOI21_X1_2110_ (
  .A({ S77 }),
  .B1({ S22694 }),
  .B2({ S22840 }),
  .ZN({ S22841 })
);
NAND2_X1 #() 
NAND2_X1_3929_ (
  .A1({ S22736 }),
  .A2({ S21015 }),
  .ZN({ S22842 })
);
NOR2_X1 #() 
NOR2_X1_995_ (
  .A1({ S25957[1035] }),
  .A2({ S22670 }),
  .ZN({ S22843 })
);
NAND2_X1 #() 
NAND2_X1_3930_ (
  .A1({ S22843 }),
  .A2({ S22686 }),
  .ZN({ S22844 })
);
NAND3_X1 #() 
NAND3_X1_4169_ (
  .A1({ S22844 }),
  .A2({ S25957[1037] }),
  .A3({ S22760 }),
  .ZN({ S22845 })
);
OAI21_X1 #() 
OAI21_X1_2008_ (
  .A({ S22845 }),
  .B1({ S22841 }),
  .B2({ S22842 }),
  .ZN({ S22846 })
);
NAND2_X1 #() 
NAND2_X1_3931_ (
  .A1({ S22846 }),
  .A2({ S22636 }),
  .ZN({ S22847 })
);
AOI22_X1 #() 
AOI22_X1_440_ (
  .A1({ S21386 }),
  .A2({ S21389 }),
  .B1({ S22629 }),
  .B2({ S22628 }),
  .ZN({ S22848 })
);
OAI21_X1 #() 
OAI21_X1_2009_ (
  .A({ S77 }),
  .B1({ S22657 }),
  .B2({ S22848 }),
  .ZN({ S22849 })
);
OAI211_X1 #() 
OAI211_X1_1356_ (
  .A({ S22849 }),
  .B({ S25957[1037] }),
  .C1({ S22720 }),
  .C2({ S77 }),
  .ZN({ S22850 })
);
NAND2_X1 #() 
NAND2_X1_3932_ (
  .A1({ S22731 }),
  .A2({ S85 }),
  .ZN({ S22851 })
);
NOR2_X1 #() 
NOR2_X1_996_ (
  .A1({ S22851 }),
  .A2({ S77 }),
  .ZN({ S22852 })
);
NOR2_X1 #() 
NOR2_X1_997_ (
  .A1({ S22697 }),
  .A2({ S25957[1033] }),
  .ZN({ S22853 })
);
OAI21_X1 #() 
OAI21_X1_2010_ (
  .A({ S21015 }),
  .B1({ S22852 }),
  .B2({ S22853 }),
  .ZN({ S22854 })
);
NAND2_X1 #() 
NAND2_X1_3933_ (
  .A1({ S22854 }),
  .A2({ S22850 }),
  .ZN({ S22855 })
);
NAND2_X1 #() 
NAND2_X1_3934_ (
  .A1({ S22855 }),
  .A2({ S25957[1036] }),
  .ZN({ S22856 })
);
AND2_X1 #() 
AND2_X1_245_ (
  .A1({ S22856 }),
  .A2({ S22847 }),
  .ZN({ S22857 })
);
AOI21_X1 #() 
AOI21_X1_2111_ (
  .A({ S25957[1032] }),
  .B1({ S21186 }),
  .B2({ S21185 }),
  .ZN({ S22858 })
);
AOI22_X1 #() 
AOI22_X1_441_ (
  .A1({ S22843 }),
  .A2({ S22711 }),
  .B1({ S22686 }),
  .B2({ S22858 }),
  .ZN({ S22859 })
);
NAND2_X1 #() 
NAND2_X1_3935_ (
  .A1({ S22859 }),
  .A2({ S25957[1036] }),
  .ZN({ S22860 })
);
NAND4_X1 #() 
NAND4_X1_454_ (
  .A1({ S21181 }),
  .A2({ S21184 }),
  .A3({ S22663 }),
  .A4({ S22632 }),
  .ZN({ S22861 })
);
NAND3_X1 #() 
NAND3_X1_4170_ (
  .A1({ S22677 }),
  .A2({ S22648 }),
  .A3({ S22861 }),
  .ZN({ S22862 })
);
NAND2_X1 #() 
NAND2_X1_3936_ (
  .A1({ S22862 }),
  .A2({ S22636 }),
  .ZN({ S22863 })
);
AOI21_X1 #() 
AOI21_X1_2112_ (
  .A({ S21015 }),
  .B1({ S22860 }),
  .B2({ S22863 }),
  .ZN({ S22864 })
);
INV_X1 #() 
INV_X1_1304_ (
  .A({ S22864 }),
  .ZN({ S22865 })
);
NAND2_X1 #() 
NAND2_X1_3937_ (
  .A1({ S22744 }),
  .A2({ S22801 }),
  .ZN({ S22866 })
);
NAND4_X1 #() 
NAND4_X1_455_ (
  .A1({ S22686 }),
  .A2({ S22683 }),
  .A3({ S21181 }),
  .A4({ S21184 }),
  .ZN({ S22867 })
);
NAND2_X1 #() 
NAND2_X1_3938_ (
  .A1({ S22779 }),
  .A2({ S22648 }),
  .ZN({ S22868 })
);
NAND2_X1 #() 
NAND2_X1_3939_ (
  .A1({ S22868 }),
  .A2({ S77 }),
  .ZN({ S22869 })
);
NAND2_X1 #() 
NAND2_X1_3940_ (
  .A1({ S22869 }),
  .A2({ S22867 }),
  .ZN({ S22870 })
);
OAI21_X1 #() 
OAI21_X1_2011_ (
  .A({ S21015 }),
  .B1({ S22870 }),
  .B2({ S22636 }),
  .ZN({ S22871 })
);
INV_X1 #() 
INV_X1_1305_ (
  .A({ S22871 }),
  .ZN({ S22872 })
);
AOI21_X1 #() 
AOI21_X1_2113_ (
  .A({ S22635 }),
  .B1({ S22872 }),
  .B2({ S22866 }),
  .ZN({ S22873 })
);
AOI21_X1 #() 
AOI21_X1_2114_ (
  .A({ S22726 }),
  .B1({ S22865 }),
  .B2({ S22873 }),
  .ZN({ S22874 })
);
OAI21_X1 #() 
OAI21_X1_2012_ (
  .A({ S22874 }),
  .B1({ S22857 }),
  .B2({ S25957[1038] }),
  .ZN({ S22875 })
);
AOI21_X1 #() 
AOI21_X1_2115_ (
  .A({ S22644 }),
  .B1({ S85 }),
  .B2({ S22632 }),
  .ZN({ S22876 })
);
NOR2_X1 #() 
NOR2_X1_998_ (
  .A1({ S22647 }),
  .A2({ S25957[1032] }),
  .ZN({ S22877 })
);
OAI21_X1 #() 
OAI21_X1_2013_ (
  .A({ S25957[1035] }),
  .B1({ S22876 }),
  .B2({ S22877 }),
  .ZN({ S22878 })
);
NAND3_X1 #() 
NAND3_X1_4171_ (
  .A1({ S22878 }),
  .A2({ S25957[1036] }),
  .A3({ S22820 }),
  .ZN({ S22879 })
);
NAND2_X1 #() 
NAND2_X1_3941_ (
  .A1({ S25957[1035] }),
  .A2({ S22633 }),
  .ZN({ S22880 })
);
NAND4_X1 #() 
NAND4_X1_456_ (
  .A1({ S22665 }),
  .A2({ S22683 }),
  .A3({ S21185 }),
  .A4({ S21186 }),
  .ZN({ S22881 })
);
NAND3_X1 #() 
NAND3_X1_4172_ (
  .A1({ S22880 }),
  .A2({ S22636 }),
  .A3({ S22881 }),
  .ZN({ S22882 })
);
NAND3_X1 #() 
NAND3_X1_4173_ (
  .A1({ S22879 }),
  .A2({ S25957[1037] }),
  .A3({ S22882 }),
  .ZN({ S22883 })
);
NAND2_X1 #() 
NAND2_X1_3942_ (
  .A1({ S22804 }),
  .A2({ S25957[1035] }),
  .ZN({ S22884 })
);
NOR2_X1 #() 
NOR2_X1_999_ (
  .A1({ S22877 }),
  .A2({ S25957[1035] }),
  .ZN({ S22885 })
);
NAND2_X1 #() 
NAND2_X1_3943_ (
  .A1({ S22885 }),
  .A2({ S22648 }),
  .ZN({ S22886 })
);
AOI21_X1 #() 
AOI21_X1_2116_ (
  .A({ S25957[1036] }),
  .B1({ S22886 }),
  .B2({ S22884 }),
  .ZN({ S22887 })
);
NAND2_X1 #() 
NAND2_X1_3944_ (
  .A1({ S22788 }),
  .A2({ S25957[1035] }),
  .ZN({ S22888 })
);
NAND3_X1 #() 
NAND3_X1_4174_ (
  .A1({ S25957[1033] }),
  .A2({ S25957[1032] }),
  .A3({ S25957[1034] }),
  .ZN({ S22889 })
);
NAND3_X1 #() 
NAND3_X1_4175_ (
  .A1({ S77 }),
  .A2({ S22889 }),
  .A3({ S22767 }),
  .ZN({ S22890 })
);
AND3_X1 #() 
AND3_X1_149_ (
  .A1({ S22890 }),
  .A2({ S22888 }),
  .A3({ S25957[1036] }),
  .ZN({ S22891 })
);
OAI21_X1 #() 
OAI21_X1_2014_ (
  .A({ S21015 }),
  .B1({ S22887 }),
  .B2({ S22891 }),
  .ZN({ S22892 })
);
NAND2_X1 #() 
NAND2_X1_3945_ (
  .A1({ S22892 }),
  .A2({ S22883 }),
  .ZN({ S22893 })
);
INV_X1 #() 
INV_X1_1306_ (
  .A({ S22760 }),
  .ZN({ S22894 })
);
NOR2_X1 #() 
NOR2_X1_1000_ (
  .A1({ S22648 }),
  .A2({ S22634 }),
  .ZN({ S22895 })
);
AOI22_X1 #() 
AOI22_X1_442_ (
  .A1({ S22894 }),
  .A2({ S25957[1032] }),
  .B1({ S77 }),
  .B2({ S22895 }),
  .ZN({ S22896 })
);
NAND3_X1 #() 
NAND3_X1_4176_ (
  .A1({ S22702 }),
  .A2({ S25957[1035] }),
  .A3({ S22682 }),
  .ZN({ S22897 })
);
NAND2_X1 #() 
NAND2_X1_3946_ (
  .A1({ S85 }),
  .A2({ S22632 }),
  .ZN({ S22898 })
);
AOI22_X1 #() 
AOI22_X1_443_ (
  .A1({ S21184 }),
  .A2({ S21181 }),
  .B1({ S22633 }),
  .B2({ S22644 }),
  .ZN({ S22899 })
);
NAND2_X1 #() 
NAND2_X1_3947_ (
  .A1({ S22899 }),
  .A2({ S22898 }),
  .ZN({ S22900 })
);
NAND3_X1 #() 
NAND3_X1_4177_ (
  .A1({ S22897 }),
  .A2({ S22900 }),
  .A3({ S25957[1036] }),
  .ZN({ S22901 })
);
OAI21_X1 #() 
OAI21_X1_2015_ (
  .A({ S22901 }),
  .B1({ S25957[1036] }),
  .B2({ S22896 }),
  .ZN({ S22902 })
);
AOI21_X1 #() 
AOI21_X1_2117_ (
  .A({ S25957[1036] }),
  .B1({ S22808 }),
  .B2({ S22684 }),
  .ZN({ S22903 })
);
OAI21_X1 #() 
OAI21_X1_2016_ (
  .A({ S22903 }),
  .B1({ S22771 }),
  .B2({ S22809 }),
  .ZN({ S22904 })
);
OAI21_X1 #() 
OAI21_X1_2017_ (
  .A({ S25957[1036] }),
  .B1({ S22885 }),
  .B2({ S22768 }),
  .ZN({ S22905 })
);
NAND3_X1 #() 
NAND3_X1_4178_ (
  .A1({ S22904 }),
  .A2({ S25957[1037] }),
  .A3({ S22905 }),
  .ZN({ S22906 })
);
OAI21_X1 #() 
OAI21_X1_2018_ (
  .A({ S22906 }),
  .B1({ S25957[1037] }),
  .B2({ S22902 }),
  .ZN({ S22907 })
);
NAND2_X1 #() 
NAND2_X1_3948_ (
  .A1({ S22907 }),
  .A2({ S22635 }),
  .ZN({ S22908 })
);
OAI211_X1 #() 
OAI211_X1_1357_ (
  .A({ S22908 }),
  .B({ S22726 }),
  .C1({ S22635 }),
  .C2({ S22893 }),
  .ZN({ S22909 })
);
NAND3_X1 #() 
NAND3_X1_4179_ (
  .A1({ S22909 }),
  .A2({ S22875 }),
  .A3({ S20386 }),
  .ZN({ S22910 })
);
AOI21_X1 #() 
AOI21_X1_2118_ (
  .A({ S22864 }),
  .B1({ S22866 }),
  .B2({ S22872 }),
  .ZN({ S22911 })
);
NAND3_X1 #() 
NAND3_X1_4180_ (
  .A1({ S22856 }),
  .A2({ S22847 }),
  .A3({ S22635 }),
  .ZN({ S22912 })
);
OAI211_X1 #() 
OAI211_X1_1358_ (
  .A({ S22912 }),
  .B({ S25957[1039] }),
  .C1({ S22911 }),
  .C2({ S22635 }),
  .ZN({ S22913 })
);
NAND2_X1 #() 
NAND2_X1_3949_ (
  .A1({ S22893 }),
  .A2({ S25957[1038] }),
  .ZN({ S22914 })
);
OAI211_X1 #() 
OAI211_X1_1359_ (
  .A({ S22906 }),
  .B({ S22635 }),
  .C1({ S25957[1037] }),
  .C2({ S22902 }),
  .ZN({ S22915 })
);
NAND3_X1 #() 
NAND3_X1_4181_ (
  .A1({ S22914 }),
  .A2({ S22726 }),
  .A3({ S22915 }),
  .ZN({ S22916 })
);
NAND3_X1 #() 
NAND3_X1_4182_ (
  .A1({ S22913 }),
  .A2({ S22916 }),
  .A3({ S25957[1237] }),
  .ZN({ S22917 })
);
NAND3_X1 #() 
NAND3_X1_4183_ (
  .A1({ S22910 }),
  .A2({ S22917 }),
  .A3({ S22838 }),
  .ZN({ S22918 })
);
NAND2_X1 #() 
NAND2_X1_3950_ (
  .A1({ S22910 }),
  .A2({ S22917 }),
  .ZN({ S25957[981] })
);
NAND2_X1 #() 
NAND2_X1_3951_ (
  .A1({ S25957[981] }),
  .A2({ S25957[1077] }),
  .ZN({ S22919 })
);
NAND3_X1 #() 
NAND3_X1_4184_ (
  .A1({ S22919 }),
  .A2({ S25957[1045] }),
  .A3({ S22918 }),
  .ZN({ S22920 })
);
INV_X1 #() 
INV_X1_1307_ (
  .A({ S25957[1045] }),
  .ZN({ S22921 })
);
NAND2_X1 #() 
NAND2_X1_3952_ (
  .A1({ S25957[981] }),
  .A2({ S22838 }),
  .ZN({ S22922 })
);
NAND3_X1 #() 
NAND3_X1_4185_ (
  .A1({ S22910 }),
  .A2({ S22917 }),
  .A3({ S25957[1077] }),
  .ZN({ S22923 })
);
NAND3_X1 #() 
NAND3_X1_4186_ (
  .A1({ S22922 }),
  .A2({ S22921 }),
  .A3({ S22923 }),
  .ZN({ S22924 })
);
AND2_X1 #() 
AND2_X1_246_ (
  .A1({ S22924 }),
  .A2({ S22920 }),
  .ZN({ S25957[917] })
);
NOR2_X1 #() 
NOR2_X1_1001_ (
  .A1({ S20466 }),
  .A2({ S20465 }),
  .ZN({ S25957[1076] })
);
AOI21_X1 #() 
AOI21_X1_2119_ (
  .A({ S25957[1035] }),
  .B1({ S22693 }),
  .B2({ S22704 }),
  .ZN({ S22925 })
);
NAND2_X1 #() 
NAND2_X1_3953_ (
  .A1({ S25957[1035] }),
  .A2({ S22670 }),
  .ZN({ S22926 })
);
NAND3_X1 #() 
NAND3_X1_4187_ (
  .A1({ S22888 }),
  .A2({ S22926 }),
  .A3({ S22636 }),
  .ZN({ S22927 })
);
OAI211_X1 #() 
OAI211_X1_1360_ (
  .A({ S21181 }),
  .B({ S21184 }),
  .C1({ S22647 }),
  .C2({ S25957[1032] }),
  .ZN({ S22928 })
);
NAND2_X1 #() 
NAND2_X1_3954_ (
  .A1({ S22663 }),
  .A2({ S22632 }),
  .ZN({ S22929 })
);
NAND2_X1 #() 
NAND2_X1_3955_ (
  .A1({ S22686 }),
  .A2({ S85 }),
  .ZN({ S22930 })
);
OAI21_X1 #() 
OAI21_X1_2019_ (
  .A({ S77 }),
  .B1({ S22930 }),
  .B2({ S22929 }),
  .ZN({ S22931 })
);
OAI211_X1 #() 
OAI211_X1_1361_ (
  .A({ S22931 }),
  .B({ S25957[1036] }),
  .C1({ S22657 }),
  .C2({ S22928 }),
  .ZN({ S22932 })
);
OAI211_X1 #() 
OAI211_X1_1362_ (
  .A({ S22932 }),
  .B({ S25957[1037] }),
  .C1({ S22925 }),
  .C2({ S22927 }),
  .ZN({ S22933 })
);
NOR2_X1 #() 
NOR2_X1_1002_ (
  .A1({ S22663 }),
  .A2({ S25957[1032] }),
  .ZN({ S22934 })
);
OAI21_X1 #() 
OAI21_X1_2020_ (
  .A({ S25957[1035] }),
  .B1({ S22934 }),
  .B2({ S22687 }),
  .ZN({ S22935 })
);
OAI21_X1 #() 
OAI21_X1_2021_ (
  .A({ S22935 }),
  .B1({ S22934 }),
  .B2({ S22736 }),
  .ZN({ S22936 })
);
NAND2_X1 #() 
NAND2_X1_3956_ (
  .A1({ S22648 }),
  .A2({ S22634 }),
  .ZN({ S22937 })
);
NOR2_X1 #() 
NOR2_X1_1003_ (
  .A1({ S77 }),
  .A2({ S22937 }),
  .ZN({ S22938 })
);
NAND3_X1 #() 
NAND3_X1_4188_ (
  .A1({ S85 }),
  .A2({ S22645 }),
  .A3({ S22648 }),
  .ZN({ S22939 })
);
NAND4_X1 #() 
NAND4_X1_457_ (
  .A1({ S21185 }),
  .A2({ S21186 }),
  .A3({ S22634 }),
  .A4({ S22644 }),
  .ZN({ S22940 })
);
OAI211_X1 #() 
OAI211_X1_1363_ (
  .A({ S22940 }),
  .B({ S22636 }),
  .C1({ S22939 }),
  .C2({ S25957[1035] }),
  .ZN({ S22941 })
);
OAI221_X1 #() 
OAI221_X1_116_ (
  .A({ S21015 }),
  .B1({ S22941 }),
  .B2({ S22938 }),
  .C1({ S22936 }),
  .C2({ S22636 }),
  .ZN({ S22942 })
);
NAND3_X1 #() 
NAND3_X1_4189_ (
  .A1({ S22942 }),
  .A2({ S22933 }),
  .A3({ S22635 }),
  .ZN({ S22943 })
);
NAND3_X1 #() 
NAND3_X1_4190_ (
  .A1({ S77 }),
  .A2({ S22633 }),
  .A3({ S22647 }),
  .ZN({ S22944 })
);
NAND3_X1 #() 
NAND3_X1_4191_ (
  .A1({ S22729 }),
  .A2({ S22636 }),
  .A3({ S22944 }),
  .ZN({ S22945 })
);
NAND2_X1 #() 
NAND2_X1_3957_ (
  .A1({ S77 }),
  .A2({ S22653 }),
  .ZN({ S22946 })
);
NAND3_X1 #() 
NAND3_X1_4192_ (
  .A1({ S22888 }),
  .A2({ S22946 }),
  .A3({ S25957[1036] }),
  .ZN({ S22947 })
);
NAND3_X1 #() 
NAND3_X1_4193_ (
  .A1({ S22945 }),
  .A2({ S25957[1037] }),
  .A3({ S22947 }),
  .ZN({ S22948 })
);
NAND3_X1 #() 
NAND3_X1_4194_ (
  .A1({ S77 }),
  .A2({ S22660 }),
  .A3({ S22686 }),
  .ZN({ S22949 })
);
NAND3_X1 #() 
NAND3_X1_4195_ (
  .A1({ S22949 }),
  .A2({ S22733 }),
  .A3({ S22636 }),
  .ZN({ S22950 })
);
NAND2_X1 #() 
NAND2_X1_3958_ (
  .A1({ S22844 }),
  .A2({ S25957[1036] }),
  .ZN({ S22951 })
);
OAI211_X1 #() 
OAI211_X1_1364_ (
  .A({ S21015 }),
  .B({ S22950 }),
  .C1({ S22951 }),
  .C2({ S22761 }),
  .ZN({ S22952 })
);
NAND3_X1 #() 
NAND3_X1_4196_ (
  .A1({ S22952 }),
  .A2({ S25957[1038] }),
  .A3({ S22948 }),
  .ZN({ S22953 })
);
NAND3_X1 #() 
NAND3_X1_4197_ (
  .A1({ S22943 }),
  .A2({ S25957[1039] }),
  .A3({ S22953 }),
  .ZN({ S22954 })
);
INV_X1 #() 
INV_X1_1308_ (
  .A({ S22954 }),
  .ZN({ S22955 })
);
NAND3_X1 #() 
NAND3_X1_4198_ (
  .A1({ S22762 }),
  .A2({ S77 }),
  .A3({ S22686 }),
  .ZN({ S22956 })
);
NAND3_X1 #() 
NAND3_X1_4199_ (
  .A1({ S22956 }),
  .A2({ S22678 }),
  .A3({ S25957[1036] }),
  .ZN({ S22957 })
);
AOI21_X1 #() 
AOI21_X1_2120_ (
  .A({ S25957[1035] }),
  .B1({ S22648 }),
  .B2({ S22767 }),
  .ZN({ S22958 })
);
OAI21_X1 #() 
OAI21_X1_2022_ (
  .A({ S22636 }),
  .B1({ S77 }),
  .B2({ S22644 }),
  .ZN({ S22959 })
);
OAI211_X1 #() 
OAI211_X1_1365_ (
  .A({ S22957 }),
  .B({ S21015 }),
  .C1({ S22958 }),
  .C2({ S22959 }),
  .ZN({ S22960 })
);
NAND2_X1 #() 
NAND2_X1_3959_ (
  .A1({ S22665 }),
  .A2({ S25957[1034] }),
  .ZN({ S22961 })
);
AOI21_X1 #() 
AOI21_X1_2121_ (
  .A({ S25957[1035] }),
  .B1({ S22851 }),
  .B2({ S22961 }),
  .ZN({ S22962 })
);
NAND2_X1 #() 
NAND2_X1_3960_ (
  .A1({ S22884 }),
  .A2({ S22636 }),
  .ZN({ S22963 })
);
INV_X1 #() 
INV_X1_1309_ (
  .A({ S124 }),
  .ZN({ S22964 })
);
OAI21_X1 #() 
OAI21_X1_2023_ (
  .A({ S25957[1036] }),
  .B1({ S22964 }),
  .B2({ S25957[1034] }),
  .ZN({ S22965 })
);
OAI211_X1 #() 
OAI211_X1_1366_ (
  .A({ S25957[1037] }),
  .B({ S22965 }),
  .C1({ S22962 }),
  .C2({ S22963 }),
  .ZN({ S22966 })
);
AOI21_X1 #() 
AOI21_X1_2122_ (
  .A({ S22635 }),
  .B1({ S22966 }),
  .B2({ S22960 }),
  .ZN({ S22967 })
);
INV_X1 #() 
INV_X1_1310_ (
  .A({ S22967 }),
  .ZN({ S22968 })
);
NOR2_X1 #() 
NOR2_X1_1004_ (
  .A1({ S22718 }),
  .A2({ S22788 }),
  .ZN({ S22969 })
);
AOI22_X1 #() 
AOI22_X1_444_ (
  .A1({ S22665 }),
  .A2({ S22683 }),
  .B1({ S21186 }),
  .B2({ S21185 }),
  .ZN({ S22970 })
);
AOI21_X1 #() 
AOI21_X1_2123_ (
  .A({ S25957[1035] }),
  .B1({ S22762 }),
  .B2({ S22840 }),
  .ZN({ S22971 })
);
OAI21_X1 #() 
OAI21_X1_2024_ (
  .A({ S22636 }),
  .B1({ S22971 }),
  .B2({ S22970 }),
  .ZN({ S22972 })
);
OAI21_X1 #() 
OAI21_X1_2025_ (
  .A({ S22972 }),
  .B1({ S22951 }),
  .B2({ S22969 }),
  .ZN({ S22973 })
);
NAND3_X1 #() 
NAND3_X1_4200_ (
  .A1({ S22712 }),
  .A2({ S25957[1036] }),
  .A3({ S22869 }),
  .ZN({ S22974 })
);
NOR2_X1 #() 
NOR2_X1_1005_ (
  .A1({ S25957[1035] }),
  .A2({ S22632 }),
  .ZN({ S22975 })
);
OAI21_X1 #() 
OAI21_X1_2026_ (
  .A({ S22636 }),
  .B1({ S22852 }),
  .B2({ S22975 }),
  .ZN({ S22976 })
);
NAND3_X1 #() 
NAND3_X1_4201_ (
  .A1({ S22976 }),
  .A2({ S25957[1037] }),
  .A3({ S22974 }),
  .ZN({ S22977 })
);
OAI211_X1 #() 
OAI211_X1_1367_ (
  .A({ S22977 }),
  .B({ S22635 }),
  .C1({ S22973 }),
  .C2({ S25957[1037] }),
  .ZN({ S22978 })
);
AOI21_X1 #() 
AOI21_X1_2124_ (
  .A({ S25957[1039] }),
  .B1({ S22978 }),
  .B2({ S22968 }),
  .ZN({ S22979 })
);
OAI21_X1 #() 
OAI21_X1_2027_ (
  .A({ S9075 }),
  .B1({ S22955 }),
  .B2({ S22979 }),
  .ZN({ S22980 })
);
INV_X1 #() 
INV_X1_1311_ (
  .A({ S22979 }),
  .ZN({ S22981 })
);
NAND3_X1 #() 
NAND3_X1_4202_ (
  .A1({ S22981 }),
  .A2({ S25957[1236] }),
  .A3({ S22954 }),
  .ZN({ S22982 })
);
AOI21_X1 #() 
AOI21_X1_2125_ (
  .A({ S9119 }),
  .B1({ S22982 }),
  .B2({ S22980 }),
  .ZN({ S22983 })
);
AND3_X1 #() 
AND3_X1_150_ (
  .A1({ S22982 }),
  .A2({ S22980 }),
  .A3({ S9119 }),
  .ZN({ S22984 })
);
NOR2_X1 #() 
NOR2_X1_1006_ (
  .A1({ S22984 }),
  .A2({ S22983 }),
  .ZN({ S22985 })
);
INV_X1 #() 
INV_X1_1312_ (
  .A({ S22985 }),
  .ZN({ S25957[916] })
);
NAND2_X1 #() 
NAND2_X1_3961_ (
  .A1({ S20541 }),
  .A2({ S20545 }),
  .ZN({ S22986 })
);
INV_X1 #() 
INV_X1_1313_ (
  .A({ S22986 }),
  .ZN({ S25957[1075] })
);
NAND3_X1 #() 
NAND3_X1_4203_ (
  .A1({ S22898 }),
  .A2({ S77 }),
  .A3({ S22660 }),
  .ZN({ S22987 })
);
NAND3_X1 #() 
NAND3_X1_4204_ (
  .A1({ S22646 }),
  .A2({ S25957[1035] }),
  .A3({ S22937 }),
  .ZN({ S22988 })
);
AOI21_X1 #() 
AOI21_X1_2126_ (
  .A({ S25957[1036] }),
  .B1({ S22988 }),
  .B2({ S22987 }),
  .ZN({ S22989 })
);
NAND2_X1 #() 
NAND2_X1_3962_ (
  .A1({ S22665 }),
  .A2({ S22683 }),
  .ZN({ S22990 })
);
AOI21_X1 #() 
AOI21_X1_2127_ (
  .A({ S22636 }),
  .B1({ S22990 }),
  .B2({ S25957[1035] }),
  .ZN({ S22991 })
);
NAND3_X1 #() 
NAND3_X1_4205_ (
  .A1({ S77 }),
  .A2({ S22739 }),
  .A3({ S22656 }),
  .ZN({ S22992 })
);
AND2_X1 #() 
AND2_X1_247_ (
  .A1({ S22991 }),
  .A2({ S22992 }),
  .ZN({ S22993 })
);
OAI21_X1 #() 
OAI21_X1_2028_ (
  .A({ S25957[1037] }),
  .B1({ S22993 }),
  .B2({ S22989 }),
  .ZN({ S22994 })
);
NAND3_X1 #() 
NAND3_X1_4206_ (
  .A1({ S22702 }),
  .A2({ S77 }),
  .A3({ S22682 }),
  .ZN({ S22995 })
);
AOI21_X1 #() 
AOI21_X1_2128_ (
  .A({ S22636 }),
  .B1({ S22995 }),
  .B2({ S22861 }),
  .ZN({ S22996 })
);
NOR2_X1 #() 
NOR2_X1_1007_ (
  .A1({ S22959 }),
  .A2({ S22806 }),
  .ZN({ S22997 })
);
OAI21_X1 #() 
OAI21_X1_2029_ (
  .A({ S21015 }),
  .B1({ S22996 }),
  .B2({ S22997 }),
  .ZN({ S22998 })
);
NAND3_X1 #() 
NAND3_X1_4207_ (
  .A1({ S22998 }),
  .A2({ S22994 }),
  .A3({ S25957[1038] }),
  .ZN({ S22999 })
);
AOI22_X1 #() 
AOI22_X1_445_ (
  .A1({ S21185 }),
  .A2({ S21186 }),
  .B1({ S22839 }),
  .B2({ S25957[1034] }),
  .ZN({ S23000 })
);
AOI22_X1 #() 
AOI22_X1_446_ (
  .A1({ S22851 }),
  .A2({ S23000 }),
  .B1({ S77 }),
  .B2({ S22773 }),
  .ZN({ S23001 })
);
NAND2_X1 #() 
NAND2_X1_3963_ (
  .A1({ S22663 }),
  .A2({ S22648 }),
  .ZN({ S23002 })
);
AOI21_X1 #() 
AOI21_X1_2129_ (
  .A({ S22687 }),
  .B1({ S23002 }),
  .B2({ S22632 }),
  .ZN({ S23003 })
);
NAND3_X1 #() 
NAND3_X1_4208_ (
  .A1({ S22889 }),
  .A2({ S25957[1035] }),
  .A3({ S22783 }),
  .ZN({ S23004 })
);
OAI211_X1 #() 
OAI211_X1_1368_ (
  .A({ S22636 }),
  .B({ S23004 }),
  .C1({ S23003 }),
  .C2({ S25957[1035] }),
  .ZN({ S23005 })
);
OAI211_X1 #() 
OAI211_X1_1369_ (
  .A({ S23005 }),
  .B({ S25957[1037] }),
  .C1({ S23001 }),
  .C2({ S22636 }),
  .ZN({ S23006 })
);
NAND2_X1 #() 
NAND2_X1_3964_ (
  .A1({ S22693 }),
  .A2({ S25957[1035] }),
  .ZN({ S23007 })
);
NAND3_X1 #() 
NAND3_X1_4209_ (
  .A1({ S23007 }),
  .A2({ S25957[1036] }),
  .A3({ S22949 }),
  .ZN({ S23008 })
);
NOR2_X1 #() 
NOR2_X1_1008_ (
  .A1({ S22806 }),
  .A2({ S25957[1035] }),
  .ZN({ S23009 })
);
AOI21_X1 #() 
AOI21_X1_2130_ (
  .A({ S77 }),
  .B1({ S22889 }),
  .B2({ S22937 }),
  .ZN({ S23010 })
);
OAI21_X1 #() 
OAI21_X1_2030_ (
  .A({ S22636 }),
  .B1({ S23010 }),
  .B2({ S23009 }),
  .ZN({ S23011 })
);
NAND2_X1 #() 
NAND2_X1_3965_ (
  .A1({ S23011 }),
  .A2({ S23008 }),
  .ZN({ S23012 })
);
NAND2_X1 #() 
NAND2_X1_3966_ (
  .A1({ S23012 }),
  .A2({ S21015 }),
  .ZN({ S23013 })
);
NAND3_X1 #() 
NAND3_X1_4210_ (
  .A1({ S23013 }),
  .A2({ S23006 }),
  .A3({ S22635 }),
  .ZN({ S23014 })
);
NAND3_X1 #() 
NAND3_X1_4211_ (
  .A1({ S23014 }),
  .A2({ S22999 }),
  .A3({ S25957[1039] }),
  .ZN({ S23015 })
);
AND2_X1 #() 
AND2_X1_248_ (
  .A1({ S22738 }),
  .A2({ S22774 }),
  .ZN({ S23016 })
);
NOR3_X1 #() 
NOR3_X1_136_ (
  .A1({ S77 }),
  .A2({ S25957[1032] }),
  .A3({ S22696 }),
  .ZN({ S23017 })
);
NAND4_X1 #() 
NAND4_X1_458_ (
  .A1({ S22656 }),
  .A2({ S22647 }),
  .A3({ S21186 }),
  .A4({ S21185 }),
  .ZN({ S23018 })
);
NAND2_X1 #() 
NAND2_X1_3967_ (
  .A1({ S23018 }),
  .A2({ S22636 }),
  .ZN({ S23019 })
);
OAI21_X1 #() 
OAI21_X1_2031_ (
  .A({ S25957[1037] }),
  .B1({ S23019 }),
  .B2({ S23017 }),
  .ZN({ S23020 })
);
OAI21_X1 #() 
OAI21_X1_2032_ (
  .A({ S22650 }),
  .B1({ S22819 }),
  .B2({ S22681 }),
  .ZN({ S23021 })
);
NAND4_X1 #() 
NAND4_X1_459_ (
  .A1({ S21185 }),
  .A2({ S21186 }),
  .A3({ S22632 }),
  .A4({ S22648 }),
  .ZN({ S23022 })
);
AOI21_X1 #() 
AOI21_X1_2131_ (
  .A({ S25957[1037] }),
  .B1({ S23022 }),
  .B2({ S25957[1036] }),
  .ZN({ S23023 })
);
OAI21_X1 #() 
OAI21_X1_2033_ (
  .A({ S23023 }),
  .B1({ S23021 }),
  .B2({ S25957[1036] }),
  .ZN({ S23024 })
);
OAI211_X1 #() 
OAI211_X1_1370_ (
  .A({ S23024 }),
  .B({ S25957[1038] }),
  .C1({ S23016 }),
  .C2({ S23020 }),
  .ZN({ S23025 })
);
NAND3_X1 #() 
NAND3_X1_4212_ (
  .A1({ S22818 }),
  .A2({ S22660 }),
  .A3({ S22711 }),
  .ZN({ S23026 })
);
OAI211_X1 #() 
OAI211_X1_1371_ (
  .A({ S22769 }),
  .B({ S25957[1036] }),
  .C1({ S25957[1035] }),
  .C2({ S22876 }),
  .ZN({ S23027 })
);
OAI211_X1 #() 
OAI211_X1_1372_ (
  .A({ S23027 }),
  .B({ S25957[1037] }),
  .C1({ S25957[1036] }),
  .C2({ S23026 }),
  .ZN({ S23028 })
);
NOR4_X1 #() 
NOR4_X1_3_ (
  .A1({ S22703 }),
  .A2({ S22809 }),
  .A3({ S22768 }),
  .A4({ S25957[1036] }),
  .ZN({ S23029 })
);
NAND3_X1 #() 
NAND3_X1_4213_ (
  .A1({ S22898 }),
  .A2({ S25957[1035] }),
  .A3({ S22648 }),
  .ZN({ S23030 })
);
AND2_X1 #() 
AND2_X1_249_ (
  .A1({ S22820 }),
  .A2({ S23030 }),
  .ZN({ S23031 })
);
OAI21_X1 #() 
OAI21_X1_2034_ (
  .A({ S21015 }),
  .B1({ S23031 }),
  .B2({ S22636 }),
  .ZN({ S23032 })
);
OAI211_X1 #() 
OAI211_X1_1373_ (
  .A({ S22635 }),
  .B({ S23028 }),
  .C1({ S23032 }),
  .C2({ S23029 }),
  .ZN({ S23033 })
);
NAND3_X1 #() 
NAND3_X1_4214_ (
  .A1({ S23033 }),
  .A2({ S22726 }),
  .A3({ S23025 }),
  .ZN({ S23034 })
);
NAND3_X1 #() 
NAND3_X1_4215_ (
  .A1({ S23015 }),
  .A2({ S23034 }),
  .A3({ S25957[1235] }),
  .ZN({ S23035 })
);
OAI21_X1 #() 
OAI21_X1_2035_ (
  .A({ S21015 }),
  .B1({ S22959 }),
  .B2({ S22806 }),
  .ZN({ S23036 })
);
AND2_X1 #() 
AND2_X1_250_ (
  .A1({ S22988 }),
  .A2({ S22987 }),
  .ZN({ S23037 })
);
AOI21_X1 #() 
AOI21_X1_2132_ (
  .A({ S21015 }),
  .B1({ S22991 }),
  .B2({ S22992 }),
  .ZN({ S23038 })
);
OAI21_X1 #() 
OAI21_X1_2036_ (
  .A({ S23038 }),
  .B1({ S23037 }),
  .B2({ S25957[1036] }),
  .ZN({ S23039 })
);
OAI211_X1 #() 
OAI211_X1_1374_ (
  .A({ S23039 }),
  .B({ S25957[1038] }),
  .C1({ S23036 }),
  .C2({ S22996 }),
  .ZN({ S23040 })
);
NOR2_X1 #() 
NOR2_X1_1009_ (
  .A1({ S22767 }),
  .A2({ S22839 }),
  .ZN({ S23041 })
);
AOI21_X1 #() 
AOI21_X1_2133_ (
  .A({ S22636 }),
  .B1({ S22773 }),
  .B2({ S77 }),
  .ZN({ S23042 })
);
OAI21_X1 #() 
OAI21_X1_2037_ (
  .A({ S23042 }),
  .B1({ S23041 }),
  .B2({ S22769 }),
  .ZN({ S23043 })
);
NAND3_X1 #() 
NAND3_X1_4216_ (
  .A1({ S22694 }),
  .A2({ S77 }),
  .A3({ S22686 }),
  .ZN({ S23044 })
);
NAND3_X1 #() 
NAND3_X1_4217_ (
  .A1({ S22810 }),
  .A2({ S25957[1035] }),
  .A3({ S22660 }),
  .ZN({ S23045 })
);
NAND3_X1 #() 
NAND3_X1_4218_ (
  .A1({ S23044 }),
  .A2({ S23045 }),
  .A3({ S22636 }),
  .ZN({ S23046 })
);
NAND3_X1 #() 
NAND3_X1_4219_ (
  .A1({ S23043 }),
  .A2({ S25957[1037] }),
  .A3({ S23046 }),
  .ZN({ S23047 })
);
NAND3_X1 #() 
NAND3_X1_4220_ (
  .A1({ S23011 }),
  .A2({ S21015 }),
  .A3({ S23008 }),
  .ZN({ S23048 })
);
NAND3_X1 #() 
NAND3_X1_4221_ (
  .A1({ S23047 }),
  .A2({ S23048 }),
  .A3({ S22635 }),
  .ZN({ S23049 })
);
NAND3_X1 #() 
NAND3_X1_4222_ (
  .A1({ S23040 }),
  .A2({ S25957[1039] }),
  .A3({ S23049 }),
  .ZN({ S23050 })
);
AOI22_X1 #() 
AOI22_X1_447_ (
  .A1({ S22737 }),
  .A2({ S22694 }),
  .B1({ S25957[1035] }),
  .B2({ S22773 }),
  .ZN({ S23051 })
);
AOI22_X1 #() 
AOI22_X1_448_ (
  .A1({ S85 }),
  .A2({ S22663 }),
  .B1({ S21184 }),
  .B2({ S21181 }),
  .ZN({ S23052 })
);
OAI21_X1 #() 
OAI21_X1_2038_ (
  .A({ S22636 }),
  .B1({ S23017 }),
  .B2({ S23052 }),
  .ZN({ S23053 })
);
OAI211_X1 #() 
OAI211_X1_1375_ (
  .A({ S23053 }),
  .B({ S25957[1037] }),
  .C1({ S23051 }),
  .C2({ S22636 }),
  .ZN({ S23054 })
);
NAND2_X1 #() 
NAND2_X1_3968_ (
  .A1({ S22682 }),
  .A2({ S22663 }),
  .ZN({ S23055 })
);
AOI22_X1 #() 
AOI22_X1_449_ (
  .A1({ S22771 }),
  .A2({ S23055 }),
  .B1({ S22649 }),
  .B2({ S25957[1035] }),
  .ZN({ S23056 })
);
AOI22_X1 #() 
AOI22_X1_450_ (
  .A1({ S25957[1032] }),
  .A2({ S22686 }),
  .B1({ S21184 }),
  .B2({ S21181 }),
  .ZN({ S23057 })
);
NAND2_X1 #() 
NAND2_X1_3969_ (
  .A1({ S23057 }),
  .A2({ S25957[1036] }),
  .ZN({ S23058 })
);
OAI211_X1 #() 
OAI211_X1_1376_ (
  .A({ S21015 }),
  .B({ S23058 }),
  .C1({ S23056 }),
  .C2({ S25957[1036] }),
  .ZN({ S23059 })
);
NAND3_X1 #() 
NAND3_X1_4223_ (
  .A1({ S23054 }),
  .A2({ S23059 }),
  .A3({ S25957[1038] }),
  .ZN({ S23060 })
);
NAND2_X1 #() 
NAND2_X1_3970_ (
  .A1({ S22702 }),
  .A2({ S22645 }),
  .ZN({ S23061 })
);
NAND2_X1 #() 
NAND2_X1_3971_ (
  .A1({ S23061 }),
  .A2({ S77 }),
  .ZN({ S23062 })
);
OAI21_X1 #() 
OAI21_X1_2039_ (
  .A({ S25957[1035] }),
  .B1({ S22731 }),
  .B2({ S22676 }),
  .ZN({ S23063 })
);
AOI21_X1 #() 
AOI21_X1_2134_ (
  .A({ S25957[1037] }),
  .B1({ S23062 }),
  .B2({ S23063 }),
  .ZN({ S23064 })
);
NAND2_X1 #() 
NAND2_X1_3972_ (
  .A1({ S23026 }),
  .A2({ S25957[1037] }),
  .ZN({ S23065 })
);
NAND2_X1 #() 
NAND2_X1_3973_ (
  .A1({ S23065 }),
  .A2({ S22636 }),
  .ZN({ S23066 })
);
NAND4_X1 #() 
NAND4_X1_460_ (
  .A1({ S22848 }),
  .A2({ S21184 }),
  .A3({ S21181 }),
  .A4({ S22634 }),
  .ZN({ S23067 })
);
OAI211_X1 #() 
OAI211_X1_1377_ (
  .A({ S25957[1037] }),
  .B({ S23067 }),
  .C1({ S22702 }),
  .C2({ S25957[1035] }),
  .ZN({ S23068 })
);
NAND3_X1 #() 
NAND3_X1_4224_ (
  .A1({ S22820 }),
  .A2({ S23030 }),
  .A3({ S21015 }),
  .ZN({ S23069 })
);
NAND3_X1 #() 
NAND3_X1_4225_ (
  .A1({ S23069 }),
  .A2({ S23068 }),
  .A3({ S25957[1036] }),
  .ZN({ S23070 })
);
OAI211_X1 #() 
OAI211_X1_1378_ (
  .A({ S23070 }),
  .B({ S22635 }),
  .C1({ S23064 }),
  .C2({ S23066 }),
  .ZN({ S23071 })
);
NAND3_X1 #() 
NAND3_X1_4226_ (
  .A1({ S23060 }),
  .A2({ S23071 }),
  .A3({ S22726 }),
  .ZN({ S23072 })
);
NAND3_X1 #() 
NAND3_X1_4227_ (
  .A1({ S23050 }),
  .A2({ S23072 }),
  .A3({ S20537 }),
  .ZN({ S23073 })
);
NAND3_X1 #() 
NAND3_X1_4228_ (
  .A1({ S23035 }),
  .A2({ S23073 }),
  .A3({ S25957[1075] }),
  .ZN({ S23074 })
);
AOI21_X1 #() 
AOI21_X1_2135_ (
  .A({ S20537 }),
  .B1({ S23050 }),
  .B2({ S23072 }),
  .ZN({ S23075 })
);
AOI21_X1 #() 
AOI21_X1_2136_ (
  .A({ S25957[1235] }),
  .B1({ S23015 }),
  .B2({ S23034 }),
  .ZN({ S23076 })
);
OAI21_X1 #() 
OAI21_X1_2040_ (
  .A({ S22986 }),
  .B1({ S23076 }),
  .B2({ S23075 }),
  .ZN({ S23077 })
);
NAND3_X1 #() 
NAND3_X1_4229_ (
  .A1({ S23077 }),
  .A2({ S25957[1043] }),
  .A3({ S23074 }),
  .ZN({ S23078 })
);
NAND2_X1 #() 
NAND2_X1_3974_ (
  .A1({ S20539 }),
  .A2({ S20538 }),
  .ZN({ S25957[1139] })
);
NAND3_X1 #() 
NAND3_X1_4230_ (
  .A1({ S23015 }),
  .A2({ S23034 }),
  .A3({ S25957[1139] }),
  .ZN({ S23079 })
);
INV_X1 #() 
INV_X1_1314_ (
  .A({ S25957[1139] }),
  .ZN({ S23080 })
);
NAND3_X1 #() 
NAND3_X1_4231_ (
  .A1({ S23050 }),
  .A2({ S23072 }),
  .A3({ S23080 }),
  .ZN({ S23081 })
);
NAND3_X1 #() 
NAND3_X1_4232_ (
  .A1({ S23079 }),
  .A2({ S23081 }),
  .A3({ S20542 }),
  .ZN({ S23082 })
);
NAND3_X1 #() 
NAND3_X1_4233_ (
  .A1({ S23015 }),
  .A2({ S23034 }),
  .A3({ S23080 }),
  .ZN({ S23083 })
);
NAND3_X1 #() 
NAND3_X1_4234_ (
  .A1({ S23050 }),
  .A2({ S23072 }),
  .A3({ S25957[1139] }),
  .ZN({ S23084 })
);
NAND3_X1 #() 
NAND3_X1_4235_ (
  .A1({ S23083 }),
  .A2({ S23084 }),
  .A3({ S25957[1203] }),
  .ZN({ S23085 })
);
NAND3_X1 #() 
NAND3_X1_4236_ (
  .A1({ S23082 }),
  .A2({ S23085 }),
  .A3({ S74 }),
  .ZN({ S23086 })
);
NAND2_X1 #() 
NAND2_X1_3975_ (
  .A1({ S23078 }),
  .A2({ S23086 }),
  .ZN({ S86 })
);
NAND3_X1 #() 
NAND3_X1_4237_ (
  .A1({ S23077 }),
  .A2({ S74 }),
  .A3({ S23074 }),
  .ZN({ S23087 })
);
NAND3_X1 #() 
NAND3_X1_4238_ (
  .A1({ S23082 }),
  .A2({ S23085 }),
  .A3({ S25957[1043] }),
  .ZN({ S23088 })
);
NAND2_X1 #() 
NAND2_X1_3976_ (
  .A1({ S23087 }),
  .A2({ S23088 }),
  .ZN({ S25957[915] })
);
NOR2_X1 #() 
NOR2_X1_1010_ (
  .A1({ S10357 }),
  .A2({ S10368 }),
  .ZN({ S25957[1200] })
);
NAND2_X1 #() 
NAND2_X1_3977_ (
  .A1({ S20610 }),
  .A2({ S20611 }),
  .ZN({ S25957[1136] })
);
NAND2_X1 #() 
NAND2_X1_3978_ (
  .A1({ S22684 }),
  .A2({ S22682 }),
  .ZN({ S23089 })
);
NAND2_X1 #() 
NAND2_X1_3979_ (
  .A1({ S23089 }),
  .A2({ S77 }),
  .ZN({ S23090 })
);
NAND3_X1 #() 
NAND3_X1_4239_ (
  .A1({ S22711 }),
  .A2({ S25957[1035] }),
  .A3({ S22648 }),
  .ZN({ S23091 })
);
NAND3_X1 #() 
NAND3_X1_4240_ (
  .A1({ S23090 }),
  .A2({ S22636 }),
  .A3({ S23091 }),
  .ZN({ S23092 })
);
NAND2_X1 #() 
NAND2_X1_3980_ (
  .A1({ S22868 }),
  .A2({ S25957[1035] }),
  .ZN({ S23093 })
);
OAI211_X1 #() 
OAI211_X1_1379_ (
  .A({ S23093 }),
  .B({ S25957[1036] }),
  .C1({ S22655 }),
  .C2({ S25957[1035] }),
  .ZN({ S23094 })
);
NAND3_X1 #() 
NAND3_X1_4241_ (
  .A1({ S23092 }),
  .A2({ S25957[1037] }),
  .A3({ S23094 }),
  .ZN({ S23095 })
);
NAND4_X1 #() 
NAND4_X1_461_ (
  .A1({ S22884 }),
  .A2({ S22778 }),
  .A3({ S22727 }),
  .A4({ S22636 }),
  .ZN({ S23096 })
);
NAND3_X1 #() 
NAND3_X1_4242_ (
  .A1({ S22898 }),
  .A2({ S25957[1035] }),
  .A3({ S25957[1034] }),
  .ZN({ S23097 })
);
NAND3_X1 #() 
NAND3_X1_4243_ (
  .A1({ S22931 }),
  .A2({ S25957[1036] }),
  .A3({ S23097 }),
  .ZN({ S23098 })
);
NAND3_X1 #() 
NAND3_X1_4244_ (
  .A1({ S23098 }),
  .A2({ S23096 }),
  .A3({ S21015 }),
  .ZN({ S23099 })
);
NAND3_X1 #() 
NAND3_X1_4245_ (
  .A1({ S23095 }),
  .A2({ S23099 }),
  .A3({ S25957[1038] }),
  .ZN({ S23100 })
);
AND2_X1 #() 
AND2_X1_251_ (
  .A1({ S22739 }),
  .A2({ S22682 }),
  .ZN({ S23101 })
);
OAI211_X1 #() 
OAI211_X1_1380_ (
  .A({ S25957[1036] }),
  .B({ S22769 }),
  .C1({ S23101 }),
  .C2({ S25957[1035] }),
  .ZN({ S23102 })
);
NAND4_X1 #() 
NAND4_X1_462_ (
  .A1({ S22888 }),
  .A2({ S22926 }),
  .A3({ S22946 }),
  .A4({ S22636 }),
  .ZN({ S23103 })
);
NAND3_X1 #() 
NAND3_X1_4246_ (
  .A1({ S23102 }),
  .A2({ S25957[1037] }),
  .A3({ S23103 }),
  .ZN({ S23104 })
);
NAND2_X1 #() 
NAND2_X1_3981_ (
  .A1({ S22791 }),
  .A2({ S77 }),
  .ZN({ S23105 })
);
NAND2_X1 #() 
NAND2_X1_3982_ (
  .A1({ S22858 }),
  .A2({ S22663 }),
  .ZN({ S23106 })
);
AOI21_X1 #() 
AOI21_X1_2137_ (
  .A({ S25957[1036] }),
  .B1({ S23106 }),
  .B2({ S23105 }),
  .ZN({ S23107 })
);
NAND2_X1 #() 
NAND2_X1_3983_ (
  .A1({ S25957[1035] }),
  .A2({ S22663 }),
  .ZN({ S23108 })
);
OAI21_X1 #() 
OAI21_X1_2041_ (
  .A({ S77 }),
  .B1({ S22767 }),
  .B2({ S22839 }),
  .ZN({ S23109 })
);
AOI21_X1 #() 
AOI21_X1_2138_ (
  .A({ S22636 }),
  .B1({ S23109 }),
  .B2({ S23108 }),
  .ZN({ S23110 })
);
OAI21_X1 #() 
OAI21_X1_2042_ (
  .A({ S21015 }),
  .B1({ S23107 }),
  .B2({ S23110 }),
  .ZN({ S23111 })
);
NAND3_X1 #() 
NAND3_X1_4247_ (
  .A1({ S23111 }),
  .A2({ S23104 }),
  .A3({ S22635 }),
  .ZN({ S23112 })
);
NAND3_X1 #() 
NAND3_X1_4248_ (
  .A1({ S23112 }),
  .A2({ S23100 }),
  .A3({ S25957[1039] }),
  .ZN({ S23113 })
);
NAND2_X1 #() 
NAND2_X1_3984_ (
  .A1({ S22797 }),
  .A2({ S77 }),
  .ZN({ S23114 })
);
NAND2_X1 #() 
NAND2_X1_3985_ (
  .A1({ S22704 }),
  .A2({ S22683 }),
  .ZN({ S23115 })
);
AOI22_X1 #() 
AOI22_X1_451_ (
  .A1({ S21185 }),
  .A2({ S21186 }),
  .B1({ S22648 }),
  .B2({ S22634 }),
  .ZN({ S23116 })
);
AOI21_X1 #() 
AOI21_X1_2139_ (
  .A({ S22636 }),
  .B1({ S23116 }),
  .B2({ S23115 }),
  .ZN({ S23117 })
);
NAND3_X1 #() 
NAND3_X1_4249_ (
  .A1({ S22686 }),
  .A2({ S21181 }),
  .A3({ S21184 }),
  .ZN({ S23118 })
);
NAND4_X1 #() 
NAND4_X1_463_ (
  .A1({ S21185 }),
  .A2({ S21186 }),
  .A3({ S22633 }),
  .A4({ S22644 }),
  .ZN({ S23119 })
);
OAI21_X1 #() 
OAI21_X1_2043_ (
  .A({ S23119 }),
  .B1({ S23118 }),
  .B2({ S22791 }),
  .ZN({ S23120 })
);
AOI22_X1 #() 
AOI22_X1_452_ (
  .A1({ S23117 }),
  .A2({ S23114 }),
  .B1({ S23120 }),
  .B2({ S22636 }),
  .ZN({ S23121 })
);
NAND2_X1 #() 
NAND2_X1_3986_ (
  .A1({ S77 }),
  .A2({ S22937 }),
  .ZN({ S23122 })
);
NAND3_X1 #() 
NAND3_X1_4250_ (
  .A1({ S22884 }),
  .A2({ S23122 }),
  .A3({ S22636 }),
  .ZN({ S23123 })
);
NAND4_X1 #() 
NAND4_X1_464_ (
  .A1({ S22880 }),
  .A2({ S22783 }),
  .A3({ S22779 }),
  .A4({ S25957[1036] }),
  .ZN({ S23124 })
);
NAND3_X1 #() 
NAND3_X1_4251_ (
  .A1({ S23123 }),
  .A2({ S23124 }),
  .A3({ S21015 }),
  .ZN({ S23125 })
);
OAI211_X1 #() 
OAI211_X1_1381_ (
  .A({ S25957[1038] }),
  .B({ S23125 }),
  .C1({ S23121 }),
  .C2({ S21015 }),
  .ZN({ S23126 })
);
OAI21_X1 #() 
OAI21_X1_2044_ (
  .A({ S77 }),
  .B1({ S22930 }),
  .B2({ S22895 }),
  .ZN({ S23127 })
);
NAND3_X1 #() 
NAND3_X1_4252_ (
  .A1({ S23127 }),
  .A2({ S23007 }),
  .A3({ S25957[1036] }),
  .ZN({ S23128 })
);
NAND3_X1 #() 
NAND3_X1_4253_ (
  .A1({ S22711 }),
  .A2({ S22762 }),
  .A3({ S77 }),
  .ZN({ S23129 })
);
OAI21_X1 #() 
OAI21_X1_2045_ (
  .A({ S25957[1035] }),
  .B1({ S22895 }),
  .B2({ S22839 }),
  .ZN({ S23130 })
);
NAND3_X1 #() 
NAND3_X1_4254_ (
  .A1({ S23129 }),
  .A2({ S23130 }),
  .A3({ S22636 }),
  .ZN({ S23131 })
);
NAND3_X1 #() 
NAND3_X1_4255_ (
  .A1({ S23128 }),
  .A2({ S23131 }),
  .A3({ S21015 }),
  .ZN({ S23132 })
);
INV_X1 #() 
INV_X1_1315_ (
  .A({ S22900 }),
  .ZN({ S23133 })
);
OAI211_X1 #() 
OAI211_X1_1382_ (
  .A({ S22881 }),
  .B({ S25957[1036] }),
  .C1({ S22839 }),
  .C2({ S22718 }),
  .ZN({ S23134 })
);
NAND2_X1 #() 
NAND2_X1_3987_ (
  .A1({ S22660 }),
  .A2({ S22683 }),
  .ZN({ S23135 })
);
OAI21_X1 #() 
OAI21_X1_2046_ (
  .A({ S22636 }),
  .B1({ S22760 }),
  .B2({ S23135 }),
  .ZN({ S23136 })
);
OAI211_X1 #() 
OAI211_X1_1383_ (
  .A({ S23134 }),
  .B({ S25957[1037] }),
  .C1({ S23133 }),
  .C2({ S23136 }),
  .ZN({ S23137 })
);
NAND3_X1 #() 
NAND3_X1_4256_ (
  .A1({ S23132 }),
  .A2({ S23137 }),
  .A3({ S22635 }),
  .ZN({ S23138 })
);
NAND3_X1 #() 
NAND3_X1_4257_ (
  .A1({ S23126 }),
  .A2({ S23138 }),
  .A3({ S22726 }),
  .ZN({ S23139 })
);
AND3_X1 #() 
AND3_X1_151_ (
  .A1({ S23113 }),
  .A2({ S23139 }),
  .A3({ S25957[1136] }),
  .ZN({ S23140 })
);
AOI21_X1 #() 
AOI21_X1_2140_ (
  .A({ S25957[1136] }),
  .B1({ S23113 }),
  .B2({ S23139 }),
  .ZN({ S23141 })
);
OAI21_X1 #() 
OAI21_X1_2047_ (
  .A({ S25957[1200] }),
  .B1({ S23140 }),
  .B2({ S23141 }),
  .ZN({ S23142 })
);
INV_X1 #() 
INV_X1_1316_ (
  .A({ S25957[1200] }),
  .ZN({ S23143 })
);
NAND3_X1 #() 
NAND3_X1_4258_ (
  .A1({ S23113 }),
  .A2({ S23139 }),
  .A3({ S25957[1136] }),
  .ZN({ S23144 })
);
INV_X1 #() 
INV_X1_1317_ (
  .A({ S25957[1136] }),
  .ZN({ S23145 })
);
INV_X1 #() 
INV_X1_1318_ (
  .A({ S23135 }),
  .ZN({ S23146 })
);
AOI22_X1 #() 
AOI22_X1_453_ (
  .A1({ S22894 }),
  .A2({ S23146 }),
  .B1({ S22899 }),
  .B2({ S22898 }),
  .ZN({ S23147 })
);
AOI22_X1 #() 
AOI22_X1_454_ (
  .A1({ S85 }),
  .A2({ S22648 }),
  .B1({ S21184 }),
  .B2({ S21181 }),
  .ZN({ S23148 })
);
OAI21_X1 #() 
OAI21_X1_2048_ (
  .A({ S25957[1036] }),
  .B1({ S23148 }),
  .B2({ S22970 }),
  .ZN({ S23149 })
);
OAI211_X1 #() 
OAI211_X1_1384_ (
  .A({ S23149 }),
  .B({ S22635 }),
  .C1({ S23147 }),
  .C2({ S25957[1036] }),
  .ZN({ S23150 })
);
NAND4_X1 #() 
NAND4_X1_465_ (
  .A1({ S25957[1035] }),
  .A2({ S22889 }),
  .A3({ S22645 }),
  .A4({ S22937 }),
  .ZN({ S23151 })
);
NAND3_X1 #() 
NAND3_X1_4259_ (
  .A1({ S23151 }),
  .A2({ S25957[1036] }),
  .A3({ S23114 }),
  .ZN({ S23152 })
);
NAND2_X1 #() 
NAND2_X1_3988_ (
  .A1({ S23120 }),
  .A2({ S22636 }),
  .ZN({ S23153 })
);
NAND3_X1 #() 
NAND3_X1_4260_ (
  .A1({ S23153 }),
  .A2({ S23152 }),
  .A3({ S25957[1038] }),
  .ZN({ S23154 })
);
AOI21_X1 #() 
AOI21_X1_2141_ (
  .A({ S25957[1039] }),
  .B1({ S23150 }),
  .B2({ S23154 }),
  .ZN({ S23155 })
);
NOR2_X1 #() 
NOR2_X1_1011_ (
  .A1({ S22961 }),
  .A2({ S77 }),
  .ZN({ S23156 })
);
OAI21_X1 #() 
OAI21_X1_2049_ (
  .A({ S25957[1036] }),
  .B1({ S22971 }),
  .B2({ S23156 }),
  .ZN({ S23157 })
);
OAI21_X1 #() 
OAI21_X1_2050_ (
  .A({ S22636 }),
  .B1({ S22685 }),
  .B2({ S22969 }),
  .ZN({ S23158 })
);
NAND3_X1 #() 
NAND3_X1_4261_ (
  .A1({ S23158 }),
  .A2({ S23157 }),
  .A3({ S25957[1038] }),
  .ZN({ S23159 })
);
NAND4_X1 #() 
NAND4_X1_466_ (
  .A1({ S21185 }),
  .A2({ S21186 }),
  .A3({ S22663 }),
  .A4({ S22633 }),
  .ZN({ S23160 })
);
OAI211_X1 #() 
OAI211_X1_1385_ (
  .A({ S25957[1036] }),
  .B({ S23160 }),
  .C1({ S23057 }),
  .C2({ S23000 }),
  .ZN({ S23161 })
);
AND2_X1 #() 
AND2_X1_252_ (
  .A1({ S77 }),
  .A2({ S22653 }),
  .ZN({ S23162 })
);
AOI21_X1 #() 
AOI21_X1_2142_ (
  .A({ S77 }),
  .B1({ S22711 }),
  .B2({ S22739 }),
  .ZN({ S23163 })
);
OAI21_X1 #() 
OAI21_X1_2051_ (
  .A({ S22636 }),
  .B1({ S23163 }),
  .B2({ S23162 }),
  .ZN({ S23164 })
);
NAND3_X1 #() 
NAND3_X1_4262_ (
  .A1({ S23164 }),
  .A2({ S22635 }),
  .A3({ S23161 }),
  .ZN({ S23165 })
);
AOI21_X1 #() 
AOI21_X1_2143_ (
  .A({ S22726 }),
  .B1({ S23159 }),
  .B2({ S23165 }),
  .ZN({ S23166 })
);
OAI21_X1 #() 
OAI21_X1_2052_ (
  .A({ S25957[1037] }),
  .B1({ S23166 }),
  .B2({ S23155 }),
  .ZN({ S23167 })
);
AOI21_X1 #() 
AOI21_X1_2144_ (
  .A({ S25957[1035] }),
  .B1({ S22646 }),
  .B2({ S22937 }),
  .ZN({ S23168 })
);
INV_X1 #() 
INV_X1_1319_ (
  .A({ S23097 }),
  .ZN({ S23169 })
);
OAI21_X1 #() 
OAI21_X1_2053_ (
  .A({ S25957[1036] }),
  .B1({ S23169 }),
  .B2({ S23168 }),
  .ZN({ S23170 })
);
NOR2_X1 #() 
NOR2_X1_1012_ (
  .A1({ S22818 }),
  .A2({ S23135 }),
  .ZN({ S23171 })
);
OAI21_X1 #() 
OAI21_X1_2054_ (
  .A({ S22636 }),
  .B1({ S23171 }),
  .B2({ S22885 }),
  .ZN({ S23172 })
);
NAND3_X1 #() 
NAND3_X1_4263_ (
  .A1({ S23170 }),
  .A2({ S25957[1038] }),
  .A3({ S23172 }),
  .ZN({ S23173 })
);
AOI22_X1 #() 
AOI22_X1_455_ (
  .A1({ S22858 }),
  .A2({ S22663 }),
  .B1({ S22791 }),
  .B2({ S77 }),
  .ZN({ S23174 })
);
OAI211_X1 #() 
OAI211_X1_1386_ (
  .A({ S25957[1036] }),
  .B({ S22782 }),
  .C1({ S22851 }),
  .C2({ S25957[1035] }),
  .ZN({ S23175 })
);
OAI211_X1 #() 
OAI211_X1_1387_ (
  .A({ S23175 }),
  .B({ S22635 }),
  .C1({ S25957[1036] }),
  .C2({ S23174 }),
  .ZN({ S23176 })
);
AOI21_X1 #() 
AOI21_X1_2145_ (
  .A({ S22726 }),
  .B1({ S23173 }),
  .B2({ S23176 }),
  .ZN({ S23177 })
);
AOI22_X1 #() 
AOI22_X1_456_ (
  .A1({ S22682 }),
  .A2({ S22653 }),
  .B1({ S21184 }),
  .B2({ S21181 }),
  .ZN({ S23178 })
);
AOI21_X1 #() 
AOI21_X1_2146_ (
  .A({ S77 }),
  .B1({ S85 }),
  .B2({ S22889 }),
  .ZN({ S23179 })
);
OAI21_X1 #() 
OAI21_X1_2055_ (
  .A({ S22636 }),
  .B1({ S23179 }),
  .B2({ S23178 }),
  .ZN({ S23180 })
);
AOI21_X1 #() 
AOI21_X1_2147_ (
  .A({ S77 }),
  .B1({ S22898 }),
  .B2({ S22644 }),
  .ZN({ S23181 })
);
AOI22_X1 #() 
AOI22_X1_457_ (
  .A1({ S22889 }),
  .A2({ S22937 }),
  .B1({ S21184 }),
  .B2({ S21181 }),
  .ZN({ S23182 })
);
OAI21_X1 #() 
OAI21_X1_2056_ (
  .A({ S25957[1036] }),
  .B1({ S23181 }),
  .B2({ S23182 }),
  .ZN({ S23183 })
);
NAND3_X1 #() 
NAND3_X1_4264_ (
  .A1({ S23183 }),
  .A2({ S23180 }),
  .A3({ S22635 }),
  .ZN({ S23184 })
);
OAI21_X1 #() 
OAI21_X1_2057_ (
  .A({ S25957[1036] }),
  .B1({ S22780 }),
  .B2({ S22858 }),
  .ZN({ S23185 })
);
AOI22_X1 #() 
AOI22_X1_458_ (
  .A1({ S23146 }),
  .A2({ S22671 }),
  .B1({ S77 }),
  .B2({ S22937 }),
  .ZN({ S23186 })
);
OAI211_X1 #() 
OAI211_X1_1388_ (
  .A({ S25957[1038] }),
  .B({ S23185 }),
  .C1({ S23186 }),
  .C2({ S25957[1036] }),
  .ZN({ S23187 })
);
AOI21_X1 #() 
AOI21_X1_2148_ (
  .A({ S25957[1039] }),
  .B1({ S23184 }),
  .B2({ S23187 }),
  .ZN({ S23188 })
);
OAI21_X1 #() 
OAI21_X1_2058_ (
  .A({ S21015 }),
  .B1({ S23177 }),
  .B2({ S23188 }),
  .ZN({ S23189 })
);
NAND3_X1 #() 
NAND3_X1_4265_ (
  .A1({ S23189 }),
  .A2({ S23167 }),
  .A3({ S23145 }),
  .ZN({ S23190 })
);
NAND3_X1 #() 
NAND3_X1_4266_ (
  .A1({ S23190 }),
  .A2({ S23143 }),
  .A3({ S23144 }),
  .ZN({ S23191 })
);
NAND3_X1 #() 
NAND3_X1_4267_ (
  .A1({ S23142 }),
  .A2({ S23191 }),
  .A3({ S25957[1040] }),
  .ZN({ S23192 })
);
AOI21_X1 #() 
AOI21_X1_2149_ (
  .A({ S20616 }),
  .B1({ S20617 }),
  .B2({ S20618 }),
  .ZN({ S23193 })
);
AND3_X1 #() 
AND3_X1_152_ (
  .A1({ S20618 }),
  .A2({ S20617 }),
  .A3({ S20616 }),
  .ZN({ S23194 })
);
NOR2_X1 #() 
NOR2_X1_1013_ (
  .A1({ S23194 }),
  .A2({ S23193 }),
  .ZN({ S23195 })
);
NOR2_X1 #() 
NOR2_X1_1014_ (
  .A1({ S20609 }),
  .A2({ S20612 }),
  .ZN({ S25957[1072] })
);
INV_X1 #() 
INV_X1_1320_ (
  .A({ S25957[1232] }),
  .ZN({ S23196 })
);
AND3_X1 #() 
AND3_X1_153_ (
  .A1({ S23113 }),
  .A2({ S23139 }),
  .A3({ S23196 }),
  .ZN({ S23197 })
);
AOI21_X1 #() 
AOI21_X1_2150_ (
  .A({ S23196 }),
  .B1({ S23113 }),
  .B2({ S23139 }),
  .ZN({ S23198 })
);
OAI21_X1 #() 
OAI21_X1_2059_ (
  .A({ S25957[1072] }),
  .B1({ S23197 }),
  .B2({ S23198 }),
  .ZN({ S23199 })
);
INV_X1 #() 
INV_X1_1321_ (
  .A({ S25957[1072] }),
  .ZN({ S23200 })
);
NAND3_X1 #() 
NAND3_X1_4268_ (
  .A1({ S23113 }),
  .A2({ S23139 }),
  .A3({ S23196 }),
  .ZN({ S23201 })
);
NAND3_X1 #() 
NAND3_X1_4269_ (
  .A1({ S23189 }),
  .A2({ S23167 }),
  .A3({ S25957[1232] }),
  .ZN({ S23202 })
);
NAND3_X1 #() 
NAND3_X1_4270_ (
  .A1({ S23202 }),
  .A2({ S23200 }),
  .A3({ S23201 }),
  .ZN({ S23203 })
);
NAND3_X1 #() 
NAND3_X1_4271_ (
  .A1({ S23199 }),
  .A2({ S23203 }),
  .A3({ S23195 }),
  .ZN({ S23204 })
);
NAND2_X1 #() 
NAND2_X1_3989_ (
  .A1({ S23192 }),
  .A2({ S23204 }),
  .ZN({ S25957[912] })
);
NOR2_X1 #() 
NOR2_X1_1015_ (
  .A1({ S20671 }),
  .A2({ S20674 }),
  .ZN({ S25957[1073] })
);
OAI211_X1 #() 
OAI211_X1_1389_ (
  .A({ S25957[1036] }),
  .B({ S23160 }),
  .C1({ S22928 }),
  .C2({ S22876 }),
  .ZN({ S23205 })
);
NAND4_X1 #() 
NAND4_X1_467_ (
  .A1({ S22660 }),
  .A2({ S21184 }),
  .A3({ S21181 }),
  .A4({ S22632 }),
  .ZN({ S23206 })
);
OAI211_X1 #() 
OAI211_X1_1390_ (
  .A({ S23206 }),
  .B({ S22636 }),
  .C1({ S23022 }),
  .C2({ S22690 }),
  .ZN({ S23207 })
);
NAND3_X1 #() 
NAND3_X1_4272_ (
  .A1({ S23205 }),
  .A2({ S21015 }),
  .A3({ S23207 }),
  .ZN({ S23208 })
);
NAND2_X1 #() 
NAND2_X1_3990_ (
  .A1({ S84 }),
  .A2({ S22644 }),
  .ZN({ S23209 })
);
AOI21_X1 #() 
AOI21_X1_2151_ (
  .A({ S77 }),
  .B1({ S23209 }),
  .B2({ S22694 }),
  .ZN({ S23210 })
);
NAND3_X1 #() 
NAND3_X1_4273_ (
  .A1({ S22713 }),
  .A2({ S25957[1036] }),
  .A3({ S22861 }),
  .ZN({ S23211 })
);
OAI21_X1 #() 
OAI21_X1_2060_ (
  .A({ S22636 }),
  .B1({ S25957[1035] }),
  .B2({ S22934 }),
  .ZN({ S23212 })
);
OAI211_X1 #() 
OAI211_X1_1391_ (
  .A({ S23211 }),
  .B({ S25957[1037] }),
  .C1({ S23210 }),
  .C2({ S23212 }),
  .ZN({ S23213 })
);
NAND3_X1 #() 
NAND3_X1_4274_ (
  .A1({ S23208 }),
  .A2({ S23213 }),
  .A3({ S25957[1038] }),
  .ZN({ S23214 })
);
OAI211_X1 #() 
OAI211_X1_1392_ (
  .A({ S25957[1036] }),
  .B({ S22798 }),
  .C1({ S22780 }),
  .C2({ S25957[1035] }),
  .ZN({ S23215 })
);
OAI211_X1 #() 
OAI211_X1_1393_ (
  .A({ S23215 }),
  .B({ S21015 }),
  .C1({ S22941 }),
  .C2({ S22705 }),
  .ZN({ S23216 })
);
NAND3_X1 #() 
NAND3_X1_4275_ (
  .A1({ S23018 }),
  .A2({ S22867 }),
  .A3({ S22636 }),
  .ZN({ S23217 })
);
AOI21_X1 #() 
AOI21_X1_2152_ (
  .A({ S77 }),
  .B1({ S22702 }),
  .B2({ S22645 }),
  .ZN({ S23218 })
);
OAI21_X1 #() 
OAI21_X1_2061_ (
  .A({ S25957[1036] }),
  .B1({ S22708 }),
  .B2({ S25957[1035] }),
  .ZN({ S23219 })
);
OAI211_X1 #() 
OAI211_X1_1394_ (
  .A({ S23217 }),
  .B({ S25957[1037] }),
  .C1({ S23218 }),
  .C2({ S23219 }),
  .ZN({ S23220 })
);
NAND3_X1 #() 
NAND3_X1_4276_ (
  .A1({ S23216 }),
  .A2({ S22635 }),
  .A3({ S23220 }),
  .ZN({ S23221 })
);
NAND3_X1 #() 
NAND3_X1_4277_ (
  .A1({ S23221 }),
  .A2({ S23214 }),
  .A3({ S25957[1039] }),
  .ZN({ S23222 })
);
AOI21_X1 #() 
AOI21_X1_2153_ (
  .A({ S25957[1035] }),
  .B1({ S22762 }),
  .B2({ S22645 }),
  .ZN({ S23223 })
);
OAI21_X1 #() 
OAI21_X1_2062_ (
  .A({ S25957[1036] }),
  .B1({ S22666 }),
  .B2({ S22718 }),
  .ZN({ S23224 })
);
NAND4_X1 #() 
NAND4_X1_468_ (
  .A1({ S22760 }),
  .A2({ S22840 }),
  .A3({ S22648 }),
  .A4({ S22636 }),
  .ZN({ S23225 })
);
OAI211_X1 #() 
OAI211_X1_1395_ (
  .A({ S23225 }),
  .B({ S25957[1037] }),
  .C1({ S23224 }),
  .C2({ S23223 }),
  .ZN({ S23226 })
);
NAND3_X1 #() 
NAND3_X1_4278_ (
  .A1({ S22840 }),
  .A2({ S77 }),
  .A3({ S22889 }),
  .ZN({ S23227 })
);
NAND3_X1 #() 
NAND3_X1_4279_ (
  .A1({ S23151 }),
  .A2({ S23227 }),
  .A3({ S25957[1036] }),
  .ZN({ S23228 })
);
NAND3_X1 #() 
NAND3_X1_4280_ (
  .A1({ S23097 }),
  .A2({ S22805 }),
  .A3({ S22636 }),
  .ZN({ S23229 })
);
NAND3_X1 #() 
NAND3_X1_4281_ (
  .A1({ S23228 }),
  .A2({ S23229 }),
  .A3({ S21015 }),
  .ZN({ S23230 })
);
NAND3_X1 #() 
NAND3_X1_4282_ (
  .A1({ S23230 }),
  .A2({ S25957[1038] }),
  .A3({ S23226 }),
  .ZN({ S23231 })
);
AOI21_X1 #() 
AOI21_X1_2154_ (
  .A({ S22636 }),
  .B1({ S23045 }),
  .B2({ S22944 }),
  .ZN({ S23232 })
);
OAI21_X1 #() 
OAI21_X1_2063_ (
  .A({ S25957[1037] }),
  .B1({ S23232 }),
  .B2({ S22721 }),
  .ZN({ S23233 })
);
OAI21_X1 #() 
OAI21_X1_2064_ (
  .A({ S22688 }),
  .B1({ S22819 }),
  .B2({ S22681 }),
  .ZN({ S23234 })
);
NAND3_X1 #() 
NAND3_X1_4283_ (
  .A1({ S22678 }),
  .A2({ S22949 }),
  .A3({ S25957[1036] }),
  .ZN({ S23235 })
);
OAI211_X1 #() 
OAI211_X1_1396_ (
  .A({ S23235 }),
  .B({ S21015 }),
  .C1({ S23234 }),
  .C2({ S25957[1036] }),
  .ZN({ S23236 })
);
NAND3_X1 #() 
NAND3_X1_4284_ (
  .A1({ S23233 }),
  .A2({ S23236 }),
  .A3({ S22635 }),
  .ZN({ S23237 })
);
NAND3_X1 #() 
NAND3_X1_4285_ (
  .A1({ S23237 }),
  .A2({ S22726 }),
  .A3({ S23231 }),
  .ZN({ S23238 })
);
AND3_X1 #() 
AND3_X1_154_ (
  .A1({ S23238 }),
  .A2({ S23222 }),
  .A3({ S25957[1233] }),
  .ZN({ S23239 })
);
AOI21_X1 #() 
AOI21_X1_2155_ (
  .A({ S25957[1233] }),
  .B1({ S23238 }),
  .B2({ S23222 }),
  .ZN({ S23240 })
);
OAI21_X1 #() 
OAI21_X1_2065_ (
  .A({ S25957[1073] }),
  .B1({ S23239 }),
  .B2({ S23240 }),
  .ZN({ S23241 })
);
INV_X1 #() 
INV_X1_1322_ (
  .A({ S25957[1073] }),
  .ZN({ S23242 })
);
NAND3_X1 #() 
NAND3_X1_4286_ (
  .A1({ S23238 }),
  .A2({ S25957[1233] }),
  .A3({ S23222 }),
  .ZN({ S23243 })
);
NAND2_X1 #() 
NAND2_X1_3991_ (
  .A1({ S23230 }),
  .A2({ S23226 }),
  .ZN({ S23244 })
);
NAND2_X1 #() 
NAND2_X1_3992_ (
  .A1({ S23244 }),
  .A2({ S25957[1038] }),
  .ZN({ S23245 })
);
NAND2_X1 #() 
NAND2_X1_3993_ (
  .A1({ S23045 }),
  .A2({ S22944 }),
  .ZN({ S23246 })
);
NAND2_X1 #() 
NAND2_X1_3994_ (
  .A1({ S23246 }),
  .A2({ S25957[1036] }),
  .ZN({ S23247 })
);
NAND3_X1 #() 
NAND3_X1_4287_ (
  .A1({ S22722 }),
  .A2({ S23247 }),
  .A3({ S25957[1037] }),
  .ZN({ S23248 })
);
NAND2_X1 #() 
NAND2_X1_3995_ (
  .A1({ S22660 }),
  .A2({ S22686 }),
  .ZN({ S23249 })
);
NOR2_X1 #() 
NOR2_X1_1016_ (
  .A1({ S23249 }),
  .A2({ S25957[1035] }),
  .ZN({ S23250 })
);
OAI21_X1 #() 
OAI21_X1_2066_ (
  .A({ S25957[1036] }),
  .B1({ S22789 }),
  .B2({ S23250 }),
  .ZN({ S23251 })
);
NAND2_X1 #() 
NAND2_X1_3996_ (
  .A1({ S23234 }),
  .A2({ S22636 }),
  .ZN({ S23252 })
);
NAND3_X1 #() 
NAND3_X1_4288_ (
  .A1({ S23252 }),
  .A2({ S23251 }),
  .A3({ S21015 }),
  .ZN({ S23253 })
);
NAND3_X1 #() 
NAND3_X1_4289_ (
  .A1({ S23248 }),
  .A2({ S23253 }),
  .A3({ S22635 }),
  .ZN({ S23254 })
);
NAND3_X1 #() 
NAND3_X1_4290_ (
  .A1({ S23245 }),
  .A2({ S23254 }),
  .A3({ S22726 }),
  .ZN({ S23255 })
);
NAND2_X1 #() 
NAND2_X1_3997_ (
  .A1({ S23221 }),
  .A2({ S23214 }),
  .ZN({ S23256 })
);
NAND2_X1 #() 
NAND2_X1_3998_ (
  .A1({ S23256 }),
  .A2({ S25957[1039] }),
  .ZN({ S23257 })
);
NAND3_X1 #() 
NAND3_X1_4291_ (
  .A1({ S23255 }),
  .A2({ S23257 }),
  .A3({ S20621 }),
  .ZN({ S23258 })
);
NAND3_X1 #() 
NAND3_X1_4292_ (
  .A1({ S23258 }),
  .A2({ S23242 }),
  .A3({ S23243 }),
  .ZN({ S23259 })
);
NAND3_X1 #() 
NAND3_X1_4293_ (
  .A1({ S23241 }),
  .A2({ S23259 }),
  .A3({ S25957[1041] }),
  .ZN({ S23260 })
);
OAI21_X1 #() 
OAI21_X1_2067_ (
  .A({ S20676 }),
  .B1({ S20671 }),
  .B2({ S20674 }),
  .ZN({ S23261 })
);
NAND3_X1 #() 
NAND3_X1_4294_ (
  .A1({ S20677 }),
  .A2({ S20678 }),
  .A3({ S25957[1169] }),
  .ZN({ S23262 })
);
NAND2_X1 #() 
NAND2_X1_3999_ (
  .A1({ S23261 }),
  .A2({ S23262 }),
  .ZN({ S23263 })
);
NAND2_X1 #() 
NAND2_X1_4000_ (
  .A1({ S20669 }),
  .A2({ S20668 }),
  .ZN({ S25957[1137] })
);
NAND3_X1 #() 
NAND3_X1_4295_ (
  .A1({ S23238 }),
  .A2({ S25957[1137] }),
  .A3({ S23222 }),
  .ZN({ S23264 })
);
INV_X1 #() 
INV_X1_1323_ (
  .A({ S25957[1137] }),
  .ZN({ S23265 })
);
NAND3_X1 #() 
NAND3_X1_4296_ (
  .A1({ S23255 }),
  .A2({ S23257 }),
  .A3({ S23265 }),
  .ZN({ S23266 })
);
NAND3_X1 #() 
NAND3_X1_4297_ (
  .A1({ S23266 }),
  .A2({ S25957[1201] }),
  .A3({ S23264 }),
  .ZN({ S23267 })
);
NAND3_X1 #() 
NAND3_X1_4298_ (
  .A1({ S23238 }),
  .A2({ S23265 }),
  .A3({ S23222 }),
  .ZN({ S23268 })
);
NAND3_X1 #() 
NAND3_X1_4299_ (
  .A1({ S23255 }),
  .A2({ S23257 }),
  .A3({ S25957[1137] }),
  .ZN({ S23269 })
);
NAND3_X1 #() 
NAND3_X1_4300_ (
  .A1({ S23269 }),
  .A2({ S20620 }),
  .A3({ S23268 }),
  .ZN({ S23270 })
);
NAND3_X1 #() 
NAND3_X1_4301_ (
  .A1({ S23267 }),
  .A2({ S23270 }),
  .A3({ S23263 }),
  .ZN({ S23271 })
);
NAND2_X1 #() 
NAND2_X1_4001_ (
  .A1({ S23260 }),
  .A2({ S23271 }),
  .ZN({ S25957[913] })
);
NAND2_X1 #() 
NAND2_X1_4002_ (
  .A1({ S11393 }),
  .A2({ S11421 }),
  .ZN({ S23272 })
);
INV_X1 #() 
INV_X1_1324_ (
  .A({ S23272 }),
  .ZN({ S25957[1234] })
);
NAND3_X1 #() 
NAND3_X1_4302_ (
  .A1({ S22733 }),
  .A2({ S22636 }),
  .A3({ S22940 }),
  .ZN({ S23273 })
);
NOR2_X1 #() 
NOR2_X1_1017_ (
  .A1({ S22650 }),
  .A2({ S22810 }),
  .ZN({ S23274 })
);
OAI21_X1 #() 
OAI21_X1_2068_ (
  .A({ S25957[1036] }),
  .B1({ S22697 }),
  .B2({ S25957[1033] }),
  .ZN({ S23275 })
);
OAI21_X1 #() 
OAI21_X1_2069_ (
  .A({ S23273 }),
  .B1({ S23274 }),
  .B2({ S23275 }),
  .ZN({ S23276 })
);
NAND2_X1 #() 
NAND2_X1_4003_ (
  .A1({ S22961 }),
  .A2({ S25957[1035] }),
  .ZN({ S23277 })
);
OAI211_X1 #() 
OAI211_X1_1397_ (
  .A({ S22636 }),
  .B({ S22664 }),
  .C1({ S23277 }),
  .C2({ S23041 }),
  .ZN({ S23278 })
);
NAND2_X1 #() 
NAND2_X1_4004_ (
  .A1({ S23249 }),
  .A2({ S25957[1035] }),
  .ZN({ S23279 })
);
NAND3_X1 #() 
NAND3_X1_4303_ (
  .A1({ S23090 }),
  .A2({ S25957[1036] }),
  .A3({ S23279 }),
  .ZN({ S23280 })
);
NAND3_X1 #() 
NAND3_X1_4304_ (
  .A1({ S23280 }),
  .A2({ S25957[1037] }),
  .A3({ S23278 }),
  .ZN({ S23281 })
);
OAI211_X1 #() 
OAI211_X1_1398_ (
  .A({ S23281 }),
  .B({ S25957[1038] }),
  .C1({ S25957[1037] }),
  .C2({ S23276 }),
  .ZN({ S23282 })
);
NAND3_X1 #() 
NAND3_X1_4305_ (
  .A1({ S25957[1035] }),
  .A2({ S25957[1032] }),
  .A3({ S22686 }),
  .ZN({ S23283 })
);
OAI211_X1 #() 
OAI211_X1_1399_ (
  .A({ S23283 }),
  .B({ S25957[1036] }),
  .C1({ S22819 }),
  .C2({ S22681 }),
  .ZN({ S23284 })
);
NAND2_X1 #() 
NAND2_X1_4005_ (
  .A1({ S25957[1035] }),
  .A2({ S84 }),
  .ZN({ S23285 })
);
NAND2_X1 #() 
NAND2_X1_4006_ (
  .A1({ S22762 }),
  .A2({ S77 }),
  .ZN({ S23286 })
);
NAND2_X1 #() 
NAND2_X1_4007_ (
  .A1({ S22930 }),
  .A2({ S25957[1035] }),
  .ZN({ S23287 })
);
NAND3_X1 #() 
NAND3_X1_4306_ (
  .A1({ S23287 }),
  .A2({ S23286 }),
  .A3({ S23285 }),
  .ZN({ S23288 })
);
OAI211_X1 #() 
OAI211_X1_1400_ (
  .A({ S23284 }),
  .B({ S25957[1037] }),
  .C1({ S25957[1036] }),
  .C2({ S23288 }),
  .ZN({ S23289 })
);
NAND4_X1 #() 
NAND4_X1_469_ (
  .A1({ S22683 }),
  .A2({ S21184 }),
  .A3({ S21181 }),
  .A4({ S25957[1033] }),
  .ZN({ S23290 })
);
NAND3_X1 #() 
NAND3_X1_4307_ (
  .A1({ S22778 }),
  .A2({ S25957[1036] }),
  .A3({ S23290 }),
  .ZN({ S23291 })
);
OAI211_X1 #() 
OAI211_X1_1401_ (
  .A({ S23291 }),
  .B({ S21015 }),
  .C1({ S22784 }),
  .C2({ S25957[1036] }),
  .ZN({ S23292 })
);
NAND3_X1 #() 
NAND3_X1_4308_ (
  .A1({ S23289 }),
  .A2({ S23292 }),
  .A3({ S22635 }),
  .ZN({ S23293 })
);
NAND3_X1 #() 
NAND3_X1_4309_ (
  .A1({ S23282 }),
  .A2({ S23293 }),
  .A3({ S25957[1039] }),
  .ZN({ S23294 })
);
NAND3_X1 #() 
NAND3_X1_4310_ (
  .A1({ S25957[1035] }),
  .A2({ S22686 }),
  .A3({ S22656 }),
  .ZN({ S23295 })
);
AOI21_X1 #() 
AOI21_X1_2156_ (
  .A({ S22636 }),
  .B1({ S23295 }),
  .B2({ S23022 }),
  .ZN({ S23296 })
);
NAND2_X1 #() 
NAND2_X1_4008_ (
  .A1({ S22647 }),
  .A2({ S25957[1032] }),
  .ZN({ S23297 })
);
NAND2_X1 #() 
NAND2_X1_4009_ (
  .A1({ S77 }),
  .A2({ S23297 }),
  .ZN({ S23298 })
);
NAND3_X1 #() 
NAND3_X1_4311_ (
  .A1({ S22693 }),
  .A2({ S22694 }),
  .A3({ S25957[1035] }),
  .ZN({ S23299 })
);
AOI21_X1 #() 
AOI21_X1_2157_ (
  .A({ S25957[1036] }),
  .B1({ S23299 }),
  .B2({ S23298 }),
  .ZN({ S23300 })
);
OAI21_X1 #() 
OAI21_X1_2070_ (
  .A({ S25957[1037] }),
  .B1({ S23300 }),
  .B2({ S23296 }),
  .ZN({ S23301 })
);
NAND3_X1 #() 
NAND3_X1_4312_ (
  .A1({ S25957[1035] }),
  .A2({ S22783 }),
  .A3({ S22648 }),
  .ZN({ S23302 })
);
NAND2_X1 #() 
NAND2_X1_4010_ (
  .A1({ S22660 }),
  .A2({ S22663 }),
  .ZN({ S23303 })
);
OAI21_X1 #() 
OAI21_X1_2071_ (
  .A({ S77 }),
  .B1({ S23303 }),
  .B2({ S22731 }),
  .ZN({ S23304 })
);
AOI21_X1 #() 
AOI21_X1_2158_ (
  .A({ S22636 }),
  .B1({ S23304 }),
  .B2({ S23302 }),
  .ZN({ S23305 })
);
NAND3_X1 #() 
NAND3_X1_4313_ (
  .A1({ S22646 }),
  .A2({ S77 }),
  .A3({ S22937 }),
  .ZN({ S23306 })
);
AND3_X1 #() 
AND3_X1_155_ (
  .A1({ S23306 }),
  .A2({ S23290 }),
  .A3({ S22636 }),
  .ZN({ S23307 })
);
OAI21_X1 #() 
OAI21_X1_2072_ (
  .A({ S21015 }),
  .B1({ S23305 }),
  .B2({ S23307 }),
  .ZN({ S23308 })
);
NAND3_X1 #() 
NAND3_X1_4314_ (
  .A1({ S23308 }),
  .A2({ S23301 }),
  .A3({ S25957[1038] }),
  .ZN({ S23309 })
);
AOI21_X1 #() 
AOI21_X1_2159_ (
  .A({ S25957[1036] }),
  .B1({ S22877 }),
  .B2({ S77 }),
  .ZN({ S23310 })
);
NAND3_X1 #() 
NAND3_X1_4315_ (
  .A1({ S25957[1035] }),
  .A2({ S22889 }),
  .A3({ S22767 }),
  .ZN({ S23311 })
);
NAND2_X1 #() 
NAND2_X1_4011_ (
  .A1({ S23310 }),
  .A2({ S23311 }),
  .ZN({ S23312 })
);
NAND3_X1 #() 
NAND3_X1_4316_ (
  .A1({ S22840 }),
  .A2({ S25957[1035] }),
  .A3({ S22648 }),
  .ZN({ S23313 })
);
NAND3_X1 #() 
NAND3_X1_4317_ (
  .A1({ S23044 }),
  .A2({ S23313 }),
  .A3({ S25957[1036] }),
  .ZN({ S23314 })
);
NAND3_X1 #() 
NAND3_X1_4318_ (
  .A1({ S23314 }),
  .A2({ S25957[1037] }),
  .A3({ S23312 }),
  .ZN({ S23315 })
);
AOI21_X1 #() 
AOI21_X1_2160_ (
  .A({ S25957[1036] }),
  .B1({ S23089 }),
  .B2({ S77 }),
  .ZN({ S23316 })
);
NAND3_X1 #() 
NAND3_X1_4319_ (
  .A1({ S22939 }),
  .A2({ S25957[1035] }),
  .A3({ S22686 }),
  .ZN({ S23317 })
);
OAI21_X1 #() 
OAI21_X1_2073_ (
  .A({ S23290 }),
  .B1({ S22736 }),
  .B2({ S22934 }),
  .ZN({ S23318 })
);
AOI22_X1 #() 
AOI22_X1_459_ (
  .A1({ S23316 }),
  .A2({ S23317 }),
  .B1({ S23318 }),
  .B2({ S25957[1036] }),
  .ZN({ S23319 })
);
OAI211_X1 #() 
OAI211_X1_1402_ (
  .A({ S23315 }),
  .B({ S22635 }),
  .C1({ S23319 }),
  .C2({ S25957[1037] }),
  .ZN({ S23320 })
);
NAND3_X1 #() 
NAND3_X1_4320_ (
  .A1({ S23309 }),
  .A2({ S22726 }),
  .A3({ S23320 }),
  .ZN({ S23321 })
);
NAND3_X1 #() 
NAND3_X1_4321_ (
  .A1({ S23321 }),
  .A2({ S23294 }),
  .A3({ S25957[1234] }),
  .ZN({ S23322 })
);
NAND2_X1 #() 
NAND2_X1_4012_ (
  .A1({ S23276 }),
  .A2({ S21015 }),
  .ZN({ S23323 })
);
NOR2_X1 #() 
NOR2_X1_1018_ (
  .A1({ S22868 }),
  .A2({ S77 }),
  .ZN({ S23324 })
);
AOI22_X1 #() 
AOI22_X1_460_ (
  .A1({ S23324 }),
  .A2({ S22851 }),
  .B1({ S22663 }),
  .B2({ S77 }),
  .ZN({ S23325 })
);
OAI21_X1 #() 
OAI21_X1_2074_ (
  .A({ S25957[1036] }),
  .B1({ S22685 }),
  .B2({ S22719 }),
  .ZN({ S23326 })
);
OAI211_X1 #() 
OAI211_X1_1403_ (
  .A({ S23326 }),
  .B({ S25957[1037] }),
  .C1({ S23325 }),
  .C2({ S25957[1036] }),
  .ZN({ S23327 })
);
NAND3_X1 #() 
NAND3_X1_4322_ (
  .A1({ S23323 }),
  .A2({ S23327 }),
  .A3({ S25957[1038] }),
  .ZN({ S23328 })
);
OAI21_X1 #() 
OAI21_X1_2075_ (
  .A({ S23283 }),
  .B1({ S22819 }),
  .B2({ S22681 }),
  .ZN({ S23329 })
);
NAND2_X1 #() 
NAND2_X1_4013_ (
  .A1({ S23329 }),
  .A2({ S25957[1036] }),
  .ZN({ S23330 })
);
NAND2_X1 #() 
NAND2_X1_4014_ (
  .A1({ S23288 }),
  .A2({ S22636 }),
  .ZN({ S23331 })
);
NAND3_X1 #() 
NAND3_X1_4323_ (
  .A1({ S23330 }),
  .A2({ S23331 }),
  .A3({ S25957[1037] }),
  .ZN({ S23332 })
);
AND3_X1 #() 
AND3_X1_156_ (
  .A1({ S22926 }),
  .A2({ S22778 }),
  .A3({ S25957[1036] }),
  .ZN({ S23333 })
);
OAI211_X1 #() 
OAI211_X1_1404_ (
  .A({ S21015 }),
  .B({ S22782 }),
  .C1({ S23333 }),
  .C2({ S23310 }),
  .ZN({ S23334 })
);
NAND3_X1 #() 
NAND3_X1_4324_ (
  .A1({ S23332 }),
  .A2({ S23334 }),
  .A3({ S22635 }),
  .ZN({ S23335 })
);
NAND3_X1 #() 
NAND3_X1_4325_ (
  .A1({ S23328 }),
  .A2({ S23335 }),
  .A3({ S25957[1039] }),
  .ZN({ S23336 })
);
NOR2_X1 #() 
NOR2_X1_1019_ (
  .A1({ S23057 }),
  .A2({ S22636 }),
  .ZN({ S23337 })
);
AOI22_X1 #() 
AOI22_X1_461_ (
  .A1({ S22728 }),
  .A2({ S22783 }),
  .B1({ S77 }),
  .B2({ S22696 }),
  .ZN({ S23338 })
);
NAND4_X1 #() 
NAND4_X1_470_ (
  .A1({ S25957[1037] }),
  .A2({ S25957[1035] }),
  .A3({ S22686 }),
  .A4({ S22656 }),
  .ZN({ S23339 })
);
OAI211_X1 #() 
OAI211_X1_1405_ (
  .A({ S23339 }),
  .B({ S23337 }),
  .C1({ S23338 }),
  .C2({ S25957[1037] }),
  .ZN({ S23340 })
);
NOR2_X1 #() 
NOR2_X1_1020_ (
  .A1({ S22778 }),
  .A2({ S22633 }),
  .ZN({ S23341 })
);
NOR3_X1 #() 
NOR3_X1_137_ (
  .A1({ S23341 }),
  .A2({ S22695 }),
  .A3({ S21015 }),
  .ZN({ S23342 })
);
NAND3_X1 #() 
NAND3_X1_4326_ (
  .A1({ S23306 }),
  .A2({ S21015 }),
  .A3({ S23290 }),
  .ZN({ S23343 })
);
NAND2_X1 #() 
NAND2_X1_4015_ (
  .A1({ S23343 }),
  .A2({ S22636 }),
  .ZN({ S23344 })
);
OAI211_X1 #() 
OAI211_X1_1406_ (
  .A({ S23340 }),
  .B({ S25957[1038] }),
  .C1({ S23342 }),
  .C2({ S23344 }),
  .ZN({ S23345 })
);
AND2_X1 #() 
AND2_X1_253_ (
  .A1({ S23314 }),
  .A2({ S23312 }),
  .ZN({ S23346 })
);
NAND2_X1 #() 
NAND2_X1_4016_ (
  .A1({ S23318 }),
  .A2({ S25957[1036] }),
  .ZN({ S23347 })
);
NAND2_X1 #() 
NAND2_X1_4017_ (
  .A1({ S23316 }),
  .A2({ S23317 }),
  .ZN({ S23348 })
);
NAND3_X1 #() 
NAND3_X1_4327_ (
  .A1({ S23348 }),
  .A2({ S21015 }),
  .A3({ S23347 }),
  .ZN({ S23349 })
);
OAI211_X1 #() 
OAI211_X1_1407_ (
  .A({ S23349 }),
  .B({ S22635 }),
  .C1({ S23346 }),
  .C2({ S21015 }),
  .ZN({ S23350 })
);
NAND3_X1 #() 
NAND3_X1_4328_ (
  .A1({ S23350 }),
  .A2({ S23345 }),
  .A3({ S22726 }),
  .ZN({ S23351 })
);
NAND3_X1 #() 
NAND3_X1_4329_ (
  .A1({ S23336 }),
  .A2({ S23351 }),
  .A3({ S23272 }),
  .ZN({ S23352 })
);
AOI21_X1 #() 
AOI21_X1_2161_ (
  .A({ S25957[1170] }),
  .B1({ S23352 }),
  .B2({ S23322 }),
  .ZN({ S23353 })
);
AND3_X1 #() 
AND3_X1_157_ (
  .A1({ S23352 }),
  .A2({ S23322 }),
  .A3({ S25957[1170] }),
  .ZN({ S23354 })
);
NOR2_X1 #() 
NOR2_X1_1021_ (
  .A1({ S23354 }),
  .A2({ S23353 }),
  .ZN({ S25957[914] })
);
NAND3_X1 #() 
NAND3_X1_4330_ (
  .A1({ S21907 }),
  .A2({ S21908 }),
  .A3({ S25956[0] }),
  .ZN({ S23355 })
);
NAND3_X1 #() 
NAND3_X1_4331_ (
  .A1({ S21902 }),
  .A2({ S21905 }),
  .A3({ S11550 }),
  .ZN({ S23356 })
);
NAND3_X1 #() 
NAND3_X1_4332_ (
  .A1({ S21979 }),
  .A2({ S21980 }),
  .A3({ S25956[1] }),
  .ZN({ S23357 })
);
NAND3_X1 #() 
NAND3_X1_4333_ (
  .A1({ S21974 }),
  .A2({ S21977 }),
  .A3({ S11539 }),
  .ZN({ S23358 })
);
NAND4_X1 #() 
NAND4_X1_471_ (
  .A1({ S23355 }),
  .A2({ S23356 }),
  .A3({ S23357 }),
  .A4({ S23358 }),
  .ZN({ S23359 })
);
INV_X1 #() 
INV_X1_1325_ (
  .A({ S23359 }),
  .ZN({ S87 })
);
NAND2_X1 #() 
NAND2_X1_4018_ (
  .A1({ S23355 }),
  .A2({ S23356 }),
  .ZN({ S23360 })
);
NAND2_X1 #() 
NAND2_X1_4019_ (
  .A1({ S23357 }),
  .A2({ S23358 }),
  .ZN({ S23361 })
);
NAND2_X1 #() 
NAND2_X1_4020_ (
  .A1({ S23360 }),
  .A2({ S23361 }),
  .ZN({ S88 })
);
XNOR2_X1 #() 
XNOR2_X1_170_ (
  .A({ S25957[1135] }),
  .B({ S11581 }),
  .ZN({ S25957[1071] })
);
AOI21_X1 #() 
AOI21_X1_2162_ (
  .A({ S25956[37] }),
  .B1({ S21646 }),
  .B2({ S21647 }),
  .ZN({ S23362 })
);
AND3_X1 #() 
AND3_X1_158_ (
  .A1({ S21646 }),
  .A2({ S25956[37] }),
  .A3({ S21647 }),
  .ZN({ S23363 })
);
OAI21_X1 #() 
OAI21_X1_2076_ (
  .A({ S20784 }),
  .B1({ S23363 }),
  .B2({ S23362 }),
  .ZN({ S23364 })
);
INV_X1 #() 
INV_X1_1326_ (
  .A({ S23362 }),
  .ZN({ S23365 })
);
NAND2_X1 #() 
NAND2_X1_4021_ (
  .A1({ S25957[1125] }),
  .A2({ S25956[37] }),
  .ZN({ S23366 })
);
NAND3_X1 #() 
NAND3_X1_4334_ (
  .A1({ S23365 }),
  .A2({ S25957[1157] }),
  .A3({ S23366 }),
  .ZN({ S23367 })
);
NAND2_X1 #() 
NAND2_X1_4022_ (
  .A1({ S23367 }),
  .A2({ S23364 }),
  .ZN({ S23368 })
);
NAND3_X1 #() 
NAND3_X1_4335_ (
  .A1({ S25957[1026] }),
  .A2({ S23355 }),
  .A3({ S23356 }),
  .ZN({ S23369 })
);
NAND2_X1 #() 
NAND2_X1_4023_ (
  .A1({ S25957[1026] }),
  .A2({ S23361 }),
  .ZN({ S23370 })
);
NAND2_X1 #() 
NAND2_X1_4024_ (
  .A1({ S23370 }),
  .A2({ S23359 }),
  .ZN({ S23371 })
);
NAND2_X1 #() 
NAND2_X1_4025_ (
  .A1({ S23371 }),
  .A2({ S23369 }),
  .ZN({ S23372 })
);
AOI21_X1 #() 
AOI21_X1_2163_ (
  .A({ S25957[1024] }),
  .B1({ S23361 }),
  .B2({ S25957[1026] }),
  .ZN({ S23373 })
);
OAI21_X1 #() 
OAI21_X1_2077_ (
  .A({ S25957[1028] }),
  .B1({ S23373 }),
  .B2({ S25957[1027] }),
  .ZN({ S23374 })
);
AOI21_X1 #() 
AOI21_X1_2164_ (
  .A({ S23374 }),
  .B1({ S23372 }),
  .B2({ S25957[1027] }),
  .ZN({ S23375 })
);
NAND2_X1 #() 
NAND2_X1_4026_ (
  .A1({ S23359 }),
  .A2({ S25957[1026] }),
  .ZN({ S23376 })
);
NAND2_X1 #() 
NAND2_X1_4027_ (
  .A1({ S23376 }),
  .A2({ S80 }),
  .ZN({ S23377 })
);
NAND3_X1 #() 
NAND3_X1_4336_ (
  .A1({ S22027 }),
  .A2({ S22030 }),
  .A3({ S25956[2] }),
  .ZN({ S23378 })
);
NAND3_X1 #() 
NAND3_X1_4337_ (
  .A1({ S22032 }),
  .A2({ S22033 }),
  .A3({ S11642 }),
  .ZN({ S23379 })
);
NAND4_X1 #() 
NAND4_X1_472_ (
  .A1({ S23378 }),
  .A2({ S23379 }),
  .A3({ S23357 }),
  .A4({ S23358 }),
  .ZN({ S23380 })
);
NAND2_X1 #() 
NAND2_X1_4028_ (
  .A1({ S23378 }),
  .A2({ S23379 }),
  .ZN({ S23381 })
);
NAND4_X1 #() 
NAND4_X1_473_ (
  .A1({ S23381 }),
  .A2({ S23361 }),
  .A3({ S23356 }),
  .A4({ S23355 }),
  .ZN({ S23382 })
);
AOI21_X1 #() 
AOI21_X1_2165_ (
  .A({ S80 }),
  .B1({ S23382 }),
  .B2({ S23380 }),
  .ZN({ S23383 })
);
NOR2_X1 #() 
NOR2_X1_1022_ (
  .A1({ S23383 }),
  .A2({ S25957[1028] }),
  .ZN({ S23384 })
);
AOI211_X1 #() 
AOI211_X1_67_ (
  .A({ S23368 }),
  .B({ S23375 }),
  .C1({ S23377 }),
  .C2({ S23384 }),
  .ZN({ S23385 })
);
NAND2_X1 #() 
NAND2_X1_4029_ (
  .A1({ S23381 }),
  .A2({ S23361 }),
  .ZN({ S23386 })
);
NAND2_X1 #() 
NAND2_X1_4030_ (
  .A1({ S23360 }),
  .A2({ S25957[1026] }),
  .ZN({ S23387 })
);
NAND2_X1 #() 
NAND2_X1_4031_ (
  .A1({ S23387 }),
  .A2({ S23386 }),
  .ZN({ S23388 })
);
NAND2_X1 #() 
NAND2_X1_4032_ (
  .A1({ S23388 }),
  .A2({ S25957[1027] }),
  .ZN({ S23389 })
);
NAND3_X1 #() 
NAND3_X1_4338_ (
  .A1({ S25957[1024] }),
  .A2({ S25957[1025] }),
  .A3({ S25957[1026] }),
  .ZN({ S23390 })
);
AOI22_X1 #() 
AOI22_X1_462_ (
  .A1({ S23378 }),
  .A2({ S23379 }),
  .B1({ S23358 }),
  .B2({ S23357 }),
  .ZN({ S23391 })
);
AOI21_X1 #() 
AOI21_X1_2166_ (
  .A({ S25957[1027] }),
  .B1({ S23391 }),
  .B2({ S25957[1024] }),
  .ZN({ S23392 })
);
AOI21_X1 #() 
AOI21_X1_2167_ (
  .A({ S25957[1028] }),
  .B1({ S23392 }),
  .B2({ S23390 }),
  .ZN({ S23393 })
);
NAND3_X1 #() 
NAND3_X1_4339_ (
  .A1({ S21744 }),
  .A2({ S21745 }),
  .A3({ S20774 }),
  .ZN({ S23394 })
);
NAND3_X1 #() 
NAND3_X1_4340_ (
  .A1({ S21739 }),
  .A2({ S21742 }),
  .A3({ S25957[1156] }),
  .ZN({ S23395 })
);
NAND2_X1 #() 
NAND2_X1_4033_ (
  .A1({ S23394 }),
  .A2({ S23395 }),
  .ZN({ S23396 })
);
OAI211_X1 #() 
OAI211_X1_1408_ (
  .A({ S23355 }),
  .B({ S23356 }),
  .C1({ S21981 }),
  .C2({ S21978 }),
  .ZN({ S23397 })
);
OAI211_X1 #() 
OAI211_X1_1409_ (
  .A({ S23357 }),
  .B({ S23358 }),
  .C1({ S21909 }),
  .C2({ S21906 }),
  .ZN({ S23398 })
);
NAND3_X1 #() 
NAND3_X1_4341_ (
  .A1({ S23398 }),
  .A2({ S23381 }),
  .A3({ S23397 }),
  .ZN({ S23399 })
);
AOI21_X1 #() 
AOI21_X1_2168_ (
  .A({ S80 }),
  .B1({ S23399 }),
  .B2({ S23376 }),
  .ZN({ S23400 })
);
NAND2_X1 #() 
NAND2_X1_4034_ (
  .A1({ S23360 }),
  .A2({ S23381 }),
  .ZN({ S23401 })
);
NAND3_X1 #() 
NAND3_X1_4342_ (
  .A1({ S23398 }),
  .A2({ S25957[1026] }),
  .A3({ S23397 }),
  .ZN({ S23402 })
);
NAND2_X1 #() 
NAND2_X1_4035_ (
  .A1({ S23402 }),
  .A2({ S23401 }),
  .ZN({ S23403 })
);
AOI211_X1 #() 
AOI211_X1_68_ (
  .A({ S23396 }),
  .B({ S23400 }),
  .C1({ S80 }),
  .C2({ S23403 }),
  .ZN({ S23404 })
);
AOI21_X1 #() 
AOI21_X1_2169_ (
  .A({ S23404 }),
  .B1({ S23393 }),
  .B2({ S23389 }),
  .ZN({ S23405 })
);
NOR2_X1 #() 
NOR2_X1_1023_ (
  .A1({ S23405 }),
  .A2({ S25957[1029] }),
  .ZN({ S23406 })
);
OAI21_X1 #() 
OAI21_X1_2078_ (
  .A({ S25957[1030] }),
  .B1({ S23406 }),
  .B2({ S23385 }),
  .ZN({ S23407 })
);
NOR2_X1 #() 
NOR2_X1_1024_ (
  .A1({ S25957[1024] }),
  .A2({ S23380 }),
  .ZN({ S23408 })
);
NAND3_X1 #() 
NAND3_X1_4343_ (
  .A1({ S25957[1024] }),
  .A2({ S25957[1025] }),
  .A3({ S23381 }),
  .ZN({ S23409 })
);
NAND3_X1 #() 
NAND3_X1_4344_ (
  .A1({ S88 }),
  .A2({ S25957[1026] }),
  .A3({ S23359 }),
  .ZN({ S23410 })
);
NAND3_X1 #() 
NAND3_X1_4345_ (
  .A1({ S23410 }),
  .A2({ S80 }),
  .A3({ S23409 }),
  .ZN({ S23411 })
);
OAI211_X1 #() 
OAI211_X1_1410_ (
  .A({ S23411 }),
  .B({ S25957[1028] }),
  .C1({ S80 }),
  .C2({ S23408 }),
  .ZN({ S23412 })
);
XNOR2_X1 #() 
XNOR2_X1_171_ (
  .A({ S23360 }),
  .B({ S23361 }),
  .ZN({ S23413 })
);
NAND3_X1 #() 
NAND3_X1_4346_ (
  .A1({ S23413 }),
  .A2({ S80 }),
  .A3({ S25957[1026] }),
  .ZN({ S23414 })
);
NOR2_X1 #() 
NOR2_X1_1025_ (
  .A1({ S80 }),
  .A2({ S23381 }),
  .ZN({ S23415 })
);
NAND2_X1 #() 
NAND2_X1_4036_ (
  .A1({ S23415 }),
  .A2({ S23359 }),
  .ZN({ S23416 })
);
NAND3_X1 #() 
NAND3_X1_4347_ (
  .A1({ S23414 }),
  .A2({ S23396 }),
  .A3({ S23416 }),
  .ZN({ S23417 })
);
AND2_X1 #() 
AND2_X1_254_ (
  .A1({ S23417 }),
  .A2({ S23368 }),
  .ZN({ S23418 })
);
NAND2_X1 #() 
NAND2_X1_4037_ (
  .A1({ S23359 }),
  .A2({ S23381 }),
  .ZN({ S23419 })
);
INV_X1 #() 
INV_X1_1327_ (
  .A({ S23419 }),
  .ZN({ S23420 })
);
NAND2_X1 #() 
NAND2_X1_4038_ (
  .A1({ S23380 }),
  .A2({ S80 }),
  .ZN({ S23421 })
);
NAND4_X1 #() 
NAND4_X1_474_ (
  .A1({ S22031 }),
  .A2({ S22034 }),
  .A3({ S23357 }),
  .A4({ S23358 }),
  .ZN({ S23422 })
);
NAND3_X1 #() 
NAND3_X1_4348_ (
  .A1({ S23397 }),
  .A2({ S25957[1027] }),
  .A3({ S23422 }),
  .ZN({ S23423 })
);
OAI21_X1 #() 
OAI21_X1_2079_ (
  .A({ S23423 }),
  .B1({ S23420 }),
  .B2({ S23421 }),
  .ZN({ S23424 })
);
AOI21_X1 #() 
AOI21_X1_2170_ (
  .A({ S80 }),
  .B1({ S23381 }),
  .B2({ S23361 }),
  .ZN({ S23425 })
);
NAND2_X1 #() 
NAND2_X1_4039_ (
  .A1({ S23425 }),
  .A2({ S23369 }),
  .ZN({ S23426 })
);
NAND3_X1 #() 
NAND3_X1_4349_ (
  .A1({ S80 }),
  .A2({ S23355 }),
  .A3({ S23356 }),
  .ZN({ S23427 })
);
INV_X1 #() 
INV_X1_1328_ (
  .A({ S23427 }),
  .ZN({ S23428 })
);
NOR2_X1 #() 
NOR2_X1_1026_ (
  .A1({ S23428 }),
  .A2({ S23396 }),
  .ZN({ S23429 })
);
AOI22_X1 #() 
AOI22_X1_463_ (
  .A1({ S23424 }),
  .A2({ S23396 }),
  .B1({ S23426 }),
  .B2({ S23429 }),
  .ZN({ S23430 })
);
AOI22_X1 #() 
AOI22_X1_464_ (
  .A1({ S23418 }),
  .A2({ S23412 }),
  .B1({ S25957[1029] }),
  .B2({ S23430 }),
  .ZN({ S23431 })
);
OAI211_X1 #() 
OAI211_X1_1411_ (
  .A({ S23407 }),
  .B({ S21512 }),
  .C1({ S25957[1030] }),
  .C2({ S23431 }),
  .ZN({ S23432 })
);
NAND3_X1 #() 
NAND3_X1_4350_ (
  .A1({ S23397 }),
  .A2({ S25957[1027] }),
  .A3({ S23381 }),
  .ZN({ S23433 })
);
AND2_X1 #() 
AND2_X1_255_ (
  .A1({ S23433 }),
  .A2({ S25957[1028] }),
  .ZN({ S23434 })
);
NAND2_X1 #() 
NAND2_X1_4040_ (
  .A1({ S23359 }),
  .A2({ S23380 }),
  .ZN({ S23435 })
);
INV_X1 #() 
INV_X1_1329_ (
  .A({ S23435 }),
  .ZN({ S23436 })
);
NAND2_X1 #() 
NAND2_X1_4041_ (
  .A1({ S23415 }),
  .A2({ S25957[1024] }),
  .ZN({ S23437 })
);
OAI211_X1 #() 
OAI211_X1_1412_ (
  .A({ S23434 }),
  .B({ S23437 }),
  .C1({ S23436 }),
  .C2({ S25957[1027] }),
  .ZN({ S23438 })
);
OAI21_X1 #() 
OAI21_X1_2080_ (
  .A({ S23397 }),
  .B1({ S25957[1024] }),
  .B2({ S23380 }),
  .ZN({ S23439 })
);
NAND2_X1 #() 
NAND2_X1_4042_ (
  .A1({ S23439 }),
  .A2({ S25957[1027] }),
  .ZN({ S23440 })
);
OAI21_X1 #() 
OAI21_X1_2081_ (
  .A({ S23440 }),
  .B1({ S23372 }),
  .B2({ S25957[1027] }),
  .ZN({ S23441 })
);
OAI211_X1 #() 
OAI211_X1_1413_ (
  .A({ S23438 }),
  .B({ S25957[1029] }),
  .C1({ S25957[1028] }),
  .C2({ S23441 }),
  .ZN({ S23442 })
);
NOR2_X1 #() 
NOR2_X1_1027_ (
  .A1({ S23371 }),
  .A2({ S80 }),
  .ZN({ S23443 })
);
AOI21_X1 #() 
AOI21_X1_2171_ (
  .A({ S25957[1027] }),
  .B1({ S23360 }),
  .B2({ S25957[1025] }),
  .ZN({ S23444 })
);
NOR2_X1 #() 
NOR2_X1_1028_ (
  .A1({ S23443 }),
  .A2({ S23444 }),
  .ZN({ S23445 })
);
NOR2_X1 #() 
NOR2_X1_1029_ (
  .A1({ S23445 }),
  .A2({ S23396 }),
  .ZN({ S23446 })
);
NAND4_X1 #() 
NAND4_X1_475_ (
  .A1({ S23355 }),
  .A2({ S23356 }),
  .A3({ S22031 }),
  .A4({ S22034 }),
  .ZN({ S23447 })
);
NOR2_X1 #() 
NOR2_X1_1030_ (
  .A1({ S23391 }),
  .A2({ S25957[1024] }),
  .ZN({ S23448 })
);
NAND2_X1 #() 
NAND2_X1_4043_ (
  .A1({ S23448 }),
  .A2({ S23380 }),
  .ZN({ S23449 })
);
OAI21_X1 #() 
OAI21_X1_2082_ (
  .A({ S23396 }),
  .B1({ S80 }),
  .B2({ S23397 }),
  .ZN({ S23450 })
);
AOI21_X1 #() 
AOI21_X1_2172_ (
  .A({ S23450 }),
  .B1({ S23449 }),
  .B2({ S23447 }),
  .ZN({ S23451 })
);
OAI21_X1 #() 
OAI21_X1_2083_ (
  .A({ S23368 }),
  .B1({ S23446 }),
  .B2({ S23451 }),
  .ZN({ S23452 })
);
NAND3_X1 #() 
NAND3_X1_4351_ (
  .A1({ S23452 }),
  .A2({ S23442 }),
  .A3({ S25957[1030] }),
  .ZN({ S23453 })
);
NAND3_X1 #() 
NAND3_X1_4352_ (
  .A1({ S88 }),
  .A2({ S23381 }),
  .A3({ S23359 }),
  .ZN({ S23454 })
);
NAND2_X1 #() 
NAND2_X1_4044_ (
  .A1({ S23397 }),
  .A2({ S25957[1026] }),
  .ZN({ S23455 })
);
AOI21_X1 #() 
AOI21_X1_2173_ (
  .A({ S25957[1027] }),
  .B1({ S23454 }),
  .B2({ S23455 }),
  .ZN({ S23456 })
);
NOR3_X1 #() 
NOR3_X1_138_ (
  .A1({ S23456 }),
  .A2({ S23425 }),
  .A3({ S25957[1028] }),
  .ZN({ S23457 })
);
INV_X1 #() 
INV_X1_1330_ (
  .A({ S23380 }),
  .ZN({ S23458 })
);
NAND3_X1 #() 
NAND3_X1_4353_ (
  .A1({ S23402 }),
  .A2({ S23454 }),
  .A3({ S25957[1027] }),
  .ZN({ S23459 })
);
NAND2_X1 #() 
NAND2_X1_4045_ (
  .A1({ S23447 }),
  .A2({ S80 }),
  .ZN({ S23460 })
);
OAI21_X1 #() 
OAI21_X1_2084_ (
  .A({ S23459 }),
  .B1({ S23458 }),
  .B2({ S23460 }),
  .ZN({ S23461 })
);
OAI21_X1 #() 
OAI21_X1_2085_ (
  .A({ S23368 }),
  .B1({ S23461 }),
  .B2({ S23396 }),
  .ZN({ S23462 })
);
NOR2_X1 #() 
NOR2_X1_1031_ (
  .A1({ S23360 }),
  .A2({ S23381 }),
  .ZN({ S23463 })
);
NAND2_X1 #() 
NAND2_X1_4046_ (
  .A1({ S25957[1025] }),
  .A2({ S80 }),
  .ZN({ S23464 })
);
OAI21_X1 #() 
OAI21_X1_2086_ (
  .A({ S25957[1027] }),
  .B1({ S23463 }),
  .B2({ S23361 }),
  .ZN({ S23465 })
);
OAI211_X1 #() 
OAI211_X1_1414_ (
  .A({ S23465 }),
  .B({ S25957[1028] }),
  .C1({ S23463 }),
  .C2({ S23464 }),
  .ZN({ S23466 })
);
NAND3_X1 #() 
NAND3_X1_4354_ (
  .A1({ S23360 }),
  .A2({ S23381 }),
  .A3({ S23361 }),
  .ZN({ S23467 })
);
NAND2_X1 #() 
NAND2_X1_4047_ (
  .A1({ S23467 }),
  .A2({ S80 }),
  .ZN({ S23468 })
);
NAND3_X1 #() 
NAND3_X1_4355_ (
  .A1({ S23468 }),
  .A2({ S23396 }),
  .A3({ S23359 }),
  .ZN({ S23469 })
);
NAND3_X1 #() 
NAND3_X1_4356_ (
  .A1({ S23466 }),
  .A2({ S25957[1029] }),
  .A3({ S23469 }),
  .ZN({ S23470 })
);
OAI211_X1 #() 
OAI211_X1_1415_ (
  .A({ S21581 }),
  .B({ S23470 }),
  .C1({ S23462 }),
  .C2({ S23457 }),
  .ZN({ S23471 })
);
NAND3_X1 #() 
NAND3_X1_4357_ (
  .A1({ S23453 }),
  .A2({ S23471 }),
  .A3({ S25957[1031] }),
  .ZN({ S23472 })
);
NAND2_X1 #() 
NAND2_X1_4048_ (
  .A1({ S23432 }),
  .A2({ S23472 }),
  .ZN({ S23473 })
);
NOR2_X1 #() 
NOR2_X1_1032_ (
  .A1({ S23473 }),
  .A2({ S12802 }),
  .ZN({ S23474 })
);
NAND2_X1 #() 
NAND2_X1_4049_ (
  .A1({ S23473 }),
  .A2({ S12802 }),
  .ZN({ S23475 })
);
INV_X1 #() 
INV_X1_1331_ (
  .A({ S23475 }),
  .ZN({ S23476 })
);
OAI21_X1 #() 
OAI21_X1_2087_ (
  .A({ S25957[1071] }),
  .B1({ S23476 }),
  .B2({ S23474 }),
  .ZN({ S23477 })
);
INV_X1 #() 
INV_X1_1332_ (
  .A({ S25957[1071] }),
  .ZN({ S23478 })
);
NOR2_X1 #() 
NOR2_X1_1033_ (
  .A1({ S23476 }),
  .A2({ S23474 }),
  .ZN({ S25957[975] })
);
NAND2_X1 #() 
NAND2_X1_4050_ (
  .A1({ S25957[975] }),
  .A2({ S23478 }),
  .ZN({ S23479 })
);
NAND3_X1 #() 
NAND3_X1_4358_ (
  .A1({ S23479 }),
  .A2({ S25957[1039] }),
  .A3({ S23477 }),
  .ZN({ S23480 })
);
NAND2_X1 #() 
NAND2_X1_4051_ (
  .A1({ S23479 }),
  .A2({ S23477 }),
  .ZN({ S25957[943] })
);
NAND2_X1 #() 
NAND2_X1_4052_ (
  .A1({ S25957[943] }),
  .A2({ S22726 }),
  .ZN({ S23481 })
);
NAND2_X1 #() 
NAND2_X1_4053_ (
  .A1({ S23481 }),
  .A2({ S23480 }),
  .ZN({ S25957[911] })
);
XOR2_X1 #() 
XOR2_X1_73_ (
  .A({ S25957[1102] }),
  .B({ S25957[1198] }),
  .Z({ S25957[1070] })
);
NAND3_X1 #() 
NAND3_X1_4359_ (
  .A1({ S23387 }),
  .A2({ S23380 }),
  .A3({ S23447 }),
  .ZN({ S23482 })
);
AOI21_X1 #() 
AOI21_X1_2174_ (
  .A({ S23396 }),
  .B1({ S23482 }),
  .B2({ S25957[1027] }),
  .ZN({ S23483 })
);
INV_X1 #() 
INV_X1_1333_ (
  .A({ S23483 }),
  .ZN({ S23484 })
);
AOI21_X1 #() 
AOI21_X1_2175_ (
  .A({ S25957[1027] }),
  .B1({ S23454 }),
  .B2({ S23369 }),
  .ZN({ S23485 })
);
OAI211_X1 #() 
OAI211_X1_1416_ (
  .A({ S23393 }),
  .B({ S23437 }),
  .C1({ S23436 }),
  .C2({ S80 }),
  .ZN({ S23486 })
);
OAI211_X1 #() 
OAI211_X1_1417_ (
  .A({ S23486 }),
  .B({ S23368 }),
  .C1({ S23484 }),
  .C2({ S23485 }),
  .ZN({ S23487 })
);
AOI21_X1 #() 
AOI21_X1_2176_ (
  .A({ S80 }),
  .B1({ S23455 }),
  .B2({ S23447 }),
  .ZN({ S23488 })
);
NAND2_X1 #() 
NAND2_X1_4054_ (
  .A1({ S23396 }),
  .A2({ S23464 }),
  .ZN({ S23489 })
);
INV_X1 #() 
INV_X1_1334_ (
  .A({ S23422 }),
  .ZN({ S23490 })
);
AOI21_X1 #() 
AOI21_X1_2177_ (
  .A({ S23396 }),
  .B1({ S25957[1027] }),
  .B2({ S23490 }),
  .ZN({ S23491 })
);
AOI22_X1 #() 
AOI22_X1_465_ (
  .A1({ S23356 }),
  .A2({ S23355 }),
  .B1({ S23357 }),
  .B2({ S23358 }),
  .ZN({ S23492 })
);
OAI21_X1 #() 
OAI21_X1_2088_ (
  .A({ S80 }),
  .B1({ S23492 }),
  .B2({ S23381 }),
  .ZN({ S23493 })
);
NAND2_X1 #() 
NAND2_X1_4055_ (
  .A1({ S23491 }),
  .A2({ S23493 }),
  .ZN({ S23494 })
);
OAI221_X1 #() 
OAI221_X1_117_ (
  .A({ S25957[1029] }),
  .B1({ S23489 }),
  .B2({ S23443 }),
  .C1({ S23494 }),
  .C2({ S23488 }),
  .ZN({ S23495 })
);
NAND3_X1 #() 
NAND3_X1_4360_ (
  .A1({ S23487 }),
  .A2({ S25957[1030] }),
  .A3({ S23495 }),
  .ZN({ S23496 })
);
NAND2_X1 #() 
NAND2_X1_4056_ (
  .A1({ S23458 }),
  .A2({ S25957[1027] }),
  .ZN({ S23497 })
);
AOI21_X1 #() 
AOI21_X1_2178_ (
  .A({ S25957[1026] }),
  .B1({ S23356 }),
  .B2({ S23355 }),
  .ZN({ S23498 })
);
NOR2_X1 #() 
NOR2_X1_1034_ (
  .A1({ S25957[1027] }),
  .A2({ S23361 }),
  .ZN({ S23499 })
);
NAND2_X1 #() 
NAND2_X1_4057_ (
  .A1({ S23499 }),
  .A2({ S23498 }),
  .ZN({ S23500 })
);
NAND4_X1 #() 
NAND4_X1_476_ (
  .A1({ S23414 }),
  .A2({ S25957[1028] }),
  .A3({ S23497 }),
  .A4({ S23500 }),
  .ZN({ S23501 })
);
INV_X1 #() 
INV_X1_1335_ (
  .A({ S23425 }),
  .ZN({ S23502 })
);
NAND3_X1 #() 
NAND3_X1_4361_ (
  .A1({ S23398 }),
  .A2({ S23397 }),
  .A3({ S23422 }),
  .ZN({ S23503 })
);
NAND2_X1 #() 
NAND2_X1_4058_ (
  .A1({ S23503 }),
  .A2({ S80 }),
  .ZN({ S23504 })
);
OAI211_X1 #() 
OAI211_X1_1418_ (
  .A({ S23504 }),
  .B({ S23396 }),
  .C1({ S23435 }),
  .C2({ S23502 }),
  .ZN({ S23505 })
);
NAND3_X1 #() 
NAND3_X1_4362_ (
  .A1({ S23501 }),
  .A2({ S25957[1029] }),
  .A3({ S23505 }),
  .ZN({ S23506 })
);
NAND2_X1 #() 
NAND2_X1_4059_ (
  .A1({ S23397 }),
  .A2({ S23381 }),
  .ZN({ S23507 })
);
OAI21_X1 #() 
OAI21_X1_2089_ (
  .A({ S23465 }),
  .B1({ S25957[1027] }),
  .B2({ S23507 }),
  .ZN({ S23508 })
);
NAND3_X1 #() 
NAND3_X1_4363_ (
  .A1({ S25957[1025] }),
  .A2({ S23360 }),
  .A3({ S25957[1026] }),
  .ZN({ S23509 })
);
AOI21_X1 #() 
AOI21_X1_2179_ (
  .A({ S80 }),
  .B1({ S23509 }),
  .B2({ S23447 }),
  .ZN({ S23510 })
);
OAI21_X1 #() 
OAI21_X1_2090_ (
  .A({ S23396 }),
  .B1({ S23485 }),
  .B2({ S23510 }),
  .ZN({ S23511 })
);
OAI21_X1 #() 
OAI21_X1_2091_ (
  .A({ S23511 }),
  .B1({ S23396 }),
  .B2({ S23508 }),
  .ZN({ S23512 })
);
NAND2_X1 #() 
NAND2_X1_4060_ (
  .A1({ S23512 }),
  .A2({ S23368 }),
  .ZN({ S23513 })
);
NAND3_X1 #() 
NAND3_X1_4364_ (
  .A1({ S23513 }),
  .A2({ S21581 }),
  .A3({ S23506 }),
  .ZN({ S23514 })
);
NAND3_X1 #() 
NAND3_X1_4365_ (
  .A1({ S23514 }),
  .A2({ S25957[1031] }),
  .A3({ S23496 }),
  .ZN({ S23515 })
);
NAND2_X1 #() 
NAND2_X1_4061_ (
  .A1({ S88 }),
  .A2({ S23447 }),
  .ZN({ S23516 })
);
NAND3_X1 #() 
NAND3_X1_4366_ (
  .A1({ S23376 }),
  .A2({ S80 }),
  .A3({ S23447 }),
  .ZN({ S23517 })
);
OAI21_X1 #() 
OAI21_X1_2092_ (
  .A({ S23517 }),
  .B1({ S80 }),
  .B2({ S23516 }),
  .ZN({ S23518 })
);
NOR2_X1 #() 
NOR2_X1_1035_ (
  .A1({ S23518 }),
  .A2({ S23396 }),
  .ZN({ S23519 })
);
NAND2_X1 #() 
NAND2_X1_4062_ (
  .A1({ S23447 }),
  .A2({ S25957[1025] }),
  .ZN({ S23520 })
);
AOI21_X1 #() 
AOI21_X1_2180_ (
  .A({ S25957[1028] }),
  .B1({ S23437 }),
  .B2({ S23520 }),
  .ZN({ S23521 })
);
OAI21_X1 #() 
OAI21_X1_2093_ (
  .A({ S25957[1029] }),
  .B1({ S23519 }),
  .B2({ S23521 }),
  .ZN({ S23522 })
);
NAND2_X1 #() 
NAND2_X1_4063_ (
  .A1({ S23410 }),
  .A2({ S80 }),
  .ZN({ S23523 })
);
NOR2_X1 #() 
NOR2_X1_1036_ (
  .A1({ S23488 }),
  .A2({ S25957[1028] }),
  .ZN({ S23524 })
);
NAND2_X1 #() 
NAND2_X1_4064_ (
  .A1({ S23524 }),
  .A2({ S23523 }),
  .ZN({ S23525 })
);
INV_X1 #() 
INV_X1_1336_ (
  .A({ S23448 }),
  .ZN({ S23526 })
);
OAI21_X1 #() 
OAI21_X1_2094_ (
  .A({ S23491 }),
  .B1({ S23526 }),
  .B2({ S25957[1027] }),
  .ZN({ S23527 })
);
NAND3_X1 #() 
NAND3_X1_4367_ (
  .A1({ S23525 }),
  .A2({ S23368 }),
  .A3({ S23527 }),
  .ZN({ S23528 })
);
AOI21_X1 #() 
AOI21_X1_2181_ (
  .A({ S21581 }),
  .B1({ S23522 }),
  .B2({ S23528 }),
  .ZN({ S23529 })
);
NAND2_X1 #() 
NAND2_X1_4065_ (
  .A1({ S23460 }),
  .A2({ S25957[1028] }),
  .ZN({ S23530 })
);
NAND3_X1 #() 
NAND3_X1_4368_ (
  .A1({ S23360 }),
  .A2({ S25957[1026] }),
  .A3({ S23361 }),
  .ZN({ S23531 })
);
NAND2_X1 #() 
NAND2_X1_4066_ (
  .A1({ S23531 }),
  .A2({ S25957[1027] }),
  .ZN({ S23532 })
);
NOR2_X1 #() 
NOR2_X1_1037_ (
  .A1({ S23532 }),
  .A2({ S87 }),
  .ZN({ S23533 })
);
NAND2_X1 #() 
NAND2_X1_4067_ (
  .A1({ S23370 }),
  .A2({ S25957[1027] }),
  .ZN({ S23534 })
);
NAND2_X1 #() 
NAND2_X1_4068_ (
  .A1({ S23392 }),
  .A2({ S23380 }),
  .ZN({ S23535 })
);
OAI21_X1 #() 
OAI21_X1_2095_ (
  .A({ S23535 }),
  .B1({ S23490 }),
  .B2({ S23534 }),
  .ZN({ S23536 })
);
OAI22_X1 #() 
OAI22_X1_106_ (
  .A1({ S23536 }),
  .A2({ S25957[1028] }),
  .B1({ S23530 }),
  .B2({ S23533 }),
  .ZN({ S23537 })
);
NOR3_X1 #() 
NOR3_X1_139_ (
  .A1({ S23383 }),
  .A2({ S23392 }),
  .A3({ S23396 }),
  .ZN({ S23538 })
);
NAND2_X1 #() 
NAND2_X1_4069_ (
  .A1({ S23386 }),
  .A2({ S23447 }),
  .ZN({ S23539 })
);
OAI21_X1 #() 
OAI21_X1_2096_ (
  .A({ S25957[1027] }),
  .B1({ S23408 }),
  .B2({ S23539 }),
  .ZN({ S23540 })
);
OAI21_X1 #() 
OAI21_X1_2097_ (
  .A({ S23368 }),
  .B1({ S23540 }),
  .B2({ S25957[1028] }),
  .ZN({ S23541 })
);
OAI21_X1 #() 
OAI21_X1_2098_ (
  .A({ S21581 }),
  .B1({ S23541 }),
  .B2({ S23538 }),
  .ZN({ S23542 })
);
AOI21_X1 #() 
AOI21_X1_2182_ (
  .A({ S23542 }),
  .B1({ S23537 }),
  .B2({ S25957[1029] }),
  .ZN({ S23543 })
);
OAI21_X1 #() 
OAI21_X1_2099_ (
  .A({ S21512 }),
  .B1({ S23529 }),
  .B2({ S23543 }),
  .ZN({ S23544 })
);
NAND2_X1 #() 
NAND2_X1_4070_ (
  .A1({ S23515 }),
  .A2({ S23544 }),
  .ZN({ S23545 })
);
NOR2_X1 #() 
NOR2_X1_1038_ (
  .A1({ S23545 }),
  .A2({ S20876 }),
  .ZN({ S23546 })
);
AOI21_X1 #() 
AOI21_X1_2183_ (
  .A({ S25957[1230] }),
  .B1({ S23515 }),
  .B2({ S23544 }),
  .ZN({ S23547 })
);
NOR2_X1 #() 
NOR2_X1_1039_ (
  .A1({ S23546 }),
  .A2({ S23547 }),
  .ZN({ S25957[974] })
);
INV_X1 #() 
INV_X1_1337_ (
  .A({ S25957[974] }),
  .ZN({ S23548 })
);
NAND2_X1 #() 
NAND2_X1_4071_ (
  .A1({ S23548 }),
  .A2({ S20130 }),
  .ZN({ S23549 })
);
NAND2_X1 #() 
NAND2_X1_4072_ (
  .A1({ S25957[974] }),
  .A2({ S25957[1166] }),
  .ZN({ S23550 })
);
NAND2_X1 #() 
NAND2_X1_4073_ (
  .A1({ S23549 }),
  .A2({ S23550 }),
  .ZN({ S23551 })
);
INV_X1 #() 
INV_X1_1338_ (
  .A({ S23551 }),
  .ZN({ S25957[910] })
);
NAND2_X1 #() 
NAND2_X1_4074_ (
  .A1({ S21010 }),
  .A2({ S21009 }),
  .ZN({ S25957[1069] })
);
INV_X1 #() 
INV_X1_1339_ (
  .A({ S25957[1069] }),
  .ZN({ S23552 })
);
NAND2_X1 #() 
NAND2_X1_4075_ (
  .A1({ S14362 }),
  .A2({ S14391 }),
  .ZN({ S25957[1229] })
);
NAND2_X1 #() 
NAND2_X1_4076_ (
  .A1({ S25957[1027] }),
  .A2({ S23361 }),
  .ZN({ S23553 })
);
AOI21_X1 #() 
AOI21_X1_2184_ (
  .A({ S25957[1027] }),
  .B1({ S23370 }),
  .B2({ S23359 }),
  .ZN({ S23554 })
);
INV_X1 #() 
INV_X1_1340_ (
  .A({ S23554 }),
  .ZN({ S23555 })
);
NAND3_X1 #() 
NAND3_X1_4369_ (
  .A1({ S23555 }),
  .A2({ S23396 }),
  .A3({ S23553 }),
  .ZN({ S23556 })
);
NAND2_X1 #() 
NAND2_X1_4077_ (
  .A1({ S25957[1027] }),
  .A2({ S25957[1026] }),
  .ZN({ S23557 })
);
NAND3_X1 #() 
NAND3_X1_4370_ (
  .A1({ S23557 }),
  .A2({ S23397 }),
  .A3({ S23387 }),
  .ZN({ S23558 })
);
AND2_X1 #() 
AND2_X1_256_ (
  .A1({ S23558 }),
  .A2({ S23416 }),
  .ZN({ S23559 })
);
OAI21_X1 #() 
OAI21_X1_2100_ (
  .A({ S23556 }),
  .B1({ S23559 }),
  .B2({ S23396 }),
  .ZN({ S23560 })
);
NAND2_X1 #() 
NAND2_X1_4078_ (
  .A1({ S23560 }),
  .A2({ S25957[1029] }),
  .ZN({ S23561 })
);
NAND2_X1 #() 
NAND2_X1_4079_ (
  .A1({ S23409 }),
  .A2({ S80 }),
  .ZN({ S23562 })
);
OAI211_X1 #() 
OAI211_X1_1419_ (
  .A({ S23402 }),
  .B({ S25957[1027] }),
  .C1({ S25957[1026] }),
  .C2({ S23492 }),
  .ZN({ S23563 })
);
AOI21_X1 #() 
AOI21_X1_2185_ (
  .A({ S25957[1028] }),
  .B1({ S23563 }),
  .B2({ S23562 }),
  .ZN({ S23564 })
);
INV_X1 #() 
INV_X1_1341_ (
  .A({ S23460 }),
  .ZN({ S23565 })
);
NOR2_X1 #() 
NOR2_X1_1040_ (
  .A1({ S23454 }),
  .A2({ S80 }),
  .ZN({ S23566 })
);
AOI21_X1 #() 
AOI21_X1_2186_ (
  .A({ S23566 }),
  .B1({ S23565 }),
  .B2({ S23361 }),
  .ZN({ S23567 })
);
NAND2_X1 #() 
NAND2_X1_4080_ (
  .A1({ S23567 }),
  .A2({ S25957[1028] }),
  .ZN({ S23568 })
);
NAND2_X1 #() 
NAND2_X1_4081_ (
  .A1({ S23568 }),
  .A2({ S23368 }),
  .ZN({ S23569 })
);
OAI21_X1 #() 
OAI21_X1_2101_ (
  .A({ S23561 }),
  .B1({ S23569 }),
  .B2({ S23564 }),
  .ZN({ S23570 })
);
NAND2_X1 #() 
NAND2_X1_4082_ (
  .A1({ S23570 }),
  .A2({ S21581 }),
  .ZN({ S23571 })
);
NOR2_X1 #() 
NOR2_X1_1041_ (
  .A1({ S23448 }),
  .A2({ S80 }),
  .ZN({ S23572 })
);
AOI21_X1 #() 
AOI21_X1_2187_ (
  .A({ S25957[1027] }),
  .B1({ S23507 }),
  .B2({ S23509 }),
  .ZN({ S23573 })
);
NOR3_X1 #() 
NOR3_X1_140_ (
  .A1({ S23573 }),
  .A2({ S23572 }),
  .A3({ S23396 }),
  .ZN({ S23574 })
);
AOI21_X1 #() 
AOI21_X1_2188_ (
  .A({ S25957[1028] }),
  .B1({ S23463 }),
  .B2({ S25957[1027] }),
  .ZN({ S23575 })
);
NAND3_X1 #() 
NAND3_X1_4371_ (
  .A1({ S88 }),
  .A2({ S23386 }),
  .A3({ S80 }),
  .ZN({ S23576 })
);
NAND3_X1 #() 
NAND3_X1_4372_ (
  .A1({ S23359 }),
  .A2({ S23380 }),
  .A3({ S25957[1027] }),
  .ZN({ S23577 })
);
AND3_X1 #() 
AND3_X1_159_ (
  .A1({ S23575 }),
  .A2({ S23576 }),
  .A3({ S23577 }),
  .ZN({ S23578 })
);
OR3_X1 #() 
OR3_X1_26_ (
  .A1({ S23574 }),
  .A2({ S23578 }),
  .A3({ S23368 }),
  .ZN({ S23579 })
);
AND2_X1 #() 
AND2_X1_257_ (
  .A1({ S23524 }),
  .A2({ S23414 }),
  .ZN({ S23580 })
);
NAND2_X1 #() 
NAND2_X1_4083_ (
  .A1({ S23369 }),
  .A2({ S23370 }),
  .ZN({ S23581 })
);
NAND3_X1 #() 
NAND3_X1_4373_ (
  .A1({ S23386 }),
  .A2({ S25957[1027] }),
  .A3({ S23447 }),
  .ZN({ S23582 })
);
NAND2_X1 #() 
NAND2_X1_4084_ (
  .A1({ S23582 }),
  .A2({ S25957[1028] }),
  .ZN({ S23583 })
);
AOI21_X1 #() 
AOI21_X1_2189_ (
  .A({ S23583 }),
  .B1({ S23581 }),
  .B2({ S80 }),
  .ZN({ S23584 })
);
NOR2_X1 #() 
NOR2_X1_1042_ (
  .A1({ S23580 }),
  .A2({ S23584 }),
  .ZN({ S23585 })
);
NAND2_X1 #() 
NAND2_X1_4085_ (
  .A1({ S23585 }),
  .A2({ S23368 }),
  .ZN({ S23586 })
);
NAND3_X1 #() 
NAND3_X1_4374_ (
  .A1({ S23586 }),
  .A2({ S25957[1030] }),
  .A3({ S23579 }),
  .ZN({ S23587 })
);
NAND3_X1 #() 
NAND3_X1_4375_ (
  .A1({ S23571 }),
  .A2({ S23587 }),
  .A3({ S25957[1031] }),
  .ZN({ S23588 })
);
AOI21_X1 #() 
AOI21_X1_2190_ (
  .A({ S80 }),
  .B1({ S23355 }),
  .B2({ S23356 }),
  .ZN({ S23589 })
);
AOI21_X1 #() 
AOI21_X1_2191_ (
  .A({ S23589 }),
  .B1({ S23444 }),
  .B2({ S23447 }),
  .ZN({ S23590 })
);
NAND3_X1 #() 
NAND3_X1_4376_ (
  .A1({ S25957[1025] }),
  .A2({ S23360 }),
  .A3({ S23381 }),
  .ZN({ S23591 })
);
NAND3_X1 #() 
NAND3_X1_4377_ (
  .A1({ S23402 }),
  .A2({ S25957[1027] }),
  .A3({ S23591 }),
  .ZN({ S23592 })
);
NAND4_X1 #() 
NAND4_X1_477_ (
  .A1({ S23401 }),
  .A2({ S23370 }),
  .A3({ S80 }),
  .A4({ S23422 }),
  .ZN({ S23593 })
);
NAND3_X1 #() 
NAND3_X1_4378_ (
  .A1({ S23592 }),
  .A2({ S25957[1028] }),
  .A3({ S23593 }),
  .ZN({ S23594 })
);
OAI211_X1 #() 
OAI211_X1_1420_ (
  .A({ S23594 }),
  .B({ S25957[1029] }),
  .C1({ S25957[1028] }),
  .C2({ S23590 }),
  .ZN({ S23595 })
);
NAND4_X1 #() 
NAND4_X1_478_ (
  .A1({ S23398 }),
  .A2({ S23401 }),
  .A3({ S23397 }),
  .A4({ S80 }),
  .ZN({ S23596 })
);
NAND3_X1 #() 
NAND3_X1_4379_ (
  .A1({ S23402 }),
  .A2({ S25957[1027] }),
  .A3({ S23382 }),
  .ZN({ S23597 })
);
AOI21_X1 #() 
AOI21_X1_2192_ (
  .A({ S23396 }),
  .B1({ S23597 }),
  .B2({ S23596 }),
  .ZN({ S23598 })
);
NOR2_X1 #() 
NOR2_X1_1043_ (
  .A1({ S25957[1027] }),
  .A2({ S25957[1026] }),
  .ZN({ S23599 })
);
INV_X1 #() 
INV_X1_1342_ (
  .A({ S23599 }),
  .ZN({ S23600 })
);
NAND2_X1 #() 
NAND2_X1_4086_ (
  .A1({ S23600 }),
  .A2({ S23369 }),
  .ZN({ S23601 })
);
AOI21_X1 #() 
AOI21_X1_2193_ (
  .A({ S80 }),
  .B1({ S23359 }),
  .B2({ S23381 }),
  .ZN({ S23602 })
);
AOI211_X1 #() 
AOI211_X1_69_ (
  .A({ S23396 }),
  .B({ S23602 }),
  .C1({ S23498 }),
  .C2({ S23499 }),
  .ZN({ S23603 })
);
AOI21_X1 #() 
AOI21_X1_2194_ (
  .A({ S23603 }),
  .B1({ S23601 }),
  .B2({ S23521 }),
  .ZN({ S23604 })
);
NOR2_X1 #() 
NOR2_X1_1044_ (
  .A1({ S23464 }),
  .A2({ S23369 }),
  .ZN({ S23605 })
);
OAI21_X1 #() 
OAI21_X1_2102_ (
  .A({ S23368 }),
  .B1({ S23450 }),
  .B2({ S23605 }),
  .ZN({ S23606 })
);
OAI22_X1 #() 
OAI22_X1_107_ (
  .A1({ S23604 }),
  .A2({ S23368 }),
  .B1({ S23598 }),
  .B2({ S23606 }),
  .ZN({ S23607 })
);
NAND3_X1 #() 
NAND3_X1_4380_ (
  .A1({ S23376 }),
  .A2({ S25957[1027] }),
  .A3({ S23447 }),
  .ZN({ S23608 })
);
NAND3_X1 #() 
NAND3_X1_4381_ (
  .A1({ S23591 }),
  .A2({ S80 }),
  .A3({ S23369 }),
  .ZN({ S23609 })
);
NAND2_X1 #() 
NAND2_X1_4087_ (
  .A1({ S23608 }),
  .A2({ S23609 }),
  .ZN({ S23610 })
);
NAND3_X1 #() 
NAND3_X1_4382_ (
  .A1({ S23390 }),
  .A2({ S80 }),
  .A3({ S23419 }),
  .ZN({ S23611 })
);
AOI22_X1 #() 
AOI22_X1_466_ (
  .A1({ S23396 }),
  .A2({ S23610 }),
  .B1({ S23434 }),
  .B2({ S23611 }),
  .ZN({ S23612 })
);
AOI21_X1 #() 
AOI21_X1_2195_ (
  .A({ S21581 }),
  .B1({ S23612 }),
  .B2({ S23368 }),
  .ZN({ S23613 })
);
AOI22_X1 #() 
AOI22_X1_467_ (
  .A1({ S23607 }),
  .A2({ S21581 }),
  .B1({ S23595 }),
  .B2({ S23613 }),
  .ZN({ S23614 })
);
OAI211_X1 #() 
OAI211_X1_1421_ (
  .A({ S23588 }),
  .B({ S25957[1229] }),
  .C1({ S25957[1031] }),
  .C2({ S23614 }),
  .ZN({ S23615 })
);
INV_X1 #() 
INV_X1_1343_ (
  .A({ S25957[1229] }),
  .ZN({ S23616 })
);
OAI21_X1 #() 
OAI21_X1_2103_ (
  .A({ S25957[1029] }),
  .B1({ S23574 }),
  .B2({ S23578 }),
  .ZN({ S23617 })
);
OAI211_X1 #() 
OAI211_X1_1422_ (
  .A({ S25957[1030] }),
  .B({ S23617 }),
  .C1({ S23585 }),
  .C2({ S25957[1029] }),
  .ZN({ S23618 })
);
OAI211_X1 #() 
OAI211_X1_1423_ (
  .A({ S21581 }),
  .B({ S23561 }),
  .C1({ S23569 }),
  .C2({ S23564 }),
  .ZN({ S23619 })
);
AOI21_X1 #() 
AOI21_X1_2196_ (
  .A({ S21512 }),
  .B1({ S23618 }),
  .B2({ S23619 }),
  .ZN({ S23620 })
);
NOR2_X1 #() 
NOR2_X1_1045_ (
  .A1({ S23614 }),
  .A2({ S25957[1031] }),
  .ZN({ S23621 })
);
OAI21_X1 #() 
OAI21_X1_2104_ (
  .A({ S23616 }),
  .B1({ S23621 }),
  .B2({ S23620 }),
  .ZN({ S23622 })
);
NAND2_X1 #() 
NAND2_X1_4088_ (
  .A1({ S23622 }),
  .A2({ S23615 }),
  .ZN({ S23623 })
);
NAND2_X1 #() 
NAND2_X1_4089_ (
  .A1({ S23623 }),
  .A2({ S23552 }),
  .ZN({ S23624 })
);
NAND3_X1 #() 
NAND3_X1_4383_ (
  .A1({ S23622 }),
  .A2({ S23615 }),
  .A3({ S25957[1069] }),
  .ZN({ S23625 })
);
NAND3_X1 #() 
NAND3_X1_4384_ (
  .A1({ S23624 }),
  .A2({ S21015 }),
  .A3({ S23625 }),
  .ZN({ S23626 })
);
NAND2_X1 #() 
NAND2_X1_4090_ (
  .A1({ S23623 }),
  .A2({ S25957[1069] }),
  .ZN({ S23627 })
);
NAND3_X1 #() 
NAND3_X1_4385_ (
  .A1({ S23622 }),
  .A2({ S23615 }),
  .A3({ S23552 }),
  .ZN({ S23628 })
);
NAND3_X1 #() 
NAND3_X1_4386_ (
  .A1({ S23627 }),
  .A2({ S25957[1037] }),
  .A3({ S23628 }),
  .ZN({ S23629 })
);
NAND2_X1 #() 
NAND2_X1_4091_ (
  .A1({ S23626 }),
  .A2({ S23629 }),
  .ZN({ S25957[909] })
);
NAND2_X1 #() 
NAND2_X1_4092_ (
  .A1({ S21085 }),
  .A2({ S21089 }),
  .ZN({ S23630 })
);
XNOR2_X1 #() 
XNOR2_X1_172_ (
  .A({ S23630 }),
  .B({ S25957[1196] }),
  .ZN({ S25957[1068] })
);
NAND2_X1 #() 
NAND2_X1_4093_ (
  .A1({ S21088 }),
  .A2({ S21087 }),
  .ZN({ S25957[1132] })
);
INV_X1 #() 
INV_X1_1344_ (
  .A({ S25957[1132] }),
  .ZN({ S23631 })
);
NAND3_X1 #() 
NAND3_X1_4387_ (
  .A1({ S23387 }),
  .A2({ S23386 }),
  .A3({ S80 }),
  .ZN({ S23632 })
);
NAND2_X1 #() 
NAND2_X1_4094_ (
  .A1({ S23632 }),
  .A2({ S23423 }),
  .ZN({ S23633 })
);
NOR2_X1 #() 
NOR2_X1_1046_ (
  .A1({ S23554 }),
  .A2({ S23396 }),
  .ZN({ S23634 })
);
NOR2_X1 #() 
NOR2_X1_1047_ (
  .A1({ S25957[1025] }),
  .A2({ S80 }),
  .ZN({ S23635 })
);
NAND2_X1 #() 
NAND2_X1_4095_ (
  .A1({ S23635 }),
  .A2({ S23447 }),
  .ZN({ S23636 })
);
NAND2_X1 #() 
NAND2_X1_4096_ (
  .A1({ S23634 }),
  .A2({ S23636 }),
  .ZN({ S23637 })
);
OAI21_X1 #() 
OAI21_X1_2105_ (
  .A({ S23637 }),
  .B1({ S25957[1028] }),
  .B2({ S23633 }),
  .ZN({ S23638 })
);
NAND2_X1 #() 
NAND2_X1_4097_ (
  .A1({ S23531 }),
  .A2({ S80 }),
  .ZN({ S23639 })
);
NAND3_X1 #() 
NAND3_X1_4388_ (
  .A1({ S23639 }),
  .A2({ S23433 }),
  .A3({ S25957[1028] }),
  .ZN({ S23640 })
);
NAND3_X1 #() 
NAND3_X1_4389_ (
  .A1({ S23422 }),
  .A2({ S80 }),
  .A3({ S23360 }),
  .ZN({ S23641 })
);
NAND3_X1 #() 
NAND3_X1_4390_ (
  .A1({ S23426 }),
  .A2({ S23396 }),
  .A3({ S23641 }),
  .ZN({ S23642 })
);
NAND3_X1 #() 
NAND3_X1_4391_ (
  .A1({ S23642 }),
  .A2({ S25957[1029] }),
  .A3({ S23640 }),
  .ZN({ S23643 })
);
OAI211_X1 #() 
OAI211_X1_1424_ (
  .A({ S25957[1030] }),
  .B({ S23643 }),
  .C1({ S23638 }),
  .C2({ S25957[1029] }),
  .ZN({ S23644 })
);
AOI21_X1 #() 
AOI21_X1_2197_ (
  .A({ S25957[1027] }),
  .B1({ S23399 }),
  .B2({ S23376 }),
  .ZN({ S23645 })
);
NAND4_X1 #() 
NAND4_X1_479_ (
  .A1({ S25957[1027] }),
  .A2({ S25957[1025] }),
  .A3({ S23360 }),
  .A4({ S25957[1026] }),
  .ZN({ S23646 })
);
NAND2_X1 #() 
NAND2_X1_4098_ (
  .A1({ S23433 }),
  .A2({ S23646 }),
  .ZN({ S23647 })
);
NOR3_X1 #() 
NOR3_X1_141_ (
  .A1({ S23645 }),
  .A2({ S23647 }),
  .A3({ S25957[1028] }),
  .ZN({ S23648 })
);
OAI21_X1 #() 
OAI21_X1_2106_ (
  .A({ S23591 }),
  .B1({ S23599 }),
  .B2({ S23397 }),
  .ZN({ S23649 })
);
AOI21_X1 #() 
AOI21_X1_2198_ (
  .A({ S23368 }),
  .B1({ S23649 }),
  .B2({ S25957[1028] }),
  .ZN({ S23650 })
);
INV_X1 #() 
INV_X1_1345_ (
  .A({ S23650 }),
  .ZN({ S23651 })
);
NAND3_X1 #() 
NAND3_X1_4392_ (
  .A1({ S23409 }),
  .A2({ S80 }),
  .A3({ S23509 }),
  .ZN({ S23652 })
);
AOI21_X1 #() 
AOI21_X1_2199_ (
  .A({ S80 }),
  .B1({ S25957[1024] }),
  .B2({ S25957[1026] }),
  .ZN({ S23653 })
);
NAND3_X1 #() 
NAND3_X1_4393_ (
  .A1({ S23653 }),
  .A2({ S23422 }),
  .A3({ S23370 }),
  .ZN({ S23654 })
);
NAND3_X1 #() 
NAND3_X1_4394_ (
  .A1({ S23654 }),
  .A2({ S25957[1028] }),
  .A3({ S23652 }),
  .ZN({ S23655 })
);
OAI21_X1 #() 
OAI21_X1_2107_ (
  .A({ S80 }),
  .B1({ S23408 }),
  .B2({ S23539 }),
  .ZN({ S23656 })
);
AOI21_X1 #() 
AOI21_X1_2200_ (
  .A({ S25957[1028] }),
  .B1({ S23653 }),
  .B2({ S23361 }),
  .ZN({ S23657 })
);
AOI21_X1 #() 
AOI21_X1_2201_ (
  .A({ S25957[1029] }),
  .B1({ S23656 }),
  .B2({ S23657 }),
  .ZN({ S23658 })
);
NAND2_X1 #() 
NAND2_X1_4099_ (
  .A1({ S23658 }),
  .A2({ S23655 }),
  .ZN({ S23659 })
);
OAI211_X1 #() 
OAI211_X1_1425_ (
  .A({ S23659 }),
  .B({ S21581 }),
  .C1({ S23648 }),
  .C2({ S23651 }),
  .ZN({ S23660 })
);
NAND3_X1 #() 
NAND3_X1_4395_ (
  .A1({ S23660 }),
  .A2({ S23644 }),
  .A3({ S25957[1031] }),
  .ZN({ S23661 })
);
NAND3_X1 #() 
NAND3_X1_4396_ (
  .A1({ S23437 }),
  .A2({ S25957[1028] }),
  .A3({ S23553 }),
  .ZN({ S23662 })
);
INV_X1 #() 
INV_X1_1346_ (
  .A({ S23493 }),
  .ZN({ S23663 })
);
AOI21_X1 #() 
AOI21_X1_2202_ (
  .A({ S23662 }),
  .B1({ S23386 }),
  .B2({ S23663 }),
  .ZN({ S23664 })
);
INV_X1 #() 
INV_X1_1347_ (
  .A({ S125 }),
  .ZN({ S23665 })
);
OAI21_X1 #() 
OAI21_X1_2108_ (
  .A({ S25957[1028] }),
  .B1({ S23665 }),
  .B2({ S25957[1026] }),
  .ZN({ S23666 })
);
OAI21_X1 #() 
OAI21_X1_2109_ (
  .A({ S25957[1026] }),
  .B1({ S25957[1024] }),
  .B2({ S23361 }),
  .ZN({ S23667 })
);
AOI21_X1 #() 
AOI21_X1_2203_ (
  .A({ S25957[1027] }),
  .B1({ S23454 }),
  .B2({ S23667 }),
  .ZN({ S23668 })
);
NAND2_X1 #() 
NAND2_X1_4100_ (
  .A1({ S23608 }),
  .A2({ S23396 }),
  .ZN({ S23669 })
);
OAI211_X1 #() 
OAI211_X1_1426_ (
  .A({ S25957[1029] }),
  .B({ S23666 }),
  .C1({ S23669 }),
  .C2({ S23668 }),
  .ZN({ S23670 })
);
AOI21_X1 #() 
AOI21_X1_2204_ (
  .A({ S25957[1027] }),
  .B1({ S23419 }),
  .B2({ S23369 }),
  .ZN({ S23671 })
);
NAND2_X1 #() 
NAND2_X1_4101_ (
  .A1({ S23557 }),
  .A2({ S23396 }),
  .ZN({ S23672 })
);
OAI21_X1 #() 
OAI21_X1_2110_ (
  .A({ S23368 }),
  .B1({ S23671 }),
  .B2({ S23672 }),
  .ZN({ S23673 })
);
OAI211_X1 #() 
OAI211_X1_1427_ (
  .A({ S23670 }),
  .B({ S25957[1030] }),
  .C1({ S23664 }),
  .C2({ S23673 }),
  .ZN({ S23674 })
);
NOR3_X1 #() 
NOR3_X1_142_ (
  .A1({ S23458 }),
  .A2({ S23391 }),
  .A3({ S25957[1024] }),
  .ZN({ S23675 })
);
NAND2_X1 #() 
NAND2_X1_4102_ (
  .A1({ S23653 }),
  .A2({ S88 }),
  .ZN({ S23676 })
);
OAI21_X1 #() 
OAI21_X1_2111_ (
  .A({ S23676 }),
  .B1({ S23675 }),
  .B2({ S23460 }),
  .ZN({ S23677 })
);
NAND2_X1 #() 
NAND2_X1_4103_ (
  .A1({ S23677 }),
  .A2({ S23396 }),
  .ZN({ S23678 })
);
NAND2_X1 #() 
NAND2_X1_4104_ (
  .A1({ S23653 }),
  .A2({ S23507 }),
  .ZN({ S23679 })
);
AOI21_X1 #() 
AOI21_X1_2205_ (
  .A({ S25957[1029] }),
  .B1({ S23634 }),
  .B2({ S23679 }),
  .ZN({ S23680 })
);
NOR2_X1 #() 
NOR2_X1_1048_ (
  .A1({ S23359 }),
  .A2({ S25957[1027] }),
  .ZN({ S23681 })
);
OAI21_X1 #() 
OAI21_X1_2112_ (
  .A({ S23396 }),
  .B1({ S23566 }),
  .B2({ S23681 }),
  .ZN({ S23682 })
);
INV_X1 #() 
INV_X1_1348_ (
  .A({ S23383 }),
  .ZN({ S23683 })
);
AOI21_X1 #() 
AOI21_X1_2206_ (
  .A({ S23396 }),
  .B1({ S23581 }),
  .B2({ S80 }),
  .ZN({ S23684 })
);
AOI21_X1 #() 
AOI21_X1_2207_ (
  .A({ S23368 }),
  .B1({ S23683 }),
  .B2({ S23684 }),
  .ZN({ S23685 })
);
AOI22_X1 #() 
AOI22_X1_468_ (
  .A1({ S23678 }),
  .A2({ S23680 }),
  .B1({ S23685 }),
  .B2({ S23682 }),
  .ZN({ S23686 })
);
OAI211_X1 #() 
OAI211_X1_1428_ (
  .A({ S23674 }),
  .B({ S21512 }),
  .C1({ S23686 }),
  .C2({ S25957[1030] }),
  .ZN({ S23687 })
);
NAND3_X1 #() 
NAND3_X1_4397_ (
  .A1({ S23661 }),
  .A2({ S23687 }),
  .A3({ S23631 }),
  .ZN({ S23688 })
);
INV_X1 #() 
INV_X1_1349_ (
  .A({ S23668 }),
  .ZN({ S23689 })
);
INV_X1 #() 
INV_X1_1350_ (
  .A({ S23669 }),
  .ZN({ S23690 })
);
NAND2_X1 #() 
NAND2_X1_4105_ (
  .A1({ S23666 }),
  .A2({ S25957[1029] }),
  .ZN({ S23691 })
);
AOI21_X1 #() 
AOI21_X1_2208_ (
  .A({ S23691 }),
  .B1({ S23690 }),
  .B2({ S23689 }),
  .ZN({ S23692 })
);
NOR2_X1 #() 
NOR2_X1_1049_ (
  .A1({ S23664 }),
  .A2({ S23673 }),
  .ZN({ S23693 })
);
OAI21_X1 #() 
OAI21_X1_2113_ (
  .A({ S25957[1030] }),
  .B1({ S23693 }),
  .B2({ S23692 }),
  .ZN({ S23694 })
);
NAND2_X1 #() 
NAND2_X1_4106_ (
  .A1({ S23678 }),
  .A2({ S23680 }),
  .ZN({ S23695 })
);
NAND2_X1 #() 
NAND2_X1_4107_ (
  .A1({ S23685 }),
  .A2({ S23682 }),
  .ZN({ S23696 })
);
NAND3_X1 #() 
NAND3_X1_4398_ (
  .A1({ S23695 }),
  .A2({ S23696 }),
  .A3({ S21581 }),
  .ZN({ S23697 })
);
NAND3_X1 #() 
NAND3_X1_4399_ (
  .A1({ S23694 }),
  .A2({ S23697 }),
  .A3({ S21512 }),
  .ZN({ S23698 })
);
OR3_X1 #() 
OR3_X1_27_ (
  .A1({ S23645 }),
  .A2({ S23647 }),
  .A3({ S25957[1028] }),
  .ZN({ S23699 })
);
AOI22_X1 #() 
AOI22_X1_469_ (
  .A1({ S23699 }),
  .A2({ S23650 }),
  .B1({ S23655 }),
  .B2({ S23658 }),
  .ZN({ S23700 })
);
AOI21_X1 #() 
AOI21_X1_2209_ (
  .A({ S23554 }),
  .B1({ S23635 }),
  .B2({ S23447 }),
  .ZN({ S23701 })
);
NAND2_X1 #() 
NAND2_X1_4108_ (
  .A1({ S23633 }),
  .A2({ S23396 }),
  .ZN({ S23702 })
);
OAI211_X1 #() 
OAI211_X1_1429_ (
  .A({ S23702 }),
  .B({ S23368 }),
  .C1({ S23701 }),
  .C2({ S23396 }),
  .ZN({ S23703 })
);
NAND2_X1 #() 
NAND2_X1_4109_ (
  .A1({ S23642 }),
  .A2({ S23640 }),
  .ZN({ S23704 })
);
NAND2_X1 #() 
NAND2_X1_4110_ (
  .A1({ S23704 }),
  .A2({ S25957[1029] }),
  .ZN({ S23705 })
);
NAND3_X1 #() 
NAND3_X1_4400_ (
  .A1({ S23703 }),
  .A2({ S23705 }),
  .A3({ S25957[1030] }),
  .ZN({ S23706 })
);
OAI211_X1 #() 
OAI211_X1_1430_ (
  .A({ S23706 }),
  .B({ S25957[1031] }),
  .C1({ S23700 }),
  .C2({ S25957[1030] }),
  .ZN({ S23707 })
);
NAND3_X1 #() 
NAND3_X1_4401_ (
  .A1({ S23707 }),
  .A2({ S25957[1132] }),
  .A3({ S23698 }),
  .ZN({ S23708 })
);
AOI21_X1 #() 
AOI21_X1_2210_ (
  .A({ S23630 }),
  .B1({ S23708 }),
  .B2({ S23688 }),
  .ZN({ S23709 })
);
INV_X1 #() 
INV_X1_1351_ (
  .A({ S23630 }),
  .ZN({ S25957[1100] })
);
NAND3_X1 #() 
NAND3_X1_4402_ (
  .A1({ S23661 }),
  .A2({ S23687 }),
  .A3({ S25957[1132] }),
  .ZN({ S23710 })
);
NAND3_X1 #() 
NAND3_X1_4403_ (
  .A1({ S23707 }),
  .A2({ S23631 }),
  .A3({ S23698 }),
  .ZN({ S23711 })
);
AOI21_X1 #() 
AOI21_X1_2211_ (
  .A({ S25957[1100] }),
  .B1({ S23711 }),
  .B2({ S23710 }),
  .ZN({ S23712 })
);
OAI21_X1 #() 
OAI21_X1_2114_ (
  .A({ S25957[1164] }),
  .B1({ S23709 }),
  .B2({ S23712 }),
  .ZN({ S23713 })
);
NAND3_X1 #() 
NAND3_X1_4404_ (
  .A1({ S23711 }),
  .A2({ S23710 }),
  .A3({ S25957[1100] }),
  .ZN({ S23714 })
);
NAND3_X1 #() 
NAND3_X1_4405_ (
  .A1({ S23708 }),
  .A2({ S23688 }),
  .A3({ S23630 }),
  .ZN({ S23715 })
);
NAND3_X1 #() 
NAND3_X1_4406_ (
  .A1({ S23714 }),
  .A2({ S23715 }),
  .A3({ S20131 }),
  .ZN({ S23716 })
);
NAND2_X1 #() 
NAND2_X1_4111_ (
  .A1({ S23713 }),
  .A2({ S23716 }),
  .ZN({ S25957[908] })
);
NAND2_X1 #() 
NAND2_X1_4112_ (
  .A1({ S21182 }),
  .A2({ S21183 }),
  .ZN({ S23717 })
);
INV_X1 #() 
INV_X1_1352_ (
  .A({ S23717 }),
  .ZN({ S25957[1067] })
);
NAND3_X1 #() 
NAND3_X1_4407_ (
  .A1({ S23410 }),
  .A2({ S80 }),
  .A3({ S23507 }),
  .ZN({ S23718 })
);
AOI21_X1 #() 
AOI21_X1_2212_ (
  .A({ S23396 }),
  .B1({ S23435 }),
  .B2({ S25957[1027] }),
  .ZN({ S23719 })
);
NOR2_X1 #() 
NOR2_X1_1050_ (
  .A1({ S23672 }),
  .A2({ S23516 }),
  .ZN({ S23720 })
);
AOI21_X1 #() 
AOI21_X1_2213_ (
  .A({ S23720 }),
  .B1({ S23719 }),
  .B2({ S23718 }),
  .ZN({ S23721 })
);
NAND3_X1 #() 
NAND3_X1_4408_ (
  .A1({ S23398 }),
  .A2({ S25957[1027] }),
  .A3({ S23447 }),
  .ZN({ S23722 })
);
NAND2_X1 #() 
NAND2_X1_4113_ (
  .A1({ S23439 }),
  .A2({ S80 }),
  .ZN({ S23723 })
);
NAND3_X1 #() 
NAND3_X1_4409_ (
  .A1({ S23723 }),
  .A2({ S25957[1028] }),
  .A3({ S23722 }),
  .ZN({ S23724 })
);
OAI211_X1 #() 
OAI211_X1_1431_ (
  .A({ S80 }),
  .B({ S23397 }),
  .C1({ S23391 }),
  .C2({ S25957[1024] }),
  .ZN({ S23725 })
);
OAI211_X1 #() 
OAI211_X1_1432_ (
  .A({ S23396 }),
  .B({ S23725 }),
  .C1({ S23502 }),
  .C2({ S23482 }),
  .ZN({ S23726 })
);
NAND3_X1 #() 
NAND3_X1_4410_ (
  .A1({ S23724 }),
  .A2({ S23726 }),
  .A3({ S25957[1029] }),
  .ZN({ S23727 })
);
OAI211_X1 #() 
OAI211_X1_1433_ (
  .A({ S23727 }),
  .B({ S25957[1030] }),
  .C1({ S23721 }),
  .C2({ S25957[1029] }),
  .ZN({ S23728 })
);
NAND3_X1 #() 
NAND3_X1_4411_ (
  .A1({ S23410 }),
  .A2({ S80 }),
  .A3({ S23386 }),
  .ZN({ S23729 })
);
NAND4_X1 #() 
NAND4_X1_480_ (
  .A1({ S23387 }),
  .A2({ S23447 }),
  .A3({ S25957[1025] }),
  .A4({ S25957[1027] }),
  .ZN({ S23730 })
);
AND2_X1 #() 
AND2_X1_258_ (
  .A1({ S23730 }),
  .A2({ S23396 }),
  .ZN({ S23731 })
);
NAND3_X1 #() 
NAND3_X1_4412_ (
  .A1({ S23454 }),
  .A2({ S25957[1027] }),
  .A3({ S23531 }),
  .ZN({ S23732 })
);
AOI21_X1 #() 
AOI21_X1_2214_ (
  .A({ S23396 }),
  .B1({ S23482 }),
  .B2({ S80 }),
  .ZN({ S23733 })
);
AOI22_X1 #() 
AOI22_X1_470_ (
  .A1({ S23731 }),
  .A2({ S23729 }),
  .B1({ S23733 }),
  .B2({ S23732 }),
  .ZN({ S23734 })
);
NAND3_X1 #() 
NAND3_X1_4413_ (
  .A1({ S23539 }),
  .A2({ S25957[1027] }),
  .A3({ S23397 }),
  .ZN({ S23735 })
);
NAND2_X1 #() 
NAND2_X1_4114_ (
  .A1({ S23388 }),
  .A2({ S80 }),
  .ZN({ S23736 })
);
NAND3_X1 #() 
NAND3_X1_4414_ (
  .A1({ S23735 }),
  .A2({ S23736 }),
  .A3({ S25957[1028] }),
  .ZN({ S23737 })
);
NAND3_X1 #() 
NAND3_X1_4415_ (
  .A1({ S23415 }),
  .A2({ S23398 }),
  .A3({ S23397 }),
  .ZN({ S23738 })
);
NAND3_X1 #() 
NAND3_X1_4416_ (
  .A1({ S88 }),
  .A2({ S80 }),
  .A3({ S23447 }),
  .ZN({ S23739 })
);
AOI21_X1 #() 
AOI21_X1_2215_ (
  .A({ S25957[1028] }),
  .B1({ S23635 }),
  .B2({ S23381 }),
  .ZN({ S23740 })
);
NAND3_X1 #() 
NAND3_X1_4417_ (
  .A1({ S23740 }),
  .A2({ S23738 }),
  .A3({ S23739 }),
  .ZN({ S23741 })
);
NAND3_X1 #() 
NAND3_X1_4418_ (
  .A1({ S23737 }),
  .A2({ S23741 }),
  .A3({ S23368 }),
  .ZN({ S23742 })
);
OAI211_X1 #() 
OAI211_X1_1434_ (
  .A({ S21581 }),
  .B({ S23742 }),
  .C1({ S23734 }),
  .C2({ S23368 }),
  .ZN({ S23743 })
);
NAND3_X1 #() 
NAND3_X1_4419_ (
  .A1({ S23743 }),
  .A2({ S23728 }),
  .A3({ S25957[1031] }),
  .ZN({ S23744 })
);
NAND3_X1 #() 
NAND3_X1_4420_ (
  .A1({ S23428 }),
  .A2({ S23422 }),
  .A3({ S23370 }),
  .ZN({ S23745 })
);
NAND3_X1 #() 
NAND3_X1_4421_ (
  .A1({ S23745 }),
  .A2({ S23575 }),
  .A3({ S23433 }),
  .ZN({ S23746 })
);
OAI21_X1 #() 
OAI21_X1_2115_ (
  .A({ S80 }),
  .B1({ S23391 }),
  .B2({ S23360 }),
  .ZN({ S23747 })
);
AOI21_X1 #() 
AOI21_X1_2216_ (
  .A({ S25957[1029] }),
  .B1({ S23747 }),
  .B2({ S25957[1028] }),
  .ZN({ S23748 })
);
NAND2_X1 #() 
NAND2_X1_4115_ (
  .A1({ S23746 }),
  .A2({ S23748 }),
  .ZN({ S23749 })
);
NAND2_X1 #() 
NAND2_X1_4116_ (
  .A1({ S23483 }),
  .A2({ S23411 }),
  .ZN({ S23750 })
);
NAND3_X1 #() 
NAND3_X1_4422_ (
  .A1({ S23397 }),
  .A2({ S80 }),
  .A3({ S23422 }),
  .ZN({ S23751 })
);
AOI21_X1 #() 
AOI21_X1_2217_ (
  .A({ S25957[1028] }),
  .B1({ S23589 }),
  .B2({ S23380 }),
  .ZN({ S23752 })
);
NAND2_X1 #() 
NAND2_X1_4117_ (
  .A1({ S23752 }),
  .A2({ S23751 }),
  .ZN({ S23753 })
);
NAND3_X1 #() 
NAND3_X1_4423_ (
  .A1({ S23750 }),
  .A2({ S25957[1029] }),
  .A3({ S23753 }),
  .ZN({ S23754 })
);
NAND3_X1 #() 
NAND3_X1_4424_ (
  .A1({ S23754 }),
  .A2({ S25957[1030] }),
  .A3({ S23749 }),
  .ZN({ S23755 })
);
NAND2_X1 #() 
NAND2_X1_4118_ (
  .A1({ S23396 }),
  .A2({ S80 }),
  .ZN({ S23756 })
);
NAND3_X1 #() 
NAND3_X1_4425_ (
  .A1({ S23419 }),
  .A2({ S23396 }),
  .A3({ S23369 }),
  .ZN({ S23757 })
);
AOI22_X1 #() 
AOI22_X1_471_ (
  .A1({ S23403 }),
  .A2({ S80 }),
  .B1({ S23757 }),
  .B2({ S23756 }),
  .ZN({ S23758 })
);
OAI211_X1 #() 
OAI211_X1_1435_ (
  .A({ S88 }),
  .B({ S25957[1027] }),
  .C1({ S25957[1026] }),
  .C2({ S23359 }),
  .ZN({ S23759 })
);
NAND3_X1 #() 
NAND3_X1_4426_ (
  .A1({ S23759 }),
  .A2({ S23593 }),
  .A3({ S25957[1028] }),
  .ZN({ S23760 })
);
NAND2_X1 #() 
NAND2_X1_4119_ (
  .A1({ S23760 }),
  .A2({ S23368 }),
  .ZN({ S23761 })
);
NAND4_X1 #() 
NAND4_X1_481_ (
  .A1({ S23534 }),
  .A2({ S23422 }),
  .A3({ S25957[1024] }),
  .A4({ S23396 }),
  .ZN({ S23762 })
);
OAI211_X1 #() 
OAI211_X1_1436_ (
  .A({ S25957[1028] }),
  .B({ S25957[1026] }),
  .C1({ S23681 }),
  .C2({ S23492 }),
  .ZN({ S23763 })
);
NAND3_X1 #() 
NAND3_X1_4427_ (
  .A1({ S23763 }),
  .A2({ S23762 }),
  .A3({ S25957[1029] }),
  .ZN({ S23764 })
);
OAI211_X1 #() 
OAI211_X1_1437_ (
  .A({ S21581 }),
  .B({ S23764 }),
  .C1({ S23758 }),
  .C2({ S23761 }),
  .ZN({ S23765 })
);
NAND3_X1 #() 
NAND3_X1_4428_ (
  .A1({ S23755 }),
  .A2({ S21512 }),
  .A3({ S23765 }),
  .ZN({ S23766 })
);
AND3_X1 #() 
AND3_X1_160_ (
  .A1({ S23744 }),
  .A2({ S23766 }),
  .A3({ S21173 }),
  .ZN({ S23767 })
);
AOI21_X1 #() 
AOI21_X1_2218_ (
  .A({ S21173 }),
  .B1({ S23744 }),
  .B2({ S23766 }),
  .ZN({ S23768 })
);
OAI21_X1 #() 
OAI21_X1_2116_ (
  .A({ S25957[1067] }),
  .B1({ S23767 }),
  .B2({ S23768 }),
  .ZN({ S23769 })
);
NAND3_X1 #() 
NAND3_X1_4429_ (
  .A1({ S23744 }),
  .A2({ S23766 }),
  .A3({ S21173 }),
  .ZN({ S23770 })
);
NAND2_X1 #() 
NAND2_X1_4120_ (
  .A1({ S23755 }),
  .A2({ S23765 }),
  .ZN({ S23771 })
);
NAND2_X1 #() 
NAND2_X1_4121_ (
  .A1({ S23771 }),
  .A2({ S21512 }),
  .ZN({ S23772 })
);
NAND2_X1 #() 
NAND2_X1_4122_ (
  .A1({ S23718 }),
  .A2({ S23719 }),
  .ZN({ S23773 })
);
INV_X1 #() 
INV_X1_1353_ (
  .A({ S23720 }),
  .ZN({ S23774 })
);
AOI21_X1 #() 
AOI21_X1_2219_ (
  .A({ S25957[1029] }),
  .B1({ S23773 }),
  .B2({ S23774 }),
  .ZN({ S23775 })
);
INV_X1 #() 
INV_X1_1354_ (
  .A({ S23727 }),
  .ZN({ S23776 })
);
OAI21_X1 #() 
OAI21_X1_2117_ (
  .A({ S25957[1030] }),
  .B1({ S23776 }),
  .B2({ S23775 }),
  .ZN({ S23777 })
);
NAND2_X1 #() 
NAND2_X1_4123_ (
  .A1({ S23731 }),
  .A2({ S23729 }),
  .ZN({ S23778 })
);
NAND2_X1 #() 
NAND2_X1_4124_ (
  .A1({ S23733 }),
  .A2({ S23732 }),
  .ZN({ S23779 })
);
AOI21_X1 #() 
AOI21_X1_2220_ (
  .A({ S23368 }),
  .B1({ S23778 }),
  .B2({ S23779 }),
  .ZN({ S23780 })
);
INV_X1 #() 
INV_X1_1355_ (
  .A({ S23742 }),
  .ZN({ S23781 })
);
OAI21_X1 #() 
OAI21_X1_2118_ (
  .A({ S21581 }),
  .B1({ S23780 }),
  .B2({ S23781 }),
  .ZN({ S23782 })
);
NAND3_X1 #() 
NAND3_X1_4430_ (
  .A1({ S23782 }),
  .A2({ S25957[1031] }),
  .A3({ S23777 }),
  .ZN({ S23783 })
);
NAND3_X1 #() 
NAND3_X1_4431_ (
  .A1({ S23783 }),
  .A2({ S23772 }),
  .A3({ S25957[1227] }),
  .ZN({ S23784 })
);
NAND3_X1 #() 
NAND3_X1_4432_ (
  .A1({ S23784 }),
  .A2({ S23717 }),
  .A3({ S23770 }),
  .ZN({ S23785 })
);
NAND3_X1 #() 
NAND3_X1_4433_ (
  .A1({ S23769 }),
  .A2({ S23785 }),
  .A3({ S25957[1035] }),
  .ZN({ S23786 })
);
NAND2_X1 #() 
NAND2_X1_4125_ (
  .A1({ S21175 }),
  .A2({ S21174 }),
  .ZN({ S25957[1131] })
);
AND3_X1 #() 
AND3_X1_161_ (
  .A1({ S23744 }),
  .A2({ S23766 }),
  .A3({ S25957[1131] }),
  .ZN({ S23787 })
);
AOI21_X1 #() 
AOI21_X1_2221_ (
  .A({ S25957[1131] }),
  .B1({ S23744 }),
  .B2({ S23766 }),
  .ZN({ S23788 })
);
OAI21_X1 #() 
OAI21_X1_2119_ (
  .A({ S25957[1195] }),
  .B1({ S23787 }),
  .B2({ S23788 }),
  .ZN({ S23789 })
);
NAND3_X1 #() 
NAND3_X1_4434_ (
  .A1({ S23744 }),
  .A2({ S23766 }),
  .A3({ S25957[1131] }),
  .ZN({ S23790 })
);
INV_X1 #() 
INV_X1_1356_ (
  .A({ S25957[1131] }),
  .ZN({ S23791 })
);
NAND3_X1 #() 
NAND3_X1_4435_ (
  .A1({ S23783 }),
  .A2({ S23772 }),
  .A3({ S23791 }),
  .ZN({ S23792 })
);
NAND3_X1 #() 
NAND3_X1_4436_ (
  .A1({ S23792 }),
  .A2({ S21094 }),
  .A3({ S23790 }),
  .ZN({ S23793 })
);
NAND3_X1 #() 
NAND3_X1_4437_ (
  .A1({ S23789 }),
  .A2({ S23793 }),
  .A3({ S77 }),
  .ZN({ S23794 })
);
NAND2_X1 #() 
NAND2_X1_4126_ (
  .A1({ S23786 }),
  .A2({ S23794 }),
  .ZN({ S89 })
);
NAND3_X1 #() 
NAND3_X1_4438_ (
  .A1({ S23769 }),
  .A2({ S23785 }),
  .A3({ S77 }),
  .ZN({ S23795 })
);
NAND3_X1 #() 
NAND3_X1_4439_ (
  .A1({ S23789 }),
  .A2({ S23793 }),
  .A3({ S25957[1035] }),
  .ZN({ S23796 })
);
NAND2_X1 #() 
NAND2_X1_4127_ (
  .A1({ S23795 }),
  .A2({ S23796 }),
  .ZN({ S25957[907] })
);
NAND2_X1 #() 
NAND2_X1_4128_ (
  .A1({ S23391 }),
  .A2({ S80 }),
  .ZN({ S23797 })
);
NAND3_X1 #() 
NAND3_X1_4440_ (
  .A1({ S23733 }),
  .A2({ S23797 }),
  .A3({ S23738 }),
  .ZN({ S23798 })
);
AOI21_X1 #() 
AOI21_X1_2222_ (
  .A({ S25957[1028] }),
  .B1({ S80 }),
  .B2({ S23401 }),
  .ZN({ S23799 })
);
NAND3_X1 #() 
NAND3_X1_4441_ (
  .A1({ S23376 }),
  .A2({ S23447 }),
  .A3({ S23464 }),
  .ZN({ S23800 })
);
AOI21_X1 #() 
AOI21_X1_2223_ (
  .A({ S25957[1029] }),
  .B1({ S23799 }),
  .B2({ S23800 }),
  .ZN({ S23801 })
);
NAND2_X1 #() 
NAND2_X1_4129_ (
  .A1({ S23415 }),
  .A2({ S23398 }),
  .ZN({ S23802 })
);
OAI211_X1 #() 
OAI211_X1_1438_ (
  .A({ S25957[1028] }),
  .B({ S23802 }),
  .C1({ S23675 }),
  .C2({ S23460 }),
  .ZN({ S23803 })
);
NAND3_X1 #() 
NAND3_X1_4442_ (
  .A1({ S23399 }),
  .A2({ S80 }),
  .A3({ S23370 }),
  .ZN({ S23804 })
);
AOI21_X1 #() 
AOI21_X1_2224_ (
  .A({ S25957[1028] }),
  .B1({ S23653 }),
  .B2({ S23507 }),
  .ZN({ S23805 })
);
AOI21_X1 #() 
AOI21_X1_2225_ (
  .A({ S23368 }),
  .B1({ S23804 }),
  .B2({ S23805 }),
  .ZN({ S23806 })
);
AOI22_X1 #() 
AOI22_X1_472_ (
  .A1({ S23806 }),
  .A2({ S23803 }),
  .B1({ S23798 }),
  .B2({ S23801 }),
  .ZN({ S23807 })
);
OAI211_X1 #() 
OAI211_X1_1439_ (
  .A({ S25957[1028] }),
  .B({ S23497 }),
  .C1({ S23413 }),
  .C2({ S23600 }),
  .ZN({ S23808 })
);
NAND2_X1 #() 
NAND2_X1_4130_ (
  .A1({ S25957[1027] }),
  .A2({ S23360 }),
  .ZN({ S23809 })
);
NOR2_X1 #() 
NOR2_X1_1051_ (
  .A1({ S23809 }),
  .A2({ S23458 }),
  .ZN({ S23810 })
);
AOI21_X1 #() 
AOI21_X1_2226_ (
  .A({ S25957[1027] }),
  .B1({ S23509 }),
  .B2({ S23447 }),
  .ZN({ S23811 })
);
OAI21_X1 #() 
OAI21_X1_2120_ (
  .A({ S23396 }),
  .B1({ S23811 }),
  .B2({ S23810 }),
  .ZN({ S23812 })
);
NAND3_X1 #() 
NAND3_X1_4443_ (
  .A1({ S23812 }),
  .A2({ S23808 }),
  .A3({ S23368 }),
  .ZN({ S23813 })
);
NAND3_X1 #() 
NAND3_X1_4444_ (
  .A1({ S23639 }),
  .A2({ S23433 }),
  .A3({ S23646 }),
  .ZN({ S23814 })
);
NAND2_X1 #() 
NAND2_X1_4131_ (
  .A1({ S23814 }),
  .A2({ S23396 }),
  .ZN({ S23815 })
);
NAND2_X1 #() 
NAND2_X1_4132_ (
  .A1({ S23747 }),
  .A2({ S23532 }),
  .ZN({ S23816 })
);
NAND3_X1 #() 
NAND3_X1_4445_ (
  .A1({ S23380 }),
  .A2({ S80 }),
  .A3({ S23360 }),
  .ZN({ S23817 })
);
AND2_X1 #() 
AND2_X1_259_ (
  .A1({ S23817 }),
  .A2({ S25957[1028] }),
  .ZN({ S23818 })
);
NAND2_X1 #() 
NAND2_X1_4133_ (
  .A1({ S23816 }),
  .A2({ S23818 }),
  .ZN({ S23819 })
);
NAND3_X1 #() 
NAND3_X1_4446_ (
  .A1({ S23815 }),
  .A2({ S23819 }),
  .A3({ S25957[1029] }),
  .ZN({ S23820 })
);
NAND3_X1 #() 
NAND3_X1_4447_ (
  .A1({ S23820 }),
  .A2({ S23813 }),
  .A3({ S21581 }),
  .ZN({ S23821 })
);
OAI211_X1 #() 
OAI211_X1_1440_ (
  .A({ S23821 }),
  .B({ S25957[1031] }),
  .C1({ S23807 }),
  .C2({ S21581 }),
  .ZN({ S23822 })
);
NAND2_X1 #() 
NAND2_X1_4134_ (
  .A1({ S23402 }),
  .A2({ S23602 }),
  .ZN({ S23823 })
);
OAI21_X1 #() 
OAI21_X1_2121_ (
  .A({ S80 }),
  .B1({ S23391 }),
  .B2({ S25957[1024] }),
  .ZN({ S23824 })
);
NAND3_X1 #() 
NAND3_X1_4448_ (
  .A1({ S23823 }),
  .A2({ S25957[1028] }),
  .A3({ S23824 }),
  .ZN({ S23825 })
);
NAND2_X1 #() 
NAND2_X1_4135_ (
  .A1({ S23540 }),
  .A2({ S23799 }),
  .ZN({ S23826 })
);
NAND3_X1 #() 
NAND3_X1_4449_ (
  .A1({ S23825 }),
  .A2({ S23826 }),
  .A3({ S25957[1029] }),
  .ZN({ S23827 })
);
NAND3_X1 #() 
NAND3_X1_4450_ (
  .A1({ S23608 }),
  .A2({ S23396 }),
  .A3({ S23576 }),
  .ZN({ S23828 })
);
NAND4_X1 #() 
NAND4_X1_482_ (
  .A1({ S23591 }),
  .A2({ S23809 }),
  .A3({ S25957[1028] }),
  .A4({ S23370 }),
  .ZN({ S23829 })
);
NAND2_X1 #() 
NAND2_X1_4136_ (
  .A1({ S23828 }),
  .A2({ S23829 }),
  .ZN({ S23830 })
);
NAND2_X1 #() 
NAND2_X1_4137_ (
  .A1({ S23830 }),
  .A2({ S23368 }),
  .ZN({ S23831 })
);
NAND3_X1 #() 
NAND3_X1_4451_ (
  .A1({ S23831 }),
  .A2({ S23827 }),
  .A3({ S25957[1030] }),
  .ZN({ S23832 })
);
NAND3_X1 #() 
NAND3_X1_4452_ (
  .A1({ S23382 }),
  .A2({ S23531 }),
  .A3({ S80 }),
  .ZN({ S23833 })
);
OAI211_X1 #() 
OAI211_X1_1441_ (
  .A({ S88 }),
  .B({ S25957[1027] }),
  .C1({ S23360 }),
  .C2({ S23380 }),
  .ZN({ S23834 })
);
AOI21_X1 #() 
AOI21_X1_2227_ (
  .A({ S25957[1029] }),
  .B1({ S23833 }),
  .B2({ S23834 }),
  .ZN({ S23835 })
);
NAND4_X1 #() 
NAND4_X1_483_ (
  .A1({ S23387 }),
  .A2({ S23447 }),
  .A3({ S23361 }),
  .A4({ S25957[1027] }),
  .ZN({ S23836 })
);
AND3_X1 #() 
AND3_X1_162_ (
  .A1({ S23596 }),
  .A2({ S25957[1029] }),
  .A3({ S23836 }),
  .ZN({ S23837 })
);
OAI21_X1 #() 
OAI21_X1_2122_ (
  .A({ S23396 }),
  .B1({ S23837 }),
  .B2({ S23835 }),
  .ZN({ S23838 })
);
AOI21_X1 #() 
AOI21_X1_2228_ (
  .A({ S23368 }),
  .B1({ S23444 }),
  .B2({ S23447 }),
  .ZN({ S23839 })
);
NAND3_X1 #() 
NAND3_X1_4453_ (
  .A1({ S23410 }),
  .A2({ S80 }),
  .A3({ S23422 }),
  .ZN({ S23840 })
);
AOI21_X1 #() 
AOI21_X1_2229_ (
  .A({ S25957[1029] }),
  .B1({ S23399 }),
  .B2({ S25957[1027] }),
  .ZN({ S23841 })
);
AOI22_X1 #() 
AOI22_X1_473_ (
  .A1({ S23841 }),
  .A2({ S23840 }),
  .B1({ S23839 }),
  .B2({ S23676 }),
  .ZN({ S23842 })
);
OAI211_X1 #() 
OAI211_X1_1442_ (
  .A({ S23838 }),
  .B({ S21581 }),
  .C1({ S23396 }),
  .C2({ S23842 }),
  .ZN({ S23843 })
);
NAND3_X1 #() 
NAND3_X1_4454_ (
  .A1({ S23843 }),
  .A2({ S21512 }),
  .A3({ S23832 }),
  .ZN({ S23844 })
);
AOI21_X1 #() 
AOI21_X1_2230_ (
  .A({ S21187 }),
  .B1({ S23844 }),
  .B2({ S23822 }),
  .ZN({ S23845 })
);
NAND2_X1 #() 
NAND2_X1_4138_ (
  .A1({ S23798 }),
  .A2({ S23801 }),
  .ZN({ S23846 })
);
NAND2_X1 #() 
NAND2_X1_4139_ (
  .A1({ S23806 }),
  .A2({ S23803 }),
  .ZN({ S23847 })
);
NAND3_X1 #() 
NAND3_X1_4455_ (
  .A1({ S23847 }),
  .A2({ S23846 }),
  .A3({ S25957[1030] }),
  .ZN({ S23848 })
);
AOI22_X1 #() 
AOI22_X1_474_ (
  .A1({ S23814 }),
  .A2({ S23396 }),
  .B1({ S23816 }),
  .B2({ S23818 }),
  .ZN({ S23849 })
);
NAND3_X1 #() 
NAND3_X1_4456_ (
  .A1({ S23667 }),
  .A2({ S80 }),
  .A3({ S23401 }),
  .ZN({ S23850 })
);
NAND2_X1 #() 
NAND2_X1_4140_ (
  .A1({ S23850 }),
  .A2({ S23752 }),
  .ZN({ S23851 })
);
NAND2_X1 #() 
NAND2_X1_4141_ (
  .A1({ S23380 }),
  .A2({ S25957[1027] }),
  .ZN({ S23852 })
);
NAND2_X1 #() 
NAND2_X1_4142_ (
  .A1({ S23454 }),
  .A2({ S80 }),
  .ZN({ S23853 })
);
NAND3_X1 #() 
NAND3_X1_4457_ (
  .A1({ S23853 }),
  .A2({ S25957[1028] }),
  .A3({ S23852 }),
  .ZN({ S23854 })
);
NAND3_X1 #() 
NAND3_X1_4458_ (
  .A1({ S23854 }),
  .A2({ S23851 }),
  .A3({ S23368 }),
  .ZN({ S23855 })
);
OAI211_X1 #() 
OAI211_X1_1443_ (
  .A({ S23855 }),
  .B({ S21581 }),
  .C1({ S23849 }),
  .C2({ S23368 }),
  .ZN({ S23856 })
);
NAND3_X1 #() 
NAND3_X1_4459_ (
  .A1({ S23848 }),
  .A2({ S23856 }),
  .A3({ S25957[1031] }),
  .ZN({ S23857 })
);
AOI21_X1 #() 
AOI21_X1_2231_ (
  .A({ S23396 }),
  .B1({ S23402 }),
  .B2({ S23602 }),
  .ZN({ S23858 })
);
AOI22_X1 #() 
AOI22_X1_475_ (
  .A1({ S23858 }),
  .A2({ S23824 }),
  .B1({ S23540 }),
  .B2({ S23799 }),
  .ZN({ S23859 })
);
NAND3_X1 #() 
NAND3_X1_4460_ (
  .A1({ S23828 }),
  .A2({ S23368 }),
  .A3({ S23829 }),
  .ZN({ S23860 })
);
OAI211_X1 #() 
OAI211_X1_1444_ (
  .A({ S25957[1030] }),
  .B({ S23860 }),
  .C1({ S23859 }),
  .C2({ S23368 }),
  .ZN({ S23861 })
);
NAND2_X1 #() 
NAND2_X1_4143_ (
  .A1({ S23444 }),
  .A2({ S23447 }),
  .ZN({ S23862 })
);
NAND3_X1 #() 
NAND3_X1_4461_ (
  .A1({ S23862 }),
  .A2({ S23676 }),
  .A3({ S25957[1028] }),
  .ZN({ S23863 })
);
NAND3_X1 #() 
NAND3_X1_4462_ (
  .A1({ S23596 }),
  .A2({ S23836 }),
  .A3({ S23396 }),
  .ZN({ S23864 })
);
NAND3_X1 #() 
NAND3_X1_4463_ (
  .A1({ S23863 }),
  .A2({ S25957[1029] }),
  .A3({ S23864 }),
  .ZN({ S23865 })
);
NAND2_X1 #() 
NAND2_X1_4144_ (
  .A1({ S23399 }),
  .A2({ S25957[1027] }),
  .ZN({ S23866 })
);
AOI21_X1 #() 
AOI21_X1_2232_ (
  .A({ S23396 }),
  .B1({ S23840 }),
  .B2({ S23866 }),
  .ZN({ S23867 })
);
AND3_X1 #() 
AND3_X1_163_ (
  .A1({ S23833 }),
  .A2({ S23834 }),
  .A3({ S23396 }),
  .ZN({ S23868 })
);
OAI21_X1 #() 
OAI21_X1_2123_ (
  .A({ S23368 }),
  .B1({ S23867 }),
  .B2({ S23868 }),
  .ZN({ S23869 })
);
NAND3_X1 #() 
NAND3_X1_4464_ (
  .A1({ S23869 }),
  .A2({ S21581 }),
  .A3({ S23865 }),
  .ZN({ S23870 })
);
NAND3_X1 #() 
NAND3_X1_4465_ (
  .A1({ S23870 }),
  .A2({ S21512 }),
  .A3({ S23861 }),
  .ZN({ S23871 })
);
AOI21_X1 #() 
AOI21_X1_2233_ (
  .A({ S25957[1224] }),
  .B1({ S23871 }),
  .B2({ S23857 }),
  .ZN({ S23872 })
);
OAI21_X1 #() 
OAI21_X1_2124_ (
  .A({ S25957[1160] }),
  .B1({ S23872 }),
  .B2({ S23845 }),
  .ZN({ S23873 })
);
NAND3_X1 #() 
NAND3_X1_4466_ (
  .A1({ S23871 }),
  .A2({ S23857 }),
  .A3({ S25957[1224] }),
  .ZN({ S23874 })
);
NAND3_X1 #() 
NAND3_X1_4467_ (
  .A1({ S23844 }),
  .A2({ S23822 }),
  .A3({ S21187 }),
  .ZN({ S23875 })
);
NAND3_X1 #() 
NAND3_X1_4468_ (
  .A1({ S23874 }),
  .A2({ S23875 }),
  .A3({ S20144 }),
  .ZN({ S23876 })
);
NAND2_X1 #() 
NAND2_X1_4145_ (
  .A1({ S23873 }),
  .A2({ S23876 }),
  .ZN({ S25957[904] })
);
NOR2_X1 #() 
NOR2_X1_1052_ (
  .A1({ S17241 }),
  .A2({ S17284 }),
  .ZN({ S25957[1193] })
);
NAND2_X1 #() 
NAND2_X1_4146_ (
  .A1({ S21309 }),
  .A2({ S21312 }),
  .ZN({ S25957[1097] })
);
XOR2_X1 #() 
XOR2_X1_74_ (
  .A({ S25957[1097] }),
  .B({ S25957[1193] }),
  .Z({ S25957[1065] })
);
AOI21_X1 #() 
AOI21_X1_2234_ (
  .A({ S80 }),
  .B1({ S23410 }),
  .B2({ S23409 }),
  .ZN({ S23877 })
);
NAND3_X1 #() 
NAND3_X1_4469_ (
  .A1({ S23377 }),
  .A2({ S23577 }),
  .A3({ S25957[1028] }),
  .ZN({ S23878 })
);
NAND3_X1 #() 
NAND3_X1_4470_ (
  .A1({ S23421 }),
  .A2({ S23396 }),
  .A3({ S23427 }),
  .ZN({ S23879 })
);
OAI211_X1 #() 
OAI211_X1_1445_ (
  .A({ S23878 }),
  .B({ S25957[1029] }),
  .C1({ S23877 }),
  .C2({ S23879 }),
  .ZN({ S23880 })
);
NAND2_X1 #() 
NAND2_X1_4147_ (
  .A1({ S23592 }),
  .A2({ S23818 }),
  .ZN({ S23881 })
);
NOR2_X1 #() 
NOR2_X1_1053_ (
  .A1({ S23391 }),
  .A2({ S23360 }),
  .ZN({ S23882 })
);
NAND3_X1 #() 
NAND3_X1_4471_ (
  .A1({ S23387 }),
  .A2({ S25957[1027] }),
  .A3({ S23359 }),
  .ZN({ S23883 })
);
OAI211_X1 #() 
OAI211_X1_1446_ (
  .A({ S23883 }),
  .B({ S23396 }),
  .C1({ S23468 }),
  .C2({ S23882 }),
  .ZN({ S23884 })
);
NAND3_X1 #() 
NAND3_X1_4472_ (
  .A1({ S23881 }),
  .A2({ S23368 }),
  .A3({ S23884 }),
  .ZN({ S23885 })
);
NAND3_X1 #() 
NAND3_X1_4473_ (
  .A1({ S23885 }),
  .A2({ S25957[1030] }),
  .A3({ S23880 }),
  .ZN({ S23886 })
);
NAND3_X1 #() 
NAND3_X1_4474_ (
  .A1({ S23582 }),
  .A2({ S23751 }),
  .A3({ S23396 }),
  .ZN({ S23887 })
);
AOI21_X1 #() 
AOI21_X1_2235_ (
  .A({ S80 }),
  .B1({ S23402 }),
  .B2({ S23401 }),
  .ZN({ S23888 })
);
OAI211_X1 #() 
OAI211_X1_1447_ (
  .A({ S25957[1029] }),
  .B({ S23887 }),
  .C1({ S23888 }),
  .C2({ S23374 }),
  .ZN({ S23889 })
);
NAND2_X1 #() 
NAND2_X1_4148_ (
  .A1({ S23656 }),
  .A2({ S23396 }),
  .ZN({ S23890 })
);
NAND3_X1 #() 
NAND3_X1_4475_ (
  .A1({ S23591 }),
  .A2({ S80 }),
  .A3({ S23370 }),
  .ZN({ S23891 })
);
AOI21_X1 #() 
AOI21_X1_2236_ (
  .A({ S25957[1029] }),
  .B1({ S23491 }),
  .B2({ S23891 }),
  .ZN({ S23892 })
);
OAI21_X1 #() 
OAI21_X1_2125_ (
  .A({ S23892 }),
  .B1({ S23890 }),
  .B2({ S23400 }),
  .ZN({ S23893 })
);
NAND3_X1 #() 
NAND3_X1_4476_ (
  .A1({ S23893 }),
  .A2({ S23889 }),
  .A3({ S21581 }),
  .ZN({ S23894 })
);
NAND3_X1 #() 
NAND3_X1_4477_ (
  .A1({ S23894 }),
  .A2({ S23886 }),
  .A3({ S25957[1031] }),
  .ZN({ S23895 })
);
INV_X1 #() 
INV_X1_1357_ (
  .A({ S23447 }),
  .ZN({ S23896 })
);
NAND4_X1 #() 
NAND4_X1_484_ (
  .A1({ S23398 }),
  .A2({ S23369 }),
  .A3({ S23397 }),
  .A4({ S25957[1027] }),
  .ZN({ S23897 })
);
OAI211_X1 #() 
OAI211_X1_1448_ (
  .A({ S23897 }),
  .B({ S25957[1028] }),
  .C1({ S23896 }),
  .C2({ S23639 }),
  .ZN({ S23898 })
);
OAI211_X1 #() 
OAI211_X1_1449_ (
  .A({ S80 }),
  .B({ S23447 }),
  .C1({ S23391 }),
  .C2({ S25957[1024] }),
  .ZN({ S23899 })
);
NAND3_X1 #() 
NAND3_X1_4478_ (
  .A1({ S23465 }),
  .A2({ S23899 }),
  .A3({ S23396 }),
  .ZN({ S23900 })
);
NAND3_X1 #() 
NAND3_X1_4479_ (
  .A1({ S23898 }),
  .A2({ S23900 }),
  .A3({ S25957[1029] }),
  .ZN({ S23901 })
);
NAND3_X1 #() 
NAND3_X1_4480_ (
  .A1({ S23390 }),
  .A2({ S80 }),
  .A3({ S23467 }),
  .ZN({ S23902 })
);
NAND3_X1 #() 
NAND3_X1_4481_ (
  .A1({ S23823 }),
  .A2({ S25957[1028] }),
  .A3({ S23902 }),
  .ZN({ S23903 })
);
NAND3_X1 #() 
NAND3_X1_4482_ (
  .A1({ S23517 }),
  .A2({ S23396 }),
  .A3({ S23738 }),
  .ZN({ S23904 })
);
NAND3_X1 #() 
NAND3_X1_4483_ (
  .A1({ S23903 }),
  .A2({ S23368 }),
  .A3({ S23904 }),
  .ZN({ S23905 })
);
NAND3_X1 #() 
NAND3_X1_4484_ (
  .A1({ S23905 }),
  .A2({ S25957[1030] }),
  .A3({ S23901 }),
  .ZN({ S23906 })
);
AOI21_X1 #() 
AOI21_X1_2237_ (
  .A({ S23396 }),
  .B1({ S23730 }),
  .B2({ S23641 }),
  .ZN({ S23907 })
);
OAI21_X1 #() 
OAI21_X1_2126_ (
  .A({ S25957[1029] }),
  .B1({ S23907 }),
  .B2({ S23393 }),
  .ZN({ S23908 })
);
NAND2_X1 #() 
NAND2_X1_4149_ (
  .A1({ S23745 }),
  .A2({ S23740 }),
  .ZN({ S23909 })
);
NAND3_X1 #() 
NAND3_X1_4485_ (
  .A1({ S23465 }),
  .A2({ S25957[1028] }),
  .A3({ S23632 }),
  .ZN({ S23910 })
);
NAND3_X1 #() 
NAND3_X1_4486_ (
  .A1({ S23909 }),
  .A2({ S23910 }),
  .A3({ S23368 }),
  .ZN({ S23911 })
);
NAND3_X1 #() 
NAND3_X1_4487_ (
  .A1({ S23908 }),
  .A2({ S23911 }),
  .A3({ S21581 }),
  .ZN({ S23912 })
);
NAND3_X1 #() 
NAND3_X1_4488_ (
  .A1({ S23906 }),
  .A2({ S21512 }),
  .A3({ S23912 }),
  .ZN({ S23913 })
);
NAND3_X1 #() 
NAND3_X1_4489_ (
  .A1({ S23895 }),
  .A2({ S23913 }),
  .A3({ S25957[1225] }),
  .ZN({ S23914 })
);
NAND2_X1 #() 
NAND2_X1_4150_ (
  .A1({ S23895 }),
  .A2({ S23913 }),
  .ZN({ S23915 })
);
NAND2_X1 #() 
NAND2_X1_4151_ (
  .A1({ S23915 }),
  .A2({ S21266 }),
  .ZN({ S23916 })
);
NAND3_X1 #() 
NAND3_X1_4490_ (
  .A1({ S23916 }),
  .A2({ S25957[1065] }),
  .A3({ S23914 }),
  .ZN({ S23917 })
);
INV_X1 #() 
INV_X1_1358_ (
  .A({ S25957[1065] }),
  .ZN({ S23918 })
);
AND3_X1 #() 
AND3_X1_164_ (
  .A1({ S23895 }),
  .A2({ S23913 }),
  .A3({ S25957[1225] }),
  .ZN({ S23919 })
);
AOI21_X1 #() 
AOI21_X1_2238_ (
  .A({ S25957[1225] }),
  .B1({ S23895 }),
  .B2({ S23913 }),
  .ZN({ S23920 })
);
OAI21_X1 #() 
OAI21_X1_2127_ (
  .A({ S23918 }),
  .B1({ S23919 }),
  .B2({ S23920 }),
  .ZN({ S23921 })
);
NAND3_X1 #() 
NAND3_X1_4491_ (
  .A1({ S23921 }),
  .A2({ S23917 }),
  .A3({ S22634 }),
  .ZN({ S23922 })
);
OAI21_X1 #() 
OAI21_X1_2128_ (
  .A({ S25957[1065] }),
  .B1({ S23919 }),
  .B2({ S23920 }),
  .ZN({ S23923 })
);
NAND3_X1 #() 
NAND3_X1_4492_ (
  .A1({ S23916 }),
  .A2({ S23918 }),
  .A3({ S23914 }),
  .ZN({ S23924 })
);
NAND3_X1 #() 
NAND3_X1_4493_ (
  .A1({ S23923 }),
  .A2({ S23924 }),
  .A3({ S25957[1033] }),
  .ZN({ S23925 })
);
NAND2_X1 #() 
NAND2_X1_4152_ (
  .A1({ S23922 }),
  .A2({ S23925 }),
  .ZN({ S25957[905] })
);
NOR2_X1 #() 
NOR2_X1_1054_ (
  .A1({ S21382 }),
  .A2({ S21385 }),
  .ZN({ S25957[1066] })
);
INV_X1 #() 
INV_X1_1359_ (
  .A({ S25957[1066] }),
  .ZN({ S23926 })
);
AOI21_X1 #() 
AOI21_X1_2239_ (
  .A({ S23368 }),
  .B1({ S23428 }),
  .B2({ S23422 }),
  .ZN({ S23927 })
);
NAND4_X1 #() 
NAND4_X1_485_ (
  .A1({ S23455 }),
  .A2({ S23447 }),
  .A3({ S23386 }),
  .A4({ S80 }),
  .ZN({ S23928 })
);
NAND3_X1 #() 
NAND3_X1_4494_ (
  .A1({ S23447 }),
  .A2({ S25957[1027] }),
  .A3({ S25957[1025] }),
  .ZN({ S23929 })
);
AND2_X1 #() 
AND2_X1_260_ (
  .A1({ S23929 }),
  .A2({ S23368 }),
  .ZN({ S23930 })
);
AOI22_X1 #() 
AOI22_X1_476_ (
  .A1({ S23459 }),
  .A2({ S23927 }),
  .B1({ S23930 }),
  .B2({ S23928 }),
  .ZN({ S23931 })
);
OAI211_X1 #() 
OAI211_X1_1450_ (
  .A({ S23369 }),
  .B({ S25957[1027] }),
  .C1({ S25957[1024] }),
  .C2({ S23422 }),
  .ZN({ S23932 })
);
NAND2_X1 #() 
NAND2_X1_4153_ (
  .A1({ S23458 }),
  .A2({ S80 }),
  .ZN({ S23933 })
);
AOI21_X1 #() 
AOI21_X1_2240_ (
  .A({ S25957[1029] }),
  .B1({ S23932 }),
  .B2({ S23933 }),
  .ZN({ S23934 })
);
NAND3_X1 #() 
NAND3_X1_4495_ (
  .A1({ S25957[1029] }),
  .A2({ S23425 }),
  .A3({ S23397 }),
  .ZN({ S23935 })
);
NAND2_X1 #() 
NAND2_X1_4154_ (
  .A1({ S23935 }),
  .A2({ S23747 }),
  .ZN({ S23936 })
);
OAI21_X1 #() 
OAI21_X1_2129_ (
  .A({ S25957[1028] }),
  .B1({ S23934 }),
  .B2({ S23936 }),
  .ZN({ S23937 })
);
OAI211_X1 #() 
OAI211_X1_1451_ (
  .A({ S23937 }),
  .B({ S25957[1030] }),
  .C1({ S23931 }),
  .C2({ S25957[1028] }),
  .ZN({ S23938 })
);
AOI21_X1 #() 
AOI21_X1_2241_ (
  .A({ S23396 }),
  .B1({ S23652 }),
  .B2({ S23929 }),
  .ZN({ S23939 })
);
OAI211_X1 #() 
OAI211_X1_1452_ (
  .A({ S80 }),
  .B({ S23380 }),
  .C1({ S23419 }),
  .C2({ S23492 }),
  .ZN({ S23940 })
);
AOI21_X1 #() 
AOI21_X1_2242_ (
  .A({ S25957[1028] }),
  .B1({ S23540 }),
  .B2({ S23940 }),
  .ZN({ S23941 })
);
OAI21_X1 #() 
OAI21_X1_2130_ (
  .A({ S23368 }),
  .B1({ S23941 }),
  .B2({ S23939 }),
  .ZN({ S23942 })
);
AOI21_X1 #() 
AOI21_X1_2243_ (
  .A({ S23396 }),
  .B1({ S23653 }),
  .B2({ S23467 }),
  .ZN({ S23943 })
);
NAND2_X1 #() 
NAND2_X1_4155_ (
  .A1({ S23943 }),
  .A2({ S23729 }),
  .ZN({ S23944 })
);
NAND3_X1 #() 
NAND3_X1_4496_ (
  .A1({ S23390 }),
  .A2({ S25957[1027] }),
  .A3({ S23419 }),
  .ZN({ S23945 })
);
AOI21_X1 #() 
AOI21_X1_2244_ (
  .A({ S25957[1028] }),
  .B1({ S23499 }),
  .B2({ S23498 }),
  .ZN({ S23946 })
);
AOI21_X1 #() 
AOI21_X1_2245_ (
  .A({ S23368 }),
  .B1({ S23946 }),
  .B2({ S23945 }),
  .ZN({ S23947 })
);
AOI21_X1 #() 
AOI21_X1_2246_ (
  .A({ S25957[1030] }),
  .B1({ S23947 }),
  .B2({ S23944 }),
  .ZN({ S23948 })
);
NAND2_X1 #() 
NAND2_X1_4156_ (
  .A1({ S23942 }),
  .A2({ S23948 }),
  .ZN({ S23949 })
);
NAND3_X1 #() 
NAND3_X1_4497_ (
  .A1({ S23949 }),
  .A2({ S23938 }),
  .A3({ S21512 }),
  .ZN({ S23950 })
);
NAND3_X1 #() 
NAND3_X1_4498_ (
  .A1({ S23804 }),
  .A2({ S25957[1028] }),
  .A3({ S23389 }),
  .ZN({ S23951 })
);
NAND3_X1 #() 
NAND3_X1_4499_ (
  .A1({ S23454 }),
  .A2({ S23667 }),
  .A3({ S25957[1027] }),
  .ZN({ S23952 })
);
NAND3_X1 #() 
NAND3_X1_4500_ (
  .A1({ S23952 }),
  .A2({ S23396 }),
  .A3({ S23421 }),
  .ZN({ S23953 })
);
NAND3_X1 #() 
NAND3_X1_4501_ (
  .A1({ S23951 }),
  .A2({ S23953 }),
  .A3({ S25957[1029] }),
  .ZN({ S23954 })
);
INV_X1 #() 
INV_X1_1360_ (
  .A({ S23954 }),
  .ZN({ S23955 })
);
NAND2_X1 #() 
NAND2_X1_4157_ (
  .A1({ S23425 }),
  .A2({ S25957[1024] }),
  .ZN({ S23956 })
);
NAND3_X1 #() 
NAND3_X1_4502_ (
  .A1({ S23745 }),
  .A2({ S25957[1028] }),
  .A3({ S23956 }),
  .ZN({ S23957 })
);
NAND3_X1 #() 
NAND3_X1_4503_ (
  .A1({ S23398 }),
  .A2({ S25957[1027] }),
  .A3({ S23381 }),
  .ZN({ S23958 })
);
NAND4_X1 #() 
NAND4_X1_486_ (
  .A1({ S23738 }),
  .A2({ S23958 }),
  .A3({ S23493 }),
  .A4({ S23396 }),
  .ZN({ S23959 })
);
NAND3_X1 #() 
NAND3_X1_4504_ (
  .A1({ S23957 }),
  .A2({ S23959 }),
  .A3({ S25957[1029] }),
  .ZN({ S23960 })
);
NAND3_X1 #() 
NAND3_X1_4505_ (
  .A1({ S23500 }),
  .A2({ S23396 }),
  .A3({ S23497 }),
  .ZN({ S23961 })
);
OAI211_X1 #() 
OAI211_X1_1453_ (
  .A({ S23929 }),
  .B({ S25957[1028] }),
  .C1({ S25957[1027] }),
  .C2({ S23490 }),
  .ZN({ S23962 })
);
NAND3_X1 #() 
NAND3_X1_4506_ (
  .A1({ S23961 }),
  .A2({ S23368 }),
  .A3({ S23962 }),
  .ZN({ S23963 })
);
NAND3_X1 #() 
NAND3_X1_4507_ (
  .A1({ S23960 }),
  .A2({ S23963 }),
  .A3({ S21581 }),
  .ZN({ S23964 })
);
NAND3_X1 #() 
NAND3_X1_4508_ (
  .A1({ S23447 }),
  .A2({ S80 }),
  .A3({ S23361 }),
  .ZN({ S23965 })
);
AND2_X1 #() 
AND2_X1_261_ (
  .A1({ S23965 }),
  .A2({ S25957[1028] }),
  .ZN({ S23966 })
);
NAND3_X1 #() 
NAND3_X1_4509_ (
  .A1({ S23454 }),
  .A2({ S25957[1027] }),
  .A3({ S23455 }),
  .ZN({ S23967 })
);
AND2_X1 #() 
AND2_X1_262_ (
  .A1({ S23967 }),
  .A2({ S23966 }),
  .ZN({ S23968 })
);
NAND3_X1 #() 
NAND3_X1_4510_ (
  .A1({ S23423 }),
  .A2({ S23396 }),
  .A3({ S23797 }),
  .ZN({ S23969 })
);
NAND2_X1 #() 
NAND2_X1_4158_ (
  .A1({ S23969 }),
  .A2({ S23368 }),
  .ZN({ S23970 })
);
OAI21_X1 #() 
OAI21_X1_2131_ (
  .A({ S25957[1030] }),
  .B1({ S23968 }),
  .B2({ S23970 }),
  .ZN({ S23971 })
);
OAI211_X1 #() 
OAI211_X1_1454_ (
  .A({ S25957[1031] }),
  .B({ S23964 }),
  .C1({ S23955 }),
  .C2({ S23971 }),
  .ZN({ S23972 })
);
NAND3_X1 #() 
NAND3_X1_4511_ (
  .A1({ S23950 }),
  .A2({ S23972 }),
  .A3({ S25957[1226] }),
  .ZN({ S23973 })
);
NAND2_X1 #() 
NAND2_X1_4159_ (
  .A1({ S23967 }),
  .A2({ S23966 }),
  .ZN({ S23974 })
);
NAND3_X1 #() 
NAND3_X1_4512_ (
  .A1({ S23974 }),
  .A2({ S23368 }),
  .A3({ S23969 }),
  .ZN({ S23975 })
);
NAND2_X1 #() 
NAND2_X1_4160_ (
  .A1({ S23954 }),
  .A2({ S23975 }),
  .ZN({ S23976 })
);
NAND2_X1 #() 
NAND2_X1_4161_ (
  .A1({ S23976 }),
  .A2({ S25957[1030] }),
  .ZN({ S23977 })
);
NAND2_X1 #() 
NAND2_X1_4162_ (
  .A1({ S23960 }),
  .A2({ S23963 }),
  .ZN({ S23978 })
);
NAND2_X1 #() 
NAND2_X1_4163_ (
  .A1({ S23978 }),
  .A2({ S21581 }),
  .ZN({ S23979 })
);
NAND3_X1 #() 
NAND3_X1_4513_ (
  .A1({ S23977 }),
  .A2({ S25957[1031] }),
  .A3({ S23979 }),
  .ZN({ S23980 })
);
NAND2_X1 #() 
NAND2_X1_4164_ (
  .A1({ S23425 }),
  .A2({ S23397 }),
  .ZN({ S23981 })
);
NAND2_X1 #() 
NAND2_X1_4165_ (
  .A1({ S23981 }),
  .A2({ S23747 }),
  .ZN({ S23982 })
);
NAND2_X1 #() 
NAND2_X1_4166_ (
  .A1({ S23982 }),
  .A2({ S25957[1028] }),
  .ZN({ S23983 })
);
AOI21_X1 #() 
AOI21_X1_2247_ (
  .A({ S25957[1028] }),
  .B1({ S23428 }),
  .B2({ S23422 }),
  .ZN({ S23984 })
);
NAND2_X1 #() 
NAND2_X1_4167_ (
  .A1({ S23459 }),
  .A2({ S23984 }),
  .ZN({ S23985 })
);
AOI21_X1 #() 
AOI21_X1_2248_ (
  .A({ S23368 }),
  .B1({ S23985 }),
  .B2({ S23983 }),
  .ZN({ S23986 })
);
AND4_X1 #() 
AND4_X1_10_ (
  .A1({ S25957[1028] }),
  .A2({ S23932 }),
  .A3({ S23933 }),
  .A4({ S23747 }),
  .ZN({ S23987 })
);
NAND2_X1 #() 
NAND2_X1_4168_ (
  .A1({ S23398 }),
  .A2({ S23381 }),
  .ZN({ S23988 })
);
AOI21_X1 #() 
AOI21_X1_2249_ (
  .A({ S25957[1027] }),
  .B1({ S23988 }),
  .B2({ S23455 }),
  .ZN({ S23989 })
);
NAND3_X1 #() 
NAND3_X1_4514_ (
  .A1({ S23398 }),
  .A2({ S25957[1027] }),
  .A3({ S23380 }),
  .ZN({ S23990 })
);
NAND2_X1 #() 
NAND2_X1_4169_ (
  .A1({ S23990 }),
  .A2({ S23396 }),
  .ZN({ S23991 })
);
OAI21_X1 #() 
OAI21_X1_2132_ (
  .A({ S23368 }),
  .B1({ S23989 }),
  .B2({ S23991 }),
  .ZN({ S23992 })
);
NOR2_X1 #() 
NOR2_X1_1055_ (
  .A1({ S23992 }),
  .A2({ S23987 }),
  .ZN({ S23993 })
);
OAI21_X1 #() 
OAI21_X1_2133_ (
  .A({ S25957[1030] }),
  .B1({ S23993 }),
  .B2({ S23986 }),
  .ZN({ S23994 })
);
AOI22_X1 #() 
AOI22_X1_477_ (
  .A1({ S23943 }),
  .A2({ S23729 }),
  .B1({ S23946 }),
  .B2({ S23945 }),
  .ZN({ S23995 })
);
NAND2_X1 #() 
NAND2_X1_4170_ (
  .A1({ S23958 }),
  .A2({ S23646 }),
  .ZN({ S23996 })
);
AOI21_X1 #() 
AOI21_X1_2250_ (
  .A({ S25957[1029] }),
  .B1({ S23996 }),
  .B2({ S23396 }),
  .ZN({ S23997 })
);
AOI22_X1 #() 
AOI22_X1_478_ (
  .A1({ S23421 }),
  .A2({ S23427 }),
  .B1({ S23490 }),
  .B2({ S25957[1024] }),
  .ZN({ S23998 })
);
INV_X1 #() 
INV_X1_1361_ (
  .A({ S23929 }),
  .ZN({ S23999 })
);
OAI21_X1 #() 
OAI21_X1_2134_ (
  .A({ S25957[1028] }),
  .B1({ S23998 }),
  .B2({ S23999 }),
  .ZN({ S24000 })
);
NAND4_X1 #() 
NAND4_X1_487_ (
  .A1({ S23454 }),
  .A2({ S23380 }),
  .A3({ S80 }),
  .A4({ S23396 }),
  .ZN({ S24001 })
);
NAND3_X1 #() 
NAND3_X1_4515_ (
  .A1({ S23997 }),
  .A2({ S24000 }),
  .A3({ S24001 }),
  .ZN({ S24002 })
);
OAI211_X1 #() 
OAI211_X1_1455_ (
  .A({ S24002 }),
  .B({ S21581 }),
  .C1({ S23368 }),
  .C2({ S23995 }),
  .ZN({ S24003 })
);
NAND3_X1 #() 
NAND3_X1_4516_ (
  .A1({ S23994 }),
  .A2({ S24003 }),
  .A3({ S21512 }),
  .ZN({ S24004 })
);
NAND3_X1 #() 
NAND3_X1_4517_ (
  .A1({ S23980 }),
  .A2({ S22637 }),
  .A3({ S24004 }),
  .ZN({ S24005 })
);
NAND3_X1 #() 
NAND3_X1_4518_ (
  .A1({ S24005 }),
  .A2({ S23926 }),
  .A3({ S23973 }),
  .ZN({ S24006 })
);
AND3_X1 #() 
AND3_X1_165_ (
  .A1({ S23950 }),
  .A2({ S23972 }),
  .A3({ S25957[1226] }),
  .ZN({ S24007 })
);
AOI21_X1 #() 
AOI21_X1_2251_ (
  .A({ S25957[1226] }),
  .B1({ S23950 }),
  .B2({ S23972 }),
  .ZN({ S24008 })
);
OAI21_X1 #() 
OAI21_X1_2135_ (
  .A({ S25957[1066] }),
  .B1({ S24007 }),
  .B2({ S24008 }),
  .ZN({ S24009 })
);
NAND3_X1 #() 
NAND3_X1_4519_ (
  .A1({ S24009 }),
  .A2({ S24006 }),
  .A3({ S25957[1034] }),
  .ZN({ S24010 })
);
OAI21_X1 #() 
OAI21_X1_2136_ (
  .A({ S23926 }),
  .B1({ S24007 }),
  .B2({ S24008 }),
  .ZN({ S24011 })
);
NAND3_X1 #() 
NAND3_X1_4520_ (
  .A1({ S24005 }),
  .A2({ S25957[1066] }),
  .A3({ S23973 }),
  .ZN({ S24012 })
);
NAND3_X1 #() 
NAND3_X1_4521_ (
  .A1({ S24011 }),
  .A2({ S24012 }),
  .A3({ S22644 }),
  .ZN({ S24013 })
);
NAND2_X1 #() 
NAND2_X1_4171_ (
  .A1({ S24010 }),
  .A2({ S24013 }),
  .ZN({ S25957[906] })
);
NAND3_X1 #() 
NAND3_X1_4522_ (
  .A1({ S22562 }),
  .A2({ S25957[1241] }),
  .A3({ S22560 }),
  .ZN({ S24014 })
);
INV_X1 #() 
INV_X1_1362_ (
  .A({ S25957[1241] }),
  .ZN({ S24015 })
);
NAND3_X1 #() 
NAND3_X1_4523_ (
  .A1({ S22565 }),
  .A2({ S24015 }),
  .A3({ S22564 }),
  .ZN({ S24016 })
);
NAND3_X1 #() 
NAND3_X1_4524_ (
  .A1({ S24014 }),
  .A2({ S24016 }),
  .A3({ S25956[25] }),
  .ZN({ S24017 })
);
NAND3_X1 #() 
NAND3_X1_4525_ (
  .A1({ S22562 }),
  .A2({ S24015 }),
  .A3({ S22560 }),
  .ZN({ S24018 })
);
NAND3_X1 #() 
NAND3_X1_4526_ (
  .A1({ S22565 }),
  .A2({ S25957[1241] }),
  .A3({ S22564 }),
  .ZN({ S24019 })
);
NAND3_X1 #() 
NAND3_X1_4527_ (
  .A1({ S24018 }),
  .A2({ S24019 }),
  .A3({ S18383 }),
  .ZN({ S24020 })
);
AND4_X1 #() 
AND4_X1_11_ (
  .A1({ S22518 }),
  .A2({ S24017 }),
  .A3({ S24020 }),
  .A4({ S22521 }),
  .ZN({ S90 })
);
NAND2_X1 #() 
NAND2_X1_4172_ (
  .A1({ S22518 }),
  .A2({ S22521 }),
  .ZN({ S24021 })
);
NAND2_X1 #() 
NAND2_X1_4173_ (
  .A1({ S24017 }),
  .A2({ S24020 }),
  .ZN({ S24022 })
);
NAND2_X1 #() 
NAND2_X1_4174_ (
  .A1({ S24022 }),
  .A2({ S24021 }),
  .ZN({ S91 })
);
INV_X1 #() 
INV_X1_1363_ (
  .A({ S25957[1191] }),
  .ZN({ S24023 })
);
NAND3_X1 #() 
NAND3_X1_4528_ (
  .A1({ S22621 }),
  .A2({ S22627 }),
  .A3({ S25957[1048] }),
  .ZN({ S24024 })
);
NAND4_X1 #() 
NAND4_X1_488_ (
  .A1({ S22567 }),
  .A2({ S22570 }),
  .A3({ S22518 }),
  .A4({ S22521 }),
  .ZN({ S24025 })
);
NAND3_X1 #() 
NAND3_X1_4529_ (
  .A1({ S24021 }),
  .A2({ S24017 }),
  .A3({ S24020 }),
  .ZN({ S24026 })
);
NAND2_X1 #() 
NAND2_X1_4175_ (
  .A1({ S24026 }),
  .A2({ S24025 }),
  .ZN({ S24027 })
);
AOI21_X1 #() 
AOI21_X1_2252_ (
  .A({ S25957[1051] }),
  .B1({ S24027 }),
  .B2({ S25957[1050] }),
  .ZN({ S24028 })
);
NAND2_X1 #() 
NAND2_X1_4176_ (
  .A1({ S24028 }),
  .A2({ S24024 }),
  .ZN({ S24029 })
);
AOI21_X1 #() 
AOI21_X1_2253_ (
  .A({ S21411 }),
  .B1({ S22625 }),
  .B2({ S22626 }),
  .ZN({ S24030 })
);
NOR3_X1 #() 
NOR3_X1_143_ (
  .A1({ S22620 }),
  .A2({ S22619 }),
  .A3({ S25957[1178] }),
  .ZN({ S24031 })
);
NAND4_X1 #() 
NAND4_X1_489_ (
  .A1({ S24017 }),
  .A2({ S24020 }),
  .A3({ S22518 }),
  .A4({ S22521 }),
  .ZN({ S24032 })
);
OAI21_X1 #() 
OAI21_X1_2137_ (
  .A({ S24032 }),
  .B1({ S24031 }),
  .B2({ S24030 }),
  .ZN({ S24033 })
);
NAND4_X1 #() 
NAND4_X1_490_ (
  .A1({ S24026 }),
  .A2({ S22621 }),
  .A3({ S24025 }),
  .A4({ S22627 }),
  .ZN({ S24034 })
);
AOI21_X1 #() 
AOI21_X1_2254_ (
  .A({ S83 }),
  .B1({ S24033 }),
  .B2({ S24034 }),
  .ZN({ S24035 })
);
INV_X1 #() 
INV_X1_1364_ (
  .A({ S24035 }),
  .ZN({ S24036 })
);
NAND3_X1 #() 
NAND3_X1_4530_ (
  .A1({ S24036 }),
  .A2({ S25957[1052] }),
  .A3({ S24029 }),
  .ZN({ S24037 })
);
NAND2_X1 #() 
NAND2_X1_4177_ (
  .A1({ S25957[1050] }),
  .A2({ S25957[1048] }),
  .ZN({ S24038 })
);
NAND3_X1 #() 
NAND3_X1_4531_ (
  .A1({ S22621 }),
  .A2({ S22627 }),
  .A3({ S25957[1049] }),
  .ZN({ S24039 })
);
NAND3_X1 #() 
NAND3_X1_4532_ (
  .A1({ S24038 }),
  .A2({ S25957[1051] }),
  .A3({ S24039 }),
  .ZN({ S24040 })
);
NAND3_X1 #() 
NAND3_X1_4533_ (
  .A1({ S22621 }),
  .A2({ S24025 }),
  .A3({ S22627 }),
  .ZN({ S24041 })
);
NAND2_X1 #() 
NAND2_X1_4178_ (
  .A1({ S24033 }),
  .A2({ S24041 }),
  .ZN({ S24042 })
);
AOI21_X1 #() 
AOI21_X1_2255_ (
  .A({ S25957[1052] }),
  .B1({ S24042 }),
  .B2({ S83 }),
  .ZN({ S24043 })
);
NAND2_X1 #() 
NAND2_X1_4179_ (
  .A1({ S24043 }),
  .A2({ S24040 }),
  .ZN({ S24044 })
);
NAND3_X1 #() 
NAND3_X1_4534_ (
  .A1({ S24037 }),
  .A2({ S24044 }),
  .A3({ S22294 }),
  .ZN({ S24045 })
);
NAND2_X1 #() 
NAND2_X1_4180_ (
  .A1({ S22357 }),
  .A2({ S22360 }),
  .ZN({ S24046 })
);
NAND3_X1 #() 
NAND3_X1_4535_ (
  .A1({ S90 }),
  .A2({ S22621 }),
  .A3({ S22627 }),
  .ZN({ S24047 })
);
AND2_X1 #() 
AND2_X1_263_ (
  .A1({ S24022 }),
  .A2({ S24021 }),
  .ZN({ S24048 })
);
OAI21_X1 #() 
OAI21_X1_2138_ (
  .A({ S24048 }),
  .B1({ S24031 }),
  .B2({ S24030 }),
  .ZN({ S24049 })
);
NAND3_X1 #() 
NAND3_X1_4536_ (
  .A1({ S24049 }),
  .A2({ S25957[1051] }),
  .A3({ S24047 }),
  .ZN({ S24050 })
);
NAND3_X1 #() 
NAND3_X1_4537_ (
  .A1({ S22621 }),
  .A2({ S22627 }),
  .A3({ S24021 }),
  .ZN({ S24051 })
);
NOR2_X1 #() 
NOR2_X1_1056_ (
  .A1({ S25957[1048] }),
  .A2({ S24022 }),
  .ZN({ S24052 })
);
OAI21_X1 #() 
OAI21_X1_2139_ (
  .A({ S24052 }),
  .B1({ S24031 }),
  .B2({ S24030 }),
  .ZN({ S24053 })
);
NAND3_X1 #() 
NAND3_X1_4538_ (
  .A1({ S24053 }),
  .A2({ S83 }),
  .A3({ S24051 }),
  .ZN({ S24054 })
);
AND2_X1 #() 
AND2_X1_264_ (
  .A1({ S24054 }),
  .A2({ S24050 }),
  .ZN({ S24055 })
);
AOI22_X1 #() 
AOI22_X1_479_ (
  .A1({ S22621 }),
  .A2({ S22627 }),
  .B1({ S25957[1049] }),
  .B2({ S25957[1048] }),
  .ZN({ S24056 })
);
NOR2_X1 #() 
NOR2_X1_1057_ (
  .A1({ S24056 }),
  .A2({ S25957[1051] }),
  .ZN({ S24057 })
);
NAND2_X1 #() 
NAND2_X1_4181_ (
  .A1({ S25957[1050] }),
  .A2({ S24022 }),
  .ZN({ S24058 })
);
NAND2_X1 #() 
NAND2_X1_4182_ (
  .A1({ S24058 }),
  .A2({ S24041 }),
  .ZN({ S24059 })
);
NOR2_X1 #() 
NOR2_X1_1058_ (
  .A1({ S24059 }),
  .A2({ S83 }),
  .ZN({ S24060 })
);
OAI21_X1 #() 
OAI21_X1_2140_ (
  .A({ S24046 }),
  .B1({ S24060 }),
  .B2({ S24057 }),
  .ZN({ S24061 })
);
OAI211_X1 #() 
OAI211_X1_1456_ (
  .A({ S24061 }),
  .B({ S25957[1053] }),
  .C1({ S24046 }),
  .C2({ S24055 }),
  .ZN({ S24062 })
);
AOI21_X1 #() 
AOI21_X1_2256_ (
  .A({ S22219 }),
  .B1({ S24062 }),
  .B2({ S24045 }),
  .ZN({ S24063 })
);
NAND2_X1 #() 
NAND2_X1_4183_ (
  .A1({ S91 }),
  .A2({ S24032 }),
  .ZN({ S24064 })
);
NAND2_X1 #() 
NAND2_X1_4184_ (
  .A1({ S25957[1050] }),
  .A2({ S24064 }),
  .ZN({ S24065 })
);
NOR2_X1 #() 
NOR2_X1_1059_ (
  .A1({ S24065 }),
  .A2({ S25957[1051] }),
  .ZN({ S24066 })
);
OAI21_X1 #() 
OAI21_X1_2141_ (
  .A({ S24046 }),
  .B1({ S24033 }),
  .B2({ S83 }),
  .ZN({ S24067 })
);
NAND2_X1 #() 
NAND2_X1_4185_ (
  .A1({ S24028 }),
  .A2({ S24047 }),
  .ZN({ S24068 })
);
INV_X1 #() 
INV_X1_1365_ (
  .A({ S24068 }),
  .ZN({ S24069 })
);
AOI21_X1 #() 
AOI21_X1_2257_ (
  .A({ S24026 }),
  .B1({ S22627 }),
  .B2({ S22621 }),
  .ZN({ S24070 })
);
OAI21_X1 #() 
OAI21_X1_2142_ (
  .A({ S25957[1052] }),
  .B1({ S24070 }),
  .B2({ S83 }),
  .ZN({ S24071 })
);
OAI22_X1 #() 
OAI22_X1_108_ (
  .A1({ S24069 }),
  .A2({ S24071 }),
  .B1({ S24067 }),
  .B2({ S24066 }),
  .ZN({ S24072 })
);
NAND2_X1 #() 
NAND2_X1_4186_ (
  .A1({ S24072 }),
  .A2({ S22294 }),
  .ZN({ S24073 })
);
NAND3_X1 #() 
NAND3_X1_4539_ (
  .A1({ S22621 }),
  .A2({ S22627 }),
  .A3({ S24022 }),
  .ZN({ S24074 })
);
AOI21_X1 #() 
AOI21_X1_2258_ (
  .A({ S24021 }),
  .B1({ S22621 }),
  .B2({ S22627 }),
  .ZN({ S24075 })
);
NOR2_X1 #() 
NOR2_X1_1060_ (
  .A1({ S24075 }),
  .A2({ S83 }),
  .ZN({ S24076 })
);
AOI21_X1 #() 
AOI21_X1_2259_ (
  .A({ S24021 }),
  .B1({ S22437 }),
  .B2({ S22434 }),
  .ZN({ S24077 })
);
AOI21_X1 #() 
AOI21_X1_2260_ (
  .A({ S24077 }),
  .B1({ S24076 }),
  .B2({ S24074 }),
  .ZN({ S24078 })
);
AOI21_X1 #() 
AOI21_X1_2261_ (
  .A({ S25957[1051] }),
  .B1({ S24058 }),
  .B2({ S24047 }),
  .ZN({ S24079 })
);
NAND3_X1 #() 
NAND3_X1_4540_ (
  .A1({ S24039 }),
  .A2({ S25957[1051] }),
  .A3({ S24025 }),
  .ZN({ S24080 })
);
NAND2_X1 #() 
NAND2_X1_4187_ (
  .A1({ S24080 }),
  .A2({ S24046 }),
  .ZN({ S24081 })
);
OAI221_X1 #() 
OAI221_X1_118_ (
  .A({ S25957[1053] }),
  .B1({ S24081 }),
  .B2({ S24079 }),
  .C1({ S24078 }),
  .C2({ S24046 }),
  .ZN({ S24082 })
);
AOI21_X1 #() 
AOI21_X1_2262_ (
  .A({ S25957[1054] }),
  .B1({ S24073 }),
  .B2({ S24082 }),
  .ZN({ S24083 })
);
OAI21_X1 #() 
OAI21_X1_2143_ (
  .A({ S22150 }),
  .B1({ S24063 }),
  .B2({ S24083 }),
  .ZN({ S24084 })
);
NAND2_X1 #() 
NAND2_X1_4188_ (
  .A1({ S83 }),
  .A2({ S25957[1049] }),
  .ZN({ S24085 })
);
NOR2_X1 #() 
NOR2_X1_1061_ (
  .A1({ S24075 }),
  .A2({ S24085 }),
  .ZN({ S24086 })
);
NOR2_X1 #() 
NOR2_X1_1062_ (
  .A1({ S83 }),
  .A2({ S25957[1049] }),
  .ZN({ S24087 })
);
AOI21_X1 #() 
AOI21_X1_2263_ (
  .A({ S24087 }),
  .B1({ S24075 }),
  .B2({ S25957[1051] }),
  .ZN({ S24088 })
);
NAND2_X1 #() 
NAND2_X1_4189_ (
  .A1({ S24088 }),
  .A2({ S25957[1052] }),
  .ZN({ S24089 })
);
NAND3_X1 #() 
NAND3_X1_4541_ (
  .A1({ S24048 }),
  .A2({ S22621 }),
  .A3({ S22627 }),
  .ZN({ S24090 })
);
INV_X1 #() 
INV_X1_1366_ (
  .A({ S24090 }),
  .ZN({ S24091 })
);
NOR2_X1 #() 
NOR2_X1_1063_ (
  .A1({ S90 }),
  .A2({ S83 }),
  .ZN({ S24092 })
);
OAI21_X1 #() 
OAI21_X1_2144_ (
  .A({ S24046 }),
  .B1({ S24091 }),
  .B2({ S24092 }),
  .ZN({ S24093 })
);
OAI211_X1 #() 
OAI211_X1_1457_ (
  .A({ S24093 }),
  .B({ S25957[1053] }),
  .C1({ S24089 }),
  .C2({ S24086 }),
  .ZN({ S24094 })
);
AOI21_X1 #() 
AOI21_X1_2264_ (
  .A({ S24022 }),
  .B1({ S22621 }),
  .B2({ S22627 }),
  .ZN({ S24095 })
);
AOI22_X1 #() 
AOI22_X1_480_ (
  .A1({ S24026 }),
  .A2({ S24025 }),
  .B1({ S22621 }),
  .B2({ S22627 }),
  .ZN({ S24096 })
);
INV_X1 #() 
INV_X1_1367_ (
  .A({ S24034 }),
  .ZN({ S24097 })
);
OAI21_X1 #() 
OAI21_X1_2145_ (
  .A({ S25957[1051] }),
  .B1({ S24097 }),
  .B2({ S24096 }),
  .ZN({ S24098 })
);
NAND2_X1 #() 
NAND2_X1_4190_ (
  .A1({ S24024 }),
  .A2({ S83 }),
  .ZN({ S24099 })
);
OAI21_X1 #() 
OAI21_X1_2146_ (
  .A({ S24098 }),
  .B1({ S24095 }),
  .B2({ S24099 }),
  .ZN({ S24100 })
);
NAND2_X1 #() 
NAND2_X1_4191_ (
  .A1({ S24074 }),
  .A2({ S25957[1051] }),
  .ZN({ S24101 })
);
NAND4_X1 #() 
NAND4_X1_491_ (
  .A1({ S22621 }),
  .A2({ S91 }),
  .A3({ S22627 }),
  .A4({ S24032 }),
  .ZN({ S24102 })
);
INV_X1 #() 
INV_X1_1368_ (
  .A({ S24102 }),
  .ZN({ S24103 })
);
AOI22_X1 #() 
AOI22_X1_481_ (
  .A1({ S22621 }),
  .A2({ S22627 }),
  .B1({ S24022 }),
  .B2({ S25957[1048] }),
  .ZN({ S24104 })
);
OAI21_X1 #() 
OAI21_X1_2147_ (
  .A({ S83 }),
  .B1({ S24103 }),
  .B2({ S24104 }),
  .ZN({ S24105 })
);
NAND3_X1 #() 
NAND3_X1_4542_ (
  .A1({ S24105 }),
  .A2({ S24046 }),
  .A3({ S24101 }),
  .ZN({ S24106 })
);
OAI211_X1 #() 
OAI211_X1_1458_ (
  .A({ S22294 }),
  .B({ S24106 }),
  .C1({ S24100 }),
  .C2({ S24046 }),
  .ZN({ S24107 })
);
AOI21_X1 #() 
AOI21_X1_2265_ (
  .A({ S25957[1054] }),
  .B1({ S24107 }),
  .B2({ S24094 }),
  .ZN({ S24108 })
);
NAND3_X1 #() 
NAND3_X1_4543_ (
  .A1({ S22621 }),
  .A2({ S91 }),
  .A3({ S22627 }),
  .ZN({ S24109 })
);
NOR2_X1 #() 
NOR2_X1_1064_ (
  .A1({ S24025 }),
  .A2({ S83 }),
  .ZN({ S24110 })
);
AOI21_X1 #() 
AOI21_X1_2266_ (
  .A({ S24110 }),
  .B1({ S24049 }),
  .B2({ S24109 }),
  .ZN({ S24111 })
);
NAND2_X1 #() 
NAND2_X1_4192_ (
  .A1({ S24026 }),
  .A2({ S83 }),
  .ZN({ S24112 })
);
NAND2_X1 #() 
NAND2_X1_4193_ (
  .A1({ S24058 }),
  .A2({ S25957[1051] }),
  .ZN({ S24113 })
);
NOR2_X1 #() 
NOR2_X1_1065_ (
  .A1({ S24113 }),
  .A2({ S90 }),
  .ZN({ S24114 })
);
INV_X1 #() 
INV_X1_1369_ (
  .A({ S24114 }),
  .ZN({ S24115 })
);
NAND3_X1 #() 
NAND3_X1_4544_ (
  .A1({ S24115 }),
  .A2({ S25957[1052] }),
  .A3({ S24112 }),
  .ZN({ S24116 })
);
OAI211_X1 #() 
OAI211_X1_1459_ (
  .A({ S24116 }),
  .B({ S22294 }),
  .C1({ S25957[1052] }),
  .C2({ S24111 }),
  .ZN({ S24117 })
);
NAND2_X1 #() 
NAND2_X1_4194_ (
  .A1({ S24051 }),
  .A2({ S91 }),
  .ZN({ S24118 })
);
INV_X1 #() 
INV_X1_1370_ (
  .A({ S24118 }),
  .ZN({ S24119 })
);
NAND2_X1 #() 
NAND2_X1_4195_ (
  .A1({ S24038 }),
  .A2({ S24074 }),
  .ZN({ S24120 })
);
OAI21_X1 #() 
OAI21_X1_2148_ (
  .A({ S24046 }),
  .B1({ S24120 }),
  .B2({ S24112 }),
  .ZN({ S24121 })
);
AOI21_X1 #() 
AOI21_X1_2267_ (
  .A({ S24121 }),
  .B1({ S24119 }),
  .B2({ S24092 }),
  .ZN({ S24122 })
);
NAND4_X1 #() 
NAND4_X1_492_ (
  .A1({ S25957[1051] }),
  .A2({ S22621 }),
  .A3({ S24025 }),
  .A4({ S22627 }),
  .ZN({ S24123 })
);
NAND2_X1 #() 
NAND2_X1_4196_ (
  .A1({ S24123 }),
  .A2({ S25957[1052] }),
  .ZN({ S24124 })
);
NAND3_X1 #() 
NAND3_X1_4545_ (
  .A1({ S25957[1050] }),
  .A2({ S25957[1051] }),
  .A3({ S25957[1048] }),
  .ZN({ S24125 })
);
NAND3_X1 #() 
NAND3_X1_4546_ (
  .A1({ S24051 }),
  .A2({ S83 }),
  .A3({ S25957[1049] }),
  .ZN({ S24126 })
);
NAND2_X1 #() 
NAND2_X1_4197_ (
  .A1({ S24126 }),
  .A2({ S24125 }),
  .ZN({ S24127 })
);
OAI21_X1 #() 
OAI21_X1_2149_ (
  .A({ S25957[1053] }),
  .B1({ S24127 }),
  .B2({ S24124 }),
  .ZN({ S24128 })
);
OAI21_X1 #() 
OAI21_X1_2150_ (
  .A({ S24117 }),
  .B1({ S24128 }),
  .B2({ S24122 }),
  .ZN({ S24129 })
);
AOI21_X1 #() 
AOI21_X1_2268_ (
  .A({ S24108 }),
  .B1({ S24129 }),
  .B2({ S25957[1054] }),
  .ZN({ S24130 })
);
OAI21_X1 #() 
OAI21_X1_2151_ (
  .A({ S24084 }),
  .B1({ S24130 }),
  .B2({ S22150 }),
  .ZN({ S24131 })
);
XNOR2_X1 #() 
XNOR2_X1_173_ (
  .A({ S24131 }),
  .B({ S25957[1127] }),
  .ZN({ S25957[999] })
);
NAND2_X1 #() 
NAND2_X1_4198_ (
  .A1({ S25957[999] }),
  .A2({ S24023 }),
  .ZN({ S24132 })
);
NOR2_X1 #() 
NOR2_X1_1066_ (
  .A1({ S25957[999] }),
  .A2({ S24023 }),
  .ZN({ S24133 })
);
INV_X1 #() 
INV_X1_1371_ (
  .A({ S24133 }),
  .ZN({ S24134 })
);
NAND3_X1 #() 
NAND3_X1_4547_ (
  .A1({ S24134 }),
  .A2({ S21512 }),
  .A3({ S24132 }),
  .ZN({ S24135 })
);
NAND2_X1 #() 
NAND2_X1_4199_ (
  .A1({ S24134 }),
  .A2({ S24132 }),
  .ZN({ S25957[935] })
);
NAND2_X1 #() 
NAND2_X1_4200_ (
  .A1({ S25957[935] }),
  .A2({ S25957[1031] }),
  .ZN({ S24136 })
);
NAND2_X1 #() 
NAND2_X1_4201_ (
  .A1({ S24136 }),
  .A2({ S24135 }),
  .ZN({ S24137 })
);
INV_X1 #() 
INV_X1_1372_ (
  .A({ S24137 }),
  .ZN({ S25957[903] })
);
XOR2_X1 #() 
XOR2_X1_75_ (
  .A({ S25957[1094] }),
  .B({ S25957[1190] }),
  .Z({ S25957[1062] })
);
NAND2_X1 #() 
NAND2_X1_4202_ (
  .A1({ S25957[1050] }),
  .A2({ S24077 }),
  .ZN({ S24138 })
);
OAI21_X1 #() 
OAI21_X1_2152_ (
  .A({ S24138 }),
  .B1({ S24102 }),
  .B2({ S25957[1051] }),
  .ZN({ S24139 })
);
NAND2_X1 #() 
NAND2_X1_4203_ (
  .A1({ S25957[1050] }),
  .A2({ S24025 }),
  .ZN({ S24140 })
);
NAND2_X1 #() 
NAND2_X1_4204_ (
  .A1({ S24140 }),
  .A2({ S24024 }),
  .ZN({ S24141 })
);
NAND2_X1 #() 
NAND2_X1_4205_ (
  .A1({ S24141 }),
  .A2({ S25957[1051] }),
  .ZN({ S24142 })
);
NAND2_X1 #() 
NAND2_X1_4206_ (
  .A1({ S24142 }),
  .A2({ S25957[1052] }),
  .ZN({ S24143 })
);
AND3_X1 #() 
AND3_X1_166_ (
  .A1({ S22621 }),
  .A2({ S24025 }),
  .A3({ S22627 }),
  .ZN({ S24144 })
);
OAI21_X1 #() 
OAI21_X1_2153_ (
  .A({ S83 }),
  .B1({ S24144 }),
  .B2({ S24056 }),
  .ZN({ S24145 })
);
NAND2_X1 #() 
NAND2_X1_4207_ (
  .A1({ S25957[1050] }),
  .A2({ S91 }),
  .ZN({ S24146 })
);
AND2_X1 #() 
AND2_X1_265_ (
  .A1({ S24146 }),
  .A2({ S24047 }),
  .ZN({ S24147 })
);
OAI21_X1 #() 
OAI21_X1_2154_ (
  .A({ S24145 }),
  .B1({ S24147 }),
  .B2({ S83 }),
  .ZN({ S24148 })
);
OAI22_X1 #() 
OAI22_X1_109_ (
  .A1({ S24148 }),
  .A2({ S25957[1052] }),
  .B1({ S24143 }),
  .B2({ S24139 }),
  .ZN({ S24149 })
);
NAND3_X1 #() 
NAND3_X1_4548_ (
  .A1({ S24140 }),
  .A2({ S25957[1051] }),
  .A3({ S24109 }),
  .ZN({ S24150 })
);
NAND3_X1 #() 
NAND3_X1_4549_ (
  .A1({ S25957[1050] }),
  .A2({ S83 }),
  .A3({ S91 }),
  .ZN({ S24151 })
);
NAND3_X1 #() 
NAND3_X1_4550_ (
  .A1({ S24150 }),
  .A2({ S25957[1052] }),
  .A3({ S24151 }),
  .ZN({ S24152 })
);
NAND2_X1 #() 
NAND2_X1_4208_ (
  .A1({ S24115 }),
  .A2({ S24085 }),
  .ZN({ S24153 })
);
AOI21_X1 #() 
AOI21_X1_2269_ (
  .A({ S22294 }),
  .B1({ S24153 }),
  .B2({ S24046 }),
  .ZN({ S24154 })
);
AOI22_X1 #() 
AOI22_X1_482_ (
  .A1({ S24154 }),
  .A2({ S24152 }),
  .B1({ S24149 }),
  .B2({ S22294 }),
  .ZN({ S24155 })
);
AOI21_X1 #() 
AOI21_X1_2270_ (
  .A({ S83 }),
  .B1({ S24053 }),
  .B2({ S24024 }),
  .ZN({ S24156 })
);
OAI21_X1 #() 
OAI21_X1_2155_ (
  .A({ S24046 }),
  .B1({ S24139 }),
  .B2({ S24156 }),
  .ZN({ S24157 })
);
OAI211_X1 #() 
OAI211_X1_1460_ (
  .A({ S24088 }),
  .B({ S25957[1052] }),
  .C1({ S25957[1051] }),
  .C2({ S24041 }),
  .ZN({ S24158 })
);
NAND3_X1 #() 
NAND3_X1_4551_ (
  .A1({ S24157 }),
  .A2({ S22294 }),
  .A3({ S24158 }),
  .ZN({ S24159 })
);
AND3_X1 #() 
AND3_X1_167_ (
  .A1({ S24026 }),
  .A2({ S22621 }),
  .A3({ S22627 }),
  .ZN({ S24160 })
);
AOI21_X1 #() 
AOI21_X1_2271_ (
  .A({ S25957[1052] }),
  .B1({ S24160 }),
  .B2({ S25957[1051] }),
  .ZN({ S24161 })
);
NAND2_X1 #() 
NAND2_X1_4209_ (
  .A1({ S24024 }),
  .A2({ S24064 }),
  .ZN({ S24162 })
);
NAND2_X1 #() 
NAND2_X1_4210_ (
  .A1({ S24095 }),
  .A2({ S25957[1051] }),
  .ZN({ S24163 })
);
OAI211_X1 #() 
OAI211_X1_1461_ (
  .A({ S24161 }),
  .B({ S24163 }),
  .C1({ S25957[1051] }),
  .C2({ S24162 }),
  .ZN({ S24164 })
);
OAI21_X1 #() 
OAI21_X1_2156_ (
  .A({ S25957[1049] }),
  .B1({ S24031 }),
  .B2({ S24030 }),
  .ZN({ S24165 })
);
NOR2_X1 #() 
NOR2_X1_1067_ (
  .A1({ S24165 }),
  .A2({ S83 }),
  .ZN({ S24166 })
);
NOR2_X1 #() 
NOR2_X1_1068_ (
  .A1({ S24051 }),
  .A2({ S24085 }),
  .ZN({ S24167 })
);
NOR2_X1 #() 
NOR2_X1_1069_ (
  .A1({ S24166 }),
  .A2({ S24167 }),
  .ZN({ S24168 })
);
INV_X1 #() 
INV_X1_1373_ (
  .A({ S24168 }),
  .ZN({ S24169 })
);
OAI21_X1 #() 
OAI21_X1_2157_ (
  .A({ S25957[1052] }),
  .B1({ S24169 }),
  .B2({ S24066 }),
  .ZN({ S24170 })
);
NAND3_X1 #() 
NAND3_X1_4552_ (
  .A1({ S24170 }),
  .A2({ S25957[1053] }),
  .A3({ S24164 }),
  .ZN({ S24171 })
);
NAND2_X1 #() 
NAND2_X1_4211_ (
  .A1({ S24171 }),
  .A2({ S24159 }),
  .ZN({ S24172 })
);
AOI21_X1 #() 
AOI21_X1_2272_ (
  .A({ S22150 }),
  .B1({ S24172 }),
  .B2({ S22219 }),
  .ZN({ S24173 })
);
OAI21_X1 #() 
OAI21_X1_2158_ (
  .A({ S24173 }),
  .B1({ S22219 }),
  .B2({ S24155 }),
  .ZN({ S24174 })
);
NAND2_X1 #() 
NAND2_X1_4212_ (
  .A1({ S24024 }),
  .A2({ S25957[1051] }),
  .ZN({ S24175 })
);
NOR2_X1 #() 
NOR2_X1_1070_ (
  .A1({ S24175 }),
  .A2({ S24048 }),
  .ZN({ S24176 })
);
AOI21_X1 #() 
AOI21_X1_2273_ (
  .A({ S24176 }),
  .B1({ S24057 }),
  .B2({ S24024 }),
  .ZN({ S24177 })
);
NAND3_X1 #() 
NAND3_X1_4553_ (
  .A1({ S24024 }),
  .A2({ S83 }),
  .A3({ S25957[1049] }),
  .ZN({ S24178 })
);
NAND2_X1 #() 
NAND2_X1_4213_ (
  .A1({ S24178 }),
  .A2({ S24046 }),
  .ZN({ S24179 })
);
OAI221_X1 #() 
OAI221_X1_119_ (
  .A({ S25957[1053] }),
  .B1({ S24179 }),
  .B2({ S24176 }),
  .C1({ S24177 }),
  .C2({ S24046 }),
  .ZN({ S24180 })
);
NAND3_X1 #() 
NAND3_X1_4554_ (
  .A1({ S24074 }),
  .A2({ S83 }),
  .A3({ S24021 }),
  .ZN({ S24181 })
);
NAND4_X1 #() 
NAND4_X1_493_ (
  .A1({ S22621 }),
  .A2({ S25957[1051] }),
  .A3({ S22627 }),
  .A4({ S25957[1049] }),
  .ZN({ S24182 })
);
AND2_X1 #() 
AND2_X1_266_ (
  .A1({ S24182 }),
  .A2({ S25957[1052] }),
  .ZN({ S24183 })
);
AOI21_X1 #() 
AOI21_X1_2274_ (
  .A({ S83 }),
  .B1({ S24140 }),
  .B2({ S24024 }),
  .ZN({ S24184 })
);
NOR3_X1 #() 
NOR3_X1_144_ (
  .A1({ S24184 }),
  .A2({ S24028 }),
  .A3({ S25957[1052] }),
  .ZN({ S24185 })
);
AOI21_X1 #() 
AOI21_X1_2275_ (
  .A({ S24185 }),
  .B1({ S24183 }),
  .B2({ S24181 }),
  .ZN({ S24186 })
);
NAND2_X1 #() 
NAND2_X1_4214_ (
  .A1({ S24186 }),
  .A2({ S22294 }),
  .ZN({ S24187 })
);
AOI21_X1 #() 
AOI21_X1_2276_ (
  .A({ S22219 }),
  .B1({ S24187 }),
  .B2({ S24180 }),
  .ZN({ S24188 })
);
AOI21_X1 #() 
AOI21_X1_2277_ (
  .A({ S91 }),
  .B1({ S22621 }),
  .B2({ S22627 }),
  .ZN({ S24189 })
);
NOR2_X1 #() 
NOR2_X1_1071_ (
  .A1({ S24189 }),
  .A2({ S83 }),
  .ZN({ S24190 })
);
INV_X1 #() 
INV_X1_1374_ (
  .A({ S24190 }),
  .ZN({ S24191 })
);
OAI211_X1 #() 
OAI211_X1_1462_ (
  .A({ S25957[1052] }),
  .B({ S24099 }),
  .C1({ S24191 }),
  .C2({ S90 }),
  .ZN({ S24192 })
);
INV_X1 #() 
INV_X1_1375_ (
  .A({ S24039 }),
  .ZN({ S24193 })
);
NAND2_X1 #() 
NAND2_X1_4215_ (
  .A1({ S24059 }),
  .A2({ S83 }),
  .ZN({ S24194 })
);
OAI21_X1 #() 
OAI21_X1_2159_ (
  .A({ S24194 }),
  .B1({ S24193 }),
  .B2({ S24113 }),
  .ZN({ S24195 })
);
OAI211_X1 #() 
OAI211_X1_1463_ (
  .A({ S24192 }),
  .B({ S25957[1053] }),
  .C1({ S24195 }),
  .C2({ S25957[1052] }),
  .ZN({ S24196 })
);
INV_X1 #() 
INV_X1_1376_ (
  .A({ S24025 }),
  .ZN({ S24197 })
);
NAND3_X1 #() 
NAND3_X1_4555_ (
  .A1({ S24197 }),
  .A2({ S22621 }),
  .A3({ S22627 }),
  .ZN({ S24198 })
);
NAND2_X1 #() 
NAND2_X1_4216_ (
  .A1({ S24198 }),
  .A2({ S83 }),
  .ZN({ S24199 })
);
NAND2_X1 #() 
NAND2_X1_4217_ (
  .A1({ S24199 }),
  .A2({ S25957[1052] }),
  .ZN({ S24200 })
);
OAI211_X1 #() 
OAI211_X1_1464_ (
  .A({ S25957[1051] }),
  .B({ S24046 }),
  .C1({ S24160 }),
  .C2({ S24070 }),
  .ZN({ S24201 })
);
OAI21_X1 #() 
OAI21_X1_2160_ (
  .A({ S24201 }),
  .B1({ S24060 }),
  .B2({ S24200 }),
  .ZN({ S24202 })
);
NAND2_X1 #() 
NAND2_X1_4218_ (
  .A1({ S24202 }),
  .A2({ S22294 }),
  .ZN({ S24203 })
);
AOI21_X1 #() 
AOI21_X1_2278_ (
  .A({ S25957[1054] }),
  .B1({ S24203 }),
  .B2({ S24196 }),
  .ZN({ S24204 })
);
OAI21_X1 #() 
OAI21_X1_2161_ (
  .A({ S22150 }),
  .B1({ S24188 }),
  .B2({ S24204 }),
  .ZN({ S24205 })
);
NAND2_X1 #() 
NAND2_X1_4219_ (
  .A1({ S24174 }),
  .A2({ S24205 }),
  .ZN({ S24206 })
);
NOR2_X1 #() 
NOR2_X1_1072_ (
  .A1({ S24206 }),
  .A2({ S21513 }),
  .ZN({ S24207 })
);
NAND2_X1 #() 
NAND2_X1_4220_ (
  .A1({ S24206 }),
  .A2({ S21513 }),
  .ZN({ S24208 })
);
INV_X1 #() 
INV_X1_1377_ (
  .A({ S24208 }),
  .ZN({ S24209 })
);
NOR2_X1 #() 
NOR2_X1_1073_ (
  .A1({ S24209 }),
  .A2({ S24207 }),
  .ZN({ S25957[966] })
);
NOR2_X1 #() 
NOR2_X1_1074_ (
  .A1({ S25957[966] }),
  .A2({ S25957[1158] }),
  .ZN({ S24210 })
);
INV_X1 #() 
INV_X1_1378_ (
  .A({ S25957[966] }),
  .ZN({ S24211 })
);
NOR2_X1 #() 
NOR2_X1_1075_ (
  .A1({ S24211 }),
  .A2({ S19194 }),
  .ZN({ S24212 })
);
NOR2_X1 #() 
NOR2_X1_1076_ (
  .A1({ S24212 }),
  .A2({ S24210 }),
  .ZN({ S25957[902] })
);
NOR2_X1 #() 
NOR2_X1_1077_ (
  .A1({ S23363 }),
  .A2({ S23362 }),
  .ZN({ S25957[1061] })
);
INV_X1 #() 
INV_X1_1379_ (
  .A({ S25957[1061] }),
  .ZN({ S24213 })
);
INV_X1 #() 
INV_X1_1380_ (
  .A({ S24138 }),
  .ZN({ S24214 })
);
AOI21_X1 #() 
AOI21_X1_2279_ (
  .A({ S25957[1048] }),
  .B1({ S83 }),
  .B2({ S25957[1049] }),
  .ZN({ S24215 })
);
OAI21_X1 #() 
OAI21_X1_2162_ (
  .A({ S24046 }),
  .B1({ S24214 }),
  .B2({ S24215 }),
  .ZN({ S24216 })
);
NAND3_X1 #() 
NAND3_X1_4556_ (
  .A1({ S24058 }),
  .A2({ S83 }),
  .A3({ S24041 }),
  .ZN({ S24217 })
);
INV_X1 #() 
INV_X1_1381_ (
  .A({ S24217 }),
  .ZN({ S24218 })
);
NAND4_X1 #() 
NAND4_X1_494_ (
  .A1({ S22621 }),
  .A2({ S22627 }),
  .A3({ S24021 }),
  .A4({ S25957[1049] }),
  .ZN({ S24219 })
);
NAND3_X1 #() 
NAND3_X1_4557_ (
  .A1({ S24065 }),
  .A2({ S25957[1051] }),
  .A3({ S24219 }),
  .ZN({ S24220 })
);
NAND2_X1 #() 
NAND2_X1_4221_ (
  .A1({ S24220 }),
  .A2({ S25957[1052] }),
  .ZN({ S24221 })
);
OAI211_X1 #() 
OAI211_X1_1465_ (
  .A({ S24216 }),
  .B({ S25957[1053] }),
  .C1({ S24221 }),
  .C2({ S24218 }),
  .ZN({ S24222 })
);
NAND2_X1 #() 
NAND2_X1_4222_ (
  .A1({ S24033 }),
  .A2({ S24047 }),
  .ZN({ S24223 })
);
AOI21_X1 #() 
AOI21_X1_2280_ (
  .A({ S24124 }),
  .B1({ S24223 }),
  .B2({ S83 }),
  .ZN({ S24224 })
);
NAND3_X1 #() 
NAND3_X1_4558_ (
  .A1({ S24033 }),
  .A2({ S25957[1051] }),
  .A3({ S24024 }),
  .ZN({ S24225 })
);
AOI21_X1 #() 
AOI21_X1_2281_ (
  .A({ S25957[1048] }),
  .B1({ S22621 }),
  .B2({ S22627 }),
  .ZN({ S24226 })
);
OAI21_X1 #() 
OAI21_X1_2163_ (
  .A({ S83 }),
  .B1({ S24160 }),
  .B2({ S24226 }),
  .ZN({ S24227 })
);
AOI21_X1 #() 
AOI21_X1_2282_ (
  .A({ S25957[1052] }),
  .B1({ S24227 }),
  .B2({ S24225 }),
  .ZN({ S24228 })
);
OR3_X1 #() 
OR3_X1_28_ (
  .A1({ S24228 }),
  .A2({ S24224 }),
  .A3({ S25957[1053] }),
  .ZN({ S24229 })
);
NAND3_X1 #() 
NAND3_X1_4559_ (
  .A1({ S24229 }),
  .A2({ S25957[1054] }),
  .A3({ S24222 }),
  .ZN({ S24230 })
);
AOI21_X1 #() 
AOI21_X1_2283_ (
  .A({ S25957[1052] }),
  .B1({ S24075 }),
  .B2({ S25957[1051] }),
  .ZN({ S24231 })
);
OAI21_X1 #() 
OAI21_X1_2164_ (
  .A({ S24231 }),
  .B1({ S24226 }),
  .B2({ S24178 }),
  .ZN({ S24232 })
);
NAND3_X1 #() 
NAND3_X1_4560_ (
  .A1({ S22621 }),
  .A2({ S22627 }),
  .A3({ S24032 }),
  .ZN({ S24233 })
);
NAND2_X1 #() 
NAND2_X1_4223_ (
  .A1({ S24219 }),
  .A2({ S83 }),
  .ZN({ S24234 })
);
OAI211_X1 #() 
OAI211_X1_1466_ (
  .A({ S24234 }),
  .B({ S25957[1052] }),
  .C1({ S83 }),
  .C2({ S24233 }),
  .ZN({ S24235 })
);
NAND3_X1 #() 
NAND3_X1_4561_ (
  .A1({ S24232 }),
  .A2({ S24235 }),
  .A3({ S25957[1053] }),
  .ZN({ S24236 })
);
NOR2_X1 #() 
NOR2_X1_1078_ (
  .A1({ S24031 }),
  .A2({ S24030 }),
  .ZN({ S24237 })
);
NAND2_X1 #() 
NAND2_X1_4224_ (
  .A1({ S90 }),
  .A2({ S83 }),
  .ZN({ S24238 })
);
NOR2_X1 #() 
NOR2_X1_1079_ (
  .A1({ S24237 }),
  .A2({ S24238 }),
  .ZN({ S24239 })
);
OAI21_X1 #() 
OAI21_X1_2165_ (
  .A({ S24046 }),
  .B1({ S24239 }),
  .B2({ S24110 }),
  .ZN({ S24240 })
);
AOI22_X1 #() 
AOI22_X1_483_ (
  .A1({ S22621 }),
  .A2({ S22627 }),
  .B1({ S91 }),
  .B2({ S24032 }),
  .ZN({ S24241 })
);
NOR2_X1 #() 
NOR2_X1_1080_ (
  .A1({ S25957[1050] }),
  .A2({ S24025 }),
  .ZN({ S24242 })
);
NOR3_X1 #() 
NOR3_X1_145_ (
  .A1({ S24242 }),
  .A2({ S24241 }),
  .A3({ S83 }),
  .ZN({ S24243 })
);
NAND3_X1 #() 
NAND3_X1_4562_ (
  .A1({ S24051 }),
  .A2({ S83 }),
  .A3({ S24064 }),
  .ZN({ S24244 })
);
NAND2_X1 #() 
NAND2_X1_4225_ (
  .A1({ S24244 }),
  .A2({ S25957[1052] }),
  .ZN({ S24245 })
);
OAI21_X1 #() 
OAI21_X1_2166_ (
  .A({ S24240 }),
  .B1({ S24243 }),
  .B2({ S24245 }),
  .ZN({ S24246 })
);
NAND2_X1 #() 
NAND2_X1_4226_ (
  .A1({ S24246 }),
  .A2({ S22294 }),
  .ZN({ S24247 })
);
AOI21_X1 #() 
AOI21_X1_2284_ (
  .A({ S25957[1054] }),
  .B1({ S24247 }),
  .B2({ S24236 }),
  .ZN({ S24248 })
);
INV_X1 #() 
INV_X1_1382_ (
  .A({ S24248 }),
  .ZN({ S24249 })
);
AOI21_X1 #() 
AOI21_X1_2285_ (
  .A({ S25957[1055] }),
  .B1({ S24249 }),
  .B2({ S24230 }),
  .ZN({ S24250 })
);
NAND2_X1 #() 
NAND2_X1_4227_ (
  .A1({ S25957[1050] }),
  .A2({ S24026 }),
  .ZN({ S24251 })
);
AOI21_X1 #() 
AOI21_X1_2286_ (
  .A({ S83 }),
  .B1({ S24251 }),
  .B2({ S24233 }),
  .ZN({ S24252 })
);
NAND2_X1 #() 
NAND2_X1_4228_ (
  .A1({ S24138 }),
  .A2({ S24085 }),
  .ZN({ S24253 })
);
OAI21_X1 #() 
OAI21_X1_2167_ (
  .A({ S24046 }),
  .B1({ S24252 }),
  .B2({ S24253 }),
  .ZN({ S24254 })
);
OAI221_X1 #() 
OAI221_X1_120_ (
  .A({ S25957[1052] }),
  .B1({ S24144 }),
  .B2({ S24112 }),
  .C1({ S24101 }),
  .C2({ S25957[1048] }),
  .ZN({ S24255 })
);
NAND3_X1 #() 
NAND3_X1_4563_ (
  .A1({ S24254 }),
  .A2({ S25957[1053] }),
  .A3({ S24255 }),
  .ZN({ S24256 })
);
NAND3_X1 #() 
NAND3_X1_4564_ (
  .A1({ S24026 }),
  .A2({ S22621 }),
  .A3({ S22627 }),
  .ZN({ S24257 })
);
OAI211_X1 #() 
OAI211_X1_1467_ (
  .A({ S24257 }),
  .B({ S25957[1052] }),
  .C1({ S25957[1051] }),
  .C2({ S24026 }),
  .ZN({ S24258 })
);
OAI21_X1 #() 
OAI21_X1_2168_ (
  .A({ S24046 }),
  .B1({ S24184 }),
  .B2({ S24066 }),
  .ZN({ S24259 })
);
NAND3_X1 #() 
NAND3_X1_4565_ (
  .A1({ S24259 }),
  .A2({ S24258 }),
  .A3({ S22294 }),
  .ZN({ S24260 })
);
NAND3_X1 #() 
NAND3_X1_4566_ (
  .A1({ S24256 }),
  .A2({ S24260 }),
  .A3({ S25957[1054] }),
  .ZN({ S24261 })
);
NAND2_X1 #() 
NAND2_X1_4229_ (
  .A1({ S24047 }),
  .A2({ S83 }),
  .ZN({ S24262 })
);
INV_X1 #() 
INV_X1_1383_ (
  .A({ S24262 }),
  .ZN({ S24263 })
);
NAND2_X1 #() 
NAND2_X1_4230_ (
  .A1({ S24027 }),
  .A2({ S25957[1050] }),
  .ZN({ S24264 })
);
AOI21_X1 #() 
AOI21_X1_2287_ (
  .A({ S83 }),
  .B1({ S24264 }),
  .B2({ S24090 }),
  .ZN({ S24265 })
);
OAI21_X1 #() 
OAI21_X1_2169_ (
  .A({ S24046 }),
  .B1({ S24265 }),
  .B2({ S24263 }),
  .ZN({ S24266 })
);
NOR2_X1 #() 
NOR2_X1_1081_ (
  .A1({ S24102 }),
  .A2({ S83 }),
  .ZN({ S24267 })
);
OAI21_X1 #() 
OAI21_X1_2170_ (
  .A({ S25957[1052] }),
  .B1({ S24099 }),
  .B2({ S25957[1049] }),
  .ZN({ S24268 })
);
OAI21_X1 #() 
OAI21_X1_2171_ (
  .A({ S24266 }),
  .B1({ S24267 }),
  .B2({ S24268 }),
  .ZN({ S24269 })
);
INV_X1 #() 
INV_X1_1384_ (
  .A({ S24074 }),
  .ZN({ S24270 })
);
NAND2_X1 #() 
NAND2_X1_4231_ (
  .A1({ S25957[1051] }),
  .A2({ S24022 }),
  .ZN({ S24271 })
);
OAI21_X1 #() 
OAI21_X1_2172_ (
  .A({ S24271 }),
  .B1({ S24270 }),
  .B2({ S24112 }),
  .ZN({ S24272 })
);
NAND2_X1 #() 
NAND2_X1_4232_ (
  .A1({ S24272 }),
  .A2({ S24046 }),
  .ZN({ S24273 })
);
NAND2_X1 #() 
NAND2_X1_4233_ (
  .A1({ S24051 }),
  .A2({ S83 }),
  .ZN({ S24274 })
);
NAND3_X1 #() 
NAND3_X1_4567_ (
  .A1({ S24033 }),
  .A2({ S25957[1051] }),
  .A3({ S24041 }),
  .ZN({ S24275 })
);
NAND2_X1 #() 
NAND2_X1_4234_ (
  .A1({ S24275 }),
  .A2({ S24274 }),
  .ZN({ S24276 })
);
NAND3_X1 #() 
NAND3_X1_4568_ (
  .A1({ S24276 }),
  .A2({ S25957[1052] }),
  .A3({ S24238 }),
  .ZN({ S24277 })
);
NAND3_X1 #() 
NAND3_X1_4569_ (
  .A1({ S24277 }),
  .A2({ S25957[1053] }),
  .A3({ S24273 }),
  .ZN({ S24278 })
);
OAI211_X1 #() 
OAI211_X1_1468_ (
  .A({ S24278 }),
  .B({ S22219 }),
  .C1({ S24269 }),
  .C2({ S25957[1053] }),
  .ZN({ S24279 })
);
AOI21_X1 #() 
AOI21_X1_2288_ (
  .A({ S22150 }),
  .B1({ S24279 }),
  .B2({ S24261 }),
  .ZN({ S24280 })
);
OAI21_X1 #() 
OAI21_X1_2173_ (
  .A({ S25957[1221] }),
  .B1({ S24250 }),
  .B2({ S24280 }),
  .ZN({ S24281 })
);
OAI21_X1 #() 
OAI21_X1_2174_ (
  .A({ S24216 }),
  .B1({ S24221 }),
  .B2({ S24218 }),
  .ZN({ S24282 })
);
NAND2_X1 #() 
NAND2_X1_4235_ (
  .A1({ S24282 }),
  .A2({ S25957[1053] }),
  .ZN({ S24283 })
);
OAI21_X1 #() 
OAI21_X1_2175_ (
  .A({ S22294 }),
  .B1({ S24228 }),
  .B2({ S24224 }),
  .ZN({ S24284 })
);
AOI21_X1 #() 
AOI21_X1_2289_ (
  .A({ S22219 }),
  .B1({ S24283 }),
  .B2({ S24284 }),
  .ZN({ S24285 })
);
OAI21_X1 #() 
OAI21_X1_2176_ (
  .A({ S22150 }),
  .B1({ S24285 }),
  .B2({ S24248 }),
  .ZN({ S24286 })
);
NAND2_X1 #() 
NAND2_X1_4236_ (
  .A1({ S24279 }),
  .A2({ S24261 }),
  .ZN({ S24287 })
);
NAND2_X1 #() 
NAND2_X1_4237_ (
  .A1({ S24287 }),
  .A2({ S25957[1055] }),
  .ZN({ S24288 })
);
NAND3_X1 #() 
NAND3_X1_4570_ (
  .A1({ S24288 }),
  .A2({ S21649 }),
  .A3({ S24286 }),
  .ZN({ S24289 })
);
NAND3_X1 #() 
NAND3_X1_4571_ (
  .A1({ S24281 }),
  .A2({ S24289 }),
  .A3({ S24213 }),
  .ZN({ S24290 })
);
AOI21_X1 #() 
AOI21_X1_2290_ (
  .A({ S21649 }),
  .B1({ S24288 }),
  .B2({ S24286 }),
  .ZN({ S24291 })
);
NOR3_X1 #() 
NOR3_X1_146_ (
  .A1({ S24250 }),
  .A2({ S24280 }),
  .A3({ S25957[1221] }),
  .ZN({ S24292 })
);
OAI21_X1 #() 
OAI21_X1_2177_ (
  .A({ S25957[1061] }),
  .B1({ S24292 }),
  .B2({ S24291 }),
  .ZN({ S24293 })
);
NAND3_X1 #() 
NAND3_X1_4572_ (
  .A1({ S24293 }),
  .A2({ S23368 }),
  .A3({ S24290 }),
  .ZN({ S24294 })
);
OAI21_X1 #() 
OAI21_X1_2178_ (
  .A({ S24213 }),
  .B1({ S24292 }),
  .B2({ S24291 }),
  .ZN({ S24295 })
);
NAND3_X1 #() 
NAND3_X1_4573_ (
  .A1({ S24281 }),
  .A2({ S24289 }),
  .A3({ S25957[1061] }),
  .ZN({ S24296 })
);
NAND3_X1 #() 
NAND3_X1_4574_ (
  .A1({ S24295 }),
  .A2({ S25957[1029] }),
  .A3({ S24296 }),
  .ZN({ S24297 })
);
NAND2_X1 #() 
NAND2_X1_4238_ (
  .A1({ S24294 }),
  .A2({ S24297 }),
  .ZN({ S25957[901] })
);
NAND2_X1 #() 
NAND2_X1_4239_ (
  .A1({ S21739 }),
  .A2({ S21742 }),
  .ZN({ S24298 })
);
INV_X1 #() 
INV_X1_1385_ (
  .A({ S24298 }),
  .ZN({ S25957[1060] })
);
AOI21_X1 #() 
AOI21_X1_2291_ (
  .A({ S25957[1051] }),
  .B1({ S24033 }),
  .B2({ S24034 }),
  .ZN({ S24299 })
);
OAI21_X1 #() 
OAI21_X1_2179_ (
  .A({ S83 }),
  .B1({ S24160 }),
  .B2({ S24104 }),
  .ZN({ S24300 })
);
NAND3_X1 #() 
NAND3_X1_4575_ (
  .A1({ S24219 }),
  .A2({ S25957[1051] }),
  .A3({ S24025 }),
  .ZN({ S24301 })
);
NAND3_X1 #() 
NAND3_X1_4576_ (
  .A1({ S24300 }),
  .A2({ S25957[1052] }),
  .A3({ S24301 }),
  .ZN({ S24302 })
);
NAND2_X1 #() 
NAND2_X1_4240_ (
  .A1({ S24052 }),
  .A2({ S25957[1051] }),
  .ZN({ S24303 })
);
NAND3_X1 #() 
NAND3_X1_4577_ (
  .A1({ S24123 }),
  .A2({ S24303 }),
  .A3({ S24046 }),
  .ZN({ S24304 })
);
OAI211_X1 #() 
OAI211_X1_1469_ (
  .A({ S24302 }),
  .B({ S25957[1053] }),
  .C1({ S24299 }),
  .C2({ S24304 }),
  .ZN({ S24305 })
);
AOI21_X1 #() 
AOI21_X1_2292_ (
  .A({ S25957[1051] }),
  .B1({ S24053 }),
  .B2({ S24257 }),
  .ZN({ S24306 })
);
NOR2_X1 #() 
NOR2_X1_1082_ (
  .A1({ S25957[1052] }),
  .A2({ S24087 }),
  .ZN({ S24307 })
);
NOR2_X1 #() 
NOR2_X1_1083_ (
  .A1({ S25957[1052] }),
  .A2({ S24021 }),
  .ZN({ S24308 })
);
AOI21_X1 #() 
AOI21_X1_2293_ (
  .A({ S24307 }),
  .B1({ S25957[1050] }),
  .B2({ S24308 }),
  .ZN({ S24309 })
);
NAND3_X1 #() 
NAND3_X1_4578_ (
  .A1({ S24053 }),
  .A2({ S83 }),
  .A3({ S24047 }),
  .ZN({ S24310 })
);
NAND3_X1 #() 
NAND3_X1_4579_ (
  .A1({ S24251 }),
  .A2({ S25957[1051] }),
  .A3({ S24039 }),
  .ZN({ S24311 })
);
NAND3_X1 #() 
NAND3_X1_4580_ (
  .A1({ S24311 }),
  .A2({ S24310 }),
  .A3({ S25957[1052] }),
  .ZN({ S24312 })
);
OAI211_X1 #() 
OAI211_X1_1470_ (
  .A({ S24312 }),
  .B({ S22294 }),
  .C1({ S24306 }),
  .C2({ S24309 }),
  .ZN({ S24313 })
);
NAND3_X1 #() 
NAND3_X1_4581_ (
  .A1({ S24305 }),
  .A2({ S24313 }),
  .A3({ S22219 }),
  .ZN({ S24314 })
);
NOR2_X1 #() 
NOR2_X1_1084_ (
  .A1({ S24189 }),
  .A2({ S25957[1051] }),
  .ZN({ S24315 })
);
NAND3_X1 #() 
NAND3_X1_4582_ (
  .A1({ S24039 }),
  .A2({ S83 }),
  .A3({ S24021 }),
  .ZN({ S24316 })
);
OAI211_X1 #() 
OAI211_X1_1471_ (
  .A({ S24046 }),
  .B({ S24316 }),
  .C1({ S24120 }),
  .C2({ S83 }),
  .ZN({ S24317 })
);
OAI211_X1 #() 
OAI211_X1_1472_ (
  .A({ S24317 }),
  .B({ S25957[1053] }),
  .C1({ S24124 }),
  .C2({ S24315 }),
  .ZN({ S24318 })
);
NOR2_X1 #() 
NOR2_X1_1085_ (
  .A1({ S24226 }),
  .A2({ S25957[1051] }),
  .ZN({ S24319 })
);
NAND2_X1 #() 
NAND2_X1_4241_ (
  .A1({ S24319 }),
  .A2({ S24074 }),
  .ZN({ S24320 })
);
NAND3_X1 #() 
NAND3_X1_4583_ (
  .A1({ S24320 }),
  .A2({ S24046 }),
  .A3({ S24080 }),
  .ZN({ S24321 })
);
INV_X1 #() 
INV_X1_1386_ (
  .A({ S24112 }),
  .ZN({ S24322 })
);
AOI21_X1 #() 
AOI21_X1_2294_ (
  .A({ S24046 }),
  .B1({ S24322 }),
  .B2({ S24074 }),
  .ZN({ S24323 })
);
OAI21_X1 #() 
OAI21_X1_2180_ (
  .A({ S24323 }),
  .B1({ S25957[1049] }),
  .B2({ S24175 }),
  .ZN({ S24324 })
);
NAND3_X1 #() 
NAND3_X1_4584_ (
  .A1({ S24321 }),
  .A2({ S24324 }),
  .A3({ S22294 }),
  .ZN({ S24325 })
);
NAND3_X1 #() 
NAND3_X1_4585_ (
  .A1({ S24318 }),
  .A2({ S24325 }),
  .A3({ S25957[1054] }),
  .ZN({ S24326 })
);
NAND3_X1 #() 
NAND3_X1_4586_ (
  .A1({ S24326 }),
  .A2({ S24314 }),
  .A3({ S25957[1055] }),
  .ZN({ S24327 })
);
AOI21_X1 #() 
AOI21_X1_2295_ (
  .A({ S83 }),
  .B1({ S24024 }),
  .B2({ S24026 }),
  .ZN({ S24328 })
);
AOI21_X1 #() 
AOI21_X1_2296_ (
  .A({ S25957[1051] }),
  .B1({ S24146 }),
  .B2({ S24090 }),
  .ZN({ S24329 })
);
OAI21_X1 #() 
OAI21_X1_2181_ (
  .A({ S24046 }),
  .B1({ S24329 }),
  .B2({ S24328 }),
  .ZN({ S24330 })
);
NAND3_X1 #() 
NAND3_X1_4587_ (
  .A1({ S24038 }),
  .A2({ S25957[1051] }),
  .A3({ S24041 }),
  .ZN({ S24331 })
);
AOI21_X1 #() 
AOI21_X1_2297_ (
  .A({ S25957[1053] }),
  .B1({ S24323 }),
  .B2({ S24331 }),
  .ZN({ S24332 })
);
OAI221_X1 #() 
OAI221_X1_121_ (
  .A({ S25957[1052] }),
  .B1({ S24112 }),
  .B2({ S24237 }),
  .C1({ S24059 }),
  .C2({ S83 }),
  .ZN({ S24333 })
);
OAI21_X1 #() 
OAI21_X1_2182_ (
  .A({ S24238 }),
  .B1({ S24102 }),
  .B2({ S83 }),
  .ZN({ S24334 })
);
AOI21_X1 #() 
AOI21_X1_2298_ (
  .A({ S22294 }),
  .B1({ S24334 }),
  .B2({ S24046 }),
  .ZN({ S24335 })
);
AOI22_X1 #() 
AOI22_X1_484_ (
  .A1({ S24333 }),
  .A2({ S24335 }),
  .B1({ S24330 }),
  .B2({ S24332 }),
  .ZN({ S24336 })
);
AOI21_X1 #() 
AOI21_X1_2299_ (
  .A({ S24046 }),
  .B1({ S24237 }),
  .B2({ S126 }),
  .ZN({ S24337 })
);
NAND2_X1 #() 
NAND2_X1_4242_ (
  .A1({ S25957[1050] }),
  .A2({ S25957[1051] }),
  .ZN({ S24338 })
);
OAI211_X1 #() 
OAI211_X1_1473_ (
  .A({ S24046 }),
  .B({ S24338 }),
  .C1({ S24262 }),
  .C2({ S24226 }),
  .ZN({ S24339 })
);
NAND2_X1 #() 
NAND2_X1_4243_ (
  .A1({ S24165 }),
  .A2({ S83 }),
  .ZN({ S24340 })
);
NOR2_X1 #() 
NOR2_X1_1086_ (
  .A1({ S24120 }),
  .A2({ S24340 }),
  .ZN({ S24341 })
);
OAI211_X1 #() 
OAI211_X1_1474_ (
  .A({ S22294 }),
  .B({ S24339 }),
  .C1({ S24341 }),
  .C2({ S24089 }),
  .ZN({ S24342 })
);
AOI21_X1 #() 
AOI21_X1_2300_ (
  .A({ S25957[1051] }),
  .B1({ S24251 }),
  .B2({ S24102 }),
  .ZN({ S24343 })
);
NAND2_X1 #() 
NAND2_X1_4244_ (
  .A1({ S24225 }),
  .A2({ S24046 }),
  .ZN({ S24344 })
);
OAI21_X1 #() 
OAI21_X1_2183_ (
  .A({ S25957[1053] }),
  .B1({ S24344 }),
  .B2({ S24343 }),
  .ZN({ S24345 })
);
OAI211_X1 #() 
OAI211_X1_1475_ (
  .A({ S24342 }),
  .B({ S25957[1054] }),
  .C1({ S24337 }),
  .C2({ S24345 }),
  .ZN({ S24346 })
);
OAI211_X1 #() 
OAI211_X1_1476_ (
  .A({ S24346 }),
  .B({ S22150 }),
  .C1({ S24336 }),
  .C2({ S25957[1054] }),
  .ZN({ S24347 })
);
NAND3_X1 #() 
NAND3_X1_4588_ (
  .A1({ S24347 }),
  .A2({ S24327 }),
  .A3({ S19311 }),
  .ZN({ S24348 })
);
NAND2_X1 #() 
NAND2_X1_4245_ (
  .A1({ S24347 }),
  .A2({ S24327 }),
  .ZN({ S24349 })
);
NAND2_X1 #() 
NAND2_X1_4246_ (
  .A1({ S24349 }),
  .A2({ S25957[1220] }),
  .ZN({ S24350 })
);
NAND3_X1 #() 
NAND3_X1_4589_ (
  .A1({ S24350 }),
  .A2({ S24298 }),
  .A3({ S24348 }),
  .ZN({ S24351 })
);
NAND2_X1 #() 
NAND2_X1_4247_ (
  .A1({ S24350 }),
  .A2({ S24348 }),
  .ZN({ S25957[964] })
);
NAND2_X1 #() 
NAND2_X1_4248_ (
  .A1({ S25957[964] }),
  .A2({ S25957[1060] }),
  .ZN({ S24352 })
);
NAND3_X1 #() 
NAND3_X1_4590_ (
  .A1({ S24352 }),
  .A2({ S23396 }),
  .A3({ S24351 }),
  .ZN({ S24353 })
);
NAND2_X1 #() 
NAND2_X1_4249_ (
  .A1({ S21736 }),
  .A2({ S21737 }),
  .ZN({ S25957[1124] })
);
NAND3_X1 #() 
NAND3_X1_4591_ (
  .A1({ S24347 }),
  .A2({ S24327 }),
  .A3({ S25957[1124] }),
  .ZN({ S24354 })
);
INV_X1 #() 
INV_X1_1387_ (
  .A({ S24354 }),
  .ZN({ S24355 })
);
AOI21_X1 #() 
AOI21_X1_2301_ (
  .A({ S25957[1124] }),
  .B1({ S24347 }),
  .B2({ S24327 }),
  .ZN({ S24356 })
);
OAI21_X1 #() 
OAI21_X1_2184_ (
  .A({ S25957[1188] }),
  .B1({ S24355 }),
  .B2({ S24356 }),
  .ZN({ S24357 })
);
INV_X1 #() 
INV_X1_1388_ (
  .A({ S24356 }),
  .ZN({ S24358 })
);
NAND3_X1 #() 
NAND3_X1_4592_ (
  .A1({ S24358 }),
  .A2({ S21657 }),
  .A3({ S24354 }),
  .ZN({ S24359 })
);
NAND3_X1 #() 
NAND3_X1_4593_ (
  .A1({ S24357 }),
  .A2({ S24359 }),
  .A3({ S25957[1028] }),
  .ZN({ S24360 })
);
NAND2_X1 #() 
NAND2_X1_4250_ (
  .A1({ S24353 }),
  .A2({ S24360 }),
  .ZN({ S25957[900] })
);
NOR2_X1 #() 
NOR2_X1_1087_ (
  .A1({ S19371 }),
  .A2({ S19372 }),
  .ZN({ S25957[1187] })
);
INV_X1 #() 
INV_X1_1389_ (
  .A({ S25957[1187] }),
  .ZN({ S24361 })
);
NAND2_X1 #() 
NAND2_X1_4251_ (
  .A1({ S21830 }),
  .A2({ S21831 }),
  .ZN({ S25957[1123] })
);
OAI21_X1 #() 
OAI21_X1_2185_ (
  .A({ S25957[1051] }),
  .B1({ S24103 }),
  .B2({ S24189 }),
  .ZN({ S24362 })
);
OAI211_X1 #() 
OAI211_X1_1477_ (
  .A({ S24362 }),
  .B({ S25957[1052] }),
  .C1({ S25957[1051] }),
  .C2({ S24141 }),
  .ZN({ S24363 })
);
OAI21_X1 #() 
OAI21_X1_2186_ (
  .A({ S24021 }),
  .B1({ S24031 }),
  .B2({ S24030 }),
  .ZN({ S24364 })
);
NAND4_X1 #() 
NAND4_X1_495_ (
  .A1({ S24364 }),
  .A2({ S24024 }),
  .A3({ S25957[1049] }),
  .A4({ S25957[1051] }),
  .ZN({ S24365 })
);
NAND2_X1 #() 
NAND2_X1_4252_ (
  .A1({ S24028 }),
  .A2({ S24074 }),
  .ZN({ S24366 })
);
NAND2_X1 #() 
NAND2_X1_4253_ (
  .A1({ S24366 }),
  .A2({ S24365 }),
  .ZN({ S24367 })
);
NAND2_X1 #() 
NAND2_X1_4254_ (
  .A1({ S24367 }),
  .A2({ S24046 }),
  .ZN({ S24368 })
);
NAND3_X1 #() 
NAND3_X1_4594_ (
  .A1({ S24368 }),
  .A2({ S24363 }),
  .A3({ S25957[1053] }),
  .ZN({ S24369 })
);
NAND2_X1 #() 
NAND2_X1_4255_ (
  .A1({ S24034 }),
  .A2({ S25957[1051] }),
  .ZN({ S24370 })
);
INV_X1 #() 
INV_X1_1390_ (
  .A({ S24370 }),
  .ZN({ S24371 })
);
NAND4_X1 #() 
NAND4_X1_496_ (
  .A1({ S22621 }),
  .A2({ S22627 }),
  .A3({ S83 }),
  .A4({ S25957[1049] }),
  .ZN({ S24372 })
);
NAND3_X1 #() 
NAND3_X1_4595_ (
  .A1({ S24138 }),
  .A2({ S25957[1052] }),
  .A3({ S24372 }),
  .ZN({ S24373 })
);
AOI21_X1 #() 
AOI21_X1_2302_ (
  .A({ S83 }),
  .B1({ S24264 }),
  .B2({ S24039 }),
  .ZN({ S24374 })
);
OAI21_X1 #() 
OAI21_X1_2187_ (
  .A({ S24046 }),
  .B1({ S24075 }),
  .B2({ S24112 }),
  .ZN({ S24375 })
);
OAI22_X1 #() 
OAI22_X1_110_ (
  .A1({ S24374 }),
  .A2({ S24375 }),
  .B1({ S24371 }),
  .B2({ S24373 }),
  .ZN({ S24376 })
);
NAND2_X1 #() 
NAND2_X1_4256_ (
  .A1({ S24376 }),
  .A2({ S22294 }),
  .ZN({ S24377 })
);
NAND3_X1 #() 
NAND3_X1_4596_ (
  .A1({ S24369 }),
  .A2({ S22219 }),
  .A3({ S24377 }),
  .ZN({ S24378 })
);
NAND3_X1 #() 
NAND3_X1_4597_ (
  .A1({ S24024 }),
  .A2({ S25957[1051] }),
  .A3({ S24026 }),
  .ZN({ S24379 })
);
NAND3_X1 #() 
NAND3_X1_4598_ (
  .A1({ S24051 }),
  .A2({ S24027 }),
  .A3({ S83 }),
  .ZN({ S24380 })
);
AOI21_X1 #() 
AOI21_X1_2303_ (
  .A({ S24046 }),
  .B1({ S24379 }),
  .B2({ S24380 }),
  .ZN({ S24381 })
);
NAND2_X1 #() 
NAND2_X1_4257_ (
  .A1({ S24319 }),
  .A2({ S24064 }),
  .ZN({ S24382 })
);
NAND3_X1 #() 
NAND3_X1_4599_ (
  .A1({ S24140 }),
  .A2({ S25957[1051] }),
  .A3({ S24257 }),
  .ZN({ S24383 })
);
AOI21_X1 #() 
AOI21_X1_2304_ (
  .A({ S25957[1052] }),
  .B1({ S24382 }),
  .B2({ S24383 }),
  .ZN({ S24384 })
);
OAI21_X1 #() 
OAI21_X1_2188_ (
  .A({ S25957[1053] }),
  .B1({ S24384 }),
  .B2({ S24381 }),
  .ZN({ S24385 })
);
NAND2_X1 #() 
NAND2_X1_4258_ (
  .A1({ S24165 }),
  .A2({ S24092 }),
  .ZN({ S24386 })
);
NAND3_X1 #() 
NAND3_X1_4600_ (
  .A1({ S24065 }),
  .A2({ S24198 }),
  .A3({ S83 }),
  .ZN({ S24387 })
);
AOI21_X1 #() 
AOI21_X1_2305_ (
  .A({ S24046 }),
  .B1({ S24387 }),
  .B2({ S24386 }),
  .ZN({ S24388 })
);
NAND4_X1 #() 
NAND4_X1_497_ (
  .A1({ S24338 }),
  .A2({ S24024 }),
  .A3({ S91 }),
  .A4({ S24046 }),
  .ZN({ S24389 })
);
INV_X1 #() 
INV_X1_1391_ (
  .A({ S24389 }),
  .ZN({ S24390 })
);
OAI21_X1 #() 
OAI21_X1_2189_ (
  .A({ S22294 }),
  .B1({ S24388 }),
  .B2({ S24390 }),
  .ZN({ S24391 })
);
NAND3_X1 #() 
NAND3_X1_4601_ (
  .A1({ S24385 }),
  .A2({ S25957[1054] }),
  .A3({ S24391 }),
  .ZN({ S24392 })
);
NAND3_X1 #() 
NAND3_X1_4602_ (
  .A1({ S24378 }),
  .A2({ S24392 }),
  .A3({ S25957[1055] }),
  .ZN({ S24393 })
);
NAND3_X1 #() 
NAND3_X1_4603_ (
  .A1({ S24142 }),
  .A2({ S24068 }),
  .A3({ S25957[1052] }),
  .ZN({ S24394 })
);
NAND3_X1 #() 
NAND3_X1_4604_ (
  .A1({ S24039 }),
  .A2({ S83 }),
  .A3({ S24025 }),
  .ZN({ S24395 })
);
OAI211_X1 #() 
OAI211_X1_1478_ (
  .A({ S24046 }),
  .B({ S24395 }),
  .C1({ S24119 }),
  .C2({ S83 }),
  .ZN({ S24396 })
);
NAND3_X1 #() 
NAND3_X1_4605_ (
  .A1({ S24394 }),
  .A2({ S24396 }),
  .A3({ S25957[1053] }),
  .ZN({ S24397 })
);
NAND2_X1 #() 
NAND2_X1_4259_ (
  .A1({ S24032 }),
  .A2({ S83 }),
  .ZN({ S24398 })
);
OR2_X1 #() 
OR2_X1_59_ (
  .A1({ S24075 }),
  .A2({ S24398 }),
  .ZN({ S24399 })
);
NAND2_X1 #() 
NAND2_X1_4260_ (
  .A1({ S24399 }),
  .A2({ S25957[1052] }),
  .ZN({ S24400 })
);
NAND3_X1 #() 
NAND3_X1_4606_ (
  .A1({ S24033 }),
  .A2({ S24041 }),
  .A3({ S83 }),
  .ZN({ S24401 })
);
NAND3_X1 #() 
NAND3_X1_4607_ (
  .A1({ S24401 }),
  .A2({ S24231 }),
  .A3({ S24123 }),
  .ZN({ S24402 })
);
NAND3_X1 #() 
NAND3_X1_4608_ (
  .A1({ S24402 }),
  .A2({ S22294 }),
  .A3({ S24400 }),
  .ZN({ S24403 })
);
NAND3_X1 #() 
NAND3_X1_4609_ (
  .A1({ S24397 }),
  .A2({ S25957[1054] }),
  .A3({ S24403 }),
  .ZN({ S24404 })
);
OAI211_X1 #() 
OAI211_X1_1479_ (
  .A({ S25957[1051] }),
  .B({ S91 }),
  .C1({ S25957[1050] }),
  .C2({ S24032 }),
  .ZN({ S24405 })
);
AOI21_X1 #() 
AOI21_X1_2306_ (
  .A({ S24046 }),
  .B1({ S24217 }),
  .B2({ S24405 }),
  .ZN({ S24406 })
);
NAND3_X1 #() 
NAND3_X1_4610_ (
  .A1({ S24364 }),
  .A2({ S25957[1051] }),
  .A3({ S24047 }),
  .ZN({ S24407 })
);
AOI21_X1 #() 
AOI21_X1_2307_ (
  .A({ S25957[1052] }),
  .B1({ S24029 }),
  .B2({ S24407 }),
  .ZN({ S24408 })
);
OAI21_X1 #() 
OAI21_X1_2190_ (
  .A({ S22294 }),
  .B1({ S24408 }),
  .B2({ S24406 }),
  .ZN({ S24409 })
);
OAI21_X1 #() 
OAI21_X1_2191_ (
  .A({ S25957[1052] }),
  .B1({ S24239 }),
  .B2({ S24189 }),
  .ZN({ S24410 })
);
NAND3_X1 #() 
NAND3_X1_4611_ (
  .A1({ S24113 }),
  .A2({ S24039 }),
  .A3({ S24308 }),
  .ZN({ S24411 })
);
NAND3_X1 #() 
NAND3_X1_4612_ (
  .A1({ S24411 }),
  .A2({ S24410 }),
  .A3({ S25957[1053] }),
  .ZN({ S24412 })
);
NAND3_X1 #() 
NAND3_X1_4613_ (
  .A1({ S24409 }),
  .A2({ S22219 }),
  .A3({ S24412 }),
  .ZN({ S24413 })
);
NAND3_X1 #() 
NAND3_X1_4614_ (
  .A1({ S24413 }),
  .A2({ S24404 }),
  .A3({ S22150 }),
  .ZN({ S24414 })
);
NAND3_X1 #() 
NAND3_X1_4615_ (
  .A1({ S24393 }),
  .A2({ S25957[1123] }),
  .A3({ S24414 }),
  .ZN({ S24415 })
);
INV_X1 #() 
INV_X1_1392_ (
  .A({ S25957[1123] }),
  .ZN({ S24416 })
);
NAND2_X1 #() 
NAND2_X1_4261_ (
  .A1({ S24397 }),
  .A2({ S24403 }),
  .ZN({ S24417 })
);
NAND2_X1 #() 
NAND2_X1_4262_ (
  .A1({ S24417 }),
  .A2({ S25957[1054] }),
  .ZN({ S24418 })
);
NAND2_X1 #() 
NAND2_X1_4263_ (
  .A1({ S24411 }),
  .A2({ S24410 }),
  .ZN({ S24419 })
);
NAND2_X1 #() 
NAND2_X1_4264_ (
  .A1({ S24419 }),
  .A2({ S25957[1053] }),
  .ZN({ S24420 })
);
INV_X1 #() 
INV_X1_1393_ (
  .A({ S24406 }),
  .ZN({ S24421 })
);
INV_X1 #() 
INV_X1_1394_ (
  .A({ S24408 }),
  .ZN({ S24422 })
);
NAND3_X1 #() 
NAND3_X1_4616_ (
  .A1({ S24422 }),
  .A2({ S22294 }),
  .A3({ S24421 }),
  .ZN({ S24423 })
);
NAND3_X1 #() 
NAND3_X1_4617_ (
  .A1({ S24423 }),
  .A2({ S22219 }),
  .A3({ S24420 }),
  .ZN({ S24424 })
);
NAND3_X1 #() 
NAND3_X1_4618_ (
  .A1({ S24418 }),
  .A2({ S24424 }),
  .A3({ S22150 }),
  .ZN({ S24425 })
);
INV_X1 #() 
INV_X1_1395_ (
  .A({ S24388 }),
  .ZN({ S24426 })
);
NAND3_X1 #() 
NAND3_X1_4619_ (
  .A1({ S24426 }),
  .A2({ S22294 }),
  .A3({ S24389 }),
  .ZN({ S24427 })
);
INV_X1 #() 
INV_X1_1396_ (
  .A({ S24381 }),
  .ZN({ S24428 })
);
AND2_X1 #() 
AND2_X1_267_ (
  .A1({ S24382 }),
  .A2({ S24383 }),
  .ZN({ S24429 })
);
OAI211_X1 #() 
OAI211_X1_1480_ (
  .A({ S25957[1053] }),
  .B({ S24428 }),
  .C1({ S24429 }),
  .C2({ S25957[1052] }),
  .ZN({ S24430 })
);
NAND3_X1 #() 
NAND3_X1_4620_ (
  .A1({ S24430 }),
  .A2({ S24427 }),
  .A3({ S25957[1054] }),
  .ZN({ S24431 })
);
NAND2_X1 #() 
NAND2_X1_4265_ (
  .A1({ S24141 }),
  .A2({ S83 }),
  .ZN({ S24432 })
);
OAI211_X1 #() 
OAI211_X1_1481_ (
  .A({ S24432 }),
  .B({ S25957[1052] }),
  .C1({ S24191 }),
  .C2({ S24103 }),
  .ZN({ S24433 })
);
NAND3_X1 #() 
NAND3_X1_4621_ (
  .A1({ S24366 }),
  .A2({ S24046 }),
  .A3({ S24365 }),
  .ZN({ S24434 })
);
NAND3_X1 #() 
NAND3_X1_4622_ (
  .A1({ S24433 }),
  .A2({ S25957[1053] }),
  .A3({ S24434 }),
  .ZN({ S24435 })
);
OAI221_X1 #() 
OAI221_X1_122_ (
  .A({ S22294 }),
  .B1({ S24371 }),
  .B2({ S24373 }),
  .C1({ S24374 }),
  .C2({ S24375 }),
  .ZN({ S24436 })
);
NAND3_X1 #() 
NAND3_X1_4623_ (
  .A1({ S24435 }),
  .A2({ S24436 }),
  .A3({ S22219 }),
  .ZN({ S24437 })
);
NAND3_X1 #() 
NAND3_X1_4624_ (
  .A1({ S24431 }),
  .A2({ S24437 }),
  .A3({ S25957[1055] }),
  .ZN({ S24438 })
);
NAND3_X1 #() 
NAND3_X1_4625_ (
  .A1({ S24425 }),
  .A2({ S24438 }),
  .A3({ S24416 }),
  .ZN({ S24439 })
);
NAND3_X1 #() 
NAND3_X1_4626_ (
  .A1({ S24439 }),
  .A2({ S24415 }),
  .A3({ S24361 }),
  .ZN({ S24440 })
);
NAND3_X1 #() 
NAND3_X1_4627_ (
  .A1({ S24393 }),
  .A2({ S24416 }),
  .A3({ S24414 }),
  .ZN({ S24441 })
);
NAND3_X1 #() 
NAND3_X1_4628_ (
  .A1({ S24425 }),
  .A2({ S24438 }),
  .A3({ S25957[1123] }),
  .ZN({ S24442 })
);
NAND3_X1 #() 
NAND3_X1_4629_ (
  .A1({ S24442 }),
  .A2({ S24441 }),
  .A3({ S25957[1187] }),
  .ZN({ S24443 })
);
NAND3_X1 #() 
NAND3_X1_4630_ (
  .A1({ S24440 }),
  .A2({ S24443 }),
  .A3({ S80 }),
  .ZN({ S24444 })
);
NAND2_X1 #() 
NAND2_X1_4266_ (
  .A1({ S21828 }),
  .A2({ S21832 }),
  .ZN({ S24445 })
);
XNOR2_X1 #() 
XNOR2_X1_174_ (
  .A({ S24445 }),
  .B({ S25957[1187] }),
  .ZN({ S25957[1059] })
);
NAND3_X1 #() 
NAND3_X1_4631_ (
  .A1({ S24393 }),
  .A2({ S25957[1219] }),
  .A3({ S24414 }),
  .ZN({ S24446 })
);
NAND3_X1 #() 
NAND3_X1_4632_ (
  .A1({ S24425 }),
  .A2({ S24438 }),
  .A3({ S21829 }),
  .ZN({ S24447 })
);
NAND3_X1 #() 
NAND3_X1_4633_ (
  .A1({ S24447 }),
  .A2({ S24446 }),
  .A3({ S25957[1059] }),
  .ZN({ S24448 })
);
INV_X1 #() 
INV_X1_1397_ (
  .A({ S25957[1059] }),
  .ZN({ S24449 })
);
AOI21_X1 #() 
AOI21_X1_2308_ (
  .A({ S21829 }),
  .B1({ S24425 }),
  .B2({ S24438 }),
  .ZN({ S24450 })
);
AOI21_X1 #() 
AOI21_X1_2309_ (
  .A({ S25957[1219] }),
  .B1({ S24393 }),
  .B2({ S24414 }),
  .ZN({ S24451 })
);
OAI21_X1 #() 
OAI21_X1_2192_ (
  .A({ S24449 }),
  .B1({ S24450 }),
  .B2({ S24451 }),
  .ZN({ S24452 })
);
NAND3_X1 #() 
NAND3_X1_4634_ (
  .A1({ S24452 }),
  .A2({ S25957[1027] }),
  .A3({ S24448 }),
  .ZN({ S24453 })
);
NAND2_X1 #() 
NAND2_X1_4267_ (
  .A1({ S24453 }),
  .A2({ S24444 }),
  .ZN({ S92 })
);
NAND3_X1 #() 
NAND3_X1_4635_ (
  .A1({ S24452 }),
  .A2({ S80 }),
  .A3({ S24448 }),
  .ZN({ S24454 })
);
NAND3_X1 #() 
NAND3_X1_4636_ (
  .A1({ S24440 }),
  .A2({ S24443 }),
  .A3({ S25957[1027] }),
  .ZN({ S24455 })
);
NAND2_X1 #() 
NAND2_X1_4268_ (
  .A1({ S24454 }),
  .A2({ S24455 }),
  .ZN({ S25957[899] })
);
NOR2_X1 #() 
NOR2_X1_1088_ (
  .A1({ S19428 }),
  .A2({ S19429 }),
  .ZN({ S25957[1184] })
);
NAND2_X1 #() 
NAND2_X1_4269_ (
  .A1({ S21907 }),
  .A2({ S21908 }),
  .ZN({ S24456 })
);
XNOR2_X1 #() 
XNOR2_X1_175_ (
  .A({ S24456 }),
  .B({ S25957[1184] }),
  .ZN({ S25957[1056] })
);
INV_X1 #() 
INV_X1_1398_ (
  .A({ S25957[1056] }),
  .ZN({ S24457 })
);
NAND3_X1 #() 
NAND3_X1_4637_ (
  .A1({ S24049 }),
  .A2({ S83 }),
  .A3({ S24109 }),
  .ZN({ S24458 })
);
OAI211_X1 #() 
OAI211_X1_1482_ (
  .A({ S24458 }),
  .B({ S25957[1052] }),
  .C1({ S83 }),
  .C2({ S24251 }),
  .ZN({ S24459 })
);
NAND4_X1 #() 
NAND4_X1_498_ (
  .A1({ S24058 }),
  .A2({ S24047 }),
  .A3({ S83 }),
  .A4({ S91 }),
  .ZN({ S24460 })
);
NAND3_X1 #() 
NAND3_X1_4638_ (
  .A1({ S24460 }),
  .A2({ S24331 }),
  .A3({ S24046 }),
  .ZN({ S24461 })
);
NAND3_X1 #() 
NAND3_X1_4639_ (
  .A1({ S24459 }),
  .A2({ S24461 }),
  .A3({ S25957[1053] }),
  .ZN({ S24462 })
);
AOI21_X1 #() 
AOI21_X1_2310_ (
  .A({ S25957[1052] }),
  .B1({ S24225 }),
  .B2({ S24234 }),
  .ZN({ S24463 })
);
NAND3_X1 #() 
NAND3_X1_4640_ (
  .A1({ S25957[1050] }),
  .A2({ S24064 }),
  .A3({ S25957[1051] }),
  .ZN({ S24464 })
);
AOI21_X1 #() 
AOI21_X1_2311_ (
  .A({ S24046 }),
  .B1({ S24300 }),
  .B2({ S24464 }),
  .ZN({ S24465 })
);
OAI21_X1 #() 
OAI21_X1_2193_ (
  .A({ S22294 }),
  .B1({ S24465 }),
  .B2({ S24463 }),
  .ZN({ S24466 })
);
AOI21_X1 #() 
AOI21_X1_2312_ (
  .A({ S22219 }),
  .B1({ S24466 }),
  .B2({ S24462 }),
  .ZN({ S24467 })
);
AOI21_X1 #() 
AOI21_X1_2313_ (
  .A({ S83 }),
  .B1({ S24051 }),
  .B2({ S91 }),
  .ZN({ S24468 })
);
AOI21_X1 #() 
AOI21_X1_2314_ (
  .A({ S25957[1051] }),
  .B1({ S24053 }),
  .B2({ S24024 }),
  .ZN({ S24469 })
);
OAI21_X1 #() 
OAI21_X1_2194_ (
  .A({ S24046 }),
  .B1({ S24469 }),
  .B2({ S24468 }),
  .ZN({ S24470 })
);
OAI211_X1 #() 
OAI211_X1_1483_ (
  .A({ S24163 }),
  .B({ S25957[1052] }),
  .C1({ S25957[1051] }),
  .C2({ S24102 }),
  .ZN({ S24471 })
);
NAND3_X1 #() 
NAND3_X1_4641_ (
  .A1({ S24470 }),
  .A2({ S22294 }),
  .A3({ S24471 }),
  .ZN({ S24472 })
);
OAI211_X1 #() 
OAI211_X1_1484_ (
  .A({ S24123 }),
  .B({ S24303 }),
  .C1({ S24189 }),
  .C2({ S25957[1051] }),
  .ZN({ S24473 })
);
NAND2_X1 #() 
NAND2_X1_4270_ (
  .A1({ S24473 }),
  .A2({ S24046 }),
  .ZN({ S24474 })
);
NAND3_X1 #() 
NAND3_X1_4642_ (
  .A1({ S24198 }),
  .A2({ S24364 }),
  .A3({ S83 }),
  .ZN({ S24475 })
);
NOR2_X1 #() 
NOR2_X1_1089_ (
  .A1({ S24189 }),
  .A2({ S24046 }),
  .ZN({ S24476 })
);
NAND2_X1 #() 
NAND2_X1_4271_ (
  .A1({ S24475 }),
  .A2({ S24476 }),
  .ZN({ S24477 })
);
NAND3_X1 #() 
NAND3_X1_4643_ (
  .A1({ S24474 }),
  .A2({ S24477 }),
  .A3({ S25957[1053] }),
  .ZN({ S24478 })
);
AND3_X1 #() 
AND3_X1_168_ (
  .A1({ S24472 }),
  .A2({ S22219 }),
  .A3({ S24478 }),
  .ZN({ S24479 })
);
OAI21_X1 #() 
OAI21_X1_2195_ (
  .A({ S25957[1055] }),
  .B1({ S24467 }),
  .B2({ S24479 }),
  .ZN({ S24480 })
);
NOR2_X1 #() 
NOR2_X1_1090_ (
  .A1({ S24226 }),
  .A2({ S24112 }),
  .ZN({ S24481 })
);
NAND2_X1 #() 
NAND2_X1_4272_ (
  .A1({ S24233 }),
  .A2({ S25957[1051] }),
  .ZN({ S24482 })
);
OAI21_X1 #() 
OAI21_X1_2196_ (
  .A({ S25957[1052] }),
  .B1({ S24482 }),
  .B2({ S24241 }),
  .ZN({ S24483 })
);
NOR2_X1 #() 
NOR2_X1_1091_ (
  .A1({ S24483 }),
  .A2({ S24481 }),
  .ZN({ S24484 })
);
AOI21_X1 #() 
AOI21_X1_2315_ (
  .A({ S83 }),
  .B1({ S24053 }),
  .B2({ S24257 }),
  .ZN({ S24485 })
);
NAND2_X1 #() 
NAND2_X1_4273_ (
  .A1({ S24274 }),
  .A2({ S24046 }),
  .ZN({ S24486 })
);
NOR2_X1 #() 
NOR2_X1_1092_ (
  .A1({ S24485 }),
  .A2({ S24486 }),
  .ZN({ S24487 })
);
OAI21_X1 #() 
OAI21_X1_2197_ (
  .A({ S25957[1053] }),
  .B1({ S24484 }),
  .B2({ S24487 }),
  .ZN({ S24488 })
);
NAND3_X1 #() 
NAND3_X1_4644_ (
  .A1({ S24165 }),
  .A2({ S24074 }),
  .A3({ S24047 }),
  .ZN({ S24489 })
);
OAI211_X1 #() 
OAI211_X1_1485_ (
  .A({ S24489 }),
  .B({ S25957[1052] }),
  .C1({ S83 }),
  .C2({ S25957[1048] }),
  .ZN({ S24490 })
);
OAI211_X1 #() 
OAI211_X1_1486_ (
  .A({ S24490 }),
  .B({ S22294 }),
  .C1({ S24253 }),
  .C2({ S24344 }),
  .ZN({ S24491 })
);
NAND3_X1 #() 
NAND3_X1_4645_ (
  .A1({ S24488 }),
  .A2({ S24491 }),
  .A3({ S25957[1054] }),
  .ZN({ S24492 })
);
NAND2_X1 #() 
NAND2_X1_4274_ (
  .A1({ S24039 }),
  .A2({ S83 }),
  .ZN({ S24493 })
);
OAI211_X1 #() 
OAI211_X1_1487_ (
  .A({ S24370 }),
  .B({ S25957[1052] }),
  .C1({ S24096 }),
  .C2({ S24493 }),
  .ZN({ S24494 })
);
NAND3_X1 #() 
NAND3_X1_4646_ (
  .A1({ S24024 }),
  .A2({ S25957[1051] }),
  .A3({ S24064 }),
  .ZN({ S24495 })
);
OAI21_X1 #() 
OAI21_X1_2198_ (
  .A({ S83 }),
  .B1({ S24242 }),
  .B2({ S24189 }),
  .ZN({ S24496 })
);
NAND3_X1 #() 
NAND3_X1_4647_ (
  .A1({ S24496 }),
  .A2({ S24046 }),
  .A3({ S24495 }),
  .ZN({ S24497 })
);
NAND3_X1 #() 
NAND3_X1_4648_ (
  .A1({ S24497 }),
  .A2({ S24494 }),
  .A3({ S22294 }),
  .ZN({ S24498 })
);
NOR2_X1 #() 
NOR2_X1_1093_ (
  .A1({ S24099 }),
  .A2({ S24052 }),
  .ZN({ S24499 })
);
OR2_X1 #() 
OR2_X1_60_ (
  .A1({ S24328 }),
  .A2({ S24046 }),
  .ZN({ S24500 })
);
NAND3_X1 #() 
NAND3_X1_4649_ (
  .A1({ S24150 }),
  .A2({ S24046 }),
  .A3({ S24244 }),
  .ZN({ S24501 })
);
OAI211_X1 #() 
OAI211_X1_1488_ (
  .A({ S24501 }),
  .B({ S25957[1053] }),
  .C1({ S24500 }),
  .C2({ S24499 }),
  .ZN({ S24502 })
);
NAND3_X1 #() 
NAND3_X1_4650_ (
  .A1({ S24498 }),
  .A2({ S24502 }),
  .A3({ S22219 }),
  .ZN({ S24503 })
);
NAND3_X1 #() 
NAND3_X1_4651_ (
  .A1({ S24492 }),
  .A2({ S24503 }),
  .A3({ S22150 }),
  .ZN({ S24504 })
);
NAND3_X1 #() 
NAND3_X1_4652_ (
  .A1({ S24480 }),
  .A2({ S25957[1216] }),
  .A3({ S24504 }),
  .ZN({ S24505 })
);
NAND3_X1 #() 
NAND3_X1_4653_ (
  .A1({ S24470 }),
  .A2({ S22219 }),
  .A3({ S24471 }),
  .ZN({ S24506 })
);
OAI21_X1 #() 
OAI21_X1_2199_ (
  .A({ S24234 }),
  .B1({ S24175 }),
  .B2({ S24056 }),
  .ZN({ S24507 })
);
NAND2_X1 #() 
NAND2_X1_4275_ (
  .A1({ S24507 }),
  .A2({ S24046 }),
  .ZN({ S24508 })
);
AOI21_X1 #() 
AOI21_X1_2316_ (
  .A({ S25957[1051] }),
  .B1({ S24140 }),
  .B2({ S24257 }),
  .ZN({ S24509 })
);
INV_X1 #() 
INV_X1_1399_ (
  .A({ S24464 }),
  .ZN({ S24510 })
);
OAI21_X1 #() 
OAI21_X1_2200_ (
  .A({ S25957[1052] }),
  .B1({ S24509 }),
  .B2({ S24510 }),
  .ZN({ S24511 })
);
NAND3_X1 #() 
NAND3_X1_4654_ (
  .A1({ S24511 }),
  .A2({ S24508 }),
  .A3({ S25957[1054] }),
  .ZN({ S24512 })
);
AOI21_X1 #() 
AOI21_X1_2317_ (
  .A({ S22150 }),
  .B1({ S24512 }),
  .B2({ S24506 }),
  .ZN({ S24513 })
);
NAND3_X1 #() 
NAND3_X1_4655_ (
  .A1({ S24058 }),
  .A2({ S83 }),
  .A3({ S24219 }),
  .ZN({ S24514 })
);
NAND4_X1 #() 
NAND4_X1_499_ (
  .A1({ S24514 }),
  .A2({ S24024 }),
  .A3({ S24032 }),
  .A4({ S25957[1052] }),
  .ZN({ S24515 })
);
OAI21_X1 #() 
OAI21_X1_2201_ (
  .A({ S83 }),
  .B1({ S24075 }),
  .B2({ S25957[1049] }),
  .ZN({ S24516 })
);
AND2_X1 #() 
AND2_X1_268_ (
  .A1({ S24225 }),
  .A2({ S24516 }),
  .ZN({ S24517 })
);
OAI211_X1 #() 
OAI211_X1_1489_ (
  .A({ S24515 }),
  .B({ S25957[1054] }),
  .C1({ S24517 }),
  .C2({ S25957[1052] }),
  .ZN({ S24518 })
);
OAI21_X1 #() 
OAI21_X1_2202_ (
  .A({ S24370 }),
  .B1({ S24493 }),
  .B2({ S24096 }),
  .ZN({ S24519 })
);
NAND2_X1 #() 
NAND2_X1_4276_ (
  .A1({ S24519 }),
  .A2({ S25957[1052] }),
  .ZN({ S24520 })
);
NAND2_X1 #() 
NAND2_X1_4277_ (
  .A1({ S24162 }),
  .A2({ S25957[1051] }),
  .ZN({ S24521 })
);
OAI211_X1 #() 
OAI211_X1_1490_ (
  .A({ S24521 }),
  .B({ S24046 }),
  .C1({ S24199 }),
  .C2({ S24189 }),
  .ZN({ S24522 })
);
NAND3_X1 #() 
NAND3_X1_4656_ (
  .A1({ S24520 }),
  .A2({ S24522 }),
  .A3({ S22219 }),
  .ZN({ S24523 })
);
AOI21_X1 #() 
AOI21_X1_2318_ (
  .A({ S25957[1055] }),
  .B1({ S24518 }),
  .B2({ S24523 }),
  .ZN({ S24524 })
);
OAI21_X1 #() 
OAI21_X1_2203_ (
  .A({ S22294 }),
  .B1({ S24524 }),
  .B2({ S24513 }),
  .ZN({ S24525 })
);
NAND3_X1 #() 
NAND3_X1_4657_ (
  .A1({ S24474 }),
  .A2({ S24477 }),
  .A3({ S22219 }),
  .ZN({ S24526 })
);
NAND2_X1 #() 
NAND2_X1_4278_ (
  .A1({ S24460 }),
  .A2({ S24331 }),
  .ZN({ S24527 })
);
NAND2_X1 #() 
NAND2_X1_4279_ (
  .A1({ S24527 }),
  .A2({ S24046 }),
  .ZN({ S24528 })
);
NOR2_X1 #() 
NOR2_X1_1094_ (
  .A1({ S24251 }),
  .A2({ S83 }),
  .ZN({ S24529 })
);
OAI21_X1 #() 
OAI21_X1_2204_ (
  .A({ S25957[1052] }),
  .B1({ S24329 }),
  .B2({ S24529 }),
  .ZN({ S24530 })
);
NAND3_X1 #() 
NAND3_X1_4658_ (
  .A1({ S24528 }),
  .A2({ S24530 }),
  .A3({ S25957[1054] }),
  .ZN({ S24531 })
);
AOI21_X1 #() 
AOI21_X1_2319_ (
  .A({ S22150 }),
  .B1({ S24531 }),
  .B2({ S24526 }),
  .ZN({ S24532 })
);
OAI21_X1 #() 
OAI21_X1_2205_ (
  .A({ S25957[1052] }),
  .B1({ S24499 }),
  .B2({ S24328 }),
  .ZN({ S24533 })
);
NAND2_X1 #() 
NAND2_X1_4280_ (
  .A1({ S24150 }),
  .A2({ S24244 }),
  .ZN({ S24534 })
);
NAND2_X1 #() 
NAND2_X1_4281_ (
  .A1({ S24534 }),
  .A2({ S24046 }),
  .ZN({ S24535 })
);
NAND3_X1 #() 
NAND3_X1_4659_ (
  .A1({ S24535 }),
  .A2({ S24533 }),
  .A3({ S22219 }),
  .ZN({ S24536 })
);
OAI221_X1 #() 
OAI221_X1_123_ (
  .A({ S25957[1054] }),
  .B1({ S24485 }),
  .B2({ S24486 }),
  .C1({ S24483 }),
  .C2({ S24481 }),
  .ZN({ S24537 })
);
AOI21_X1 #() 
AOI21_X1_2320_ (
  .A({ S25957[1055] }),
  .B1({ S24536 }),
  .B2({ S24537 }),
  .ZN({ S24538 })
);
OAI21_X1 #() 
OAI21_X1_2206_ (
  .A({ S25957[1053] }),
  .B1({ S24532 }),
  .B2({ S24538 }),
  .ZN({ S24539 })
);
NAND3_X1 #() 
NAND3_X1_4660_ (
  .A1({ S24539 }),
  .A2({ S24525 }),
  .A3({ S21837 }),
  .ZN({ S24540 })
);
NAND3_X1 #() 
NAND3_X1_4661_ (
  .A1({ S24540 }),
  .A2({ S24505 }),
  .A3({ S24457 }),
  .ZN({ S24541 })
);
AOI21_X1 #() 
AOI21_X1_2321_ (
  .A({ S21837 }),
  .B1({ S24539 }),
  .B2({ S24525 }),
  .ZN({ S24542 })
);
AOI21_X1 #() 
AOI21_X1_2322_ (
  .A({ S25957[1216] }),
  .B1({ S24480 }),
  .B2({ S24504 }),
  .ZN({ S24543 })
);
OAI21_X1 #() 
OAI21_X1_2207_ (
  .A({ S25957[1056] }),
  .B1({ S24542 }),
  .B2({ S24543 }),
  .ZN({ S24544 })
);
NAND3_X1 #() 
NAND3_X1_4662_ (
  .A1({ S24544 }),
  .A2({ S25957[1024] }),
  .A3({ S24541 }),
  .ZN({ S24545 })
);
NAND2_X1 #() 
NAND2_X1_4282_ (
  .A1({ S21904 }),
  .A2({ S21903 }),
  .ZN({ S25957[1120] })
);
NAND2_X1 #() 
NAND2_X1_4283_ (
  .A1({ S24466 }),
  .A2({ S24462 }),
  .ZN({ S24546 })
);
AOI22_X1 #() 
AOI22_X1_485_ (
  .A1({ S24473 }),
  .A2({ S24046 }),
  .B1({ S24475 }),
  .B2({ S24476 }),
  .ZN({ S24547 })
);
AOI21_X1 #() 
AOI21_X1_2323_ (
  .A({ S25957[1054] }),
  .B1({ S24547 }),
  .B2({ S25957[1053] }),
  .ZN({ S24548 })
);
AOI22_X1 #() 
AOI22_X1_486_ (
  .A1({ S24546 }),
  .A2({ S25957[1054] }),
  .B1({ S24472 }),
  .B2({ S24548 }),
  .ZN({ S24549 })
);
OAI211_X1 #() 
OAI211_X1_1491_ (
  .A({ S25957[1120] }),
  .B({ S24504 }),
  .C1({ S24549 }),
  .C2({ S22150 }),
  .ZN({ S24550 })
);
INV_X1 #() 
INV_X1_1400_ (
  .A({ S25957[1120] }),
  .ZN({ S24551 })
);
NAND3_X1 #() 
NAND3_X1_4663_ (
  .A1({ S24539 }),
  .A2({ S24525 }),
  .A3({ S24551 }),
  .ZN({ S24552 })
);
NAND3_X1 #() 
NAND3_X1_4664_ (
  .A1({ S24552 }),
  .A2({ S24550 }),
  .A3({ S25957[1184] }),
  .ZN({ S24553 })
);
INV_X1 #() 
INV_X1_1401_ (
  .A({ S25957[1184] }),
  .ZN({ S24554 })
);
NAND3_X1 #() 
NAND3_X1_4665_ (
  .A1({ S24480 }),
  .A2({ S24551 }),
  .A3({ S24504 }),
  .ZN({ S24555 })
);
NAND3_X1 #() 
NAND3_X1_4666_ (
  .A1({ S24539 }),
  .A2({ S24525 }),
  .A3({ S25957[1120] }),
  .ZN({ S24556 })
);
NAND3_X1 #() 
NAND3_X1_4667_ (
  .A1({ S24556 }),
  .A2({ S24555 }),
  .A3({ S24554 }),
  .ZN({ S24557 })
);
NAND3_X1 #() 
NAND3_X1_4668_ (
  .A1({ S24557 }),
  .A2({ S24553 }),
  .A3({ S23360 }),
  .ZN({ S24558 })
);
NAND2_X1 #() 
NAND2_X1_4284_ (
  .A1({ S24545 }),
  .A2({ S24558 }),
  .ZN({ S25957[896] })
);
NAND2_X1 #() 
NAND2_X1_4285_ (
  .A1({ S21979 }),
  .A2({ S21980 }),
  .ZN({ S24559 })
);
INV_X1 #() 
INV_X1_1402_ (
  .A({ S24559 }),
  .ZN({ S25957[1089] })
);
NAND2_X1 #() 
NAND2_X1_4286_ (
  .A1({ S21976 }),
  .A2({ S21975 }),
  .ZN({ S25957[1121] })
);
INV_X1 #() 
INV_X1_1403_ (
  .A({ S25957[1121] }),
  .ZN({ S24560 })
);
NAND3_X1 #() 
NAND3_X1_4669_ (
  .A1({ S24264 }),
  .A2({ S25957[1051] }),
  .A3({ S24024 }),
  .ZN({ S24561 })
);
AOI21_X1 #() 
AOI21_X1_2324_ (
  .A({ S24046 }),
  .B1({ S24561 }),
  .B2({ S24054 }),
  .ZN({ S24562 })
);
NAND2_X1 #() 
NAND2_X1_4287_ (
  .A1({ S24257 }),
  .A2({ S25957[1051] }),
  .ZN({ S24563 })
);
AOI21_X1 #() 
AOI21_X1_2325_ (
  .A({ S25957[1052] }),
  .B1({ S24395 }),
  .B2({ S24563 }),
  .ZN({ S24564 })
);
OAI21_X1 #() 
OAI21_X1_2208_ (
  .A({ S25957[1053] }),
  .B1({ S24562 }),
  .B2({ S24564 }),
  .ZN({ S24565 })
);
OAI21_X1 #() 
OAI21_X1_2209_ (
  .A({ S83 }),
  .B1({ S24160 }),
  .B2({ S24070 }),
  .ZN({ S24566 })
);
NAND3_X1 #() 
NAND3_X1_4670_ (
  .A1({ S24036 }),
  .A2({ S24046 }),
  .A3({ S24566 }),
  .ZN({ S24567 })
);
AOI21_X1 #() 
AOI21_X1_2326_ (
  .A({ S25957[1053] }),
  .B1({ S24183 }),
  .B2({ S24514 }),
  .ZN({ S24568 })
);
NAND2_X1 #() 
NAND2_X1_4288_ (
  .A1({ S24567 }),
  .A2({ S24568 }),
  .ZN({ S24569 })
);
NAND3_X1 #() 
NAND3_X1_4671_ (
  .A1({ S24565 }),
  .A2({ S24569 }),
  .A3({ S22219 }),
  .ZN({ S24570 })
);
NAND2_X1 #() 
NAND2_X1_4289_ (
  .A1({ S24118 }),
  .A2({ S83 }),
  .ZN({ S24571 })
);
NAND3_X1 #() 
NAND3_X1_4672_ (
  .A1({ S24220 }),
  .A2({ S24571 }),
  .A3({ S25957[1052] }),
  .ZN({ S24572 })
);
NAND3_X1 #() 
NAND3_X1_4673_ (
  .A1({ S24237 }),
  .A2({ S83 }),
  .A3({ S24197 }),
  .ZN({ S24573 })
);
NAND3_X1 #() 
NAND3_X1_4674_ (
  .A1({ S24364 }),
  .A2({ S25957[1051] }),
  .A3({ S24032 }),
  .ZN({ S24574 })
);
NAND4_X1 #() 
NAND4_X1_500_ (
  .A1({ S24574 }),
  .A2({ S24573 }),
  .A3({ S24181 }),
  .A4({ S24046 }),
  .ZN({ S24575 })
);
NAND3_X1 #() 
NAND3_X1_4675_ (
  .A1({ S24572 }),
  .A2({ S24575 }),
  .A3({ S22294 }),
  .ZN({ S24576 })
);
NAND2_X1 #() 
NAND2_X1_4290_ (
  .A1({ S24033 }),
  .A2({ S83 }),
  .ZN({ S24577 })
);
NAND3_X1 #() 
NAND3_X1_4676_ (
  .A1({ S24577 }),
  .A2({ S24386 }),
  .A3({ S25957[1052] }),
  .ZN({ S24578 })
);
NAND3_X1 #() 
NAND3_X1_4677_ (
  .A1({ S24065 }),
  .A2({ S25957[1051] }),
  .A3({ S24233 }),
  .ZN({ S24579 })
);
AOI21_X1 #() 
AOI21_X1_2327_ (
  .A({ S25957[1052] }),
  .B1({ S24053 }),
  .B2({ S83 }),
  .ZN({ S24580 })
);
NAND2_X1 #() 
NAND2_X1_4291_ (
  .A1({ S24579 }),
  .A2({ S24580 }),
  .ZN({ S24581 })
);
NAND3_X1 #() 
NAND3_X1_4678_ (
  .A1({ S24581 }),
  .A2({ S24578 }),
  .A3({ S25957[1053] }),
  .ZN({ S24582 })
);
NAND3_X1 #() 
NAND3_X1_4679_ (
  .A1({ S24576 }),
  .A2({ S25957[1054] }),
  .A3({ S24582 }),
  .ZN({ S24583 })
);
NAND3_X1 #() 
NAND3_X1_4680_ (
  .A1({ S24570 }),
  .A2({ S25957[1055] }),
  .A3({ S24583 }),
  .ZN({ S24584 })
);
NAND3_X1 #() 
NAND3_X1_4681_ (
  .A1({ S24038 }),
  .A2({ S25957[1051] }),
  .A3({ S24064 }),
  .ZN({ S24585 })
);
NAND3_X1 #() 
NAND3_X1_4682_ (
  .A1({ S24049 }),
  .A2({ S83 }),
  .A3({ S24024 }),
  .ZN({ S24586 })
);
NAND3_X1 #() 
NAND3_X1_4683_ (
  .A1({ S24585 }),
  .A2({ S24586 }),
  .A3({ S25957[1052] }),
  .ZN({ S24587 })
);
NAND3_X1 #() 
NAND3_X1_4684_ (
  .A1({ S24364 }),
  .A2({ S24024 }),
  .A3({ S24039 }),
  .ZN({ S24588 })
);
AOI21_X1 #() 
AOI21_X1_2328_ (
  .A({ S22294 }),
  .B1({ S24588 }),
  .B2({ S24307 }),
  .ZN({ S24589 })
);
NAND2_X1 #() 
NAND2_X1_4292_ (
  .A1({ S24587 }),
  .A2({ S24589 }),
  .ZN({ S24590 })
);
AOI21_X1 #() 
AOI21_X1_2329_ (
  .A({ S25957[1051] }),
  .B1({ S24033 }),
  .B2({ S24109 }),
  .ZN({ S24591 })
);
OAI211_X1 #() 
OAI211_X1_1492_ (
  .A({ S24464 }),
  .B({ S24046 }),
  .C1({ S24099 }),
  .C2({ S24056 }),
  .ZN({ S24592 })
);
OAI211_X1 #() 
OAI211_X1_1493_ (
  .A({ S24592 }),
  .B({ S22294 }),
  .C1({ S24483 }),
  .C2({ S24591 }),
  .ZN({ S24593 })
);
NAND3_X1 #() 
NAND3_X1_4685_ (
  .A1({ S24593 }),
  .A2({ S24590 }),
  .A3({ S25957[1054] }),
  .ZN({ S24594 })
);
OAI21_X1 #() 
OAI21_X1_2210_ (
  .A({ S24046 }),
  .B1({ S25957[1050] }),
  .B2({ S24271 }),
  .ZN({ S24595 })
);
AOI21_X1 #() 
AOI21_X1_2330_ (
  .A({ S24595 }),
  .B1({ S24057 }),
  .B2({ S24041 }),
  .ZN({ S24596 })
);
AOI21_X1 #() 
AOI21_X1_2331_ (
  .A({ S24046 }),
  .B1({ S24365 }),
  .B2({ S24316 }),
  .ZN({ S24597 })
);
OAI21_X1 #() 
OAI21_X1_2211_ (
  .A({ S25957[1053] }),
  .B1({ S24597 }),
  .B2({ S24043 }),
  .ZN({ S24598 })
);
NAND2_X1 #() 
NAND2_X1_4293_ (
  .A1({ S24125 }),
  .A2({ S24271 }),
  .ZN({ S24599 })
);
OAI21_X1 #() 
OAI21_X1_2212_ (
  .A({ S22294 }),
  .B1({ S24373 }),
  .B2({ S24599 }),
  .ZN({ S24600 })
);
OAI211_X1 #() 
OAI211_X1_1494_ (
  .A({ S24598 }),
  .B({ S22219 }),
  .C1({ S24600 }),
  .C2({ S24596 }),
  .ZN({ S24601 })
);
NAND3_X1 #() 
NAND3_X1_4686_ (
  .A1({ S24601 }),
  .A2({ S22150 }),
  .A3({ S24594 }),
  .ZN({ S24602 })
);
NAND3_X1 #() 
NAND3_X1_4687_ (
  .A1({ S24602 }),
  .A2({ S24584 }),
  .A3({ S24560 }),
  .ZN({ S24603 })
);
NAND3_X1 #() 
NAND3_X1_4688_ (
  .A1({ S24593 }),
  .A2({ S24590 }),
  .A3({ S22150 }),
  .ZN({ S24604 })
);
NAND3_X1 #() 
NAND3_X1_4689_ (
  .A1({ S24576 }),
  .A2({ S25957[1055] }),
  .A3({ S24582 }),
  .ZN({ S24605 })
);
NAND2_X1 #() 
NAND2_X1_4294_ (
  .A1({ S24605 }),
  .A2({ S24604 }),
  .ZN({ S24606 })
);
NAND2_X1 #() 
NAND2_X1_4295_ (
  .A1({ S24606 }),
  .A2({ S25957[1054] }),
  .ZN({ S24607 })
);
NAND4_X1 #() 
NAND4_X1_501_ (
  .A1({ S22621 }),
  .A2({ S22627 }),
  .A3({ S83 }),
  .A4({ S24022 }),
  .ZN({ S24608 })
);
NAND3_X1 #() 
NAND3_X1_4690_ (
  .A1({ S24126 }),
  .A2({ S24182 }),
  .A3({ S24608 }),
  .ZN({ S24609 })
);
NAND2_X1 #() 
NAND2_X1_4296_ (
  .A1({ S24609 }),
  .A2({ S25957[1052] }),
  .ZN({ S24610 })
);
OAI21_X1 #() 
OAI21_X1_2213_ (
  .A({ S24046 }),
  .B1({ S24035 }),
  .B2({ S24306 }),
  .ZN({ S24611 })
);
NAND3_X1 #() 
NAND3_X1_4691_ (
  .A1({ S24611 }),
  .A2({ S24610 }),
  .A3({ S22294 }),
  .ZN({ S24612 })
);
AOI21_X1 #() 
AOI21_X1_2332_ (
  .A({ S25957[1051] }),
  .B1({ S25957[1050] }),
  .B2({ S24052 }),
  .ZN({ S24613 })
);
INV_X1 #() 
INV_X1_1404_ (
  .A({ S24175 }),
  .ZN({ S24614 })
);
AOI22_X1 #() 
AOI22_X1_487_ (
  .A1({ S24614 }),
  .A2({ S24264 }),
  .B1({ S24613 }),
  .B2({ S24051 }),
  .ZN({ S24615 })
);
NAND3_X1 #() 
NAND3_X1_4692_ (
  .A1({ S24165 }),
  .A2({ S83 }),
  .A3({ S91 }),
  .ZN({ S24616 })
);
AOI21_X1 #() 
AOI21_X1_2333_ (
  .A({ S22294 }),
  .B1({ S24161 }),
  .B2({ S24616 }),
  .ZN({ S24617 })
);
OAI21_X1 #() 
OAI21_X1_2214_ (
  .A({ S24617 }),
  .B1({ S24615 }),
  .B2({ S24046 }),
  .ZN({ S24618 })
);
AOI21_X1 #() 
AOI21_X1_2334_ (
  .A({ S22150 }),
  .B1({ S24612 }),
  .B2({ S24618 }),
  .ZN({ S24619 })
);
NOR2_X1 #() 
NOR2_X1_1095_ (
  .A1({ S24373 }),
  .A2({ S24599 }),
  .ZN({ S24620 })
);
OAI21_X1 #() 
OAI21_X1_2215_ (
  .A({ S22294 }),
  .B1({ S24620 }),
  .B2({ S24596 }),
  .ZN({ S24621 })
);
AND3_X1 #() 
AND3_X1_169_ (
  .A1({ S24039 }),
  .A2({ S24021 }),
  .A3({ S83 }),
  .ZN({ S24622 })
);
OAI21_X1 #() 
OAI21_X1_2216_ (
  .A({ S90 }),
  .B1({ S24031 }),
  .B2({ S24030 }),
  .ZN({ S24623 })
);
AOI21_X1 #() 
AOI21_X1_2335_ (
  .A({ S83 }),
  .B1({ S24623 }),
  .B2({ S24219 }),
  .ZN({ S24624 })
);
OAI21_X1 #() 
OAI21_X1_2217_ (
  .A({ S25957[1052] }),
  .B1({ S24624 }),
  .B2({ S24622 }),
  .ZN({ S24625 })
);
AOI21_X1 #() 
AOI21_X1_2336_ (
  .A({ S22294 }),
  .B1({ S24145 }),
  .B2({ S24046 }),
  .ZN({ S24626 })
);
NAND2_X1 #() 
NAND2_X1_4297_ (
  .A1({ S24626 }),
  .A2({ S24625 }),
  .ZN({ S24627 })
);
AOI21_X1 #() 
AOI21_X1_2337_ (
  .A({ S25957[1055] }),
  .B1({ S24621 }),
  .B2({ S24627 }),
  .ZN({ S24628 })
);
OAI21_X1 #() 
OAI21_X1_2218_ (
  .A({ S22219 }),
  .B1({ S24619 }),
  .B2({ S24628 }),
  .ZN({ S24629 })
);
NAND3_X1 #() 
NAND3_X1_4693_ (
  .A1({ S24629 }),
  .A2({ S24607 }),
  .A3({ S25957[1121] }),
  .ZN({ S24630 })
);
NAND3_X1 #() 
NAND3_X1_4694_ (
  .A1({ S24630 }),
  .A2({ S25957[1089] }),
  .A3({ S24603 }),
  .ZN({ S24631 })
);
NAND3_X1 #() 
NAND3_X1_4695_ (
  .A1({ S24602 }),
  .A2({ S24584 }),
  .A3({ S25957[1121] }),
  .ZN({ S24632 })
);
NAND3_X1 #() 
NAND3_X1_4696_ (
  .A1({ S24629 }),
  .A2({ S24607 }),
  .A3({ S24560 }),
  .ZN({ S24633 })
);
NAND3_X1 #() 
NAND3_X1_4697_ (
  .A1({ S24633 }),
  .A2({ S24559 }),
  .A3({ S24632 }),
  .ZN({ S24634 })
);
NAND3_X1 #() 
NAND3_X1_4698_ (
  .A1({ S24631 }),
  .A2({ S24634 }),
  .A3({ S25957[1153] }),
  .ZN({ S24635 })
);
NAND3_X1 #() 
NAND3_X1_4699_ (
  .A1({ S24633 }),
  .A2({ S25957[1089] }),
  .A3({ S24632 }),
  .ZN({ S24636 })
);
NAND3_X1 #() 
NAND3_X1_4700_ (
  .A1({ S24630 }),
  .A2({ S24559 }),
  .A3({ S24603 }),
  .ZN({ S24637 })
);
NAND3_X1 #() 
NAND3_X1_4701_ (
  .A1({ S24636 }),
  .A2({ S24637 }),
  .A3({ S20761 }),
  .ZN({ S24638 })
);
NAND2_X1 #() 
NAND2_X1_4298_ (
  .A1({ S24635 }),
  .A2({ S24638 }),
  .ZN({ S25957[897] })
);
NAND3_X1 #() 
NAND3_X1_4702_ (
  .A1({ S24251 }),
  .A2({ S24102 }),
  .A3({ S25957[1051] }),
  .ZN({ S24639 })
);
NAND3_X1 #() 
NAND3_X1_4703_ (
  .A1({ S24639 }),
  .A2({ S24046 }),
  .A3({ S24340 }),
  .ZN({ S24640 })
);
NAND3_X1 #() 
NAND3_X1_4704_ (
  .A1({ S24460 }),
  .A2({ S24040 }),
  .A3({ S25957[1052] }),
  .ZN({ S24641 })
);
NAND3_X1 #() 
NAND3_X1_4705_ (
  .A1({ S24641 }),
  .A2({ S25957[1053] }),
  .A3({ S24640 }),
  .ZN({ S24642 })
);
NAND3_X1 #() 
NAND3_X1_4706_ (
  .A1({ S24080 }),
  .A2({ S24046 }),
  .A3({ S24608 }),
  .ZN({ S24643 })
);
NOR3_X1 #() 
NOR3_X1_147_ (
  .A1({ S24103 }),
  .A2({ S24104 }),
  .A3({ S83 }),
  .ZN({ S24644 })
);
OAI211_X1 #() 
OAI211_X1_1495_ (
  .A({ S22294 }),
  .B({ S24643 }),
  .C1({ S24644 }),
  .C2({ S24268 }),
  .ZN({ S24645 })
);
NAND3_X1 #() 
NAND3_X1_4707_ (
  .A1({ S24642 }),
  .A2({ S24645 }),
  .A3({ S25957[1054] }),
  .ZN({ S24646 })
);
NAND3_X1 #() 
NAND3_X1_4708_ (
  .A1({ S24074 }),
  .A2({ S25957[1051] }),
  .A3({ S25957[1048] }),
  .ZN({ S24647 })
);
AOI21_X1 #() 
AOI21_X1_2338_ (
  .A({ S24046 }),
  .B1({ S24401 }),
  .B2({ S24647 }),
  .ZN({ S24648 })
);
NAND3_X1 #() 
NAND3_X1_4709_ (
  .A1({ S24074 }),
  .A2({ S24027 }),
  .A3({ S25957[1051] }),
  .ZN({ S24649 })
);
INV_X1 #() 
INV_X1_1405_ (
  .A({ S24649 }),
  .ZN({ S24650 })
);
NAND2_X1 #() 
NAND2_X1_4299_ (
  .A1({ S24151 }),
  .A2({ S24046 }),
  .ZN({ S24651 })
);
NOR2_X1 #() 
NOR2_X1_1096_ (
  .A1({ S24650 }),
  .A2({ S24651 }),
  .ZN({ S24652 })
);
OAI21_X1 #() 
OAI21_X1_2219_ (
  .A({ S25957[1053] }),
  .B1({ S24652 }),
  .B2({ S24648 }),
  .ZN({ S24653 })
);
NAND3_X1 #() 
NAND3_X1_4710_ (
  .A1({ S24237 }),
  .A2({ S83 }),
  .A3({ S24052 }),
  .ZN({ S24654 })
);
AOI21_X1 #() 
AOI21_X1_2339_ (
  .A({ S25957[1052] }),
  .B1({ S24654 }),
  .B2({ S24163 }),
  .ZN({ S24655 })
);
NAND3_X1 #() 
NAND3_X1_4711_ (
  .A1({ S24024 }),
  .A2({ S25957[1051] }),
  .A3({ S25957[1049] }),
  .ZN({ S24656 })
);
AOI21_X1 #() 
AOI21_X1_2340_ (
  .A({ S24046 }),
  .B1({ S24656 }),
  .B2({ S24493 }),
  .ZN({ S24657 })
);
OAI21_X1 #() 
OAI21_X1_2220_ (
  .A({ S22294 }),
  .B1({ S24655 }),
  .B2({ S24657 }),
  .ZN({ S24658 })
);
NAND3_X1 #() 
NAND3_X1_4712_ (
  .A1({ S24653 }),
  .A2({ S22219 }),
  .A3({ S24658 }),
  .ZN({ S24659 })
);
NAND3_X1 #() 
NAND3_X1_4713_ (
  .A1({ S24659 }),
  .A2({ S24646 }),
  .A3({ S25957[1055] }),
  .ZN({ S24660 })
);
NAND3_X1 #() 
NAND3_X1_4714_ (
  .A1({ S24074 }),
  .A2({ S25957[1051] }),
  .A3({ S24025 }),
  .ZN({ S24661 })
);
OAI21_X1 #() 
OAI21_X1_2221_ (
  .A({ S24661 }),
  .B1({ S24075 }),
  .B2({ S24398 }),
  .ZN({ S24662 })
);
AOI21_X1 #() 
AOI21_X1_2341_ (
  .A({ S25957[1052] }),
  .B1({ S24319 }),
  .B2({ S24041 }),
  .ZN({ S24663 })
);
AOI22_X1 #() 
AOI22_X1_488_ (
  .A1({ S24663 }),
  .A2({ S24098 }),
  .B1({ S24662 }),
  .B2({ S25957[1052] }),
  .ZN({ S24664 })
);
NOR2_X1 #() 
NOR2_X1_1097_ (
  .A1({ S24237 }),
  .A2({ S24025 }),
  .ZN({ S24665 })
);
NAND3_X1 #() 
NAND3_X1_4715_ (
  .A1({ S24038 }),
  .A2({ S25957[1051] }),
  .A3({ S24219 }),
  .ZN({ S24666 })
);
OAI211_X1 #() 
OAI211_X1_1496_ (
  .A({ S24666 }),
  .B({ S25957[1052] }),
  .C1({ S24665 }),
  .C2({ S24262 }),
  .ZN({ S24667 })
);
NAND3_X1 #() 
NAND3_X1_4716_ (
  .A1({ S24165 }),
  .A2({ S25957[1051] }),
  .A3({ S24219 }),
  .ZN({ S24668 })
);
NAND3_X1 #() 
NAND3_X1_4717_ (
  .A1({ S24300 }),
  .A2({ S24046 }),
  .A3({ S24668 }),
  .ZN({ S24669 })
);
NAND3_X1 #() 
NAND3_X1_4718_ (
  .A1({ S24667 }),
  .A2({ S24669 }),
  .A3({ S22294 }),
  .ZN({ S24670 })
);
OAI211_X1 #() 
OAI211_X1_1497_ (
  .A({ S24670 }),
  .B({ S25957[1054] }),
  .C1({ S24664 }),
  .C2({ S22294 }),
  .ZN({ S24671 })
);
NAND3_X1 #() 
NAND3_X1_4719_ (
  .A1({ S24038 }),
  .A2({ S24090 }),
  .A3({ S25957[1051] }),
  .ZN({ S24672 })
);
NAND3_X1 #() 
NAND3_X1_4720_ (
  .A1({ S24366 }),
  .A2({ S24672 }),
  .A3({ S25957[1052] }),
  .ZN({ S24673 })
);
NAND3_X1 #() 
NAND3_X1_4721_ (
  .A1({ S24623 }),
  .A2({ S25957[1051] }),
  .A3({ S24233 }),
  .ZN({ S24674 })
);
NAND3_X1 #() 
NAND3_X1_4722_ (
  .A1({ S24674 }),
  .A2({ S24046 }),
  .A3({ S24654 }),
  .ZN({ S24675 })
);
NAND3_X1 #() 
NAND3_X1_4723_ (
  .A1({ S24673 }),
  .A2({ S24675 }),
  .A3({ S25957[1053] }),
  .ZN({ S24676 })
);
AOI21_X1 #() 
AOI21_X1_2342_ (
  .A({ S24046 }),
  .B1({ S24310 }),
  .B2({ S24656 }),
  .ZN({ S24677 })
);
NAND4_X1 #() 
NAND4_X1_502_ (
  .A1({ S24165 }),
  .A2({ S24102 }),
  .A3({ S24046 }),
  .A4({ S83 }),
  .ZN({ S24678 })
);
NAND2_X1 #() 
NAND2_X1_4300_ (
  .A1({ S24201 }),
  .A2({ S24678 }),
  .ZN({ S24679 })
);
OAI21_X1 #() 
OAI21_X1_2222_ (
  .A({ S22294 }),
  .B1({ S24679 }),
  .B2({ S24677 }),
  .ZN({ S24680 })
);
NAND3_X1 #() 
NAND3_X1_4724_ (
  .A1({ S24680 }),
  .A2({ S24676 }),
  .A3({ S22219 }),
  .ZN({ S24681 })
);
NAND3_X1 #() 
NAND3_X1_4725_ (
  .A1({ S24671 }),
  .A2({ S24681 }),
  .A3({ S22150 }),
  .ZN({ S24682 })
);
NAND3_X1 #() 
NAND3_X1_4726_ (
  .A1({ S24682 }),
  .A2({ S25957[1218] }),
  .A3({ S24660 }),
  .ZN({ S24683 })
);
OAI21_X1 #() 
OAI21_X1_2223_ (
  .A({ S24643 }),
  .B1({ S24644 }),
  .B2({ S24268 }),
  .ZN({ S24684 })
);
NAND2_X1 #() 
NAND2_X1_4301_ (
  .A1({ S24684 }),
  .A2({ S22294 }),
  .ZN({ S24685 })
);
AOI21_X1 #() 
AOI21_X1_2343_ (
  .A({ S83 }),
  .B1({ S24364 }),
  .B2({ S24074 }),
  .ZN({ S24686 })
);
AOI21_X1 #() 
AOI21_X1_2344_ (
  .A({ S25957[1051] }),
  .B1({ S24165 }),
  .B2({ S24102 }),
  .ZN({ S24687 })
);
OAI21_X1 #() 
OAI21_X1_2224_ (
  .A({ S25957[1052] }),
  .B1({ S24687 }),
  .B2({ S24686 }),
  .ZN({ S24688 })
);
NAND2_X1 #() 
NAND2_X1_4302_ (
  .A1({ S24639 }),
  .A2({ S24340 }),
  .ZN({ S24689 })
);
NAND2_X1 #() 
NAND2_X1_4303_ (
  .A1({ S24689 }),
  .A2({ S24046 }),
  .ZN({ S24690 })
);
NAND3_X1 #() 
NAND3_X1_4727_ (
  .A1({ S24690 }),
  .A2({ S24688 }),
  .A3({ S25957[1053] }),
  .ZN({ S24691 })
);
NAND3_X1 #() 
NAND3_X1_4728_ (
  .A1({ S24685 }),
  .A2({ S24691 }),
  .A3({ S25957[1054] }),
  .ZN({ S24692 })
);
NAND3_X1 #() 
NAND3_X1_4729_ (
  .A1({ S24668 }),
  .A2({ S25957[1052] }),
  .A3({ S24372 }),
  .ZN({ S24693 })
);
OAI211_X1 #() 
OAI211_X1_1498_ (
  .A({ S24693 }),
  .B({ S22294 }),
  .C1({ S24168 }),
  .C2({ S25957[1052] }),
  .ZN({ S24694 })
);
OAI21_X1 #() 
OAI21_X1_2225_ (
  .A({ S25957[1053] }),
  .B1({ S24650 }),
  .B2({ S24651 }),
  .ZN({ S24695 })
);
OAI211_X1 #() 
OAI211_X1_1499_ (
  .A({ S24694 }),
  .B({ S22219 }),
  .C1({ S24648 }),
  .C2({ S24695 }),
  .ZN({ S24696 })
);
NAND3_X1 #() 
NAND3_X1_4730_ (
  .A1({ S24692 }),
  .A2({ S24696 }),
  .A3({ S25957[1055] }),
  .ZN({ S24697 })
);
NAND2_X1 #() 
NAND2_X1_4304_ (
  .A1({ S24319 }),
  .A2({ S24041 }),
  .ZN({ S24698 })
);
NAND3_X1 #() 
NAND3_X1_4731_ (
  .A1({ S24098 }),
  .A2({ S24698 }),
  .A3({ S25957[1053] }),
  .ZN({ S24699 })
);
AOI21_X1 #() 
AOI21_X1_2345_ (
  .A({ S83 }),
  .B1({ S24024 }),
  .B2({ S25957[1049] }),
  .ZN({ S24700 })
);
OAI21_X1 #() 
OAI21_X1_2226_ (
  .A({ S22294 }),
  .B1({ S24509 }),
  .B2({ S24700 }),
  .ZN({ S24701 })
);
NAND3_X1 #() 
NAND3_X1_4732_ (
  .A1({ S24699 }),
  .A2({ S24046 }),
  .A3({ S24701 }),
  .ZN({ S24702 })
);
NOR2_X1 #() 
NOR2_X1_1098_ (
  .A1({ S24665 }),
  .A2({ S24262 }),
  .ZN({ S24703 })
);
AOI21_X1 #() 
AOI21_X1_2346_ (
  .A({ S83 }),
  .B1({ S24364 }),
  .B2({ S24257 }),
  .ZN({ S24704 })
);
OAI21_X1 #() 
OAI21_X1_2227_ (
  .A({ S22294 }),
  .B1({ S24703 }),
  .B2({ S24704 }),
  .ZN({ S24705 })
);
OAI21_X1 #() 
OAI21_X1_2228_ (
  .A({ S24101 }),
  .B1({ S24075 }),
  .B2({ S24398 }),
  .ZN({ S24706 })
);
NOR2_X1 #() 
NOR2_X1_1099_ (
  .A1({ S22294 }),
  .A2({ S24110 }),
  .ZN({ S24707 })
);
AOI21_X1 #() 
AOI21_X1_2347_ (
  .A({ S24046 }),
  .B1({ S24707 }),
  .B2({ S24706 }),
  .ZN({ S24708 })
);
NAND2_X1 #() 
NAND2_X1_4305_ (
  .A1({ S24705 }),
  .A2({ S24708 }),
  .ZN({ S24709 })
);
NAND3_X1 #() 
NAND3_X1_4733_ (
  .A1({ S24702 }),
  .A2({ S24709 }),
  .A3({ S25957[1054] }),
  .ZN({ S24710 })
);
AOI21_X1 #() 
AOI21_X1_2348_ (
  .A({ S25957[1053] }),
  .B1({ S24485 }),
  .B2({ S24046 }),
  .ZN({ S24711 })
);
NAND2_X1 #() 
NAND2_X1_4306_ (
  .A1({ S24310 }),
  .A2({ S24656 }),
  .ZN({ S24712 })
);
NAND2_X1 #() 
NAND2_X1_4307_ (
  .A1({ S24712 }),
  .A2({ S25957[1052] }),
  .ZN({ S24713 })
);
NAND3_X1 #() 
NAND3_X1_4734_ (
  .A1({ S24713 }),
  .A2({ S24711 }),
  .A3({ S24678 }),
  .ZN({ S24714 })
);
AOI21_X1 #() 
AOI21_X1_2349_ (
  .A({ S25957[1052] }),
  .B1({ S24674 }),
  .B2({ S24654 }),
  .ZN({ S24715 })
);
AOI22_X1 #() 
AOI22_X1_489_ (
  .A1({ S24588 }),
  .A2({ S25957[1051] }),
  .B1({ S24028 }),
  .B2({ S24074 }),
  .ZN({ S24716 })
);
OAI21_X1 #() 
OAI21_X1_2229_ (
  .A({ S25957[1053] }),
  .B1({ S24716 }),
  .B2({ S24046 }),
  .ZN({ S24717 })
);
OAI211_X1 #() 
OAI211_X1_1500_ (
  .A({ S24714 }),
  .B({ S22219 }),
  .C1({ S24717 }),
  .C2({ S24715 }),
  .ZN({ S24718 })
);
NAND3_X1 #() 
NAND3_X1_4735_ (
  .A1({ S24718 }),
  .A2({ S24710 }),
  .A3({ S22150 }),
  .ZN({ S24719 })
);
NAND3_X1 #() 
NAND3_X1_4736_ (
  .A1({ S24719 }),
  .A2({ S24697 }),
  .A3({ S19534 }),
  .ZN({ S24720 })
);
AOI21_X1 #() 
AOI21_X1_2350_ (
  .A({ S25957[1154] }),
  .B1({ S24720 }),
  .B2({ S24683 }),
  .ZN({ S24721 })
);
AND3_X1 #() 
AND3_X1_170_ (
  .A1({ S24720 }),
  .A2({ S24683 }),
  .A3({ S25957[1154] }),
  .ZN({ S24722 })
);
NOR2_X1 #() 
NOR2_X1_1100_ (
  .A1({ S24722 }),
  .A2({ S24721 }),
  .ZN({ S25957[898] })
);
NAND3_X1 #() 
NAND3_X1_4737_ (
  .A1({ S23261 }),
  .A2({ S25957[1040] }),
  .A3({ S23262 }),
  .ZN({ S24723 })
);
INV_X1 #() 
INV_X1_1406_ (
  .A({ S24723 }),
  .ZN({ S93 })
);
NAND3_X1 #() 
NAND3_X1_4738_ (
  .A1({ S20675 }),
  .A2({ S23195 }),
  .A3({ S20679 }),
  .ZN({ S94 })
);
XNOR2_X1 #() 
XNOR2_X1_176_ (
  .A({ S22148 }),
  .B({ S25957[1215] }),
  .ZN({ S25957[1087] })
);
NAND3_X1 #() 
NAND3_X1_4739_ (
  .A1({ S23261 }),
  .A2({ S23262 }),
  .A3({ S25957[1042] }),
  .ZN({ S24724 })
);
AOI21_X1 #() 
AOI21_X1_2351_ (
  .A({ S25957[1170] }),
  .B1({ S20753 }),
  .B2({ S20754 }),
  .ZN({ S24725 })
);
AND3_X1 #() 
AND3_X1_171_ (
  .A1({ S20754 }),
  .A2({ S20753 }),
  .A3({ S25957[1170] }),
  .ZN({ S24726 })
);
NOR2_X1 #() 
NOR2_X1_1101_ (
  .A1({ S24726 }),
  .A2({ S24725 }),
  .ZN({ S24727 })
);
NAND3_X1 #() 
NAND3_X1_4740_ (
  .A1({ S94 }),
  .A2({ S24723 }),
  .A3({ S24727 }),
  .ZN({ S24728 })
);
AOI21_X1 #() 
AOI21_X1_2352_ (
  .A({ S25957[1043] }),
  .B1({ S24728 }),
  .B2({ S24724 }),
  .ZN({ S24729 })
);
AOI21_X1 #() 
AOI21_X1_2353_ (
  .A({ S25957[1042] }),
  .B1({ S23261 }),
  .B2({ S23262 }),
  .ZN({ S24730 })
);
NAND2_X1 #() 
NAND2_X1_4308_ (
  .A1({ S24730 }),
  .A2({ S25957[1043] }),
  .ZN({ S24731 })
);
NAND2_X1 #() 
NAND2_X1_4309_ (
  .A1({ S23195 }),
  .A2({ S25957[1042] }),
  .ZN({ S24732 })
);
NAND2_X1 #() 
NAND2_X1_4310_ (
  .A1({ S24732 }),
  .A2({ S74 }),
  .ZN({ S24733 })
);
AOI211_X1 #() 
AOI211_X1_70_ (
  .A({ S25957[1044] }),
  .B({ S24729 }),
  .C1({ S24731 }),
  .C2({ S24733 }),
  .ZN({ S24734 })
);
AOI22_X1 #() 
AOI22_X1_490_ (
  .A1({ S20619 }),
  .A2({ S20613 }),
  .B1({ S20752 }),
  .B2({ S20755 }),
  .ZN({ S24735 })
);
NAND2_X1 #() 
NAND2_X1_4311_ (
  .A1({ S25957[1041] }),
  .A2({ S74 }),
  .ZN({ S24736 })
);
OAI21_X1 #() 
OAI21_X1_2230_ (
  .A({ S25957[1043] }),
  .B1({ S23263 }),
  .B2({ S24735 }),
  .ZN({ S24737 })
);
NAND2_X1 #() 
NAND2_X1_4312_ (
  .A1({ S24737 }),
  .A2({ S25957[1044] }),
  .ZN({ S24738 })
);
INV_X1 #() 
INV_X1_1407_ (
  .A({ S24738 }),
  .ZN({ S24739 })
);
OAI21_X1 #() 
OAI21_X1_2231_ (
  .A({ S24739 }),
  .B1({ S24735 }),
  .B2({ S24736 }),
  .ZN({ S24740 })
);
NAND4_X1 #() 
NAND4_X1_503_ (
  .A1({ S20613 }),
  .A2({ S20752 }),
  .A3({ S20619 }),
  .A4({ S20755 }),
  .ZN({ S24741 })
);
NAND2_X1 #() 
NAND2_X1_4313_ (
  .A1({ S74 }),
  .A2({ S24741 }),
  .ZN({ S24742 })
);
OAI211_X1 #() 
OAI211_X1_1501_ (
  .A({ S24736 }),
  .B({ S24742 }),
  .C1({ S24723 }),
  .C2({ S74 }),
  .ZN({ S24743 })
);
OAI211_X1 #() 
OAI211_X1_1502_ (
  .A({ S24740 }),
  .B({ S25957[1045] }),
  .C1({ S25957[1044] }),
  .C2({ S24743 }),
  .ZN({ S24744 })
);
NAND3_X1 #() 
NAND3_X1_4741_ (
  .A1({ S94 }),
  .A2({ S24723 }),
  .A3({ S25957[1042] }),
  .ZN({ S24745 })
);
NAND3_X1 #() 
NAND3_X1_4742_ (
  .A1({ S23261 }),
  .A2({ S23195 }),
  .A3({ S23262 }),
  .ZN({ S24746 })
);
NAND3_X1 #() 
NAND3_X1_4743_ (
  .A1({ S20675 }),
  .A2({ S25957[1040] }),
  .A3({ S20679 }),
  .ZN({ S24747 })
);
NAND3_X1 #() 
NAND3_X1_4744_ (
  .A1({ S24746 }),
  .A2({ S24747 }),
  .A3({ S24727 }),
  .ZN({ S24748 })
);
AOI21_X1 #() 
AOI21_X1_2354_ (
  .A({ S74 }),
  .B1({ S24745 }),
  .B2({ S24748 }),
  .ZN({ S24749 })
);
INV_X1 #() 
INV_X1_1408_ (
  .A({ S24724 }),
  .ZN({ S24750 })
);
AOI22_X1 #() 
AOI22_X1_491_ (
  .A1({ S24727 }),
  .A2({ S25957[1040] }),
  .B1({ S20549 }),
  .B2({ S20546 }),
  .ZN({ S24751 })
);
INV_X1 #() 
INV_X1_1409_ (
  .A({ S24751 }),
  .ZN({ S24752 })
);
OAI21_X1 #() 
OAI21_X1_2232_ (
  .A({ S25957[1044] }),
  .B1({ S24752 }),
  .B2({ S24750 }),
  .ZN({ S24753 })
);
OAI21_X1 #() 
OAI21_X1_2233_ (
  .A({ S22921 }),
  .B1({ S24749 }),
  .B2({ S24753 }),
  .ZN({ S24754 })
);
OAI211_X1 #() 
OAI211_X1_1503_ (
  .A({ S24744 }),
  .B({ S22832 }),
  .C1({ S24734 }),
  .C2({ S24754 }),
  .ZN({ S24755 })
);
INV_X1 #() 
INV_X1_1410_ (
  .A({ S24746 }),
  .ZN({ S24756 })
);
AOI21_X1 #() 
AOI21_X1_2355_ (
  .A({ S74 }),
  .B1({ S23263 }),
  .B2({ S25957[1042] }),
  .ZN({ S24757 })
);
NAND2_X1 #() 
NAND2_X1_4314_ (
  .A1({ S24757 }),
  .A2({ S24723 }),
  .ZN({ S24758 })
);
OAI21_X1 #() 
OAI21_X1_2234_ (
  .A({ S24758 }),
  .B1({ S25957[1043] }),
  .B2({ S24756 }),
  .ZN({ S24759 })
);
NAND4_X1 #() 
NAND4_X1_504_ (
  .A1({ S20675 }),
  .A2({ S23195 }),
  .A3({ S20679 }),
  .A4({ S25957[1042] }),
  .ZN({ S24760 })
);
NAND3_X1 #() 
NAND3_X1_4745_ (
  .A1({ S23261 }),
  .A2({ S24727 }),
  .A3({ S23262 }),
  .ZN({ S24761 })
);
NAND2_X1 #() 
NAND2_X1_4315_ (
  .A1({ S24727 }),
  .A2({ S25957[1040] }),
  .ZN({ S24762 })
);
NAND3_X1 #() 
NAND3_X1_4746_ (
  .A1({ S24760 }),
  .A2({ S24761 }),
  .A3({ S24762 }),
  .ZN({ S24763 })
);
INV_X1 #() 
INV_X1_1411_ (
  .A({ S24747 }),
  .ZN({ S24764 })
);
AOI21_X1 #() 
AOI21_X1_2356_ (
  .A({ S25957[1044] }),
  .B1({ S24764 }),
  .B2({ S25957[1043] }),
  .ZN({ S24765 })
);
AOI22_X1 #() 
AOI22_X1_492_ (
  .A1({ S24759 }),
  .A2({ S25957[1044] }),
  .B1({ S24763 }),
  .B2({ S24765 }),
  .ZN({ S24766 })
);
NOR2_X1 #() 
NOR2_X1_1102_ (
  .A1({ S24727 }),
  .A2({ S25957[1040] }),
  .ZN({ S24767 })
);
NOR2_X1 #() 
NOR2_X1_1103_ (
  .A1({ S24767 }),
  .A2({ S74 }),
  .ZN({ S24768 })
);
NAND4_X1 #() 
NAND4_X1_505_ (
  .A1({ S20675 }),
  .A2({ S24727 }),
  .A3({ S25957[1040] }),
  .A4({ S20679 }),
  .ZN({ S24769 })
);
NAND2_X1 #() 
NAND2_X1_4316_ (
  .A1({ S24768 }),
  .A2({ S24769 }),
  .ZN({ S24770 })
);
OAI211_X1 #() 
OAI211_X1_1504_ (
  .A({ S24770 }),
  .B({ S25957[1044] }),
  .C1({ S23263 }),
  .C2({ S24742 }),
  .ZN({ S24771 })
);
NAND4_X1 #() 
NAND4_X1_506_ (
  .A1({ S23261 }),
  .A2({ S23195 }),
  .A3({ S23262 }),
  .A4({ S25957[1042] }),
  .ZN({ S24772 })
);
AOI21_X1 #() 
AOI21_X1_2357_ (
  .A({ S74 }),
  .B1({ S24772 }),
  .B2({ S24747 }),
  .ZN({ S24773 })
);
OAI21_X1 #() 
OAI21_X1_2235_ (
  .A({ S9119 }),
  .B1({ S20466 }),
  .B2({ S20465 }),
  .ZN({ S24774 })
);
NAND3_X1 #() 
NAND3_X1_4747_ (
  .A1({ S20471 }),
  .A2({ S25957[1172] }),
  .A3({ S20472 }),
  .ZN({ S24775 })
);
NAND2_X1 #() 
NAND2_X1_4317_ (
  .A1({ S24774 }),
  .A2({ S24775 }),
  .ZN({ S24776 })
);
NAND3_X1 #() 
NAND3_X1_4748_ (
  .A1({ S20675 }),
  .A2({ S24727 }),
  .A3({ S20679 }),
  .ZN({ S24777 })
);
NAND2_X1 #() 
NAND2_X1_4318_ (
  .A1({ S24777 }),
  .A2({ S24747 }),
  .ZN({ S24778 })
);
INV_X1 #() 
INV_X1_1412_ (
  .A({ S24778 }),
  .ZN({ S24779 })
);
OAI211_X1 #() 
OAI211_X1_1505_ (
  .A({ S23262 }),
  .B({ S23261 }),
  .C1({ S23195 }),
  .C2({ S25957[1042] }),
  .ZN({ S24780 })
);
NAND2_X1 #() 
NAND2_X1_4319_ (
  .A1({ S24779 }),
  .A2({ S24780 }),
  .ZN({ S24781 })
);
OAI21_X1 #() 
OAI21_X1_2236_ (
  .A({ S24776 }),
  .B1({ S24781 }),
  .B2({ S25957[1043] }),
  .ZN({ S24782 })
);
OAI211_X1 #() 
OAI211_X1_1506_ (
  .A({ S25957[1045] }),
  .B({ S24771 }),
  .C1({ S24782 }),
  .C2({ S24773 }),
  .ZN({ S24783 })
);
OAI211_X1 #() 
OAI211_X1_1507_ (
  .A({ S24783 }),
  .B({ S25957[1046] }),
  .C1({ S24766 }),
  .C2({ S25957[1045] }),
  .ZN({ S24784 })
);
NAND3_X1 #() 
NAND3_X1_4749_ (
  .A1({ S24784 }),
  .A2({ S24755 }),
  .A3({ S25957[1047] }),
  .ZN({ S24785 })
);
INV_X1 #() 
INV_X1_1413_ (
  .A({ S24772 }),
  .ZN({ S24786 })
);
NOR2_X1 #() 
NOR2_X1_1104_ (
  .A1({ S24786 }),
  .A2({ S24742 }),
  .ZN({ S24787 })
);
AOI211_X1 #() 
AOI211_X1_71_ (
  .A({ S24776 }),
  .B({ S24787 }),
  .C1({ S24781 }),
  .C2({ S25957[1043] }),
  .ZN({ S24788 })
);
NAND3_X1 #() 
NAND3_X1_4750_ (
  .A1({ S24769 }),
  .A2({ S25957[1043] }),
  .A3({ S24724 }),
  .ZN({ S24789 })
);
NAND2_X1 #() 
NAND2_X1_4320_ (
  .A1({ S24723 }),
  .A2({ S25957[1042] }),
  .ZN({ S24790 })
);
INV_X1 #() 
INV_X1_1414_ (
  .A({ S24790 }),
  .ZN({ S24791 })
);
NAND2_X1 #() 
NAND2_X1_4321_ (
  .A1({ S24791 }),
  .A2({ S74 }),
  .ZN({ S24792 })
);
AOI21_X1 #() 
AOI21_X1_2358_ (
  .A({ S25957[1044] }),
  .B1({ S24792 }),
  .B2({ S24789 }),
  .ZN({ S24793 })
);
OAI21_X1 #() 
OAI21_X1_2237_ (
  .A({ S25957[1045] }),
  .B1({ S24788 }),
  .B2({ S24793 }),
  .ZN({ S24794 })
);
AOI21_X1 #() 
AOI21_X1_2359_ (
  .A({ S74 }),
  .B1({ S24748 }),
  .B2({ S24790 }),
  .ZN({ S24795 })
);
INV_X1 #() 
INV_X1_1415_ (
  .A({ S24741 }),
  .ZN({ S24796 })
);
NAND3_X1 #() 
NAND3_X1_4751_ (
  .A1({ S20675 }),
  .A2({ S20679 }),
  .A3({ S25957[1042] }),
  .ZN({ S24797 })
);
NAND2_X1 #() 
NAND2_X1_4322_ (
  .A1({ S25957[1040] }),
  .A2({ S25957[1042] }),
  .ZN({ S24798 })
);
AOI22_X1 #() 
AOI22_X1_493_ (
  .A1({ S24797 }),
  .A2({ S24798 }),
  .B1({ S23263 }),
  .B2({ S25957[1040] }),
  .ZN({ S24799 })
);
OAI21_X1 #() 
OAI21_X1_2238_ (
  .A({ S74 }),
  .B1({ S24799 }),
  .B2({ S24796 }),
  .ZN({ S24800 })
);
NAND2_X1 #() 
NAND2_X1_4323_ (
  .A1({ S24800 }),
  .A2({ S25957[1044] }),
  .ZN({ S24801 })
);
AOI21_X1 #() 
AOI21_X1_2360_ (
  .A({ S74 }),
  .B1({ S24777 }),
  .B2({ S24732 }),
  .ZN({ S24802 })
);
NAND4_X1 #() 
NAND4_X1_507_ (
  .A1({ S24761 }),
  .A2({ S24797 }),
  .A3({ S24732 }),
  .A4({ S24741 }),
  .ZN({ S24803 })
);
AOI21_X1 #() 
AOI21_X1_2361_ (
  .A({ S25957[1044] }),
  .B1({ S24803 }),
  .B2({ S74 }),
  .ZN({ S24804 })
);
INV_X1 #() 
INV_X1_1416_ (
  .A({ S24804 }),
  .ZN({ S24805 })
);
OAI221_X1 #() 
OAI221_X1_124_ (
  .A({ S22921 }),
  .B1({ S24805 }),
  .B2({ S24802 }),
  .C1({ S24801 }),
  .C2({ S24795 }),
  .ZN({ S24806 })
);
AOI21_X1 #() 
AOI21_X1_2362_ (
  .A({ S22832 }),
  .B1({ S24794 }),
  .B2({ S24806 }),
  .ZN({ S24807 })
);
NOR2_X1 #() 
NOR2_X1_1105_ (
  .A1({ S24735 }),
  .A2({ S74 }),
  .ZN({ S24808 })
);
AOI22_X1 #() 
AOI22_X1_494_ (
  .A1({ S20549 }),
  .A2({ S20546 }),
  .B1({ S20613 }),
  .B2({ S20619 }),
  .ZN({ S24809 })
);
AOI211_X1 #() 
AOI211_X1_72_ (
  .A({ S24809 }),
  .B({ S24776 }),
  .C1({ S24808 }),
  .C2({ S24777 }),
  .ZN({ S24810 })
);
NAND2_X1 #() 
NAND2_X1_4324_ (
  .A1({ S24777 }),
  .A2({ S24741 }),
  .ZN({ S24811 })
);
NAND2_X1 #() 
NAND2_X1_4325_ (
  .A1({ S24724 }),
  .A2({ S74 }),
  .ZN({ S24812 })
);
NAND3_X1 #() 
NAND3_X1_4752_ (
  .A1({ S24761 }),
  .A2({ S24747 }),
  .A3({ S25957[1043] }),
  .ZN({ S24813 })
);
OAI21_X1 #() 
OAI21_X1_2239_ (
  .A({ S24813 }),
  .B1({ S24811 }),
  .B2({ S24812 }),
  .ZN({ S24814 })
);
AOI211_X1 #() 
AOI211_X1_73_ (
  .A({ S22921 }),
  .B({ S24810 }),
  .C1({ S24776 }),
  .C2({ S24814 }),
  .ZN({ S24815 })
);
NAND4_X1 #() 
NAND4_X1_508_ (
  .A1({ S24746 }),
  .A2({ S24747 }),
  .A3({ S74 }),
  .A4({ S25957[1042] }),
  .ZN({ S24816 })
);
INV_X1 #() 
INV_X1_1417_ (
  .A({ S24816 }),
  .ZN({ S24817 })
);
AOI211_X1 #() 
AOI211_X1_74_ (
  .A({ S25957[1044] }),
  .B({ S24817 }),
  .C1({ S25957[1043] }),
  .C2({ S24791 }),
  .ZN({ S24818 })
);
NOR2_X1 #() 
NOR2_X1_1106_ (
  .A1({ S23195 }),
  .A2({ S25957[1042] }),
  .ZN({ S24819 })
);
AOI21_X1 #() 
AOI21_X1_2363_ (
  .A({ S25957[1043] }),
  .B1({ S24819 }),
  .B2({ S25957[1041] }),
  .ZN({ S24820 })
);
NAND2_X1 #() 
NAND2_X1_4326_ (
  .A1({ S24820 }),
  .A2({ S24745 }),
  .ZN({ S24821 })
);
AOI21_X1 #() 
AOI21_X1_2364_ (
  .A({ S24776 }),
  .B1({ S24772 }),
  .B2({ S25957[1043] }),
  .ZN({ S24822 })
);
AOI211_X1 #() 
AOI211_X1_75_ (
  .A({ S25957[1045] }),
  .B({ S24818 }),
  .C1({ S24821 }),
  .C2({ S24822 }),
  .ZN({ S24823 })
);
NOR3_X1 #() 
NOR3_X1_148_ (
  .A1({ S24823 }),
  .A2({ S24815 }),
  .A3({ S25957[1046] }),
  .ZN({ S24824 })
);
OAI21_X1 #() 
OAI21_X1_2240_ (
  .A({ S20242 }),
  .B1({ S24824 }),
  .B2({ S24807 }),
  .ZN({ S24825 })
);
NAND2_X1 #() 
NAND2_X1_4327_ (
  .A1({ S24825 }),
  .A2({ S24785 }),
  .ZN({ S24826 })
);
NAND2_X1 #() 
NAND2_X1_4328_ (
  .A1({ S24826 }),
  .A2({ S22145 }),
  .ZN({ S24827 })
);
INV_X1 #() 
INV_X1_1418_ (
  .A({ S24827 }),
  .ZN({ S24828 })
);
NOR2_X1 #() 
NOR2_X1_1107_ (
  .A1({ S24826 }),
  .A2({ S22145 }),
  .ZN({ S24829 })
);
OAI21_X1 #() 
OAI21_X1_2241_ (
  .A({ S25957[1087] }),
  .B1({ S24828 }),
  .B2({ S24829 }),
  .ZN({ S24830 })
);
INV_X1 #() 
INV_X1_1419_ (
  .A({ S25957[1087] }),
  .ZN({ S24831 })
);
NOR2_X1 #() 
NOR2_X1_1108_ (
  .A1({ S24828 }),
  .A2({ S24829 }),
  .ZN({ S25957[991] })
);
NAND2_X1 #() 
NAND2_X1_4329_ (
  .A1({ S25957[991] }),
  .A2({ S24831 }),
  .ZN({ S24832 })
);
NAND3_X1 #() 
NAND3_X1_4753_ (
  .A1({ S24832 }),
  .A2({ S22150 }),
  .A3({ S24830 }),
  .ZN({ S24833 })
);
NAND2_X1 #() 
NAND2_X1_4330_ (
  .A1({ S24832 }),
  .A2({ S24830 }),
  .ZN({ S25957[959] })
);
NAND2_X1 #() 
NAND2_X1_4331_ (
  .A1({ S25957[959] }),
  .A2({ S25957[1055] }),
  .ZN({ S24834 })
);
NAND2_X1 #() 
NAND2_X1_4332_ (
  .A1({ S24834 }),
  .A2({ S24833 }),
  .ZN({ S24835 })
);
INV_X1 #() 
INV_X1_1420_ (
  .A({ S24835 }),
  .ZN({ S25957[927] })
);
XOR2_X1 #() 
XOR2_X1_76_ (
  .A({ S25957[1118] }),
  .B({ S25957[1214] }),
  .Z({ S25957[1086] })
);
NAND2_X1 #() 
NAND2_X1_4333_ (
  .A1({ S24751 }),
  .A2({ S24746 }),
  .ZN({ S24836 })
);
NAND4_X1 #() 
NAND4_X1_509_ (
  .A1({ S23261 }),
  .A2({ S23195 }),
  .A3({ S24727 }),
  .A4({ S23262 }),
  .ZN({ S24837 })
);
NAND2_X1 #() 
NAND2_X1_4334_ (
  .A1({ S24837 }),
  .A2({ S24797 }),
  .ZN({ S24838 })
);
OAI221_X1 #() 
OAI221_X1_125_ (
  .A({ S24776 }),
  .B1({ S24838 }),
  .B2({ S74 }),
  .C1({ S24836 }),
  .C2({ S24764 }),
  .ZN({ S24839 })
);
NAND3_X1 #() 
NAND3_X1_4754_ (
  .A1({ S25957[1042] }),
  .A2({ S20546 }),
  .A3({ S20549 }),
  .ZN({ S24840 })
);
OAI22_X1 #() 
OAI22_X1_111_ (
  .A1({ S24837 }),
  .A2({ S25957[1043] }),
  .B1({ S23263 }),
  .B2({ S24840 }),
  .ZN({ S24841 })
);
OAI21_X1 #() 
OAI21_X1_2242_ (
  .A({ S25957[1044] }),
  .B1({ S24817 }),
  .B2({ S24841 }),
  .ZN({ S24842 })
);
AOI21_X1 #() 
AOI21_X1_2365_ (
  .A({ S22921 }),
  .B1({ S24839 }),
  .B2({ S24842 }),
  .ZN({ S24843 })
);
AOI22_X1 #() 
AOI22_X1_495_ (
  .A1({ S23195 }),
  .A2({ S25957[1042] }),
  .B1({ S20549 }),
  .B2({ S20546 }),
  .ZN({ S24844 })
);
AOI21_X1 #() 
AOI21_X1_2366_ (
  .A({ S74 }),
  .B1({ S24772 }),
  .B2({ S24762 }),
  .ZN({ S24845 })
);
AOI21_X1 #() 
AOI21_X1_2367_ (
  .A({ S24845 }),
  .B1({ S24844 }),
  .B2({ S24748 }),
  .ZN({ S24846 })
);
NAND2_X1 #() 
NAND2_X1_4335_ (
  .A1({ S24747 }),
  .A2({ S24727 }),
  .ZN({ S24847 })
);
OAI21_X1 #() 
OAI21_X1_2243_ (
  .A({ S24739 }),
  .B1({ S25957[1043] }),
  .B2({ S24847 }),
  .ZN({ S24848 })
);
OAI21_X1 #() 
OAI21_X1_2244_ (
  .A({ S24848 }),
  .B1({ S24846 }),
  .B2({ S25957[1044] }),
  .ZN({ S24849 })
);
AOI21_X1 #() 
AOI21_X1_2368_ (
  .A({ S24843 }),
  .B1({ S24849 }),
  .B2({ S22921 }),
  .ZN({ S24850 })
);
NOR2_X1 #() 
NOR2_X1_1109_ (
  .A1({ S24819 }),
  .A2({ S74 }),
  .ZN({ S24851 })
);
AOI21_X1 #() 
AOI21_X1_2369_ (
  .A({ S25957[1043] }),
  .B1({ S24724 }),
  .B2({ S24798 }),
  .ZN({ S24852 })
);
AOI211_X1 #() 
AOI211_X1_76_ (
  .A({ S24776 }),
  .B({ S24852 }),
  .C1({ S24778 }),
  .C2({ S24851 }),
  .ZN({ S24853 })
);
AOI21_X1 #() 
AOI21_X1_2370_ (
  .A({ S25957[1044] }),
  .B1({ S24758 }),
  .B2({ S24736 }),
  .ZN({ S24854 })
);
OAI21_X1 #() 
OAI21_X1_2245_ (
  .A({ S25957[1045] }),
  .B1({ S24853 }),
  .B2({ S24854 }),
  .ZN({ S24855 })
);
AND3_X1 #() 
AND3_X1_172_ (
  .A1({ S24809 }),
  .A2({ S24761 }),
  .A3({ S24797 }),
  .ZN({ S24856 })
);
INV_X1 #() 
INV_X1_1421_ (
  .A({ S24797 }),
  .ZN({ S24857 })
);
NOR2_X1 #() 
NOR2_X1_1110_ (
  .A1({ S74 }),
  .A2({ S25957[1040] }),
  .ZN({ S24858 })
);
NAND2_X1 #() 
NAND2_X1_4336_ (
  .A1({ S24857 }),
  .A2({ S24858 }),
  .ZN({ S24859 })
);
NAND2_X1 #() 
NAND2_X1_4337_ (
  .A1({ S24859 }),
  .A2({ S24776 }),
  .ZN({ S24860 })
);
AOI211_X1 #() 
AOI211_X1_77_ (
  .A({ S24856 }),
  .B({ S24860 }),
  .C1({ S24811 }),
  .C2({ S25957[1043] }),
  .ZN({ S24861 })
);
NAND2_X1 #() 
NAND2_X1_4338_ (
  .A1({ S24748 }),
  .A2({ S24844 }),
  .ZN({ S24862 })
);
NAND3_X1 #() 
NAND3_X1_4755_ (
  .A1({ S24724 }),
  .A2({ S24732 }),
  .A3({ S24762 }),
  .ZN({ S24863 })
);
NAND2_X1 #() 
NAND2_X1_4339_ (
  .A1({ S24863 }),
  .A2({ S25957[1043] }),
  .ZN({ S24864 })
);
AOI21_X1 #() 
AOI21_X1_2371_ (
  .A({ S24776 }),
  .B1({ S24862 }),
  .B2({ S24864 }),
  .ZN({ S24865 })
);
OAI21_X1 #() 
OAI21_X1_2246_ (
  .A({ S22921 }),
  .B1({ S24861 }),
  .B2({ S24865 }),
  .ZN({ S24866 })
);
NAND2_X1 #() 
NAND2_X1_4340_ (
  .A1({ S24866 }),
  .A2({ S24855 }),
  .ZN({ S24867 })
);
NAND2_X1 #() 
NAND2_X1_4341_ (
  .A1({ S24867 }),
  .A2({ S25957[1046] }),
  .ZN({ S24868 })
);
OAI211_X1 #() 
OAI211_X1_1508_ (
  .A({ S24868 }),
  .B({ S25957[1047] }),
  .C1({ S25957[1046] }),
  .C2({ S24850 }),
  .ZN({ S24869 })
);
NAND3_X1 #() 
NAND3_X1_4756_ (
  .A1({ S24777 }),
  .A2({ S74 }),
  .A3({ S23195 }),
  .ZN({ S24870 })
);
INV_X1 #() 
INV_X1_1422_ (
  .A({ S24761 }),
  .ZN({ S24871 })
);
NAND2_X1 #() 
NAND2_X1_4342_ (
  .A1({ S24871 }),
  .A2({ S25957[1043] }),
  .ZN({ S24872 })
);
NAND3_X1 #() 
NAND3_X1_4757_ (
  .A1({ S24872 }),
  .A2({ S25957[1044] }),
  .A3({ S24870 }),
  .ZN({ S24873 })
);
AOI21_X1 #() 
AOI21_X1_2372_ (
  .A({ S24727 }),
  .B1({ S24746 }),
  .B2({ S24747 }),
  .ZN({ S24874 })
);
OAI211_X1 #() 
OAI211_X1_1509_ (
  .A({ S24864 }),
  .B({ S24776 }),
  .C1({ S25957[1043] }),
  .C2({ S24874 }),
  .ZN({ S24875 })
);
AOI21_X1 #() 
AOI21_X1_2373_ (
  .A({ S25957[1045] }),
  .B1({ S24875 }),
  .B2({ S24873 }),
  .ZN({ S24876 })
);
NAND2_X1 #() 
NAND2_X1_4343_ (
  .A1({ S24790 }),
  .A2({ S24751 }),
  .ZN({ S24877 })
);
NAND2_X1 #() 
NAND2_X1_4344_ (
  .A1({ S24746 }),
  .A2({ S24798 }),
  .ZN({ S24878 })
);
AOI21_X1 #() 
AOI21_X1_2374_ (
  .A({ S24776 }),
  .B1({ S24878 }),
  .B2({ S25957[1043] }),
  .ZN({ S24879 })
);
NAND2_X1 #() 
NAND2_X1_4345_ (
  .A1({ S25957[1043] }),
  .A2({ S24735 }),
  .ZN({ S24880 })
);
AOI21_X1 #() 
AOI21_X1_2375_ (
  .A({ S25957[1044] }),
  .B1({ S24880 }),
  .B2({ S24780 }),
  .ZN({ S24881 })
);
AOI211_X1 #() 
AOI211_X1_78_ (
  .A({ S22921 }),
  .B({ S24881 }),
  .C1({ S24877 }),
  .C2({ S24879 }),
  .ZN({ S24882 })
);
OR2_X1 #() 
OR2_X1_61_ (
  .A1({ S24882 }),
  .A2({ S22832 }),
  .ZN({ S24883 })
);
NAND2_X1 #() 
NAND2_X1_4346_ (
  .A1({ S24752 }),
  .A2({ S25957[1044] }),
  .ZN({ S24884 })
);
NAND2_X1 #() 
NAND2_X1_4347_ (
  .A1({ S24723 }),
  .A2({ S24727 }),
  .ZN({ S24885 })
);
AOI21_X1 #() 
AOI21_X1_2376_ (
  .A({ S74 }),
  .B1({ S24745 }),
  .B2({ S24885 }),
  .ZN({ S24886 })
);
NAND2_X1 #() 
NAND2_X1_4348_ (
  .A1({ S24797 }),
  .A2({ S25957[1043] }),
  .ZN({ S24887 })
);
NAND2_X1 #() 
NAND2_X1_4349_ (
  .A1({ S24769 }),
  .A2({ S74 }),
  .ZN({ S24888 })
);
OAI22_X1 #() 
OAI22_X1_112_ (
  .A1({ S24888 }),
  .A2({ S24750 }),
  .B1({ S24887 }),
  .B2({ S24871 }),
  .ZN({ S24889 })
);
OAI22_X1 #() 
OAI22_X1_113_ (
  .A1({ S24889 }),
  .A2({ S25957[1044] }),
  .B1({ S24884 }),
  .B2({ S24886 }),
  .ZN({ S24890 })
);
NAND2_X1 #() 
NAND2_X1_4350_ (
  .A1({ S24890 }),
  .A2({ S25957[1045] }),
  .ZN({ S24891 })
);
NAND2_X1 #() 
NAND2_X1_4351_ (
  .A1({ S24730 }),
  .A2({ S24809 }),
  .ZN({ S24892 })
);
AOI21_X1 #() 
AOI21_X1_2377_ (
  .A({ S24776 }),
  .B1({ S24789 }),
  .B2({ S24892 }),
  .ZN({ S24893 })
);
NOR2_X1 #() 
NOR2_X1_1111_ (
  .A1({ S25957[1044] }),
  .A2({ S74 }),
  .ZN({ S24894 })
);
NAND3_X1 #() 
NAND3_X1_4758_ (
  .A1({ S24772 }),
  .A2({ S24777 }),
  .A3({ S24762 }),
  .ZN({ S24895 })
);
NAND2_X1 #() 
NAND2_X1_4352_ (
  .A1({ S24895 }),
  .A2({ S24894 }),
  .ZN({ S24896 })
);
NAND2_X1 #() 
NAND2_X1_4353_ (
  .A1({ S24896 }),
  .A2({ S22921 }),
  .ZN({ S24897 })
);
OAI211_X1 #() 
OAI211_X1_1510_ (
  .A({ S24891 }),
  .B({ S22832 }),
  .C1({ S24893 }),
  .C2({ S24897 }),
  .ZN({ S24898 })
);
OAI211_X1 #() 
OAI211_X1_1511_ (
  .A({ S20242 }),
  .B({ S24898 }),
  .C1({ S24883 }),
  .C2({ S24876 }),
  .ZN({ S24899 })
);
AOI21_X1 #() 
AOI21_X1_2378_ (
  .A({ S22151 }),
  .B1({ S24869 }),
  .B2({ S24899 }),
  .ZN({ S24900 })
);
NAND2_X1 #() 
NAND2_X1_4354_ (
  .A1({ S24869 }),
  .A2({ S24899 }),
  .ZN({ S24901 })
);
NOR2_X1 #() 
NOR2_X1_1112_ (
  .A1({ S24901 }),
  .A2({ S25957[1246] }),
  .ZN({ S24902 })
);
NOR2_X1 #() 
NOR2_X1_1113_ (
  .A1({ S24902 }),
  .A2({ S24900 }),
  .ZN({ S25957[990] })
);
XNOR2_X1 #() 
XNOR2_X1_177_ (
  .A({ S25957[990] }),
  .B({ S21433 }),
  .ZN({ S25957[926] })
);
NAND2_X1 #() 
NAND2_X1_4355_ (
  .A1({ S22287 }),
  .A2({ S22289 }),
  .ZN({ S24903 })
);
XNOR2_X1 #() 
XNOR2_X1_178_ (
  .A({ S24903 }),
  .B({ S25957[1213] }),
  .ZN({ S25957[1085] })
);
NAND2_X1 #() 
NAND2_X1_4356_ (
  .A1({ S24777 }),
  .A2({ S24762 }),
  .ZN({ S24904 })
);
NAND2_X1 #() 
NAND2_X1_4357_ (
  .A1({ S24797 }),
  .A2({ S24798 }),
  .ZN({ S24905 })
);
NAND2_X1 #() 
NAND2_X1_4358_ (
  .A1({ S24905 }),
  .A2({ S74 }),
  .ZN({ S24906 })
);
OAI21_X1 #() 
OAI21_X1_2247_ (
  .A({ S24906 }),
  .B1({ S74 }),
  .B2({ S24904 }),
  .ZN({ S24907 })
);
NAND2_X1 #() 
NAND2_X1_4359_ (
  .A1({ S24864 }),
  .A2({ S24816 }),
  .ZN({ S24908 })
);
MUX2_X1 #() 
MUX2_X1_16_ (
  .A({ S24908 }),
  .B({ S24907 }),
  .S({ S25957[1044] }),
  .Z({ S24909 })
);
NAND2_X1 #() 
NAND2_X1_4360_ (
  .A1({ S24847 }),
  .A2({ S24772 }),
  .ZN({ S24910 })
);
AOI21_X1 #() 
AOI21_X1_2379_ (
  .A({ S24776 }),
  .B1({ S24858 }),
  .B2({ S24777 }),
  .ZN({ S24911 })
);
OAI21_X1 #() 
OAI21_X1_2248_ (
  .A({ S24911 }),
  .B1({ S24910 }),
  .B2({ S25957[1043] }),
  .ZN({ S24912 })
);
OAI21_X1 #() 
OAI21_X1_2249_ (
  .A({ S24894 }),
  .B1({ S24811 }),
  .B2({ S24905 }),
  .ZN({ S24913 })
);
NAND2_X1 #() 
NAND2_X1_4361_ (
  .A1({ S23263 }),
  .A2({ S24798 }),
  .ZN({ S24914 })
);
NAND3_X1 #() 
NAND3_X1_4759_ (
  .A1({ S24914 }),
  .A2({ S24776 }),
  .A3({ S74 }),
  .ZN({ S24915 })
);
NAND4_X1 #() 
NAND4_X1_510_ (
  .A1({ S24912 }),
  .A2({ S25957[1045] }),
  .A3({ S24913 }),
  .A4({ S24915 }),
  .ZN({ S24916 })
);
OAI211_X1 #() 
OAI211_X1_1512_ (
  .A({ S25957[1046] }),
  .B({ S24916 }),
  .C1({ S24909 }),
  .C2({ S25957[1045] }),
  .ZN({ S24917 })
);
NAND3_X1 #() 
NAND3_X1_4760_ (
  .A1({ S24811 }),
  .A2({ S25957[1043] }),
  .A3({ S94 }),
  .ZN({ S24918 })
);
AOI21_X1 #() 
AOI21_X1_2380_ (
  .A({ S24776 }),
  .B1({ S24751 }),
  .B2({ S23263 }),
  .ZN({ S24919 })
);
NAND2_X1 #() 
NAND2_X1_4362_ (
  .A1({ S24918 }),
  .A2({ S24919 }),
  .ZN({ S24920 })
);
NAND2_X1 #() 
NAND2_X1_4363_ (
  .A1({ S24796 }),
  .A2({ S23263 }),
  .ZN({ S24921 })
);
NAND2_X1 #() 
NAND2_X1_4364_ (
  .A1({ S24745 }),
  .A2({ S24921 }),
  .ZN({ S24922 })
);
AOI21_X1 #() 
AOI21_X1_2381_ (
  .A({ S24820 }),
  .B1({ S24922 }),
  .B2({ S25957[1043] }),
  .ZN({ S24923 })
);
OAI21_X1 #() 
OAI21_X1_2250_ (
  .A({ S24920 }),
  .B1({ S24923 }),
  .B2({ S25957[1044] }),
  .ZN({ S24924 })
);
OAI21_X1 #() 
OAI21_X1_2251_ (
  .A({ S74 }),
  .B1({ S24764 }),
  .B2({ S24767 }),
  .ZN({ S24925 })
);
OAI21_X1 #() 
OAI21_X1_2252_ (
  .A({ S24925 }),
  .B1({ S74 }),
  .B2({ S24803 }),
  .ZN({ S24926 })
);
NAND2_X1 #() 
NAND2_X1_4365_ (
  .A1({ S25957[1043] }),
  .A2({ S23263 }),
  .ZN({ S24927 })
);
NAND3_X1 #() 
NAND3_X1_4761_ (
  .A1({ S24746 }),
  .A2({ S24777 }),
  .A3({ S74 }),
  .ZN({ S24928 })
);
AOI21_X1 #() 
AOI21_X1_2382_ (
  .A({ S25957[1044] }),
  .B1({ S24928 }),
  .B2({ S24927 }),
  .ZN({ S24929 })
);
AOI21_X1 #() 
AOI21_X1_2383_ (
  .A({ S24929 }),
  .B1({ S24926 }),
  .B2({ S25957[1044] }),
  .ZN({ S24930 })
);
AOI21_X1 #() 
AOI21_X1_2384_ (
  .A({ S25957[1046] }),
  .B1({ S24930 }),
  .B2({ S25957[1045] }),
  .ZN({ S24931 })
);
OAI21_X1 #() 
OAI21_X1_2253_ (
  .A({ S24931 }),
  .B1({ S25957[1045] }),
  .B2({ S24924 }),
  .ZN({ S24932 })
);
NAND3_X1 #() 
NAND3_X1_4762_ (
  .A1({ S24932 }),
  .A2({ S25957[1047] }),
  .A3({ S24917 }),
  .ZN({ S24933 })
);
NOR2_X1 #() 
NOR2_X1_1114_ (
  .A1({ S23263 }),
  .A2({ S24741 }),
  .ZN({ S24934 })
);
NOR3_X1 #() 
NOR3_X1_149_ (
  .A1({ S24799 }),
  .A2({ S24934 }),
  .A3({ S74 }),
  .ZN({ S24935 })
);
OAI21_X1 #() 
OAI21_X1_2254_ (
  .A({ S24836 }),
  .B1({ S74 }),
  .B2({ S25957[1040] }),
  .ZN({ S24936 })
);
NAND2_X1 #() 
NAND2_X1_4366_ (
  .A1({ S24936 }),
  .A2({ S24776 }),
  .ZN({ S24937 })
);
NAND3_X1 #() 
NAND3_X1_4763_ (
  .A1({ S24847 }),
  .A2({ S74 }),
  .A3({ S24797 }),
  .ZN({ S24938 })
);
NAND2_X1 #() 
NAND2_X1_4367_ (
  .A1({ S24938 }),
  .A2({ S25957[1044] }),
  .ZN({ S24939 })
);
OAI211_X1 #() 
OAI211_X1_1513_ (
  .A({ S24937 }),
  .B({ S25957[1045] }),
  .C1({ S24935 }),
  .C2({ S24939 }),
  .ZN({ S24940 })
);
NAND3_X1 #() 
NAND3_X1_4764_ (
  .A1({ S24747 }),
  .A2({ S25957[1043] }),
  .A3({ S24727 }),
  .ZN({ S24941 })
);
NAND4_X1 #() 
NAND4_X1_511_ (
  .A1({ S23261 }),
  .A2({ S25957[1040] }),
  .A3({ S25957[1042] }),
  .A4({ S23262 }),
  .ZN({ S24942 })
);
NAND3_X1 #() 
NAND3_X1_4765_ (
  .A1({ S24942 }),
  .A2({ S24777 }),
  .A3({ S24741 }),
  .ZN({ S24943 })
);
OAI211_X1 #() 
OAI211_X1_1514_ (
  .A({ S25957[1044] }),
  .B({ S24941 }),
  .C1({ S24943 }),
  .C2({ S25957[1043] }),
  .ZN({ S24944 })
);
NOR2_X1 #() 
NOR2_X1_1115_ (
  .A1({ S24723 }),
  .A2({ S74 }),
  .ZN({ S24945 })
);
NAND2_X1 #() 
NAND2_X1_4368_ (
  .A1({ S24837 }),
  .A2({ S74 }),
  .ZN({ S24946 })
);
NAND4_X1 #() 
NAND4_X1_512_ (
  .A1({ S24797 }),
  .A2({ S25957[1043] }),
  .A3({ S24732 }),
  .A4({ S24762 }),
  .ZN({ S24947 })
);
NAND2_X1 #() 
NAND2_X1_4369_ (
  .A1({ S24947 }),
  .A2({ S24946 }),
  .ZN({ S24948 })
);
OAI211_X1 #() 
OAI211_X1_1515_ (
  .A({ S24948 }),
  .B({ S24776 }),
  .C1({ S24798 }),
  .C2({ S24945 }),
  .ZN({ S24949 })
);
NAND3_X1 #() 
NAND3_X1_4766_ (
  .A1({ S24949 }),
  .A2({ S22921 }),
  .A3({ S24944 }),
  .ZN({ S24950 })
);
NAND3_X1 #() 
NAND3_X1_4767_ (
  .A1({ S24950 }),
  .A2({ S24940 }),
  .A3({ S25957[1046] }),
  .ZN({ S24951 })
);
OAI21_X1 #() 
OAI21_X1_2255_ (
  .A({ S24946 }),
  .B1({ S74 }),
  .B2({ S24885 }),
  .ZN({ S24952 })
);
NAND2_X1 #() 
NAND2_X1_4370_ (
  .A1({ S24952 }),
  .A2({ S25957[1044] }),
  .ZN({ S24953 })
);
NAND2_X1 #() 
NAND2_X1_4371_ (
  .A1({ S24880 }),
  .A2({ S24733 }),
  .ZN({ S24954 })
);
NAND2_X1 #() 
NAND2_X1_4372_ (
  .A1({ S24881 }),
  .A2({ S24954 }),
  .ZN({ S24955 })
);
AOI21_X1 #() 
AOI21_X1_2385_ (
  .A({ S22921 }),
  .B1({ S24953 }),
  .B2({ S24955 }),
  .ZN({ S24956 })
);
AOI21_X1 #() 
AOI21_X1_2386_ (
  .A({ S25957[1044] }),
  .B1({ S24724 }),
  .B2({ S74 }),
  .ZN({ S24957 })
);
OAI211_X1 #() 
OAI211_X1_1516_ (
  .A({ S24957 }),
  .B({ S25957[1040] }),
  .C1({ S23263 }),
  .C2({ S74 }),
  .ZN({ S24958 })
);
NAND3_X1 #() 
NAND3_X1_4768_ (
  .A1({ S24745 }),
  .A2({ S74 }),
  .A3({ S24885 }),
  .ZN({ S24959 })
);
NAND3_X1 #() 
NAND3_X1_4769_ (
  .A1({ S24746 }),
  .A2({ S24747 }),
  .A3({ S25957[1042] }),
  .ZN({ S24960 })
);
NAND3_X1 #() 
NAND3_X1_4770_ (
  .A1({ S24960 }),
  .A2({ S25957[1043] }),
  .A3({ S24769 }),
  .ZN({ S24961 })
);
NAND3_X1 #() 
NAND3_X1_4771_ (
  .A1({ S24959 }),
  .A2({ S24961 }),
  .A3({ S25957[1044] }),
  .ZN({ S24962 })
);
AOI21_X1 #() 
AOI21_X1_2387_ (
  .A({ S25957[1045] }),
  .B1({ S24962 }),
  .B2({ S24958 }),
  .ZN({ S24963 })
);
OAI21_X1 #() 
OAI21_X1_2256_ (
  .A({ S22832 }),
  .B1({ S24963 }),
  .B2({ S24956 }),
  .ZN({ S24964 })
);
NAND3_X1 #() 
NAND3_X1_4772_ (
  .A1({ S24964 }),
  .A2({ S24951 }),
  .A3({ S20242 }),
  .ZN({ S24965 })
);
NAND3_X1 #() 
NAND3_X1_4773_ (
  .A1({ S24933 }),
  .A2({ S22288 }),
  .A3({ S24965 }),
  .ZN({ S24966 })
);
INV_X1 #() 
INV_X1_1423_ (
  .A({ S24966 }),
  .ZN({ S24967 })
);
AOI21_X1 #() 
AOI21_X1_2388_ (
  .A({ S22288 }),
  .B1({ S24933 }),
  .B2({ S24965 }),
  .ZN({ S24968 })
);
OAI21_X1 #() 
OAI21_X1_2257_ (
  .A({ S25957[1085] }),
  .B1({ S24967 }),
  .B2({ S24968 }),
  .ZN({ S24969 })
);
INV_X1 #() 
INV_X1_1424_ (
  .A({ S25957[1085] }),
  .ZN({ S24970 })
);
NOR2_X1 #() 
NOR2_X1_1116_ (
  .A1({ S24967 }),
  .A2({ S24968 }),
  .ZN({ S25957[989] })
);
NAND2_X1 #() 
NAND2_X1_4373_ (
  .A1({ S25957[989] }),
  .A2({ S24970 }),
  .ZN({ S24971 })
);
NAND3_X1 #() 
NAND3_X1_4774_ (
  .A1({ S24971 }),
  .A2({ S25957[1053] }),
  .A3({ S24969 }),
  .ZN({ S24972 })
);
OAI21_X1 #() 
OAI21_X1_2258_ (
  .A({ S24970 }),
  .B1({ S24967 }),
  .B2({ S24968 }),
  .ZN({ S24973 })
);
INV_X1 #() 
INV_X1_1425_ (
  .A({ S24968 }),
  .ZN({ S24974 })
);
NAND3_X1 #() 
NAND3_X1_4775_ (
  .A1({ S24974 }),
  .A2({ S25957[1085] }),
  .A3({ S24966 }),
  .ZN({ S24975 })
);
NAND3_X1 #() 
NAND3_X1_4776_ (
  .A1({ S24973 }),
  .A2({ S24975 }),
  .A3({ S22294 }),
  .ZN({ S24976 })
);
NAND2_X1 #() 
NAND2_X1_4374_ (
  .A1({ S24972 }),
  .A2({ S24976 }),
  .ZN({ S25957[925] })
);
INV_X1 #() 
INV_X1_1426_ (
  .A({ S25957[1212] }),
  .ZN({ S24977 })
);
NAND2_X1 #() 
NAND2_X1_4375_ (
  .A1({ S22352 }),
  .A2({ S22356 }),
  .ZN({ S24978 })
);
INV_X1 #() 
INV_X1_1427_ (
  .A({ S24978 }),
  .ZN({ S25957[1116] })
);
NAND2_X1 #() 
NAND2_X1_4376_ (
  .A1({ S25957[1116] }),
  .A2({ S24977 }),
  .ZN({ S24979 })
);
NAND2_X1 #() 
NAND2_X1_4377_ (
  .A1({ S24978 }),
  .A2({ S25957[1212] }),
  .ZN({ S24980 })
);
NAND2_X1 #() 
NAND2_X1_4378_ (
  .A1({ S24979 }),
  .A2({ S24980 }),
  .ZN({ S25957[1084] })
);
NAND2_X1 #() 
NAND2_X1_4379_ (
  .A1({ S24748 }),
  .A2({ S24790 }),
  .ZN({ S24981 })
);
NAND2_X1 #() 
NAND2_X1_4380_ (
  .A1({ S24981 }),
  .A2({ S74 }),
  .ZN({ S24982 })
);
NAND3_X1 #() 
NAND3_X1_4777_ (
  .A1({ S25957[1043] }),
  .A2({ S25957[1041] }),
  .A3({ S23195 }),
  .ZN({ S24983 })
);
AND3_X1 #() 
AND3_X1_173_ (
  .A1({ S24941 }),
  .A2({ S24983 }),
  .A3({ S24776 }),
  .ZN({ S24984 })
);
NAND2_X1 #() 
NAND2_X1_4381_ (
  .A1({ S24982 }),
  .A2({ S24984 }),
  .ZN({ S24985 })
);
NAND2_X1 #() 
NAND2_X1_4382_ (
  .A1({ S24724 }),
  .A2({ S24732 }),
  .ZN({ S24986 })
);
OAI21_X1 #() 
OAI21_X1_2259_ (
  .A({ S74 }),
  .B1({ S24904 }),
  .B2({ S24986 }),
  .ZN({ S24987 })
);
NOR2_X1 #() 
NOR2_X1_1117_ (
  .A1({ S24945 }),
  .A2({ S24776 }),
  .ZN({ S24988 })
);
NAND3_X1 #() 
NAND3_X1_4778_ (
  .A1({ S24987 }),
  .A2({ S24813 }),
  .A3({ S24988 }),
  .ZN({ S24989 })
);
NAND3_X1 #() 
NAND3_X1_4779_ (
  .A1({ S24985 }),
  .A2({ S25957[1045] }),
  .A3({ S24989 }),
  .ZN({ S24990 })
);
NAND3_X1 #() 
NAND3_X1_4780_ (
  .A1({ S25957[1043] }),
  .A2({ S23263 }),
  .A3({ S24798 }),
  .ZN({ S24991 })
);
NAND2_X1 #() 
NAND2_X1_4383_ (
  .A1({ S25957[1043] }),
  .A2({ S24776 }),
  .ZN({ S24992 })
);
NAND4_X1 #() 
NAND4_X1_513_ (
  .A1({ S24772 }),
  .A2({ S24762 }),
  .A3({ S24777 }),
  .A4({ S24776 }),
  .ZN({ S24993 })
);
NAND2_X1 #() 
NAND2_X1_4384_ (
  .A1({ S24993 }),
  .A2({ S24992 }),
  .ZN({ S24994 })
);
NAND2_X1 #() 
NAND2_X1_4385_ (
  .A1({ S24994 }),
  .A2({ S24991 }),
  .ZN({ S24995 })
);
OAI21_X1 #() 
OAI21_X1_2260_ (
  .A({ S74 }),
  .B1({ S24811 }),
  .B2({ S24905 }),
  .ZN({ S24996 })
);
NAND2_X1 #() 
NAND2_X1_4386_ (
  .A1({ S24777 }),
  .A2({ S24732 }),
  .ZN({ S24997 })
);
AOI21_X1 #() 
AOI21_X1_2389_ (
  .A({ S24776 }),
  .B1({ S24757 }),
  .B2({ S24997 }),
  .ZN({ S24998 })
);
AOI21_X1 #() 
AOI21_X1_2390_ (
  .A({ S25957[1045] }),
  .B1({ S24996 }),
  .B2({ S24998 }),
  .ZN({ S24999 })
);
NAND2_X1 #() 
NAND2_X1_4387_ (
  .A1({ S24999 }),
  .A2({ S24995 }),
  .ZN({ S25000 })
);
NAND3_X1 #() 
NAND3_X1_4781_ (
  .A1({ S24990 }),
  .A2({ S22832 }),
  .A3({ S25000 }),
  .ZN({ S25001 })
);
NAND2_X1 #() 
NAND2_X1_4388_ (
  .A1({ S24760 }),
  .A2({ S74 }),
  .ZN({ S25002 })
);
NAND3_X1 #() 
NAND3_X1_4782_ (
  .A1({ S25002 }),
  .A2({ S24941 }),
  .A3({ S25957[1044] }),
  .ZN({ S25003 })
);
NAND2_X1 #() 
NAND2_X1_4389_ (
  .A1({ S24777 }),
  .A2({ S25957[1043] }),
  .ZN({ S25004 })
);
NAND3_X1 #() 
NAND3_X1_4783_ (
  .A1({ S24761 }),
  .A2({ S74 }),
  .A3({ S23195 }),
  .ZN({ S25005 })
);
OAI211_X1 #() 
OAI211_X1_1517_ (
  .A({ S25005 }),
  .B({ S24776 }),
  .C1({ S25004 }),
  .C2({ S24735 }),
  .ZN({ S25006 })
);
NAND3_X1 #() 
NAND3_X1_4784_ (
  .A1({ S25006 }),
  .A2({ S25003 }),
  .A3({ S25957[1045] }),
  .ZN({ S25007 })
);
OAI211_X1 #() 
OAI211_X1_1518_ (
  .A({ S24813 }),
  .B({ S24776 }),
  .C1({ S25957[1043] }),
  .C2({ S24997 }),
  .ZN({ S25008 })
);
OAI211_X1 #() 
OAI211_X1_1519_ (
  .A({ S24928 }),
  .B({ S25957[1044] }),
  .C1({ S24819 }),
  .C2({ S24927 }),
  .ZN({ S25009 })
);
NAND3_X1 #() 
NAND3_X1_4785_ (
  .A1({ S25009 }),
  .A2({ S25008 }),
  .A3({ S22921 }),
  .ZN({ S25010 })
);
NAND3_X1 #() 
NAND3_X1_4786_ (
  .A1({ S25010 }),
  .A2({ S25007 }),
  .A3({ S25957[1046] }),
  .ZN({ S25011 })
);
NAND3_X1 #() 
NAND3_X1_4787_ (
  .A1({ S25001 }),
  .A2({ S25957[1047] }),
  .A3({ S25011 }),
  .ZN({ S25012 })
);
NAND2_X1 #() 
NAND2_X1_4390_ (
  .A1({ S24808 }),
  .A2({ S94 }),
  .ZN({ S25013 })
);
NAND4_X1 #() 
NAND4_X1_514_ (
  .A1({ S24760 }),
  .A2({ S74 }),
  .A3({ S24761 }),
  .A4({ S24762 }),
  .ZN({ S25014 })
);
AOI21_X1 #() 
AOI21_X1_2391_ (
  .A({ S25957[1045] }),
  .B1({ S25014 }),
  .B2({ S25013 }),
  .ZN({ S25015 })
);
NAND3_X1 #() 
NAND3_X1_4788_ (
  .A1({ S25957[1041] }),
  .A2({ S74 }),
  .A3({ S25957[1040] }),
  .ZN({ S25016 })
);
AOI21_X1 #() 
AOI21_X1_2392_ (
  .A({ S22921 }),
  .B1({ S24918 }),
  .B2({ S25016 }),
  .ZN({ S25017 })
);
OAI21_X1 #() 
OAI21_X1_2261_ (
  .A({ S24776 }),
  .B1({ S25017 }),
  .B2({ S25015 }),
  .ZN({ S25018 })
);
NAND4_X1 #() 
NAND4_X1_515_ (
  .A1({ S24761 }),
  .A2({ S25957[1043] }),
  .A3({ S24741 }),
  .A4({ S24798 }),
  .ZN({ S25019 })
);
AND2_X1 #() 
AND2_X1_269_ (
  .A1({ S24928 }),
  .A2({ S22921 }),
  .ZN({ S25020 })
);
AOI21_X1 #() 
AOI21_X1_2393_ (
  .A({ S22921 }),
  .B1({ S24757 }),
  .B2({ S24847 }),
  .ZN({ S25021 })
);
AOI22_X1 #() 
AOI22_X1_496_ (
  .A1({ S25021 }),
  .A2({ S24906 }),
  .B1({ S25020 }),
  .B2({ S25019 }),
  .ZN({ S25022 })
);
OAI211_X1 #() 
OAI211_X1_1520_ (
  .A({ S25018 }),
  .B({ S22832 }),
  .C1({ S25022 }),
  .C2({ S24776 }),
  .ZN({ S25023 })
);
AOI21_X1 #() 
AOI21_X1_2394_ (
  .A({ S25957[1042] }),
  .B1({ S24746 }),
  .B2({ S24747 }),
  .ZN({ S25024 })
);
OAI21_X1 #() 
OAI21_X1_2262_ (
  .A({ S74 }),
  .B1({ S25024 }),
  .B2({ S24905 }),
  .ZN({ S25025 })
);
AOI21_X1 #() 
AOI21_X1_2395_ (
  .A({ S25957[1044] }),
  .B1({ S24851 }),
  .B2({ S24790 }),
  .ZN({ S25026 })
);
INV_X1 #() 
INV_X1_1428_ (
  .A({ S127 }),
  .ZN({ S25027 })
);
OAI21_X1 #() 
OAI21_X1_2263_ (
  .A({ S25957[1044] }),
  .B1({ S25027 }),
  .B2({ S25957[1042] }),
  .ZN({ S25028 })
);
NAND2_X1 #() 
NAND2_X1_4391_ (
  .A1({ S25028 }),
  .A2({ S25957[1045] }),
  .ZN({ S25029 })
);
AOI21_X1 #() 
AOI21_X1_2396_ (
  .A({ S25029 }),
  .B1({ S25025 }),
  .B2({ S25026 }),
  .ZN({ S25030 })
);
INV_X1 #() 
INV_X1_1429_ (
  .A({ S25030 }),
  .ZN({ S25031 })
);
NAND3_X1 #() 
NAND3_X1_4789_ (
  .A1({ S24724 }),
  .A2({ S74 }),
  .A3({ S24798 }),
  .ZN({ S25032 })
);
OAI211_X1 #() 
OAI211_X1_1521_ (
  .A({ S25957[1044] }),
  .B({ S24737 }),
  .C1({ S25032 }),
  .C2({ S24730 }),
  .ZN({ S25033 })
);
AND2_X1 #() 
AND2_X1_270_ (
  .A1({ S24776 }),
  .A2({ S24840 }),
  .ZN({ S25034 })
);
NAND2_X1 #() 
NAND2_X1_4392_ (
  .A1({ S24819 }),
  .A2({ S25957[1041] }),
  .ZN({ S25035 })
);
NAND2_X1 #() 
NAND2_X1_4393_ (
  .A1({ S25035 }),
  .A2({ S24844 }),
  .ZN({ S25036 })
);
AOI21_X1 #() 
AOI21_X1_2397_ (
  .A({ S25957[1045] }),
  .B1({ S25036 }),
  .B2({ S25034 }),
  .ZN({ S25037 })
);
AOI21_X1 #() 
AOI21_X1_2398_ (
  .A({ S22832 }),
  .B1({ S25037 }),
  .B2({ S25033 }),
  .ZN({ S25038 })
);
AOI21_X1 #() 
AOI21_X1_2399_ (
  .A({ S25957[1047] }),
  .B1({ S25031 }),
  .B2({ S25038 }),
  .ZN({ S25039 })
);
NAND2_X1 #() 
NAND2_X1_4394_ (
  .A1({ S25023 }),
  .A2({ S25039 }),
  .ZN({ S25040 })
);
NAND3_X1 #() 
NAND3_X1_4790_ (
  .A1({ S25012 }),
  .A2({ S25040 }),
  .A3({ S25957[1244] }),
  .ZN({ S25041 })
);
NAND2_X1 #() 
NAND2_X1_4395_ (
  .A1({ S25010 }),
  .A2({ S25007 }),
  .ZN({ S25042 })
);
NAND2_X1 #() 
NAND2_X1_4396_ (
  .A1({ S25042 }),
  .A2({ S25957[1046] }),
  .ZN({ S25043 })
);
AOI21_X1 #() 
AOI21_X1_2400_ (
  .A({ S22921 }),
  .B1({ S24982 }),
  .B2({ S24984 }),
  .ZN({ S25044 })
);
AOI22_X1 #() 
AOI22_X1_497_ (
  .A1({ S25044 }),
  .A2({ S24989 }),
  .B1({ S24999 }),
  .B2({ S24995 }),
  .ZN({ S25045 })
);
OAI211_X1 #() 
OAI211_X1_1522_ (
  .A({ S25957[1047] }),
  .B({ S25043 }),
  .C1({ S25045 }),
  .C2({ S25957[1046] }),
  .ZN({ S25046 })
);
AND2_X1 #() 
AND2_X1_271_ (
  .A1({ S25037 }),
  .A2({ S25033 }),
  .ZN({ S25047 })
);
OAI21_X1 #() 
OAI21_X1_2264_ (
  .A({ S25957[1046] }),
  .B1({ S25047 }),
  .B2({ S25030 }),
  .ZN({ S25048 })
);
OAI211_X1 #() 
OAI211_X1_1523_ (
  .A({ S24789 }),
  .B({ S25957[1044] }),
  .C1({ S25957[1043] }),
  .C2({ S24905 }),
  .ZN({ S25049 })
);
OAI211_X1 #() 
OAI211_X1_1524_ (
  .A({ S25016 }),
  .B({ S24776 }),
  .C1({ S24728 }),
  .C2({ S74 }),
  .ZN({ S25050 })
);
AND3_X1 #() 
AND3_X1_174_ (
  .A1({ S25049 }),
  .A2({ S25050 }),
  .A3({ S25957[1045] }),
  .ZN({ S25051 })
);
NAND2_X1 #() 
NAND2_X1_4397_ (
  .A1({ S25014 }),
  .A2({ S25013 }),
  .ZN({ S25052 })
);
NAND2_X1 #() 
NAND2_X1_4398_ (
  .A1({ S25052 }),
  .A2({ S24776 }),
  .ZN({ S25053 })
);
NAND3_X1 #() 
NAND3_X1_4791_ (
  .A1({ S25019 }),
  .A2({ S24928 }),
  .A3({ S25957[1044] }),
  .ZN({ S25054 })
);
AOI21_X1 #() 
AOI21_X1_2401_ (
  .A({ S25957[1045] }),
  .B1({ S25053 }),
  .B2({ S25054 }),
  .ZN({ S25055 })
);
OAI21_X1 #() 
OAI21_X1_2265_ (
  .A({ S22832 }),
  .B1({ S25055 }),
  .B2({ S25051 }),
  .ZN({ S25056 })
);
NAND3_X1 #() 
NAND3_X1_4792_ (
  .A1({ S25056 }),
  .A2({ S20242 }),
  .A3({ S25048 }),
  .ZN({ S25057 })
);
NAND3_X1 #() 
NAND3_X1_4793_ (
  .A1({ S25046 }),
  .A2({ S25057 }),
  .A3({ S22353 }),
  .ZN({ S25058 })
);
NAND4_X1 #() 
NAND4_X1_516_ (
  .A1({ S25058 }),
  .A2({ S25041 }),
  .A3({ S24980 }),
  .A4({ S24979 }),
  .ZN({ S25059 })
);
AOI21_X1 #() 
AOI21_X1_2402_ (
  .A({ S22353 }),
  .B1({ S25046 }),
  .B2({ S25057 }),
  .ZN({ S25060 })
);
AOI21_X1 #() 
AOI21_X1_2403_ (
  .A({ S25957[1244] }),
  .B1({ S25012 }),
  .B2({ S25040 }),
  .ZN({ S25061 })
);
OAI21_X1 #() 
OAI21_X1_2266_ (
  .A({ S25957[1084] }),
  .B1({ S25060 }),
  .B2({ S25061 }),
  .ZN({ S25062 })
);
NAND3_X1 #() 
NAND3_X1_4794_ (
  .A1({ S25062 }),
  .A2({ S24046 }),
  .A3({ S25059 }),
  .ZN({ S25063 })
);
NAND2_X1 #() 
NAND2_X1_4399_ (
  .A1({ S22354 }),
  .A2({ S22355 }),
  .ZN({ S25957[1148] })
);
NAND3_X1 #() 
NAND3_X1_4795_ (
  .A1({ S25012 }),
  .A2({ S25040 }),
  .A3({ S25957[1148] }),
  .ZN({ S25064 })
);
INV_X1 #() 
INV_X1_1430_ (
  .A({ S25957[1148] }),
  .ZN({ S25065 })
);
NAND3_X1 #() 
NAND3_X1_4796_ (
  .A1({ S25046 }),
  .A2({ S25057 }),
  .A3({ S25065 }),
  .ZN({ S25066 })
);
NAND3_X1 #() 
NAND3_X1_4797_ (
  .A1({ S25066 }),
  .A2({ S25064 }),
  .A3({ S25957[1212] }),
  .ZN({ S25067 })
);
NAND3_X1 #() 
NAND3_X1_4798_ (
  .A1({ S25012 }),
  .A2({ S25040 }),
  .A3({ S25065 }),
  .ZN({ S25068 })
);
NAND3_X1 #() 
NAND3_X1_4799_ (
  .A1({ S25046 }),
  .A2({ S25057 }),
  .A3({ S25957[1148] }),
  .ZN({ S25069 })
);
NAND3_X1 #() 
NAND3_X1_4800_ (
  .A1({ S25069 }),
  .A2({ S25068 }),
  .A3({ S24977 }),
  .ZN({ S25070 })
);
NAND3_X1 #() 
NAND3_X1_4801_ (
  .A1({ S25067 }),
  .A2({ S25070 }),
  .A3({ S25957[1052] }),
  .ZN({ S25071 })
);
NAND2_X1 #() 
NAND2_X1_4400_ (
  .A1({ S25063 }),
  .A2({ S25071 }),
  .ZN({ S25072 })
);
INV_X1 #() 
INV_X1_1431_ (
  .A({ S25072 }),
  .ZN({ S25957[924] })
);
NOR2_X1 #() 
NOR2_X1_1118_ (
  .A1({ S19950 }),
  .A2({ S19954 }),
  .ZN({ S25957[1211] })
);
INV_X1 #() 
INV_X1_1432_ (
  .A({ S25957[1211] }),
  .ZN({ S25073 })
);
NAND2_X1 #() 
NAND2_X1_4401_ (
  .A1({ S22432 }),
  .A2({ S22431 }),
  .ZN({ S25957[1147] })
);
AOI21_X1 #() 
AOI21_X1_2404_ (
  .A({ S24776 }),
  .B1({ S24808 }),
  .B2({ S94 }),
  .ZN({ S25074 })
);
OAI21_X1 #() 
OAI21_X1_2267_ (
  .A({ S25074 }),
  .B1({ S24874 }),
  .B2({ S24888 }),
  .ZN({ S25075 })
);
NAND4_X1 #() 
NAND4_X1_517_ (
  .A1({ S24746 }),
  .A2({ S24747 }),
  .A3({ S74 }),
  .A4({ S24732 }),
  .ZN({ S25076 })
);
OAI21_X1 #() 
OAI21_X1_2268_ (
  .A({ S25076 }),
  .B1({ S25004 }),
  .B2({ S24863 }),
  .ZN({ S25077 })
);
AOI21_X1 #() 
AOI21_X1_2405_ (
  .A({ S22832 }),
  .B1({ S25077 }),
  .B2({ S24776 }),
  .ZN({ S25078 })
);
NAND3_X1 #() 
NAND3_X1_4802_ (
  .A1({ S24745 }),
  .A2({ S74 }),
  .A3({ S24777 }),
  .ZN({ S25079 })
);
AOI21_X1 #() 
AOI21_X1_2406_ (
  .A({ S74 }),
  .B1({ S24767 }),
  .B2({ S23263 }),
  .ZN({ S25080 })
);
NAND2_X1 #() 
NAND2_X1_4402_ (
  .A1({ S25080 }),
  .A2({ S24728 }),
  .ZN({ S25081 })
);
AOI21_X1 #() 
AOI21_X1_2407_ (
  .A({ S24776 }),
  .B1({ S24863 }),
  .B2({ S74 }),
  .ZN({ S25082 })
);
NAND4_X1 #() 
NAND4_X1_518_ (
  .A1({ S25957[1043] }),
  .A2({ S25957[1041] }),
  .A3({ S24732 }),
  .A4({ S24762 }),
  .ZN({ S25083 })
);
AND2_X1 #() 
AND2_X1_272_ (
  .A1({ S25083 }),
  .A2({ S24776 }),
  .ZN({ S25084 })
);
AOI22_X1 #() 
AOI22_X1_498_ (
  .A1({ S25084 }),
  .A2({ S25079 }),
  .B1({ S25082 }),
  .B2({ S25081 }),
  .ZN({ S25085 })
);
AOI22_X1 #() 
AOI22_X1_499_ (
  .A1({ S25085 }),
  .A2({ S22832 }),
  .B1({ S25078 }),
  .B2({ S25075 }),
  .ZN({ S25086 })
);
NAND3_X1 #() 
NAND3_X1_4803_ (
  .A1({ S24761 }),
  .A2({ S74 }),
  .A3({ S24798 }),
  .ZN({ S25087 })
);
OAI211_X1 #() 
OAI211_X1_1525_ (
  .A({ S25957[1044] }),
  .B({ S25087 }),
  .C1({ S24748 }),
  .C2({ S74 }),
  .ZN({ S25088 })
);
NAND4_X1 #() 
NAND4_X1_519_ (
  .A1({ S24746 }),
  .A2({ S24747 }),
  .A3({ S25957[1043] }),
  .A4({ S25957[1042] }),
  .ZN({ S25089 })
);
NAND2_X1 #() 
NAND2_X1_4403_ (
  .A1({ S24751 }),
  .A2({ S94 }),
  .ZN({ S25090 })
);
NAND4_X1 #() 
NAND4_X1_520_ (
  .A1({ S25089 }),
  .A2({ S25090 }),
  .A3({ S24776 }),
  .A4({ S24731 }),
  .ZN({ S25091 })
);
AOI21_X1 #() 
AOI21_X1_2408_ (
  .A({ S25957[1046] }),
  .B1({ S25091 }),
  .B2({ S25088 }),
  .ZN({ S25092 })
);
OAI21_X1 #() 
OAI21_X1_2269_ (
  .A({ S25957[1043] }),
  .B1({ S24796 }),
  .B2({ S23263 }),
  .ZN({ S25093 })
);
OAI21_X1 #() 
OAI21_X1_2270_ (
  .A({ S25093 }),
  .B1({ S24799 }),
  .B2({ S24888 }),
  .ZN({ S25094 })
);
NAND2_X1 #() 
NAND2_X1_4404_ (
  .A1({ S25034 }),
  .A2({ S24878 }),
  .ZN({ S25095 })
);
NAND2_X1 #() 
NAND2_X1_4405_ (
  .A1({ S25095 }),
  .A2({ S25957[1046] }),
  .ZN({ S25096 })
);
AOI21_X1 #() 
AOI21_X1_2409_ (
  .A({ S25096 }),
  .B1({ S25094 }),
  .B2({ S25957[1044] }),
  .ZN({ S25097 })
);
OAI21_X1 #() 
OAI21_X1_2271_ (
  .A({ S22921 }),
  .B1({ S25097 }),
  .B2({ S25092 }),
  .ZN({ S25098 })
);
OAI211_X1 #() 
OAI211_X1_1526_ (
  .A({ S25098 }),
  .B({ S25957[1047] }),
  .C1({ S25086 }),
  .C2({ S22921 }),
  .ZN({ S25099 })
);
OAI21_X1 #() 
OAI21_X1_2272_ (
  .A({ S94 }),
  .B1({ S24723 }),
  .B2({ S25957[1042] }),
  .ZN({ S25100 })
);
OAI211_X1 #() 
OAI211_X1_1527_ (
  .A({ S24938 }),
  .B({ S25957[1044] }),
  .C1({ S74 }),
  .C2({ S25100 }),
  .ZN({ S25101 })
);
AOI21_X1 #() 
AOI21_X1_2410_ (
  .A({ S74 }),
  .B1({ S24885 }),
  .B2({ S24798 }),
  .ZN({ S25102 })
);
INV_X1 #() 
INV_X1_1433_ (
  .A({ S25102 }),
  .ZN({ S25103 })
);
NAND3_X1 #() 
NAND3_X1_4804_ (
  .A1({ S24800 }),
  .A2({ S25103 }),
  .A3({ S24776 }),
  .ZN({ S25104 })
);
NAND3_X1 #() 
NAND3_X1_4805_ (
  .A1({ S25104 }),
  .A2({ S25101 }),
  .A3({ S22921 }),
  .ZN({ S25105 })
);
AOI21_X1 #() 
AOI21_X1_2411_ (
  .A({ S25080 }),
  .B1({ S24960 }),
  .B2({ S74 }),
  .ZN({ S25106 })
);
NAND2_X1 #() 
NAND2_X1_4406_ (
  .A1({ S24761 }),
  .A2({ S25957[1040] }),
  .ZN({ S25107 })
);
OAI21_X1 #() 
OAI21_X1_2273_ (
  .A({ S24776 }),
  .B1({ S24757 }),
  .B2({ S25107 }),
  .ZN({ S25108 })
);
OAI21_X1 #() 
OAI21_X1_2274_ (
  .A({ S25108 }),
  .B1({ S25106 }),
  .B2({ S24776 }),
  .ZN({ S25109 })
);
NAND2_X1 #() 
NAND2_X1_4407_ (
  .A1({ S25109 }),
  .A2({ S25957[1045] }),
  .ZN({ S25110 })
);
NAND3_X1 #() 
NAND3_X1_4806_ (
  .A1({ S25105 }),
  .A2({ S25110 }),
  .A3({ S22832 }),
  .ZN({ S25111 })
);
NAND3_X1 #() 
NAND3_X1_4807_ (
  .A1({ S24821 }),
  .A2({ S25957[1044] }),
  .A3({ S24864 }),
  .ZN({ S25112 })
);
NAND3_X1 #() 
NAND3_X1_4808_ (
  .A1({ S24761 }),
  .A2({ S24747 }),
  .A3({ S74 }),
  .ZN({ S25113 })
);
AOI21_X1 #() 
AOI21_X1_2412_ (
  .A({ S25957[1044] }),
  .B1({ S24858 }),
  .B2({ S24724 }),
  .ZN({ S25114 })
);
AOI21_X1 #() 
AOI21_X1_2413_ (
  .A({ S22921 }),
  .B1({ S25114 }),
  .B2({ S25113 }),
  .ZN({ S25115 })
);
NAND3_X1 #() 
NAND3_X1_4809_ (
  .A1({ S24809 }),
  .A2({ S24761 }),
  .A3({ S24797 }),
  .ZN({ S25116 })
);
NAND3_X1 #() 
NAND3_X1_4810_ (
  .A1({ S24770 }),
  .A2({ S24776 }),
  .A3({ S25116 }),
  .ZN({ S25117 })
);
NAND3_X1 #() 
NAND3_X1_4811_ (
  .A1({ S24723 }),
  .A2({ S74 }),
  .A3({ S24798 }),
  .ZN({ S25118 })
);
AOI21_X1 #() 
AOI21_X1_2414_ (
  .A({ S25957[1045] }),
  .B1({ S25118 }),
  .B2({ S25957[1044] }),
  .ZN({ S25119 })
);
AOI22_X1 #() 
AOI22_X1_500_ (
  .A1({ S25112 }),
  .A2({ S25115 }),
  .B1({ S25117 }),
  .B2({ S25119 }),
  .ZN({ S25120 })
);
AOI21_X1 #() 
AOI21_X1_2415_ (
  .A({ S25957[1047] }),
  .B1({ S25120 }),
  .B2({ S25957[1046] }),
  .ZN({ S25121 })
);
NAND2_X1 #() 
NAND2_X1_4408_ (
  .A1({ S25111 }),
  .A2({ S25121 }),
  .ZN({ S25122 })
);
NAND3_X1 #() 
NAND3_X1_4812_ (
  .A1({ S25099 }),
  .A2({ S25122 }),
  .A3({ S25957[1147] }),
  .ZN({ S25123 })
);
INV_X1 #() 
INV_X1_1434_ (
  .A({ S25957[1147] }),
  .ZN({ S25124 })
);
NAND2_X1 #() 
NAND2_X1_4409_ (
  .A1({ S24770 }),
  .A2({ S25116 }),
  .ZN({ S25125 })
);
NAND2_X1 #() 
NAND2_X1_4410_ (
  .A1({ S25125 }),
  .A2({ S24776 }),
  .ZN({ S25126 })
);
AOI21_X1 #() 
AOI21_X1_2416_ (
  .A({ S25957[1043] }),
  .B1({ S24777 }),
  .B2({ S25957[1040] }),
  .ZN({ S25127 })
);
NAND2_X1 #() 
NAND2_X1_4411_ (
  .A1({ S25127 }),
  .A2({ S25957[1044] }),
  .ZN({ S25128 })
);
NAND3_X1 #() 
NAND3_X1_4813_ (
  .A1({ S25126 }),
  .A2({ S25957[1046] }),
  .A3({ S25128 }),
  .ZN({ S25129 })
);
AOI21_X1 #() 
AOI21_X1_2417_ (
  .A({ S25957[1043] }),
  .B1({ S24960 }),
  .B2({ S24741 }),
  .ZN({ S25130 })
);
OAI21_X1 #() 
OAI21_X1_2275_ (
  .A({ S24776 }),
  .B1({ S25130 }),
  .B2({ S25102 }),
  .ZN({ S25131 })
);
NAND2_X1 #() 
NAND2_X1_4412_ (
  .A1({ S25100 }),
  .A2({ S25957[1043] }),
  .ZN({ S25132 })
);
AND2_X1 #() 
AND2_X1_273_ (
  .A1({ S24724 }),
  .A2({ S74 }),
  .ZN({ S25133 })
);
AOI21_X1 #() 
AOI21_X1_2418_ (
  .A({ S24776 }),
  .B1({ S25133 }),
  .B2({ S24769 }),
  .ZN({ S25134 })
);
AOI21_X1 #() 
AOI21_X1_2419_ (
  .A({ S25957[1046] }),
  .B1({ S25134 }),
  .B2({ S25132 }),
  .ZN({ S25135 })
);
NAND2_X1 #() 
NAND2_X1_4413_ (
  .A1({ S25135 }),
  .A2({ S25131 }),
  .ZN({ S25136 })
);
AOI21_X1 #() 
AOI21_X1_2420_ (
  .A({ S25957[1045] }),
  .B1({ S25136 }),
  .B2({ S25129 }),
  .ZN({ S25137 })
);
AOI22_X1 #() 
AOI22_X1_501_ (
  .A1({ S24820 }),
  .A2({ S24745 }),
  .B1({ S24863 }),
  .B2({ S25957[1043] }),
  .ZN({ S25138 })
);
AOI21_X1 #() 
AOI21_X1_2421_ (
  .A({ S25957[1043] }),
  .B1({ S94 }),
  .B2({ S24724 }),
  .ZN({ S25139 })
);
AOI21_X1 #() 
AOI21_X1_2422_ (
  .A({ S74 }),
  .B1({ S24760 }),
  .B2({ S24741 }),
  .ZN({ S25140 })
);
OAI21_X1 #() 
OAI21_X1_2276_ (
  .A({ S24776 }),
  .B1({ S25140 }),
  .B2({ S25139 }),
  .ZN({ S25141 })
);
OAI211_X1 #() 
OAI211_X1_1528_ (
  .A({ S25141 }),
  .B({ S25957[1046] }),
  .C1({ S25138 }),
  .C2({ S24776 }),
  .ZN({ S25142 })
);
OAI211_X1 #() 
OAI211_X1_1529_ (
  .A({ S22832 }),
  .B({ S25108 }),
  .C1({ S25106 }),
  .C2({ S24776 }),
  .ZN({ S25143 })
);
AOI21_X1 #() 
AOI21_X1_2423_ (
  .A({ S22921 }),
  .B1({ S25142 }),
  .B2({ S25143 }),
  .ZN({ S25144 })
);
OAI21_X1 #() 
OAI21_X1_2277_ (
  .A({ S20242 }),
  .B1({ S25137 }),
  .B2({ S25144 }),
  .ZN({ S25145 })
);
NAND2_X1 #() 
NAND2_X1_4414_ (
  .A1({ S25094 }),
  .A2({ S25957[1044] }),
  .ZN({ S25146 })
);
NAND3_X1 #() 
NAND3_X1_4814_ (
  .A1({ S25146 }),
  .A2({ S22921 }),
  .A3({ S25095 }),
  .ZN({ S25147 })
);
NAND2_X1 #() 
NAND2_X1_4415_ (
  .A1({ S25077 }),
  .A2({ S24776 }),
  .ZN({ S25148 })
);
NAND3_X1 #() 
NAND3_X1_4815_ (
  .A1({ S25148 }),
  .A2({ S25957[1045] }),
  .A3({ S25075 }),
  .ZN({ S25149 })
);
NAND3_X1 #() 
NAND3_X1_4816_ (
  .A1({ S25147 }),
  .A2({ S25957[1046] }),
  .A3({ S25149 }),
  .ZN({ S25150 })
);
NOR2_X1 #() 
NOR2_X1_1119_ (
  .A1({ S24733 }),
  .A2({ S24730 }),
  .ZN({ S25151 })
);
NAND3_X1 #() 
NAND3_X1_4817_ (
  .A1({ S25089 }),
  .A2({ S25090 }),
  .A3({ S24731 }),
  .ZN({ S25152 })
);
NAND2_X1 #() 
NAND2_X1_4416_ (
  .A1({ S25152 }),
  .A2({ S24776 }),
  .ZN({ S25153 })
);
NAND2_X1 #() 
NAND2_X1_4417_ (
  .A1({ S24748 }),
  .A2({ S25957[1043] }),
  .ZN({ S25154 })
);
NAND2_X1 #() 
NAND2_X1_4418_ (
  .A1({ S25154 }),
  .A2({ S25957[1044] }),
  .ZN({ S25155 })
);
OAI211_X1 #() 
OAI211_X1_1530_ (
  .A({ S25153 }),
  .B({ S22921 }),
  .C1({ S25151 }),
  .C2({ S25155 }),
  .ZN({ S25156 })
);
NAND2_X1 #() 
NAND2_X1_4419_ (
  .A1({ S25085 }),
  .A2({ S25957[1045] }),
  .ZN({ S25157 })
);
NAND3_X1 #() 
NAND3_X1_4818_ (
  .A1({ S25157 }),
  .A2({ S25156 }),
  .A3({ S22832 }),
  .ZN({ S25158 })
);
NAND3_X1 #() 
NAND3_X1_4819_ (
  .A1({ S25158 }),
  .A2({ S25150 }),
  .A3({ S25957[1047] }),
  .ZN({ S25159 })
);
NAND3_X1 #() 
NAND3_X1_4820_ (
  .A1({ S25145 }),
  .A2({ S25159 }),
  .A3({ S25124 }),
  .ZN({ S25160 })
);
NAND3_X1 #() 
NAND3_X1_4821_ (
  .A1({ S25160 }),
  .A2({ S25123 }),
  .A3({ S25073 }),
  .ZN({ S25161 })
);
NAND3_X1 #() 
NAND3_X1_4822_ (
  .A1({ S25099 }),
  .A2({ S25122 }),
  .A3({ S25124 }),
  .ZN({ S25162 })
);
NAND3_X1 #() 
NAND3_X1_4823_ (
  .A1({ S25145 }),
  .A2({ S25159 }),
  .A3({ S25957[1147] }),
  .ZN({ S25163 })
);
NAND3_X1 #() 
NAND3_X1_4824_ (
  .A1({ S25163 }),
  .A2({ S25162 }),
  .A3({ S25957[1211] }),
  .ZN({ S25164 })
);
NAND3_X1 #() 
NAND3_X1_4825_ (
  .A1({ S25161 }),
  .A2({ S25164 }),
  .A3({ S83 }),
  .ZN({ S25165 })
);
NAND2_X1 #() 
NAND2_X1_4420_ (
  .A1({ S22429 }),
  .A2({ S22433 }),
  .ZN({ S25166 })
);
INV_X1 #() 
INV_X1_1435_ (
  .A({ S25166 }),
  .ZN({ S25957[1115] })
);
NAND2_X1 #() 
NAND2_X1_4421_ (
  .A1({ S25957[1115] }),
  .A2({ S25957[1211] }),
  .ZN({ S25167 })
);
NAND2_X1 #() 
NAND2_X1_4422_ (
  .A1({ S25166 }),
  .A2({ S25073 }),
  .ZN({ S25168 })
);
NAND2_X1 #() 
NAND2_X1_4423_ (
  .A1({ S25167 }),
  .A2({ S25168 }),
  .ZN({ S25169 })
);
INV_X1 #() 
INV_X1_1436_ (
  .A({ S25169 }),
  .ZN({ S25957[1083] })
);
NAND3_X1 #() 
NAND3_X1_4826_ (
  .A1({ S25099 }),
  .A2({ S25122 }),
  .A3({ S25957[1243] }),
  .ZN({ S25170 })
);
NAND3_X1 #() 
NAND3_X1_4827_ (
  .A1({ S25145 }),
  .A2({ S25159 }),
  .A3({ S22430 }),
  .ZN({ S25171 })
);
NAND3_X1 #() 
NAND3_X1_4828_ (
  .A1({ S25171 }),
  .A2({ S25170 }),
  .A3({ S25957[1083] }),
  .ZN({ S25172 })
);
AOI21_X1 #() 
AOI21_X1_2424_ (
  .A({ S22430 }),
  .B1({ S25145 }),
  .B2({ S25159 }),
  .ZN({ S25173 })
);
AOI21_X1 #() 
AOI21_X1_2425_ (
  .A({ S25957[1243] }),
  .B1({ S25099 }),
  .B2({ S25122 }),
  .ZN({ S25174 })
);
OAI21_X1 #() 
OAI21_X1_2278_ (
  .A({ S25169 }),
  .B1({ S25173 }),
  .B2({ S25174 }),
  .ZN({ S25175 })
);
NAND3_X1 #() 
NAND3_X1_4829_ (
  .A1({ S25175 }),
  .A2({ S25957[1051] }),
  .A3({ S25172 }),
  .ZN({ S25176 })
);
NAND2_X1 #() 
NAND2_X1_4424_ (
  .A1({ S25176 }),
  .A2({ S25165 }),
  .ZN({ S95 })
);
NAND3_X1 #() 
NAND3_X1_4830_ (
  .A1({ S25175 }),
  .A2({ S83 }),
  .A3({ S25172 }),
  .ZN({ S25177 })
);
NAND3_X1 #() 
NAND3_X1_4831_ (
  .A1({ S25161 }),
  .A2({ S25164 }),
  .A3({ S25957[1051] }),
  .ZN({ S25178 })
);
NAND2_X1 #() 
NAND2_X1_4425_ (
  .A1({ S25177 }),
  .A2({ S25178 }),
  .ZN({ S25957[923] })
);
NAND2_X1 #() 
NAND2_X1_4426_ (
  .A1({ S20021 }),
  .A2({ S20022 }),
  .ZN({ S25179 })
);
INV_X1 #() 
INV_X1_1437_ (
  .A({ S25179 }),
  .ZN({ S25957[1208] })
);
NAND2_X1 #() 
NAND2_X1_4427_ (
  .A1({ S22513 }),
  .A2({ S22517 }),
  .ZN({ S25180 })
);
INV_X1 #() 
INV_X1_1438_ (
  .A({ S25180 }),
  .ZN({ S25957[1112] })
);
NAND2_X1 #() 
NAND2_X1_4428_ (
  .A1({ S25957[1112] }),
  .A2({ S25957[1208] }),
  .ZN({ S25181 })
);
NAND2_X1 #() 
NAND2_X1_4429_ (
  .A1({ S25180 }),
  .A2({ S25179 }),
  .ZN({ S25182 })
);
NAND2_X1 #() 
NAND2_X1_4430_ (
  .A1({ S25181 }),
  .A2({ S25182 }),
  .ZN({ S25183 })
);
INV_X1 #() 
INV_X1_1439_ (
  .A({ S25183 }),
  .ZN({ S25957[1080] })
);
NAND2_X1 #() 
NAND2_X1_4431_ (
  .A1({ S25019 }),
  .A2({ S24776 }),
  .ZN({ S25184 })
);
NAND3_X1 #() 
NAND3_X1_4832_ (
  .A1({ S24746 }),
  .A2({ S25957[1043] }),
  .A3({ S25957[1042] }),
  .ZN({ S25185 })
);
NAND3_X1 #() 
NAND3_X1_4833_ (
  .A1({ S25014 }),
  .A2({ S25957[1044] }),
  .A3({ S25185 }),
  .ZN({ S25186 })
);
OAI21_X1 #() 
OAI21_X1_2279_ (
  .A({ S25186 }),
  .B1({ S24729 }),
  .B2({ S25184 }),
  .ZN({ S25187 })
);
NAND2_X1 #() 
NAND2_X1_4432_ (
  .A1({ S25187 }),
  .A2({ S25957[1045] }),
  .ZN({ S25188 })
);
NAND2_X1 #() 
NAND2_X1_4433_ (
  .A1({ S24746 }),
  .A2({ S24727 }),
  .ZN({ S25189 })
);
NAND2_X1 #() 
NAND2_X1_4434_ (
  .A1({ S24747 }),
  .A2({ S25957[1042] }),
  .ZN({ S25190 })
);
AOI21_X1 #() 
AOI21_X1_2426_ (
  .A({ S25957[1043] }),
  .B1({ S25189 }),
  .B2({ S25190 }),
  .ZN({ S25191 })
);
INV_X1 #() 
INV_X1_1440_ (
  .A({ S25089 }),
  .ZN({ S25192 })
);
OAI21_X1 #() 
OAI21_X1_2280_ (
  .A({ S25957[1044] }),
  .B1({ S25191 }),
  .B2({ S25192 }),
  .ZN({ S25193 })
);
AOI21_X1 #() 
AOI21_X1_2427_ (
  .A({ S25957[1045] }),
  .B1({ S24948 }),
  .B2({ S24776 }),
  .ZN({ S25194 })
);
NAND2_X1 #() 
NAND2_X1_4435_ (
  .A1({ S25193 }),
  .A2({ S25194 }),
  .ZN({ S25195 })
);
NAND3_X1 #() 
NAND3_X1_4834_ (
  .A1({ S25188 }),
  .A2({ S25957[1046] }),
  .A3({ S25195 }),
  .ZN({ S25196 })
);
NAND2_X1 #() 
NAND2_X1_4436_ (
  .A1({ S24736 }),
  .A2({ S24733 }),
  .ZN({ S25197 })
);
AOI21_X1 #() 
AOI21_X1_2428_ (
  .A({ S25197 }),
  .B1({ S24910 }),
  .B2({ S25957[1043] }),
  .ZN({ S25198 })
);
OAI211_X1 #() 
OAI211_X1_1531_ (
  .A({ S24859 }),
  .B({ S25957[1044] }),
  .C1({ S24786 }),
  .C2({ S24888 }),
  .ZN({ S25199 })
);
OAI211_X1 #() 
OAI211_X1_1532_ (
  .A({ S25199 }),
  .B({ S25957[1045] }),
  .C1({ S25198 }),
  .C2({ S25957[1044] }),
  .ZN({ S25200 })
);
OAI221_X1 #() 
OAI221_X1_126_ (
  .A({ S25957[1044] }),
  .B1({ S24840 }),
  .B2({ S23263 }),
  .C1({ S24728 }),
  .C2({ S25957[1043] }),
  .ZN({ S25201 })
);
NAND4_X1 #() 
NAND4_X1_521_ (
  .A1({ S24797 }),
  .A2({ S74 }),
  .A3({ S24798 }),
  .A4({ S24741 }),
  .ZN({ S25202 })
);
INV_X1 #() 
INV_X1_1441_ (
  .A({ S25202 }),
  .ZN({ S25203 })
);
OAI21_X1 #() 
OAI21_X1_2281_ (
  .A({ S24776 }),
  .B1({ S25203 }),
  .B2({ S25140 }),
  .ZN({ S25204 })
);
NAND3_X1 #() 
NAND3_X1_4835_ (
  .A1({ S25204 }),
  .A2({ S25201 }),
  .A3({ S22921 }),
  .ZN({ S25205 })
);
NAND3_X1 #() 
NAND3_X1_4836_ (
  .A1({ S25200 }),
  .A2({ S22832 }),
  .A3({ S25205 }),
  .ZN({ S25206 })
);
NAND3_X1 #() 
NAND3_X1_4837_ (
  .A1({ S25196 }),
  .A2({ S25206 }),
  .A3({ S25957[1047] }),
  .ZN({ S25207 })
);
AOI21_X1 #() 
AOI21_X1_2429_ (
  .A({ S25957[1044] }),
  .B1({ S24851 }),
  .B2({ S24778 }),
  .ZN({ S25208 })
);
AOI22_X1 #() 
AOI22_X1_502_ (
  .A1({ S25208 }),
  .A2({ S24959 }),
  .B1({ S25074 }),
  .B2({ S24836 }),
  .ZN({ S25209 })
);
NAND2_X1 #() 
NAND2_X1_4437_ (
  .A1({ S24730 }),
  .A2({ S74 }),
  .ZN({ S25210 })
);
AND2_X1 #() 
AND2_X1_274_ (
  .A1({ S24816 }),
  .A2({ S25210 }),
  .ZN({ S25211 })
);
AOI21_X1 #() 
AOI21_X1_2430_ (
  .A({ S24776 }),
  .B1({ S25211 }),
  .B2({ S25154 }),
  .ZN({ S25212 })
);
AOI21_X1 #() 
AOI21_X1_2431_ (
  .A({ S74 }),
  .B1({ S24942 }),
  .B2({ S94 }),
  .ZN({ S25213 })
);
AOI21_X1 #() 
AOI21_X1_2432_ (
  .A({ S25957[1043] }),
  .B1({ S24760 }),
  .B2({ S24769 }),
  .ZN({ S25214 })
);
OAI21_X1 #() 
OAI21_X1_2282_ (
  .A({ S24776 }),
  .B1({ S25214 }),
  .B2({ S25213 }),
  .ZN({ S25215 })
);
NAND2_X1 #() 
NAND2_X1_4438_ (
  .A1({ S25215 }),
  .A2({ S22921 }),
  .ZN({ S25216 })
);
OAI22_X1 #() 
OAI22_X1_114_ (
  .A1({ S25212 }),
  .A2({ S25216 }),
  .B1({ S25209 }),
  .B2({ S22921 }),
  .ZN({ S25217 })
);
OAI21_X1 #() 
OAI21_X1_2283_ (
  .A({ S25957[1044] }),
  .B1({ S24838 }),
  .B2({ S24858 }),
  .ZN({ S25218 })
);
AOI22_X1 #() 
AOI22_X1_503_ (
  .A1({ S24851 }),
  .A2({ S24790 }),
  .B1({ S24914 }),
  .B2({ S74 }),
  .ZN({ S25219 })
);
OAI211_X1 #() 
OAI211_X1_1533_ (
  .A({ S25218 }),
  .B({ S22921 }),
  .C1({ S25219 }),
  .C2({ S25957[1044] }),
  .ZN({ S25220 })
);
NAND3_X1 #() 
NAND3_X1_4838_ (
  .A1({ S24745 }),
  .A2({ S25957[1043] }),
  .A3({ S25035 }),
  .ZN({ S25221 })
);
AOI21_X1 #() 
AOI21_X1_2433_ (
  .A({ S24776 }),
  .B1({ S25221 }),
  .B2({ S24870 }),
  .ZN({ S25222 })
);
AOI22_X1 #() 
AOI22_X1_504_ (
  .A1({ S24774 }),
  .A2({ S24775 }),
  .B1({ S20549 }),
  .B2({ S20546 }),
  .ZN({ S25223 })
);
AOI21_X1 #() 
AOI21_X1_2434_ (
  .A({ S22921 }),
  .B1({ S25223 }),
  .B2({ S24796 }),
  .ZN({ S25224 })
);
OAI21_X1 #() 
OAI21_X1_2284_ (
  .A({ S25224 }),
  .B1({ S24895 }),
  .B2({ S24992 }),
  .ZN({ S25225 })
);
OAI211_X1 #() 
OAI211_X1_1534_ (
  .A({ S25220 }),
  .B({ S25957[1046] }),
  .C1({ S25222 }),
  .C2({ S25225 }),
  .ZN({ S25226 })
);
OAI211_X1 #() 
OAI211_X1_1535_ (
  .A({ S20242 }),
  .B({ S25226 }),
  .C1({ S25217 }),
  .C2({ S25957[1046] }),
  .ZN({ S25227 })
);
AOI21_X1 #() 
AOI21_X1_2435_ (
  .A({ S25957[1240] }),
  .B1({ S25227 }),
  .B2({ S25207 }),
  .ZN({ S25228 })
);
AOI21_X1 #() 
AOI21_X1_2436_ (
  .A({ S25957[1043] }),
  .B1({ S24767 }),
  .B2({ S25957[1041] }),
  .ZN({ S25229 })
);
AOI22_X1 #() 
AOI22_X1_505_ (
  .A1({ S25229 }),
  .A2({ S24769 }),
  .B1({ S24857 }),
  .B2({ S24858 }),
  .ZN({ S25230 })
);
NAND4_X1 #() 
NAND4_X1_522_ (
  .A1({ S25002 }),
  .A2({ S24941 }),
  .A3({ S24983 }),
  .A4({ S24776 }),
  .ZN({ S25231 })
);
OAI211_X1 #() 
OAI211_X1_1536_ (
  .A({ S25957[1045] }),
  .B({ S25231 }),
  .C1({ S25230 }),
  .C2({ S24776 }),
  .ZN({ S25232 })
);
NAND2_X1 #() 
NAND2_X1_4439_ (
  .A1({ S24724 }),
  .A2({ S25957[1043] }),
  .ZN({ S25233 })
);
OAI211_X1 #() 
OAI211_X1_1537_ (
  .A({ S25957[1044] }),
  .B({ S25233 }),
  .C1({ S25024 }),
  .C2({ S25957[1043] }),
  .ZN({ S25234 })
);
AOI21_X1 #() 
AOI21_X1_2437_ (
  .A({ S25957[1045] }),
  .B1({ S25114 }),
  .B2({ S25202 }),
  .ZN({ S25235 })
);
NAND2_X1 #() 
NAND2_X1_4440_ (
  .A1({ S25235 }),
  .A2({ S25234 }),
  .ZN({ S25236 })
);
NAND3_X1 #() 
NAND3_X1_4839_ (
  .A1({ S25232 }),
  .A2({ S22832 }),
  .A3({ S25236 }),
  .ZN({ S25237 })
);
AOI22_X1 #() 
AOI22_X1_506_ (
  .A1({ S25187 }),
  .A2({ S25957[1045] }),
  .B1({ S25193 }),
  .B2({ S25194 }),
  .ZN({ S25238 })
);
OAI211_X1 #() 
OAI211_X1_1538_ (
  .A({ S25957[1047] }),
  .B({ S25237 }),
  .C1({ S25238 }),
  .C2({ S22832 }),
  .ZN({ S25239 })
);
NAND2_X1 #() 
NAND2_X1_4441_ (
  .A1({ S25208 }),
  .A2({ S24959 }),
  .ZN({ S25240 })
);
AOI21_X1 #() 
AOI21_X1_2438_ (
  .A({ S22921 }),
  .B1({ S25074 }),
  .B2({ S24836 }),
  .ZN({ S25241 })
);
NAND2_X1 #() 
NAND2_X1_4442_ (
  .A1({ S25241 }),
  .A2({ S25240 }),
  .ZN({ S25242 })
);
NAND4_X1 #() 
NAND4_X1_523_ (
  .A1({ S25154 }),
  .A2({ S25210 }),
  .A3({ S24816 }),
  .A4({ S25957[1044] }),
  .ZN({ S25243 })
);
NAND2_X1 #() 
NAND2_X1_4443_ (
  .A1({ S24942 }),
  .A2({ S94 }),
  .ZN({ S25244 })
);
NAND2_X1 #() 
NAND2_X1_4444_ (
  .A1({ S25244 }),
  .A2({ S25957[1043] }),
  .ZN({ S25245 })
);
OAI211_X1 #() 
OAI211_X1_1539_ (
  .A({ S23263 }),
  .B({ S74 }),
  .C1({ S24767 }),
  .C2({ S24819 }),
  .ZN({ S25246 })
);
NAND3_X1 #() 
NAND3_X1_4840_ (
  .A1({ S25245 }),
  .A2({ S24776 }),
  .A3({ S25246 }),
  .ZN({ S25247 })
);
NAND3_X1 #() 
NAND3_X1_4841_ (
  .A1({ S25243 }),
  .A2({ S22921 }),
  .A3({ S25247 }),
  .ZN({ S25248 })
);
NAND3_X1 #() 
NAND3_X1_4842_ (
  .A1({ S25248 }),
  .A2({ S22832 }),
  .A3({ S25242 }),
  .ZN({ S25249 })
);
NAND2_X1 #() 
NAND2_X1_4445_ (
  .A1({ S24914 }),
  .A2({ S74 }),
  .ZN({ S25250 })
);
NAND3_X1 #() 
NAND3_X1_4843_ (
  .A1({ S25250 }),
  .A2({ S24947 }),
  .A3({ S24776 }),
  .ZN({ S25251 })
);
OAI221_X1 #() 
OAI221_X1_127_ (
  .A({ S25957[1044] }),
  .B1({ S25957[1040] }),
  .B2({ S74 }),
  .C1({ S24904 }),
  .C2({ S24750 }),
  .ZN({ S25252 })
);
AOI21_X1 #() 
AOI21_X1_2439_ (
  .A({ S25957[1045] }),
  .B1({ S25252 }),
  .B2({ S25251 }),
  .ZN({ S25253 })
);
NAND2_X1 #() 
NAND2_X1_4446_ (
  .A1({ S25221 }),
  .A2({ S24870 }),
  .ZN({ S25254 })
);
AOI21_X1 #() 
AOI21_X1_2440_ (
  .A({ S25225 }),
  .B1({ S25254 }),
  .B2({ S25957[1044] }),
  .ZN({ S25255 })
);
OAI21_X1 #() 
OAI21_X1_2285_ (
  .A({ S25957[1046] }),
  .B1({ S25255 }),
  .B2({ S25253 }),
  .ZN({ S25256 })
);
NAND3_X1 #() 
NAND3_X1_4844_ (
  .A1({ S25256 }),
  .A2({ S20242 }),
  .A3({ S25249 }),
  .ZN({ S25257 })
);
AOI21_X1 #() 
AOI21_X1_2441_ (
  .A({ S22514 }),
  .B1({ S25239 }),
  .B2({ S25257 }),
  .ZN({ S25258 })
);
OAI21_X1 #() 
OAI21_X1_2286_ (
  .A({ S25957[1080] }),
  .B1({ S25228 }),
  .B2({ S25258 }),
  .ZN({ S25259 })
);
NAND3_X1 #() 
NAND3_X1_4845_ (
  .A1({ S25239 }),
  .A2({ S25257 }),
  .A3({ S22514 }),
  .ZN({ S25260 })
);
NAND3_X1 #() 
NAND3_X1_4846_ (
  .A1({ S25227 }),
  .A2({ S25207 }),
  .A3({ S25957[1240] }),
  .ZN({ S25261 })
);
NAND3_X1 #() 
NAND3_X1_4847_ (
  .A1({ S25261 }),
  .A2({ S25260 }),
  .A3({ S25183 }),
  .ZN({ S25262 })
);
NAND3_X1 #() 
NAND3_X1_4848_ (
  .A1({ S25259 }),
  .A2({ S24021 }),
  .A3({ S25262 }),
  .ZN({ S25263 })
);
OAI21_X1 #() 
OAI21_X1_2287_ (
  .A({ S25183 }),
  .B1({ S25228 }),
  .B2({ S25258 }),
  .ZN({ S25264 })
);
NAND3_X1 #() 
NAND3_X1_4849_ (
  .A1({ S25261 }),
  .A2({ S25260 }),
  .A3({ S25957[1080] }),
  .ZN({ S25265 })
);
NAND3_X1 #() 
NAND3_X1_4850_ (
  .A1({ S25264 }),
  .A2({ S25957[1048] }),
  .A3({ S25265 }),
  .ZN({ S25266 })
);
NAND2_X1 #() 
NAND2_X1_4447_ (
  .A1({ S25263 }),
  .A2({ S25266 }),
  .ZN({ S25957[920] })
);
NAND3_X1 #() 
NAND3_X1_4851_ (
  .A1({ S24723 }),
  .A2({ S25957[1043] }),
  .A3({ S24732 }),
  .ZN({ S25267 })
);
NAND4_X1 #() 
NAND4_X1_524_ (
  .A1({ S25267 }),
  .A2({ S24870 }),
  .A3({ S24892 }),
  .A4({ S24776 }),
  .ZN({ S25268 })
);
INV_X1 #() 
INV_X1_1442_ (
  .A({ S25268 }),
  .ZN({ S25269 })
);
AOI21_X1 #() 
AOI21_X1_2442_ (
  .A({ S24934 }),
  .B1({ S24905 }),
  .B2({ S24747 }),
  .ZN({ S25270 })
);
OAI21_X1 #() 
OAI21_X1_2288_ (
  .A({ S25957[1044] }),
  .B1({ S24812 }),
  .B2({ S25957[1040] }),
  .ZN({ S25271 })
);
AOI21_X1 #() 
AOI21_X1_2443_ (
  .A({ S25271 }),
  .B1({ S25270 }),
  .B2({ S25957[1043] }),
  .ZN({ S25272 })
);
OAI21_X1 #() 
OAI21_X1_2289_ (
  .A({ S22921 }),
  .B1({ S25272 }),
  .B2({ S25269 }),
  .ZN({ S25273 })
);
AOI21_X1 #() 
AOI21_X1_2444_ (
  .A({ S74 }),
  .B1({ S24745 }),
  .B2({ S25035 }),
  .ZN({ S25274 })
);
OAI211_X1 #() 
OAI211_X1_1540_ (
  .A({ S25093 }),
  .B({ S25957[1044] }),
  .C1({ S24857 }),
  .C2({ S24733 }),
  .ZN({ S25275 })
);
INV_X1 #() 
INV_X1_1443_ (
  .A({ S24809 }),
  .ZN({ S25276 })
);
NAND3_X1 #() 
NAND3_X1_4852_ (
  .A1({ S24812 }),
  .A2({ S24776 }),
  .A3({ S25276 }),
  .ZN({ S25277 })
);
OAI21_X1 #() 
OAI21_X1_2290_ (
  .A({ S25275 }),
  .B1({ S25274 }),
  .B2({ S25277 }),
  .ZN({ S25278 })
);
NAND2_X1 #() 
NAND2_X1_4448_ (
  .A1({ S25278 }),
  .A2({ S25957[1045] }),
  .ZN({ S25279 })
);
NAND3_X1 #() 
NAND3_X1_4853_ (
  .A1({ S25273 }),
  .A2({ S25957[1046] }),
  .A3({ S25279 }),
  .ZN({ S25280 })
);
NAND3_X1 #() 
NAND3_X1_4854_ (
  .A1({ S24837 }),
  .A2({ S74 }),
  .A3({ S24797 }),
  .ZN({ S25281 })
);
NAND3_X1 #() 
NAND3_X1_4855_ (
  .A1({ S24872 }),
  .A2({ S25281 }),
  .A3({ S25957[1044] }),
  .ZN({ S25282 })
);
INV_X1 #() 
INV_X1_1444_ (
  .A({ S25282 }),
  .ZN({ S25283 })
);
AOI22_X1 #() 
AOI22_X1_507_ (
  .A1({ S24981 }),
  .A2({ S25957[1043] }),
  .B1({ S24993 }),
  .B2({ S24992 }),
  .ZN({ S25284 })
);
OAI21_X1 #() 
OAI21_X1_2291_ (
  .A({ S22921 }),
  .B1({ S25284 }),
  .B2({ S25283 }),
  .ZN({ S25285 })
);
AOI21_X1 #() 
AOI21_X1_2445_ (
  .A({ S74 }),
  .B1({ S24960 }),
  .B2({ S24741 }),
  .ZN({ S25286 })
);
OAI21_X1 #() 
OAI21_X1_2292_ (
  .A({ S25957[1044] }),
  .B1({ S25286 }),
  .B2({ S24787 }),
  .ZN({ S25287 })
);
OAI21_X1 #() 
OAI21_X1_2293_ (
  .A({ S25113 }),
  .B1({ S24904 }),
  .B2({ S74 }),
  .ZN({ S25288 })
);
AOI21_X1 #() 
AOI21_X1_2446_ (
  .A({ S22921 }),
  .B1({ S25288 }),
  .B2({ S24776 }),
  .ZN({ S25289 })
);
NAND2_X1 #() 
NAND2_X1_4449_ (
  .A1({ S25287 }),
  .A2({ S25289 }),
  .ZN({ S25290 })
);
NAND3_X1 #() 
NAND3_X1_4856_ (
  .A1({ S25285 }),
  .A2({ S25290 }),
  .A3({ S22832 }),
  .ZN({ S25291 })
);
NAND3_X1 #() 
NAND3_X1_4857_ (
  .A1({ S25280 }),
  .A2({ S25291 }),
  .A3({ S25957[1047] }),
  .ZN({ S25292 })
);
NOR2_X1 #() 
NOR2_X1_1120_ (
  .A1({ S23263 }),
  .A2({ S24762 }),
  .ZN({ S25293 })
);
NOR2_X1 #() 
NOR2_X1_1121_ (
  .A1({ S24874 }),
  .A2({ S25293 }),
  .ZN({ S25294 })
);
NAND3_X1 #() 
NAND3_X1_4858_ (
  .A1({ S24921 }),
  .A2({ S74 }),
  .A3({ S24942 }),
  .ZN({ S25295 })
);
OAI211_X1 #() 
OAI211_X1_1541_ (
  .A({ S25957[1044] }),
  .B({ S25295 }),
  .C1({ S25294 }),
  .C2({ S74 }),
  .ZN({ S25296 })
);
NAND4_X1 #() 
NAND4_X1_525_ (
  .A1({ S24927 }),
  .A2({ S24921 }),
  .A3({ S24798 }),
  .A4({ S24776 }),
  .ZN({ S25297 })
);
AOI21_X1 #() 
AOI21_X1_2447_ (
  .A({ S25957[1044] }),
  .B1({ S24790 }),
  .B2({ S24751 }),
  .ZN({ S25298 })
);
AOI21_X1 #() 
AOI21_X1_2448_ (
  .A({ S25957[1045] }),
  .B1({ S25298 }),
  .B2({ S25089 }),
  .ZN({ S25299 })
);
AOI21_X1 #() 
AOI21_X1_2449_ (
  .A({ S24776 }),
  .B1({ S24751 }),
  .B2({ S24760 }),
  .ZN({ S25300 })
);
AOI21_X1 #() 
AOI21_X1_2450_ (
  .A({ S22921 }),
  .B1({ S25132 }),
  .B2({ S25300 }),
  .ZN({ S25301 })
);
AOI22_X1 #() 
AOI22_X1_508_ (
  .A1({ S25296 }),
  .A2({ S25299 }),
  .B1({ S25297 }),
  .B2({ S25301 }),
  .ZN({ S25302 })
);
OAI21_X1 #() 
OAI21_X1_2294_ (
  .A({ S24776 }),
  .B1({ S24777 }),
  .B2({ S74 }),
  .ZN({ S25303 })
);
OAI22_X1 #() 
OAI22_X1_115_ (
  .A1({ S24738 }),
  .A2({ S25151 }),
  .B1({ S24856 }),
  .B2({ S25303 }),
  .ZN({ S25304 })
);
NAND2_X1 #() 
NAND2_X1_4450_ (
  .A1({ S25304 }),
  .A2({ S22921 }),
  .ZN({ S25305 })
);
AOI21_X1 #() 
AOI21_X1_2451_ (
  .A({ S24776 }),
  .B1({ S25083 }),
  .B2({ S25005 }),
  .ZN({ S25306 })
);
INV_X1 #() 
INV_X1_1445_ (
  .A({ S25306 }),
  .ZN({ S25307 })
);
NAND3_X1 #() 
NAND3_X1_4859_ (
  .A1({ S24805 }),
  .A2({ S25307 }),
  .A3({ S25957[1045] }),
  .ZN({ S25308 })
);
NAND3_X1 #() 
NAND3_X1_4860_ (
  .A1({ S25308 }),
  .A2({ S25305 }),
  .A3({ S22832 }),
  .ZN({ S25309 })
);
OAI211_X1 #() 
OAI211_X1_1542_ (
  .A({ S25309 }),
  .B({ S20242 }),
  .C1({ S25302 }),
  .C2({ S22832 }),
  .ZN({ S25310 })
);
AOI21_X1 #() 
AOI21_X1_2452_ (
  .A({ S25957[1241] }),
  .B1({ S25292 }),
  .B2({ S25310 }),
  .ZN({ S25311 })
);
AND2_X1 #() 
AND2_X1_275_ (
  .A1({ S24993 }),
  .A2({ S24992 }),
  .ZN({ S25312 })
);
OAI21_X1 #() 
OAI21_X1_2295_ (
  .A({ S25282 }),
  .B1({ S25312 }),
  .B2({ S24795 }),
  .ZN({ S25313 })
);
AOI22_X1 #() 
AOI22_X1_509_ (
  .A1({ S25313 }),
  .A2({ S22921 }),
  .B1({ S25287 }),
  .B2({ S25289 }),
  .ZN({ S25314 })
);
NAND2_X1 #() 
NAND2_X1_4451_ (
  .A1({ S25268 }),
  .A2({ S22921 }),
  .ZN({ S25315 })
);
OAI211_X1 #() 
OAI211_X1_1543_ (
  .A({ S25275 }),
  .B({ S25957[1045] }),
  .C1({ S25274 }),
  .C2({ S25277 }),
  .ZN({ S25316 })
);
OAI211_X1 #() 
OAI211_X1_1544_ (
  .A({ S25316 }),
  .B({ S25957[1046] }),
  .C1({ S25272 }),
  .C2({ S25315 }),
  .ZN({ S25317 })
);
OAI211_X1 #() 
OAI211_X1_1545_ (
  .A({ S25957[1047] }),
  .B({ S25317 }),
  .C1({ S25314 }),
  .C2({ S25957[1046] }),
  .ZN({ S25318 })
);
AOI22_X1 #() 
AOI22_X1_510_ (
  .A1({ S24736 }),
  .A2({ S24742 }),
  .B1({ S24735 }),
  .B2({ S25957[1041] }),
  .ZN({ S25319 })
);
NOR3_X1 #() 
NOR3_X1_150_ (
  .A1({ S25274 }),
  .A2({ S25319 }),
  .A3({ S24776 }),
  .ZN({ S25320 })
);
NAND2_X1 #() 
NAND2_X1_4452_ (
  .A1({ S25298 }),
  .A2({ S25089 }),
  .ZN({ S25321 })
);
NAND2_X1 #() 
NAND2_X1_4453_ (
  .A1({ S25321 }),
  .A2({ S22921 }),
  .ZN({ S25322 })
);
NAND2_X1 #() 
NAND2_X1_4454_ (
  .A1({ S25132 }),
  .A2({ S25300 }),
  .ZN({ S25323 })
);
NAND3_X1 #() 
NAND3_X1_4861_ (
  .A1({ S25323 }),
  .A2({ S25957[1045] }),
  .A3({ S25297 }),
  .ZN({ S25324 })
);
OAI211_X1 #() 
OAI211_X1_1546_ (
  .A({ S25957[1046] }),
  .B({ S25324 }),
  .C1({ S25320 }),
  .C2({ S25322 }),
  .ZN({ S25325 })
);
OAI21_X1 #() 
OAI21_X1_2296_ (
  .A({ S25957[1045] }),
  .B1({ S24804 }),
  .B2({ S25306 }),
  .ZN({ S25326 })
);
OAI211_X1 #() 
OAI211_X1_1547_ (
  .A({ S25326 }),
  .B({ S22832 }),
  .C1({ S25957[1045] }),
  .C2({ S25304 }),
  .ZN({ S25327 })
);
NAND3_X1 #() 
NAND3_X1_4862_ (
  .A1({ S25325 }),
  .A2({ S25327 }),
  .A3({ S20242 }),
  .ZN({ S25328 })
);
AOI21_X1 #() 
AOI21_X1_2453_ (
  .A({ S24015 }),
  .B1({ S25318 }),
  .B2({ S25328 }),
  .ZN({ S25329 })
);
OAI21_X1 #() 
OAI21_X1_2297_ (
  .A({ S21399 }),
  .B1({ S25329 }),
  .B2({ S25311 }),
  .ZN({ S25330 })
);
AOI21_X1 #() 
AOI21_X1_2454_ (
  .A({ S25957[1046] }),
  .B1({ S25285 }),
  .B2({ S25290 }),
  .ZN({ S25331 })
);
NAND2_X1 #() 
NAND2_X1_4455_ (
  .A1({ S25317 }),
  .A2({ S25957[1047] }),
  .ZN({ S25332 })
);
OAI211_X1 #() 
OAI211_X1_1548_ (
  .A({ S25328 }),
  .B({ S24015 }),
  .C1({ S25332 }),
  .C2({ S25331 }),
  .ZN({ S25333 })
);
NAND3_X1 #() 
NAND3_X1_4863_ (
  .A1({ S25292 }),
  .A2({ S25310 }),
  .A3({ S25957[1241] }),
  .ZN({ S25334 })
);
NAND3_X1 #() 
NAND3_X1_4864_ (
  .A1({ S25334 }),
  .A2({ S25333 }),
  .A3({ S25957[1177] }),
  .ZN({ S25335 })
);
NAND2_X1 #() 
NAND2_X1_4456_ (
  .A1({ S25330 }),
  .A2({ S25335 }),
  .ZN({ S25957[921] })
);
NOR2_X1 #() 
NOR2_X1_1122_ (
  .A1({ S22623 }),
  .A2({ S22624 }),
  .ZN({ S25957[1114] })
);
NAND2_X1 #() 
NAND2_X1_4457_ (
  .A1({ S22614 }),
  .A2({ S22612 }),
  .ZN({ S25957[1146] })
);
INV_X1 #() 
INV_X1_1446_ (
  .A({ S25957[1146] }),
  .ZN({ S25336 })
);
AOI21_X1 #() 
AOI21_X1_2455_ (
  .A({ S24750 }),
  .B1({ S24811 }),
  .B2({ S94 }),
  .ZN({ S25337 })
);
NOR2_X1 #() 
NOR2_X1_1123_ (
  .A1({ S24802 }),
  .A2({ S24776 }),
  .ZN({ S25338 })
);
OAI21_X1 #() 
OAI21_X1_2298_ (
  .A({ S25338 }),
  .B1({ S25337 }),
  .B2({ S25957[1043] }),
  .ZN({ S25339 })
);
NAND2_X1 #() 
NAND2_X1_4458_ (
  .A1({ S24746 }),
  .A2({ S25957[1042] }),
  .ZN({ S25340 })
);
NAND3_X1 #() 
NAND3_X1_4865_ (
  .A1({ S24728 }),
  .A2({ S25957[1043] }),
  .A3({ S25340 }),
  .ZN({ S25341 })
);
AOI21_X1 #() 
AOI21_X1_2456_ (
  .A({ S22921 }),
  .B1({ S25341 }),
  .B2({ S24957 }),
  .ZN({ S25342 })
);
NAND2_X1 #() 
NAND2_X1_4459_ (
  .A1({ S25342 }),
  .A2({ S25339 }),
  .ZN({ S25343 })
);
NAND3_X1 #() 
NAND3_X1_4866_ (
  .A1({ S24728 }),
  .A2({ S25957[1043] }),
  .A3({ S25190 }),
  .ZN({ S25344 })
);
NAND2_X1 #() 
NAND2_X1_4460_ (
  .A1({ S25344 }),
  .A2({ S24919 }),
  .ZN({ S25345 })
);
AOI21_X1 #() 
AOI21_X1_2457_ (
  .A({ S25957[1044] }),
  .B1({ S24730 }),
  .B2({ S74 }),
  .ZN({ S25346 })
);
AOI21_X1 #() 
AOI21_X1_2458_ (
  .A({ S25957[1045] }),
  .B1({ S25346 }),
  .B2({ S24813 }),
  .ZN({ S25347 })
);
NAND2_X1 #() 
NAND2_X1_4461_ (
  .A1({ S25345 }),
  .A2({ S25347 }),
  .ZN({ S25348 })
);
NAND3_X1 #() 
NAND3_X1_4867_ (
  .A1({ S25343 }),
  .A2({ S25957[1046] }),
  .A3({ S25348 }),
  .ZN({ S25349 })
);
NAND3_X1 #() 
NAND3_X1_4868_ (
  .A1({ S24777 }),
  .A2({ S25957[1043] }),
  .A3({ S25957[1040] }),
  .ZN({ S25350 })
);
NAND3_X1 #() 
NAND3_X1_4869_ (
  .A1({ S25116 }),
  .A2({ S25350 }),
  .A3({ S25957[1044] }),
  .ZN({ S25351 })
);
OAI211_X1 #() 
OAI211_X1_1549_ (
  .A({ S24746 }),
  .B({ S25957[1043] }),
  .C1({ S24747 }),
  .C2({ S24727 }),
  .ZN({ S25352 })
);
NAND3_X1 #() 
NAND3_X1_4870_ (
  .A1({ S25352 }),
  .A2({ S24776 }),
  .A3({ S25032 }),
  .ZN({ S25353 })
);
NAND3_X1 #() 
NAND3_X1_4871_ (
  .A1({ S25353 }),
  .A2({ S25957[1045] }),
  .A3({ S25351 }),
  .ZN({ S25354 })
);
NAND2_X1 #() 
NAND2_X1_4462_ (
  .A1({ S24761 }),
  .A2({ S74 }),
  .ZN({ S25355 })
);
NAND3_X1 #() 
NAND3_X1_4872_ (
  .A1({ S25957[1043] }),
  .A2({ S25957[1041] }),
  .A3({ S24762 }),
  .ZN({ S25356 })
);
NAND3_X1 #() 
NAND3_X1_4873_ (
  .A1({ S25356 }),
  .A2({ S25355 }),
  .A3({ S25957[1044] }),
  .ZN({ S25357 })
);
OAI211_X1 #() 
OAI211_X1_1550_ (
  .A({ S25357 }),
  .B({ S22921 }),
  .C1({ S24841 }),
  .C2({ S25957[1044] }),
  .ZN({ S25358 })
);
NAND3_X1 #() 
NAND3_X1_4874_ (
  .A1({ S25354 }),
  .A2({ S25358 }),
  .A3({ S22832 }),
  .ZN({ S25359 })
);
NAND3_X1 #() 
NAND3_X1_4875_ (
  .A1({ S25349 }),
  .A2({ S25957[1047] }),
  .A3({ S25359 }),
  .ZN({ S25360 })
);
AOI21_X1 #() 
AOI21_X1_2459_ (
  .A({ S24776 }),
  .B1({ S24996 }),
  .B2({ S25356 }),
  .ZN({ S25361 })
);
NAND2_X1 #() 
NAND2_X1_4463_ (
  .A1({ S24728 }),
  .A2({ S24724 }),
  .ZN({ S25362 })
);
INV_X1 #() 
INV_X1_1447_ (
  .A({ S25223 }),
  .ZN({ S25363 })
);
OAI21_X1 #() 
OAI21_X1_2299_ (
  .A({ S24896 }),
  .B1({ S25362 }),
  .B2({ S25363 }),
  .ZN({ S25364 })
);
OAI21_X1 #() 
OAI21_X1_2300_ (
  .A({ S22921 }),
  .B1({ S25361 }),
  .B2({ S25364 }),
  .ZN({ S25365 })
);
AOI21_X1 #() 
AOI21_X1_2460_ (
  .A({ S24776 }),
  .B1({ S24921 }),
  .B2({ S24808 }),
  .ZN({ S25366 })
);
NAND2_X1 #() 
NAND2_X1_4464_ (
  .A1({ S25079 }),
  .A2({ S25366 }),
  .ZN({ S25367 })
);
AOI221_X4 #() 
AOI221_X4_1_ (
  .A({ S22921 }),
  .B1({ S25223 }),
  .B2({ S24837 }),
  .C1({ S24943 }),
  .C2({ S24894 }),
  .ZN({ S25368 })
);
AOI21_X1 #() 
AOI21_X1_2461_ (
  .A({ S25957[1046] }),
  .B1({ S25368 }),
  .B2({ S25367 }),
  .ZN({ S25369 })
);
NAND2_X1 #() 
NAND2_X1_4465_ (
  .A1({ S25365 }),
  .A2({ S25369 }),
  .ZN({ S25370 })
);
NAND3_X1 #() 
NAND3_X1_4876_ (
  .A1({ S24728 }),
  .A2({ S24960 }),
  .A3({ S25957[1043] }),
  .ZN({ S25371 })
);
AOI21_X1 #() 
AOI21_X1_2462_ (
  .A({ S25957[1044] }),
  .B1({ S24809 }),
  .B2({ S24761 }),
  .ZN({ S25372 })
);
OAI21_X1 #() 
OAI21_X1_2301_ (
  .A({ S25118 }),
  .B1({ S24778 }),
  .B2({ S74 }),
  .ZN({ S25373 })
);
AOI22_X1 #() 
AOI22_X1_511_ (
  .A1({ S25372 }),
  .A2({ S25371 }),
  .B1({ S25373 }),
  .B2({ S25957[1044] }),
  .ZN({ S25374 })
);
NAND2_X1 #() 
NAND2_X1_4466_ (
  .A1({ S24863 }),
  .A2({ S74 }),
  .ZN({ S25375 })
);
AOI21_X1 #() 
AOI21_X1_2463_ (
  .A({ S25957[1044] }),
  .B1({ S24780 }),
  .B2({ S25957[1043] }),
  .ZN({ S25376 })
);
NAND3_X1 #() 
NAND3_X1_4877_ (
  .A1({ S25375 }),
  .A2({ S25210 }),
  .A3({ S25376 }),
  .ZN({ S25377 })
);
OAI21_X1 #() 
OAI21_X1_2302_ (
  .A({ S74 }),
  .B1({ S24811 }),
  .B2({ S24986 }),
  .ZN({ S25378 })
);
AOI21_X1 #() 
AOI21_X1_2464_ (
  .A({ S24776 }),
  .B1({ S24808 }),
  .B2({ S24837 }),
  .ZN({ S25379 })
);
NAND2_X1 #() 
NAND2_X1_4467_ (
  .A1({ S25378 }),
  .A2({ S25379 }),
  .ZN({ S25380 })
);
NAND3_X1 #() 
NAND3_X1_4878_ (
  .A1({ S25380 }),
  .A2({ S25377 }),
  .A3({ S22921 }),
  .ZN({ S25381 })
);
OAI211_X1 #() 
OAI211_X1_1551_ (
  .A({ S25381 }),
  .B({ S25957[1046] }),
  .C1({ S25374 }),
  .C2({ S22921 }),
  .ZN({ S25382 })
);
NAND3_X1 #() 
NAND3_X1_4879_ (
  .A1({ S25370 }),
  .A2({ S25382 }),
  .A3({ S20242 }),
  .ZN({ S25383 })
);
NAND3_X1 #() 
NAND3_X1_4880_ (
  .A1({ S25383 }),
  .A2({ S25336 }),
  .A3({ S25360 }),
  .ZN({ S25384 })
);
INV_X1 #() 
INV_X1_1448_ (
  .A({ S25372 }),
  .ZN({ S25385 })
);
AOI21_X1 #() 
AOI21_X1_2465_ (
  .A({ S74 }),
  .B1({ S23263 }),
  .B2({ S24732 }),
  .ZN({ S25386 })
);
OAI21_X1 #() 
OAI21_X1_2303_ (
  .A({ S25957[1044] }),
  .B1({ S25127 }),
  .B2({ S25386 }),
  .ZN({ S25387 })
);
OAI21_X1 #() 
OAI21_X1_2304_ (
  .A({ S25387 }),
  .B1({ S24749 }),
  .B2({ S25385 }),
  .ZN({ S25388 })
);
AOI21_X1 #() 
AOI21_X1_2466_ (
  .A({ S25957[1045] }),
  .B1({ S24987 }),
  .B2({ S25376 }),
  .ZN({ S25389 })
);
AOI22_X1 #() 
AOI22_X1_512_ (
  .A1({ S25388 }),
  .A2({ S25957[1045] }),
  .B1({ S25389 }),
  .B2({ S25380 }),
  .ZN({ S25390 })
);
AOI22_X1 #() 
AOI22_X1_513_ (
  .A1({ S25390 }),
  .A2({ S25957[1046] }),
  .B1({ S25365 }),
  .B2({ S25369 }),
  .ZN({ S25391 })
);
AOI22_X1 #() 
AOI22_X1_514_ (
  .A1({ S25342 }),
  .A2({ S25339 }),
  .B1({ S25347 }),
  .B2({ S25345 }),
  .ZN({ S25392 })
);
NAND2_X1 #() 
NAND2_X1_4468_ (
  .A1({ S25354 }),
  .A2({ S25358 }),
  .ZN({ S25393 })
);
NAND2_X1 #() 
NAND2_X1_4469_ (
  .A1({ S25393 }),
  .A2({ S22832 }),
  .ZN({ S25394 })
);
OAI211_X1 #() 
OAI211_X1_1552_ (
  .A({ S25394 }),
  .B({ S25957[1047] }),
  .C1({ S22832 }),
  .C2({ S25392 }),
  .ZN({ S25395 })
);
OAI211_X1 #() 
OAI211_X1_1553_ (
  .A({ S25395 }),
  .B({ S25957[1146] }),
  .C1({ S25391 }),
  .C2({ S25957[1047] }),
  .ZN({ S25396 })
);
NAND3_X1 #() 
NAND3_X1_4881_ (
  .A1({ S25396 }),
  .A2({ S25957[1114] }),
  .A3({ S25384 }),
  .ZN({ S25397 })
);
INV_X1 #() 
INV_X1_1449_ (
  .A({ S25957[1114] }),
  .ZN({ S25398 })
);
NAND3_X1 #() 
NAND3_X1_4882_ (
  .A1({ S25383 }),
  .A2({ S25957[1146] }),
  .A3({ S25360 }),
  .ZN({ S25399 })
);
OAI211_X1 #() 
OAI211_X1_1554_ (
  .A({ S25395 }),
  .B({ S25336 }),
  .C1({ S25391 }),
  .C2({ S25957[1047] }),
  .ZN({ S25400 })
);
NAND3_X1 #() 
NAND3_X1_4883_ (
  .A1({ S25400 }),
  .A2({ S25398 }),
  .A3({ S25399 }),
  .ZN({ S25401 })
);
NAND3_X1 #() 
NAND3_X1_4884_ (
  .A1({ S25397 }),
  .A2({ S25401 }),
  .A3({ S21411 }),
  .ZN({ S25402 })
);
NAND3_X1 #() 
NAND3_X1_4885_ (
  .A1({ S25396 }),
  .A2({ S25398 }),
  .A3({ S25384 }),
  .ZN({ S25403 })
);
NAND3_X1 #() 
NAND3_X1_4886_ (
  .A1({ S25400 }),
  .A2({ S25957[1114] }),
  .A3({ S25399 }),
  .ZN({ S25404 })
);
NAND3_X1 #() 
NAND3_X1_4887_ (
  .A1({ S25403 }),
  .A2({ S25404 }),
  .A3({ S25957[1178] }),
  .ZN({ S25405 })
);
NAND2_X1 #() 
NAND2_X1_4470_ (
  .A1({ S25402 }),
  .A2({ S25405 }),
  .ZN({ S25957[922] })
);
AOI21_X1 #() 
AOI21_X1_2467_ (
  .A({ S20144 }),
  .B1({ S23874 }),
  .B2({ S23875 }),
  .ZN({ S25406 })
);
AND3_X1 #() 
AND3_X1_175_ (
  .A1({ S23874 }),
  .A2({ S23875 }),
  .A3({ S20144 }),
  .ZN({ S25407 })
);
NOR2_X1 #() 
NOR2_X1_1124_ (
  .A1({ S25407 }),
  .A2({ S25406 }),
  .ZN({ S25408 })
);
AOI21_X1 #() 
AOI21_X1_2468_ (
  .A({ S25408 }),
  .B1({ S23922 }),
  .B2({ S23925 }),
  .ZN({ S96 })
);
NAND3_X1 #() 
NAND3_X1_4888_ (
  .A1({ S25408 }),
  .A2({ S23922 }),
  .A3({ S23925 }),
  .ZN({ S97 })
);
INV_X1 #() 
INV_X1_1450_ (
  .A({ S25957[1196] }),
  .ZN({ S25409 })
);
NAND2_X1 #() 
NAND2_X1_4471_ (
  .A1({ S23708 }),
  .A2({ S23688 }),
  .ZN({ S25957[1004] })
);
NAND2_X1 #() 
NAND2_X1_4472_ (
  .A1({ S25957[1004] }),
  .A2({ S25409 }),
  .ZN({ S25410 })
);
NAND3_X1 #() 
NAND3_X1_4889_ (
  .A1({ S23708 }),
  .A2({ S23688 }),
  .A3({ S25957[1196] }),
  .ZN({ S25411 })
);
NAND3_X1 #() 
NAND3_X1_4890_ (
  .A1({ S25410 }),
  .A2({ S25411 }),
  .A3({ S22636 }),
  .ZN({ S25412 })
);
NAND3_X1 #() 
NAND3_X1_4891_ (
  .A1({ S23708 }),
  .A2({ S23688 }),
  .A3({ S25409 }),
  .ZN({ S25413 })
);
NAND2_X1 #() 
NAND2_X1_4473_ (
  .A1({ S25957[1004] }),
  .A2({ S25957[1196] }),
  .ZN({ S25414 })
);
NAND3_X1 #() 
NAND3_X1_4892_ (
  .A1({ S25414 }),
  .A2({ S25957[1036] }),
  .A3({ S25413 }),
  .ZN({ S25415 })
);
NAND2_X1 #() 
NAND2_X1_4474_ (
  .A1({ S25412 }),
  .A2({ S25415 }),
  .ZN({ S25416 })
);
NAND2_X1 #() 
NAND2_X1_4475_ (
  .A1({ S25957[906] }),
  .A2({ S25957[905] }),
  .ZN({ S25417 })
);
INV_X1 #() 
INV_X1_1451_ (
  .A({ S25417 }),
  .ZN({ S25418 })
);
AOI21_X1 #() 
AOI21_X1_2469_ (
  .A({ S25957[1033] }),
  .B1({ S23923 }),
  .B2({ S23924 }),
  .ZN({ S25419 })
);
AOI21_X1 #() 
AOI21_X1_2470_ (
  .A({ S22634 }),
  .B1({ S23921 }),
  .B2({ S23917 }),
  .ZN({ S25420 })
);
OAI21_X1 #() 
OAI21_X1_2305_ (
  .A({ S25408 }),
  .B1({ S25419 }),
  .B2({ S25420 }),
  .ZN({ S25421 })
);
NAND3_X1 #() 
NAND3_X1_4893_ (
  .A1({ S23922 }),
  .A2({ S23925 }),
  .A3({ S25957[904] }),
  .ZN({ S25422 })
);
AOI21_X1 #() 
AOI21_X1_2471_ (
  .A({ S25957[906] }),
  .B1({ S25421 }),
  .B2({ S25422 }),
  .ZN({ S25423 })
);
OAI21_X1 #() 
OAI21_X1_2306_ (
  .A({ S89 }),
  .B1({ S25423 }),
  .B2({ S25418 }),
  .ZN({ S25424 })
);
NOR2_X1 #() 
NOR2_X1_1125_ (
  .A1({ S25957[906] }),
  .A2({ S25957[905] }),
  .ZN({ S25425 })
);
NAND2_X1 #() 
NAND2_X1_4476_ (
  .A1({ S25425 }),
  .A2({ S25957[907] }),
  .ZN({ S25426 })
);
NAND3_X1 #() 
NAND3_X1_4894_ (
  .A1({ S24009 }),
  .A2({ S24006 }),
  .A3({ S22644 }),
  .ZN({ S25427 })
);
NAND3_X1 #() 
NAND3_X1_4895_ (
  .A1({ S24011 }),
  .A2({ S24012 }),
  .A3({ S25957[1034] }),
  .ZN({ S25428 })
);
NAND3_X1 #() 
NAND3_X1_4896_ (
  .A1({ S25408 }),
  .A2({ S25427 }),
  .A3({ S25428 }),
  .ZN({ S25429 })
);
NAND2_X1 #() 
NAND2_X1_4477_ (
  .A1({ S25429 }),
  .A2({ S89 }),
  .ZN({ S25430 })
);
AOI21_X1 #() 
AOI21_X1_2472_ (
  .A({ S25957[908] }),
  .B1({ S25426 }),
  .B2({ S25430 }),
  .ZN({ S25431 })
);
NAND2_X1 #() 
NAND2_X1_4478_ (
  .A1({ S25431 }),
  .A2({ S25424 }),
  .ZN({ S25432 })
);
NAND3_X1 #() 
NAND3_X1_4897_ (
  .A1({ S24010 }),
  .A2({ S24013 }),
  .A3({ S25957[904] }),
  .ZN({ S25433 })
);
NAND2_X1 #() 
NAND2_X1_4479_ (
  .A1({ S25433 }),
  .A2({ S89 }),
  .ZN({ S25434 })
);
NAND3_X1 #() 
NAND3_X1_4898_ (
  .A1({ S25421 }),
  .A2({ S25957[906] }),
  .A3({ S25422 }),
  .ZN({ S25435 })
);
NAND2_X1 #() 
NAND2_X1_4480_ (
  .A1({ S25427 }),
  .A2({ S25428 }),
  .ZN({ S25436 })
);
OAI21_X1 #() 
OAI21_X1_2307_ (
  .A({ S25957[904] }),
  .B1({ S25419 }),
  .B2({ S25420 }),
  .ZN({ S25437 })
);
NAND3_X1 #() 
NAND3_X1_4899_ (
  .A1({ S25437 }),
  .A2({ S25436 }),
  .A3({ S97 }),
  .ZN({ S25438 })
);
NAND3_X1 #() 
NAND3_X1_4900_ (
  .A1({ S25435 }),
  .A2({ S25438 }),
  .A3({ S25957[907] }),
  .ZN({ S25439 })
);
OAI21_X1 #() 
OAI21_X1_2308_ (
  .A({ S25439 }),
  .B1({ S25418 }),
  .B2({ S25434 }),
  .ZN({ S25440 })
);
OAI21_X1 #() 
OAI21_X1_2309_ (
  .A({ S25432 }),
  .B1({ S25440 }),
  .B2({ S25416 }),
  .ZN({ S25441 })
);
NAND3_X1 #() 
NAND3_X1_4901_ (
  .A1({ S25427 }),
  .A2({ S25428 }),
  .A3({ S25957[904] }),
  .ZN({ S25442 })
);
AOI22_X1 #() 
AOI22_X1_515_ (
  .A1({ S23794 }),
  .A2({ S23786 }),
  .B1({ S23922 }),
  .B2({ S23925 }),
  .ZN({ S25443 })
);
NOR2_X1 #() 
NOR2_X1_1126_ (
  .A1({ S25419 }),
  .A2({ S25420 }),
  .ZN({ S25444 })
);
NAND2_X1 #() 
NAND2_X1_4481_ (
  .A1({ S25444 }),
  .A2({ S25957[907] }),
  .ZN({ S25445 })
);
NAND3_X1 #() 
NAND3_X1_4902_ (
  .A1({ S25957[906] }),
  .A2({ S25957[907] }),
  .A3({ S25957[904] }),
  .ZN({ S25446 })
);
NAND3_X1 #() 
NAND3_X1_4903_ (
  .A1({ S25445 }),
  .A2({ S25446 }),
  .A3({ S25957[908] }),
  .ZN({ S25447 })
);
AOI21_X1 #() 
AOI21_X1_2473_ (
  .A({ S25447 }),
  .B1({ S25443 }),
  .B2({ S25442 }),
  .ZN({ S25448 })
);
OAI21_X1 #() 
OAI21_X1_2310_ (
  .A({ S89 }),
  .B1({ S97 }),
  .B2({ S25957[906] }),
  .ZN({ S25449 })
);
AOI21_X1 #() 
AOI21_X1_2474_ (
  .A({ S25957[908] }),
  .B1({ S96 }),
  .B2({ S25957[907] }),
  .ZN({ S25450 })
);
NAND2_X1 #() 
NAND2_X1_4482_ (
  .A1({ S25450 }),
  .A2({ S25449 }),
  .ZN({ S25451 })
);
NAND2_X1 #() 
NAND2_X1_4483_ (
  .A1({ S25451 }),
  .A2({ S25957[909] }),
  .ZN({ S25452 })
);
OAI221_X1 #() 
OAI221_X1_128_ (
  .A({ S23551 }),
  .B1({ S25448 }),
  .B2({ S25452 }),
  .C1({ S25441 }),
  .C2({ S25957[909] }),
  .ZN({ S25453 })
);
NOR2_X1 #() 
NOR2_X1_1127_ (
  .A1({ S89 }),
  .A2({ S25957[905] }),
  .ZN({ S25454 })
);
NAND2_X1 #() 
NAND2_X1_4484_ (
  .A1({ S97 }),
  .A2({ S25957[906] }),
  .ZN({ S25455 })
);
AOI21_X1 #() 
AOI21_X1_2475_ (
  .A({ S25957[904] }),
  .B1({ S25427 }),
  .B2({ S25428 }),
  .ZN({ S25456 })
);
NAND2_X1 #() 
NAND2_X1_4485_ (
  .A1({ S25456 }),
  .A2({ S25444 }),
  .ZN({ S25457 })
);
NAND2_X1 #() 
NAND2_X1_4486_ (
  .A1({ S25457 }),
  .A2({ S25455 }),
  .ZN({ S25458 })
);
AOI21_X1 #() 
AOI21_X1_2476_ (
  .A({ S25458 }),
  .B1({ S25454 }),
  .B2({ S25957[904] }),
  .ZN({ S25459 })
);
AOI21_X1 #() 
AOI21_X1_2477_ (
  .A({ S25957[904] }),
  .B1({ S23922 }),
  .B2({ S23925 }),
  .ZN({ S25460 })
);
NOR2_X1 #() 
NOR2_X1_1128_ (
  .A1({ S25460 }),
  .A2({ S25957[907] }),
  .ZN({ S25461 })
);
INV_X1 #() 
INV_X1_1452_ (
  .A({ S25461 }),
  .ZN({ S25462 })
);
NAND4_X1 #() 
NAND4_X1_526_ (
  .A1({ S25427 }),
  .A2({ S25428 }),
  .A3({ S23922 }),
  .A4({ S23925 }),
  .ZN({ S25463 })
);
NAND2_X1 #() 
NAND2_X1_4487_ (
  .A1({ S25463 }),
  .A2({ S25957[907] }),
  .ZN({ S25464 })
);
INV_X1 #() 
INV_X1_1453_ (
  .A({ S25464 }),
  .ZN({ S25465 })
);
NAND2_X1 #() 
NAND2_X1_4488_ (
  .A1({ S25465 }),
  .A2({ S25437 }),
  .ZN({ S25466 })
);
NAND3_X1 #() 
NAND3_X1_4904_ (
  .A1({ S25466 }),
  .A2({ S25957[908] }),
  .A3({ S25462 }),
  .ZN({ S25467 })
);
OAI21_X1 #() 
OAI21_X1_2311_ (
  .A({ S25467 }),
  .B1({ S25459 }),
  .B2({ S25957[908] }),
  .ZN({ S25468 })
);
NAND3_X1 #() 
NAND3_X1_4905_ (
  .A1({ S25408 }),
  .A2({ S24010 }),
  .A3({ S24013 }),
  .ZN({ S25469 })
);
NOR2_X1 #() 
NOR2_X1_1129_ (
  .A1({ S25442 }),
  .A2({ S89 }),
  .ZN({ S25470 })
);
NAND3_X1 #() 
NAND3_X1_4906_ (
  .A1({ S25422 }),
  .A2({ S25436 }),
  .A3({ S25957[907] }),
  .ZN({ S25471 })
);
NAND2_X1 #() 
NAND2_X1_4489_ (
  .A1({ S25471 }),
  .A2({ S25957[908] }),
  .ZN({ S25472 })
);
AOI211_X1 #() 
AOI211_X1_79_ (
  .A({ S25470 }),
  .B({ S25472 }),
  .C1({ S25443 }),
  .C2({ S25469 }),
  .ZN({ S25473 })
);
NAND2_X1 #() 
NAND2_X1_4490_ (
  .A1({ S25437 }),
  .A2({ S97 }),
  .ZN({ S25474 })
);
AOI22_X1 #() 
AOI22_X1_516_ (
  .A1({ S25436 }),
  .A2({ S25957[905] }),
  .B1({ S23796 }),
  .B2({ S23795 }),
  .ZN({ S25475 })
);
INV_X1 #() 
INV_X1_1454_ (
  .A({ S25475 }),
  .ZN({ S25476 })
);
NAND2_X1 #() 
NAND2_X1_4491_ (
  .A1({ S25437 }),
  .A2({ S25429 }),
  .ZN({ S25477 })
);
AOI21_X1 #() 
AOI21_X1_2478_ (
  .A({ S25957[907] }),
  .B1({ S25957[905] }),
  .B2({ S25957[906] }),
  .ZN({ S25478 })
);
NAND2_X1 #() 
NAND2_X1_4492_ (
  .A1({ S25478 }),
  .A2({ S25477 }),
  .ZN({ S25479 })
);
OAI21_X1 #() 
OAI21_X1_2312_ (
  .A({ S25479 }),
  .B1({ S25474 }),
  .B2({ S25476 }),
  .ZN({ S25480 })
);
OAI21_X1 #() 
OAI21_X1_2313_ (
  .A({ S25957[909] }),
  .B1({ S25480 }),
  .B2({ S25957[908] }),
  .ZN({ S25481 })
);
OAI221_X1 #() 
OAI221_X1_129_ (
  .A({ S25957[910] }),
  .B1({ S25481 }),
  .B2({ S25473 }),
  .C1({ S25957[909] }),
  .C2({ S25468 }),
  .ZN({ S25482 })
);
AND3_X1 #() 
AND3_X1_176_ (
  .A1({ S25453 }),
  .A2({ S25482 }),
  .A3({ S25957[911] }),
  .ZN({ S25483 })
);
AND2_X1 #() 
AND2_X1_276_ (
  .A1({ S23629 }),
  .A2({ S23626 }),
  .ZN({ S25484 })
);
NAND2_X1 #() 
NAND2_X1_4493_ (
  .A1({ S25437 }),
  .A2({ S25957[906] }),
  .ZN({ S25485 })
);
NAND2_X1 #() 
NAND2_X1_4494_ (
  .A1({ S25422 }),
  .A2({ S25436 }),
  .ZN({ S25486 })
);
NAND2_X1 #() 
NAND2_X1_4495_ (
  .A1({ S25485 }),
  .A2({ S25486 }),
  .ZN({ S25487 })
);
AOI21_X1 #() 
AOI21_X1_2479_ (
  .A({ S25957[908] }),
  .B1({ S25487 }),
  .B2({ S89 }),
  .ZN({ S25488 })
);
INV_X1 #() 
INV_X1_1455_ (
  .A({ S25488 }),
  .ZN({ S25489 })
);
AOI21_X1 #() 
AOI21_X1_2480_ (
  .A({ S25489 }),
  .B1({ S25475 }),
  .B2({ S25442 }),
  .ZN({ S25490 })
);
NAND3_X1 #() 
NAND3_X1_4907_ (
  .A1({ S25437 }),
  .A2({ S25957[906] }),
  .A3({ S97 }),
  .ZN({ S25491 })
);
INV_X1 #() 
INV_X1_1456_ (
  .A({ S25434 }),
  .ZN({ S25492 })
);
NAND3_X1 #() 
NAND3_X1_4908_ (
  .A1({ S25421 }),
  .A2({ S25436 }),
  .A3({ S25422 }),
  .ZN({ S25493 })
);
AOI21_X1 #() 
AOI21_X1_2481_ (
  .A({ S89 }),
  .B1({ S25493 }),
  .B2({ S25485 }),
  .ZN({ S25494 })
);
AOI211_X1 #() 
AOI211_X1_80_ (
  .A({ S25416 }),
  .B({ S25494 }),
  .C1({ S25491 }),
  .C2({ S25492 }),
  .ZN({ S25495 })
);
OAI21_X1 #() 
OAI21_X1_2314_ (
  .A({ S25484 }),
  .B1({ S25490 }),
  .B2({ S25495 }),
  .ZN({ S25496 })
);
NAND2_X1 #() 
NAND2_X1_4496_ (
  .A1({ S25460 }),
  .A2({ S25957[906] }),
  .ZN({ S25497 })
);
NOR2_X1 #() 
NOR2_X1_1130_ (
  .A1({ S25456 }),
  .A2({ S25957[907] }),
  .ZN({ S25498 })
);
NAND2_X1 #() 
NAND2_X1_4497_ (
  .A1({ S25498 }),
  .A2({ S25497 }),
  .ZN({ S25499 })
);
NAND3_X1 #() 
NAND3_X1_4909_ (
  .A1({ S25437 }),
  .A2({ S25957[907] }),
  .A3({ S25429 }),
  .ZN({ S25500 })
);
NOR2_X1 #() 
NOR2_X1_1131_ (
  .A1({ S25436 }),
  .A2({ S89 }),
  .ZN({ S25501 })
);
AOI21_X1 #() 
AOI21_X1_2482_ (
  .A({ S25416 }),
  .B1({ S25501 }),
  .B2({ S25957[905] }),
  .ZN({ S25502 })
);
NAND3_X1 #() 
NAND3_X1_4910_ (
  .A1({ S25502 }),
  .A2({ S25499 }),
  .A3({ S25500 }),
  .ZN({ S25503 })
);
AND2_X1 #() 
AND2_X1_277_ (
  .A1({ S25422 }),
  .A2({ S25436 }),
  .ZN({ S25504 })
);
NAND3_X1 #() 
NAND3_X1_4911_ (
  .A1({ S25463 }),
  .A2({ S89 }),
  .A3({ S25429 }),
  .ZN({ S25505 })
);
OAI211_X1 #() 
OAI211_X1_1555_ (
  .A({ S25416 }),
  .B({ S25505 }),
  .C1({ S25504 }),
  .C2({ S25464 }),
  .ZN({ S25506 })
);
AND2_X1 #() 
AND2_X1_278_ (
  .A1({ S25503 }),
  .A2({ S25506 }),
  .ZN({ S25507 })
);
AOI21_X1 #() 
AOI21_X1_2483_ (
  .A({ S23551 }),
  .B1({ S25507 }),
  .B2({ S25957[909] }),
  .ZN({ S25508 })
);
NAND2_X1 #() 
NAND2_X1_4498_ (
  .A1({ S25437 }),
  .A2({ S25436 }),
  .ZN({ S25509 })
);
AOI22_X1 #() 
AOI22_X1_517_ (
  .A1({ S25509 }),
  .A2({ S25478 }),
  .B1({ S25475 }),
  .B2({ S25422 }),
  .ZN({ S25510 })
);
NAND2_X1 #() 
NAND2_X1_4499_ (
  .A1({ S25442 }),
  .A2({ S25957[907] }),
  .ZN({ S25511 })
);
NAND2_X1 #() 
NAND2_X1_4500_ (
  .A1({ S89 }),
  .A2({ S25957[904] }),
  .ZN({ S25512 })
);
OAI211_X1 #() 
OAI211_X1_1556_ (
  .A({ S25957[908] }),
  .B({ S25512 }),
  .C1({ S25425 }),
  .C2({ S25511 }),
  .ZN({ S25513 })
);
OAI211_X1 #() 
OAI211_X1_1557_ (
  .A({ S25957[909] }),
  .B({ S25513 }),
  .C1({ S25510 }),
  .C2({ S25957[908] }),
  .ZN({ S25514 })
);
NAND2_X1 #() 
NAND2_X1_4501_ (
  .A1({ S96 }),
  .A2({ S25436 }),
  .ZN({ S25515 })
);
NAND3_X1 #() 
NAND3_X1_4912_ (
  .A1({ S25491 }),
  .A2({ S89 }),
  .A3({ S25515 }),
  .ZN({ S25516 })
);
AOI21_X1 #() 
AOI21_X1_2484_ (
  .A({ S25416 }),
  .B1({ S25497 }),
  .B2({ S25957[907] }),
  .ZN({ S25517 })
);
NAND4_X1 #() 
NAND4_X1_527_ (
  .A1({ S25421 }),
  .A2({ S25422 }),
  .A3({ S89 }),
  .A4({ S25957[906] }),
  .ZN({ S25518 })
);
AOI21_X1 #() 
AOI21_X1_2485_ (
  .A({ S25957[908] }),
  .B1({ S25501 }),
  .B2({ S25437 }),
  .ZN({ S25519 })
);
AOI22_X1 #() 
AOI22_X1_518_ (
  .A1({ S25516 }),
  .A2({ S25517 }),
  .B1({ S25519 }),
  .B2({ S25518 }),
  .ZN({ S25520 })
);
AOI21_X1 #() 
AOI21_X1_2486_ (
  .A({ S25957[910] }),
  .B1({ S25520 }),
  .B2({ S25484 }),
  .ZN({ S25521 })
);
AOI22_X1 #() 
AOI22_X1_519_ (
  .A1({ S25496 }),
  .A2({ S25508 }),
  .B1({ S25521 }),
  .B2({ S25514 }),
  .ZN({ S25522 })
);
NOR2_X1 #() 
NOR2_X1_1132_ (
  .A1({ S25522 }),
  .A2({ S25957[911] }),
  .ZN({ S25523 })
);
NOR3_X1 #() 
NOR3_X1_151_ (
  .A1({ S25523 }),
  .A2({ S25483 }),
  .A3({ S20239 }),
  .ZN({ S25524 })
);
NOR2_X1 #() 
NOR2_X1_1133_ (
  .A1({ S25523 }),
  .A2({ S25483 }),
  .ZN({ S25525 })
);
NOR2_X1 #() 
NOR2_X1_1134_ (
  .A1({ S25525 }),
  .A2({ S25957[1111] }),
  .ZN({ S25526 })
);
NOR2_X1 #() 
NOR2_X1_1135_ (
  .A1({ S25526 }),
  .A2({ S25524 }),
  .ZN({ S25957[855] })
);
INV_X1 #() 
INV_X1_1457_ (
  .A({ S25957[855] }),
  .ZN({ S25527 })
);
NAND2_X1 #() 
NAND2_X1_4502_ (
  .A1({ S25527 }),
  .A2({ S25957[1047] }),
  .ZN({ S25528 })
);
NAND2_X1 #() 
NAND2_X1_4503_ (
  .A1({ S25957[855] }),
  .A2({ S20242 }),
  .ZN({ S25529 })
);
NAND2_X1 #() 
NAND2_X1_4504_ (
  .A1({ S25528 }),
  .A2({ S25529 }),
  .ZN({ S25957[791] })
);
AOI21_X1 #() 
AOI21_X1_2487_ (
  .A({ S25957[906] }),
  .B1({ S25437 }),
  .B2({ S97 }),
  .ZN({ S25530 })
);
NAND2_X1 #() 
NAND2_X1_4505_ (
  .A1({ S25469 }),
  .A2({ S97 }),
  .ZN({ S25531 })
);
OAI22_X1 #() 
OAI22_X1_116_ (
  .A1({ S25530 }),
  .A2({ S25430 }),
  .B1({ S25531 }),
  .B2({ S25511 }),
  .ZN({ S25532 })
);
OAI211_X1 #() 
OAI211_X1_1558_ (
  .A({ S25445 }),
  .B({ S25446 }),
  .C1({ S25486 }),
  .C2({ S25957[907] }),
  .ZN({ S25533 })
);
AOI21_X1 #() 
AOI21_X1_2488_ (
  .A({ S25957[909] }),
  .B1({ S25533 }),
  .B2({ S25957[908] }),
  .ZN({ S25534 })
);
OAI21_X1 #() 
OAI21_X1_2315_ (
  .A({ S25534 }),
  .B1({ S25957[908] }),
  .B2({ S25532 }),
  .ZN({ S25535 })
);
NAND3_X1 #() 
NAND3_X1_4913_ (
  .A1({ S25436 }),
  .A2({ S23922 }),
  .A3({ S23925 }),
  .ZN({ S25536 })
);
NAND2_X1 #() 
NAND2_X1_4506_ (
  .A1({ S25536 }),
  .A2({ S25957[907] }),
  .ZN({ S25537 })
);
AOI22_X1 #() 
AOI22_X1_520_ (
  .A1({ S25436 }),
  .A2({ S25408 }),
  .B1({ S23922 }),
  .B2({ S23925 }),
  .ZN({ S25538 })
);
NAND2_X1 #() 
NAND2_X1_4507_ (
  .A1({ S97 }),
  .A2({ S25436 }),
  .ZN({ S25539 })
);
NAND2_X1 #() 
NAND2_X1_4508_ (
  .A1({ S25491 }),
  .A2({ S25539 }),
  .ZN({ S25540 })
);
AOI21_X1 #() 
AOI21_X1_2489_ (
  .A({ S25957[908] }),
  .B1({ S25540 }),
  .B2({ S89 }),
  .ZN({ S25541 })
);
OAI21_X1 #() 
OAI21_X1_2316_ (
  .A({ S25541 }),
  .B1({ S25537 }),
  .B2({ S25538 }),
  .ZN({ S25542 })
);
NAND2_X1 #() 
NAND2_X1_4509_ (
  .A1({ S25443 }),
  .A2({ S25456 }),
  .ZN({ S25543 })
);
NAND3_X1 #() 
NAND3_X1_4914_ (
  .A1({ S25502 }),
  .A2({ S25518 }),
  .A3({ S25543 }),
  .ZN({ S25544 })
);
NAND3_X1 #() 
NAND3_X1_4915_ (
  .A1({ S25542 }),
  .A2({ S25957[909] }),
  .A3({ S25544 }),
  .ZN({ S25545 })
);
AOI21_X1 #() 
AOI21_X1_2490_ (
  .A({ S25957[910] }),
  .B1({ S25545 }),
  .B2({ S25535 }),
  .ZN({ S25546 })
);
AOI21_X1 #() 
AOI21_X1_2491_ (
  .A({ S25957[904] }),
  .B1({ S24010 }),
  .B2({ S24013 }),
  .ZN({ S25547 })
);
NOR2_X1 #() 
NOR2_X1_1136_ (
  .A1({ S25547 }),
  .A2({ S25957[907] }),
  .ZN({ S25548 })
);
NAND2_X1 #() 
NAND2_X1_4510_ (
  .A1({ S25422 }),
  .A2({ S25957[906] }),
  .ZN({ S25549 })
);
NAND2_X1 #() 
NAND2_X1_4511_ (
  .A1({ S25549 }),
  .A2({ S25433 }),
  .ZN({ S25550 })
);
NAND2_X1 #() 
NAND2_X1_4512_ (
  .A1({ S25550 }),
  .A2({ S25957[907] }),
  .ZN({ S25551 })
);
INV_X1 #() 
INV_X1_1458_ (
  .A({ S25551 }),
  .ZN({ S25552 })
);
AOI21_X1 #() 
AOI21_X1_2492_ (
  .A({ S25552 }),
  .B1({ S25548 }),
  .B2({ S25493 }),
  .ZN({ S25553 })
);
INV_X1 #() 
INV_X1_1459_ (
  .A({ S25442 }),
  .ZN({ S25554 })
);
NAND4_X1 #() 
NAND4_X1_528_ (
  .A1({ S25486 }),
  .A2({ S25463 }),
  .A3({ S25429 }),
  .A4({ S89 }),
  .ZN({ S25555 })
);
NAND2_X1 #() 
NAND2_X1_4513_ (
  .A1({ S25469 }),
  .A2({ S25957[905] }),
  .ZN({ S25556 })
);
NAND2_X1 #() 
NAND2_X1_4514_ (
  .A1({ S25556 }),
  .A2({ S25957[907] }),
  .ZN({ S25557 })
);
OAI211_X1 #() 
OAI211_X1_1559_ (
  .A({ S25555 }),
  .B({ S25416 }),
  .C1({ S25557 }),
  .C2({ S25554 }),
  .ZN({ S25558 })
);
OAI211_X1 #() 
OAI211_X1_1560_ (
  .A({ S25558 }),
  .B({ S25484 }),
  .C1({ S25553 }),
  .C2({ S25416 }),
  .ZN({ S25559 })
);
NAND3_X1 #() 
NAND3_X1_4916_ (
  .A1({ S25454 }),
  .A2({ S25433 }),
  .A3({ S25429 }),
  .ZN({ S25560 })
);
OAI211_X1 #() 
OAI211_X1_1561_ (
  .A({ S25560 }),
  .B({ S25957[908] }),
  .C1({ S25957[907] }),
  .C2({ S25455 }),
  .ZN({ S25561 })
);
INV_X1 #() 
INV_X1_1460_ (
  .A({ S25443 }),
  .ZN({ S25562 })
);
NAND2_X1 #() 
NAND2_X1_4515_ (
  .A1({ S25466 }),
  .A2({ S25562 }),
  .ZN({ S25563 })
);
AOI21_X1 #() 
AOI21_X1_2493_ (
  .A({ S25484 }),
  .B1({ S25563 }),
  .B2({ S25416 }),
  .ZN({ S25564 })
);
AOI21_X1 #() 
AOI21_X1_2494_ (
  .A({ S23551 }),
  .B1({ S25564 }),
  .B2({ S25561 }),
  .ZN({ S25565 })
);
AND2_X1 #() 
AND2_X1_279_ (
  .A1({ S25559 }),
  .A2({ S25565 }),
  .ZN({ S25566 })
);
OAI21_X1 #() 
OAI21_X1_2317_ (
  .A({ S25957[911] }),
  .B1({ S25566 }),
  .B2({ S25546 }),
  .ZN({ S25567 })
);
AND2_X1 #() 
AND2_X1_280_ (
  .A1({ S23481 }),
  .A2({ S23480 }),
  .ZN({ S25568 })
);
AOI21_X1 #() 
AOI21_X1_2495_ (
  .A({ S25957[907] }),
  .B1({ S25421 }),
  .B2({ S25429 }),
  .ZN({ S25569 })
);
NAND2_X1 #() 
NAND2_X1_4516_ (
  .A1({ S25436 }),
  .A2({ S25957[905] }),
  .ZN({ S25570 })
);
OAI21_X1 #() 
OAI21_X1_2318_ (
  .A({ S25957[908] }),
  .B1({ S25570 }),
  .B2({ S89 }),
  .ZN({ S25571 })
);
NOR2_X1 #() 
NOR2_X1_1137_ (
  .A1({ S25571 }),
  .A2({ S25569 }),
  .ZN({ S25572 })
);
NAND4_X1 #() 
NAND4_X1_529_ (
  .A1({ S25463 }),
  .A2({ S25429 }),
  .A3({ S25433 }),
  .A4({ S89 }),
  .ZN({ S25573 })
);
NAND2_X1 #() 
NAND2_X1_4517_ (
  .A1({ S25421 }),
  .A2({ S25442 }),
  .ZN({ S25574 })
);
AOI21_X1 #() 
AOI21_X1_2496_ (
  .A({ S25416 }),
  .B1({ S25574 }),
  .B2({ S25957[907] }),
  .ZN({ S25575 })
);
NAND2_X1 #() 
NAND2_X1_4518_ (
  .A1({ S25433 }),
  .A2({ S25957[905] }),
  .ZN({ S25576 })
);
AOI21_X1 #() 
AOI21_X1_2497_ (
  .A({ S25957[908] }),
  .B1({ S25446 }),
  .B2({ S25576 }),
  .ZN({ S25577 })
);
AOI21_X1 #() 
AOI21_X1_2498_ (
  .A({ S25577 }),
  .B1({ S25575 }),
  .B2({ S25573 }),
  .ZN({ S25578 })
);
NOR2_X1 #() 
NOR2_X1_1138_ (
  .A1({ S25455 }),
  .A2({ S96 }),
  .ZN({ S25579 })
);
OAI211_X1 #() 
OAI211_X1_1562_ (
  .A({ S25551 }),
  .B({ S25416 }),
  .C1({ S25957[907] }),
  .C2({ S25579 }),
  .ZN({ S25580 })
);
NAND2_X1 #() 
NAND2_X1_4519_ (
  .A1({ S25580 }),
  .A2({ S25484 }),
  .ZN({ S25581 })
);
OAI221_X1 #() 
OAI221_X1_130_ (
  .A({ S25957[910] }),
  .B1({ S25578 }),
  .B2({ S25484 }),
  .C1({ S25581 }),
  .C2({ S25572 }),
  .ZN({ S25582 })
);
NAND3_X1 #() 
NAND3_X1_4917_ (
  .A1({ S25444 }),
  .A2({ S25957[904] }),
  .A3({ S25436 }),
  .ZN({ S25583 })
);
NAND3_X1 #() 
NAND3_X1_4918_ (
  .A1({ S25583 }),
  .A2({ S25957[907] }),
  .A3({ S25417 }),
  .ZN({ S25584 })
);
OAI21_X1 #() 
OAI21_X1_2319_ (
  .A({ S25584 }),
  .B1({ S25957[907] }),
  .B2({ S25583 }),
  .ZN({ S25585 })
);
NOR2_X1 #() 
NOR2_X1_1139_ (
  .A1({ S25421 }),
  .A2({ S25436 }),
  .ZN({ S25586 })
);
NOR2_X1 #() 
NOR2_X1_1140_ (
  .A1({ S25460 }),
  .A2({ S25957[906] }),
  .ZN({ S25587 })
);
OAI211_X1 #() 
OAI211_X1_1563_ (
  .A({ S25957[907] }),
  .B({ S25416 }),
  .C1({ S25586 }),
  .C2({ S25587 }),
  .ZN({ S25588 })
);
INV_X1 #() 
INV_X1_1461_ (
  .A({ S25588 }),
  .ZN({ S25589 })
);
AOI21_X1 #() 
AOI21_X1_2499_ (
  .A({ S25589 }),
  .B1({ S25585 }),
  .B2({ S25957[908] }),
  .ZN({ S25590 })
);
INV_X1 #() 
INV_X1_1462_ (
  .A({ S25570 }),
  .ZN({ S25591 })
);
NOR2_X1 #() 
NOR2_X1_1141_ (
  .A1({ S25422 }),
  .A2({ S25957[906] }),
  .ZN({ S25592 })
);
INV_X1 #() 
INV_X1_1463_ (
  .A({ S25478 }),
  .ZN({ S25593 })
);
OAI22_X1 #() 
OAI22_X1_117_ (
  .A1({ S25593 }),
  .A2({ S25592 }),
  .B1({ S25591 }),
  .B2({ S25464 }),
  .ZN({ S25594 })
);
AOI21_X1 #() 
AOI21_X1_2500_ (
  .A({ S25416 }),
  .B1({ S25433 }),
  .B2({ S89 }),
  .ZN({ S25595 })
);
INV_X1 #() 
INV_X1_1464_ (
  .A({ S25509 }),
  .ZN({ S25596 })
);
OAI21_X1 #() 
OAI21_X1_2320_ (
  .A({ S25957[907] }),
  .B1({ S25596 }),
  .B2({ S25579 }),
  .ZN({ S25597 })
);
AOI21_X1 #() 
AOI21_X1_2501_ (
  .A({ S25484 }),
  .B1({ S25597 }),
  .B2({ S25595 }),
  .ZN({ S25598 })
);
OAI21_X1 #() 
OAI21_X1_2321_ (
  .A({ S25598 }),
  .B1({ S25957[908] }),
  .B2({ S25594 }),
  .ZN({ S25599 })
);
OAI211_X1 #() 
OAI211_X1_1564_ (
  .A({ S25599 }),
  .B({ S23551 }),
  .C1({ S25957[909] }),
  .C2({ S25590 }),
  .ZN({ S25600 })
);
NAND3_X1 #() 
NAND3_X1_4919_ (
  .A1({ S25600 }),
  .A2({ S25568 }),
  .A3({ S25582 }),
  .ZN({ S25601 })
);
NAND2_X1 #() 
NAND2_X1_4520_ (
  .A1({ S25567 }),
  .A2({ S25601 }),
  .ZN({ S25602 })
);
OR2_X1 #() 
OR2_X1_62_ (
  .A1({ S25602 }),
  .A2({ S25957[1110] }),
  .ZN({ S25603 })
);
NAND2_X1 #() 
NAND2_X1_4521_ (
  .A1({ S25602 }),
  .A2({ S25957[1110] }),
  .ZN({ S25604 })
);
AOI21_X1 #() 
AOI21_X1_2502_ (
  .A({ S25957[1046] }),
  .B1({ S25603 }),
  .B2({ S25604 }),
  .ZN({ S25605 })
);
NAND2_X1 #() 
NAND2_X1_4522_ (
  .A1({ S25603 }),
  .A2({ S25604 }),
  .ZN({ S25957[854] })
);
NOR2_X1 #() 
NOR2_X1_1142_ (
  .A1({ S25957[854] }),
  .A2({ S22832 }),
  .ZN({ S25606 })
);
NOR2_X1 #() 
NOR2_X1_1143_ (
  .A1({ S25606 }),
  .A2({ S25605 }),
  .ZN({ S25607 })
);
INV_X1 #() 
INV_X1_1465_ (
  .A({ S25607 }),
  .ZN({ S25957[790] })
);
NAND2_X1 #() 
NAND2_X1_4523_ (
  .A1({ S22920 }),
  .A2({ S22924 }),
  .ZN({ S25608 })
);
NAND2_X1 #() 
NAND2_X1_4524_ (
  .A1({ S20387 }),
  .A2({ S20388 }),
  .ZN({ S25957[1141] })
);
NAND2_X1 #() 
NAND2_X1_4525_ (
  .A1({ S22909 }),
  .A2({ S22875 }),
  .ZN({ S25609 })
);
XNOR2_X1 #() 
XNOR2_X1_179_ (
  .A({ S25609 }),
  .B({ S25957[1141] }),
  .ZN({ S25957[1013] })
);
NAND2_X1 #() 
NAND2_X1_4526_ (
  .A1({ S25460 }),
  .A2({ S25436 }),
  .ZN({ S25610 })
);
NAND3_X1 #() 
NAND3_X1_4920_ (
  .A1({ S25435 }),
  .A2({ S25957[907] }),
  .A3({ S25610 }),
  .ZN({ S25611 })
);
NAND2_X1 #() 
NAND2_X1_4527_ (
  .A1({ S25957[907] }),
  .A2({ S25408 }),
  .ZN({ S25612 })
);
NAND2_X1 #() 
NAND2_X1_4528_ (
  .A1({ S25461 }),
  .A2({ S25433 }),
  .ZN({ S25613 })
);
AOI21_X1 #() 
AOI21_X1_2503_ (
  .A({ S25957[908] }),
  .B1({ S25613 }),
  .B2({ S25612 }),
  .ZN({ S25614 })
);
NAND3_X1 #() 
NAND3_X1_4921_ (
  .A1({ S25486 }),
  .A2({ S89 }),
  .A3({ S25463 }),
  .ZN({ S25615 })
);
AND2_X1 #() 
AND2_X1_281_ (
  .A1({ S25615 }),
  .A2({ S25957[908] }),
  .ZN({ S25616 })
);
AOI211_X1 #() 
AOI211_X1_81_ (
  .A({ S25484 }),
  .B({ S25614 }),
  .C1({ S25611 }),
  .C2({ S25616 }),
  .ZN({ S25617 })
);
NAND2_X1 #() 
NAND2_X1_4529_ (
  .A1({ S25610 }),
  .A2({ S89 }),
  .ZN({ S25618 })
);
NAND4_X1 #() 
NAND4_X1_530_ (
  .A1({ S25463 }),
  .A2({ S25429 }),
  .A3({ S25433 }),
  .A4({ S25957[907] }),
  .ZN({ S25619 })
);
AOI21_X1 #() 
AOI21_X1_2504_ (
  .A({ S25957[908] }),
  .B1({ S25618 }),
  .B2({ S25619 }),
  .ZN({ S25620 })
);
INV_X1 #() 
INV_X1_1466_ (
  .A({ S25620 }),
  .ZN({ S25621 })
);
NAND3_X1 #() 
NAND3_X1_4922_ (
  .A1({ S25433 }),
  .A2({ S25957[907] }),
  .A3({ S25957[905] }),
  .ZN({ S25622 })
);
AOI21_X1 #() 
AOI21_X1_2505_ (
  .A({ S25621 }),
  .B1({ S25554 }),
  .B2({ S25622 }),
  .ZN({ S25623 })
);
AOI21_X1 #() 
AOI21_X1_2506_ (
  .A({ S25957[907] }),
  .B1({ S25485 }),
  .B2({ S25515 }),
  .ZN({ S25624 })
);
OAI21_X1 #() 
OAI21_X1_2322_ (
  .A({ S25484 }),
  .B1({ S25624 }),
  .B2({ S25472 }),
  .ZN({ S25625 })
);
OAI21_X1 #() 
OAI21_X1_2323_ (
  .A({ S25957[910] }),
  .B1({ S25623 }),
  .B2({ S25625 }),
  .ZN({ S25626 })
);
OAI21_X1 #() 
OAI21_X1_2324_ (
  .A({ S25577 }),
  .B1({ S25470 }),
  .B2({ S25548 }),
  .ZN({ S25627 })
);
OAI211_X1 #() 
OAI211_X1_1565_ (
  .A({ S25957[908] }),
  .B({ S25543 }),
  .C1({ S25596 }),
  .C2({ S89 }),
  .ZN({ S25628 })
);
NAND3_X1 #() 
NAND3_X1_4923_ (
  .A1({ S25627 }),
  .A2({ S25628 }),
  .A3({ S25957[909] }),
  .ZN({ S25629 })
);
NAND3_X1 #() 
NAND3_X1_4924_ (
  .A1({ S25435 }),
  .A2({ S25957[907] }),
  .A3({ S25583 }),
  .ZN({ S25630 })
);
NAND2_X1 #() 
NAND2_X1_4530_ (
  .A1({ S25477 }),
  .A2({ S25461 }),
  .ZN({ S25631 })
);
NAND3_X1 #() 
NAND3_X1_4925_ (
  .A1({ S25630 }),
  .A2({ S25957[908] }),
  .A3({ S25631 }),
  .ZN({ S25632 })
);
NOR2_X1 #() 
NOR2_X1_1144_ (
  .A1({ S25478 }),
  .A2({ S25957[908] }),
  .ZN({ S25633 })
);
OAI211_X1 #() 
OAI211_X1_1566_ (
  .A({ S25633 }),
  .B({ S25957[904] }),
  .C1({ S25454 }),
  .C2({ S89 }),
  .ZN({ S25634 })
);
NAND3_X1 #() 
NAND3_X1_4926_ (
  .A1({ S25634 }),
  .A2({ S25632 }),
  .A3({ S25484 }),
  .ZN({ S25635 })
);
NAND3_X1 #() 
NAND3_X1_4927_ (
  .A1({ S25635 }),
  .A2({ S23551 }),
  .A3({ S25629 }),
  .ZN({ S25636 })
);
OAI211_X1 #() 
OAI211_X1_1567_ (
  .A({ S25568 }),
  .B({ S25636 }),
  .C1({ S25626 }),
  .C2({ S25617 }),
  .ZN({ S25637 })
);
AOI211_X1 #() 
AOI211_X1_82_ (
  .A({ S25443 }),
  .B({ S25554 }),
  .C1({ S25556 }),
  .C2({ S25957[907] }),
  .ZN({ S25638 })
);
OAI221_X1 #() 
OAI221_X1_131_ (
  .A({ S25957[908] }),
  .B1({ S25537 }),
  .B2({ S25957[904] }),
  .C1({ S25504 }),
  .C2({ S25462 }),
  .ZN({ S25639 })
);
OAI21_X1 #() 
OAI21_X1_2325_ (
  .A({ S25639 }),
  .B1({ S25638 }),
  .B2({ S25957[908] }),
  .ZN({ S25640 })
);
AOI21_X1 #() 
AOI21_X1_2507_ (
  .A({ S25957[908] }),
  .B1({ S25551 }),
  .B2({ S25518 }),
  .ZN({ S25641 })
);
NAND2_X1 #() 
NAND2_X1_4531_ (
  .A1({ S25421 }),
  .A2({ S25957[906] }),
  .ZN({ S25642 })
);
NAND2_X1 #() 
NAND2_X1_4532_ (
  .A1({ S25460 }),
  .A2({ S25957[907] }),
  .ZN({ S25643 })
);
AOI21_X1 #() 
AOI21_X1_2508_ (
  .A({ S25416 }),
  .B1({ S25642 }),
  .B2({ S25643 }),
  .ZN({ S25644 })
);
OR3_X1 #() 
OR3_X1_29_ (
  .A1({ S25641 }),
  .A2({ S25644 }),
  .A3({ S25957[909] }),
  .ZN({ S25645 })
);
OAI211_X1 #() 
OAI211_X1_1568_ (
  .A({ S25645 }),
  .B({ S25957[910] }),
  .C1({ S25640 }),
  .C2({ S25484 }),
  .ZN({ S25646 })
);
NAND2_X1 #() 
NAND2_X1_4533_ (
  .A1({ S25429 }),
  .A2({ S25422 }),
  .ZN({ S25647 })
);
OAI221_X1 #() 
OAI221_X1_132_ (
  .A({ S25957[908] }),
  .B1({ S25501 }),
  .B2({ S25647 }),
  .C1({ S89 }),
  .C2({ S25485 }),
  .ZN({ S25648 })
);
OAI21_X1 #() 
OAI21_X1_2326_ (
  .A({ S25445 }),
  .B1({ S25462 }),
  .B2({ S25425 }),
  .ZN({ S25649 })
);
NAND2_X1 #() 
NAND2_X1_4534_ (
  .A1({ S25649 }),
  .A2({ S25416 }),
  .ZN({ S25650 })
);
AOI21_X1 #() 
AOI21_X1_2509_ (
  .A({ S25484 }),
  .B1({ S25650 }),
  .B2({ S25648 }),
  .ZN({ S25651 })
);
INV_X1 #() 
INV_X1_1467_ (
  .A({ S25515 }),
  .ZN({ S25652 })
);
NOR2_X1 #() 
NOR2_X1_1145_ (
  .A1({ S25652 }),
  .A2({ S25957[907] }),
  .ZN({ S25653 })
);
AOI21_X1 #() 
AOI21_X1_2510_ (
  .A({ S89 }),
  .B1({ S25491 }),
  .B2({ S25457 }),
  .ZN({ S25654 })
);
OAI21_X1 #() 
OAI21_X1_2327_ (
  .A({ S25416 }),
  .B1({ S25653 }),
  .B2({ S25654 }),
  .ZN({ S25655 })
);
NAND2_X1 #() 
NAND2_X1_4535_ (
  .A1({ S25423 }),
  .A2({ S25957[907] }),
  .ZN({ S25656 })
);
NOR2_X1 #() 
NOR2_X1_1146_ (
  .A1({ S25416 }),
  .A2({ S25444 }),
  .ZN({ S25657 })
);
OAI21_X1 #() 
OAI21_X1_2328_ (
  .A({ S25656 }),
  .B1({ S25595 }),
  .B2({ S25657 }),
  .ZN({ S25658 })
);
AOI21_X1 #() 
AOI21_X1_2511_ (
  .A({ S25957[909] }),
  .B1({ S25655 }),
  .B2({ S25658 }),
  .ZN({ S25659 })
);
OAI21_X1 #() 
OAI21_X1_2329_ (
  .A({ S23551 }),
  .B1({ S25659 }),
  .B2({ S25651 }),
  .ZN({ S25660 })
);
NAND3_X1 #() 
NAND3_X1_4928_ (
  .A1({ S25646 }),
  .A2({ S25957[911] }),
  .A3({ S25660 }),
  .ZN({ S25661 })
);
NAND2_X1 #() 
NAND2_X1_4536_ (
  .A1({ S25661 }),
  .A2({ S25637 }),
  .ZN({ S25662 })
);
NAND2_X1 #() 
NAND2_X1_4537_ (
  .A1({ S25662 }),
  .A2({ S25957[1013] }),
  .ZN({ S25663 })
);
INV_X1 #() 
INV_X1_1468_ (
  .A({ S25957[1013] }),
  .ZN({ S25664 })
);
NAND3_X1 #() 
NAND3_X1_4929_ (
  .A1({ S25661 }),
  .A2({ S25637 }),
  .A3({ S25664 }),
  .ZN({ S25665 })
);
NAND2_X1 #() 
NAND2_X1_4538_ (
  .A1({ S25663 }),
  .A2({ S25665 }),
  .ZN({ S25666 })
);
NOR2_X1 #() 
NOR2_X1_1147_ (
  .A1({ S25666 }),
  .A2({ S22838 }),
  .ZN({ S25667 })
);
AOI21_X1 #() 
AOI21_X1_2512_ (
  .A({ S25957[1077] }),
  .B1({ S25663 }),
  .B2({ S25665 }),
  .ZN({ S25668 })
);
OAI21_X1 #() 
OAI21_X1_2330_ (
  .A({ S25608 }),
  .B1({ S25667 }),
  .B2({ S25668 }),
  .ZN({ S25669 })
);
INV_X1 #() 
INV_X1_1469_ (
  .A({ S25666 }),
  .ZN({ S25957[885] })
);
NAND2_X1 #() 
NAND2_X1_4539_ (
  .A1({ S25957[885] }),
  .A2({ S25957[1077] }),
  .ZN({ S25670 })
);
INV_X1 #() 
INV_X1_1470_ (
  .A({ S25668 }),
  .ZN({ S25671 })
);
NAND3_X1 #() 
NAND3_X1_4930_ (
  .A1({ S25670 }),
  .A2({ S25957[917] }),
  .A3({ S25671 }),
  .ZN({ S25672 })
);
NAND2_X1 #() 
NAND2_X1_4540_ (
  .A1({ S25672 }),
  .A2({ S25669 }),
  .ZN({ S25673 })
);
INV_X1 #() 
INV_X1_1471_ (
  .A({ S25673 }),
  .ZN({ S25957[789] })
);
INV_X1 #() 
INV_X1_1472_ (
  .A({ S22980 }),
  .ZN({ S25674 })
);
INV_X1 #() 
INV_X1_1473_ (
  .A({ S22982 }),
  .ZN({ S25675 })
);
NOR2_X1 #() 
NOR2_X1_1148_ (
  .A1({ S25675 }),
  .A2({ S25674 }),
  .ZN({ S25957[980] })
);
XNOR2_X1 #() 
XNOR2_X1_180_ (
  .A({ S25957[980] }),
  .B({ S25957[1076] }),
  .ZN({ S25676 })
);
INV_X1 #() 
INV_X1_1474_ (
  .A({ S25676 }),
  .ZN({ S25957[948] })
);
NAND2_X1 #() 
NAND2_X1_4541_ (
  .A1({ S20460 }),
  .A2({ S20449 }),
  .ZN({ S25957[1140] })
);
NAND2_X1 #() 
NAND2_X1_4542_ (
  .A1({ S22981 }),
  .A2({ S22954 }),
  .ZN({ S25677 })
);
XNOR2_X1 #() 
XNOR2_X1_181_ (
  .A({ S25677 }),
  .B({ S25957[1140] }),
  .ZN({ S25957[1012] })
);
INV_X1 #() 
INV_X1_1475_ (
  .A({ S25957[1012] }),
  .ZN({ S25678 })
);
INV_X1 #() 
INV_X1_1476_ (
  .A({ S25422 }),
  .ZN({ S25679 })
);
NAND2_X1 #() 
NAND2_X1_4543_ (
  .A1({ S25610 }),
  .A2({ S25957[907] }),
  .ZN({ S25680 })
);
INV_X1 #() 
INV_X1_1477_ (
  .A({ S25549 }),
  .ZN({ S25681 })
);
OAI21_X1 #() 
OAI21_X1_2331_ (
  .A({ S89 }),
  .B1({ S25681 }),
  .B2({ S25587 }),
  .ZN({ S25682 })
);
OAI211_X1 #() 
OAI211_X1_1569_ (
  .A({ S25682 }),
  .B({ S25957[908] }),
  .C1({ S25679 }),
  .C2({ S25680 }),
  .ZN({ S25683 })
);
NAND2_X1 #() 
NAND2_X1_4544_ (
  .A1({ S25463 }),
  .A2({ S25429 }),
  .ZN({ S25684 })
);
OAI21_X1 #() 
OAI21_X1_2332_ (
  .A({ S89 }),
  .B1({ S25530 }),
  .B2({ S25684 }),
  .ZN({ S25685 })
);
NAND4_X1 #() 
NAND4_X1_531_ (
  .A1({ S25685 }),
  .A2({ S25643 }),
  .A3({ S25471 }),
  .A4({ S25416 }),
  .ZN({ S25686 })
);
NAND3_X1 #() 
NAND3_X1_4931_ (
  .A1({ S25686 }),
  .A2({ S25683 }),
  .A3({ S25957[909] }),
  .ZN({ S25687 })
);
NAND3_X1 #() 
NAND3_X1_4932_ (
  .A1({ S25444 }),
  .A2({ S25442 }),
  .A3({ S25957[907] }),
  .ZN({ S25688 })
);
NAND2_X1 #() 
NAND2_X1_4545_ (
  .A1({ S25421 }),
  .A2({ S25436 }),
  .ZN({ S25689 })
);
AOI21_X1 #() 
AOI21_X1_2513_ (
  .A({ S25957[907] }),
  .B1({ S25689 }),
  .B2({ S25497 }),
  .ZN({ S25690 })
);
NOR2_X1 #() 
NOR2_X1_1149_ (
  .A1({ S25690 }),
  .A2({ S25957[908] }),
  .ZN({ S25691 })
);
NAND2_X1 #() 
NAND2_X1_4546_ (
  .A1({ S25691 }),
  .A2({ S25688 }),
  .ZN({ S25692 })
);
OAI21_X1 #() 
OAI21_X1_2333_ (
  .A({ S89 }),
  .B1({ S25556 }),
  .B2({ S25554 }),
  .ZN({ S25693 })
);
AOI21_X1 #() 
AOI21_X1_2514_ (
  .A({ S89 }),
  .B1({ S25957[904] }),
  .B2({ S25957[906] }),
  .ZN({ S25694 })
);
NAND3_X1 #() 
NAND3_X1_4933_ (
  .A1({ S25694 }),
  .A2({ S25463 }),
  .A3({ S25570 }),
  .ZN({ S25695 })
);
NAND3_X1 #() 
NAND3_X1_4934_ (
  .A1({ S25695 }),
  .A2({ S25693 }),
  .A3({ S25957[908] }),
  .ZN({ S25696 })
);
NAND3_X1 #() 
NAND3_X1_4935_ (
  .A1({ S25692 }),
  .A2({ S25484 }),
  .A3({ S25696 }),
  .ZN({ S25697 })
);
NAND3_X1 #() 
NAND3_X1_4936_ (
  .A1({ S25697 }),
  .A2({ S25687 }),
  .A3({ S23551 }),
  .ZN({ S25698 })
);
OAI21_X1 #() 
OAI21_X1_2334_ (
  .A({ S89 }),
  .B1({ S97 }),
  .B2({ S25436 }),
  .ZN({ S25699 })
);
NAND3_X1 #() 
NAND3_X1_4937_ (
  .A1({ S25699 }),
  .A2({ S25957[908] }),
  .A3({ S25471 }),
  .ZN({ S25700 })
);
NAND3_X1 #() 
NAND3_X1_4938_ (
  .A1({ S25570 }),
  .A2({ S89 }),
  .A3({ S25408 }),
  .ZN({ S25701 })
);
OAI21_X1 #() 
OAI21_X1_2335_ (
  .A({ S25701 }),
  .B1({ S25511 }),
  .B2({ S25425 }),
  .ZN({ S25702 })
);
OAI211_X1 #() 
OAI211_X1_1570_ (
  .A({ S25957[909] }),
  .B({ S25700 }),
  .C1({ S25702 }),
  .C2({ S25957[908] }),
  .ZN({ S25703 })
);
NAND2_X1 #() 
NAND2_X1_4547_ (
  .A1({ S25433 }),
  .A2({ S25957[907] }),
  .ZN({ S25704 })
);
OAI221_X1 #() 
OAI221_X1_133_ (
  .A({ S25957[908] }),
  .B1({ S25704 }),
  .B2({ S25957[905] }),
  .C1({ S25462 }),
  .C2({ S25425 }),
  .ZN({ S25705 })
);
NAND2_X1 #() 
NAND2_X1_4548_ (
  .A1({ S25548 }),
  .A2({ S25536 }),
  .ZN({ S25706 })
);
AOI21_X1 #() 
AOI21_X1_2515_ (
  .A({ S25957[908] }),
  .B1({ S25475 }),
  .B2({ S25422 }),
  .ZN({ S25707 })
);
NAND2_X1 #() 
NAND2_X1_4549_ (
  .A1({ S25707 }),
  .A2({ S25706 }),
  .ZN({ S25708 })
);
NAND3_X1 #() 
NAND3_X1_4939_ (
  .A1({ S25705 }),
  .A2({ S25484 }),
  .A3({ S25708 }),
  .ZN({ S25709 })
);
NAND3_X1 #() 
NAND3_X1_4940_ (
  .A1({ S25709 }),
  .A2({ S25703 }),
  .A3({ S25957[910] }),
  .ZN({ S25710 })
);
NAND3_X1 #() 
NAND3_X1_4941_ (
  .A1({ S25698 }),
  .A2({ S25957[911] }),
  .A3({ S25710 }),
  .ZN({ S25711 })
);
INV_X1 #() 
INV_X1_1478_ (
  .A({ S25711 }),
  .ZN({ S25712 })
);
NOR2_X1 #() 
NOR2_X1_1150_ (
  .A1({ S25501 }),
  .A2({ S25957[908] }),
  .ZN({ S25713 })
);
OAI21_X1 #() 
OAI21_X1_2336_ (
  .A({ S25713 }),
  .B1({ S25652 }),
  .B2({ S25430 }),
  .ZN({ S25714 })
);
NAND2_X1 #() 
NAND2_X1_4550_ (
  .A1({ S25455 }),
  .A2({ S89 }),
  .ZN({ S25715 })
);
NOR2_X1 #() 
NOR2_X1_1151_ (
  .A1({ S25715 }),
  .A2({ S25425 }),
  .ZN({ S25716 })
);
OAI21_X1 #() 
OAI21_X1_2337_ (
  .A({ S25714 }),
  .B1({ S25447 }),
  .B2({ S25716 }),
  .ZN({ S25717 })
);
AOI21_X1 #() 
AOI21_X1_2516_ (
  .A({ S25416 }),
  .B1({ S128 }),
  .B2({ S25436 }),
  .ZN({ S25718 })
);
AOI21_X1 #() 
AOI21_X1_2517_ (
  .A({ S25957[907] }),
  .B1({ S25438 }),
  .B2({ S25642 }),
  .ZN({ S25719 })
);
NAND2_X1 #() 
NAND2_X1_4551_ (
  .A1({ S25619 }),
  .A2({ S25416 }),
  .ZN({ S25720 })
);
OAI21_X1 #() 
OAI21_X1_2338_ (
  .A({ S25957[909] }),
  .B1({ S25719 }),
  .B2({ S25720 }),
  .ZN({ S25721 })
);
OAI22_X1 #() 
OAI22_X1_118_ (
  .A1({ S25717 }),
  .A2({ S25957[909] }),
  .B1({ S25721 }),
  .B2({ S25718 }),
  .ZN({ S25722 })
);
NAND2_X1 #() 
NAND2_X1_4552_ (
  .A1({ S25722 }),
  .A2({ S25957[910] }),
  .ZN({ S25723 })
);
NAND3_X1 #() 
NAND3_X1_4942_ (
  .A1({ S25442 }),
  .A2({ S97 }),
  .A3({ S25957[907] }),
  .ZN({ S25724 })
);
NAND2_X1 #() 
NAND2_X1_4553_ (
  .A1({ S25547 }),
  .A2({ S25444 }),
  .ZN({ S25725 })
);
NAND3_X1 #() 
NAND3_X1_4943_ (
  .A1({ S25725 }),
  .A2({ S89 }),
  .A3({ S25539 }),
  .ZN({ S25726 })
);
AND2_X1 #() 
AND2_X1_282_ (
  .A1({ S25726 }),
  .A2({ S25724 }),
  .ZN({ S25727 })
);
NAND2_X1 #() 
NAND2_X1_4554_ (
  .A1({ S25694 }),
  .A2({ S25486 }),
  .ZN({ S25728 })
);
OAI211_X1 #() 
OAI211_X1_1571_ (
  .A({ S25728 }),
  .B({ S25957[908] }),
  .C1({ S25462 }),
  .C2({ S25425 }),
  .ZN({ S25729 })
);
OAI211_X1 #() 
OAI211_X1_1572_ (
  .A({ S25484 }),
  .B({ S25729 }),
  .C1({ S25727 }),
  .C2({ S25957[908] }),
  .ZN({ S25730 })
);
NAND2_X1 #() 
NAND2_X1_4555_ (
  .A1({ S25642 }),
  .A2({ S89 }),
  .ZN({ S25731 })
);
NAND3_X1 #() 
NAND3_X1_4944_ (
  .A1({ S25584 }),
  .A2({ S25731 }),
  .A3({ S25957[908] }),
  .ZN({ S25732 })
);
OAI221_X1 #() 
OAI221_X1_134_ (
  .A({ S25416 }),
  .B1({ S25512 }),
  .B2({ S25444 }),
  .C1({ S25438 }),
  .C2({ S89 }),
  .ZN({ S25733 })
);
NAND2_X1 #() 
NAND2_X1_4556_ (
  .A1({ S25733 }),
  .A2({ S25732 }),
  .ZN({ S25734 })
);
AOI21_X1 #() 
AOI21_X1_2518_ (
  .A({ S25957[910] }),
  .B1({ S25734 }),
  .B2({ S25957[909] }),
  .ZN({ S25735 })
);
NAND2_X1 #() 
NAND2_X1_4557_ (
  .A1({ S25735 }),
  .A2({ S25730 }),
  .ZN({ S25736 })
);
AOI21_X1 #() 
AOI21_X1_2519_ (
  .A({ S25957[911] }),
  .B1({ S25723 }),
  .B2({ S25736 }),
  .ZN({ S25737 })
);
OAI21_X1 #() 
OAI21_X1_2339_ (
  .A({ S25678 }),
  .B1({ S25712 }),
  .B2({ S25737 }),
  .ZN({ S25738 })
);
AND2_X1 #() 
AND2_X1_283_ (
  .A1({ S25723 }),
  .A2({ S25736 }),
  .ZN({ S25739 })
);
OAI211_X1 #() 
OAI211_X1_1573_ (
  .A({ S25711 }),
  .B({ S25957[1012] }),
  .C1({ S25739 }),
  .C2({ S25957[911] }),
  .ZN({ S25740 })
);
AOI21_X1 #() 
AOI21_X1_2520_ (
  .A({ S25957[980] }),
  .B1({ S25738 }),
  .B2({ S25740 }),
  .ZN({ S25741 })
);
INV_X1 #() 
INV_X1_1479_ (
  .A({ S25957[980] }),
  .ZN({ S25742 })
);
OAI211_X1 #() 
OAI211_X1_1574_ (
  .A({ S25711 }),
  .B({ S25678 }),
  .C1({ S25739 }),
  .C2({ S25957[911] }),
  .ZN({ S25743 })
);
OAI21_X1 #() 
OAI21_X1_2340_ (
  .A({ S25957[1012] }),
  .B1({ S25712 }),
  .B2({ S25737 }),
  .ZN({ S25744 })
);
AOI21_X1 #() 
AOI21_X1_2521_ (
  .A({ S25742 }),
  .B1({ S25744 }),
  .B2({ S25743 }),
  .ZN({ S25745 })
);
OAI21_X1 #() 
OAI21_X1_2341_ (
  .A({ S24776 }),
  .B1({ S25741 }),
  .B2({ S25745 }),
  .ZN({ S25746 })
);
NAND3_X1 #() 
NAND3_X1_4945_ (
  .A1({ S25744 }),
  .A2({ S25743 }),
  .A3({ S25742 }),
  .ZN({ S25747 })
);
NAND3_X1 #() 
NAND3_X1_4946_ (
  .A1({ S25738 }),
  .A2({ S25740 }),
  .A3({ S25957[980] }),
  .ZN({ S25748 })
);
NAND3_X1 #() 
NAND3_X1_4947_ (
  .A1({ S25747 }),
  .A2({ S25748 }),
  .A3({ S25957[1044] }),
  .ZN({ S25749 })
);
AND2_X1 #() 
AND2_X1_284_ (
  .A1({ S25746 }),
  .A2({ S25749 }),
  .ZN({ S25957[788] })
);
NAND2_X1 #() 
NAND2_X1_4558_ (
  .A1({ S23077 }),
  .A2({ S23074 }),
  .ZN({ S25750 })
);
NAND2_X1 #() 
NAND2_X1_4559_ (
  .A1({ S20536 }),
  .A2({ S20540 }),
  .ZN({ S25751 })
);
INV_X1 #() 
INV_X1_1480_ (
  .A({ S25751 }),
  .ZN({ S25957[1107] })
);
NAND2_X1 #() 
NAND2_X1_4560_ (
  .A1({ S25509 }),
  .A2({ S25442 }),
  .ZN({ S25752 })
);
AOI22_X1 #() 
AOI22_X1_521_ (
  .A1({ S25752 }),
  .A2({ S25957[907] }),
  .B1({ S25491 }),
  .B2({ S25492 }),
  .ZN({ S25753 })
);
OAI21_X1 #() 
OAI21_X1_2342_ (
  .A({ S97 }),
  .B1({ S25437 }),
  .B2({ S25957[906] }),
  .ZN({ S25754 })
);
NAND2_X1 #() 
NAND2_X1_4561_ (
  .A1({ S25754 }),
  .A2({ S25957[907] }),
  .ZN({ S25755 })
);
AOI21_X1 #() 
AOI21_X1_2522_ (
  .A({ S25416 }),
  .B1({ S25478 }),
  .B2({ S25583 }),
  .ZN({ S25756 })
);
NAND2_X1 #() 
NAND2_X1_4562_ (
  .A1({ S25756 }),
  .A2({ S25755 }),
  .ZN({ S25757 })
);
OAI211_X1 #() 
OAI211_X1_1575_ (
  .A({ S25757 }),
  .B({ S25484 }),
  .C1({ S25753 }),
  .C2({ S25957[908] }),
  .ZN({ S25758 })
);
AOI21_X1 #() 
AOI21_X1_2523_ (
  .A({ S25957[907] }),
  .B1({ S25474 }),
  .B2({ S25957[906] }),
  .ZN({ S25759 })
);
OAI21_X1 #() 
OAI21_X1_2343_ (
  .A({ S25957[907] }),
  .B1({ S97 }),
  .B2({ S25436 }),
  .ZN({ S25760 })
);
NAND2_X1 #() 
NAND2_X1_4563_ (
  .A1({ S25760 }),
  .A2({ S25957[908] }),
  .ZN({ S25761 })
);
NAND4_X1 #() 
NAND4_X1_532_ (
  .A1({ S25464 }),
  .A2({ S25570 }),
  .A3({ S25957[904] }),
  .A4({ S25416 }),
  .ZN({ S25762 })
);
OAI21_X1 #() 
OAI21_X1_2344_ (
  .A({ S25762 }),
  .B1({ S25759 }),
  .B2({ S25761 }),
  .ZN({ S25763 })
);
AOI21_X1 #() 
AOI21_X1_2524_ (
  .A({ S25957[910] }),
  .B1({ S25763 }),
  .B2({ S25957[909] }),
  .ZN({ S25764 })
);
NAND2_X1 #() 
NAND2_X1_4564_ (
  .A1({ S25764 }),
  .A2({ S25758 }),
  .ZN({ S25765 })
);
NAND3_X1 #() 
NAND3_X1_4948_ (
  .A1({ S25437 }),
  .A2({ S89 }),
  .A3({ S25442 }),
  .ZN({ S25766 })
);
NOR2_X1 #() 
NOR2_X1_1152_ (
  .A1({ S25766 }),
  .A2({ S25416 }),
  .ZN({ S25767 })
);
INV_X1 #() 
INV_X1_1481_ (
  .A({ S25767 }),
  .ZN({ S25768 })
);
OAI21_X1 #() 
OAI21_X1_2345_ (
  .A({ S89 }),
  .B1({ S25504 }),
  .B2({ S25684 }),
  .ZN({ S25769 })
);
NAND3_X1 #() 
NAND3_X1_4949_ (
  .A1({ S25769 }),
  .A2({ S25416 }),
  .A3({ S25728 }),
  .ZN({ S25770 })
);
NAND2_X1 #() 
NAND2_X1_4565_ (
  .A1({ S25770 }),
  .A2({ S25768 }),
  .ZN({ S25771 })
);
NAND3_X1 #() 
NAND3_X1_4950_ (
  .A1({ S25516 }),
  .A2({ S25551 }),
  .A3({ S25957[908] }),
  .ZN({ S25772 })
);
NAND2_X1 #() 
NAND2_X1_4566_ (
  .A1({ S25531 }),
  .A2({ S25957[907] }),
  .ZN({ S25773 })
);
NAND2_X1 #() 
NAND2_X1_4567_ (
  .A1({ S25417 }),
  .A2({ S97 }),
  .ZN({ S25774 })
);
AOI21_X1 #() 
AOI21_X1_2525_ (
  .A({ S25957[908] }),
  .B1({ S25774 }),
  .B2({ S89 }),
  .ZN({ S25775 })
);
AOI21_X1 #() 
AOI21_X1_2526_ (
  .A({ S25484 }),
  .B1({ S25775 }),
  .B2({ S25773 }),
  .ZN({ S25776 })
);
AOI22_X1 #() 
AOI22_X1_522_ (
  .A1({ S25771 }),
  .A2({ S25484 }),
  .B1({ S25772 }),
  .B2({ S25776 }),
  .ZN({ S25777 })
);
OAI211_X1 #() 
OAI211_X1_1576_ (
  .A({ S25568 }),
  .B({ S25765 }),
  .C1({ S25777 }),
  .C2({ S23551 }),
  .ZN({ S25778 })
);
NAND2_X1 #() 
NAND2_X1_4568_ (
  .A1({ S25550 }),
  .A2({ S89 }),
  .ZN({ S25779 })
);
AOI21_X1 #() 
AOI21_X1_2527_ (
  .A({ S89 }),
  .B1({ S25547 }),
  .B2({ S25444 }),
  .ZN({ S25780 })
);
NAND2_X1 #() 
NAND2_X1_4569_ (
  .A1({ S25780 }),
  .A2({ S25438 }),
  .ZN({ S25781 })
);
NAND3_X1 #() 
NAND3_X1_4951_ (
  .A1({ S25779 }),
  .A2({ S25781 }),
  .A3({ S25957[908] }),
  .ZN({ S25782 })
);
NAND4_X1 #() 
NAND4_X1_533_ (
  .A1({ S25429 }),
  .A2({ S25433 }),
  .A3({ S25957[905] }),
  .A4({ S25957[907] }),
  .ZN({ S25783 })
);
OAI211_X1 #() 
OAI211_X1_1577_ (
  .A({ S25536 }),
  .B({ S89 }),
  .C1({ S25455 }),
  .C2({ S96 }),
  .ZN({ S25784 })
);
NAND3_X1 #() 
NAND3_X1_4952_ (
  .A1({ S25784 }),
  .A2({ S25416 }),
  .A3({ S25783 }),
  .ZN({ S25785 })
);
NAND3_X1 #() 
NAND3_X1_4953_ (
  .A1({ S25782 }),
  .A2({ S25957[909] }),
  .A3({ S25785 }),
  .ZN({ S25786 })
);
NAND2_X1 #() 
NAND2_X1_4570_ (
  .A1({ S25493 }),
  .A2({ S25957[907] }),
  .ZN({ S25787 })
);
NAND3_X1 #() 
NAND3_X1_4954_ (
  .A1({ S25787 }),
  .A2({ S25706 }),
  .A3({ S25957[908] }),
  .ZN({ S25788 })
);
INV_X1 #() 
INV_X1_1482_ (
  .A({ S25435 }),
  .ZN({ S25789 })
);
NAND3_X1 #() 
NAND3_X1_4955_ (
  .A1({ S25421 }),
  .A2({ S89 }),
  .A3({ S25442 }),
  .ZN({ S25790 })
);
OAI211_X1 #() 
OAI211_X1_1578_ (
  .A({ S25416 }),
  .B({ S25790 }),
  .C1({ S25789 }),
  .C2({ S25537 }),
  .ZN({ S25791 })
);
NAND3_X1 #() 
NAND3_X1_4956_ (
  .A1({ S25791 }),
  .A2({ S25788 }),
  .A3({ S25484 }),
  .ZN({ S25792 })
);
NAND3_X1 #() 
NAND3_X1_4957_ (
  .A1({ S25786 }),
  .A2({ S25792 }),
  .A3({ S23551 }),
  .ZN({ S25793 })
);
OAI211_X1 #() 
OAI211_X1_1579_ (
  .A({ S25549 }),
  .B({ S25957[907] }),
  .C1({ S25957[906] }),
  .C2({ S25460 }),
  .ZN({ S25794 })
);
NAND4_X1 #() 
NAND4_X1_534_ (
  .A1({ S25421 }),
  .A2({ S89 }),
  .A3({ S25429 }),
  .A4({ S25422 }),
  .ZN({ S25795 })
);
AOI21_X1 #() 
AOI21_X1_2528_ (
  .A({ S25957[908] }),
  .B1({ S25794 }),
  .B2({ S25795 }),
  .ZN({ S25796 })
);
NAND3_X1 #() 
NAND3_X1_4958_ (
  .A1({ S25421 }),
  .A2({ S25957[907] }),
  .A3({ S25433 }),
  .ZN({ S25797 })
);
NAND4_X1 #() 
NAND4_X1_535_ (
  .A1({ S25570 }),
  .A2({ S25437 }),
  .A3({ S97 }),
  .A4({ S89 }),
  .ZN({ S25798 })
);
AOI21_X1 #() 
AOI21_X1_2529_ (
  .A({ S25416 }),
  .B1({ S25798 }),
  .B2({ S25797 }),
  .ZN({ S25799 })
);
NOR3_X1 #() 
NOR3_X1_152_ (
  .A1({ S25796 }),
  .A2({ S25799 }),
  .A3({ S25484 }),
  .ZN({ S25800 })
);
NAND3_X1 #() 
NAND3_X1_4959_ (
  .A1({ S25435 }),
  .A2({ S89 }),
  .A3({ S25583 }),
  .ZN({ S25801 })
);
AOI21_X1 #() 
AOI21_X1_2530_ (
  .A({ S25416 }),
  .B1({ S25801 }),
  .B2({ S25557 }),
  .ZN({ S25802 })
);
OAI211_X1 #() 
OAI211_X1_1580_ (
  .A({ S25574 }),
  .B({ S25416 }),
  .C1({ S89 }),
  .C2({ S25436 }),
  .ZN({ S25803 })
);
NAND2_X1 #() 
NAND2_X1_4571_ (
  .A1({ S25803 }),
  .A2({ S25484 }),
  .ZN({ S25804 })
);
OAI21_X1 #() 
OAI21_X1_2346_ (
  .A({ S25957[910] }),
  .B1({ S25802 }),
  .B2({ S25804 }),
  .ZN({ S25805 })
);
OAI211_X1 #() 
OAI211_X1_1581_ (
  .A({ S25793 }),
  .B({ S25957[911] }),
  .C1({ S25800 }),
  .C2({ S25805 }),
  .ZN({ S25806 })
);
NAND3_X1 #() 
NAND3_X1_4960_ (
  .A1({ S25778 }),
  .A2({ S25806 }),
  .A3({ S25957[1107] }),
  .ZN({ S25807 })
);
AND3_X1 #() 
AND3_X1_177_ (
  .A1({ S25786 }),
  .A2({ S25792 }),
  .A3({ S23551 }),
  .ZN({ S25808 })
);
NOR2_X1 #() 
NOR2_X1_1153_ (
  .A1({ S25805 }),
  .A2({ S25800 }),
  .ZN({ S25809 })
);
OAI21_X1 #() 
OAI21_X1_2347_ (
  .A({ S25957[911] }),
  .B1({ S25808 }),
  .B2({ S25809 }),
  .ZN({ S25810 })
);
OAI211_X1 #() 
OAI211_X1_1582_ (
  .A({ S25615 }),
  .B({ S25957[908] }),
  .C1({ S25754 }),
  .C2({ S89 }),
  .ZN({ S25811 })
);
NOR2_X1 #() 
NOR2_X1_1154_ (
  .A1({ S25470 }),
  .A2({ S25957[908] }),
  .ZN({ S25812 })
);
OAI211_X1 #() 
OAI211_X1_1583_ (
  .A({ S25812 }),
  .B({ S25500 }),
  .C1({ S25579 }),
  .C2({ S25434 }),
  .ZN({ S25813 })
);
NAND3_X1 #() 
NAND3_X1_4961_ (
  .A1({ S25813 }),
  .A2({ S25484 }),
  .A3({ S25811 }),
  .ZN({ S25814 })
);
OAI211_X1 #() 
OAI211_X1_1584_ (
  .A({ S25957[909] }),
  .B({ S25762 }),
  .C1({ S25759 }),
  .C2({ S25761 }),
  .ZN({ S25815 })
);
AOI21_X1 #() 
AOI21_X1_2531_ (
  .A({ S25957[910] }),
  .B1({ S25814 }),
  .B2({ S25815 }),
  .ZN({ S25816 })
);
AND2_X1 #() 
AND2_X1_285_ (
  .A1({ S25471 }),
  .A2({ S25446 }),
  .ZN({ S25817 })
);
AOI21_X1 #() 
AOI21_X1_2532_ (
  .A({ S25957[908] }),
  .B1({ S25817 }),
  .B2({ S25555 }),
  .ZN({ S25818 })
);
OAI21_X1 #() 
OAI21_X1_2348_ (
  .A({ S25484 }),
  .B1({ S25818 }),
  .B2({ S25767 }),
  .ZN({ S25819 })
);
NAND2_X1 #() 
NAND2_X1_4572_ (
  .A1({ S25570 }),
  .A2({ S89 }),
  .ZN({ S25820 })
);
OAI211_X1 #() 
OAI211_X1_1585_ (
  .A({ S25773 }),
  .B({ S25416 }),
  .C1({ S25679 }),
  .C2({ S25820 }),
  .ZN({ S25821 })
);
NAND3_X1 #() 
NAND3_X1_4962_ (
  .A1({ S25772 }),
  .A2({ S25957[909] }),
  .A3({ S25821 }),
  .ZN({ S25822 })
);
AOI21_X1 #() 
AOI21_X1_2533_ (
  .A({ S23551 }),
  .B1({ S25819 }),
  .B2({ S25822 }),
  .ZN({ S25823 })
);
OAI21_X1 #() 
OAI21_X1_2349_ (
  .A({ S25568 }),
  .B1({ S25823 }),
  .B2({ S25816 }),
  .ZN({ S25824 })
);
NAND3_X1 #() 
NAND3_X1_4963_ (
  .A1({ S25810 }),
  .A2({ S25824 }),
  .A3({ S25751 }),
  .ZN({ S25825 })
);
AOI21_X1 #() 
AOI21_X1_2534_ (
  .A({ S25750 }),
  .B1({ S25825 }),
  .B2({ S25807 }),
  .ZN({ S25826 })
);
AND3_X1 #() 
AND3_X1_178_ (
  .A1({ S25825 }),
  .A2({ S25807 }),
  .A3({ S25750 }),
  .ZN({ S25827 })
);
OAI21_X1 #() 
OAI21_X1_2350_ (
  .A({ S86 }),
  .B1({ S25827 }),
  .B2({ S25826 }),
  .ZN({ S25828 })
);
INV_X1 #() 
INV_X1_1483_ (
  .A({ S25750 }),
  .ZN({ S25957[947] })
);
AOI21_X1 #() 
AOI21_X1_2535_ (
  .A({ S25751 }),
  .B1({ S25810 }),
  .B2({ S25824 }),
  .ZN({ S25829 })
);
AOI21_X1 #() 
AOI21_X1_2536_ (
  .A({ S25957[1107] }),
  .B1({ S25778 }),
  .B2({ S25806 }),
  .ZN({ S25830 })
);
OAI21_X1 #() 
OAI21_X1_2351_ (
  .A({ S25957[947] }),
  .B1({ S25829 }),
  .B2({ S25830 }),
  .ZN({ S25831 })
);
NAND3_X1 #() 
NAND3_X1_4964_ (
  .A1({ S25825 }),
  .A2({ S25807 }),
  .A3({ S25750 }),
  .ZN({ S25832 })
);
NAND3_X1 #() 
NAND3_X1_4965_ (
  .A1({ S25831 }),
  .A2({ S25957[915] }),
  .A3({ S25832 }),
  .ZN({ S25833 })
);
NAND2_X1 #() 
NAND2_X1_4573_ (
  .A1({ S25828 }),
  .A2({ S25833 }),
  .ZN({ S98 })
);
AND2_X1 #() 
AND2_X1_286_ (
  .A1({ S25828 }),
  .A2({ S25833 }),
  .ZN({ S25957[787] })
);
NAND2_X1 #() 
NAND2_X1_4574_ (
  .A1({ S23199 }),
  .A2({ S23203 }),
  .ZN({ S25834 })
);
INV_X1 #() 
INV_X1_1484_ (
  .A({ S25834 }),
  .ZN({ S25957[944] })
);
XNOR2_X1 #() 
XNOR2_X1_182_ (
  .A({ S25957[1136] }),
  .B({ S23196 }),
  .ZN({ S25957[1104] })
);
INV_X1 #() 
INV_X1_1485_ (
  .A({ S25957[1104] }),
  .ZN({ S25835 })
);
NAND2_X1 #() 
NAND2_X1_4575_ (
  .A1({ S25766 }),
  .A2({ S25760 }),
  .ZN({ S25836 })
);
AOI21_X1 #() 
AOI21_X1_2537_ (
  .A({ S25416 }),
  .B1({ S25531 }),
  .B2({ S89 }),
  .ZN({ S25837 })
);
NAND3_X1 #() 
NAND3_X1_4966_ (
  .A1({ S25699 }),
  .A2({ S25471 }),
  .A3({ S25643 }),
  .ZN({ S25838 })
);
AOI22_X1 #() 
AOI22_X1_523_ (
  .A1({ S25837 }),
  .A2({ S25836 }),
  .B1({ S25838 }),
  .B2({ S25416 }),
  .ZN({ S25839 })
);
NAND4_X1 #() 
NAND4_X1_536_ (
  .A1({ S25469 }),
  .A2({ S25442 }),
  .A3({ S97 }),
  .A4({ S89 }),
  .ZN({ S25840 })
);
AOI21_X1 #() 
AOI21_X1_2538_ (
  .A({ S25957[908] }),
  .B1({ S25773 }),
  .B2({ S25840 }),
  .ZN({ S25841 })
);
NAND3_X1 #() 
NAND3_X1_4967_ (
  .A1({ S25957[906] }),
  .A2({ S25957[907] }),
  .A3({ S25957[905] }),
  .ZN({ S25842 })
);
NAND4_X1 #() 
NAND4_X1_537_ (
  .A1({ S25437 }),
  .A2({ S97 }),
  .A3({ S89 }),
  .A4({ S25436 }),
  .ZN({ S25843 })
);
AND3_X1 #() 
AND3_X1_179_ (
  .A1({ S25843 }),
  .A2({ S25842 }),
  .A3({ S25957[908] }),
  .ZN({ S25844 })
);
OAI21_X1 #() 
OAI21_X1_2352_ (
  .A({ S25484 }),
  .B1({ S25844 }),
  .B2({ S25841 }),
  .ZN({ S25845 })
);
OAI211_X1 #() 
OAI211_X1_1586_ (
  .A({ S25845 }),
  .B({ S23551 }),
  .C1({ S25484 }),
  .C2({ S25839 }),
  .ZN({ S25846 })
);
AOI21_X1 #() 
AOI21_X1_2539_ (
  .A({ S25408 }),
  .B1({ S25427 }),
  .B2({ S25428 }),
  .ZN({ S25847 })
);
AOI21_X1 #() 
AOI21_X1_2540_ (
  .A({ S25847 }),
  .B1({ S25422 }),
  .B2({ S25957[906] }),
  .ZN({ S25848 })
);
NAND3_X1 #() 
NAND3_X1_4968_ (
  .A1({ S25444 }),
  .A2({ S89 }),
  .A3({ S25436 }),
  .ZN({ S25849 })
);
NAND4_X1 #() 
NAND4_X1_538_ (
  .A1({ S25421 }),
  .A2({ S25422 }),
  .A3({ S25957[907] }),
  .A4({ S25957[906] }),
  .ZN({ S25850 })
);
OAI211_X1 #() 
OAI211_X1_1587_ (
  .A({ S25849 }),
  .B({ S25850 }),
  .C1({ S25848 }),
  .C2({ S25957[907] }),
  .ZN({ S25851 })
);
AOI21_X1 #() 
AOI21_X1_2541_ (
  .A({ S25620 }),
  .B1({ S25851 }),
  .B2({ S25957[908] }),
  .ZN({ S25852 })
);
AOI21_X1 #() 
AOI21_X1_2542_ (
  .A({ S25957[907] }),
  .B1({ S25438 }),
  .B2({ S25417 }),
  .ZN({ S25853 })
);
NAND2_X1 #() 
NAND2_X1_4576_ (
  .A1({ S25728 }),
  .A2({ S25416 }),
  .ZN({ S25854 })
);
NAND3_X1 #() 
NAND3_X1_4969_ (
  .A1({ S25421 }),
  .A2({ S25957[907] }),
  .A3({ S25957[906] }),
  .ZN({ S25855 })
);
NAND3_X1 #() 
NAND3_X1_4970_ (
  .A1({ S25726 }),
  .A2({ S25957[908] }),
  .A3({ S25855 }),
  .ZN({ S25856 })
);
OAI211_X1 #() 
OAI211_X1_1588_ (
  .A({ S25856 }),
  .B({ S25957[909] }),
  .C1({ S25854 }),
  .C2({ S25853 }),
  .ZN({ S25857 })
);
OAI211_X1 #() 
OAI211_X1_1589_ (
  .A({ S25957[910] }),
  .B({ S25857 }),
  .C1({ S25852 }),
  .C2({ S25957[909] }),
  .ZN({ S25858 })
);
NAND3_X1 #() 
NAND3_X1_4971_ (
  .A1({ S25858 }),
  .A2({ S25957[911] }),
  .A3({ S25846 }),
  .ZN({ S25859 })
);
NAND3_X1 #() 
NAND3_X1_4972_ (
  .A1({ S25491 }),
  .A2({ S25957[907] }),
  .A3({ S25539 }),
  .ZN({ S25860 })
);
NOR2_X1 #() 
NOR2_X1_1155_ (
  .A1({ S97 }),
  .A2({ S25436 }),
  .ZN({ S25861 })
);
OAI21_X1 #() 
OAI21_X1_2353_ (
  .A({ S89 }),
  .B1({ S25861 }),
  .B2({ S25592 }),
  .ZN({ S25862 })
);
NAND3_X1 #() 
NAND3_X1_4973_ (
  .A1({ S25860 }),
  .A2({ S25862 }),
  .A3({ S25416 }),
  .ZN({ S25863 })
);
NAND4_X1 #() 
NAND4_X1_539_ (
  .A1({ S25787 }),
  .A2({ S25849 }),
  .A3({ S25518 }),
  .A4({ S25957[908] }),
  .ZN({ S25864 })
);
NAND3_X1 #() 
NAND3_X1_4974_ (
  .A1({ S25863 }),
  .A2({ S25864 }),
  .A3({ S25484 }),
  .ZN({ S25865 })
);
NAND3_X1 #() 
NAND3_X1_4975_ (
  .A1({ S25613 }),
  .A2({ S25957[908] }),
  .A3({ S25724 }),
  .ZN({ S25866 })
);
NAND3_X1 #() 
NAND3_X1_4976_ (
  .A1({ S25631 }),
  .A2({ S25416 }),
  .A3({ S25560 }),
  .ZN({ S25867 })
);
NAND3_X1 #() 
NAND3_X1_4977_ (
  .A1({ S25867 }),
  .A2({ S25866 }),
  .A3({ S25957[909] }),
  .ZN({ S25868 })
);
NAND3_X1 #() 
NAND3_X1_4978_ (
  .A1({ S25865 }),
  .A2({ S23551 }),
  .A3({ S25868 }),
  .ZN({ S25869 })
);
OAI21_X1 #() 
OAI21_X1_2354_ (
  .A({ S25957[907] }),
  .B1({ S25586 }),
  .B2({ S25587 }),
  .ZN({ S25870 })
);
NAND2_X1 #() 
NAND2_X1_4577_ (
  .A1({ S96 }),
  .A2({ S25957[906] }),
  .ZN({ S25871 })
);
NAND4_X1 #() 
NAND4_X1_540_ (
  .A1({ S25509 }),
  .A2({ S25871 }),
  .A3({ S25957[907] }),
  .A4({ S97 }),
  .ZN({ S25872 })
);
AOI21_X1 #() 
AOI21_X1_2543_ (
  .A({ S25416 }),
  .B1({ S25461 }),
  .B2({ S25429 }),
  .ZN({ S25873 })
);
NOR2_X1 #() 
NOR2_X1_1156_ (
  .A1({ S25498 }),
  .A2({ S25957[908] }),
  .ZN({ S25874 })
);
AOI22_X1 #() 
AOI22_X1_524_ (
  .A1({ S25874 }),
  .A2({ S25870 }),
  .B1({ S25872 }),
  .B2({ S25873 }),
  .ZN({ S25875 })
);
NAND4_X1 #() 
NAND4_X1_541_ (
  .A1({ S25610 }),
  .A2({ S25612 }),
  .A3({ S25957[908] }),
  .A4({ S25463 }),
  .ZN({ S25876 })
);
NAND3_X1 #() 
NAND3_X1_4979_ (
  .A1({ S25536 }),
  .A2({ S89 }),
  .A3({ S97 }),
  .ZN({ S25877 })
);
NAND3_X1 #() 
NAND3_X1_4980_ (
  .A1({ S25877 }),
  .A2({ S25416 }),
  .A3({ S25619 }),
  .ZN({ S25878 })
);
NAND3_X1 #() 
NAND3_X1_4981_ (
  .A1({ S25878 }),
  .A2({ S25484 }),
  .A3({ S25876 }),
  .ZN({ S25879 })
);
OAI211_X1 #() 
OAI211_X1_1590_ (
  .A({ S25957[910] }),
  .B({ S25879 }),
  .C1({ S25875 }),
  .C2({ S25484 }),
  .ZN({ S25880 })
);
NAND3_X1 #() 
NAND3_X1_4982_ (
  .A1({ S25880 }),
  .A2({ S25869 }),
  .A3({ S25568 }),
  .ZN({ S25881 })
);
NAND3_X1 #() 
NAND3_X1_4983_ (
  .A1({ S25859 }),
  .A2({ S25881 }),
  .A3({ S25835 }),
  .ZN({ S25882 })
);
AOI21_X1 #() 
AOI21_X1_2544_ (
  .A({ S25416 }),
  .B1({ S25682 }),
  .B2({ S25850 }),
  .ZN({ S25883 })
);
NOR3_X1 #() 
NOR3_X1_153_ (
  .A1({ S25883 }),
  .A2({ S25620 }),
  .A3({ S25957[909] }),
  .ZN({ S25884 })
);
AOI21_X1 #() 
AOI21_X1_2545_ (
  .A({ S25957[908] }),
  .B1({ S25424 }),
  .B2({ S25728 }),
  .ZN({ S25885 })
);
AOI21_X1 #() 
AOI21_X1_2546_ (
  .A({ S89 }),
  .B1({ S25463 }),
  .B2({ S25442 }),
  .ZN({ S25886 })
);
AOI21_X1 #() 
AOI21_X1_2547_ (
  .A({ S25886 }),
  .B1({ S25458 }),
  .B2({ S89 }),
  .ZN({ S25887 })
);
OAI21_X1 #() 
OAI21_X1_2355_ (
  .A({ S25957[909] }),
  .B1({ S25887 }),
  .B2({ S25416 }),
  .ZN({ S25888 })
);
OAI21_X1 #() 
OAI21_X1_2356_ (
  .A({ S25957[910] }),
  .B1({ S25888 }),
  .B2({ S25885 }),
  .ZN({ S25889 })
);
NAND2_X1 #() 
NAND2_X1_4578_ (
  .A1({ S25836 }),
  .A2({ S25837 }),
  .ZN({ S25890 })
);
NAND2_X1 #() 
NAND2_X1_4579_ (
  .A1({ S25838 }),
  .A2({ S25416 }),
  .ZN({ S25891 })
);
NAND3_X1 #() 
NAND3_X1_4984_ (
  .A1({ S25891 }),
  .A2({ S25890 }),
  .A3({ S25957[909] }),
  .ZN({ S25892 })
);
NAND2_X1 #() 
NAND2_X1_4580_ (
  .A1({ S25502 }),
  .A2({ S25843 }),
  .ZN({ S25893 })
);
NAND2_X1 #() 
NAND2_X1_4581_ (
  .A1({ S25893 }),
  .A2({ S25484 }),
  .ZN({ S25894 })
);
OAI211_X1 #() 
OAI211_X1_1591_ (
  .A({ S25892 }),
  .B({ S23551 }),
  .C1({ S25841 }),
  .C2({ S25894 }),
  .ZN({ S25895 })
);
OAI211_X1 #() 
OAI211_X1_1592_ (
  .A({ S25957[911] }),
  .B({ S25895 }),
  .C1({ S25889 }),
  .C2({ S25884 }),
  .ZN({ S25896 })
);
NAND2_X1 #() 
NAND2_X1_4582_ (
  .A1({ S25878 }),
  .A2({ S25876 }),
  .ZN({ S25897 })
);
NAND2_X1 #() 
NAND2_X1_4583_ (
  .A1({ S25897 }),
  .A2({ S25484 }),
  .ZN({ S25898 })
);
AND2_X1 #() 
AND2_X1_287_ (
  .A1({ S25872 }),
  .A2({ S25873 }),
  .ZN({ S25899 })
);
NAND2_X1 #() 
NAND2_X1_4584_ (
  .A1({ S25870 }),
  .A2({ S25874 }),
  .ZN({ S25900 })
);
NAND2_X1 #() 
NAND2_X1_4585_ (
  .A1({ S25900 }),
  .A2({ S25957[909] }),
  .ZN({ S25901 })
);
OAI211_X1 #() 
OAI211_X1_1593_ (
  .A({ S25898 }),
  .B({ S25957[910] }),
  .C1({ S25901 }),
  .C2({ S25899 }),
  .ZN({ S25902 })
);
NAND2_X1 #() 
NAND2_X1_4586_ (
  .A1({ S25867 }),
  .A2({ S25866 }),
  .ZN({ S25903 })
);
NAND2_X1 #() 
NAND2_X1_4587_ (
  .A1({ S25903 }),
  .A2({ S25957[909] }),
  .ZN({ S25904 })
);
NAND3_X1 #() 
NAND3_X1_4985_ (
  .A1({ S25787 }),
  .A2({ S25518 }),
  .A3({ S25849 }),
  .ZN({ S25905 })
);
NAND2_X1 #() 
NAND2_X1_4588_ (
  .A1({ S25905 }),
  .A2({ S25957[908] }),
  .ZN({ S25906 })
);
NAND3_X1 #() 
NAND3_X1_4986_ (
  .A1({ S25871 }),
  .A2({ S25957[907] }),
  .A3({ S97 }),
  .ZN({ S25907 })
);
NAND3_X1 #() 
NAND3_X1_4987_ (
  .A1({ S25583 }),
  .A2({ S25725 }),
  .A3({ S89 }),
  .ZN({ S25908 })
);
NAND3_X1 #() 
NAND3_X1_4988_ (
  .A1({ S25908 }),
  .A2({ S25907 }),
  .A3({ S25416 }),
  .ZN({ S25909 })
);
NAND3_X1 #() 
NAND3_X1_4989_ (
  .A1({ S25906 }),
  .A2({ S25484 }),
  .A3({ S25909 }),
  .ZN({ S25910 })
);
NAND3_X1 #() 
NAND3_X1_4990_ (
  .A1({ S25910 }),
  .A2({ S25904 }),
  .A3({ S23551 }),
  .ZN({ S25911 })
);
NAND3_X1 #() 
NAND3_X1_4991_ (
  .A1({ S25911 }),
  .A2({ S25902 }),
  .A3({ S25568 }),
  .ZN({ S25912 })
);
NAND3_X1 #() 
NAND3_X1_4992_ (
  .A1({ S25912 }),
  .A2({ S25896 }),
  .A3({ S25957[1104] }),
  .ZN({ S25913 })
);
NAND3_X1 #() 
NAND3_X1_4993_ (
  .A1({ S25913 }),
  .A2({ S25882 }),
  .A3({ S25957[944] }),
  .ZN({ S25914 })
);
AOI21_X1 #() 
AOI21_X1_2548_ (
  .A({ S25957[1104] }),
  .B1({ S25912 }),
  .B2({ S25896 }),
  .ZN({ S25915 })
);
AOI21_X1 #() 
AOI21_X1_2549_ (
  .A({ S25835 }),
  .B1({ S25859 }),
  .B2({ S25881 }),
  .ZN({ S25916 })
);
OAI21_X1 #() 
OAI21_X1_2357_ (
  .A({ S25834 }),
  .B1({ S25915 }),
  .B2({ S25916 }),
  .ZN({ S25917 })
);
NAND3_X1 #() 
NAND3_X1_4994_ (
  .A1({ S25917 }),
  .A2({ S25957[912] }),
  .A3({ S25914 }),
  .ZN({ S25918 })
);
NAND3_X1 #() 
NAND3_X1_4995_ (
  .A1({ S23199 }),
  .A2({ S23203 }),
  .A3({ S25957[1040] }),
  .ZN({ S25919 })
);
NAND3_X1 #() 
NAND3_X1_4996_ (
  .A1({ S23142 }),
  .A2({ S23191 }),
  .A3({ S23195 }),
  .ZN({ S25920 })
);
NAND2_X1 #() 
NAND2_X1_4589_ (
  .A1({ S25920 }),
  .A2({ S25919 }),
  .ZN({ S25921 })
);
OAI21_X1 #() 
OAI21_X1_2358_ (
  .A({ S25957[944] }),
  .B1({ S25915 }),
  .B2({ S25916 }),
  .ZN({ S25922 })
);
NAND3_X1 #() 
NAND3_X1_4997_ (
  .A1({ S25913 }),
  .A2({ S25882 }),
  .A3({ S25834 }),
  .ZN({ S25923 })
);
NAND3_X1 #() 
NAND3_X1_4998_ (
  .A1({ S25922 }),
  .A2({ S25921 }),
  .A3({ S25923 }),
  .ZN({ S25924 })
);
NAND2_X1 #() 
NAND2_X1_4590_ (
  .A1({ S25918 }),
  .A2({ S25924 }),
  .ZN({ S25957[784] })
);
NAND2_X1 #() 
NAND2_X1_4591_ (
  .A1({ S23241 }),
  .A2({ S23259 }),
  .ZN({ S25957[945] })
);
INV_X1 #() 
INV_X1_1486_ (
  .A({ S25957[945] }),
  .ZN({ S25925 })
);
NAND2_X1 #() 
NAND2_X1_4592_ (
  .A1({ S20672 }),
  .A2({ S20673 }),
  .ZN({ S25926 })
);
INV_X1 #() 
INV_X1_1487_ (
  .A({ S25926 }),
  .ZN({ S25957[1105] })
);
INV_X1 #() 
INV_X1_1488_ (
  .A({ S25457 }),
  .ZN({ S25927 })
);
OAI21_X1 #() 
OAI21_X1_2359_ (
  .A({ S25500 }),
  .B1({ S25927 }),
  .B2({ S25766 }),
  .ZN({ S25928 })
);
AOI21_X1 #() 
AOI21_X1_2550_ (
  .A({ S25957[909] }),
  .B1({ S25611 }),
  .B2({ S25837 }),
  .ZN({ S25929 })
);
OAI21_X1 #() 
OAI21_X1_2360_ (
  .A({ S25929 }),
  .B1({ S25957[908] }),
  .B2({ S25928 }),
  .ZN({ S25930 })
);
AOI21_X1 #() 
AOI21_X1_2551_ (
  .A({ S89 }),
  .B1({ S25491 }),
  .B2({ S25515 }),
  .ZN({ S25931 })
);
OAI21_X1 #() 
OAI21_X1_2361_ (
  .A({ S25416 }),
  .B1({ S25586 }),
  .B2({ S25957[907] }),
  .ZN({ S25932 })
);
NAND3_X1 #() 
NAND3_X1_4999_ (
  .A1({ S25557 }),
  .A2({ S25957[908] }),
  .A3({ S25505 }),
  .ZN({ S25933 })
);
OAI211_X1 #() 
OAI211_X1_1594_ (
  .A({ S25933 }),
  .B({ S25957[909] }),
  .C1({ S25931 }),
  .C2({ S25932 }),
  .ZN({ S25934 })
);
NAND3_X1 #() 
NAND3_X1_5000_ (
  .A1({ S25930 }),
  .A2({ S25957[910] }),
  .A3({ S25934 }),
  .ZN({ S25935 })
);
NOR2_X1 #() 
NOR2_X1_1157_ (
  .A1({ S25579 }),
  .A2({ S25704 }),
  .ZN({ S25936 })
);
NAND2_X1 #() 
NAND2_X1_4593_ (
  .A1({ S25499 }),
  .A2({ S25957[908] }),
  .ZN({ S25937 })
);
OAI21_X1 #() 
OAI21_X1_2362_ (
  .A({ S25957[907] }),
  .B1({ S25460 }),
  .B2({ S25957[906] }),
  .ZN({ S25938 })
);
OAI211_X1 #() 
OAI211_X1_1595_ (
  .A({ S25416 }),
  .B({ S25938 }),
  .C1({ S25820 }),
  .C2({ S25679 }),
  .ZN({ S25939 })
);
OAI211_X1 #() 
OAI211_X1_1596_ (
  .A({ S25957[909] }),
  .B({ S25939 }),
  .C1({ S25937 }),
  .C2({ S25936 }),
  .ZN({ S25940 })
);
NOR3_X1 #() 
NOR3_X1_154_ (
  .A1({ S25494 }),
  .A2({ S25690 }),
  .A3({ S25957[908] }),
  .ZN({ S25941 })
);
AOI21_X1 #() 
AOI21_X1_2552_ (
  .A({ S25957[907] }),
  .B1({ S25556 }),
  .B2({ S25536 }),
  .ZN({ S25942 })
);
OAI21_X1 #() 
OAI21_X1_2363_ (
  .A({ S25484 }),
  .B1({ S25942 }),
  .B2({ S25571 }),
  .ZN({ S25943 })
);
OAI211_X1 #() 
OAI211_X1_1597_ (
  .A({ S25940 }),
  .B({ S23551 }),
  .C1({ S25943 }),
  .C2({ S25941 }),
  .ZN({ S25944 })
);
AND3_X1 #() 
AND3_X1_180_ (
  .A1({ S25944 }),
  .A2({ S25935 }),
  .A3({ S25957[911] }),
  .ZN({ S25945 })
);
NOR2_X1 #() 
NOR2_X1_1158_ (
  .A1({ S25430 }),
  .A2({ S25425 }),
  .ZN({ S25946 })
);
NAND3_X1 #() 
NAND3_X1_5001_ (
  .A1({ S25555 }),
  .A2({ S25416 }),
  .A3({ S25426 }),
  .ZN({ S25947 })
);
OAI211_X1 #() 
OAI211_X1_1598_ (
  .A({ S25947 }),
  .B({ S25484 }),
  .C1({ S25447 }),
  .C2({ S25946 }),
  .ZN({ S25948 })
);
AOI21_X1 #() 
AOI21_X1_2553_ (
  .A({ S25416 }),
  .B1({ S25701 }),
  .B2({ S25783 }),
  .ZN({ S25949 })
);
OAI21_X1 #() 
OAI21_X1_2364_ (
  .A({ S25957[909] }),
  .B1({ S25488 }),
  .B2({ S25949 }),
  .ZN({ S25950 })
);
NAND2_X1 #() 
NAND2_X1_4594_ (
  .A1({ S25950 }),
  .A2({ S25948 }),
  .ZN({ S25951 })
);
NAND2_X1 #() 
NAND2_X1_4595_ (
  .A1({ S25951 }),
  .A2({ S23551 }),
  .ZN({ S25952 })
);
NOR2_X1 #() 
NOR2_X1_1159_ (
  .A1({ S25437 }),
  .A2({ S25436 }),
  .ZN({ S25953 })
);
OAI21_X1 #() 
OAI21_X1_2365_ (
  .A({ S25957[908] }),
  .B1({ S25953 }),
  .B2({ S25449 }),
  .ZN({ S25954 })
);
NAND3_X1 #() 
NAND3_X1_5002_ (
  .A1({ S25850 }),
  .A2({ S25573 }),
  .A3({ S25416 }),
  .ZN({ S25955 })
);
OAI211_X1 #() 
OAI211_X1_1599_ (
  .A({ S25484 }),
  .B({ S25955 }),
  .C1({ S25954 }),
  .C2({ S25931 }),
  .ZN({ S236 })
);
INV_X1 #() 
INV_X1_1489_ (
  .A({ S236 }),
  .ZN({ S237 })
);
AND3_X1 #() 
AND3_X1_181_ (
  .A1({ S25408 }),
  .A2({ S23922 }),
  .A3({ S23925 }),
  .ZN({ S238 })
);
AOI21_X1 #() 
AOI21_X1_2554_ (
  .A({ S238 }),
  .B1({ S96 }),
  .B2({ S25436 }),
  .ZN({ S239 })
);
OAI211_X1 #() 
OAI211_X1_1600_ (
  .A({ S89 }),
  .B({ S25433 }),
  .C1({ S97 }),
  .C2({ S25436 }),
  .ZN({ S240 })
);
OAI21_X1 #() 
OAI21_X1_2366_ (
  .A({ S240 }),
  .B1({ S239 }),
  .B2({ S89 }),
  .ZN({ S241 })
);
NAND2_X1 #() 
NAND2_X1_4596_ (
  .A1({ S241 }),
  .A2({ S25957[908] }),
  .ZN({ S242 })
);
OAI21_X1 #() 
OAI21_X1_2367_ (
  .A({ S25444 }),
  .B1({ S25456 }),
  .B2({ S25957[907] }),
  .ZN({ S243 })
);
AOI21_X1 #() 
AOI21_X1_2555_ (
  .A({ S25957[908] }),
  .B1({ S243 }),
  .B2({ S25442 }),
  .ZN({ S244 })
);
INV_X1 #() 
INV_X1_1490_ (
  .A({ S244 }),
  .ZN({ S245 })
);
AOI21_X1 #() 
AOI21_X1_2556_ (
  .A({ S25484 }),
  .B1({ S242 }),
  .B2({ S245 }),
  .ZN({ S246 })
);
OAI21_X1 #() 
OAI21_X1_2368_ (
  .A({ S25957[910] }),
  .B1({ S246 }),
  .B2({ S237 }),
  .ZN({ S247 })
);
AOI21_X1 #() 
AOI21_X1_2557_ (
  .A({ S25957[911] }),
  .B1({ S247 }),
  .B2({ S25952 }),
  .ZN({ S248 })
);
OAI21_X1 #() 
OAI21_X1_2369_ (
  .A({ S25957[1105] }),
  .B1({ S248 }),
  .B2({ S25945 }),
  .ZN({ S249 })
);
NAND3_X1 #() 
NAND3_X1_5003_ (
  .A1({ S25944 }),
  .A2({ S25935 }),
  .A3({ S25957[911] }),
  .ZN({ S250 })
);
AOI21_X1 #() 
AOI21_X1_2558_ (
  .A({ S25957[910] }),
  .B1({ S25950 }),
  .B2({ S25948 }),
  .ZN({ S251 })
);
AOI21_X1 #() 
AOI21_X1_2559_ (
  .A({ S25416 }),
  .B1({ S25755 }),
  .B2({ S240 }),
  .ZN({ S252 })
);
OAI21_X1 #() 
OAI21_X1_2370_ (
  .A({ S25957[909] }),
  .B1({ S252 }),
  .B2({ S244 }),
  .ZN({ S253 })
);
AOI21_X1 #() 
AOI21_X1_2560_ (
  .A({ S23551 }),
  .B1({ S253 }),
  .B2({ S236 }),
  .ZN({ S254 })
);
OAI21_X1 #() 
OAI21_X1_2371_ (
  .A({ S25568 }),
  .B1({ S254 }),
  .B2({ S251 }),
  .ZN({ S255 })
);
NAND3_X1 #() 
NAND3_X1_5004_ (
  .A1({ S255 }),
  .A2({ S25926 }),
  .A3({ S250 }),
  .ZN({ S256 })
);
AOI21_X1 #() 
AOI21_X1_2561_ (
  .A({ S25925 }),
  .B1({ S249 }),
  .B2({ S256 }),
  .ZN({ S257 })
);
AOI21_X1 #() 
AOI21_X1_2562_ (
  .A({ S25926 }),
  .B1({ S255 }),
  .B2({ S250 }),
  .ZN({ S258 })
);
AND3_X1 #() 
AND3_X1_182_ (
  .A1({ S255 }),
  .A2({ S250 }),
  .A3({ S25926 }),
  .ZN({ S259 })
);
NOR3_X1 #() 
NOR3_X1_155_ (
  .A1({ S259 }),
  .A2({ S258 }),
  .A3({ S25957[945] }),
  .ZN({ S260 })
);
OAI21_X1 #() 
OAI21_X1_2372_ (
  .A({ S25957[913] }),
  .B1({ S260 }),
  .B2({ S257 }),
  .ZN({ S261 })
);
NAND3_X1 #() 
NAND3_X1_5005_ (
  .A1({ S23241 }),
  .A2({ S23259 }),
  .A3({ S23263 }),
  .ZN({ S262 })
);
NAND3_X1 #() 
NAND3_X1_5006_ (
  .A1({ S23267 }),
  .A2({ S23270 }),
  .A3({ S25957[1041] }),
  .ZN({ S263 })
);
NAND2_X1 #() 
NAND2_X1_4597_ (
  .A1({ S262 }),
  .A2({ S263 }),
  .ZN({ S264 })
);
OAI21_X1 #() 
OAI21_X1_2373_ (
  .A({ S25957[945] }),
  .B1({ S259 }),
  .B2({ S258 }),
  .ZN({ S265 })
);
NAND3_X1 #() 
NAND3_X1_5007_ (
  .A1({ S249 }),
  .A2({ S25925 }),
  .A3({ S256 }),
  .ZN({ S266 })
);
NAND3_X1 #() 
NAND3_X1_5008_ (
  .A1({ S265 }),
  .A2({ S264 }),
  .A3({ S266 }),
  .ZN({ S267 })
);
NAND2_X1 #() 
NAND2_X1_4598_ (
  .A1({ S261 }),
  .A2({ S267 }),
  .ZN({ S25957[785] })
);
NOR2_X1 #() 
NOR2_X1_1160_ (
  .A1({ S20748 }),
  .A2({ S20751 }),
  .ZN({ S268 })
);
NAND2_X1 #() 
NAND2_X1_4599_ (
  .A1({ S20728 }),
  .A2({ S20747 }),
  .ZN({ S25957[1138] })
);
NAND2_X1 #() 
NAND2_X1_4600_ (
  .A1({ S23321 }),
  .A2({ S23294 }),
  .ZN({ S269 })
);
XNOR2_X1 #() 
XNOR2_X1_183_ (
  .A({ S269 }),
  .B({ S25957[1138] }),
  .ZN({ S25957[1010] })
);
INV_X1 #() 
INV_X1_1491_ (
  .A({ S25957[1010] }),
  .ZN({ S270 })
);
NAND3_X1 #() 
NAND3_X1_5009_ (
  .A1({ S25715 }),
  .A2({ S25450 }),
  .A3({ S25688 }),
  .ZN({ S271 })
);
OAI211_X1 #() 
OAI211_X1_1601_ (
  .A({ S25957[907] }),
  .B({ S25957[904] }),
  .C1({ S25957[906] }),
  .C2({ S25957[905] }),
  .ZN({ S272 })
);
OAI211_X1 #() 
OAI211_X1_1602_ (
  .A({ S25957[908] }),
  .B({ S272 }),
  .C1({ S25505 }),
  .C2({ S25504 }),
  .ZN({ S273 })
);
NAND3_X1 #() 
NAND3_X1_5010_ (
  .A1({ S273 }),
  .A2({ S271 }),
  .A3({ S25957[909] }),
  .ZN({ S274 })
);
AOI21_X1 #() 
AOI21_X1_2563_ (
  .A({ S25957[908] }),
  .B1({ S25443 }),
  .B2({ S25456 }),
  .ZN({ S275 })
);
NAND2_X1 #() 
NAND2_X1_4601_ (
  .A1({ S275 }),
  .A2({ S25842 }),
  .ZN({ S276 })
);
NAND3_X1 #() 
NAND3_X1_5011_ (
  .A1({ S25820 }),
  .A2({ S25957[908] }),
  .A3({ S25622 }),
  .ZN({ S277 })
);
NAND3_X1 #() 
NAND3_X1_5012_ (
  .A1({ S276 }),
  .A2({ S277 }),
  .A3({ S25484 }),
  .ZN({ S278 })
);
NAND2_X1 #() 
NAND2_X1_4602_ (
  .A1({ S274 }),
  .A2({ S278 }),
  .ZN({ S279 })
);
AOI21_X1 #() 
AOI21_X1_2564_ (
  .A({ S25416 }),
  .B1({ S25475 }),
  .B2({ S25442 }),
  .ZN({ S280 })
);
NAND2_X1 #() 
NAND2_X1_4603_ (
  .A1({ S25424 }),
  .A2({ S280 }),
  .ZN({ S281 })
);
NAND3_X1 #() 
NAND3_X1_5013_ (
  .A1({ S25438 }),
  .A2({ S25957[907] }),
  .A3({ S25642 }),
  .ZN({ S282 })
);
AOI21_X1 #() 
AOI21_X1_2565_ (
  .A({ S25484 }),
  .B1({ S282 }),
  .B2({ S25633 }),
  .ZN({ S283 })
);
NAND2_X1 #() 
NAND2_X1_4604_ (
  .A1({ S283 }),
  .A2({ S281 }),
  .ZN({ S284 })
);
NAND2_X1 #() 
NAND2_X1_4605_ (
  .A1({ S25583 }),
  .A2({ S25549 }),
  .ZN({ S285 })
);
OAI22_X1 #() 
OAI22_X1_119_ (
  .A1({ S285 }),
  .A2({ S25680 }),
  .B1({ S25595 }),
  .B2({ S25657 }),
  .ZN({ S286 })
);
AOI21_X1 #() 
AOI21_X1_2566_ (
  .A({ S25957[909] }),
  .B1({ S25707 }),
  .B2({ S25849 }),
  .ZN({ S287 })
);
NAND2_X1 #() 
NAND2_X1_4606_ (
  .A1({ S287 }),
  .A2({ S286 }),
  .ZN({ S288 })
);
NAND3_X1 #() 
NAND3_X1_5014_ (
  .A1({ S284 }),
  .A2({ S25957[910] }),
  .A3({ S288 }),
  .ZN({ S289 })
);
OAI211_X1 #() 
OAI211_X1_1603_ (
  .A({ S289 }),
  .B({ S25957[911] }),
  .C1({ S25957[910] }),
  .C2({ S279 }),
  .ZN({ S290 })
);
NAND3_X1 #() 
NAND3_X1_5015_ (
  .A1({ S25509 }),
  .A2({ S25871 }),
  .A3({ S25957[907] }),
  .ZN({ S291 })
);
NAND2_X1 #() 
NAND2_X1_4607_ (
  .A1({ S291 }),
  .A2({ S275 }),
  .ZN({ S292 })
);
NAND2_X1 #() 
NAND2_X1_4608_ (
  .A1({ S25694 }),
  .A2({ S25457 }),
  .ZN({ S293 })
);
NAND3_X1 #() 
NAND3_X1_5016_ (
  .A1({ S25784 }),
  .A2({ S293 }),
  .A3({ S25957[908] }),
  .ZN({ S294 })
);
AOI21_X1 #() 
AOI21_X1_2567_ (
  .A({ S25957[910] }),
  .B1({ S294 }),
  .B2({ S292 }),
  .ZN({ S295 })
);
AOI21_X1 #() 
AOI21_X1_2568_ (
  .A({ S25957[908] }),
  .B1({ S25548 }),
  .B2({ S25486 }),
  .ZN({ S296 })
);
NAND2_X1 #() 
NAND2_X1_4609_ (
  .A1({ S25439 }),
  .A2({ S296 }),
  .ZN({ S297 })
);
OAI211_X1 #() 
OAI211_X1_1604_ (
  .A({ S25422 }),
  .B({ S25957[907] }),
  .C1({ S25957[906] }),
  .C2({ S25957[905] }),
  .ZN({ S298 })
);
NAND2_X1 #() 
NAND2_X1_4610_ (
  .A1({ S25766 }),
  .A2({ S298 }),
  .ZN({ S299 })
);
AOI21_X1 #() 
AOI21_X1_2569_ (
  .A({ S23551 }),
  .B1({ S299 }),
  .B2({ S25957[908] }),
  .ZN({ S300 })
);
AND2_X1 #() 
AND2_X1_288_ (
  .A1({ S300 }),
  .A2({ S297 }),
  .ZN({ S301 })
);
OAI21_X1 #() 
OAI21_X1_2374_ (
  .A({ S25957[909] }),
  .B1({ S301 }),
  .B2({ S295 }),
  .ZN({ S302 })
);
AOI21_X1 #() 
AOI21_X1_2570_ (
  .A({ S25957[908] }),
  .B1({ S25576 }),
  .B2({ S25957[907] }),
  .ZN({ S303 })
);
NAND2_X1 #() 
NAND2_X1_4611_ (
  .A1({ S25682 }),
  .A2({ S303 }),
  .ZN({ S304 })
);
AOI21_X1 #() 
AOI21_X1_2571_ (
  .A({ S25408 }),
  .B1({ S25570 }),
  .B2({ S25463 }),
  .ZN({ S305 })
);
NAND2_X1 #() 
NAND2_X1_4612_ (
  .A1({ S25694 }),
  .A2({ S25610 }),
  .ZN({ S306 })
);
OAI211_X1 #() 
OAI211_X1_1605_ (
  .A({ S306 }),
  .B({ S25957[908] }),
  .C1({ S305 }),
  .C2({ S25957[907] }),
  .ZN({ S307 })
);
AOI21_X1 #() 
AOI21_X1_2572_ (
  .A({ S23551 }),
  .B1({ S304 }),
  .B2({ S307 }),
  .ZN({ S308 })
);
AOI21_X1 #() 
AOI21_X1_2573_ (
  .A({ S25416 }),
  .B1({ S25693 }),
  .B2({ S25622 }),
  .ZN({ S309 })
);
NAND4_X1 #() 
NAND4_X1_542_ (
  .A1({ S25438 }),
  .A2({ S25417 }),
  .A3({ S89 }),
  .A4({ S25416 }),
  .ZN({ S310 })
);
NAND3_X1 #() 
NAND3_X1_5017_ (
  .A1({ S25588 }),
  .A2({ S23551 }),
  .A3({ S310 }),
  .ZN({ S311 })
);
NOR2_X1 #() 
NOR2_X1_1161_ (
  .A1({ S311 }),
  .A2({ S309 }),
  .ZN({ S312 })
);
OAI21_X1 #() 
OAI21_X1_2375_ (
  .A({ S25484 }),
  .B1({ S312 }),
  .B2({ S308 }),
  .ZN({ S313 })
);
NAND3_X1 #() 
NAND3_X1_5018_ (
  .A1({ S313 }),
  .A2({ S302 }),
  .A3({ S25568 }),
  .ZN({ S314 })
);
NAND3_X1 #() 
NAND3_X1_5019_ (
  .A1({ S314 }),
  .A2({ S290 }),
  .A3({ S270 }),
  .ZN({ S315 })
);
AOI22_X1 #() 
AOI22_X1_525_ (
  .A1({ S283 }),
  .A2({ S281 }),
  .B1({ S287 }),
  .B2({ S286 }),
  .ZN({ S316 })
);
NAND2_X1 #() 
NAND2_X1_4613_ (
  .A1({ S279 }),
  .A2({ S23551 }),
  .ZN({ S317 })
);
OAI211_X1 #() 
OAI211_X1_1606_ (
  .A({ S317 }),
  .B({ S25957[911] }),
  .C1({ S23551 }),
  .C2({ S316 }),
  .ZN({ S318 })
);
NAND2_X1 #() 
NAND2_X1_4614_ (
  .A1({ S299 }),
  .A2({ S25957[908] }),
  .ZN({ S319 })
);
AOI21_X1 #() 
AOI21_X1_2574_ (
  .A({ S25484 }),
  .B1({ S297 }),
  .B2({ S319 }),
  .ZN({ S320 })
);
AOI21_X1 #() 
AOI21_X1_2575_ (
  .A({ S25957[907] }),
  .B1({ S25509 }),
  .B2({ S25549 }),
  .ZN({ S321 })
);
NOR2_X1 #() 
NOR2_X1_1162_ (
  .A1({ S25421 }),
  .A2({ S25957[906] }),
  .ZN({ S322 })
);
OAI21_X1 #() 
OAI21_X1_2376_ (
  .A({ S25957[908] }),
  .B1({ S322 }),
  .B2({ S25511 }),
  .ZN({ S323 })
);
NOR2_X1 #() 
NOR2_X1_1163_ (
  .A1({ S323 }),
  .A2({ S321 }),
  .ZN({ S324 })
);
AOI21_X1 #() 
AOI21_X1_2576_ (
  .A({ S25957[907] }),
  .B1({ S25689 }),
  .B2({ S25549 }),
  .ZN({ S325 })
);
AOI22_X1 #() 
AOI22_X1_526_ (
  .A1({ S25436 }),
  .A2({ S25957[904] }),
  .B1({ S23922 }),
  .B2({ S23925 }),
  .ZN({ S326 })
);
OAI21_X1 #() 
OAI21_X1_2377_ (
  .A({ S25416 }),
  .B1({ S326 }),
  .B2({ S89 }),
  .ZN({ S327 })
);
OAI21_X1 #() 
OAI21_X1_2378_ (
  .A({ S25484 }),
  .B1({ S325 }),
  .B2({ S327 }),
  .ZN({ S328 })
);
NOR2_X1 #() 
NOR2_X1_1164_ (
  .A1({ S328 }),
  .A2({ S324 }),
  .ZN({ S329 })
);
OAI21_X1 #() 
OAI21_X1_2379_ (
  .A({ S25957[910] }),
  .B1({ S329 }),
  .B2({ S320 }),
  .ZN({ S330 })
);
INV_X1 #() 
INV_X1_1492_ (
  .A({ S25622 }),
  .ZN({ S331 })
);
AOI21_X1 #() 
AOI21_X1_2577_ (
  .A({ S25957[907] }),
  .B1({ S25538 }),
  .B2({ S25442 }),
  .ZN({ S332 })
);
OAI21_X1 #() 
OAI21_X1_2380_ (
  .A({ S25957[908] }),
  .B1({ S332 }),
  .B2({ S331 }),
  .ZN({ S333 })
);
NAND4_X1 #() 
NAND4_X1_543_ (
  .A1({ S333 }),
  .A2({ S310 }),
  .A3({ S25484 }),
  .A4({ S25588 }),
  .ZN({ S334 })
);
NAND2_X1 #() 
NAND2_X1_4615_ (
  .A1({ S294 }),
  .A2({ S292 }),
  .ZN({ S335 })
);
NAND2_X1 #() 
NAND2_X1_4616_ (
  .A1({ S335 }),
  .A2({ S25957[909] }),
  .ZN({ S336 })
);
NAND3_X1 #() 
NAND3_X1_5020_ (
  .A1({ S336 }),
  .A2({ S334 }),
  .A3({ S23551 }),
  .ZN({ S337 })
);
NAND3_X1 #() 
NAND3_X1_5021_ (
  .A1({ S330 }),
  .A2({ S337 }),
  .A3({ S25568 }),
  .ZN({ S338 })
);
NAND3_X1 #() 
NAND3_X1_5022_ (
  .A1({ S338 }),
  .A2({ S25957[1010] }),
  .A3({ S318 }),
  .ZN({ S339 })
);
AOI21_X1 #() 
AOI21_X1_2578_ (
  .A({ S268 }),
  .B1({ S315 }),
  .B2({ S339 }),
  .ZN({ S340 })
);
INV_X1 #() 
INV_X1_1493_ (
  .A({ S268 }),
  .ZN({ S25957[1074] })
);
NAND3_X1 #() 
NAND3_X1_5023_ (
  .A1({ S314 }),
  .A2({ S290 }),
  .A3({ S25957[1010] }),
  .ZN({ S341 })
);
NAND3_X1 #() 
NAND3_X1_5024_ (
  .A1({ S338 }),
  .A2({ S270 }),
  .A3({ S318 }),
  .ZN({ S342 })
);
AOI21_X1 #() 
AOI21_X1_2579_ (
  .A({ S25957[1074] }),
  .B1({ S341 }),
  .B2({ S342 }),
  .ZN({ S343 })
);
OAI21_X1 #() 
OAI21_X1_2381_ (
  .A({ S25957[914] }),
  .B1({ S340 }),
  .B2({ S343 }),
  .ZN({ S344 })
);
AOI21_X1 #() 
AOI21_X1_2580_ (
  .A({ S23272 }),
  .B1({ S23336 }),
  .B2({ S23351 }),
  .ZN({ S345 })
);
AOI21_X1 #() 
AOI21_X1_2581_ (
  .A({ S25957[1234] }),
  .B1({ S23321 }),
  .B2({ S23294 }),
  .ZN({ S346 })
);
OAI21_X1 #() 
OAI21_X1_2382_ (
  .A({ S20682 }),
  .B1({ S345 }),
  .B2({ S346 }),
  .ZN({ S347 })
);
NAND3_X1 #() 
NAND3_X1_5025_ (
  .A1({ S23352 }),
  .A2({ S23322 }),
  .A3({ S25957[1170] }),
  .ZN({ S348 })
);
NAND2_X1 #() 
NAND2_X1_4617_ (
  .A1({ S347 }),
  .A2({ S348 }),
  .ZN({ S349 })
);
NAND3_X1 #() 
NAND3_X1_5026_ (
  .A1({ S341 }),
  .A2({ S342 }),
  .A3({ S25957[1074] }),
  .ZN({ S350 })
);
NAND3_X1 #() 
NAND3_X1_5027_ (
  .A1({ S315 }),
  .A2({ S339 }),
  .A3({ S268 }),
  .ZN({ S351 })
);
NAND3_X1 #() 
NAND3_X1_5028_ (
  .A1({ S350 }),
  .A2({ S351 }),
  .A3({ S349 }),
  .ZN({ S352 })
);
NAND2_X1 #() 
NAND2_X1_4618_ (
  .A1({ S344 }),
  .A2({ S352 }),
  .ZN({ S25957[786] })
);
AOI22_X1 #() 
AOI22_X1_527_ (
  .A1({ S24545 }),
  .A2({ S24558 }),
  .B1({ S24638 }),
  .B2({ S24635 }),
  .ZN({ S99 })
);
NAND4_X1 #() 
NAND4_X1_544_ (
  .A1({ S24545 }),
  .A2({ S24558 }),
  .A3({ S24635 }),
  .A4({ S24638 }),
  .ZN({ S100 })
);
INV_X1 #() 
INV_X1_1494_ (
  .A({ S25957[902] }),
  .ZN({ S353 })
);
INV_X1 #() 
INV_X1_1495_ (
  .A({ S25957[901] }),
  .ZN({ S354 })
);
AOI21_X1 #() 
AOI21_X1_2582_ (
  .A({ S19534 }),
  .B1({ S24719 }),
  .B2({ S24697 }),
  .ZN({ S355 })
);
AOI21_X1 #() 
AOI21_X1_2583_ (
  .A({ S25957[1218] }),
  .B1({ S24682 }),
  .B2({ S24660 }),
  .ZN({ S356 })
);
OAI21_X1 #() 
OAI21_X1_2383_ (
  .A({ S20775 }),
  .B1({ S355 }),
  .B2({ S356 }),
  .ZN({ S357 })
);
NAND3_X1 #() 
NAND3_X1_5029_ (
  .A1({ S24720 }),
  .A2({ S25957[1154] }),
  .A3({ S24683 }),
  .ZN({ S358 })
);
NAND2_X1 #() 
NAND2_X1_4619_ (
  .A1({ S357 }),
  .A2({ S358 }),
  .ZN({ S359 })
);
NAND3_X1 #() 
NAND3_X1_5030_ (
  .A1({ S24545 }),
  .A2({ S24558 }),
  .A3({ S359 }),
  .ZN({ S360 })
);
NAND2_X1 #() 
NAND2_X1_4620_ (
  .A1({ S360 }),
  .A2({ S25957[897] }),
  .ZN({ S361 })
);
AOI21_X1 #() 
AOI21_X1_2584_ (
  .A({ S359 }),
  .B1({ S24545 }),
  .B2({ S24558 }),
  .ZN({ S362 })
);
NAND2_X1 #() 
NAND2_X1_4621_ (
  .A1({ S362 }),
  .A2({ S25957[899] }),
  .ZN({ S363 })
);
NAND2_X1 #() 
NAND2_X1_4622_ (
  .A1({ S25957[897] }),
  .A2({ S359 }),
  .ZN({ S364 })
);
NAND2_X1 #() 
NAND2_X1_4623_ (
  .A1({ S364 }),
  .A2({ S360 }),
  .ZN({ S365 })
);
NAND2_X1 #() 
NAND2_X1_4624_ (
  .A1({ S365 }),
  .A2({ S25957[899] }),
  .ZN({ S366 })
);
OAI211_X1 #() 
OAI211_X1_1607_ (
  .A({ S366 }),
  .B({ S363 }),
  .C1({ S361 }),
  .C2({ S25957[899] }),
  .ZN({ S367 })
);
AOI21_X1 #() 
AOI21_X1_2585_ (
  .A({ S23360 }),
  .B1({ S24557 }),
  .B2({ S24553 }),
  .ZN({ S368 })
);
AND3_X1 #() 
AND3_X1_183_ (
  .A1({ S24557 }),
  .A2({ S24553 }),
  .A3({ S23360 }),
  .ZN({ S369 })
);
OAI21_X1 #() 
OAI21_X1_2384_ (
  .A({ S25957[897] }),
  .B1({ S369 }),
  .B2({ S368 }),
  .ZN({ S370 })
);
NAND2_X1 #() 
NAND2_X1_4625_ (
  .A1({ S370 }),
  .A2({ S100 }),
  .ZN({ S371 })
);
NAND2_X1 #() 
NAND2_X1_4626_ (
  .A1({ S360 }),
  .A2({ S25957[899] }),
  .ZN({ S372 })
);
OAI211_X1 #() 
OAI211_X1_1608_ (
  .A({ S24635 }),
  .B({ S24638 }),
  .C1({ S369 }),
  .C2({ S368 }),
  .ZN({ S373 })
);
AOI22_X1 #() 
AOI22_X1_528_ (
  .A1({ S25957[897] }),
  .A2({ S25957[898] }),
  .B1({ S24453 }),
  .B2({ S24444 }),
  .ZN({ S374 })
);
NAND3_X1 #() 
NAND3_X1_5031_ (
  .A1({ S374 }),
  .A2({ S373 }),
  .A3({ S360 }),
  .ZN({ S375 })
);
OAI21_X1 #() 
OAI21_X1_2385_ (
  .A({ S375 }),
  .B1({ S371 }),
  .B2({ S372 }),
  .ZN({ S376 })
);
MUX2_X1 #() 
MUX2_X1_17_ (
  .A({ S376 }),
  .B({ S367 }),
  .S({ S25957[900] }),
  .Z({ S377 })
);
AOI21_X1 #() 
AOI21_X1_2586_ (
  .A({ S25957[898] }),
  .B1({ S24638 }),
  .B2({ S24635 }),
  .ZN({ S378 })
);
NOR2_X1 #() 
NOR2_X1_1165_ (
  .A1({ S378 }),
  .A2({ S92 }),
  .ZN({ S379 })
);
INV_X1 #() 
INV_X1_1496_ (
  .A({ S379 }),
  .ZN({ S380 })
);
NAND3_X1 #() 
NAND3_X1_5032_ (
  .A1({ S25957[898] }),
  .A2({ S24635 }),
  .A3({ S24638 }),
  .ZN({ S381 })
);
NOR2_X1 #() 
NOR2_X1_1166_ (
  .A1({ S25957[896] }),
  .A2({ S381 }),
  .ZN({ S382 })
);
OAI21_X1 #() 
OAI21_X1_2386_ (
  .A({ S359 }),
  .B1({ S369 }),
  .B2({ S368 }),
  .ZN({ S383 })
);
NAND2_X1 #() 
NAND2_X1_4627_ (
  .A1({ S383 }),
  .A2({ S364 }),
  .ZN({ S384 })
);
OAI21_X1 #() 
OAI21_X1_2387_ (
  .A({ S92 }),
  .B1({ S25957[896] }),
  .B2({ S381 }),
  .ZN({ S385 })
);
OAI22_X1 #() 
OAI22_X1_120_ (
  .A1({ S380 }),
  .A2({ S382 }),
  .B1({ S385 }),
  .B2({ S384 }),
  .ZN({ S386 })
);
NAND3_X1 #() 
NAND3_X1_5033_ (
  .A1({ S25957[897] }),
  .A2({ S24545 }),
  .A3({ S24558 }),
  .ZN({ S387 })
);
INV_X1 #() 
INV_X1_1497_ (
  .A({ S387 }),
  .ZN({ S388 })
);
NOR2_X1 #() 
NOR2_X1_1167_ (
  .A1({ S388 }),
  .A2({ S25957[899] }),
  .ZN({ S389 })
);
NAND3_X1 #() 
NAND3_X1_5034_ (
  .A1({ S24635 }),
  .A2({ S24638 }),
  .A3({ S359 }),
  .ZN({ S390 })
);
AOI21_X1 #() 
AOI21_X1_2587_ (
  .A({ S92 }),
  .B1({ S387 }),
  .B2({ S390 }),
  .ZN({ S391 })
);
OAI21_X1 #() 
OAI21_X1_2388_ (
  .A({ S25957[900] }),
  .B1({ S389 }),
  .B2({ S391 }),
  .ZN({ S392 })
);
OAI211_X1 #() 
OAI211_X1_1609_ (
  .A({ S392 }),
  .B({ S354 }),
  .C1({ S25957[900] }),
  .C2({ S386 }),
  .ZN({ S393 })
);
OAI21_X1 #() 
OAI21_X1_2389_ (
  .A({ S393 }),
  .B1({ S377 }),
  .B2({ S354 }),
  .ZN({ S394 })
);
NAND3_X1 #() 
NAND3_X1_5035_ (
  .A1({ S24352 }),
  .A2({ S25957[1028] }),
  .A3({ S24351 }),
  .ZN({ S395 })
);
NAND3_X1 #() 
NAND3_X1_5036_ (
  .A1({ S24357 }),
  .A2({ S24359 }),
  .A3({ S23396 }),
  .ZN({ S396 })
);
NAND2_X1 #() 
NAND2_X1_4628_ (
  .A1({ S395 }),
  .A2({ S396 }),
  .ZN({ S397 })
);
NAND2_X1 #() 
NAND2_X1_4629_ (
  .A1({ S25957[897] }),
  .A2({ S25957[898] }),
  .ZN({ S398 })
);
NAND3_X1 #() 
NAND3_X1_5037_ (
  .A1({ S373 }),
  .A2({ S387 }),
  .A3({ S359 }),
  .ZN({ S399 })
);
NAND3_X1 #() 
NAND3_X1_5038_ (
  .A1({ S370 }),
  .A2({ S100 }),
  .A3({ S25957[898] }),
  .ZN({ S400 })
);
AOI21_X1 #() 
AOI21_X1_2588_ (
  .A({ S92 }),
  .B1({ S399 }),
  .B2({ S400 }),
  .ZN({ S401 })
);
AOI21_X1 #() 
AOI21_X1_2589_ (
  .A({ S25957[898] }),
  .B1({ S24545 }),
  .B2({ S24558 }),
  .ZN({ S402 })
);
NOR2_X1 #() 
NOR2_X1_1168_ (
  .A1({ S402 }),
  .A2({ S25957[899] }),
  .ZN({ S403 })
);
AOI21_X1 #() 
AOI21_X1_2590_ (
  .A({ S401 }),
  .B1({ S398 }),
  .B2({ S403 }),
  .ZN({ S404 })
);
NAND3_X1 #() 
NAND3_X1_5039_ (
  .A1({ S24545 }),
  .A2({ S24558 }),
  .A3({ S25957[898] }),
  .ZN({ S405 })
);
NAND2_X1 #() 
NAND2_X1_4630_ (
  .A1({ S405 }),
  .A2({ S92 }),
  .ZN({ S406 })
);
AND3_X1 #() 
AND3_X1_184_ (
  .A1({ S24635 }),
  .A2({ S24638 }),
  .A3({ S359 }),
  .ZN({ S407 })
);
NAND2_X1 #() 
NAND2_X1_4631_ (
  .A1({ S407 }),
  .A2({ S25957[899] }),
  .ZN({ S408 })
);
NAND2_X1 #() 
NAND2_X1_4632_ (
  .A1({ S360 }),
  .A2({ S390 }),
  .ZN({ S409 })
);
NAND2_X1 #() 
NAND2_X1_4633_ (
  .A1({ S409 }),
  .A2({ S100 }),
  .ZN({ S410 })
);
NAND2_X1 #() 
NAND2_X1_4634_ (
  .A1({ S410 }),
  .A2({ S398 }),
  .ZN({ S411 })
);
OAI211_X1 #() 
OAI211_X1_1610_ (
  .A({ S397 }),
  .B({ S408 }),
  .C1({ S411 }),
  .C2({ S406 }),
  .ZN({ S412 })
);
OAI21_X1 #() 
OAI21_X1_2390_ (
  .A({ S412 }),
  .B1({ S404 }),
  .B2({ S397 }),
  .ZN({ S413 })
);
NAND2_X1 #() 
NAND2_X1_4635_ (
  .A1({ S92 }),
  .A2({ S25957[897] }),
  .ZN({ S414 })
);
NOR2_X1 #() 
NOR2_X1_1169_ (
  .A1({ S414 }),
  .A2({ S362 }),
  .ZN({ S415 })
);
NOR2_X1 #() 
NOR2_X1_1170_ (
  .A1({ S92 }),
  .A2({ S25957[897] }),
  .ZN({ S416 })
);
OAI21_X1 #() 
OAI21_X1_2391_ (
  .A({ S25957[898] }),
  .B1({ S369 }),
  .B2({ S368 }),
  .ZN({ S417 })
);
NOR2_X1 #() 
NOR2_X1_1171_ (
  .A1({ S417 }),
  .A2({ S92 }),
  .ZN({ S418 })
);
NOR2_X1 #() 
NOR2_X1_1172_ (
  .A1({ S418 }),
  .A2({ S416 }),
  .ZN({ S419 })
);
NAND2_X1 #() 
NAND2_X1_4636_ (
  .A1({ S419 }),
  .A2({ S25957[900] }),
  .ZN({ S420 })
);
OAI21_X1 #() 
OAI21_X1_2392_ (
  .A({ S92 }),
  .B1({ S25957[896] }),
  .B2({ S390 }),
  .ZN({ S421 })
);
NAND3_X1 #() 
NAND3_X1_5040_ (
  .A1({ S421 }),
  .A2({ S397 }),
  .A3({ S370 }),
  .ZN({ S422 })
);
OAI21_X1 #() 
OAI21_X1_2393_ (
  .A({ S422 }),
  .B1({ S420 }),
  .B2({ S415 }),
  .ZN({ S423 })
);
AOI21_X1 #() 
AOI21_X1_2591_ (
  .A({ S25957[902] }),
  .B1({ S423 }),
  .B2({ S25957[901] }),
  .ZN({ S424 })
);
OAI21_X1 #() 
OAI21_X1_2394_ (
  .A({ S424 }),
  .B1({ S413 }),
  .B2({ S25957[901] }),
  .ZN({ S425 })
);
OAI21_X1 #() 
OAI21_X1_2395_ (
  .A({ S425 }),
  .B1({ S394 }),
  .B2({ S353 }),
  .ZN({ S426 })
);
NAND2_X1 #() 
NAND2_X1_4637_ (
  .A1({ S426 }),
  .A2({ S25957[903] }),
  .ZN({ S427 })
);
NAND4_X1 #() 
NAND4_X1_545_ (
  .A1({ S364 }),
  .A2({ S405 }),
  .A3({ S360 }),
  .A4({ S381 }),
  .ZN({ S428 })
);
AOI21_X1 #() 
AOI21_X1_2592_ (
  .A({ S25957[900] }),
  .B1({ S428 }),
  .B2({ S92 }),
  .ZN({ S429 })
);
OAI21_X1 #() 
OAI21_X1_2396_ (
  .A({ S429 }),
  .B1({ S362 }),
  .B2({ S380 }),
  .ZN({ S430 })
);
NAND2_X1 #() 
NAND2_X1_4638_ (
  .A1({ S405 }),
  .A2({ S381 }),
  .ZN({ S431 })
);
INV_X1 #() 
INV_X1_1498_ (
  .A({ S431 }),
  .ZN({ S432 })
);
AOI21_X1 #() 
AOI21_X1_2593_ (
  .A({ S92 }),
  .B1({ S399 }),
  .B2({ S432 }),
  .ZN({ S433 })
);
INV_X1 #() 
INV_X1_1499_ (
  .A({ S360 }),
  .ZN({ S434 })
);
AOI21_X1 #() 
AOI21_X1_2594_ (
  .A({ S359 }),
  .B1({ S370 }),
  .B2({ S100 }),
  .ZN({ S435 })
);
OAI21_X1 #() 
OAI21_X1_2397_ (
  .A({ S92 }),
  .B1({ S435 }),
  .B2({ S434 }),
  .ZN({ S436 })
);
NAND2_X1 #() 
NAND2_X1_4639_ (
  .A1({ S436 }),
  .A2({ S25957[900] }),
  .ZN({ S437 })
);
OAI21_X1 #() 
OAI21_X1_2398_ (
  .A({ S430 }),
  .B1({ S437 }),
  .B2({ S433 }),
  .ZN({ S438 })
);
NAND3_X1 #() 
NAND3_X1_5041_ (
  .A1({ S370 }),
  .A2({ S25957[899] }),
  .A3({ S405 }),
  .ZN({ S439 })
);
INV_X1 #() 
INV_X1_1500_ (
  .A({ S439 }),
  .ZN({ S440 })
);
INV_X1 #() 
INV_X1_1501_ (
  .A({ S374 }),
  .ZN({ S441 })
);
NAND2_X1 #() 
NAND2_X1_4640_ (
  .A1({ S25957[896] }),
  .A2({ S92 }),
  .ZN({ S442 })
);
NAND2_X1 #() 
NAND2_X1_4641_ (
  .A1({ S441 }),
  .A2({ S442 }),
  .ZN({ S443 })
);
OAI21_X1 #() 
OAI21_X1_2399_ (
  .A({ S25957[900] }),
  .B1({ S398 }),
  .B2({ S92 }),
  .ZN({ S444 })
);
AOI211_X1 #() 
AOI211_X1_83_ (
  .A({ S444 }),
  .B({ S440 }),
  .C1({ S443 }),
  .C2({ S360 }),
  .ZN({ S445 })
);
NAND2_X1 #() 
NAND2_X1_4642_ (
  .A1({ S407 }),
  .A2({ S25957[896] }),
  .ZN({ S446 })
);
NAND3_X1 #() 
NAND3_X1_5042_ (
  .A1({ S446 }),
  .A2({ S25957[899] }),
  .A3({ S398 }),
  .ZN({ S447 })
);
NAND2_X1 #() 
NAND2_X1_4643_ (
  .A1({ S431 }),
  .A2({ S92 }),
  .ZN({ S448 })
);
AOI21_X1 #() 
AOI21_X1_2595_ (
  .A({ S25957[900] }),
  .B1({ S447 }),
  .B2({ S448 }),
  .ZN({ S449 })
);
OAI21_X1 #() 
OAI21_X1_2400_ (
  .A({ S25957[901] }),
  .B1({ S445 }),
  .B2({ S449 }),
  .ZN({ S450 })
);
OAI21_X1 #() 
OAI21_X1_2401_ (
  .A({ S450 }),
  .B1({ S25957[901] }),
  .B2({ S438 }),
  .ZN({ S451 })
);
NOR2_X1 #() 
NOR2_X1_1173_ (
  .A1({ S362 }),
  .A2({ S92 }),
  .ZN({ S452 })
);
NAND2_X1 #() 
NAND2_X1_4644_ (
  .A1({ S452 }),
  .A2({ S390 }),
  .ZN({ S453 })
);
AND2_X1 #() 
AND2_X1_289_ (
  .A1({ S453 }),
  .A2({ S442 }),
  .ZN({ S454 })
);
AOI21_X1 #() 
AOI21_X1_2596_ (
  .A({ S25957[900] }),
  .B1({ S379 }),
  .B2({ S373 }),
  .ZN({ S455 })
);
OAI21_X1 #() 
OAI21_X1_2402_ (
  .A({ S455 }),
  .B1({ S441 }),
  .B2({ S409 }),
  .ZN({ S456 })
);
OAI21_X1 #() 
OAI21_X1_2403_ (
  .A({ S456 }),
  .B1({ S454 }),
  .B2({ S397 }),
  .ZN({ S457 })
);
AOI21_X1 #() 
AOI21_X1_2597_ (
  .A({ S25957[899] }),
  .B1({ S378 }),
  .B2({ S25957[896] }),
  .ZN({ S458 })
);
NAND2_X1 #() 
NAND2_X1_4645_ (
  .A1({ S400 }),
  .A2({ S458 }),
  .ZN({ S459 })
);
NAND4_X1 #() 
NAND4_X1_546_ (
  .A1({ S25957[897] }),
  .A2({ S25957[898] }),
  .A3({ S24545 }),
  .A4({ S24558 }),
  .ZN({ S460 })
);
AOI21_X1 #() 
AOI21_X1_2598_ (
  .A({ S397 }),
  .B1({ S460 }),
  .B2({ S25957[899] }),
  .ZN({ S461 })
);
NAND2_X1 #() 
NAND2_X1_4646_ (
  .A1({ S435 }),
  .A2({ S92 }),
  .ZN({ S462 })
);
NOR2_X1 #() 
NOR2_X1_1174_ (
  .A1({ S92 }),
  .A2({ S359 }),
  .ZN({ S463 })
);
AOI21_X1 #() 
AOI21_X1_2599_ (
  .A({ S25957[900] }),
  .B1({ S463 }),
  .B2({ S370 }),
  .ZN({ S464 })
);
AOI22_X1 #() 
AOI22_X1_529_ (
  .A1({ S464 }),
  .A2({ S462 }),
  .B1({ S459 }),
  .B2({ S461 }),
  .ZN({ S465 })
);
MUX2_X1 #() 
MUX2_X1_18_ (
  .A({ S465 }),
  .B({ S457 }),
  .S({ S25957[901] }),
  .Z({ S466 })
);
AOI21_X1 #() 
AOI21_X1_2600_ (
  .A({ S25957[903] }),
  .B1({ S466 }),
  .B2({ S353 }),
  .ZN({ S467 })
);
OAI21_X1 #() 
OAI21_X1_2404_ (
  .A({ S467 }),
  .B1({ S353 }),
  .B2({ S451 }),
  .ZN({ S468 })
);
NAND2_X1 #() 
NAND2_X1_4647_ (
  .A1({ S468 }),
  .A2({ S427 }),
  .ZN({ S469 })
);
NOR2_X1 #() 
NOR2_X1_1175_ (
  .A1({ S469 }),
  .A2({ S20873 }),
  .ZN({ S470 })
);
NAND2_X1 #() 
NAND2_X1_4648_ (
  .A1({ S469 }),
  .A2({ S20873 }),
  .ZN({ S471 })
);
INV_X1 #() 
INV_X1_1502_ (
  .A({ S471 }),
  .ZN({ S472 })
);
NOR2_X1 #() 
NOR2_X1_1176_ (
  .A1({ S472 }),
  .A2({ S470 }),
  .ZN({ S25957[847] })
);
NAND2_X1 #() 
NAND2_X1_4649_ (
  .A1({ S25957[847] }),
  .A2({ S22726 }),
  .ZN({ S473 })
);
INV_X1 #() 
INV_X1_1503_ (
  .A({ S25957[847] }),
  .ZN({ S474 })
);
NAND2_X1 #() 
NAND2_X1_4650_ (
  .A1({ S474 }),
  .A2({ S25957[1039] }),
  .ZN({ S475 })
);
NAND2_X1 #() 
NAND2_X1_4651_ (
  .A1({ S475 }),
  .A2({ S473 }),
  .ZN({ S25957[783] })
);
XOR2_X1 #() 
XOR2_X1_77_ (
  .A({ S25957[974] }),
  .B({ S25957[1070] }),
  .Z({ S25957[942] })
);
INV_X1 #() 
INV_X1_1504_ (
  .A({ S25957[942] }),
  .ZN({ S476 })
);
XNOR2_X1 #() 
XNOR2_X1_184_ (
  .A({ S23545 }),
  .B({ S25957[1134] }),
  .ZN({ S25957[1006] })
);
NAND3_X1 #() 
NAND3_X1_5043_ (
  .A1({ S383 }),
  .A2({ S398 }),
  .A3({ S405 }),
  .ZN({ S477 })
);
NAND2_X1 #() 
NAND2_X1_4652_ (
  .A1({ S477 }),
  .A2({ S25957[899] }),
  .ZN({ S478 })
);
NAND2_X1 #() 
NAND2_X1_4653_ (
  .A1({ S400 }),
  .A2({ S92 }),
  .ZN({ S479 })
);
AOI21_X1 #() 
AOI21_X1_2601_ (
  .A({ S25957[900] }),
  .B1({ S479 }),
  .B2({ S478 }),
  .ZN({ S480 })
);
NAND2_X1 #() 
NAND2_X1_4654_ (
  .A1({ S407 }),
  .A2({ S92 }),
  .ZN({ S481 })
);
AND3_X1 #() 
AND3_X1_185_ (
  .A1({ S481 }),
  .A2({ S442 }),
  .A3({ S25957[900] }),
  .ZN({ S482 })
);
NAND2_X1 #() 
NAND2_X1_4655_ (
  .A1({ S482 }),
  .A2({ S380 }),
  .ZN({ S483 })
);
INV_X1 #() 
INV_X1_1505_ (
  .A({ S483 }),
  .ZN({ S484 })
);
OAI21_X1 #() 
OAI21_X1_2405_ (
  .A({ S354 }),
  .B1({ S484 }),
  .B2({ S480 }),
  .ZN({ S485 })
);
NAND4_X1 #() 
NAND4_X1_547_ (
  .A1({ S383 }),
  .A2({ S405 }),
  .A3({ S381 }),
  .A4({ S92 }),
  .ZN({ S486 })
);
NAND2_X1 #() 
NAND2_X1_4656_ (
  .A1({ S383 }),
  .A2({ S100 }),
  .ZN({ S487 })
);
OAI211_X1 #() 
OAI211_X1_1611_ (
  .A({ S486 }),
  .B({ S25957[900] }),
  .C1({ S92 }),
  .C2({ S487 }),
  .ZN({ S488 })
);
INV_X1 #() 
INV_X1_1506_ (
  .A({ S488 }),
  .ZN({ S489 })
);
INV_X1 #() 
INV_X1_1507_ (
  .A({ S25957[897] }),
  .ZN({ S490 })
);
NOR2_X1 #() 
NOR2_X1_1177_ (
  .A1({ S402 }),
  .A2({ S490 }),
  .ZN({ S491 })
);
INV_X1 #() 
INV_X1_1508_ (
  .A({ S491 }),
  .ZN({ S492 })
);
AOI21_X1 #() 
AOI21_X1_2602_ (
  .A({ S25957[900] }),
  .B1({ S492 }),
  .B2({ S363 }),
  .ZN({ S493 })
);
OAI21_X1 #() 
OAI21_X1_2406_ (
  .A({ S25957[901] }),
  .B1({ S489 }),
  .B2({ S493 }),
  .ZN({ S494 })
);
NAND3_X1 #() 
NAND3_X1_5044_ (
  .A1({ S485 }),
  .A2({ S25957[902] }),
  .A3({ S494 }),
  .ZN({ S495 })
);
NAND3_X1 #() 
NAND3_X1_5045_ (
  .A1({ S460 }),
  .A2({ S390 }),
  .A3({ S383 }),
  .ZN({ S496 })
);
AOI21_X1 #() 
AOI21_X1_2603_ (
  .A({ S25957[900] }),
  .B1({ S496 }),
  .B2({ S25957[899] }),
  .ZN({ S497 })
);
INV_X1 #() 
INV_X1_1509_ (
  .A({ S403 }),
  .ZN({ S498 })
);
NOR2_X1 #() 
NOR2_X1_1178_ (
  .A1({ S369 }),
  .A2({ S368 }),
  .ZN({ S499 })
);
AND3_X1 #() 
AND3_X1_186_ (
  .A1({ S25957[898] }),
  .A2({ S24638 }),
  .A3({ S24635 }),
  .ZN({ S500 })
);
NAND2_X1 #() 
NAND2_X1_4657_ (
  .A1({ S500 }),
  .A2({ S499 }),
  .ZN({ S501 })
);
NAND3_X1 #() 
NAND3_X1_5046_ (
  .A1({ S501 }),
  .A2({ S25957[899] }),
  .A3({ S370 }),
  .ZN({ S502 })
);
NAND3_X1 #() 
NAND3_X1_5047_ (
  .A1({ S502 }),
  .A2({ S498 }),
  .A3({ S25957[900] }),
  .ZN({ S503 })
);
NAND2_X1 #() 
NAND2_X1_4658_ (
  .A1({ S446 }),
  .A2({ S374 }),
  .ZN({ S504 })
);
OAI21_X1 #() 
OAI21_X1_2407_ (
  .A({ S504 }),
  .B1({ S380 }),
  .B2({ S500 }),
  .ZN({ S505 })
);
OAI21_X1 #() 
OAI21_X1_2408_ (
  .A({ S503 }),
  .B1({ S505 }),
  .B2({ S25957[900] }),
  .ZN({ S506 })
);
OAI21_X1 #() 
OAI21_X1_2409_ (
  .A({ S447 }),
  .B1({ S499 }),
  .B2({ S481 }),
  .ZN({ S507 })
);
OAI21_X1 #() 
OAI21_X1_2410_ (
  .A({ S354 }),
  .B1({ S507 }),
  .B2({ S397 }),
  .ZN({ S508 })
);
OAI221_X1 #() 
OAI221_X1_135_ (
  .A({ S353 }),
  .B1({ S506 }),
  .B2({ S354 }),
  .C1({ S508 }),
  .C2({ S497 }),
  .ZN({ S509 })
);
NAND2_X1 #() 
NAND2_X1_4659_ (
  .A1({ S509 }),
  .A2({ S495 }),
  .ZN({ S510 })
);
INV_X1 #() 
INV_X1_1510_ (
  .A({ S414 }),
  .ZN({ S511 })
);
OAI21_X1 #() 
OAI21_X1_2411_ (
  .A({ S397 }),
  .B1({ S391 }),
  .B2({ S511 }),
  .ZN({ S512 })
);
NAND3_X1 #() 
NAND3_X1_5048_ (
  .A1({ S416 }),
  .A2({ S405 }),
  .A3({ S383 }),
  .ZN({ S513 })
);
NAND2_X1 #() 
NAND2_X1_4660_ (
  .A1({ S100 }),
  .A2({ S92 }),
  .ZN({ S514 })
);
OAI211_X1 #() 
OAI211_X1_1612_ (
  .A({ S513 }),
  .B({ S25957[900] }),
  .C1({ S359 }),
  .C2({ S514 }),
  .ZN({ S515 })
);
NAND3_X1 #() 
NAND3_X1_5049_ (
  .A1({ S515 }),
  .A2({ S25957[901] }),
  .A3({ S512 }),
  .ZN({ S516 })
);
AOI21_X1 #() 
AOI21_X1_2604_ (
  .A({ S92 }),
  .B1({ S500 }),
  .B2({ S499 }),
  .ZN({ S517 })
);
AOI21_X1 #() 
AOI21_X1_2605_ (
  .A({ S517 }),
  .B1({ S428 }),
  .B2({ S92 }),
  .ZN({ S518 })
);
AOI21_X1 #() 
AOI21_X1_2606_ (
  .A({ S92 }),
  .B1({ S360 }),
  .B2({ S390 }),
  .ZN({ S519 })
);
NOR3_X1 #() 
NOR3_X1_156_ (
  .A1({ S518 }),
  .A2({ S519 }),
  .A3({ S25957[900] }),
  .ZN({ S520 })
);
INV_X1 #() 
INV_X1_1511_ (
  .A({ S406 }),
  .ZN({ S521 })
);
NAND2_X1 #() 
NAND2_X1_4661_ (
  .A1({ S399 }),
  .A2({ S521 }),
  .ZN({ S522 })
);
AOI21_X1 #() 
AOI21_X1_2607_ (
  .A({ S397 }),
  .B1({ S522 }),
  .B2({ S478 }),
  .ZN({ S523 })
);
OR2_X1 #() 
OR2_X1_63_ (
  .A1({ S523 }),
  .A2({ S25957[901] }),
  .ZN({ S524 })
);
OAI211_X1 #() 
OAI211_X1_1613_ (
  .A({ S25957[902] }),
  .B({ S516 }),
  .C1({ S524 }),
  .C2({ S520 }),
  .ZN({ S525 })
);
NAND4_X1 #() 
NAND4_X1_548_ (
  .A1({ S25957[897] }),
  .A2({ S359 }),
  .A3({ S24545 }),
  .A4({ S24558 }),
  .ZN({ S526 })
);
INV_X1 #() 
INV_X1_1512_ (
  .A({ S526 }),
  .ZN({ S527 })
);
AOI22_X1 #() 
AOI22_X1_530_ (
  .A1({ S527 }),
  .A2({ S92 }),
  .B1({ S463 }),
  .B2({ S25957[897] }),
  .ZN({ S528 })
);
AOI21_X1 #() 
AOI21_X1_2608_ (
  .A({ S397 }),
  .B1({ S528 }),
  .B2({ S462 }),
  .ZN({ S529 })
);
NAND2_X1 #() 
NAND2_X1_4662_ (
  .A1({ S526 }),
  .A2({ S25957[899] }),
  .ZN({ S530 })
);
OAI21_X1 #() 
OAI21_X1_2412_ (
  .A({ S397 }),
  .B1({ S530 }),
  .B2({ S500 }),
  .ZN({ S531 })
);
AOI21_X1 #() 
AOI21_X1_2609_ (
  .A({ S531 }),
  .B1({ S403 }),
  .B2({ S371 }),
  .ZN({ S532 })
);
OAI21_X1 #() 
OAI21_X1_2413_ (
  .A({ S25957[901] }),
  .B1({ S532 }),
  .B2({ S529 }),
  .ZN({ S533 })
);
AOI21_X1 #() 
AOI21_X1_2610_ (
  .A({ S92 }),
  .B1({ S460 }),
  .B2({ S383 }),
  .ZN({ S534 })
);
AOI21_X1 #() 
AOI21_X1_2611_ (
  .A({ S534 }),
  .B1({ S521 }),
  .B2({ S399 }),
  .ZN({ S535 })
);
NOR2_X1 #() 
NOR2_X1_1179_ (
  .A1({ S535 }),
  .A2({ S25957[900] }),
  .ZN({ S536 })
);
AOI21_X1 #() 
AOI21_X1_2612_ (
  .A({ S420 }),
  .B1({ S365 }),
  .B2({ S92 }),
  .ZN({ S537 })
);
OAI21_X1 #() 
OAI21_X1_2414_ (
  .A({ S354 }),
  .B1({ S537 }),
  .B2({ S536 }),
  .ZN({ S538 })
);
NAND2_X1 #() 
NAND2_X1_4663_ (
  .A1({ S538 }),
  .A2({ S533 }),
  .ZN({ S539 })
);
NAND2_X1 #() 
NAND2_X1_4664_ (
  .A1({ S539 }),
  .A2({ S353 }),
  .ZN({ S540 })
);
NAND2_X1 #() 
NAND2_X1_4665_ (
  .A1({ S540 }),
  .A2({ S525 }),
  .ZN({ S541 })
);
NAND2_X1 #() 
NAND2_X1_4666_ (
  .A1({ S541 }),
  .A2({ S25957[903] }),
  .ZN({ S542 })
);
OAI211_X1 #() 
OAI211_X1_1614_ (
  .A({ S542 }),
  .B({ S25957[1006] }),
  .C1({ S510 }),
  .C2({ S25957[903] }),
  .ZN({ S543 })
);
INV_X1 #() 
INV_X1_1513_ (
  .A({ S25957[1006] }),
  .ZN({ S544 })
);
NAND2_X1 #() 
NAND2_X1_4667_ (
  .A1({ S510 }),
  .A2({ S24137 }),
  .ZN({ S545 })
);
NAND3_X1 #() 
NAND3_X1_5050_ (
  .A1({ S540 }),
  .A2({ S25957[903] }),
  .A3({ S525 }),
  .ZN({ S546 })
);
NAND3_X1 #() 
NAND3_X1_5051_ (
  .A1({ S546 }),
  .A2({ S544 }),
  .A3({ S545 }),
  .ZN({ S547 })
);
NAND3_X1 #() 
NAND3_X1_5052_ (
  .A1({ S543 }),
  .A2({ S23548 }),
  .A3({ S547 }),
  .ZN({ S548 })
);
OAI211_X1 #() 
OAI211_X1_1615_ (
  .A({ S542 }),
  .B({ S544 }),
  .C1({ S510 }),
  .C2({ S25957[903] }),
  .ZN({ S549 })
);
NAND3_X1 #() 
NAND3_X1_5053_ (
  .A1({ S546 }),
  .A2({ S25957[1006] }),
  .A3({ S545 }),
  .ZN({ S550 })
);
NAND3_X1 #() 
NAND3_X1_5054_ (
  .A1({ S549 }),
  .A2({ S550 }),
  .A3({ S25957[974] }),
  .ZN({ S551 })
);
AOI21_X1 #() 
AOI21_X1_2613_ (
  .A({ S476 }),
  .B1({ S548 }),
  .B2({ S551 }),
  .ZN({ S552 })
);
INV_X1 #() 
INV_X1_1514_ (
  .A({ S552 }),
  .ZN({ S553 })
);
NAND3_X1 #() 
NAND3_X1_5055_ (
  .A1({ S548 }),
  .A2({ S551 }),
  .A3({ S476 }),
  .ZN({ S554 })
);
NAND3_X1 #() 
NAND3_X1_5056_ (
  .A1({ S553 }),
  .A2({ S554 }),
  .A3({ S23551 }),
  .ZN({ S555 })
);
AND3_X1 #() 
AND3_X1_187_ (
  .A1({ S551 }),
  .A2({ S548 }),
  .A3({ S476 }),
  .ZN({ S556 })
);
OAI21_X1 #() 
OAI21_X1_2415_ (
  .A({ S25957[910] }),
  .B1({ S556 }),
  .B2({ S552 }),
  .ZN({ S557 })
);
NAND2_X1 #() 
NAND2_X1_4668_ (
  .A1({ S555 }),
  .A2({ S557 }),
  .ZN({ S25957[782] })
);
XNOR2_X1 #() 
XNOR2_X1_185_ (
  .A({ S25957[1133] }),
  .B({ S25957[1229] }),
  .ZN({ S558 })
);
INV_X1 #() 
INV_X1_1515_ (
  .A({ S558 }),
  .ZN({ S25957[1101] })
);
NAND2_X1 #() 
NAND2_X1_4669_ (
  .A1({ S499 }),
  .A2({ S407 }),
  .ZN({ S559 })
);
AOI21_X1 #() 
AOI21_X1_2614_ (
  .A({ S92 }),
  .B1({ S400 }),
  .B2({ S559 }),
  .ZN({ S560 })
);
OAI21_X1 #() 
OAI21_X1_2416_ (
  .A({ S397 }),
  .B1({ S560 }),
  .B2({ S458 }),
  .ZN({ S561 })
);
NOR2_X1 #() 
NOR2_X1_1180_ (
  .A1({ S410 }),
  .A2({ S92 }),
  .ZN({ S562 })
);
AOI21_X1 #() 
AOI21_X1_2615_ (
  .A({ S397 }),
  .B1({ S403 }),
  .B2({ S490 }),
  .ZN({ S563 })
);
INV_X1 #() 
INV_X1_1516_ (
  .A({ S563 }),
  .ZN({ S564 })
);
OAI21_X1 #() 
OAI21_X1_2417_ (
  .A({ S561 }),
  .B1({ S562 }),
  .B2({ S564 }),
  .ZN({ S565 })
);
NAND2_X1 #() 
NAND2_X1_4670_ (
  .A1({ S99 }),
  .A2({ S92 }),
  .ZN({ S566 })
);
NAND2_X1 #() 
NAND2_X1_4671_ (
  .A1({ S360 }),
  .A2({ S92 }),
  .ZN({ S567 })
);
OAI21_X1 #() 
OAI21_X1_2418_ (
  .A({ S567 }),
  .B1({ S428 }),
  .B2({ S92 }),
  .ZN({ S568 })
);
NAND2_X1 #() 
NAND2_X1_4672_ (
  .A1({ S568 }),
  .A2({ S566 }),
  .ZN({ S569 })
);
NAND2_X1 #() 
NAND2_X1_4673_ (
  .A1({ S569 }),
  .A2({ S25957[900] }),
  .ZN({ S570 })
);
AOI21_X1 #() 
AOI21_X1_2616_ (
  .A({ S25957[899] }),
  .B1({ S370 }),
  .B2({ S381 }),
  .ZN({ S571 })
);
INV_X1 #() 
INV_X1_1517_ (
  .A({ S571 }),
  .ZN({ S572 })
);
NOR2_X1 #() 
NOR2_X1_1181_ (
  .A1({ S416 }),
  .A2({ S25957[900] }),
  .ZN({ S573 })
);
AOI21_X1 #() 
AOI21_X1_2617_ (
  .A({ S354 }),
  .B1({ S572 }),
  .B2({ S573 }),
  .ZN({ S574 })
);
AOI22_X1 #() 
AOI22_X1_531_ (
  .A1({ S565 }),
  .A2({ S354 }),
  .B1({ S570 }),
  .B2({ S574 }),
  .ZN({ S575 })
);
NAND3_X1 #() 
NAND3_X1_5057_ (
  .A1({ S387 }),
  .A2({ S364 }),
  .A3({ S360 }),
  .ZN({ S576 })
);
NOR2_X1 #() 
NOR2_X1_1182_ (
  .A1({ S576 }),
  .A2({ S25957[899] }),
  .ZN({ S577 })
);
NOR2_X1 #() 
NOR2_X1_1183_ (
  .A1({ S25957[896] }),
  .A2({ S92 }),
  .ZN({ S578 })
);
NAND2_X1 #() 
NAND2_X1_4674_ (
  .A1({ S578 }),
  .A2({ S390 }),
  .ZN({ S579 })
);
NAND2_X1 #() 
NAND2_X1_4675_ (
  .A1({ S579 }),
  .A2({ S25957[900] }),
  .ZN({ S580 })
);
NAND2_X1 #() 
NAND2_X1_4676_ (
  .A1({ S361 }),
  .A2({ S25957[899] }),
  .ZN({ S581 })
);
INV_X1 #() 
INV_X1_1518_ (
  .A({ S581 }),
  .ZN({ S582 })
);
NOR3_X1 #() 
NOR3_X1_157_ (
  .A1({ S582 }),
  .A2({ S511 }),
  .A3({ S362 }),
  .ZN({ S583 })
);
OAI221_X1 #() 
OAI221_X1_136_ (
  .A({ S25957[901] }),
  .B1({ S580 }),
  .B2({ S577 }),
  .C1({ S25957[900] }),
  .C2({ S583 }),
  .ZN({ S584 })
);
AOI21_X1 #() 
AOI21_X1_2618_ (
  .A({ S92 }),
  .B1({ S383 }),
  .B2({ S390 }),
  .ZN({ S585 })
);
NAND2_X1 #() 
NAND2_X1_4677_ (
  .A1({ S417 }),
  .A2({ S381 }),
  .ZN({ S586 })
);
OAI21_X1 #() 
OAI21_X1_2419_ (
  .A({ S25957[900] }),
  .B1({ S586 }),
  .B2({ S25957[899] }),
  .ZN({ S587 })
);
AND2_X1 #() 
AND2_X1_290_ (
  .A1({ S462 }),
  .A2({ S478 }),
  .ZN({ S588 })
);
OAI221_X1 #() 
OAI221_X1_137_ (
  .A({ S354 }),
  .B1({ S585 }),
  .B2({ S587 }),
  .C1({ S588 }),
  .C2({ S25957[900] }),
  .ZN({ S589 })
);
NAND3_X1 #() 
NAND3_X1_5058_ (
  .A1({ S584 }),
  .A2({ S589 }),
  .A3({ S25957[902] }),
  .ZN({ S590 })
);
OAI211_X1 #() 
OAI211_X1_1616_ (
  .A({ S590 }),
  .B({ S25957[903] }),
  .C1({ S25957[902] }),
  .C2({ S575 }),
  .ZN({ S591 })
);
NAND3_X1 #() 
NAND3_X1_5059_ (
  .A1({ S373 }),
  .A2({ S387 }),
  .A3({ S25957[898] }),
  .ZN({ S592 })
);
AOI21_X1 #() 
AOI21_X1_2619_ (
  .A({ S92 }),
  .B1({ S499 }),
  .B2({ S378 }),
  .ZN({ S593 })
);
NAND4_X1 #() 
NAND4_X1_549_ (
  .A1({ S364 }),
  .A2({ S360 }),
  .A3({ S92 }),
  .A4({ S381 }),
  .ZN({ S594 })
);
INV_X1 #() 
INV_X1_1519_ (
  .A({ S594 }),
  .ZN({ S595 })
);
AOI21_X1 #() 
AOI21_X1_2620_ (
  .A({ S595 }),
  .B1({ S593 }),
  .B2({ S592 }),
  .ZN({ S596 })
);
NAND2_X1 #() 
NAND2_X1_4678_ (
  .A1({ S403 }),
  .A2({ S387 }),
  .ZN({ S597 })
);
OAI211_X1 #() 
OAI211_X1_1617_ (
  .A({ S597 }),
  .B({ S397 }),
  .C1({ S92 }),
  .C2({ S25957[896] }),
  .ZN({ S598 })
);
OAI211_X1 #() 
OAI211_X1_1618_ (
  .A({ S25957[901] }),
  .B({ S598 }),
  .C1({ S596 }),
  .C2({ S397 }),
  .ZN({ S599 })
);
NAND4_X1 #() 
NAND4_X1_550_ (
  .A1({ S383 }),
  .A2({ S405 }),
  .A3({ S381 }),
  .A4({ S25957[899] }),
  .ZN({ S600 })
);
NAND2_X1 #() 
NAND2_X1_4679_ (
  .A1({ S526 }),
  .A2({ S92 }),
  .ZN({ S601 })
);
NAND2_X1 #() 
NAND2_X1_4680_ (
  .A1({ S600 }),
  .A2({ S601 }),
  .ZN({ S602 })
);
NAND2_X1 #() 
NAND2_X1_4681_ (
  .A1({ S602 }),
  .A2({ S397 }),
  .ZN({ S603 })
);
AOI21_X1 #() 
AOI21_X1_2621_ (
  .A({ S603 }),
  .B1({ S600 }),
  .B2({ S362 }),
  .ZN({ S604 })
);
INV_X1 #() 
INV_X1_1520_ (
  .A({ S366 }),
  .ZN({ S605 })
);
AOI21_X1 #() 
AOI21_X1_2622_ (
  .A({ S359 }),
  .B1({ S24638 }),
  .B2({ S24635 }),
  .ZN({ S606 })
);
NAND2_X1 #() 
NAND2_X1_4682_ (
  .A1({ S25957[896] }),
  .A2({ S606 }),
  .ZN({ S607 })
);
INV_X1 #() 
INV_X1_1521_ (
  .A({ S607 }),
  .ZN({ S608 })
);
NOR3_X1 #() 
NOR3_X1_158_ (
  .A1({ S608 }),
  .A2({ S409 }),
  .A3({ S25957[899] }),
  .ZN({ S609 })
);
NOR3_X1 #() 
NOR3_X1_159_ (
  .A1({ S609 }),
  .A2({ S605 }),
  .A3({ S397 }),
  .ZN({ S610 })
);
OAI21_X1 #() 
OAI21_X1_2420_ (
  .A({ S354 }),
  .B1({ S604 }),
  .B2({ S610 }),
  .ZN({ S611 })
);
AND2_X1 #() 
AND2_X1_291_ (
  .A1({ S611 }),
  .A2({ S599 }),
  .ZN({ S612 })
);
NAND2_X1 #() 
NAND2_X1_4683_ (
  .A1({ S490 }),
  .A2({ S25957[899] }),
  .ZN({ S613 })
);
NAND2_X1 #() 
NAND2_X1_4684_ (
  .A1({ S606 }),
  .A2({ S92 }),
  .ZN({ S614 })
);
NAND2_X1 #() 
NAND2_X1_4685_ (
  .A1({ S613 }),
  .A2({ S614 }),
  .ZN({ S615 })
);
NOR2_X1 #() 
NOR2_X1_1184_ (
  .A1({ S25957[900] }),
  .A2({ S499 }),
  .ZN({ S616 })
);
NAND2_X1 #() 
NAND2_X1_4686_ (
  .A1({ S373 }),
  .A2({ S359 }),
  .ZN({ S617 })
);
AOI21_X1 #() 
AOI21_X1_2623_ (
  .A({ S92 }),
  .B1({ S400 }),
  .B2({ S617 }),
  .ZN({ S618 })
);
OAI21_X1 #() 
OAI21_X1_2421_ (
  .A({ S92 }),
  .B1({ S382 }),
  .B2({ S99 }),
  .ZN({ S619 })
);
NAND2_X1 #() 
NAND2_X1_4687_ (
  .A1({ S619 }),
  .A2({ S25957[900] }),
  .ZN({ S620 })
);
NOR2_X1 #() 
NOR2_X1_1185_ (
  .A1({ S620 }),
  .A2({ S618 }),
  .ZN({ S621 })
);
AOI211_X1 #() 
AOI211_X1_84_ (
  .A({ S25957[901] }),
  .B({ S621 }),
  .C1({ S615 }),
  .C2({ S616 }),
  .ZN({ S622 })
);
INV_X1 #() 
INV_X1_1522_ (
  .A({ S519 }),
  .ZN({ S623 })
);
AOI21_X1 #() 
AOI21_X1_2624_ (
  .A({ S397 }),
  .B1({ S623 }),
  .B2({ S601 }),
  .ZN({ S624 })
);
NAND2_X1 #() 
NAND2_X1_4688_ (
  .A1({ S363 }),
  .A2({ S406 }),
  .ZN({ S625 })
);
AOI21_X1 #() 
AOI21_X1_2625_ (
  .A({ S624 }),
  .B1({ S493 }),
  .B2({ S625 }),
  .ZN({ S626 })
);
NAND2_X1 #() 
NAND2_X1_4689_ (
  .A1({ S626 }),
  .A2({ S25957[901] }),
  .ZN({ S627 })
);
NAND2_X1 #() 
NAND2_X1_4690_ (
  .A1({ S627 }),
  .A2({ S353 }),
  .ZN({ S628 })
);
OAI221_X1 #() 
OAI221_X1_138_ (
  .A({ S24137 }),
  .B1({ S622 }),
  .B2({ S628 }),
  .C1({ S612 }),
  .C2({ S353 }),
  .ZN({ S629 })
);
AND3_X1 #() 
AND3_X1_188_ (
  .A1({ S629 }),
  .A2({ S591 }),
  .A3({ S25957[1101] }),
  .ZN({ S630 })
);
AOI21_X1 #() 
AOI21_X1_2626_ (
  .A({ S25957[1101] }),
  .B1({ S629 }),
  .B2({ S591 }),
  .ZN({ S631 })
);
OAI21_X1 #() 
OAI21_X1_2422_ (
  .A({ S21015 }),
  .B1({ S630 }),
  .B2({ S631 }),
  .ZN({ S632 })
);
NOR2_X1 #() 
NOR2_X1_1186_ (
  .A1({ S630 }),
  .A2({ S631 }),
  .ZN({ S633 })
);
NAND2_X1 #() 
NAND2_X1_4691_ (
  .A1({ S633 }),
  .A2({ S25957[1037] }),
  .ZN({ S634 })
);
NAND2_X1 #() 
NAND2_X1_4692_ (
  .A1({ S634 }),
  .A2({ S632 }),
  .ZN({ S25957[781] })
);
NAND2_X1 #() 
NAND2_X1_4693_ (
  .A1({ S25410 }),
  .A2({ S25411 }),
  .ZN({ S25957[940] })
);
INV_X1 #() 
INV_X1_1523_ (
  .A({ S25957[1068] }),
  .ZN({ S635 })
);
INV_X1 #() 
INV_X1_1524_ (
  .A({ S25957[1004] }),
  .ZN({ S636 })
);
INV_X1 #() 
INV_X1_1525_ (
  .A({ S455 }),
  .ZN({ S637 })
);
NAND3_X1 #() 
NAND3_X1_5060_ (
  .A1({ S405 }),
  .A2({ S92 }),
  .A3({ S390 }),
  .ZN({ S638 })
);
INV_X1 #() 
INV_X1_1526_ (
  .A({ S638 }),
  .ZN({ S639 })
);
NOR2_X1 #() 
NOR2_X1_1187_ (
  .A1({ S637 }),
  .A2({ S639 }),
  .ZN({ S640 })
);
NAND3_X1 #() 
NAND3_X1_5061_ (
  .A1({ S366 }),
  .A2({ S25957[900] }),
  .A3({ S385 }),
  .ZN({ S641 })
);
NOR2_X1 #() 
NOR2_X1_1188_ (
  .A1({ S378 }),
  .A2({ S25957[899] }),
  .ZN({ S642 })
);
NAND2_X1 #() 
NAND2_X1_4694_ (
  .A1({ S642 }),
  .A2({ S499 }),
  .ZN({ S643 })
);
NAND2_X1 #() 
NAND2_X1_4695_ (
  .A1({ S453 }),
  .A2({ S643 }),
  .ZN({ S644 })
);
OAI21_X1 #() 
OAI21_X1_2423_ (
  .A({ S641 }),
  .B1({ S644 }),
  .B2({ S25957[900] }),
  .ZN({ S645 })
);
NOR2_X1 #() 
NOR2_X1_1189_ (
  .A1({ S571 }),
  .A2({ S397 }),
  .ZN({ S646 })
);
OAI21_X1 #() 
OAI21_X1_2424_ (
  .A({ S646 }),
  .B1({ S613 }),
  .B2({ S402 }),
  .ZN({ S647 })
);
NAND2_X1 #() 
NAND2_X1_4696_ (
  .A1({ S647 }),
  .A2({ S354 }),
  .ZN({ S648 })
);
OAI221_X1 #() 
OAI221_X1_139_ (
  .A({ S25957[902] }),
  .B1({ S645 }),
  .B2({ S354 }),
  .C1({ S648 }),
  .C2({ S640 }),
  .ZN({ S649 })
);
NAND2_X1 #() 
NAND2_X1_4697_ (
  .A1({ S416 }),
  .A2({ S417 }),
  .ZN({ S650 })
);
OAI211_X1 #() 
OAI211_X1_1619_ (
  .A({ S650 }),
  .B({ S397 }),
  .C1({ S601 }),
  .C2({ S586 }),
  .ZN({ S651 })
);
INV_X1 #() 
INV_X1_1527_ (
  .A({ S373 }),
  .ZN({ S652 })
);
NAND3_X1 #() 
NAND3_X1_5062_ (
  .A1({ S383 }),
  .A2({ S100 }),
  .A3({ S398 }),
  .ZN({ S653 })
);
NAND2_X1 #() 
NAND2_X1_4698_ (
  .A1({ S653 }),
  .A2({ S92 }),
  .ZN({ S654 })
);
OAI211_X1 #() 
OAI211_X1_1620_ (
  .A({ S654 }),
  .B({ S25957[900] }),
  .C1({ S652 }),
  .C2({ S530 }),
  .ZN({ S655 })
);
NAND2_X1 #() 
NAND2_X1_4699_ (
  .A1({ S405 }),
  .A2({ S390 }),
  .ZN({ S656 })
);
NAND3_X1 #() 
NAND3_X1_5063_ (
  .A1({ S656 }),
  .A2({ S25957[899] }),
  .A3({ S381 }),
  .ZN({ S657 })
);
NAND3_X1 #() 
NAND3_X1_5064_ (
  .A1({ S417 }),
  .A2({ S25957[897] }),
  .A3({ S360 }),
  .ZN({ S658 })
);
AOI21_X1 #() 
AOI21_X1_2627_ (
  .A({ S397 }),
  .B1({ S658 }),
  .B2({ S92 }),
  .ZN({ S659 })
);
AOI21_X1 #() 
AOI21_X1_2628_ (
  .A({ S25957[901] }),
  .B1({ S659 }),
  .B2({ S657 }),
  .ZN({ S660 })
);
AOI21_X1 #() 
AOI21_X1_2629_ (
  .A({ S25957[898] }),
  .B1({ S370 }),
  .B2({ S100 }),
  .ZN({ S661 })
);
OAI21_X1 #() 
OAI21_X1_2425_ (
  .A({ S92 }),
  .B1({ S661 }),
  .B2({ S431 }),
  .ZN({ S662 })
);
AOI21_X1 #() 
AOI21_X1_2630_ (
  .A({ S25957[900] }),
  .B1({ S576 }),
  .B2({ S25957[899] }),
  .ZN({ S663 })
);
AOI21_X1 #() 
AOI21_X1_2631_ (
  .A({ S354 }),
  .B1({ S662 }),
  .B2({ S663 }),
  .ZN({ S664 })
);
AOI22_X1 #() 
AOI22_X1_532_ (
  .A1({ S664 }),
  .A2({ S655 }),
  .B1({ S660 }),
  .B2({ S651 }),
  .ZN({ S665 })
);
NAND2_X1 #() 
NAND2_X1_4700_ (
  .A1({ S665 }),
  .A2({ S353 }),
  .ZN({ S666 })
);
NAND3_X1 #() 
NAND3_X1_5065_ (
  .A1({ S649 }),
  .A2({ S25957[903] }),
  .A3({ S666 }),
  .ZN({ S667 })
);
NAND2_X1 #() 
NAND2_X1_4701_ (
  .A1({ S452 }),
  .A2({ S100 }),
  .ZN({ S668 })
);
OAI21_X1 #() 
OAI21_X1_2426_ (
  .A({ S668 }),
  .B1({ S384 }),
  .B2({ S385 }),
  .ZN({ S669 })
);
NAND2_X1 #() 
NAND2_X1_4702_ (
  .A1({ S669 }),
  .A2({ S397 }),
  .ZN({ S670 })
);
NAND4_X1 #() 
NAND4_X1_551_ (
  .A1({ S417 }),
  .A2({ S364 }),
  .A3({ S360 }),
  .A4({ S25957[899] }),
  .ZN({ S671 })
);
AOI21_X1 #() 
AOI21_X1_2632_ (
  .A({ S25957[901] }),
  .B1({ S646 }),
  .B2({ S671 }),
  .ZN({ S672 })
);
INV_X1 #() 
INV_X1_1528_ (
  .A({ S447 }),
  .ZN({ S673 })
);
NAND2_X1 #() 
NAND2_X1_4703_ (
  .A1({ S566 }),
  .A2({ S397 }),
  .ZN({ S674 })
);
OAI22_X1 #() 
OAI22_X1_121_ (
  .A1({ S562 }),
  .A2({ S674 }),
  .B1({ S673 }),
  .B2({ S587 }),
  .ZN({ S675 })
);
AOI22_X1 #() 
AOI22_X1_533_ (
  .A1({ S675 }),
  .A2({ S25957[901] }),
  .B1({ S670 }),
  .B2({ S672 }),
  .ZN({ S676 })
);
NAND2_X1 #() 
NAND2_X1_4704_ (
  .A1({ S443 }),
  .A2({ S399 }),
  .ZN({ S677 })
);
AND2_X1 #() 
AND2_X1_292_ (
  .A1({ S600 }),
  .A2({ S397 }),
  .ZN({ S678 })
);
AND2_X1 #() 
AND2_X1_293_ (
  .A1({ S677 }),
  .A2({ S678 }),
  .ZN({ S679 })
);
AOI21_X1 #() 
AOI21_X1_2633_ (
  .A({ S397 }),
  .B1({ S129 }),
  .B2({ S359 }),
  .ZN({ S680 })
);
OR2_X1 #() 
OR2_X1_64_ (
  .A1({ S680 }),
  .A2({ S354 }),
  .ZN({ S681 })
);
NOR2_X1 #() 
NOR2_X1_1190_ (
  .A1({ S463 }),
  .A2({ S25957[900] }),
  .ZN({ S682 })
);
NAND2_X1 #() 
NAND2_X1_4705_ (
  .A1({ S378 }),
  .A2({ S25957[896] }),
  .ZN({ S683 })
);
NAND3_X1 #() 
NAND3_X1_5066_ (
  .A1({ S683 }),
  .A2({ S92 }),
  .A3({ S405 }),
  .ZN({ S684 })
);
NAND2_X1 #() 
NAND2_X1_4706_ (
  .A1({ S684 }),
  .A2({ S682 }),
  .ZN({ S685 })
);
OAI21_X1 #() 
OAI21_X1_2427_ (
  .A({ S92 }),
  .B1({ S382 }),
  .B2({ S378 }),
  .ZN({ S686 })
);
NAND3_X1 #() 
NAND3_X1_5067_ (
  .A1({ S419 }),
  .A2({ S25957[900] }),
  .A3({ S686 }),
  .ZN({ S687 })
);
NAND3_X1 #() 
NAND3_X1_5068_ (
  .A1({ S687 }),
  .A2({ S354 }),
  .A3({ S685 }),
  .ZN({ S688 })
);
OAI211_X1 #() 
OAI211_X1_1621_ (
  .A({ S688 }),
  .B({ S25957[902] }),
  .C1({ S679 }),
  .C2({ S681 }),
  .ZN({ S689 })
);
OAI211_X1 #() 
OAI211_X1_1622_ (
  .A({ S689 }),
  .B({ S24137 }),
  .C1({ S676 }),
  .C2({ S25957[902] }),
  .ZN({ S690 })
);
NAND3_X1 #() 
NAND3_X1_5069_ (
  .A1({ S667 }),
  .A2({ S690 }),
  .A3({ S636 }),
  .ZN({ S691 })
);
OAI21_X1 #() 
OAI21_X1_2428_ (
  .A({ S688 }),
  .B1({ S679 }),
  .B2({ S681 }),
  .ZN({ S692 })
);
NAND2_X1 #() 
NAND2_X1_4707_ (
  .A1({ S692 }),
  .A2({ S25957[902] }),
  .ZN({ S693 })
);
NAND2_X1 #() 
NAND2_X1_4708_ (
  .A1({ S670 }),
  .A2({ S672 }),
  .ZN({ S694 })
);
NAND2_X1 #() 
NAND2_X1_4709_ (
  .A1({ S675 }),
  .A2({ S25957[901] }),
  .ZN({ S695 })
);
NAND3_X1 #() 
NAND3_X1_5070_ (
  .A1({ S695 }),
  .A2({ S694 }),
  .A3({ S353 }),
  .ZN({ S696 })
);
NAND3_X1 #() 
NAND3_X1_5071_ (
  .A1({ S693 }),
  .A2({ S696 }),
  .A3({ S24137 }),
  .ZN({ S697 })
);
AOI21_X1 #() 
AOI21_X1_2634_ (
  .A({ S639 }),
  .B1({ S373 }),
  .B2({ S379 }),
  .ZN({ S698 })
);
NOR2_X1 #() 
NOR2_X1_1191_ (
  .A1({ S613 }),
  .A2({ S402 }),
  .ZN({ S699 })
);
OAI21_X1 #() 
OAI21_X1_2429_ (
  .A({ S25957[900] }),
  .B1({ S699 }),
  .B2({ S571 }),
  .ZN({ S700 })
);
OAI211_X1 #() 
OAI211_X1_1623_ (
  .A({ S354 }),
  .B({ S700 }),
  .C1({ S698 }),
  .C2({ S25957[900] }),
  .ZN({ S701 })
);
NAND2_X1 #() 
NAND2_X1_4710_ (
  .A1({ S645 }),
  .A2({ S25957[901] }),
  .ZN({ S702 })
);
NAND3_X1 #() 
NAND3_X1_5072_ (
  .A1({ S702 }),
  .A2({ S25957[902] }),
  .A3({ S701 }),
  .ZN({ S703 })
);
OAI211_X1 #() 
OAI211_X1_1624_ (
  .A({ S703 }),
  .B({ S25957[903] }),
  .C1({ S665 }),
  .C2({ S25957[902] }),
  .ZN({ S704 })
);
NAND3_X1 #() 
NAND3_X1_5073_ (
  .A1({ S697 }),
  .A2({ S704 }),
  .A3({ S25957[1004] }),
  .ZN({ S705 })
);
AOI21_X1 #() 
AOI21_X1_2635_ (
  .A({ S635 }),
  .B1({ S691 }),
  .B2({ S705 }),
  .ZN({ S706 })
);
NAND3_X1 #() 
NAND3_X1_5074_ (
  .A1({ S667 }),
  .A2({ S690 }),
  .A3({ S25957[1004] }),
  .ZN({ S707 })
);
NAND3_X1 #() 
NAND3_X1_5075_ (
  .A1({ S697 }),
  .A2({ S704 }),
  .A3({ S636 }),
  .ZN({ S708 })
);
AOI21_X1 #() 
AOI21_X1_2636_ (
  .A({ S25957[1068] }),
  .B1({ S707 }),
  .B2({ S708 }),
  .ZN({ S709 })
);
OAI21_X1 #() 
OAI21_X1_2430_ (
  .A({ S25957[908] }),
  .B1({ S706 }),
  .B2({ S709 }),
  .ZN({ S710 })
);
NAND2_X1 #() 
NAND2_X1_4711_ (
  .A1({ S691 }),
  .A2({ S705 }),
  .ZN({ S25957[876] })
);
NAND2_X1 #() 
NAND2_X1_4712_ (
  .A1({ S25957[876] }),
  .A2({ S25957[1068] }),
  .ZN({ S711 })
);
NAND3_X1 #() 
NAND3_X1_5076_ (
  .A1({ S691 }),
  .A2({ S705 }),
  .A3({ S635 }),
  .ZN({ S712 })
);
NAND3_X1 #() 
NAND3_X1_5077_ (
  .A1({ S711 }),
  .A2({ S712 }),
  .A3({ S25416 }),
  .ZN({ S713 })
);
NAND2_X1 #() 
NAND2_X1_4713_ (
  .A1({ S710 }),
  .A2({ S713 }),
  .ZN({ S25957[780] })
);
NOR2_X1 #() 
NOR2_X1_1192_ (
  .A1({ S23787 }),
  .A2({ S23788 }),
  .ZN({ S25957[1003] })
);
NAND2_X1 #() 
NAND2_X1_4714_ (
  .A1({ S410 }),
  .A2({ S517 }),
  .ZN({ S714 })
);
NAND2_X1 #() 
NAND2_X1_4715_ (
  .A1({ S477 }),
  .A2({ S92 }),
  .ZN({ S715 })
);
NAND3_X1 #() 
NAND3_X1_5078_ (
  .A1({ S714 }),
  .A2({ S25957[900] }),
  .A3({ S715 }),
  .ZN({ S716 })
);
NAND3_X1 #() 
NAND3_X1_5079_ (
  .A1({ S400 }),
  .A2({ S92 }),
  .A3({ S390 }),
  .ZN({ S717 })
);
NAND4_X1 #() 
NAND4_X1_552_ (
  .A1({ S383 }),
  .A2({ S405 }),
  .A3({ S25957[897] }),
  .A4({ S25957[899] }),
  .ZN({ S718 })
);
NAND3_X1 #() 
NAND3_X1_5080_ (
  .A1({ S717 }),
  .A2({ S397 }),
  .A3({ S718 }),
  .ZN({ S719 })
);
NAND3_X1 #() 
NAND3_X1_5081_ (
  .A1({ S716 }),
  .A2({ S719 }),
  .A3({ S25957[901] }),
  .ZN({ S720 })
);
NAND2_X1 #() 
NAND2_X1_4716_ (
  .A1({ S417 }),
  .A2({ S490 }),
  .ZN({ S721 })
);
NAND3_X1 #() 
NAND3_X1_5082_ (
  .A1({ S721 }),
  .A2({ S25957[899] }),
  .A3({ S607 }),
  .ZN({ S722 })
);
NAND2_X1 #() 
NAND2_X1_4717_ (
  .A1({ S487 }),
  .A2({ S92 }),
  .ZN({ S723 })
);
NAND3_X1 #() 
NAND3_X1_5083_ (
  .A1({ S722 }),
  .A2({ S397 }),
  .A3({ S723 }),
  .ZN({ S724 })
);
OAI21_X1 #() 
OAI21_X1_2431_ (
  .A({ S25957[900] }),
  .B1({ S661 }),
  .B2({ S92 }),
  .ZN({ S725 })
);
OAI211_X1 #() 
OAI211_X1_1625_ (
  .A({ S724 }),
  .B({ S354 }),
  .C1({ S639 }),
  .C2({ S725 }),
  .ZN({ S726 })
);
AOI21_X1 #() 
AOI21_X1_2637_ (
  .A({ S25957[902] }),
  .B1({ S720 }),
  .B2({ S726 }),
  .ZN({ S727 })
);
AOI21_X1 #() 
AOI21_X1_2638_ (
  .A({ S25957[899] }),
  .B1({ S400 }),
  .B2({ S617 }),
  .ZN({ S728 })
);
OAI21_X1 #() 
OAI21_X1_2432_ (
  .A({ S25957[900] }),
  .B1({ S728 }),
  .B2({ S582 }),
  .ZN({ S729 })
);
NAND3_X1 #() 
NAND3_X1_5084_ (
  .A1({ S682 }),
  .A2({ S100 }),
  .A3({ S383 }),
  .ZN({ S730 })
);
AOI21_X1 #() 
AOI21_X1_2639_ (
  .A({ S25957[901] }),
  .B1({ S729 }),
  .B2({ S730 }),
  .ZN({ S731 })
);
NAND3_X1 #() 
NAND3_X1_5085_ (
  .A1({ S460 }),
  .A2({ S373 }),
  .A3({ S92 }),
  .ZN({ S732 })
);
AOI21_X1 #() 
AOI21_X1_2640_ (
  .A({ S397 }),
  .B1({ S668 }),
  .B2({ S732 }),
  .ZN({ S733 })
);
INV_X1 #() 
INV_X1_1529_ (
  .A({ S371 }),
  .ZN({ S734 })
);
NAND4_X1 #() 
NAND4_X1_553_ (
  .A1({ S383 }),
  .A2({ S100 }),
  .A3({ S398 }),
  .A4({ S25957[899] }),
  .ZN({ S735 })
);
OAI211_X1 #() 
OAI211_X1_1626_ (
  .A({ S735 }),
  .B({ S397 }),
  .C1({ S734 }),
  .C2({ S406 }),
  .ZN({ S736 })
);
NAND2_X1 #() 
NAND2_X1_4718_ (
  .A1({ S736 }),
  .A2({ S25957[901] }),
  .ZN({ S737 })
);
OAI21_X1 #() 
OAI21_X1_2433_ (
  .A({ S25957[902] }),
  .B1({ S737 }),
  .B2({ S733 }),
  .ZN({ S738 })
);
OAI21_X1 #() 
OAI21_X1_2434_ (
  .A({ S25957[903] }),
  .B1({ S738 }),
  .B2({ S731 }),
  .ZN({ S739 })
);
NAND3_X1 #() 
NAND3_X1_5086_ (
  .A1({ S459 }),
  .A2({ S478 }),
  .A3({ S25957[900] }),
  .ZN({ S740 })
);
NAND2_X1 #() 
NAND2_X1_4719_ (
  .A1({ S642 }),
  .A2({ S373 }),
  .ZN({ S741 })
);
NAND2_X1 #() 
NAND2_X1_4720_ (
  .A1({ S578 }),
  .A2({ S398 }),
  .ZN({ S742 })
);
NAND3_X1 #() 
NAND3_X1_5087_ (
  .A1({ S741 }),
  .A2({ S742 }),
  .A3({ S397 }),
  .ZN({ S743 })
);
NAND3_X1 #() 
NAND3_X1_5088_ (
  .A1({ S740 }),
  .A2({ S25957[901] }),
  .A3({ S743 }),
  .ZN({ S744 })
);
OAI21_X1 #() 
OAI21_X1_2435_ (
  .A({ S92 }),
  .B1({ S499 }),
  .B2({ S407 }),
  .ZN({ S745 })
);
NOR2_X1 #() 
NOR2_X1_1193_ (
  .A1({ S745 }),
  .A2({ S397 }),
  .ZN({ S746 })
);
AOI21_X1 #() 
AOI21_X1_2641_ (
  .A({ S746 }),
  .B1({ S429 }),
  .B2({ S671 }),
  .ZN({ S747 })
);
OAI211_X1 #() 
OAI211_X1_1627_ (
  .A({ S744 }),
  .B({ S25957[902] }),
  .C1({ S25957[901] }),
  .C2({ S747 }),
  .ZN({ S748 })
);
OAI21_X1 #() 
OAI21_X1_2436_ (
  .A({ S616 }),
  .B1({ S642 }),
  .B2({ S500 }),
  .ZN({ S749 })
);
NAND2_X1 #() 
NAND2_X1_4721_ (
  .A1({ S501 }),
  .A2({ S25957[899] }),
  .ZN({ S750 })
);
OAI211_X1 #() 
OAI211_X1_1628_ (
  .A({ S750 }),
  .B({ S25957[900] }),
  .C1({ S435 }),
  .C2({ S25957[899] }),
  .ZN({ S751 })
);
NAND3_X1 #() 
NAND3_X1_5089_ (
  .A1({ S751 }),
  .A2({ S25957[901] }),
  .A3({ S749 }),
  .ZN({ S752 })
);
AOI21_X1 #() 
AOI21_X1_2642_ (
  .A({ S25957[899] }),
  .B1({ S592 }),
  .B2({ S360 }),
  .ZN({ S753 })
);
OAI211_X1 #() 
OAI211_X1_1629_ (
  .A({ S25957[899] }),
  .B({ S100 }),
  .C1({ S370 }),
  .C2({ S25957[898] }),
  .ZN({ S754 })
);
NAND3_X1 #() 
NAND3_X1_5090_ (
  .A1({ S754 }),
  .A2({ S25957[900] }),
  .A3({ S594 }),
  .ZN({ S755 })
);
NAND3_X1 #() 
NAND3_X1_5091_ (
  .A1({ S623 }),
  .A2({ S397 }),
  .A3({ S363 }),
  .ZN({ S756 })
);
OAI211_X1 #() 
OAI211_X1_1630_ (
  .A({ S354 }),
  .B({ S755 }),
  .C1({ S756 }),
  .C2({ S753 }),
  .ZN({ S757 })
);
NAND3_X1 #() 
NAND3_X1_5092_ (
  .A1({ S757 }),
  .A2({ S752 }),
  .A3({ S353 }),
  .ZN({ S758 })
);
NAND3_X1 #() 
NAND3_X1_5093_ (
  .A1({ S748 }),
  .A2({ S24137 }),
  .A3({ S758 }),
  .ZN({ S759 })
);
OAI211_X1 #() 
OAI211_X1_1631_ (
  .A({ S759 }),
  .B({ S25957[1003] }),
  .C1({ S739 }),
  .C2({ S727 }),
  .ZN({ S760 })
);
INV_X1 #() 
INV_X1_1530_ (
  .A({ S25957[1003] }),
  .ZN({ S761 })
);
AOI22_X1 #() 
AOI22_X1_534_ (
  .A1({ S458 }),
  .A2({ S400 }),
  .B1({ S477 }),
  .B2({ S25957[899] }),
  .ZN({ S762 })
);
NAND2_X1 #() 
NAND2_X1_4722_ (
  .A1({ S741 }),
  .A2({ S742 }),
  .ZN({ S763 })
);
NAND2_X1 #() 
NAND2_X1_4723_ (
  .A1({ S763 }),
  .A2({ S397 }),
  .ZN({ S764 })
);
OAI211_X1 #() 
OAI211_X1_1632_ (
  .A({ S764 }),
  .B({ S25957[901] }),
  .C1({ S397 }),
  .C2({ S762 }),
  .ZN({ S765 })
);
NAND2_X1 #() 
NAND2_X1_4724_ (
  .A1({ S429 }),
  .A2({ S671 }),
  .ZN({ S766 })
);
NOR2_X1 #() 
NOR2_X1_1194_ (
  .A1({ S746 }),
  .A2({ S25957[901] }),
  .ZN({ S767 })
);
NAND2_X1 #() 
NAND2_X1_4725_ (
  .A1({ S766 }),
  .A2({ S767 }),
  .ZN({ S768 })
);
NAND3_X1 #() 
NAND3_X1_5094_ (
  .A1({ S765 }),
  .A2({ S25957[902] }),
  .A3({ S768 }),
  .ZN({ S769 })
);
NAND2_X1 #() 
NAND2_X1_4726_ (
  .A1({ S757 }),
  .A2({ S752 }),
  .ZN({ S770 })
);
NAND2_X1 #() 
NAND2_X1_4727_ (
  .A1({ S770 }),
  .A2({ S353 }),
  .ZN({ S771 })
);
NAND3_X1 #() 
NAND3_X1_5095_ (
  .A1({ S771 }),
  .A2({ S769 }),
  .A3({ S24137 }),
  .ZN({ S772 })
);
NAND3_X1 #() 
NAND3_X1_5096_ (
  .A1({ S729 }),
  .A2({ S354 }),
  .A3({ S730 }),
  .ZN({ S773 })
);
AOI21_X1 #() 
AOI21_X1_2643_ (
  .A({ S406 }),
  .B1({ S100 }),
  .B2({ S370 }),
  .ZN({ S774 })
);
INV_X1 #() 
INV_X1_1531_ (
  .A({ S735 }),
  .ZN({ S775 })
);
OAI21_X1 #() 
OAI21_X1_2437_ (
  .A({ S397 }),
  .B1({ S774 }),
  .B2({ S775 }),
  .ZN({ S776 })
);
AOI21_X1 #() 
AOI21_X1_2644_ (
  .A({ S397 }),
  .B1({ S452 }),
  .B2({ S100 }),
  .ZN({ S777 })
);
AOI21_X1 #() 
AOI21_X1_2645_ (
  .A({ S354 }),
  .B1({ S777 }),
  .B2({ S732 }),
  .ZN({ S778 })
);
NAND2_X1 #() 
NAND2_X1_4728_ (
  .A1({ S778 }),
  .A2({ S776 }),
  .ZN({ S779 })
);
NAND3_X1 #() 
NAND3_X1_5097_ (
  .A1({ S773 }),
  .A2({ S25957[902] }),
  .A3({ S779 }),
  .ZN({ S780 })
);
NAND3_X1 #() 
NAND3_X1_5098_ (
  .A1({ S720 }),
  .A2({ S726 }),
  .A3({ S353 }),
  .ZN({ S781 })
);
NAND3_X1 #() 
NAND3_X1_5099_ (
  .A1({ S780 }),
  .A2({ S781 }),
  .A3({ S25957[903] }),
  .ZN({ S782 })
);
NAND3_X1 #() 
NAND3_X1_5100_ (
  .A1({ S772 }),
  .A2({ S782 }),
  .A3({ S761 }),
  .ZN({ S783 })
);
AOI21_X1 #() 
AOI21_X1_2646_ (
  .A({ S23717 }),
  .B1({ S783 }),
  .B2({ S760 }),
  .ZN({ S784 })
);
OAI211_X1 #() 
OAI211_X1_1633_ (
  .A({ S759 }),
  .B({ S761 }),
  .C1({ S739 }),
  .C2({ S727 }),
  .ZN({ S785 })
);
NAND3_X1 #() 
NAND3_X1_5101_ (
  .A1({ S772 }),
  .A2({ S782 }),
  .A3({ S25957[1003] }),
  .ZN({ S786 })
);
AOI21_X1 #() 
AOI21_X1_2647_ (
  .A({ S25957[1067] }),
  .B1({ S786 }),
  .B2({ S785 }),
  .ZN({ S787 })
);
OAI21_X1 #() 
OAI21_X1_2438_ (
  .A({ S25957[907] }),
  .B1({ S784 }),
  .B2({ S787 }),
  .ZN({ S788 })
);
NAND3_X1 #() 
NAND3_X1_5102_ (
  .A1({ S786 }),
  .A2({ S785 }),
  .A3({ S25957[1067] }),
  .ZN({ S789 })
);
NAND3_X1 #() 
NAND3_X1_5103_ (
  .A1({ S783 }),
  .A2({ S760 }),
  .A3({ S23717 }),
  .ZN({ S790 })
);
NAND3_X1 #() 
NAND3_X1_5104_ (
  .A1({ S789 }),
  .A2({ S790 }),
  .A3({ S89 }),
  .ZN({ S791 })
);
NAND2_X1 #() 
NAND2_X1_4729_ (
  .A1({ S788 }),
  .A2({ S791 }),
  .ZN({ S101 })
);
AOI21_X1 #() 
AOI21_X1_2648_ (
  .A({ S89 }),
  .B1({ S789 }),
  .B2({ S790 }),
  .ZN({ S792 })
);
AND3_X1 #() 
AND3_X1_189_ (
  .A1({ S790 }),
  .A2({ S789 }),
  .A3({ S89 }),
  .ZN({ S793 })
);
NOR2_X1 #() 
NOR2_X1_1195_ (
  .A1({ S793 }),
  .A2({ S792 }),
  .ZN({ S25957[779] })
);
NOR2_X1 #() 
NOR2_X1_1196_ (
  .A1({ S23872 }),
  .A2({ S23845 }),
  .ZN({ S25957[968] })
);
NAND2_X1 #() 
NAND2_X1_4730_ (
  .A1({ S21260 }),
  .A2({ S21259 }),
  .ZN({ S25957[1128] })
);
NAND2_X1 #() 
NAND2_X1_4731_ (
  .A1({ S23871 }),
  .A2({ S23857 }),
  .ZN({ S794 })
);
XNOR2_X1 #() 
XNOR2_X1_186_ (
  .A({ S794 }),
  .B({ S25957[1128] }),
  .ZN({ S25957[1000] })
);
AOI21_X1 #() 
AOI21_X1_2649_ (
  .A({ S25957[900] }),
  .B1({ S600 }),
  .B2({ S601 }),
  .ZN({ S795 })
);
NAND2_X1 #() 
NAND2_X1_4732_ (
  .A1({ S371 }),
  .A2({ S463 }),
  .ZN({ S796 })
);
NAND2_X1 #() 
NAND2_X1_4733_ (
  .A1({ S654 }),
  .A2({ S796 }),
  .ZN({ S797 })
);
AOI21_X1 #() 
AOI21_X1_2650_ (
  .A({ S795 }),
  .B1({ S797 }),
  .B2({ S25957[900] }),
  .ZN({ S798 })
);
NAND2_X1 #() 
NAND2_X1_4734_ (
  .A1({ S383 }),
  .A2({ S490 }),
  .ZN({ S799 })
);
NAND2_X1 #() 
NAND2_X1_4735_ (
  .A1({ S458 }),
  .A2({ S799 }),
  .ZN({ S800 })
);
NAND3_X1 #() 
NAND3_X1_5105_ (
  .A1({ S800 }),
  .A2({ S397 }),
  .A3({ S671 }),
  .ZN({ S801 })
);
NAND3_X1 #() 
NAND3_X1_5106_ (
  .A1({ S387 }),
  .A2({ S25957[899] }),
  .A3({ S25957[898] }),
  .ZN({ S802 })
);
OAI211_X1 #() 
OAI211_X1_1634_ (
  .A({ S802 }),
  .B({ S25957[900] }),
  .C1({ S384 }),
  .C2({ S385 }),
  .ZN({ S803 })
);
NAND3_X1 #() 
NAND3_X1_5107_ (
  .A1({ S801 }),
  .A2({ S25957[901] }),
  .A3({ S803 }),
  .ZN({ S804 })
);
OAI211_X1 #() 
OAI211_X1_1635_ (
  .A({ S25957[902] }),
  .B({ S804 }),
  .C1({ S798 }),
  .C2({ S25957[901] }),
  .ZN({ S805 })
);
NAND4_X1 #() 
NAND4_X1_554_ (
  .A1({ S417 }),
  .A2({ S100 }),
  .A3({ S92 }),
  .A4({ S360 }),
  .ZN({ S806 })
);
AOI21_X1 #() 
AOI21_X1_2651_ (
  .A({ S25957[900] }),
  .B1({ S742 }),
  .B2({ S806 }),
  .ZN({ S807 })
);
AOI21_X1 #() 
AOI21_X1_2652_ (
  .A({ S25957[899] }),
  .B1({ S499 }),
  .B2({ S490 }),
  .ZN({ S808 })
);
AOI21_X1 #() 
AOI21_X1_2653_ (
  .A({ S444 }),
  .B1({ S409 }),
  .B2({ S808 }),
  .ZN({ S809 })
);
OAI21_X1 #() 
OAI21_X1_2439_ (
  .A({ S354 }),
  .B1({ S807 }),
  .B2({ S809 }),
  .ZN({ S810 })
);
AOI22_X1 #() 
AOI22_X1_535_ (
  .A1({ S402 }),
  .A2({ S490 }),
  .B1({ S499 }),
  .B2({ S606 }),
  .ZN({ S811 })
);
OAI211_X1 #() 
OAI211_X1_1636_ (
  .A({ S750 }),
  .B({ S25957[900] }),
  .C1({ S811 }),
  .C2({ S25957[899] }),
  .ZN({ S812 })
);
NAND2_X1 #() 
NAND2_X1_4736_ (
  .A1({ S576 }),
  .A2({ S25957[899] }),
  .ZN({ S813 })
);
NAND3_X1 #() 
NAND3_X1_5108_ (
  .A1({ S813 }),
  .A2({ S397 }),
  .A3({ S385 }),
  .ZN({ S814 })
);
NAND3_X1 #() 
NAND3_X1_5109_ (
  .A1({ S814 }),
  .A2({ S812 }),
  .A3({ S25957[901] }),
  .ZN({ S815 })
);
NAND3_X1 #() 
NAND3_X1_5110_ (
  .A1({ S815 }),
  .A2({ S810 }),
  .A3({ S353 }),
  .ZN({ S816 })
);
NAND3_X1 #() 
NAND3_X1_5111_ (
  .A1({ S805 }),
  .A2({ S25957[903] }),
  .A3({ S816 }),
  .ZN({ S817 })
);
INV_X1 #() 
INV_X1_1532_ (
  .A({ S683 }),
  .ZN({ S818 })
);
AOI21_X1 #() 
AOI21_X1_2654_ (
  .A({ S359 }),
  .B1({ S373 }),
  .B2({ S387 }),
  .ZN({ S819 })
);
OAI21_X1 #() 
OAI21_X1_2440_ (
  .A({ S25957[899] }),
  .B1({ S819 }),
  .B2({ S818 }),
  .ZN({ S820 })
);
NAND4_X1 #() 
NAND4_X1_555_ (
  .A1({ S460 }),
  .A2({ S383 }),
  .A3({ S390 }),
  .A4({ S25957[899] }),
  .ZN({ S821 })
);
NAND2_X1 #() 
NAND2_X1_4737_ (
  .A1({ S434 }),
  .A2({ S92 }),
  .ZN({ S822 })
);
NAND2_X1 #() 
NAND2_X1_4738_ (
  .A1({ S821 }),
  .A2({ S822 }),
  .ZN({ S823 })
);
AOI22_X1 #() 
AOI22_X1_536_ (
  .A1({ S820 }),
  .A2({ S482 }),
  .B1({ S823 }),
  .B2({ S397 }),
  .ZN({ S824 })
);
NAND2_X1 #() 
NAND2_X1_4739_ (
  .A1({ S721 }),
  .A2({ S92 }),
  .ZN({ S825 })
);
NAND3_X1 #() 
NAND3_X1_5112_ (
  .A1({ S825 }),
  .A2({ S397 }),
  .A3({ S600 }),
  .ZN({ S826 })
);
OAI211_X1 #() 
OAI211_X1_1637_ (
  .A({ S25957[900] }),
  .B({ S381 }),
  .C1({ S92 }),
  .C2({ S25957[896] }),
  .ZN({ S827 })
);
OAI211_X1 #() 
OAI211_X1_1638_ (
  .A({ S826 }),
  .B({ S354 }),
  .C1({ S527 }),
  .C2({ S827 }),
  .ZN({ S828 })
);
OAI211_X1 #() 
OAI211_X1_1639_ (
  .A({ S828 }),
  .B({ S25957[902] }),
  .C1({ S824 }),
  .C2({ S354 }),
  .ZN({ S829 })
);
NAND3_X1 #() 
NAND3_X1_5113_ (
  .A1({ S619 }),
  .A2({ S397 }),
  .A3({ S513 }),
  .ZN({ S830 })
);
NAND2_X1 #() 
NAND2_X1_4740_ (
  .A1({ S777 }),
  .A2({ S597 }),
  .ZN({ S831 })
);
NAND3_X1 #() 
NAND3_X1_5114_ (
  .A1({ S831 }),
  .A2({ S830 }),
  .A3({ S25957[901] }),
  .ZN({ S832 })
);
AOI21_X1 #() 
AOI21_X1_2655_ (
  .A({ S25957[899] }),
  .B1({ S721 }),
  .B2({ S607 }),
  .ZN({ S833 })
);
NAND4_X1 #() 
NAND4_X1_556_ (
  .A1({ S374 }),
  .A2({ S360 }),
  .A3({ S364 }),
  .A4({ S417 }),
  .ZN({ S834 })
);
OAI211_X1 #() 
OAI211_X1_1640_ (
  .A({ S373 }),
  .B({ S25957[899] }),
  .C1({ S362 }),
  .C2({ S490 }),
  .ZN({ S835 })
);
NAND3_X1 #() 
NAND3_X1_5115_ (
  .A1({ S834 }),
  .A2({ S835 }),
  .A3({ S397 }),
  .ZN({ S836 })
);
OAI211_X1 #() 
OAI211_X1_1641_ (
  .A({ S836 }),
  .B({ S354 }),
  .C1({ S725 }),
  .C2({ S833 }),
  .ZN({ S837 })
);
NAND3_X1 #() 
NAND3_X1_5116_ (
  .A1({ S837 }),
  .A2({ S832 }),
  .A3({ S353 }),
  .ZN({ S838 })
);
NAND3_X1 #() 
NAND3_X1_5117_ (
  .A1({ S829 }),
  .A2({ S24137 }),
  .A3({ S838 }),
  .ZN({ S839 })
);
NAND3_X1 #() 
NAND3_X1_5118_ (
  .A1({ S839 }),
  .A2({ S817 }),
  .A3({ S25957[1000] }),
  .ZN({ S840 })
);
INV_X1 #() 
INV_X1_1533_ (
  .A({ S25957[1000] }),
  .ZN({ S841 })
);
AOI22_X1 #() 
AOI22_X1_537_ (
  .A1({ S431 }),
  .A2({ S100 }),
  .B1({ S25957[897] }),
  .B2({ S402 }),
  .ZN({ S842 })
);
OAI21_X1 #() 
OAI21_X1_2441_ (
  .A({ S482 }),
  .B1({ S842 }),
  .B2({ S92 }),
  .ZN({ S843 })
);
NAND2_X1 #() 
NAND2_X1_4741_ (
  .A1({ S823 }),
  .A2({ S397 }),
  .ZN({ S844 })
);
AOI21_X1 #() 
AOI21_X1_2656_ (
  .A({ S354 }),
  .B1({ S843 }),
  .B2({ S844 }),
  .ZN({ S845 })
);
OAI21_X1 #() 
OAI21_X1_2442_ (
  .A({ S354 }),
  .B1({ S827 }),
  .B2({ S527 }),
  .ZN({ S846 })
);
AOI21_X1 #() 
AOI21_X1_2657_ (
  .A({ S846 }),
  .B1({ S678 }),
  .B2({ S825 }),
  .ZN({ S847 })
);
OAI21_X1 #() 
OAI21_X1_2443_ (
  .A({ S25957[902] }),
  .B1({ S845 }),
  .B2({ S847 }),
  .ZN({ S848 })
);
NAND2_X1 #() 
NAND2_X1_4742_ (
  .A1({ S837 }),
  .A2({ S832 }),
  .ZN({ S849 })
);
NAND2_X1 #() 
NAND2_X1_4743_ (
  .A1({ S849 }),
  .A2({ S353 }),
  .ZN({ S850 })
);
NAND3_X1 #() 
NAND3_X1_5119_ (
  .A1({ S850 }),
  .A2({ S848 }),
  .A3({ S24137 }),
  .ZN({ S851 })
);
AOI22_X1 #() 
AOI22_X1_538_ (
  .A1({ S653 }),
  .A2({ S92 }),
  .B1({ S371 }),
  .B2({ S463 }),
  .ZN({ S852 })
);
OAI211_X1 #() 
OAI211_X1_1642_ (
  .A({ S603 }),
  .B({ S354 }),
  .C1({ S852 }),
  .C2({ S397 }),
  .ZN({ S853 })
);
NAND2_X1 #() 
NAND2_X1_4744_ (
  .A1({ S801 }),
  .A2({ S803 }),
  .ZN({ S854 })
);
NAND2_X1 #() 
NAND2_X1_4745_ (
  .A1({ S854 }),
  .A2({ S25957[901] }),
  .ZN({ S855 })
);
NAND3_X1 #() 
NAND3_X1_5120_ (
  .A1({ S855 }),
  .A2({ S853 }),
  .A3({ S25957[902] }),
  .ZN({ S856 })
);
NAND2_X1 #() 
NAND2_X1_4746_ (
  .A1({ S815 }),
  .A2({ S810 }),
  .ZN({ S857 })
);
NAND2_X1 #() 
NAND2_X1_4747_ (
  .A1({ S857 }),
  .A2({ S353 }),
  .ZN({ S858 })
);
NAND3_X1 #() 
NAND3_X1_5121_ (
  .A1({ S858 }),
  .A2({ S25957[903] }),
  .A3({ S856 }),
  .ZN({ S859 })
);
NAND3_X1 #() 
NAND3_X1_5122_ (
  .A1({ S851 }),
  .A2({ S859 }),
  .A3({ S841 }),
  .ZN({ S860 })
);
NAND3_X1 #() 
NAND3_X1_5123_ (
  .A1({ S860 }),
  .A2({ S25957[968] }),
  .A3({ S840 }),
  .ZN({ S861 })
);
INV_X1 #() 
INV_X1_1534_ (
  .A({ S25957[968] }),
  .ZN({ S862 })
);
NAND3_X1 #() 
NAND3_X1_5124_ (
  .A1({ S839 }),
  .A2({ S817 }),
  .A3({ S841 }),
  .ZN({ S863 })
);
NAND3_X1 #() 
NAND3_X1_5125_ (
  .A1({ S851 }),
  .A2({ S859 }),
  .A3({ S25957[1000] }),
  .ZN({ S864 })
);
NAND3_X1 #() 
NAND3_X1_5126_ (
  .A1({ S864 }),
  .A2({ S862 }),
  .A3({ S863 }),
  .ZN({ S865 })
);
NAND3_X1 #() 
NAND3_X1_5127_ (
  .A1({ S861 }),
  .A2({ S865 }),
  .A3({ S22633 }),
  .ZN({ S866 })
);
NAND3_X1 #() 
NAND3_X1_5128_ (
  .A1({ S860 }),
  .A2({ S862 }),
  .A3({ S840 }),
  .ZN({ S867 })
);
NAND3_X1 #() 
NAND3_X1_5129_ (
  .A1({ S864 }),
  .A2({ S25957[968] }),
  .A3({ S863 }),
  .ZN({ S868 })
);
NAND3_X1 #() 
NAND3_X1_5130_ (
  .A1({ S867 }),
  .A2({ S868 }),
  .A3({ S25957[1032] }),
  .ZN({ S869 })
);
NAND2_X1 #() 
NAND2_X1_4748_ (
  .A1({ S866 }),
  .A2({ S869 }),
  .ZN({ S25957[776] })
);
NOR2_X1 #() 
NOR2_X1_1197_ (
  .A1({ S23919 }),
  .A2({ S23920 }),
  .ZN({ S25957[969] })
);
INV_X1 #() 
INV_X1_1535_ (
  .A({ S25957[969] }),
  .ZN({ S870 })
);
NAND2_X1 #() 
NAND2_X1_4749_ (
  .A1({ S21311 }),
  .A2({ S21310 }),
  .ZN({ S25957[1129] })
);
XNOR2_X1 #() 
XNOR2_X1_187_ (
  .A({ S23915 }),
  .B({ S25957[1129] }),
  .ZN({ S25957[1001] })
);
INV_X1 #() 
INV_X1_1536_ (
  .A({ S25957[1001] }),
  .ZN({ S871 })
);
AOI21_X1 #() 
AOI21_X1_2658_ (
  .A({ S92 }),
  .B1({ S400 }),
  .B2({ S683 }),
  .ZN({ S872 })
);
NOR3_X1 #() 
NOR3_X1_160_ (
  .A1({ S872 }),
  .A2({ S443 }),
  .A3({ S25957[900] }),
  .ZN({ S873 })
);
NAND3_X1 #() 
NAND3_X1_5131_ (
  .A1({ S405 }),
  .A2({ S92 }),
  .A3({ S381 }),
  .ZN({ S874 })
);
NAND3_X1 #() 
NAND3_X1_5132_ (
  .A1({ S581 }),
  .A2({ S25957[900] }),
  .A3({ S874 }),
  .ZN({ S875 })
);
NAND2_X1 #() 
NAND2_X1_4750_ (
  .A1({ S875 }),
  .A2({ S25957[901] }),
  .ZN({ S876 })
);
NOR2_X1 #() 
NOR2_X1_1198_ (
  .A1({ S25957[896] }),
  .A2({ S390 }),
  .ZN({ S877 })
);
OAI211_X1 #() 
OAI211_X1_1643_ (
  .A({ S439 }),
  .B({ S397 }),
  .C1({ S745 }),
  .C2({ S877 }),
  .ZN({ S878 })
);
NAND2_X1 #() 
NAND2_X1_4751_ (
  .A1({ S374 }),
  .A2({ S499 }),
  .ZN({ S879 })
);
OAI211_X1 #() 
OAI211_X1_1644_ (
  .A({ S25957[900] }),
  .B({ S879 }),
  .C1({ S435 }),
  .C2({ S530 }),
  .ZN({ S880 })
);
NAND3_X1 #() 
NAND3_X1_5133_ (
  .A1({ S880 }),
  .A2({ S354 }),
  .A3({ S878 }),
  .ZN({ S881 })
);
OAI211_X1 #() 
OAI211_X1_1645_ (
  .A({ S881 }),
  .B({ S25957[902] }),
  .C1({ S873 }),
  .C2({ S876 }),
  .ZN({ S882 })
);
OAI21_X1 #() 
OAI21_X1_2444_ (
  .A({ S397 }),
  .B1({ S601 }),
  .B2({ S586 }),
  .ZN({ S883 })
);
NAND3_X1 #() 
NAND3_X1_5134_ (
  .A1({ S526 }),
  .A2({ S92 }),
  .A3({ S381 }),
  .ZN({ S884 })
);
AOI21_X1 #() 
AOI21_X1_2659_ (
  .A({ S397 }),
  .B1({ S25957[899] }),
  .B2({ S378 }),
  .ZN({ S885 })
);
AOI21_X1 #() 
AOI21_X1_2660_ (
  .A({ S25957[901] }),
  .B1({ S885 }),
  .B2({ S884 }),
  .ZN({ S886 })
);
OAI21_X1 #() 
OAI21_X1_2445_ (
  .A({ S886 }),
  .B1({ S433 }),
  .B2({ S883 }),
  .ZN({ S887 })
);
AOI21_X1 #() 
AOI21_X1_2661_ (
  .A({ S92 }),
  .B1({ S592 }),
  .B2({ S360 }),
  .ZN({ S888 })
);
INV_X1 #() 
INV_X1_1537_ (
  .A({ S460 }),
  .ZN({ S889 })
);
OAI21_X1 #() 
OAI21_X1_2446_ (
  .A({ S25957[900] }),
  .B1({ S889 }),
  .B2({ S567 }),
  .ZN({ S890 })
);
NAND3_X1 #() 
NAND3_X1_5135_ (
  .A1({ S383 }),
  .A2({ S25957[899] }),
  .A3({ S390 }),
  .ZN({ S891 })
);
NAND3_X1 #() 
NAND3_X1_5136_ (
  .A1({ S741 }),
  .A2({ S397 }),
  .A3({ S891 }),
  .ZN({ S892 })
);
OAI211_X1 #() 
OAI211_X1_1646_ (
  .A({ S892 }),
  .B({ S25957[901] }),
  .C1({ S888 }),
  .C2({ S890 }),
  .ZN({ S893 })
);
NAND3_X1 #() 
NAND3_X1_5137_ (
  .A1({ S893 }),
  .A2({ S887 }),
  .A3({ S353 }),
  .ZN({ S894 })
);
NAND3_X1 #() 
NAND3_X1_5138_ (
  .A1({ S882 }),
  .A2({ S25957[903] }),
  .A3({ S894 }),
  .ZN({ S895 })
);
NAND3_X1 #() 
NAND3_X1_5139_ (
  .A1({ S796 }),
  .A2({ S397 }),
  .A3({ S486 }),
  .ZN({ S896 })
);
OAI21_X1 #() 
OAI21_X1_2447_ (
  .A({ S25957[900] }),
  .B1({ S608 }),
  .B2({ S421 }),
  .ZN({ S897 })
);
OAI211_X1 #() 
OAI211_X1_1647_ (
  .A({ S896 }),
  .B({ S354 }),
  .C1({ S872 }),
  .C2({ S897 }),
  .ZN({ S898 })
);
NAND2_X1 #() 
NAND2_X1_4752_ (
  .A1({ S371 }),
  .A2({ S452 }),
  .ZN({ S899 })
);
OAI211_X1 #() 
OAI211_X1_1648_ (
  .A({ S899 }),
  .B({ S25957[900] }),
  .C1({ S382 }),
  .C2({ S498 }),
  .ZN({ S900 })
);
NAND3_X1 #() 
NAND3_X1_5140_ (
  .A1({ S573 }),
  .A2({ S417 }),
  .A3({ S559 }),
  .ZN({ S901 })
);
NAND3_X1 #() 
NAND3_X1_5141_ (
  .A1({ S900 }),
  .A2({ S25957[901] }),
  .A3({ S901 }),
  .ZN({ S902 })
);
NAND3_X1 #() 
NAND3_X1_5142_ (
  .A1({ S902 }),
  .A2({ S898 }),
  .A3({ S25957[902] }),
  .ZN({ S903 })
);
AOI21_X1 #() 
AOI21_X1_2662_ (
  .A({ S397 }),
  .B1({ S643 }),
  .B2({ S718 }),
  .ZN({ S904 })
);
OAI21_X1 #() 
OAI21_X1_2448_ (
  .A({ S25957[901] }),
  .B1({ S904 }),
  .B2({ S429 }),
  .ZN({ S905 })
);
NAND4_X1 #() 
NAND4_X1_557_ (
  .A1({ S638 }),
  .A2({ S363 }),
  .A3({ S613 }),
  .A4({ S25957[900] }),
  .ZN({ S906 })
);
OAI211_X1 #() 
OAI211_X1_1649_ (
  .A({ S397 }),
  .B({ S408 }),
  .C1({ S874 }),
  .C2({ S365 }),
  .ZN({ S907 })
);
NAND3_X1 #() 
NAND3_X1_5143_ (
  .A1({ S907 }),
  .A2({ S354 }),
  .A3({ S906 }),
  .ZN({ S908 })
);
NAND3_X1 #() 
NAND3_X1_5144_ (
  .A1({ S905 }),
  .A2({ S353 }),
  .A3({ S908 }),
  .ZN({ S909 })
);
NAND3_X1 #() 
NAND3_X1_5145_ (
  .A1({ S903 }),
  .A2({ S909 }),
  .A3({ S24137 }),
  .ZN({ S910 })
);
NAND3_X1 #() 
NAND3_X1_5146_ (
  .A1({ S910 }),
  .A2({ S895 }),
  .A3({ S871 }),
  .ZN({ S911 })
);
AOI22_X1 #() 
AOI22_X1_539_ (
  .A1({ S452 }),
  .A2({ S371 }),
  .B1({ S403 }),
  .B2({ S501 }),
  .ZN({ S912 })
);
AOI21_X1 #() 
AOI21_X1_2663_ (
  .A({ S25957[897] }),
  .B1({ S360 }),
  .B2({ S92 }),
  .ZN({ S913 })
);
OAI21_X1 #() 
OAI21_X1_2449_ (
  .A({ S397 }),
  .B1({ S913 }),
  .B2({ S362 }),
  .ZN({ S914 })
);
OAI211_X1 #() 
OAI211_X1_1650_ (
  .A({ S25957[901] }),
  .B({ S914 }),
  .C1({ S912 }),
  .C2({ S397 }),
  .ZN({ S915 })
);
AOI21_X1 #() 
AOI21_X1_2664_ (
  .A({ S25957[900] }),
  .B1({ S371 }),
  .B2({ S463 }),
  .ZN({ S916 })
);
AOI21_X1 #() 
AOI21_X1_2665_ (
  .A({ S25957[899] }),
  .B1({ S499 }),
  .B2({ S407 }),
  .ZN({ S917 })
);
AOI21_X1 #() 
AOI21_X1_2666_ (
  .A({ S397 }),
  .B1({ S917 }),
  .B2({ S607 }),
  .ZN({ S918 })
);
AOI22_X1 #() 
AOI22_X1_540_ (
  .A1({ S820 }),
  .A2({ S918 }),
  .B1({ S486 }),
  .B2({ S916 }),
  .ZN({ S919 })
);
OAI211_X1 #() 
OAI211_X1_1651_ (
  .A({ S915 }),
  .B({ S25957[902] }),
  .C1({ S919 }),
  .C2({ S25957[901] }),
  .ZN({ S920 })
);
NAND2_X1 #() 
NAND2_X1_4753_ (
  .A1({ S907 }),
  .A2({ S906 }),
  .ZN({ S921 })
);
NAND2_X1 #() 
NAND2_X1_4754_ (
  .A1({ S921 }),
  .A2({ S354 }),
  .ZN({ S922 })
);
INV_X1 #() 
INV_X1_1538_ (
  .A({ S429 }),
  .ZN({ S923 })
);
NAND2_X1 #() 
NAND2_X1_4755_ (
  .A1({ S923 }),
  .A2({ S25957[901] }),
  .ZN({ S924 })
);
OAI211_X1 #() 
OAI211_X1_1652_ (
  .A({ S922 }),
  .B({ S353 }),
  .C1({ S924 }),
  .C2({ S904 }),
  .ZN({ S925 })
);
NAND3_X1 #() 
NAND3_X1_5147_ (
  .A1({ S920 }),
  .A2({ S925 }),
  .A3({ S24137 }),
  .ZN({ S926 })
);
NAND3_X1 #() 
NAND3_X1_5148_ (
  .A1({ S581 }),
  .A2({ S25957[901] }),
  .A3({ S874 }),
  .ZN({ S927 })
);
AOI21_X1 #() 
AOI21_X1_2667_ (
  .A({ S25957[901] }),
  .B1({ S374 }),
  .B2({ S499 }),
  .ZN({ S928 })
);
OAI21_X1 #() 
OAI21_X1_2450_ (
  .A({ S928 }),
  .B1({ S435 }),
  .B2({ S530 }),
  .ZN({ S929 })
);
NAND2_X1 #() 
NAND2_X1_4756_ (
  .A1({ S929 }),
  .A2({ S927 }),
  .ZN({ S930 })
);
NAND2_X1 #() 
NAND2_X1_4757_ (
  .A1({ S930 }),
  .A2({ S25957[900] }),
  .ZN({ S931 })
);
NAND3_X1 #() 
NAND3_X1_5149_ (
  .A1({ S441 }),
  .A2({ S25957[901] }),
  .A3({ S442 }),
  .ZN({ S932 })
);
OAI211_X1 #() 
OAI211_X1_1653_ (
  .A({ S439 }),
  .B({ S354 }),
  .C1({ S745 }),
  .C2({ S877 }),
  .ZN({ S933 })
);
OAI21_X1 #() 
OAI21_X1_2451_ (
  .A({ S933 }),
  .B1({ S872 }),
  .B2({ S932 }),
  .ZN({ S934 })
);
NAND2_X1 #() 
NAND2_X1_4758_ (
  .A1({ S934 }),
  .A2({ S397 }),
  .ZN({ S935 })
);
NAND3_X1 #() 
NAND3_X1_5150_ (
  .A1({ S935 }),
  .A2({ S931 }),
  .A3({ S25957[902] }),
  .ZN({ S936 })
);
NAND2_X1 #() 
NAND2_X1_4759_ (
  .A1({ S893 }),
  .A2({ S887 }),
  .ZN({ S937 })
);
NAND2_X1 #() 
NAND2_X1_4760_ (
  .A1({ S937 }),
  .A2({ S353 }),
  .ZN({ S938 })
);
NAND3_X1 #() 
NAND3_X1_5151_ (
  .A1({ S938 }),
  .A2({ S936 }),
  .A3({ S25957[903] }),
  .ZN({ S939 })
);
NAND3_X1 #() 
NAND3_X1_5152_ (
  .A1({ S939 }),
  .A2({ S25957[1001] }),
  .A3({ S926 }),
  .ZN({ S940 })
);
NAND3_X1 #() 
NAND3_X1_5153_ (
  .A1({ S940 }),
  .A2({ S870 }),
  .A3({ S911 }),
  .ZN({ S941 })
);
NAND3_X1 #() 
NAND3_X1_5154_ (
  .A1({ S910 }),
  .A2({ S895 }),
  .A3({ S25957[1001] }),
  .ZN({ S942 })
);
NAND3_X1 #() 
NAND3_X1_5155_ (
  .A1({ S939 }),
  .A2({ S871 }),
  .A3({ S926 }),
  .ZN({ S943 })
);
NAND3_X1 #() 
NAND3_X1_5156_ (
  .A1({ S943 }),
  .A2({ S25957[969] }),
  .A3({ S942 }),
  .ZN({ S944 })
);
AOI21_X1 #() 
AOI21_X1_2668_ (
  .A({ S25957[1033] }),
  .B1({ S941 }),
  .B2({ S944 }),
  .ZN({ S945 })
);
AND3_X1 #() 
AND3_X1_190_ (
  .A1({ S944 }),
  .A2({ S941 }),
  .A3({ S25957[1033] }),
  .ZN({ S946 })
);
NOR2_X1 #() 
NOR2_X1_1199_ (
  .A1({ S946 }),
  .A2({ S945 }),
  .ZN({ S25957[777] })
);
NAND2_X1 #() 
NAND2_X1_4761_ (
  .A1({ S21384 }),
  .A2({ S21383 }),
  .ZN({ S25957[1130] })
);
NAND2_X1 #() 
NAND2_X1_4762_ (
  .A1({ S23950 }),
  .A2({ S23972 }),
  .ZN({ S947 })
);
XNOR2_X1 #() 
XNOR2_X1_188_ (
  .A({ S947 }),
  .B({ S25957[1130] }),
  .ZN({ S25957[1002] })
);
NAND4_X1 #() 
NAND4_X1_558_ (
  .A1({ S398 }),
  .A2({ S360 }),
  .A3({ S405 }),
  .A4({ S390 }),
  .ZN({ S948 })
);
AOI22_X1 #() 
AOI22_X1_541_ (
  .A1({ S948 }),
  .A2({ S92 }),
  .B1({ S593 }),
  .B2({ S417 }),
  .ZN({ S949 })
);
NAND3_X1 #() 
NAND3_X1_5157_ (
  .A1({ S383 }),
  .A2({ S25957[899] }),
  .A3({ S25957[897] }),
  .ZN({ S950 })
);
OAI211_X1 #() 
OAI211_X1_1654_ (
  .A({ S397 }),
  .B({ S950 }),
  .C1({ S441 }),
  .C2({ S487 }),
  .ZN({ S951 })
);
OAI211_X1 #() 
OAI211_X1_1655_ (
  .A({ S354 }),
  .B({ S951 }),
  .C1({ S949 }),
  .C2({ S397 }),
  .ZN({ S952 })
);
NAND2_X1 #() 
NAND2_X1_4763_ (
  .A1({ S364 }),
  .A2({ S92 }),
  .ZN({ S953 })
);
OAI21_X1 #() 
OAI21_X1_2452_ (
  .A({ S397 }),
  .B1({ S953 }),
  .B2({ S499 }),
  .ZN({ S954 })
);
AOI21_X1 #() 
AOI21_X1_2669_ (
  .A({ S25957[899] }),
  .B1({ S25957[896] }),
  .B2({ S390 }),
  .ZN({ S955 })
);
AOI21_X1 #() 
AOI21_X1_2670_ (
  .A({ S92 }),
  .B1({ S405 }),
  .B2({ S490 }),
  .ZN({ S956 })
);
OAI21_X1 #() 
OAI21_X1_2453_ (
  .A({ S25957[900] }),
  .B1({ S956 }),
  .B2({ S955 }),
  .ZN({ S957 })
);
OAI211_X1 #() 
OAI211_X1_1656_ (
  .A({ S25957[901] }),
  .B({ S957 }),
  .C1({ S401 }),
  .C2({ S954 }),
  .ZN({ S958 })
);
AND3_X1 #() 
AND3_X1_191_ (
  .A1({ S952 }),
  .A2({ S25957[902] }),
  .A3({ S958 }),
  .ZN({ S959 })
);
NAND2_X1 #() 
NAND2_X1_4764_ (
  .A1({ S496 }),
  .A2({ S25957[899] }),
  .ZN({ S960 })
);
NAND4_X1 #() 
NAND4_X1_559_ (
  .A1({ S446 }),
  .A2({ S526 }),
  .A3({ S92 }),
  .A4({ S398 }),
  .ZN({ S961 })
);
NAND3_X1 #() 
NAND3_X1_5158_ (
  .A1({ S960 }),
  .A2({ S397 }),
  .A3({ S961 }),
  .ZN({ S962 })
);
NAND2_X1 #() 
NAND2_X1_4765_ (
  .A1({ S658 }),
  .A2({ S92 }),
  .ZN({ S963 })
);
NAND3_X1 #() 
NAND3_X1_5159_ (
  .A1({ S963 }),
  .A2({ S25957[900] }),
  .A3({ S950 }),
  .ZN({ S964 })
);
NAND3_X1 #() 
NAND3_X1_5160_ (
  .A1({ S962 }),
  .A2({ S354 }),
  .A3({ S964 }),
  .ZN({ S965 })
);
NAND4_X1 #() 
NAND4_X1_560_ (
  .A1({ S607 }),
  .A2({ S360 }),
  .A3({ S390 }),
  .A4({ S25957[899] }),
  .ZN({ S966 })
);
OAI211_X1 #() 
OAI211_X1_1657_ (
  .A({ S966 }),
  .B({ S397 }),
  .C1({ S360 }),
  .C2({ S414 }),
  .ZN({ S967 })
);
NAND2_X1 #() 
NAND2_X1_4766_ (
  .A1({ S452 }),
  .A2({ S559 }),
  .ZN({ S968 })
);
NAND3_X1 #() 
NAND3_X1_5161_ (
  .A1({ S717 }),
  .A2({ S25957[900] }),
  .A3({ S968 }),
  .ZN({ S969 })
);
NAND3_X1 #() 
NAND3_X1_5162_ (
  .A1({ S969 }),
  .A2({ S25957[901] }),
  .A3({ S967 }),
  .ZN({ S970 })
);
AOI21_X1 #() 
AOI21_X1_2671_ (
  .A({ S25957[902] }),
  .B1({ S970 }),
  .B2({ S965 }),
  .ZN({ S971 })
);
OAI21_X1 #() 
OAI21_X1_2454_ (
  .A({ S24137 }),
  .B1({ S959 }),
  .B2({ S971 }),
  .ZN({ S972 })
);
NAND3_X1 #() 
NAND3_X1_5163_ (
  .A1({ S25957[896] }),
  .A2({ S25957[899] }),
  .A3({ S390 }),
  .ZN({ S973 })
);
OAI211_X1 #() 
OAI211_X1_1658_ (
  .A({ S25957[900] }),
  .B({ S973 }),
  .C1({ S874 }),
  .C2({ S365 }),
  .ZN({ S974 })
);
NAND2_X1 #() 
NAND2_X1_4767_ (
  .A1({ S374 }),
  .A2({ S417 }),
  .ZN({ S975 })
);
AOI21_X1 #() 
AOI21_X1_2672_ (
  .A({ S25957[900] }),
  .B1({ S99 }),
  .B2({ S25957[899] }),
  .ZN({ S976 })
);
NAND3_X1 #() 
NAND3_X1_5164_ (
  .A1({ S976 }),
  .A2({ S650 }),
  .A3({ S975 }),
  .ZN({ S977 })
);
NAND3_X1 #() 
NAND3_X1_5165_ (
  .A1({ S977 }),
  .A2({ S974 }),
  .A3({ S25957[901] }),
  .ZN({ S978 })
);
OAI221_X1 #() 
OAI221_X1_140_ (
  .A({ S397 }),
  .B1({ S398 }),
  .B2({ S92 }),
  .C1({ S414 }),
  .C2({ S360 }),
  .ZN({ S979 })
);
NAND3_X1 #() 
NAND3_X1_5166_ (
  .A1({ S950 }),
  .A2({ S25957[900] }),
  .A3({ S953 }),
  .ZN({ S980 })
);
NAND3_X1 #() 
NAND3_X1_5167_ (
  .A1({ S979 }),
  .A2({ S980 }),
  .A3({ S354 }),
  .ZN({ S981 })
);
NAND3_X1 #() 
NAND3_X1_5168_ (
  .A1({ S978 }),
  .A2({ S353 }),
  .A3({ S981 }),
  .ZN({ S982 })
);
NAND2_X1 #() 
NAND2_X1_4768_ (
  .A1({ S387 }),
  .A2({ S25957[898] }),
  .ZN({ S983 })
);
AOI21_X1 #() 
AOI21_X1_2673_ (
  .A({ S92 }),
  .B1({ S410 }),
  .B2({ S983 }),
  .ZN({ S984 })
);
NAND2_X1 #() 
NAND2_X1_4769_ (
  .A1({ S614 }),
  .A2({ S397 }),
  .ZN({ S985 })
);
AOI22_X1 #() 
AOI22_X1_542_ (
  .A1({ S458 }),
  .A2({ S799 }),
  .B1({ S656 }),
  .B2({ S25957[899] }),
  .ZN({ S986 })
);
OAI22_X1 #() 
OAI22_X1_122_ (
  .A1({ S984 }),
  .A2({ S985 }),
  .B1({ S986 }),
  .B2({ S397 }),
  .ZN({ S987 })
);
NAND2_X1 #() 
NAND2_X1_4770_ (
  .A1({ S987 }),
  .A2({ S25957[901] }),
  .ZN({ S988 })
);
NAND2_X1 #() 
NAND2_X1_4771_ (
  .A1({ S405 }),
  .A2({ S25957[899] }),
  .ZN({ S989 })
);
OAI21_X1 #() 
OAI21_X1_2455_ (
  .A({ S563 }),
  .B1({ S411 }),
  .B2({ S989 }),
  .ZN({ S990 })
);
AOI21_X1 #() 
AOI21_X1_2674_ (
  .A({ S25957[901] }),
  .B1({ S455 }),
  .B2({ S481 }),
  .ZN({ S991 })
);
NAND2_X1 #() 
NAND2_X1_4772_ (
  .A1({ S990 }),
  .A2({ S991 }),
  .ZN({ S992 })
);
NAND3_X1 #() 
NAND3_X1_5169_ (
  .A1({ S988 }),
  .A2({ S25957[902] }),
  .A3({ S992 }),
  .ZN({ S993 })
);
NAND3_X1 #() 
NAND3_X1_5170_ (
  .A1({ S993 }),
  .A2({ S25957[903] }),
  .A3({ S982 }),
  .ZN({ S994 })
);
NAND3_X1 #() 
NAND3_X1_5171_ (
  .A1({ S972 }),
  .A2({ S994 }),
  .A3({ S25957[1002] }),
  .ZN({ S995 })
);
INV_X1 #() 
INV_X1_1539_ (
  .A({ S25957[1002] }),
  .ZN({ S996 })
);
NAND3_X1 #() 
NAND3_X1_5172_ (
  .A1({ S952 }),
  .A2({ S25957[902] }),
  .A3({ S958 }),
  .ZN({ S997 })
);
NAND2_X1 #() 
NAND2_X1_4773_ (
  .A1({ S970 }),
  .A2({ S965 }),
  .ZN({ S998 })
);
NAND2_X1 #() 
NAND2_X1_4774_ (
  .A1({ S998 }),
  .A2({ S353 }),
  .ZN({ S999 })
);
NAND3_X1 #() 
NAND3_X1_5173_ (
  .A1({ S999 }),
  .A2({ S24137 }),
  .A3({ S997 }),
  .ZN({ S1000 })
);
AOI22_X1 #() 
AOI22_X1_543_ (
  .A1({ S987 }),
  .A2({ S25957[901] }),
  .B1({ S991 }),
  .B2({ S990 }),
  .ZN({ S1001 })
);
NAND2_X1 #() 
NAND2_X1_4775_ (
  .A1({ S978 }),
  .A2({ S981 }),
  .ZN({ S1002 })
);
NAND2_X1 #() 
NAND2_X1_4776_ (
  .A1({ S1002 }),
  .A2({ S353 }),
  .ZN({ S1003 })
);
OAI211_X1 #() 
OAI211_X1_1659_ (
  .A({ S25957[903] }),
  .B({ S1003 }),
  .C1({ S1001 }),
  .C2({ S353 }),
  .ZN({ S1004 })
);
NAND3_X1 #() 
NAND3_X1_5174_ (
  .A1({ S1000 }),
  .A2({ S996 }),
  .A3({ S1004 }),
  .ZN({ S1005 })
);
NAND3_X1 #() 
NAND3_X1_5175_ (
  .A1({ S995 }),
  .A2({ S1005 }),
  .A3({ S23926 }),
  .ZN({ S1006 })
);
NAND3_X1 #() 
NAND3_X1_5176_ (
  .A1({ S972 }),
  .A2({ S994 }),
  .A3({ S996 }),
  .ZN({ S1007 })
);
NAND3_X1 #() 
NAND3_X1_5177_ (
  .A1({ S1000 }),
  .A2({ S25957[1002] }),
  .A3({ S1004 }),
  .ZN({ S1008 })
);
NAND3_X1 #() 
NAND3_X1_5178_ (
  .A1({ S1007 }),
  .A2({ S1008 }),
  .A3({ S25957[1066] }),
  .ZN({ S1009 })
);
NAND3_X1 #() 
NAND3_X1_5179_ (
  .A1({ S1006 }),
  .A2({ S1009 }),
  .A3({ S25957[906] }),
  .ZN({ S1010 })
);
NAND3_X1 #() 
NAND3_X1_5180_ (
  .A1({ S1007 }),
  .A2({ S1008 }),
  .A3({ S23926 }),
  .ZN({ S1011 })
);
NAND3_X1 #() 
NAND3_X1_5181_ (
  .A1({ S995 }),
  .A2({ S1005 }),
  .A3({ S25957[1066] }),
  .ZN({ S1012 })
);
NAND3_X1 #() 
NAND3_X1_5182_ (
  .A1({ S1011 }),
  .A2({ S1012 }),
  .A3({ S25436 }),
  .ZN({ S1013 })
);
NAND2_X1 #() 
NAND2_X1_4777_ (
  .A1({ S1010 }),
  .A2({ S1013 }),
  .ZN({ S25957[778] })
);
AOI21_X1 #() 
AOI21_X1_2675_ (
  .A({ S25957[1048] }),
  .B1({ S25264 }),
  .B2({ S25265 }),
  .ZN({ S1014 })
);
AOI21_X1 #() 
AOI21_X1_2676_ (
  .A({ S24021 }),
  .B1({ S25259 }),
  .B2({ S25262 }),
  .ZN({ S1015 })
);
OAI21_X1 #() 
OAI21_X1_2456_ (
  .A({ S25957[921] }),
  .B1({ S1014 }),
  .B2({ S1015 }),
  .ZN({ S1016 })
);
INV_X1 #() 
INV_X1_1540_ (
  .A({ S1016 }),
  .ZN({ S102 })
);
AOI21_X1 #() 
AOI21_X1_2677_ (
  .A({ S25957[1177] }),
  .B1({ S25334 }),
  .B2({ S25333 }),
  .ZN({ S1017 })
);
AND3_X1 #() 
AND3_X1_192_ (
  .A1({ S25334 }),
  .A2({ S25333 }),
  .A3({ S25957[1177] }),
  .ZN({ S1018 })
);
NOR2_X1 #() 
NOR2_X1_1200_ (
  .A1({ S1018 }),
  .A2({ S1017 }),
  .ZN({ S1019 })
);
NAND3_X1 #() 
NAND3_X1_5183_ (
  .A1({ S1019 }),
  .A2({ S25263 }),
  .A3({ S25266 }),
  .ZN({ S103 })
);
XNOR2_X1 #() 
XNOR2_X1_189_ (
  .A({ S25957[1095] }),
  .B({ S24023 }),
  .ZN({ S25957[1063] })
);
INV_X1 #() 
INV_X1_1541_ (
  .A({ S25957[999] }),
  .ZN({ S1020 })
);
INV_X1 #() 
INV_X1_1542_ (
  .A({ S25957[926] }),
  .ZN({ S1021 })
);
AOI21_X1 #() 
AOI21_X1_2678_ (
  .A({ S25957[920] }),
  .B1({ S1019 }),
  .B2({ S25957[922] }),
  .ZN({ S1022 })
);
OAI21_X1 #() 
OAI21_X1_2457_ (
  .A({ S25957[924] }),
  .B1({ S1022 }),
  .B2({ S25957[923] }),
  .ZN({ S1023 })
);
NAND3_X1 #() 
NAND3_X1_5184_ (
  .A1({ S1019 }),
  .A2({ S25402 }),
  .A3({ S25405 }),
  .ZN({ S1024 })
);
NAND2_X1 #() 
NAND2_X1_4778_ (
  .A1({ S25957[920] }),
  .A2({ S25957[922] }),
  .ZN({ S1025 })
);
NAND3_X1 #() 
NAND3_X1_5185_ (
  .A1({ S25263 }),
  .A2({ S25266 }),
  .A3({ S25957[921] }),
  .ZN({ S1026 })
);
NAND2_X1 #() 
NAND2_X1_4779_ (
  .A1({ S1025 }),
  .A2({ S1026 }),
  .ZN({ S1027 })
);
INV_X1 #() 
INV_X1_1543_ (
  .A({ S1027 }),
  .ZN({ S1028 })
);
AOI21_X1 #() 
AOI21_X1_2679_ (
  .A({ S95 }),
  .B1({ S1028 }),
  .B2({ S1024 }),
  .ZN({ S1029 })
);
NAND2_X1 #() 
NAND2_X1_4780_ (
  .A1({ S25957[922] }),
  .A2({ S25957[921] }),
  .ZN({ S1030 })
);
AOI21_X1 #() 
AOI21_X1_2680_ (
  .A({ S25957[1178] }),
  .B1({ S25403 }),
  .B2({ S25404 }),
  .ZN({ S1031 })
);
AOI21_X1 #() 
AOI21_X1_2681_ (
  .A({ S21411 }),
  .B1({ S25397 }),
  .B2({ S25401 }),
  .ZN({ S1032 })
);
NOR2_X1 #() 
NOR2_X1_1201_ (
  .A1({ S1031 }),
  .A2({ S1032 }),
  .ZN({ S1033 })
);
AOI21_X1 #() 
AOI21_X1_2682_ (
  .A({ S25957[921] }),
  .B1({ S25266 }),
  .B2({ S25263 }),
  .ZN({ S1034 })
);
NAND2_X1 #() 
NAND2_X1_4781_ (
  .A1({ S1034 }),
  .A2({ S1033 }),
  .ZN({ S1035 })
);
NAND2_X1 #() 
NAND2_X1_4782_ (
  .A1({ S1035 }),
  .A2({ S1030 }),
  .ZN({ S1036 })
);
NAND2_X1 #() 
NAND2_X1_4783_ (
  .A1({ S1036 }),
  .A2({ S25957[923] }),
  .ZN({ S1037 })
);
NAND2_X1 #() 
NAND2_X1_4784_ (
  .A1({ S25957[922] }),
  .A2({ S1019 }),
  .ZN({ S1038 })
);
OAI211_X1 #() 
OAI211_X1_1660_ (
  .A({ S25263 }),
  .B({ S25266 }),
  .C1({ S1032 }),
  .C2({ S1031 }),
  .ZN({ S1039 })
);
NAND3_X1 #() 
NAND3_X1_5186_ (
  .A1({ S1039 }),
  .A2({ S1038 }),
  .A3({ S95 }),
  .ZN({ S1040 })
);
NAND3_X1 #() 
NAND3_X1_5187_ (
  .A1({ S1037 }),
  .A2({ S25072 }),
  .A3({ S1040 }),
  .ZN({ S1041 })
);
OAI21_X1 #() 
OAI21_X1_2458_ (
  .A({ S1041 }),
  .B1({ S1023 }),
  .B2({ S1029 }),
  .ZN({ S1042 })
);
NAND2_X1 #() 
NAND2_X1_4785_ (
  .A1({ S1016 }),
  .A2({ S25957[922] }),
  .ZN({ S1043 })
);
OAI21_X1 #() 
OAI21_X1_2459_ (
  .A({ S1019 }),
  .B1({ S1014 }),
  .B2({ S1015 }),
  .ZN({ S1044 })
);
NAND3_X1 #() 
NAND3_X1_5188_ (
  .A1({ S1044 }),
  .A2({ S1033 }),
  .A3({ S1026 }),
  .ZN({ S1045 })
);
AOI21_X1 #() 
AOI21_X1_2683_ (
  .A({ S95 }),
  .B1({ S1045 }),
  .B2({ S1043 }),
  .ZN({ S1046 })
);
NAND4_X1 #() 
NAND4_X1_561_ (
  .A1({ S25263 }),
  .A2({ S25266 }),
  .A3({ S25402 }),
  .A4({ S25405 }),
  .ZN({ S1047 })
);
NAND3_X1 #() 
NAND3_X1_5189_ (
  .A1({ S1044 }),
  .A2({ S25957[922] }),
  .A3({ S1026 }),
  .ZN({ S1048 })
);
AOI21_X1 #() 
AOI21_X1_2684_ (
  .A({ S25957[923] }),
  .B1({ S1048 }),
  .B2({ S1047 }),
  .ZN({ S1049 })
);
OR3_X1 #() 
OR3_X1_30_ (
  .A1({ S1049 }),
  .A2({ S1046 }),
  .A3({ S25072 }),
  .ZN({ S1050 })
);
NAND3_X1 #() 
NAND3_X1_5190_ (
  .A1({ S25957[921] }),
  .A2({ S25402 }),
  .A3({ S25405 }),
  .ZN({ S1051 })
);
AOI22_X1 #() 
AOI22_X1_544_ (
  .A1({ S25957[920] }),
  .A2({ S25957[922] }),
  .B1({ S25178 }),
  .B2({ S25177 }),
  .ZN({ S1052 })
);
NAND2_X1 #() 
NAND2_X1_4786_ (
  .A1({ S1052 }),
  .A2({ S1051 }),
  .ZN({ S1053 })
);
NAND3_X1 #() 
NAND3_X1_5191_ (
  .A1({ S1038 }),
  .A2({ S25957[920] }),
  .A3({ S1051 }),
  .ZN({ S1054 })
);
AOI21_X1 #() 
AOI21_X1_2685_ (
  .A({ S25957[924] }),
  .B1({ S1054 }),
  .B2({ S95 }),
  .ZN({ S1055 })
);
AOI21_X1 #() 
AOI21_X1_2686_ (
  .A({ S25957[925] }),
  .B1({ S1055 }),
  .B2({ S1053 }),
  .ZN({ S1056 })
);
AOI22_X1 #() 
AOI22_X1_545_ (
  .A1({ S1042 }),
  .A2({ S25957[925] }),
  .B1({ S1050 }),
  .B2({ S1056 }),
  .ZN({ S1057 })
);
NOR2_X1 #() 
NOR2_X1_1202_ (
  .A1({ S1057 }),
  .A2({ S1021 }),
  .ZN({ S1058 })
);
AND3_X1 #() 
AND3_X1_193_ (
  .A1({ S25957[921] }),
  .A2({ S25402 }),
  .A3({ S25405 }),
  .ZN({ S1059 })
);
NOR2_X1 #() 
NOR2_X1_1203_ (
  .A1({ S1059 }),
  .A2({ S95 }),
  .ZN({ S1060 })
);
NAND2_X1 #() 
NAND2_X1_4787_ (
  .A1({ S1060 }),
  .A2({ S1044 }),
  .ZN({ S1061 })
);
NAND2_X1 #() 
NAND2_X1_4788_ (
  .A1({ S1047 }),
  .A2({ S1024 }),
  .ZN({ S1062 })
);
INV_X1 #() 
INV_X1_1544_ (
  .A({ S1062 }),
  .ZN({ S1063 })
);
AOI22_X1 #() 
AOI22_X1_546_ (
  .A1({ S25957[922] }),
  .A2({ S25957[921] }),
  .B1({ S25176 }),
  .B2({ S25165 }),
  .ZN({ S1064 })
);
NAND2_X1 #() 
NAND2_X1_4789_ (
  .A1({ S1063 }),
  .A2({ S1064 }),
  .ZN({ S1065 })
);
AOI21_X1 #() 
AOI21_X1_2687_ (
  .A({ S25957[924] }),
  .B1({ S1061 }),
  .B2({ S1065 }),
  .ZN({ S1066 })
);
NAND2_X1 #() 
NAND2_X1_4790_ (
  .A1({ S1052 }),
  .A2({ S1024 }),
  .ZN({ S1067 })
);
AOI21_X1 #() 
AOI21_X1_2688_ (
  .A({ S25072 }),
  .B1({ S95 }),
  .B2({ S25957[920] }),
  .ZN({ S1068 })
);
AOI21_X1 #() 
AOI21_X1_2689_ (
  .A({ S1066 }),
  .B1({ S1067 }),
  .B2({ S1068 }),
  .ZN({ S1069 })
);
NAND4_X1 #() 
NAND4_X1_562_ (
  .A1({ S25957[922] }),
  .A2({ S25957[921] }),
  .A3({ S25266 }),
  .A4({ S25263 }),
  .ZN({ S1070 })
);
NAND2_X1 #() 
NAND2_X1_4791_ (
  .A1({ S1070 }),
  .A2({ S25957[923] }),
  .ZN({ S1071 })
);
AND3_X1 #() 
AND3_X1_194_ (
  .A1({ S25263 }),
  .A2({ S25266 }),
  .A3({ S25957[921] }),
  .ZN({ S1072 })
);
OAI21_X1 #() 
OAI21_X1_2460_ (
  .A({ S25957[922] }),
  .B1({ S1072 }),
  .B2({ S1034 }),
  .ZN({ S1073 })
);
AOI21_X1 #() 
AOI21_X1_2690_ (
  .A({ S25957[923] }),
  .B1({ S1059 }),
  .B2({ S25957[920] }),
  .ZN({ S1074 })
);
AOI21_X1 #() 
AOI21_X1_2691_ (
  .A({ S25072 }),
  .B1({ S1073 }),
  .B2({ S1074 }),
  .ZN({ S1075 })
);
NAND3_X1 #() 
NAND3_X1_5192_ (
  .A1({ S1039 }),
  .A2({ S1038 }),
  .A3({ S25957[923] }),
  .ZN({ S1076 })
);
NAND2_X1 #() 
NAND2_X1_4792_ (
  .A1({ S1048 }),
  .A2({ S95 }),
  .ZN({ S1077 })
);
AOI21_X1 #() 
AOI21_X1_2692_ (
  .A({ S25957[924] }),
  .B1({ S1077 }),
  .B2({ S1076 }),
  .ZN({ S1078 })
);
AOI211_X1 #() 
AOI211_X1_85_ (
  .A({ S25957[925] }),
  .B({ S1078 }),
  .C1({ S1071 }),
  .C2({ S1075 }),
  .ZN({ S1079 })
);
AOI21_X1 #() 
AOI21_X1_2693_ (
  .A({ S1079 }),
  .B1({ S1069 }),
  .B2({ S25957[925] }),
  .ZN({ S1080 })
);
AOI21_X1 #() 
AOI21_X1_2694_ (
  .A({ S1058 }),
  .B1({ S1021 }),
  .B2({ S1080 }),
  .ZN({ S1081 })
);
NAND3_X1 #() 
NAND3_X1_5193_ (
  .A1({ S24971 }),
  .A2({ S22294 }),
  .A3({ S24969 }),
  .ZN({ S1082 })
);
NAND3_X1 #() 
NAND3_X1_5194_ (
  .A1({ S24973 }),
  .A2({ S24975 }),
  .A3({ S25957[1053] }),
  .ZN({ S1083 })
);
NAND2_X1 #() 
NAND2_X1_4793_ (
  .A1({ S1082 }),
  .A2({ S1083 }),
  .ZN({ S1084 })
);
INV_X1 #() 
INV_X1_1545_ (
  .A({ S1039 }),
  .ZN({ S1085 })
);
NOR2_X1 #() 
NOR2_X1_1204_ (
  .A1({ S1085 }),
  .A2({ S25957[923] }),
  .ZN({ S1086 })
);
AOI21_X1 #() 
AOI21_X1_2695_ (
  .A({ S1019 }),
  .B1({ S25402 }),
  .B2({ S25405 }),
  .ZN({ S1087 })
);
NOR2_X1 #() 
NOR2_X1_1205_ (
  .A1({ S1014 }),
  .A2({ S1015 }),
  .ZN({ S1088 })
);
NAND2_X1 #() 
NAND2_X1_4794_ (
  .A1({ S1088 }),
  .A2({ S1051 }),
  .ZN({ S1089 })
);
NAND2_X1 #() 
NAND2_X1_4795_ (
  .A1({ S1024 }),
  .A2({ S25957[920] }),
  .ZN({ S1090 })
);
AOI21_X1 #() 
AOI21_X1_2696_ (
  .A({ S1087 }),
  .B1({ S1089 }),
  .B2({ S1090 }),
  .ZN({ S1091 })
);
NAND2_X1 #() 
NAND2_X1_4796_ (
  .A1({ S1091 }),
  .A2({ S1086 }),
  .ZN({ S1092 })
);
AOI21_X1 #() 
AOI21_X1_2697_ (
  .A({ S25957[921] }),
  .B1({ S25177 }),
  .B2({ S25178 }),
  .ZN({ S1093 })
);
NAND2_X1 #() 
NAND2_X1_4797_ (
  .A1({ S1093 }),
  .A2({ S1033 }),
  .ZN({ S1094 })
);
NAND3_X1 #() 
NAND3_X1_5195_ (
  .A1({ S1092 }),
  .A2({ S25072 }),
  .A3({ S1094 }),
  .ZN({ S1095 })
);
OAI211_X1 #() 
OAI211_X1_1661_ (
  .A({ S25402 }),
  .B({ S25405 }),
  .C1({ S1015 }),
  .C2({ S1014 }),
  .ZN({ S1096 })
);
NAND2_X1 #() 
NAND2_X1_4798_ (
  .A1({ S1096 }),
  .A2({ S95 }),
  .ZN({ S1097 })
);
INV_X1 #() 
INV_X1_1546_ (
  .A({ S1097 }),
  .ZN({ S1098 })
);
AOI21_X1 #() 
AOI21_X1_2698_ (
  .A({ S95 }),
  .B1({ S1073 }),
  .B2({ S1045 }),
  .ZN({ S1099 })
);
AOI21_X1 #() 
AOI21_X1_2699_ (
  .A({ S1099 }),
  .B1({ S1098 }),
  .B2({ S1030 }),
  .ZN({ S1100 })
);
OAI21_X1 #() 
OAI21_X1_2461_ (
  .A({ S1095 }),
  .B1({ S1100 }),
  .B2({ S25072 }),
  .ZN({ S1101 })
);
NAND2_X1 #() 
NAND2_X1_4799_ (
  .A1({ S1101 }),
  .A2({ S1084 }),
  .ZN({ S1102 })
);
OAI21_X1 #() 
OAI21_X1_2462_ (
  .A({ S95 }),
  .B1({ S1024 }),
  .B2({ S25957[920] }),
  .ZN({ S1103 })
);
NAND3_X1 #() 
NAND3_X1_5196_ (
  .A1({ S1103 }),
  .A2({ S25072 }),
  .A3({ S1016 }),
  .ZN({ S1104 })
);
INV_X1 #() 
INV_X1_1547_ (
  .A({ S1093 }),
  .ZN({ S1105 })
);
NAND3_X1 #() 
NAND3_X1_5197_ (
  .A1({ S25957[923] }),
  .A2({ S25957[920] }),
  .A3({ S25957[922] }),
  .ZN({ S1106 })
);
AND2_X1 #() 
AND2_X1_294_ (
  .A1({ S1106 }),
  .A2({ S1105 }),
  .ZN({ S1107 })
);
NOR2_X1 #() 
NOR2_X1_1206_ (
  .A1({ S25957[923] }),
  .A2({ S1019 }),
  .ZN({ S1108 })
);
AOI21_X1 #() 
AOI21_X1_2700_ (
  .A({ S25072 }),
  .B1({ S1108 }),
  .B2({ S1025 }),
  .ZN({ S1109 })
);
NAND2_X1 #() 
NAND2_X1_4800_ (
  .A1({ S1107 }),
  .A2({ S1109 }),
  .ZN({ S1110 })
);
NAND3_X1 #() 
NAND3_X1_5198_ (
  .A1({ S1110 }),
  .A2({ S25957[925] }),
  .A3({ S1104 }),
  .ZN({ S1111 })
);
NAND3_X1 #() 
NAND3_X1_5199_ (
  .A1({ S1102 }),
  .A2({ S1021 }),
  .A3({ S1111 }),
  .ZN({ S1112 })
);
AOI21_X1 #() 
AOI21_X1_2701_ (
  .A({ S95 }),
  .B1({ S1024 }),
  .B2({ S1026 }),
  .ZN({ S1113 })
);
INV_X1 #() 
INV_X1_1548_ (
  .A({ S1113 }),
  .ZN({ S1114 })
);
NAND2_X1 #() 
NAND2_X1_4801_ (
  .A1({ S1026 }),
  .A2({ S95 }),
  .ZN({ S1115 })
);
AOI21_X1 #() 
AOI21_X1_2702_ (
  .A({ S25072 }),
  .B1({ S1114 }),
  .B2({ S1115 }),
  .ZN({ S1116 })
);
AOI21_X1 #() 
AOI21_X1_2703_ (
  .A({ S25957[921] }),
  .B1({ S25402 }),
  .B2({ S25405 }),
  .ZN({ S1117 })
);
NAND2_X1 #() 
NAND2_X1_4802_ (
  .A1({ S1117 }),
  .A2({ S1088 }),
  .ZN({ S1118 })
);
NAND2_X1 #() 
NAND2_X1_4803_ (
  .A1({ S103 }),
  .A2({ S1033 }),
  .ZN({ S1119 })
);
NAND3_X1 #() 
NAND3_X1_5200_ (
  .A1({ S1118 }),
  .A2({ S95 }),
  .A3({ S1119 }),
  .ZN({ S1120 })
);
AOI21_X1 #() 
AOI21_X1_2704_ (
  .A({ S25957[924] }),
  .B1({ S1060 }),
  .B2({ S1118 }),
  .ZN({ S1121 })
);
AOI21_X1 #() 
AOI21_X1_2705_ (
  .A({ S1116 }),
  .B1({ S1120 }),
  .B2({ S1121 }),
  .ZN({ S1122 })
);
INV_X1 #() 
INV_X1_1549_ (
  .A({ S1060 }),
  .ZN({ S1123 })
);
NOR2_X1 #() 
NOR2_X1_1207_ (
  .A1({ S1072 }),
  .A2({ S1034 }),
  .ZN({ S1124 })
);
NAND2_X1 #() 
NAND2_X1_4804_ (
  .A1({ S95 }),
  .A2({ S1024 }),
  .ZN({ S1125 })
);
OAI221_X1 #() 
OAI221_X1_141_ (
  .A({ S25072 }),
  .B1({ S1027 }),
  .B2({ S1125 }),
  .C1({ S1123 }),
  .C2({ S1124 }),
  .ZN({ S1126 })
);
NAND2_X1 #() 
NAND2_X1_4805_ (
  .A1({ S1047 }),
  .A2({ S95 }),
  .ZN({ S1127 })
);
NAND2_X1 #() 
NAND2_X1_4806_ (
  .A1({ S1047 }),
  .A2({ S1051 }),
  .ZN({ S1128 })
);
AOI21_X1 #() 
AOI21_X1_2706_ (
  .A({ S25072 }),
  .B1({ S1128 }),
  .B2({ S25957[923] }),
  .ZN({ S1129 })
);
OAI211_X1 #() 
OAI211_X1_1662_ (
  .A({ S1129 }),
  .B({ S1106 }),
  .C1({ S1127 }),
  .C2({ S1019 }),
  .ZN({ S1130 })
);
NAND3_X1 #() 
NAND3_X1_5201_ (
  .A1({ S1126 }),
  .A2({ S1130 }),
  .A3({ S25957[925] }),
  .ZN({ S1131 })
);
OAI21_X1 #() 
OAI21_X1_2463_ (
  .A({ S1131 }),
  .B1({ S1122 }),
  .B2({ S25957[925] }),
  .ZN({ S1132 })
);
OAI211_X1 #() 
OAI211_X1_1663_ (
  .A({ S1112 }),
  .B({ S25957[927] }),
  .C1({ S1021 }),
  .C2({ S1132 }),
  .ZN({ S1133 })
);
OAI21_X1 #() 
OAI21_X1_2464_ (
  .A({ S1133 }),
  .B1({ S1081 }),
  .B2({ S25957[927] }),
  .ZN({ S1134 })
);
OR2_X1 #() 
OR2_X1_65_ (
  .A1({ S1134 }),
  .A2({ S1020 }),
  .ZN({ S1135 })
);
NAND2_X1 #() 
NAND2_X1_4807_ (
  .A1({ S1134 }),
  .A2({ S1020 }),
  .ZN({ S1136 })
);
NAND2_X1 #() 
NAND2_X1_4808_ (
  .A1({ S1135 }),
  .A2({ S1136 }),
  .ZN({ S1137 })
);
NOR2_X1 #() 
NOR2_X1_1208_ (
  .A1({ S1137 }),
  .A2({ S25957[1063] }),
  .ZN({ S1138 })
);
NAND2_X1 #() 
NAND2_X1_4809_ (
  .A1({ S1137 }),
  .A2({ S25957[1063] }),
  .ZN({ S1139 })
);
INV_X1 #() 
INV_X1_1550_ (
  .A({ S1139 }),
  .ZN({ S1140 })
);
NOR2_X1 #() 
NOR2_X1_1209_ (
  .A1({ S1140 }),
  .A2({ S1138 }),
  .ZN({ S1141 })
);
XNOR2_X1 #() 
XNOR2_X1_190_ (
  .A({ S1141 }),
  .B({ S25957[903] }),
  .ZN({ S25957[775] })
);
XNOR2_X1 #() 
XNOR2_X1_191_ (
  .A({ S24206 }),
  .B({ S25957[1126] }),
  .ZN({ S25957[998] })
);
INV_X1 #() 
INV_X1_1551_ (
  .A({ S25957[998] }),
  .ZN({ S1142 })
);
NAND4_X1 #() 
NAND4_X1_563_ (
  .A1({ S1096 }),
  .A2({ S1039 }),
  .A3({ S1038 }),
  .A4({ S95 }),
  .ZN({ S1143 })
);
OAI21_X1 #() 
OAI21_X1_2465_ (
  .A({ S1143 }),
  .B1({ S1028 }),
  .B2({ S95 }),
  .ZN({ S1144 })
);
NAND2_X1 #() 
NAND2_X1_4810_ (
  .A1({ S1030 }),
  .A2({ S1026 }),
  .ZN({ S1145 })
);
NAND2_X1 #() 
NAND2_X1_4811_ (
  .A1({ S1106 }),
  .A2({ S25072 }),
  .ZN({ S1146 })
);
OAI21_X1 #() 
OAI21_X1_2466_ (
  .A({ S25957[925] }),
  .B1({ S1146 }),
  .B2({ S1145 }),
  .ZN({ S1147 })
);
AOI21_X1 #() 
AOI21_X1_2707_ (
  .A({ S1147 }),
  .B1({ S1144 }),
  .B2({ S25957[924] }),
  .ZN({ S1148 })
);
NAND2_X1 #() 
NAND2_X1_4812_ (
  .A1({ S1034 }),
  .A2({ S25957[922] }),
  .ZN({ S1149 })
);
NAND2_X1 #() 
NAND2_X1_4813_ (
  .A1({ S1149 }),
  .A2({ S1070 }),
  .ZN({ S1150 })
);
NAND3_X1 #() 
NAND3_X1_5202_ (
  .A1({ S1149 }),
  .A2({ S25957[923] }),
  .A3({ S1047 }),
  .ZN({ S1151 })
);
OAI211_X1 #() 
OAI211_X1_1664_ (
  .A({ S1151 }),
  .B({ S25072 }),
  .C1({ S1150 }),
  .C2({ S25957[923] }),
  .ZN({ S1152 })
);
NAND2_X1 #() 
NAND2_X1_4814_ (
  .A1({ S1088 }),
  .A2({ S1024 }),
  .ZN({ S1153 })
);
INV_X1 #() 
INV_X1_1552_ (
  .A({ S1153 }),
  .ZN({ S1154 })
);
NAND2_X1 #() 
NAND2_X1_4815_ (
  .A1({ S1154 }),
  .A2({ S95 }),
  .ZN({ S1155 })
);
AOI21_X1 #() 
AOI21_X1_2708_ (
  .A({ S25072 }),
  .B1({ S1059 }),
  .B2({ S25957[923] }),
  .ZN({ S1156 })
);
NAND2_X1 #() 
NAND2_X1_4816_ (
  .A1({ S1155 }),
  .A2({ S1156 }),
  .ZN({ S1157 })
);
AND3_X1 #() 
AND3_X1_195_ (
  .A1({ S1152 }),
  .A2({ S1084 }),
  .A3({ S1157 }),
  .ZN({ S1158 })
);
OAI21_X1 #() 
OAI21_X1_2467_ (
  .A({ S25957[926] }),
  .B1({ S1158 }),
  .B2({ S1148 }),
  .ZN({ S1159 })
);
INV_X1 #() 
INV_X1_1553_ (
  .A({ S1024 }),
  .ZN({ S1160 })
);
NOR2_X1 #() 
NOR2_X1_1210_ (
  .A1({ S1160 }),
  .A2({ S95 }),
  .ZN({ S1161 })
);
AOI22_X1 #() 
AOI22_X1_547_ (
  .A1({ S1036 }),
  .A2({ S95 }),
  .B1({ S1161 }),
  .B2({ S1030 }),
  .ZN({ S1162 })
);
OAI21_X1 #() 
OAI21_X1_2468_ (
  .A({ S25957[923] }),
  .B1({ S103 }),
  .B2({ S1033 }),
  .ZN({ S1163 })
);
OAI21_X1 #() 
OAI21_X1_2469_ (
  .A({ S1097 }),
  .B1({ S1163 }),
  .B2({ S102 }),
  .ZN({ S1164 })
);
MUX2_X1 #() 
MUX2_X1_19_ (
  .A({ S1164 }),
  .B({ S1162 }),
  .S({ S25072 }),
  .Z({ S1165 })
);
AOI21_X1 #() 
AOI21_X1_2709_ (
  .A({ S25957[923] }),
  .B1({ S1034 }),
  .B2({ S1033 }),
  .ZN({ S1166 })
);
NAND2_X1 #() 
NAND2_X1_4817_ (
  .A1({ S1037 }),
  .A2({ S25957[924] }),
  .ZN({ S1167 })
);
NOR2_X1 #() 
NOR2_X1_1211_ (
  .A1({ S1167 }),
  .A2({ S1166 }),
  .ZN({ S1168 })
);
NAND2_X1 #() 
NAND2_X1_4818_ (
  .A1({ S1033 }),
  .A2({ S1026 }),
  .ZN({ S1169 })
);
AOI21_X1 #() 
AOI21_X1_2710_ (
  .A({ S95 }),
  .B1({ S1169 }),
  .B2({ S1070 }),
  .ZN({ S1170 })
);
AOI21_X1 #() 
AOI21_X1_2711_ (
  .A({ S1168 }),
  .B1({ S25072 }),
  .B2({ S1170 }),
  .ZN({ S1171 })
);
NAND2_X1 #() 
NAND2_X1_4819_ (
  .A1({ S1171 }),
  .A2({ S1084 }),
  .ZN({ S1172 })
);
OAI211_X1 #() 
OAI211_X1_1665_ (
  .A({ S1172 }),
  .B({ S1021 }),
  .C1({ S1165 }),
  .C2({ S1084 }),
  .ZN({ S1173 })
);
AOI21_X1 #() 
AOI21_X1_2712_ (
  .A({ S25957[927] }),
  .B1({ S1173 }),
  .B2({ S1159 }),
  .ZN({ S1174 })
);
INV_X1 #() 
INV_X1_1554_ (
  .A({ S1151 }),
  .ZN({ S1175 })
);
AOI21_X1 #() 
AOI21_X1_2713_ (
  .A({ S1175 }),
  .B1({ S1089 }),
  .B2({ S1074 }),
  .ZN({ S1176 })
);
NAND4_X1 #() 
NAND4_X1_564_ (
  .A1({ S1038 }),
  .A2({ S1051 }),
  .A3({ S25957[920] }),
  .A4({ S95 }),
  .ZN({ S1177 })
);
NOR2_X1 #() 
NOR2_X1_1212_ (
  .A1({ S95 }),
  .A2({ S25957[920] }),
  .ZN({ S1178 })
);
AOI21_X1 #() 
AOI21_X1_2714_ (
  .A({ S25957[924] }),
  .B1({ S1178 }),
  .B2({ S1030 }),
  .ZN({ S1179 })
);
NAND3_X1 #() 
NAND3_X1_5203_ (
  .A1({ S1179 }),
  .A2({ S1094 }),
  .A3({ S1177 }),
  .ZN({ S1180 })
);
OAI21_X1 #() 
OAI21_X1_2470_ (
  .A({ S1180 }),
  .B1({ S1176 }),
  .B2({ S25072 }),
  .ZN({ S1181 })
);
NAND2_X1 #() 
NAND2_X1_4820_ (
  .A1({ S103 }),
  .A2({ S25957[922] }),
  .ZN({ S1182 })
);
NAND3_X1 #() 
NAND3_X1_5204_ (
  .A1({ S1096 }),
  .A2({ S1093 }),
  .A3({ S1039 }),
  .ZN({ S1183 })
);
OAI21_X1 #() 
OAI21_X1_2471_ (
  .A({ S1183 }),
  .B1({ S25957[923] }),
  .B2({ S1182 }),
  .ZN({ S1184 })
);
OAI21_X1 #() 
OAI21_X1_2472_ (
  .A({ S25072 }),
  .B1({ S1113 }),
  .B2({ S1108 }),
  .ZN({ S1185 })
);
OAI211_X1 #() 
OAI211_X1_1666_ (
  .A({ S25957[925] }),
  .B({ S1185 }),
  .C1({ S1184 }),
  .C2({ S25072 }),
  .ZN({ S1186 })
);
OAI211_X1 #() 
OAI211_X1_1667_ (
  .A({ S25957[926] }),
  .B({ S1186 }),
  .C1({ S1181 }),
  .C2({ S25957[925] }),
  .ZN({ S1187 })
);
INV_X1 #() 
INV_X1_1555_ (
  .A({ S1124 }),
  .ZN({ S1188 })
);
NAND2_X1 #() 
NAND2_X1_4821_ (
  .A1({ S95 }),
  .A2({ S1051 }),
  .ZN({ S1189 })
);
OAI21_X1 #() 
OAI21_X1_2473_ (
  .A({ S25957[923] }),
  .B1({ S1051 }),
  .B2({ S25957[920] }),
  .ZN({ S1190 })
);
OAI22_X1 #() 
OAI22_X1_123_ (
  .A1({ S1188 }),
  .A2({ S1189 }),
  .B1({ S1190 }),
  .B2({ S1117 }),
  .ZN({ S1191 })
);
NAND2_X1 #() 
NAND2_X1_4822_ (
  .A1({ S1087 }),
  .A2({ S25957[923] }),
  .ZN({ S1192 })
);
NOR2_X1 #() 
NOR2_X1_1213_ (
  .A1({ S1051 }),
  .A2({ S25957[920] }),
  .ZN({ S1193 })
);
NAND2_X1 #() 
NAND2_X1_4823_ (
  .A1({ S1193 }),
  .A2({ S95 }),
  .ZN({ S1194 })
);
NAND2_X1 #() 
NAND2_X1_4824_ (
  .A1({ S1194 }),
  .A2({ S1192 }),
  .ZN({ S1195 })
);
NOR2_X1 #() 
NOR2_X1_1214_ (
  .A1({ S1048 }),
  .A2({ S25957[923] }),
  .ZN({ S1196 })
);
OAI21_X1 #() 
OAI21_X1_2474_ (
  .A({ S25957[924] }),
  .B1({ S1195 }),
  .B2({ S1196 }),
  .ZN({ S1197 })
);
OAI21_X1 #() 
OAI21_X1_2475_ (
  .A({ S1197 }),
  .B1({ S1191 }),
  .B2({ S25957[924] }),
  .ZN({ S1198 })
);
NAND2_X1 #() 
NAND2_X1_4825_ (
  .A1({ S1026 }),
  .A2({ S25957[922] }),
  .ZN({ S1199 })
);
NAND3_X1 #() 
NAND3_X1_5205_ (
  .A1({ S1199 }),
  .A2({ S25957[923] }),
  .A3({ S1047 }),
  .ZN({ S1200 })
);
AOI21_X1 #() 
AOI21_X1_2715_ (
  .A({ S25957[924] }),
  .B1({ S1074 }),
  .B2({ S1089 }),
  .ZN({ S1201 })
);
NAND2_X1 #() 
NAND2_X1_4826_ (
  .A1({ S1201 }),
  .A2({ S1200 }),
  .ZN({ S1202 })
);
NAND2_X1 #() 
NAND2_X1_4827_ (
  .A1({ S1044 }),
  .A2({ S1033 }),
  .ZN({ S1203 })
);
OAI21_X1 #() 
OAI21_X1_2476_ (
  .A({ S1107 }),
  .B1({ S25957[923] }),
  .B2({ S1203 }),
  .ZN({ S1204 })
);
NAND2_X1 #() 
NAND2_X1_4828_ (
  .A1({ S1204 }),
  .A2({ S25957[924] }),
  .ZN({ S1205 })
);
NAND2_X1 #() 
NAND2_X1_4829_ (
  .A1({ S1205 }),
  .A2({ S1202 }),
  .ZN({ S1206 })
);
AOI21_X1 #() 
AOI21_X1_2716_ (
  .A({ S25957[926] }),
  .B1({ S1206 }),
  .B2({ S1084 }),
  .ZN({ S1207 })
);
OAI21_X1 #() 
OAI21_X1_2477_ (
  .A({ S1207 }),
  .B1({ S1084 }),
  .B2({ S1198 }),
  .ZN({ S1208 })
);
AOI21_X1 #() 
AOI21_X1_2717_ (
  .A({ S24835 }),
  .B1({ S1208 }),
  .B2({ S1187 }),
  .ZN({ S1209 })
);
OAI21_X1 #() 
OAI21_X1_2478_ (
  .A({ S1142 }),
  .B1({ S1174 }),
  .B2({ S1209 }),
  .ZN({ S1210 })
);
INV_X1 #() 
INV_X1_1556_ (
  .A({ S1174 }),
  .ZN({ S1211 })
);
INV_X1 #() 
INV_X1_1557_ (
  .A({ S1209 }),
  .ZN({ S1212 })
);
NAND3_X1 #() 
NAND3_X1_5206_ (
  .A1({ S1211 }),
  .A2({ S1212 }),
  .A3({ S25957[998] }),
  .ZN({ S1213 })
);
NAND3_X1 #() 
NAND3_X1_5207_ (
  .A1({ S1213 }),
  .A2({ S25957[1062] }),
  .A3({ S1210 }),
  .ZN({ S1214 })
);
INV_X1 #() 
INV_X1_1558_ (
  .A({ S25957[1062] }),
  .ZN({ S1215 })
);
NAND3_X1 #() 
NAND3_X1_5208_ (
  .A1({ S1211 }),
  .A2({ S1212 }),
  .A3({ S1142 }),
  .ZN({ S1216 })
);
OAI21_X1 #() 
OAI21_X1_2479_ (
  .A({ S25957[998] }),
  .B1({ S1174 }),
  .B2({ S1209 }),
  .ZN({ S1217 })
);
NAND3_X1 #() 
NAND3_X1_5209_ (
  .A1({ S1216 }),
  .A2({ S1215 }),
  .A3({ S1217 }),
  .ZN({ S1218 })
);
AOI21_X1 #() 
AOI21_X1_2718_ (
  .A({ S25957[902] }),
  .B1({ S1214 }),
  .B2({ S1218 }),
  .ZN({ S1219 })
);
AND3_X1 #() 
AND3_X1_196_ (
  .A1({ S1218 }),
  .A2({ S1214 }),
  .A3({ S25957[902] }),
  .ZN({ S1220 })
);
NOR2_X1 #() 
NOR2_X1_1215_ (
  .A1({ S1220 }),
  .A2({ S1219 }),
  .ZN({ S25957[774] })
);
NOR2_X1 #() 
NOR2_X1_1216_ (
  .A1({ S21648 }),
  .A2({ S21652 }),
  .ZN({ S25957[1093] })
);
INV_X1 #() 
INV_X1_1559_ (
  .A({ S25957[1093] }),
  .ZN({ S1221 })
);
AOI21_X1 #() 
AOI21_X1_2719_ (
  .A({ S1019 }),
  .B1({ S25177 }),
  .B2({ S25178 }),
  .ZN({ S1222 })
);
OAI21_X1 #() 
OAI21_X1_2480_ (
  .A({ S95 }),
  .B1({ S1051 }),
  .B2({ S25957[920] }),
  .ZN({ S1223 })
);
NAND4_X1 #() 
NAND4_X1_565_ (
  .A1({ S1096 }),
  .A2({ S1039 }),
  .A3({ S1038 }),
  .A4({ S25957[923] }),
  .ZN({ S1224 })
);
AOI21_X1 #() 
AOI21_X1_2720_ (
  .A({ S25957[924] }),
  .B1({ S1224 }),
  .B2({ S1223 }),
  .ZN({ S1225 })
);
OAI21_X1 #() 
OAI21_X1_2481_ (
  .A({ S1225 }),
  .B1({ S1025 }),
  .B2({ S1222 }),
  .ZN({ S1226 })
);
NAND3_X1 #() 
NAND3_X1_5210_ (
  .A1({ S25957[920] }),
  .A2({ S25957[921] }),
  .A3({ S25957[922] }),
  .ZN({ S1227 })
);
NAND3_X1 #() 
NAND3_X1_5211_ (
  .A1({ S1063 }),
  .A2({ S95 }),
  .A3({ S1227 }),
  .ZN({ S1228 })
);
AOI21_X1 #() 
AOI21_X1_2721_ (
  .A({ S25957[925] }),
  .B1({ S1228 }),
  .B2({ S1129 }),
  .ZN({ S1229 })
);
NAND2_X1 #() 
NAND2_X1_4830_ (
  .A1({ S1229 }),
  .A2({ S1226 }),
  .ZN({ S1230 })
);
NOR2_X1 #() 
NOR2_X1_1217_ (
  .A1({ S1199 }),
  .A2({ S1034 }),
  .ZN({ S1231 })
);
NAND2_X1 #() 
NAND2_X1_4831_ (
  .A1({ S1036 }),
  .A2({ S95 }),
  .ZN({ S1232 })
);
OAI21_X1 #() 
OAI21_X1_2482_ (
  .A({ S1232 }),
  .B1({ S1231 }),
  .B2({ S1190 }),
  .ZN({ S1233 })
);
AOI21_X1 #() 
AOI21_X1_2722_ (
  .A({ S25957[923] }),
  .B1({ S1025 }),
  .B2({ S103 }),
  .ZN({ S1234 })
);
OAI21_X1 #() 
OAI21_X1_2483_ (
  .A({ S25072 }),
  .B1({ S1234 }),
  .B2({ S1178 }),
  .ZN({ S1235 })
);
OAI211_X1 #() 
OAI211_X1_1668_ (
  .A({ S25957[925] }),
  .B({ S1235 }),
  .C1({ S1233 }),
  .C2({ S25072 }),
  .ZN({ S1236 })
);
NAND2_X1 #() 
NAND2_X1_4832_ (
  .A1({ S1236 }),
  .A2({ S1230 }),
  .ZN({ S1237 })
);
NAND3_X1 #() 
NAND3_X1_5212_ (
  .A1({ S1048 }),
  .A2({ S25957[923] }),
  .A3({ S1035 }),
  .ZN({ S1238 })
);
NAND4_X1 #() 
NAND4_X1_566_ (
  .A1({ S1044 }),
  .A2({ S95 }),
  .A3({ S1024 }),
  .A4({ S1026 }),
  .ZN({ S1239 })
);
NAND3_X1 #() 
NAND3_X1_5213_ (
  .A1({ S1238 }),
  .A2({ S25957[924] }),
  .A3({ S1239 }),
  .ZN({ S1240 })
);
INV_X1 #() 
INV_X1_1560_ (
  .A({ S1222 }),
  .ZN({ S1241 })
);
NOR2_X1 #() 
NOR2_X1_1218_ (
  .A1({ S1064 }),
  .A2({ S25957[924] }),
  .ZN({ S1242 })
);
NAND3_X1 #() 
NAND3_X1_5214_ (
  .A1({ S1242 }),
  .A2({ S25957[920] }),
  .A3({ S1241 }),
  .ZN({ S1243 })
);
AND3_X1 #() 
AND3_X1_197_ (
  .A1({ S1240 }),
  .A2({ S1084 }),
  .A3({ S1243 }),
  .ZN({ S1244 })
);
OAI21_X1 #() 
OAI21_X1_2484_ (
  .A({ S1194 }),
  .B1({ S95 }),
  .B2({ S1062 }),
  .ZN({ S1245 })
);
AOI21_X1 #() 
AOI21_X1_2723_ (
  .A({ S1146 }),
  .B1({ S1086 }),
  .B2({ S1145 }),
  .ZN({ S1246 })
);
AOI21_X1 #() 
AOI21_X1_2724_ (
  .A({ S1246 }),
  .B1({ S1245 }),
  .B2({ S25957[924] }),
  .ZN({ S1247 })
);
OAI21_X1 #() 
OAI21_X1_2485_ (
  .A({ S1021 }),
  .B1({ S1247 }),
  .B2({ S1084 }),
  .ZN({ S1248 })
);
OAI221_X1 #() 
OAI221_X1_142_ (
  .A({ S24835 }),
  .B1({ S1244 }),
  .B2({ S1248 }),
  .C1({ S1021 }),
  .C2({ S1237 }),
  .ZN({ S1249 })
);
AND2_X1 #() 
AND2_X1_295_ (
  .A1({ S1026 }),
  .A2({ S25957[922] }),
  .ZN({ S1250 })
);
OAI21_X1 #() 
OAI21_X1_2486_ (
  .A({ S25957[923] }),
  .B1({ S1250 }),
  .B2({ S1062 }),
  .ZN({ S1251 })
);
AND3_X1 #() 
AND3_X1_198_ (
  .A1({ S103 }),
  .A2({ S95 }),
  .A3({ S1024 }),
  .ZN({ S1252 })
);
INV_X1 #() 
INV_X1_1561_ (
  .A({ S1252 }),
  .ZN({ S1253 })
);
AOI21_X1 #() 
AOI21_X1_2725_ (
  .A({ S25957[924] }),
  .B1({ S1251 }),
  .B2({ S1253 }),
  .ZN({ S1254 })
);
INV_X1 #() 
INV_X1_1562_ (
  .A({ S1070 }),
  .ZN({ S1255 })
);
NOR3_X1 #() 
NOR3_X1_161_ (
  .A1({ S1255 }),
  .A2({ S1128 }),
  .A3({ S25957[923] }),
  .ZN({ S1256 })
);
OAI21_X1 #() 
OAI21_X1_2487_ (
  .A({ S25957[924] }),
  .B1({ S1153 }),
  .B2({ S95 }),
  .ZN({ S1257 })
);
OAI21_X1 #() 
OAI21_X1_2488_ (
  .A({ S25957[925] }),
  .B1({ S1256 }),
  .B2({ S1257 }),
  .ZN({ S1258 })
);
OAI21_X1 #() 
OAI21_X1_2489_ (
  .A({ S25072 }),
  .B1({ S1175 }),
  .B2({ S1196 }),
  .ZN({ S1259 })
);
NOR2_X1 #() 
NOR2_X1_1219_ (
  .A1({ S1199 }),
  .A2({ S25957[923] }),
  .ZN({ S1260 })
);
AOI21_X1 #() 
AOI21_X1_2726_ (
  .A({ S1260 }),
  .B1({ S1169 }),
  .B2({ S25957[923] }),
  .ZN({ S1261 })
);
OAI211_X1 #() 
OAI211_X1_1669_ (
  .A({ S1259 }),
  .B({ S1084 }),
  .C1({ S25072 }),
  .C2({ S1261 }),
  .ZN({ S1262 })
);
OAI211_X1 #() 
OAI211_X1_1670_ (
  .A({ S1262 }),
  .B({ S25957[926] }),
  .C1({ S1254 }),
  .C2({ S1258 }),
  .ZN({ S1263 })
);
NAND2_X1 #() 
NAND2_X1_4833_ (
  .A1({ S1108 }),
  .A2({ S25957[920] }),
  .ZN({ S1264 })
);
OAI21_X1 #() 
OAI21_X1_2490_ (
  .A({ S1127 }),
  .B1({ S1054 }),
  .B2({ S95 }),
  .ZN({ S1265 })
);
AOI21_X1 #() 
AOI21_X1_2727_ (
  .A({ S25072 }),
  .B1({ S1265 }),
  .B2({ S1264 }),
  .ZN({ S1266 })
);
NAND3_X1 #() 
NAND3_X1_5215_ (
  .A1({ S1026 }),
  .A2({ S95 }),
  .A3({ S1024 }),
  .ZN({ S1267 })
);
NOR2_X1 #() 
NOR2_X1_1220_ (
  .A1({ S25957[924] }),
  .A2({ S1093 }),
  .ZN({ S1268 })
);
AOI21_X1 #() 
AOI21_X1_2728_ (
  .A({ S1266 }),
  .B1({ S1267 }),
  .B2({ S1268 }),
  .ZN({ S1269 })
);
INV_X1 #() 
INV_X1_1563_ (
  .A({ S1074 }),
  .ZN({ S1270 })
);
NAND3_X1 #() 
NAND3_X1_5216_ (
  .A1({ S1048 }),
  .A2({ S25957[923] }),
  .A3({ S1119 }),
  .ZN({ S1271 })
);
AOI21_X1 #() 
AOI21_X1_2729_ (
  .A({ S25957[924] }),
  .B1({ S1271 }),
  .B2({ S1270 }),
  .ZN({ S1272 })
);
NAND3_X1 #() 
NAND3_X1_5217_ (
  .A1({ S1016 }),
  .A2({ S1033 }),
  .A3({ S103 }),
  .ZN({ S1273 })
);
NOR2_X1 #() 
NOR2_X1_1221_ (
  .A1({ S1273 }),
  .A2({ S95 }),
  .ZN({ S1274 })
);
OAI21_X1 #() 
OAI21_X1_2491_ (
  .A({ S25957[924] }),
  .B1({ S1097 }),
  .B2({ S25957[921] }),
  .ZN({ S1275 })
);
OAI21_X1 #() 
OAI21_X1_2492_ (
  .A({ S1084 }),
  .B1({ S1275 }),
  .B2({ S1274 }),
  .ZN({ S1276 })
);
OAI221_X1 #() 
OAI221_X1_143_ (
  .A({ S1021 }),
  .B1({ S1276 }),
  .B2({ S1272 }),
  .C1({ S1269 }),
  .C2({ S1084 }),
  .ZN({ S1277 })
);
NAND3_X1 #() 
NAND3_X1_5218_ (
  .A1({ S1277 }),
  .A2({ S25957[927] }),
  .A3({ S1263 }),
  .ZN({ S1278 })
);
NAND2_X1 #() 
NAND2_X1_4834_ (
  .A1({ S1249 }),
  .A2({ S1278 }),
  .ZN({ S1279 })
);
NAND2_X1 #() 
NAND2_X1_4835_ (
  .A1({ S1279 }),
  .A2({ S1221 }),
  .ZN({ S1280 })
);
NOR2_X1 #() 
NOR2_X1_1222_ (
  .A1({ S1279 }),
  .A2({ S1221 }),
  .ZN({ S1281 })
);
INV_X1 #() 
INV_X1_1564_ (
  .A({ S1281 }),
  .ZN({ S1282 })
);
NAND3_X1 #() 
NAND3_X1_5219_ (
  .A1({ S1282 }),
  .A2({ S25957[1029] }),
  .A3({ S1280 }),
  .ZN({ S1283 })
);
INV_X1 #() 
INV_X1_1565_ (
  .A({ S1280 }),
  .ZN({ S1284 })
);
OAI21_X1 #() 
OAI21_X1_2493_ (
  .A({ S23368 }),
  .B1({ S1284 }),
  .B2({ S1281 }),
  .ZN({ S1285 })
);
NAND2_X1 #() 
NAND2_X1_4836_ (
  .A1({ S1285 }),
  .A2({ S1283 }),
  .ZN({ S25957[773] })
);
NAND2_X1 #() 
NAND2_X1_4837_ (
  .A1({ S24357 }),
  .A2({ S24359 }),
  .ZN({ S25957[932] })
);
NAND2_X1 #() 
NAND2_X1_4838_ (
  .A1({ S21740 }),
  .A2({ S21741 }),
  .ZN({ S1286 })
);
INV_X1 #() 
INV_X1_1566_ (
  .A({ S1286 }),
  .ZN({ S25957[1092] })
);
AOI21_X1 #() 
AOI21_X1_2730_ (
  .A({ S25957[923] }),
  .B1({ S1273 }),
  .B2({ S1199 }),
  .ZN({ S1287 })
);
NAND2_X1 #() 
NAND2_X1_4839_ (
  .A1({ S1224 }),
  .A2({ S25072 }),
  .ZN({ S1288 })
);
INV_X1 #() 
INV_X1_1567_ (
  .A({ S130 }),
  .ZN({ S1289 })
);
OAI21_X1 #() 
OAI21_X1_2494_ (
  .A({ S25957[924] }),
  .B1({ S1289 }),
  .B2({ S25957[922] }),
  .ZN({ S1290 })
);
OAI211_X1 #() 
OAI211_X1_1671_ (
  .A({ S25957[926] }),
  .B({ S1290 }),
  .C1({ S1288 }),
  .C2({ S1287 }),
  .ZN({ S1291 })
);
NOR2_X1 #() 
NOR2_X1_1223_ (
  .A1({ S1167 }),
  .A2({ S1260 }),
  .ZN({ S1292 })
);
INV_X1 #() 
INV_X1_1568_ (
  .A({ S1274 }),
  .ZN({ S1293 })
);
AOI21_X1 #() 
AOI21_X1_2731_ (
  .A({ S25957[924] }),
  .B1({ S1293 }),
  .B2({ S1264 }),
  .ZN({ S1294 })
);
OAI21_X1 #() 
OAI21_X1_2495_ (
  .A({ S1021 }),
  .B1({ S1292 }),
  .B2({ S1294 }),
  .ZN({ S1295 })
);
AOI21_X1 #() 
AOI21_X1_2732_ (
  .A({ S1084 }),
  .B1({ S1295 }),
  .B2({ S1291 }),
  .ZN({ S1296 })
);
NAND3_X1 #() 
NAND3_X1_5220_ (
  .A1({ S1025 }),
  .A2({ S25957[923] }),
  .A3({ S103 }),
  .ZN({ S1297 })
);
AND2_X1 #() 
AND2_X1_296_ (
  .A1({ S1120 }),
  .A2({ S1297 }),
  .ZN({ S1298 })
);
NAND2_X1 #() 
NAND2_X1_4840_ (
  .A1({ S1025 }),
  .A2({ S25957[923] }),
  .ZN({ S1299 })
);
NOR2_X1 #() 
NOR2_X1_1224_ (
  .A1({ S1299 }),
  .A2({ S1128 }),
  .ZN({ S1300 })
);
NAND2_X1 #() 
NAND2_X1_4841_ (
  .A1({ S1267 }),
  .A2({ S25957[924] }),
  .ZN({ S1301 })
);
OAI22_X1 #() 
OAI22_X1_124_ (
  .A1({ S1298 }),
  .A2({ S25957[924] }),
  .B1({ S1301 }),
  .B2({ S1300 }),
  .ZN({ S1302 })
);
NAND2_X1 #() 
NAND2_X1_4842_ (
  .A1({ S1302 }),
  .A2({ S1021 }),
  .ZN({ S1303 })
);
NAND3_X1 #() 
NAND3_X1_5221_ (
  .A1({ S1182 }),
  .A2({ S95 }),
  .A3({ S1024 }),
  .ZN({ S1304 })
);
NAND3_X1 #() 
NAND3_X1_5222_ (
  .A1({ S1107 }),
  .A2({ S25957[924] }),
  .A3({ S1304 }),
  .ZN({ S1305 })
);
AOI21_X1 #() 
AOI21_X1_2733_ (
  .A({ S25957[924] }),
  .B1({ S25957[923] }),
  .B2({ S25957[922] }),
  .ZN({ S1306 })
);
OAI21_X1 #() 
OAI21_X1_2496_ (
  .A({ S1306 }),
  .B1({ S1270 }),
  .B2({ S1085 }),
  .ZN({ S1307 })
);
NAND3_X1 #() 
NAND3_X1_5223_ (
  .A1({ S1307 }),
  .A2({ S1305 }),
  .A3({ S25957[926] }),
  .ZN({ S1308 })
);
AOI21_X1 #() 
AOI21_X1_2734_ (
  .A({ S25957[925] }),
  .B1({ S1303 }),
  .B2({ S1308 }),
  .ZN({ S1309 })
);
OAI21_X1 #() 
OAI21_X1_2497_ (
  .A({ S24835 }),
  .B1({ S1296 }),
  .B2({ S1309 }),
  .ZN({ S1310 })
);
OAI21_X1 #() 
OAI21_X1_2498_ (
  .A({ S95 }),
  .B1({ S1250 }),
  .B2({ S1062 }),
  .ZN({ S1311 })
);
INV_X1 #() 
INV_X1_1569_ (
  .A({ S1311 }),
  .ZN({ S1312 })
);
OAI21_X1 #() 
OAI21_X1_2499_ (
  .A({ S25957[924] }),
  .B1({ S1123 }),
  .B2({ S1250 }),
  .ZN({ S1313 })
);
AND2_X1 #() 
AND2_X1_297_ (
  .A1({ S1025 }),
  .A2({ S1093 }),
  .ZN({ S1314 })
);
OAI21_X1 #() 
OAI21_X1_2500_ (
  .A({ S25072 }),
  .B1({ S1250 }),
  .B2({ S1223 }),
  .ZN({ S1315 })
);
OAI221_X1 #() 
OAI221_X1_144_ (
  .A({ S1084 }),
  .B1({ S1314 }),
  .B2({ S1315 }),
  .C1({ S1312 }),
  .C2({ S1313 }),
  .ZN({ S1316 })
);
NAND3_X1 #() 
NAND3_X1_5224_ (
  .A1({ S1039 }),
  .A2({ S1016 }),
  .A3({ S1024 }),
  .ZN({ S1317 })
);
NAND2_X1 #() 
NAND2_X1_4843_ (
  .A1({ S1317 }),
  .A2({ S95 }),
  .ZN({ S1318 })
);
OAI211_X1 #() 
OAI211_X1_1672_ (
  .A({ S1318 }),
  .B({ S25957[924] }),
  .C1({ S1034 }),
  .C2({ S1190 }),
  .ZN({ S1319 })
);
INV_X1 #() 
INV_X1_1570_ (
  .A({ S1319 }),
  .ZN({ S1320 })
);
AOI21_X1 #() 
AOI21_X1_2735_ (
  .A({ S25957[923] }),
  .B1({ S1045 }),
  .B2({ S1043 }),
  .ZN({ S1321 })
);
NAND3_X1 #() 
NAND3_X1_5225_ (
  .A1({ S1044 }),
  .A2({ S25957[923] }),
  .A3({ S1033 }),
  .ZN({ S1322 })
);
OAI211_X1 #() 
OAI211_X1_1673_ (
  .A({ S1322 }),
  .B({ S25072 }),
  .C1({ S95 }),
  .C2({ S1070 }),
  .ZN({ S1323 })
);
OAI21_X1 #() 
OAI21_X1_2501_ (
  .A({ S25957[925] }),
  .B1({ S1323 }),
  .B2({ S1321 }),
  .ZN({ S1324 })
);
OAI211_X1 #() 
OAI211_X1_1674_ (
  .A({ S1316 }),
  .B({ S1021 }),
  .C1({ S1320 }),
  .C2({ S1324 }),
  .ZN({ S1325 })
);
NAND3_X1 #() 
NAND3_X1_5226_ (
  .A1({ S1088 }),
  .A2({ S95 }),
  .A3({ S1051 }),
  .ZN({ S1326 })
);
NAND3_X1 #() 
NAND3_X1_5227_ (
  .A1({ S1067 }),
  .A2({ S25072 }),
  .A3({ S1326 }),
  .ZN({ S1327 })
);
OAI21_X1 #() 
OAI21_X1_2502_ (
  .A({ S95 }),
  .B1({ S103 }),
  .B2({ S1033 }),
  .ZN({ S1328 })
);
NAND2_X1 #() 
NAND2_X1_4844_ (
  .A1({ S1129 }),
  .A2({ S1328 }),
  .ZN({ S1329 })
);
NAND3_X1 #() 
NAND3_X1_5228_ (
  .A1({ S1329 }),
  .A2({ S1327 }),
  .A3({ S25957[925] }),
  .ZN({ S1330 })
);
NOR2_X1 #() 
NOR2_X1_1225_ (
  .A1({ S1088 }),
  .A2({ S25957[922] }),
  .ZN({ S1331 })
);
NOR2_X1 #() 
NOR2_X1_1226_ (
  .A1({ S1331 }),
  .A2({ S1105 }),
  .ZN({ S1332 })
);
NAND3_X1 #() 
NAND3_X1_5229_ (
  .A1({ S1039 }),
  .A2({ S95 }),
  .A3({ S1024 }),
  .ZN({ S1333 })
);
NAND3_X1 #() 
NAND3_X1_5230_ (
  .A1({ S1061 }),
  .A2({ S25072 }),
  .A3({ S1333 }),
  .ZN({ S1334 })
);
OAI211_X1 #() 
OAI211_X1_1675_ (
  .A({ S1334 }),
  .B({ S1084 }),
  .C1({ S1332 }),
  .C2({ S1301 }),
  .ZN({ S1335 })
);
NAND3_X1 #() 
NAND3_X1_5231_ (
  .A1({ S1335 }),
  .A2({ S25957[926] }),
  .A3({ S1330 }),
  .ZN({ S1336 })
);
NAND3_X1 #() 
NAND3_X1_5232_ (
  .A1({ S1325 }),
  .A2({ S25957[927] }),
  .A3({ S1336 }),
  .ZN({ S1337 })
);
NAND3_X1 #() 
NAND3_X1_5233_ (
  .A1({ S1310 }),
  .A2({ S25957[1092] }),
  .A3({ S1337 }),
  .ZN({ S1338 })
);
INV_X1 #() 
INV_X1_1571_ (
  .A({ S1338 }),
  .ZN({ S1339 })
);
AOI21_X1 #() 
AOI21_X1_2736_ (
  .A({ S25957[1092] }),
  .B1({ S1310 }),
  .B2({ S1337 }),
  .ZN({ S1340 })
);
OAI21_X1 #() 
OAI21_X1_2503_ (
  .A({ S25957[1028] }),
  .B1({ S1339 }),
  .B2({ S1340 }),
  .ZN({ S1341 })
);
INV_X1 #() 
INV_X1_1572_ (
  .A({ S1340 }),
  .ZN({ S1342 })
);
NAND3_X1 #() 
NAND3_X1_5234_ (
  .A1({ S1342 }),
  .A2({ S23396 }),
  .A3({ S1338 }),
  .ZN({ S1343 })
);
NAND2_X1 #() 
NAND2_X1_4845_ (
  .A1({ S1341 }),
  .A2({ S1343 }),
  .ZN({ S25957[772] })
);
NAND3_X1 #() 
NAND3_X1_5235_ (
  .A1({ S1044 }),
  .A2({ S95 }),
  .A3({ S1051 }),
  .ZN({ S1344 })
);
AOI22_X1 #() 
AOI22_X1_548_ (
  .A1({ S1075 }),
  .A2({ S1151 }),
  .B1({ S1344 }),
  .B2({ S1179 }),
  .ZN({ S1345 })
);
INV_X1 #() 
INV_X1_1573_ (
  .A({ S1055 }),
  .ZN({ S1346 })
);
NAND2_X1 #() 
NAND2_X1_4846_ (
  .A1({ S1090 }),
  .A2({ S95 }),
  .ZN({ S1347 })
);
NOR2_X1 #() 
NOR2_X1_1227_ (
  .A1({ S1347 }),
  .A2({ S25072 }),
  .ZN({ S1348 })
);
NOR2_X1 #() 
NOR2_X1_1228_ (
  .A1({ S1348 }),
  .A2({ S25957[925] }),
  .ZN({ S1349 })
);
OAI21_X1 #() 
OAI21_X1_2504_ (
  .A({ S1349 }),
  .B1({ S1346 }),
  .B2({ S1300 }),
  .ZN({ S1350 })
);
OAI211_X1 #() 
OAI211_X1_1676_ (
  .A({ S1350 }),
  .B({ S25957[926] }),
  .C1({ S1345 }),
  .C2({ S1084 }),
  .ZN({ S1351 })
);
AND2_X1 #() 
AND2_X1_298_ (
  .A1({ S1077 }),
  .A2({ S1163 }),
  .ZN({ S1352 })
);
NAND2_X1 #() 
NAND2_X1_4847_ (
  .A1({ S1051 }),
  .A2({ S25957[920] }),
  .ZN({ S1353 })
);
NAND2_X1 #() 
NAND2_X1_4848_ (
  .A1({ S1353 }),
  .A2({ S95 }),
  .ZN({ S1354 })
);
NAND3_X1 #() 
NAND3_X1_5236_ (
  .A1({ S1354 }),
  .A2({ S1299 }),
  .A3({ S1241 }),
  .ZN({ S1355 })
);
AOI21_X1 #() 
AOI21_X1_2737_ (
  .A({ S1084 }),
  .B1({ S1355 }),
  .B2({ S25072 }),
  .ZN({ S1356 })
);
OAI21_X1 #() 
OAI21_X1_2505_ (
  .A({ S1356 }),
  .B1({ S1352 }),
  .B2({ S25072 }),
  .ZN({ S1357 })
);
NAND2_X1 #() 
NAND2_X1_4849_ (
  .A1({ S1059 }),
  .A2({ S25957[920] }),
  .ZN({ S1358 })
);
NAND3_X1 #() 
NAND3_X1_5237_ (
  .A1({ S1358 }),
  .A2({ S25957[923] }),
  .A3({ S1039 }),
  .ZN({ S1359 })
);
INV_X1 #() 
INV_X1_1574_ (
  .A({ S1359 }),
  .ZN({ S1360 })
);
OAI21_X1 #() 
OAI21_X1_2506_ (
  .A({ S25072 }),
  .B1({ S1360 }),
  .B2({ S1049 }),
  .ZN({ S1361 })
);
NAND2_X1 #() 
NAND2_X1_4850_ (
  .A1({ S1091 }),
  .A2({ S1052 }),
  .ZN({ S1362 })
);
AOI21_X1 #() 
AOI21_X1_2738_ (
  .A({ S25072 }),
  .B1({ S1166 }),
  .B2({ S1030 }),
  .ZN({ S1363 })
);
NAND2_X1 #() 
NAND2_X1_4851_ (
  .A1({ S1362 }),
  .A2({ S1363 }),
  .ZN({ S1364 })
);
NAND3_X1 #() 
NAND3_X1_5238_ (
  .A1({ S1361 }),
  .A2({ S1084 }),
  .A3({ S1364 }),
  .ZN({ S1365 })
);
NAND3_X1 #() 
NAND3_X1_5239_ (
  .A1({ S1365 }),
  .A2({ S1021 }),
  .A3({ S1357 }),
  .ZN({ S1366 })
);
NAND3_X1 #() 
NAND3_X1_5240_ (
  .A1({ S1366 }),
  .A2({ S1351 }),
  .A3({ S24835 }),
  .ZN({ S1367 })
);
AOI21_X1 #() 
AOI21_X1_2739_ (
  .A({ S95 }),
  .B1({ S1047 }),
  .B2({ S25957[921] }),
  .ZN({ S1368 })
);
AOI21_X1 #() 
AOI21_X1_2740_ (
  .A({ S1368 }),
  .B1({ S1166 }),
  .B2({ S1048 }),
  .ZN({ S1369 })
);
NOR2_X1 #() 
NOR2_X1_1229_ (
  .A1({ S1369 }),
  .A2({ S25072 }),
  .ZN({ S1370 })
);
NAND2_X1 #() 
NAND2_X1_4852_ (
  .A1({ S1306 }),
  .A2({ S1027 }),
  .ZN({ S1371 })
);
NAND2_X1 #() 
NAND2_X1_4853_ (
  .A1({ S1371 }),
  .A2({ S1084 }),
  .ZN({ S1372 })
);
NOR2_X1 #() 
NOR2_X1_1230_ (
  .A1({ S1034 }),
  .A2({ S25957[923] }),
  .ZN({ S1373 })
);
NAND2_X1 #() 
NAND2_X1_4854_ (
  .A1({ S1044 }),
  .A2({ S1047 }),
  .ZN({ S1374 })
);
AOI22_X1 #() 
AOI22_X1_549_ (
  .A1({ S1161 }),
  .A2({ S1374 }),
  .B1({ S1373 }),
  .B2({ S1153 }),
  .ZN({ S1375 })
);
NAND3_X1 #() 
NAND3_X1_5241_ (
  .A1({ S1070 }),
  .A2({ S95 }),
  .A3({ S1044 }),
  .ZN({ S1376 })
);
NAND3_X1 #() 
NAND3_X1_5242_ (
  .A1({ S1376 }),
  .A2({ S25957[924] }),
  .A3({ S1297 }),
  .ZN({ S1377 })
);
OAI211_X1 #() 
OAI211_X1_1677_ (
  .A({ S1377 }),
  .B({ S25957[925] }),
  .C1({ S1375 }),
  .C2({ S25957[924] }),
  .ZN({ S1378 })
);
OAI211_X1 #() 
OAI211_X1_1678_ (
  .A({ S1378 }),
  .B({ S25957[926] }),
  .C1({ S1370 }),
  .C2({ S1372 }),
  .ZN({ S1379 })
);
NAND2_X1 #() 
NAND2_X1_4855_ (
  .A1({ S1027 }),
  .A2({ S95 }),
  .ZN({ S1380 })
);
OAI21_X1 #() 
OAI21_X1_2507_ (
  .A({ S25957[923] }),
  .B1({ S1231 }),
  .B2({ S1160 }),
  .ZN({ S1381 })
);
AOI21_X1 #() 
AOI21_X1_2741_ (
  .A({ S25957[924] }),
  .B1({ S1381 }),
  .B2({ S1380 }),
  .ZN({ S1382 })
);
INV_X1 #() 
INV_X1_1575_ (
  .A({ S1333 }),
  .ZN({ S1383 })
);
NAND2_X1 #() 
NAND2_X1_4856_ (
  .A1({ S1045 }),
  .A2({ S25957[923] }),
  .ZN({ S1384 })
);
NAND2_X1 #() 
NAND2_X1_4857_ (
  .A1({ S1384 }),
  .A2({ S25957[924] }),
  .ZN({ S1385 })
);
OAI21_X1 #() 
OAI21_X1_2508_ (
  .A({ S1084 }),
  .B1({ S1385 }),
  .B2({ S1383 }),
  .ZN({ S1386 })
);
AOI21_X1 #() 
AOI21_X1_2742_ (
  .A({ S25957[922] }),
  .B1({ S1044 }),
  .B2({ S1026 }),
  .ZN({ S1387 })
);
NAND3_X1 #() 
NAND3_X1_5243_ (
  .A1({ S1149 }),
  .A2({ S95 }),
  .A3({ S1047 }),
  .ZN({ S1388 })
);
OAI211_X1 #() 
OAI211_X1_1679_ (
  .A({ S1388 }),
  .B({ S25957[924] }),
  .C1({ S1387 }),
  .C2({ S1163 }),
  .ZN({ S1389 })
);
NAND3_X1 #() 
NAND3_X1_5244_ (
  .A1({ S1096 }),
  .A2({ S1222 }),
  .A3({ S1039 }),
  .ZN({ S1390 })
);
OAI211_X1 #() 
OAI211_X1_1680_ (
  .A({ S25072 }),
  .B({ S1390 }),
  .C1({ S1150 }),
  .C2({ S1125 }),
  .ZN({ S1391 })
);
NAND3_X1 #() 
NAND3_X1_5245_ (
  .A1({ S1389 }),
  .A2({ S1391 }),
  .A3({ S25957[925] }),
  .ZN({ S1392 })
);
OAI211_X1 #() 
OAI211_X1_1681_ (
  .A({ S1021 }),
  .B({ S1392 }),
  .C1({ S1386 }),
  .C2({ S1382 }),
  .ZN({ S1393 })
);
NAND3_X1 #() 
NAND3_X1_5246_ (
  .A1({ S1393 }),
  .A2({ S1379 }),
  .A3({ S25957[927] }),
  .ZN({ S1394 })
);
AOI21_X1 #() 
AOI21_X1_2743_ (
  .A({ S24445 }),
  .B1({ S1367 }),
  .B2({ S1394 }),
  .ZN({ S1395 })
);
INV_X1 #() 
INV_X1_1576_ (
  .A({ S24445 }),
  .ZN({ S25957[1091] })
);
OAI21_X1 #() 
OAI21_X1_2509_ (
  .A({ S1378 }),
  .B1({ S1370 }),
  .B2({ S1372 }),
  .ZN({ S1396 })
);
NAND2_X1 #() 
NAND2_X1_4858_ (
  .A1({ S1396 }),
  .A2({ S25957[926] }),
  .ZN({ S1397 })
);
NAND2_X1 #() 
NAND2_X1_4859_ (
  .A1({ S1389 }),
  .A2({ S1391 }),
  .ZN({ S1398 })
);
NAND2_X1 #() 
NAND2_X1_4860_ (
  .A1({ S1398 }),
  .A2({ S25957[925] }),
  .ZN({ S1399 })
);
NAND3_X1 #() 
NAND3_X1_5247_ (
  .A1({ S1381 }),
  .A2({ S25072 }),
  .A3({ S1380 }),
  .ZN({ S1400 })
);
NAND2_X1 #() 
NAND2_X1_4861_ (
  .A1({ S1384 }),
  .A2({ S1333 }),
  .ZN({ S1401 })
);
NAND2_X1 #() 
NAND2_X1_4862_ (
  .A1({ S1401 }),
  .A2({ S25957[924] }),
  .ZN({ S1402 })
);
NAND3_X1 #() 
NAND3_X1_5248_ (
  .A1({ S1400 }),
  .A2({ S1402 }),
  .A3({ S1084 }),
  .ZN({ S1403 })
);
NAND3_X1 #() 
NAND3_X1_5249_ (
  .A1({ S1403 }),
  .A2({ S1399 }),
  .A3({ S1021 }),
  .ZN({ S1404 })
);
NAND3_X1 #() 
NAND3_X1_5250_ (
  .A1({ S1397 }),
  .A2({ S1404 }),
  .A3({ S25957[927] }),
  .ZN({ S1405 })
);
NAND2_X1 #() 
NAND2_X1_4863_ (
  .A1({ S1075 }),
  .A2({ S1151 }),
  .ZN({ S1406 })
);
AOI21_X1 #() 
AOI21_X1_2744_ (
  .A({ S1084 }),
  .B1({ S1179 }),
  .B2({ S1344 }),
  .ZN({ S1407 })
);
NAND2_X1 #() 
NAND2_X1_4864_ (
  .A1({ S1406 }),
  .A2({ S1407 }),
  .ZN({ S1408 })
);
NAND2_X1 #() 
NAND2_X1_4865_ (
  .A1({ S1203 }),
  .A2({ S1052 }),
  .ZN({ S1409 })
);
AOI21_X1 #() 
AOI21_X1_2745_ (
  .A({ S1348 }),
  .B1({ S1409 }),
  .B2({ S1055 }),
  .ZN({ S1410 })
);
OAI211_X1 #() 
OAI211_X1_1682_ (
  .A({ S1408 }),
  .B({ S25957[926] }),
  .C1({ S25957[925] }),
  .C2({ S1410 }),
  .ZN({ S1411 })
);
AOI21_X1 #() 
AOI21_X1_2746_ (
  .A({ S25957[925] }),
  .B1({ S1361 }),
  .B2({ S1364 }),
  .ZN({ S1412 })
);
NAND3_X1 #() 
NAND3_X1_5251_ (
  .A1({ S1077 }),
  .A2({ S25957[924] }),
  .A3({ S1163 }),
  .ZN({ S1413 })
);
OAI211_X1 #() 
OAI211_X1_1683_ (
  .A({ S1413 }),
  .B({ S25957[925] }),
  .C1({ S25957[924] }),
  .C2({ S1355 }),
  .ZN({ S1414 })
);
NAND2_X1 #() 
NAND2_X1_4866_ (
  .A1({ S1414 }),
  .A2({ S1021 }),
  .ZN({ S1415 })
);
OAI211_X1 #() 
OAI211_X1_1684_ (
  .A({ S1411 }),
  .B({ S24835 }),
  .C1({ S1412 }),
  .C2({ S1415 }),
  .ZN({ S1416 })
);
AOI21_X1 #() 
AOI21_X1_2747_ (
  .A({ S25957[1091] }),
  .B1({ S1405 }),
  .B2({ S1416 }),
  .ZN({ S1417 })
);
OAI21_X1 #() 
OAI21_X1_2510_ (
  .A({ S80 }),
  .B1({ S1417 }),
  .B2({ S1395 }),
  .ZN({ S1418 })
);
NAND3_X1 #() 
NAND3_X1_5252_ (
  .A1({ S1405 }),
  .A2({ S1416 }),
  .A3({ S25957[1091] }),
  .ZN({ S1419 })
);
NAND3_X1 #() 
NAND3_X1_5253_ (
  .A1({ S1367 }),
  .A2({ S24445 }),
  .A3({ S1394 }),
  .ZN({ S1420 })
);
NAND3_X1 #() 
NAND3_X1_5254_ (
  .A1({ S1419 }),
  .A2({ S1420 }),
  .A3({ S25957[1027] }),
  .ZN({ S1421 })
);
NAND2_X1 #() 
NAND2_X1_4867_ (
  .A1({ S1418 }),
  .A2({ S1421 }),
  .ZN({ S104 })
);
INV_X1 #() 
INV_X1_1577_ (
  .A({ S104 }),
  .ZN({ S25957[771] })
);
INV_X1 #() 
INV_X1_1578_ (
  .A({ S24456 }),
  .ZN({ S25957[1088] })
);
OAI211_X1 #() 
OAI211_X1_1685_ (
  .A({ S25072 }),
  .B({ S1409 }),
  .C1({ S1091 }),
  .C2({ S25957[923] }),
  .ZN({ S1422 })
);
OAI211_X1 #() 
OAI211_X1_1686_ (
  .A({ S1120 }),
  .B({ S25957[924] }),
  .C1({ S95 }),
  .C2({ S1199 }),
  .ZN({ S1423 })
);
NAND3_X1 #() 
NAND3_X1_5255_ (
  .A1({ S1422 }),
  .A2({ S1423 }),
  .A3({ S25957[925] }),
  .ZN({ S1424 })
);
NAND4_X1 #() 
NAND4_X1_567_ (
  .A1({ S1044 }),
  .A2({ S1026 }),
  .A3({ S25957[923] }),
  .A4({ S25957[922] }),
  .ZN({ S1425 })
);
AOI21_X1 #() 
AOI21_X1_2748_ (
  .A({ S25072 }),
  .B1({ S1318 }),
  .B2({ S1425 }),
  .ZN({ S1426 })
);
OAI21_X1 #() 
OAI21_X1_2511_ (
  .A({ S1084 }),
  .B1({ S1426 }),
  .B2({ S1225 }),
  .ZN({ S1427 })
);
NAND3_X1 #() 
NAND3_X1_5256_ (
  .A1({ S1427 }),
  .A2({ S1424 }),
  .A3({ S25957[926] }),
  .ZN({ S1428 })
);
OAI211_X1 #() 
OAI211_X1_1687_ (
  .A({ S1322 }),
  .B({ S1328 }),
  .C1({ S1070 }),
  .C2({ S95 }),
  .ZN({ S1429 })
);
NAND2_X1 #() 
NAND2_X1_4868_ (
  .A1({ S1347 }),
  .A2({ S1163 }),
  .ZN({ S1430 })
);
AOI21_X1 #() 
AOI21_X1_2749_ (
  .A({ S25072 }),
  .B1({ S1064 }),
  .B2({ S1088 }),
  .ZN({ S1431 })
);
AOI22_X1 #() 
AOI22_X1_550_ (
  .A1({ S1429 }),
  .A2({ S25072 }),
  .B1({ S1430 }),
  .B2({ S1431 }),
  .ZN({ S1432 })
);
NAND2_X1 #() 
NAND2_X1_4869_ (
  .A1({ S1030 }),
  .A2({ S25957[923] }),
  .ZN({ S1433 })
);
OAI211_X1 #() 
OAI211_X1_1688_ (
  .A({ S25957[924] }),
  .B({ S1433 }),
  .C1({ S1387 }),
  .C2({ S25957[923] }),
  .ZN({ S1434 })
);
NAND3_X1 #() 
NAND3_X1_5257_ (
  .A1({ S1199 }),
  .A2({ S95 }),
  .A3({ S1047 }),
  .ZN({ S1435 })
);
NAND2_X1 #() 
NAND2_X1_4870_ (
  .A1({ S1179 }),
  .A2({ S1435 }),
  .ZN({ S1436 })
);
NAND3_X1 #() 
NAND3_X1_5258_ (
  .A1({ S1434 }),
  .A2({ S1436 }),
  .A3({ S1084 }),
  .ZN({ S1437 })
);
OAI211_X1 #() 
OAI211_X1_1689_ (
  .A({ S1437 }),
  .B({ S1021 }),
  .C1({ S1432 }),
  .C2({ S1084 }),
  .ZN({ S1438 })
);
NAND3_X1 #() 
NAND3_X1_5259_ (
  .A1({ S1428 }),
  .A2({ S25957[927] }),
  .A3({ S1438 }),
  .ZN({ S1439 })
);
NAND2_X1 #() 
NAND2_X1_4871_ (
  .A1({ S1127 }),
  .A2({ S25072 }),
  .ZN({ S1440 })
);
NOR2_X1 #() 
NOR2_X1_1231_ (
  .A1({ S1170 }),
  .A2({ S1440 }),
  .ZN({ S1441 })
);
NAND3_X1 #() 
NAND3_X1_5260_ (
  .A1({ S1358 }),
  .A2({ S1149 }),
  .A3({ S1070 }),
  .ZN({ S1442 })
);
NAND3_X1 #() 
NAND3_X1_5261_ (
  .A1({ S1033 }),
  .A2({ S95 }),
  .A3({ S1019 }),
  .ZN({ S1443 })
);
NAND2_X1 #() 
NAND2_X1_4872_ (
  .A1({ S1068 }),
  .A2({ S1443 }),
  .ZN({ S1444 })
);
AOI21_X1 #() 
AOI21_X1_2750_ (
  .A({ S1444 }),
  .B1({ S1442 }),
  .B2({ S25957[923] }),
  .ZN({ S1445 })
);
OAI21_X1 #() 
OAI21_X1_2512_ (
  .A({ S25957[925] }),
  .B1({ S1445 }),
  .B2({ S1441 }),
  .ZN({ S1446 })
);
NAND2_X1 #() 
NAND2_X1_4873_ (
  .A1({ S1189 }),
  .A2({ S1088 }),
  .ZN({ S1447 })
);
NOR2_X1 #() 
NOR2_X1_1232_ (
  .A1({ S1117 }),
  .A2({ S25072 }),
  .ZN({ S1448 })
);
AOI21_X1 #() 
AOI21_X1_2751_ (
  .A({ S25957[925] }),
  .B1({ S1447 }),
  .B2({ S1448 }),
  .ZN({ S1449 })
);
OAI21_X1 #() 
OAI21_X1_2513_ (
  .A({ S1449 }),
  .B1({ S1288 }),
  .B2({ S1252 }),
  .ZN({ S1450 })
);
NAND3_X1 #() 
NAND3_X1_5262_ (
  .A1({ S1446 }),
  .A2({ S25957[926] }),
  .A3({ S1450 }),
  .ZN({ S1451 })
);
AOI21_X1 #() 
AOI21_X1_2752_ (
  .A({ S25957[923] }),
  .B1({ S1048 }),
  .B2({ S1024 }),
  .ZN({ S1452 })
);
NOR2_X1 #() 
NOR2_X1_1233_ (
  .A1({ S1385 }),
  .A2({ S1452 }),
  .ZN({ S1453 })
);
NAND3_X1 #() 
NAND3_X1_5263_ (
  .A1({ S1183 }),
  .A2({ S1239 }),
  .A3({ S25072 }),
  .ZN({ S1454 })
);
OAI211_X1 #() 
OAI211_X1_1690_ (
  .A({ S1297 }),
  .B({ S25957[924] }),
  .C1({ S1331 }),
  .C2({ S1115 }),
  .ZN({ S1455 })
);
NAND3_X1 #() 
NAND3_X1_5264_ (
  .A1({ S1455 }),
  .A2({ S1454 }),
  .A3({ S25957[925] }),
  .ZN({ S1456 })
);
AOI21_X1 #() 
AOI21_X1_2753_ (
  .A({ S25957[923] }),
  .B1({ S1118 }),
  .B2({ S1035 }),
  .ZN({ S1457 })
);
NAND4_X1 #() 
NAND4_X1_568_ (
  .A1({ S1044 }),
  .A2({ S1026 }),
  .A3({ S25957[923] }),
  .A4({ S1051 }),
  .ZN({ S1458 })
);
NAND2_X1 #() 
NAND2_X1_4874_ (
  .A1({ S1458 }),
  .A2({ S25072 }),
  .ZN({ S1459 })
);
OAI21_X1 #() 
OAI21_X1_2514_ (
  .A({ S1084 }),
  .B1({ S1459 }),
  .B2({ S1457 }),
  .ZN({ S1460 })
);
OAI211_X1 #() 
OAI211_X1_1691_ (
  .A({ S1021 }),
  .B({ S1456 }),
  .C1({ S1453 }),
  .C2({ S1460 }),
  .ZN({ S1461 })
);
NAND3_X1 #() 
NAND3_X1_5265_ (
  .A1({ S1451 }),
  .A2({ S1461 }),
  .A3({ S24835 }),
  .ZN({ S1462 })
);
NAND3_X1 #() 
NAND3_X1_5266_ (
  .A1({ S1439 }),
  .A2({ S25957[1088] }),
  .A3({ S1462 }),
  .ZN({ S1463 })
);
INV_X1 #() 
INV_X1_1579_ (
  .A({ S1047 }),
  .ZN({ S1464 })
);
OAI211_X1 #() 
OAI211_X1_1692_ (
  .A({ S1038 }),
  .B({ S95 }),
  .C1({ S1026 }),
  .C2({ S25957[922] }),
  .ZN({ S1465 })
);
OAI211_X1 #() 
OAI211_X1_1693_ (
  .A({ S1465 }),
  .B({ S25957[924] }),
  .C1({ S1076 }),
  .C2({ S1464 }),
  .ZN({ S1466 })
);
AOI21_X1 #() 
AOI21_X1_2754_ (
  .A({ S95 }),
  .B1({ S1016 }),
  .B2({ S25957[922] }),
  .ZN({ S1467 })
);
AOI21_X1 #() 
AOI21_X1_2755_ (
  .A({ S1252 }),
  .B1({ S1467 }),
  .B2({ S1096 }),
  .ZN({ S1468 })
);
OAI211_X1 #() 
OAI211_X1_1694_ (
  .A({ S1466 }),
  .B({ S1084 }),
  .C1({ S1468 }),
  .C2({ S25957[924] }),
  .ZN({ S1469 })
);
AOI21_X1 #() 
AOI21_X1_2756_ (
  .A({ S25957[924] }),
  .B1({ S95 }),
  .B2({ S1047 }),
  .ZN({ S1470 })
);
XNOR2_X1 #() 
XNOR2_X1_192_ (
  .A({ S1026 }),
  .B({ S25957[922] }),
  .ZN({ S1471 })
);
OAI21_X1 #() 
OAI21_X1_2515_ (
  .A({ S1470 }),
  .B1({ S1471 }),
  .B2({ S95 }),
  .ZN({ S1472 })
);
AOI21_X1 #() 
AOI21_X1_2757_ (
  .A({ S95 }),
  .B1({ S1073 }),
  .B2({ S1358 }),
  .ZN({ S1473 })
);
OAI211_X1 #() 
OAI211_X1_1695_ (
  .A({ S1472 }),
  .B({ S25957[925] }),
  .C1({ S1473 }),
  .C2({ S1444 }),
  .ZN({ S1474 })
);
NAND3_X1 #() 
NAND3_X1_5267_ (
  .A1({ S1474 }),
  .A2({ S25957[926] }),
  .A3({ S1469 }),
  .ZN({ S1475 })
);
AOI21_X1 #() 
AOI21_X1_2758_ (
  .A({ S25072 }),
  .B1({ S1045 }),
  .B2({ S25957[923] }),
  .ZN({ S1476 })
);
OAI21_X1 #() 
OAI21_X1_2516_ (
  .A({ S95 }),
  .B1({ S1231 }),
  .B2({ S1160 }),
  .ZN({ S1477 })
);
NAND3_X1 #() 
NAND3_X1_5268_ (
  .A1({ S1203 }),
  .A2({ S1064 }),
  .A3({ S1025 }),
  .ZN({ S1478 })
);
AOI21_X1 #() 
AOI21_X1_2759_ (
  .A({ S25957[924] }),
  .B1({ S1124 }),
  .B2({ S1060 }),
  .ZN({ S1479 })
);
AOI22_X1 #() 
AOI22_X1_551_ (
  .A1({ S1477 }),
  .A2({ S1476 }),
  .B1({ S1479 }),
  .B2({ S1478 }),
  .ZN({ S1480 })
);
NAND2_X1 #() 
NAND2_X1_4875_ (
  .A1({ S1183 }),
  .A2({ S1239 }),
  .ZN({ S1481 })
);
NAND2_X1 #() 
NAND2_X1_4876_ (
  .A1({ S1481 }),
  .A2({ S25072 }),
  .ZN({ S1482 })
);
AND3_X1 #() 
AND3_X1_199_ (
  .A1({ S1025 }),
  .A2({ S103 }),
  .A3({ S25957[923] }),
  .ZN({ S1483 })
);
OAI21_X1 #() 
OAI21_X1_2517_ (
  .A({ S25957[924] }),
  .B1({ S1483 }),
  .B2({ S1234 }),
  .ZN({ S1484 })
);
NAND3_X1 #() 
NAND3_X1_5269_ (
  .A1({ S1482 }),
  .A2({ S1484 }),
  .A3({ S25957[925] }),
  .ZN({ S1485 })
);
OAI211_X1 #() 
OAI211_X1_1696_ (
  .A({ S1485 }),
  .B({ S1021 }),
  .C1({ S1480 }),
  .C2({ S25957[925] }),
  .ZN({ S1486 })
);
NAND3_X1 #() 
NAND3_X1_5270_ (
  .A1({ S1486 }),
  .A2({ S1475 }),
  .A3({ S24835 }),
  .ZN({ S1487 })
);
AOI21_X1 #() 
AOI21_X1_2760_ (
  .A({ S25957[923] }),
  .B1({ S1374 }),
  .B2({ S1024 }),
  .ZN({ S1488 })
);
INV_X1 #() 
INV_X1_1580_ (
  .A({ S1425 }),
  .ZN({ S1489 })
);
OAI21_X1 #() 
OAI21_X1_2518_ (
  .A({ S25957[924] }),
  .B1({ S1488 }),
  .B2({ S1489 }),
  .ZN({ S1490 })
);
NAND2_X1 #() 
NAND2_X1_4877_ (
  .A1({ S1224 }),
  .A2({ S1223 }),
  .ZN({ S1491 })
);
AOI21_X1 #() 
AOI21_X1_2761_ (
  .A({ S25957[925] }),
  .B1({ S1491 }),
  .B2({ S25072 }),
  .ZN({ S1492 })
);
NAND2_X1 #() 
NAND2_X1_4878_ (
  .A1({ S1492 }),
  .A2({ S1490 }),
  .ZN({ S1493 })
);
AOI21_X1 #() 
AOI21_X1_2762_ (
  .A({ S25957[923] }),
  .B1({ S1054 }),
  .B2({ S1026 }),
  .ZN({ S1494 })
);
OAI21_X1 #() 
OAI21_X1_2519_ (
  .A({ S25072 }),
  .B1({ S1494 }),
  .B2({ S1300 }),
  .ZN({ S1495 })
);
NAND2_X1 #() 
NAND2_X1_4879_ (
  .A1({ S1096 }),
  .A2({ S1051 }),
  .ZN({ S1496 })
);
OAI22_X1 #() 
OAI22_X1_125_ (
  .A1({ S1496 }),
  .A2({ S1328 }),
  .B1({ S1199 }),
  .B2({ S95 }),
  .ZN({ S1497 })
);
NAND2_X1 #() 
NAND2_X1_4880_ (
  .A1({ S1497 }),
  .A2({ S25957[924] }),
  .ZN({ S1498 })
);
NAND3_X1 #() 
NAND3_X1_5271_ (
  .A1({ S1495 }),
  .A2({ S1498 }),
  .A3({ S25957[925] }),
  .ZN({ S1499 })
);
NAND3_X1 #() 
NAND3_X1_5272_ (
  .A1({ S1499 }),
  .A2({ S1493 }),
  .A3({ S25957[926] }),
  .ZN({ S1500 })
);
NAND2_X1 #() 
NAND2_X1_4881_ (
  .A1({ S1429 }),
  .A2({ S25072 }),
  .ZN({ S1501 })
);
AOI21_X1 #() 
AOI21_X1_2763_ (
  .A({ S1084 }),
  .B1({ S1430 }),
  .B2({ S1431 }),
  .ZN({ S1502 })
);
NAND2_X1 #() 
NAND2_X1_4882_ (
  .A1({ S1501 }),
  .A2({ S1502 }),
  .ZN({ S1503 })
);
NAND2_X1 #() 
NAND2_X1_4883_ (
  .A1({ S1434 }),
  .A2({ S1436 }),
  .ZN({ S1504 })
);
NAND2_X1 #() 
NAND2_X1_4884_ (
  .A1({ S1504 }),
  .A2({ S1084 }),
  .ZN({ S1505 })
);
NAND3_X1 #() 
NAND3_X1_5273_ (
  .A1({ S1505 }),
  .A2({ S1503 }),
  .A3({ S1021 }),
  .ZN({ S1506 })
);
NAND3_X1 #() 
NAND3_X1_5274_ (
  .A1({ S1500 }),
  .A2({ S25957[927] }),
  .A3({ S1506 }),
  .ZN({ S1507 })
);
NAND3_X1 #() 
NAND3_X1_5275_ (
  .A1({ S1507 }),
  .A2({ S1487 }),
  .A3({ S24456 }),
  .ZN({ S1508 })
);
AOI21_X1 #() 
AOI21_X1_2764_ (
  .A({ S25957[1024] }),
  .B1({ S1508 }),
  .B2({ S1463 }),
  .ZN({ S1509 })
);
AND3_X1 #() 
AND3_X1_200_ (
  .A1({ S1508 }),
  .A2({ S1463 }),
  .A3({ S25957[1024] }),
  .ZN({ S1510 })
);
NOR2_X1 #() 
NOR2_X1_1234_ (
  .A1({ S1510 }),
  .A2({ S1509 }),
  .ZN({ S25957[768] })
);
NOR2_X1 #() 
NOR2_X1_1235_ (
  .A1({ S19478 }),
  .A2({ S19482 }),
  .ZN({ S25957[1185] })
);
XNOR2_X1 #() 
XNOR2_X1_193_ (
  .A({ S24559 }),
  .B({ S25957[1185] }),
  .ZN({ S25957[1057] })
);
NAND2_X1 #() 
NAND2_X1_4885_ (
  .A1({ S24631 }),
  .A2({ S24634 }),
  .ZN({ S25957[961] })
);
NAND2_X1 #() 
NAND2_X1_4886_ (
  .A1({ S25957[961] }),
  .A2({ S25957[1057] }),
  .ZN({ S1511 })
);
INV_X1 #() 
INV_X1_1581_ (
  .A({ S1511 }),
  .ZN({ S1512 })
);
NOR2_X1 #() 
NOR2_X1_1236_ (
  .A1({ S25957[961] }),
  .A2({ S25957[1057] }),
  .ZN({ S1513 })
);
NOR2_X1 #() 
NOR2_X1_1237_ (
  .A1({ S1512 }),
  .A2({ S1513 }),
  .ZN({ S25957[929] })
);
AOI21_X1 #() 
AOI21_X1_2765_ (
  .A({ S25072 }),
  .B1({ S1390 }),
  .B2({ S1326 }),
  .ZN({ S1514 })
);
OAI21_X1 #() 
OAI21_X1_2520_ (
  .A({ S25957[925] }),
  .B1({ S1514 }),
  .B2({ S1055 }),
  .ZN({ S1515 })
);
NAND3_X1 #() 
NAND3_X1_5276_ (
  .A1({ S1177 }),
  .A2({ S25072 }),
  .A3({ S1094 }),
  .ZN({ S1516 })
);
NAND4_X1 #() 
NAND4_X1_569_ (
  .A1({ S1333 }),
  .A2({ S1106 }),
  .A3({ S1105 }),
  .A4({ S25957[924] }),
  .ZN({ S1517 })
);
NAND3_X1 #() 
NAND3_X1_5277_ (
  .A1({ S1517 }),
  .A2({ S1516 }),
  .A3({ S1084 }),
  .ZN({ S1518 })
);
NAND3_X1 #() 
NAND3_X1_5278_ (
  .A1({ S1515 }),
  .A2({ S1021 }),
  .A3({ S1518 }),
  .ZN({ S1519 })
);
AND3_X1 #() 
AND3_X1_201_ (
  .A1({ S1054 }),
  .A2({ S1026 }),
  .A3({ S1052 }),
  .ZN({ S1520 })
);
OAI21_X1 #() 
OAI21_X1_2521_ (
  .A({ S25957[924] }),
  .B1({ S1328 }),
  .B2({ S1331 }),
  .ZN({ S1521 })
);
OAI21_X1 #() 
OAI21_X1_2522_ (
  .A({ S1096 }),
  .B1({ S1160 }),
  .B2({ S25957[920] }),
  .ZN({ S1522 })
);
AOI21_X1 #() 
AOI21_X1_2766_ (
  .A({ S1084 }),
  .B1({ S1522 }),
  .B2({ S1268 }),
  .ZN({ S1523 })
);
OAI21_X1 #() 
OAI21_X1_2523_ (
  .A({ S1523 }),
  .B1({ S1520 }),
  .B2({ S1521 }),
  .ZN({ S1524 })
);
INV_X1 #() 
INV_X1_1582_ (
  .A({ S1227 }),
  .ZN({ S1525 })
);
OAI21_X1 #() 
OAI21_X1_2524_ (
  .A({ S25957[924] }),
  .B1({ S1525 }),
  .B2({ S1103 }),
  .ZN({ S1526 })
);
NAND3_X1 #() 
NAND3_X1_5279_ (
  .A1({ S1143 }),
  .A2({ S25072 }),
  .A3({ S1425 }),
  .ZN({ S1527 })
);
OAI211_X1 #() 
OAI211_X1_1697_ (
  .A({ S1527 }),
  .B({ S1084 }),
  .C1({ S1473 }),
  .C2({ S1526 }),
  .ZN({ S1528 })
);
NAND3_X1 #() 
NAND3_X1_5280_ (
  .A1({ S1528 }),
  .A2({ S25957[926] }),
  .A3({ S1524 }),
  .ZN({ S1529 })
);
NAND3_X1 #() 
NAND3_X1_5281_ (
  .A1({ S1529 }),
  .A2({ S1519 }),
  .A3({ S24835 }),
  .ZN({ S1530 })
);
AOI21_X1 #() 
AOI21_X1_2767_ (
  .A({ S95 }),
  .B1({ S1048 }),
  .B2({ S1047 }),
  .ZN({ S1531 })
);
NAND2_X1 #() 
NAND2_X1_4887_ (
  .A1({ S1169 }),
  .A2({ S25957[923] }),
  .ZN({ S1532 })
);
NAND3_X1 #() 
NAND3_X1_5282_ (
  .A1({ S1532 }),
  .A2({ S1344 }),
  .A3({ S25072 }),
  .ZN({ S1533 })
);
OAI211_X1 #() 
OAI211_X1_1698_ (
  .A({ S1533 }),
  .B({ S25957[925] }),
  .C1({ S1531 }),
  .C2({ S1023 }),
  .ZN({ S1534 })
);
AOI21_X1 #() 
AOI21_X1_2768_ (
  .A({ S25957[925] }),
  .B1({ S1465 }),
  .B2({ S1156 }),
  .ZN({ S1535 })
);
OAI21_X1 #() 
OAI21_X1_2525_ (
  .A({ S1535 }),
  .B1({ S1046 }),
  .B2({ S1315 }),
  .ZN({ S1536 })
);
NAND3_X1 #() 
NAND3_X1_5283_ (
  .A1({ S1534 }),
  .A2({ S1536 }),
  .A3({ S1021 }),
  .ZN({ S1537 })
);
OAI21_X1 #() 
OAI21_X1_2526_ (
  .A({ S1431 }),
  .B1({ S1231 }),
  .B2({ S1190 }),
  .ZN({ S1538 })
);
NOR2_X1 #() 
NOR2_X1_1238_ (
  .A1({ S1024 }),
  .A2({ S25957[920] }),
  .ZN({ S1539 })
);
NAND3_X1 #() 
NAND3_X1_5284_ (
  .A1({ S1039 }),
  .A2({ S1016 }),
  .A3({ S25957[923] }),
  .ZN({ S1540 })
);
OAI211_X1 #() 
OAI211_X1_1699_ (
  .A({ S1540 }),
  .B({ S25072 }),
  .C1({ S1347 }),
  .C2({ S1539 }),
  .ZN({ S1541 })
);
NAND3_X1 #() 
NAND3_X1_5285_ (
  .A1({ S1538 }),
  .A2({ S1084 }),
  .A3({ S1541 }),
  .ZN({ S1542 })
);
NAND2_X1 #() 
NAND2_X1_4888_ (
  .A1({ S1464 }),
  .A2({ S25957[923] }),
  .ZN({ S1543 })
);
NAND4_X1 #() 
NAND4_X1_570_ (
  .A1({ S1543 }),
  .A2({ S1040 }),
  .A3({ S1105 }),
  .A4({ S25957[924] }),
  .ZN({ S1544 })
);
OAI21_X1 #() 
OAI21_X1_2527_ (
  .A({ S25072 }),
  .B1({ S1255 }),
  .B2({ S25957[923] }),
  .ZN({ S1545 })
);
OAI211_X1 #() 
OAI211_X1_1700_ (
  .A({ S1544 }),
  .B({ S25957[925] }),
  .C1({ S1473 }),
  .C2({ S1545 }),
  .ZN({ S1546 })
);
NAND3_X1 #() 
NAND3_X1_5286_ (
  .A1({ S1546 }),
  .A2({ S1542 }),
  .A3({ S25957[926] }),
  .ZN({ S1547 })
);
NAND3_X1 #() 
NAND3_X1_5287_ (
  .A1({ S1547 }),
  .A2({ S25957[927] }),
  .A3({ S1537 }),
  .ZN({ S1548 })
);
AND3_X1 #() 
AND3_X1_202_ (
  .A1({ S1548 }),
  .A2({ S1530 }),
  .A3({ S25957[1089] }),
  .ZN({ S1549 })
);
AOI21_X1 #() 
AOI21_X1_2769_ (
  .A({ S25957[1089] }),
  .B1({ S1548 }),
  .B2({ S1530 }),
  .ZN({ S1550 })
);
OAI21_X1 #() 
OAI21_X1_2528_ (
  .A({ S25957[929] }),
  .B1({ S1549 }),
  .B2({ S1550 }),
  .ZN({ S1551 })
);
INV_X1 #() 
INV_X1_1583_ (
  .A({ S25957[929] }),
  .ZN({ S1552 })
);
NAND3_X1 #() 
NAND3_X1_5288_ (
  .A1({ S1548 }),
  .A2({ S1530 }),
  .A3({ S25957[1089] }),
  .ZN({ S1553 })
);
NAND2_X1 #() 
NAND2_X1_4889_ (
  .A1({ S1548 }),
  .A2({ S1530 }),
  .ZN({ S1554 })
);
NAND2_X1 #() 
NAND2_X1_4890_ (
  .A1({ S1554 }),
  .A2({ S24559 }),
  .ZN({ S1555 })
);
NAND3_X1 #() 
NAND3_X1_5289_ (
  .A1({ S1555 }),
  .A2({ S1552 }),
  .A3({ S1553 }),
  .ZN({ S1556 })
);
NAND3_X1 #() 
NAND3_X1_5290_ (
  .A1({ S1551 }),
  .A2({ S1556 }),
  .A3({ S25957[897] }),
  .ZN({ S1557 })
);
NAND3_X1 #() 
NAND3_X1_5291_ (
  .A1({ S1555 }),
  .A2({ S25957[929] }),
  .A3({ S1553 }),
  .ZN({ S1558 })
);
OAI21_X1 #() 
OAI21_X1_2529_ (
  .A({ S1552 }),
  .B1({ S1549 }),
  .B2({ S1550 }),
  .ZN({ S1559 })
);
NAND3_X1 #() 
NAND3_X1_5292_ (
  .A1({ S1559 }),
  .A2({ S1558 }),
  .A3({ S490 }),
  .ZN({ S1560 })
);
NAND2_X1 #() 
NAND2_X1_4891_ (
  .A1({ S1557 }),
  .A2({ S1560 }),
  .ZN({ S25957[769] })
);
NAND2_X1 #() 
NAND2_X1_4892_ (
  .A1({ S19535 }),
  .A2({ S19533 }),
  .ZN({ S25957[1186] })
);
NAND2_X1 #() 
NAND2_X1_4893_ (
  .A1({ S22032 }),
  .A2({ S22033 }),
  .ZN({ S25957[1090] })
);
XOR2_X1 #() 
XOR2_X1_78_ (
  .A({ S25957[1090] }),
  .B({ S25957[1186] }),
  .Z({ S25957[1058] })
);
NAND2_X1 #() 
NAND2_X1_4894_ (
  .A1({ S22029 }),
  .A2({ S22028 }),
  .ZN({ S25957[1122] })
);
NAND3_X1 #() 
NAND3_X1_5293_ (
  .A1({ S24682 }),
  .A2({ S25957[1122] }),
  .A3({ S24660 }),
  .ZN({ S1561 })
);
NAND4_X1 #() 
NAND4_X1_571_ (
  .A1({ S24719 }),
  .A2({ S24697 }),
  .A3({ S22029 }),
  .A4({ S22028 }),
  .ZN({ S1562 })
);
NAND2_X1 #() 
NAND2_X1_4895_ (
  .A1({ S1562 }),
  .A2({ S1561 }),
  .ZN({ S1563 })
);
NAND2_X1 #() 
NAND2_X1_4896_ (
  .A1({ S1182 }),
  .A2({ S95 }),
  .ZN({ S1564 })
);
NAND3_X1 #() 
NAND3_X1_5294_ (
  .A1({ S1149 }),
  .A2({ S25957[923] }),
  .A3({ S1026 }),
  .ZN({ S1565 })
);
AOI21_X1 #() 
AOI21_X1_2770_ (
  .A({ S25957[924] }),
  .B1({ S1565 }),
  .B2({ S1564 }),
  .ZN({ S1566 })
);
NAND3_X1 #() 
NAND3_X1_5295_ (
  .A1({ S25957[923] }),
  .A2({ S1024 }),
  .A3({ S25957[920] }),
  .ZN({ S1567 })
);
AOI21_X1 #() 
AOI21_X1_2771_ (
  .A({ S25072 }),
  .B1({ S1177 }),
  .B2({ S1567 }),
  .ZN({ S1568 })
);
OAI21_X1 #() 
OAI21_X1_2530_ (
  .A({ S25957[925] }),
  .B1({ S1566 }),
  .B2({ S1568 }),
  .ZN({ S1569 })
);
AOI21_X1 #() 
AOI21_X1_2772_ (
  .A({ S25072 }),
  .B1({ S1096 }),
  .B2({ S1222 }),
  .ZN({ S1570 })
);
NAND2_X1 #() 
NAND2_X1_4897_ (
  .A1({ S1570 }),
  .A2({ S1189 }),
  .ZN({ S1571 })
);
OAI211_X1 #() 
OAI211_X1_1701_ (
  .A({ S1571 }),
  .B({ S1084 }),
  .C1({ S1195 }),
  .C2({ S25957[924] }),
  .ZN({ S1572 })
);
NAND3_X1 #() 
NAND3_X1_5296_ (
  .A1({ S1569 }),
  .A2({ S1572 }),
  .A3({ S1021 }),
  .ZN({ S1573 })
);
NAND2_X1 #() 
NAND2_X1_4898_ (
  .A1({ S1053 }),
  .A2({ S25957[924] }),
  .ZN({ S1574 })
);
NAND3_X1 #() 
NAND3_X1_5297_ (
  .A1({ S1273 }),
  .A2({ S25957[923] }),
  .A3({ S1199 }),
  .ZN({ S1575 })
);
NAND2_X1 #() 
NAND2_X1_4899_ (
  .A1({ S1575 }),
  .A2({ S1242 }),
  .ZN({ S1576 })
);
OAI211_X1 #() 
OAI211_X1_1702_ (
  .A({ S1576 }),
  .B({ S25957[925] }),
  .C1({ S1494 }),
  .C2({ S1574 }),
  .ZN({ S1577 })
);
NOR2_X1 #() 
NOR2_X1_1239_ (
  .A1({ S1034 }),
  .A2({ S1033 }),
  .ZN({ S1578 })
);
NOR3_X1 #() 
NOR3_X1_162_ (
  .A1({ S1387 }),
  .A2({ S1578 }),
  .A3({ S95 }),
  .ZN({ S1579 })
);
NAND3_X1 #() 
NAND3_X1_5298_ (
  .A1({ S1061 }),
  .A2({ S25072 }),
  .A3({ S1443 }),
  .ZN({ S1580 })
);
OAI211_X1 #() 
OAI211_X1_1703_ (
  .A({ S1580 }),
  .B({ S1084 }),
  .C1({ S1579 }),
  .C2({ S1275 }),
  .ZN({ S1581 })
);
NAND3_X1 #() 
NAND3_X1_5299_ (
  .A1({ S1577 }),
  .A2({ S1581 }),
  .A3({ S25957[926] }),
  .ZN({ S1582 })
);
NAND3_X1 #() 
NAND3_X1_5300_ (
  .A1({ S1582 }),
  .A2({ S1573 }),
  .A3({ S25957[927] }),
  .ZN({ S1583 })
);
OAI21_X1 #() 
OAI21_X1_2531_ (
  .A({ S25072 }),
  .B1({ S1353 }),
  .B2({ S25957[923] }),
  .ZN({ S1584 })
);
AOI21_X1 #() 
AOI21_X1_2773_ (
  .A({ S1093 }),
  .B1({ S95 }),
  .B2({ S1024 }),
  .ZN({ S1585 })
);
OAI21_X1 #() 
OAI21_X1_2532_ (
  .A({ S25957[924] }),
  .B1({ S1585 }),
  .B2({ S1154 }),
  .ZN({ S1586 })
);
OAI211_X1 #() 
OAI211_X1_1704_ (
  .A({ S1586 }),
  .B({ S25957[925] }),
  .C1({ S1099 }),
  .C2({ S1584 }),
  .ZN({ S1587 })
);
INV_X1 #() 
INV_X1_1584_ (
  .A({ S1193 }),
  .ZN({ S1588 })
);
OAI211_X1 #() 
OAI211_X1_1705_ (
  .A({ S1024 }),
  .B({ S1047 }),
  .C1({ S1034 }),
  .C2({ S1033 }),
  .ZN({ S1589 })
);
AOI22_X1 #() 
AOI22_X1_552_ (
  .A1({ S1589 }),
  .A2({ S95 }),
  .B1({ S1588 }),
  .B2({ S1052 }),
  .ZN({ S1590 })
);
AOI21_X1 #() 
AOI21_X1_2774_ (
  .A({ S25957[924] }),
  .B1({ S1096 }),
  .B2({ S1222 }),
  .ZN({ S1591 })
);
OAI21_X1 #() 
OAI21_X1_2533_ (
  .A({ S1591 }),
  .B1({ S1317 }),
  .B2({ S25957[923] }),
  .ZN({ S1592 })
);
OAI211_X1 #() 
OAI211_X1_1706_ (
  .A({ S1592 }),
  .B({ S1084 }),
  .C1({ S1590 }),
  .C2({ S25072 }),
  .ZN({ S1593 })
);
AND3_X1 #() 
AND3_X1_203_ (
  .A1({ S1593 }),
  .A2({ S1587 }),
  .A3({ S25957[926] }),
  .ZN({ S1594 })
);
OAI211_X1 #() 
OAI211_X1_1707_ (
  .A({ S1025 }),
  .B({ S25957[923] }),
  .C1({ S25957[920] }),
  .C2({ S1024 }),
  .ZN({ S1595 })
);
OAI211_X1 #() 
OAI211_X1_1708_ (
  .A({ S1595 }),
  .B({ S25957[924] }),
  .C1({ S1150 }),
  .C2({ S1125 }),
  .ZN({ S1596 })
);
NAND4_X1 #() 
NAND4_X1_572_ (
  .A1({ S1227 }),
  .A2({ S1047 }),
  .A3({ S1024 }),
  .A4({ S25957[923] }),
  .ZN({ S1597 })
);
NAND3_X1 #() 
NAND3_X1_5301_ (
  .A1({ S1597 }),
  .A2({ S25072 }),
  .A3({ S1194 }),
  .ZN({ S1598 })
);
NAND3_X1 #() 
NAND3_X1_5302_ (
  .A1({ S1596 }),
  .A2({ S25957[925] }),
  .A3({ S1598 }),
  .ZN({ S1599 })
);
OAI211_X1 #() 
OAI211_X1_1709_ (
  .A({ S95 }),
  .B({ S1026 }),
  .C1({ S1353 }),
  .C2({ S1117 }),
  .ZN({ S1600 })
);
OAI211_X1 #() 
OAI211_X1_1710_ (
  .A({ S25072 }),
  .B({ S1600 }),
  .C1({ S1471 }),
  .C2({ S95 }),
  .ZN({ S1601 })
);
NAND2_X1 #() 
NAND2_X1_4900_ (
  .A1({ S1311 }),
  .A2({ S1570 }),
  .ZN({ S1602 })
);
NAND3_X1 #() 
NAND3_X1_5303_ (
  .A1({ S1601 }),
  .A2({ S1084 }),
  .A3({ S1602 }),
  .ZN({ S1603 })
);
AOI21_X1 #() 
AOI21_X1_2775_ (
  .A({ S25957[926] }),
  .B1({ S1603 }),
  .B2({ S1599 }),
  .ZN({ S1604 })
);
OAI21_X1 #() 
OAI21_X1_2534_ (
  .A({ S24835 }),
  .B1({ S1594 }),
  .B2({ S1604 }),
  .ZN({ S1605 })
);
NAND3_X1 #() 
NAND3_X1_5304_ (
  .A1({ S1605 }),
  .A2({ S1563 }),
  .A3({ S1583 }),
  .ZN({ S1606 })
);
INV_X1 #() 
INV_X1_1585_ (
  .A({ S1563 }),
  .ZN({ S25957[994] })
);
AND3_X1 #() 
AND3_X1_204_ (
  .A1({ S1582 }),
  .A2({ S1573 }),
  .A3({ S25957[927] }),
  .ZN({ S1607 })
);
NAND3_X1 #() 
NAND3_X1_5305_ (
  .A1({ S1593 }),
  .A2({ S1587 }),
  .A3({ S25957[926] }),
  .ZN({ S1608 })
);
NAND2_X1 #() 
NAND2_X1_4901_ (
  .A1({ S1603 }),
  .A2({ S1599 }),
  .ZN({ S1609 })
);
NAND2_X1 #() 
NAND2_X1_4902_ (
  .A1({ S1609 }),
  .A2({ S1021 }),
  .ZN({ S1610 })
);
AOI21_X1 #() 
AOI21_X1_2776_ (
  .A({ S25957[927] }),
  .B1({ S1610 }),
  .B2({ S1608 }),
  .ZN({ S1611 })
);
OAI21_X1 #() 
OAI21_X1_2535_ (
  .A({ S25957[994] }),
  .B1({ S1611 }),
  .B2({ S1607 }),
  .ZN({ S1612 })
);
AOI21_X1 #() 
AOI21_X1_2777_ (
  .A({ S25957[1058] }),
  .B1({ S1612 }),
  .B2({ S1606 }),
  .ZN({ S1613 })
);
INV_X1 #() 
INV_X1_1586_ (
  .A({ S25957[1058] }),
  .ZN({ S1614 })
);
OAI21_X1 #() 
OAI21_X1_2536_ (
  .A({ S1563 }),
  .B1({ S1611 }),
  .B2({ S1607 }),
  .ZN({ S1615 })
);
NAND3_X1 #() 
NAND3_X1_5306_ (
  .A1({ S1605 }),
  .A2({ S25957[994] }),
  .A3({ S1583 }),
  .ZN({ S1616 })
);
AOI21_X1 #() 
AOI21_X1_2778_ (
  .A({ S1614 }),
  .B1({ S1615 }),
  .B2({ S1616 }),
  .ZN({ S1617 })
);
OAI21_X1 #() 
OAI21_X1_2537_ (
  .A({ S359 }),
  .B1({ S1613 }),
  .B2({ S1617 }),
  .ZN({ S1618 })
);
NAND3_X1 #() 
NAND3_X1_5307_ (
  .A1({ S1615 }),
  .A2({ S1614 }),
  .A3({ S1616 }),
  .ZN({ S1619 })
);
NAND3_X1 #() 
NAND3_X1_5308_ (
  .A1({ S1612 }),
  .A2({ S25957[1058] }),
  .A3({ S1606 }),
  .ZN({ S1620 })
);
NAND3_X1 #() 
NAND3_X1_5309_ (
  .A1({ S1619 }),
  .A2({ S1620 }),
  .A3({ S25957[898] }),
  .ZN({ S1621 })
);
NAND2_X1 #() 
NAND2_X1_4903_ (
  .A1({ S1618 }),
  .A2({ S1621 }),
  .ZN({ S25957[770] })
);
NAND2_X1 #() 
NAND2_X1_4904_ (
  .A1({ S25957[912] }),
  .A2({ S25957[913] }),
  .ZN({ S1622 })
);
INV_X1 #() 
INV_X1_1587_ (
  .A({ S1622 }),
  .ZN({ S105 })
);
NAND2_X1 #() 
NAND2_X1_4905_ (
  .A1({ S25921 }),
  .A2({ S264 }),
  .ZN({ S106 })
);
INV_X1 #() 
INV_X1_1588_ (
  .A({ S22148 }),
  .ZN({ S25957[1119] })
);
NAND3_X1 #() 
NAND3_X1_5310_ (
  .A1({ S25957[914] }),
  .A2({ S25919 }),
  .A3({ S25920 }),
  .ZN({ S1623 })
);
NAND4_X1 #() 
NAND4_X1_573_ (
  .A1({ S262 }),
  .A2({ S263 }),
  .A3({ S347 }),
  .A4({ S348 }),
  .ZN({ S1624 })
);
NAND2_X1 #() 
NAND2_X1_4906_ (
  .A1({ S1623 }),
  .A2({ S1624 }),
  .ZN({ S1625 })
);
INV_X1 #() 
INV_X1_1589_ (
  .A({ S1625 }),
  .ZN({ S1626 })
);
NAND3_X1 #() 
NAND3_X1_5311_ (
  .A1({ S349 }),
  .A2({ S23260 }),
  .A3({ S23271 }),
  .ZN({ S1627 })
);
AOI22_X1 #() 
AOI22_X1_553_ (
  .A1({ S23087 }),
  .A2({ S23088 }),
  .B1({ S262 }),
  .B2({ S263 }),
  .ZN({ S1628 })
);
AOI21_X1 #() 
AOI21_X1_2779_ (
  .A({ S25957[916] }),
  .B1({ S25957[912] }),
  .B2({ S1628 }),
  .ZN({ S1629 })
);
OAI211_X1 #() 
OAI211_X1_1711_ (
  .A({ S1629 }),
  .B({ S1626 }),
  .C1({ S1627 }),
  .C2({ S25957[912] }),
  .ZN({ S1630 })
);
NAND4_X1 #() 
NAND4_X1_574_ (
  .A1({ S23192 }),
  .A2({ S23204 }),
  .A3({ S262 }),
  .A4({ S263 }),
  .ZN({ S1631 })
);
NAND2_X1 #() 
NAND2_X1_4907_ (
  .A1({ S1631 }),
  .A2({ S86 }),
  .ZN({ S1632 })
);
INV_X1 #() 
INV_X1_1590_ (
  .A({ S1632 }),
  .ZN({ S1633 })
);
NAND2_X1 #() 
NAND2_X1_4908_ (
  .A1({ S1631 }),
  .A2({ S1627 }),
  .ZN({ S1634 })
);
NAND2_X1 #() 
NAND2_X1_4909_ (
  .A1({ S1634 }),
  .A2({ S25957[915] }),
  .ZN({ S1635 })
);
INV_X1 #() 
INV_X1_1591_ (
  .A({ S1635 }),
  .ZN({ S1636 })
);
OAI21_X1 #() 
OAI21_X1_2538_ (
  .A({ S25957[916] }),
  .B1({ S1636 }),
  .B2({ S1633 }),
  .ZN({ S1637 })
);
NAND3_X1 #() 
NAND3_X1_5312_ (
  .A1({ S1637 }),
  .A2({ S1630 }),
  .A3({ S25608 }),
  .ZN({ S1638 })
);
NAND3_X1 #() 
NAND3_X1_5313_ (
  .A1({ S25957[914] }),
  .A2({ S23192 }),
  .A3({ S23204 }),
  .ZN({ S1639 })
);
NAND3_X1 #() 
NAND3_X1_5314_ (
  .A1({ S25957[912] }),
  .A2({ S264 }),
  .A3({ S349 }),
  .ZN({ S1640 })
);
NAND3_X1 #() 
NAND3_X1_5315_ (
  .A1({ S1640 }),
  .A2({ S25957[915] }),
  .A3({ S1639 }),
  .ZN({ S1641 })
);
NAND3_X1 #() 
NAND3_X1_5316_ (
  .A1({ S23192 }),
  .A2({ S23204 }),
  .A3({ S349 }),
  .ZN({ S1642 })
);
NAND2_X1 #() 
NAND2_X1_4910_ (
  .A1({ S1642 }),
  .A2({ S86 }),
  .ZN({ S1643 })
);
OAI21_X1 #() 
OAI21_X1_2539_ (
  .A({ S1641 }),
  .B1({ S264 }),
  .B2({ S1643 }),
  .ZN({ S1644 })
);
NAND2_X1 #() 
NAND2_X1_4911_ (
  .A1({ S1644 }),
  .A2({ S25957[916] }),
  .ZN({ S1645 })
);
INV_X1 #() 
INV_X1_1592_ (
  .A({ S1627 }),
  .ZN({ S1646 })
);
NAND2_X1 #() 
NAND2_X1_4912_ (
  .A1({ S1631 }),
  .A2({ S1623 }),
  .ZN({ S1647 })
);
OAI21_X1 #() 
OAI21_X1_2540_ (
  .A({ S86 }),
  .B1({ S1647 }),
  .B2({ S1646 }),
  .ZN({ S1648 })
);
NAND4_X1 #() 
NAND4_X1_575_ (
  .A1({ S25920 }),
  .A2({ S25919 }),
  .A3({ S23260 }),
  .A4({ S23271 }),
  .ZN({ S1649 })
);
NAND3_X1 #() 
NAND3_X1_5317_ (
  .A1({ S25921 }),
  .A2({ S25957[913] }),
  .A3({ S25957[914] }),
  .ZN({ S1650 })
);
NAND3_X1 #() 
NAND3_X1_5318_ (
  .A1({ S1650 }),
  .A2({ S25957[915] }),
  .A3({ S1649 }),
  .ZN({ S1651 })
);
NAND3_X1 #() 
NAND3_X1_5319_ (
  .A1({ S1648 }),
  .A2({ S22985 }),
  .A3({ S1651 }),
  .ZN({ S1652 })
);
NAND3_X1 #() 
NAND3_X1_5320_ (
  .A1({ S1645 }),
  .A2({ S25957[917] }),
  .A3({ S1652 }),
  .ZN({ S1653 })
);
NAND3_X1 #() 
NAND3_X1_5321_ (
  .A1({ S1638 }),
  .A2({ S1653 }),
  .A3({ S25957[918] }),
  .ZN({ S1654 })
);
NAND4_X1 #() 
NAND4_X1_576_ (
  .A1({ S23260 }),
  .A2({ S23271 }),
  .A3({ S347 }),
  .A4({ S348 }),
  .ZN({ S1655 })
);
NAND2_X1 #() 
NAND2_X1_4913_ (
  .A1({ S1639 }),
  .A2({ S1655 }),
  .ZN({ S1656 })
);
NAND2_X1 #() 
NAND2_X1_4914_ (
  .A1({ S1656 }),
  .A2({ S106 }),
  .ZN({ S1657 })
);
NAND3_X1 #() 
NAND3_X1_5322_ (
  .A1({ S1649 }),
  .A2({ S1631 }),
  .A3({ S349 }),
  .ZN({ S1658 })
);
AOI21_X1 #() 
AOI21_X1_2780_ (
  .A({ S86 }),
  .B1({ S1657 }),
  .B2({ S1658 }),
  .ZN({ S1659 })
);
INV_X1 #() 
INV_X1_1593_ (
  .A({ S1624 }),
  .ZN({ S1660 })
);
NAND3_X1 #() 
NAND3_X1_5323_ (
  .A1({ S25920 }),
  .A2({ S25919 }),
  .A3({ S349 }),
  .ZN({ S1661 })
);
AND2_X1 #() 
AND2_X1_299_ (
  .A1({ S1661 }),
  .A2({ S86 }),
  .ZN({ S1662 })
);
INV_X1 #() 
INV_X1_1594_ (
  .A({ S1662 }),
  .ZN({ S1663 })
);
NOR2_X1 #() 
NOR2_X1_1240_ (
  .A1({ S1663 }),
  .A2({ S1660 }),
  .ZN({ S1664 })
);
OAI21_X1 #() 
OAI21_X1_2541_ (
  .A({ S25957[916] }),
  .B1({ S1664 }),
  .B2({ S1659 }),
  .ZN({ S1665 })
);
NAND2_X1 #() 
NAND2_X1_4915_ (
  .A1({ S1642 }),
  .A2({ S1627 }),
  .ZN({ S1666 })
);
AOI22_X1 #() 
AOI22_X1_554_ (
  .A1({ S1666 }),
  .A2({ S106 }),
  .B1({ S25957[914] }),
  .B2({ S1649 }),
  .ZN({ S1667 })
);
NAND2_X1 #() 
NAND2_X1_4916_ (
  .A1({ S1667 }),
  .A2({ S86 }),
  .ZN({ S1668 })
);
OAI21_X1 #() 
OAI21_X1_2542_ (
  .A({ S22985 }),
  .B1({ S86 }),
  .B2({ S1627 }),
  .ZN({ S1669 })
);
INV_X1 #() 
INV_X1_1595_ (
  .A({ S1669 }),
  .ZN({ S1670 })
);
NAND2_X1 #() 
NAND2_X1_4917_ (
  .A1({ S1668 }),
  .A2({ S1670 }),
  .ZN({ S1671 })
);
AOI21_X1 #() 
AOI21_X1_2781_ (
  .A({ S25957[917] }),
  .B1({ S1665 }),
  .B2({ S1671 }),
  .ZN({ S1672 })
);
NOR2_X1 #() 
NOR2_X1_1241_ (
  .A1({ S25957[915] }),
  .A2({ S264 }),
  .ZN({ S1673 })
);
NAND2_X1 #() 
NAND2_X1_4918_ (
  .A1({ S25957[915] }),
  .A2({ S264 }),
  .ZN({ S1674 })
);
AOI21_X1 #() 
AOI21_X1_2782_ (
  .A({ S349 }),
  .B1({ S23204 }),
  .B2({ S23192 }),
  .ZN({ S1675 })
);
NAND2_X1 #() 
NAND2_X1_4919_ (
  .A1({ S1675 }),
  .A2({ S25957[915] }),
  .ZN({ S1676 })
);
NAND3_X1 #() 
NAND3_X1_5324_ (
  .A1({ S1676 }),
  .A2({ S25957[916] }),
  .A3({ S1674 }),
  .ZN({ S1677 })
);
AOI21_X1 #() 
AOI21_X1_2783_ (
  .A({ S1677 }),
  .B1({ S1673 }),
  .B2({ S1623 }),
  .ZN({ S1678 })
);
AND2_X1 #() 
AND2_X1_300_ (
  .A1({ S1643 }),
  .A2({ S22985 }),
  .ZN({ S1679 })
);
NAND2_X1 #() 
NAND2_X1_4920_ (
  .A1({ S25957[915] }),
  .A2({ S25921 }),
  .ZN({ S1680 })
);
NAND2_X1 #() 
NAND2_X1_4921_ (
  .A1({ S1680 }),
  .A2({ S25957[913] }),
  .ZN({ S1681 })
);
AOI211_X1 #() 
AOI211_X1_86_ (
  .A({ S25608 }),
  .B({ S1678 }),
  .C1({ S1679 }),
  .C2({ S1681 }),
  .ZN({ S1682 })
);
OAI21_X1 #() 
OAI21_X1_2543_ (
  .A({ S22836 }),
  .B1({ S1682 }),
  .B2({ S1672 }),
  .ZN({ S1683 })
);
NAND3_X1 #() 
NAND3_X1_5325_ (
  .A1({ S1683 }),
  .A2({ S25957[919] }),
  .A3({ S1654 }),
  .ZN({ S1684 })
);
NAND2_X1 #() 
NAND2_X1_4922_ (
  .A1({ S22756 }),
  .A2({ S22755 }),
  .ZN({ S1685 })
);
NAND3_X1 #() 
NAND3_X1_5326_ (
  .A1({ S349 }),
  .A2({ S262 }),
  .A3({ S263 }),
  .ZN({ S1686 })
);
NOR2_X1 #() 
NOR2_X1_1242_ (
  .A1({ S1686 }),
  .A2({ S25921 }),
  .ZN({ S1687 })
);
NAND3_X1 #() 
NAND3_X1_5327_ (
  .A1({ S25921 }),
  .A2({ S264 }),
  .A3({ S25957[914] }),
  .ZN({ S1688 })
);
NAND2_X1 #() 
NAND2_X1_4923_ (
  .A1({ S1688 }),
  .A2({ S25957[915] }),
  .ZN({ S1689 })
);
NOR2_X1 #() 
NOR2_X1_1243_ (
  .A1({ S1689 }),
  .A2({ S1687 }),
  .ZN({ S1690 })
);
OAI21_X1 #() 
OAI21_X1_2544_ (
  .A({ S1642 }),
  .B1({ S1624 }),
  .B2({ S25957[912] }),
  .ZN({ S1691 })
);
OAI21_X1 #() 
OAI21_X1_2545_ (
  .A({ S25957[916] }),
  .B1({ S1691 }),
  .B2({ S25957[915] }),
  .ZN({ S1692 })
);
NAND2_X1 #() 
NAND2_X1_4924_ (
  .A1({ S1640 }),
  .A2({ S1624 }),
  .ZN({ S1693 })
);
NAND2_X1 #() 
NAND2_X1_4925_ (
  .A1({ S1693 }),
  .A2({ S25957[915] }),
  .ZN({ S1694 })
);
NAND3_X1 #() 
NAND3_X1_5328_ (
  .A1({ S1639 }),
  .A2({ S1655 }),
  .A3({ S86 }),
  .ZN({ S1695 })
);
NAND3_X1 #() 
NAND3_X1_5329_ (
  .A1({ S1694 }),
  .A2({ S22985 }),
  .A3({ S1695 }),
  .ZN({ S1696 })
);
OAI211_X1 #() 
OAI211_X1_1712_ (
  .A({ S1696 }),
  .B({ S25957[917] }),
  .C1({ S1690 }),
  .C2({ S1692 }),
  .ZN({ S1697 })
);
NOR2_X1 #() 
NOR2_X1_1244_ (
  .A1({ S1675 }),
  .A2({ S86 }),
  .ZN({ S1698 })
);
NAND2_X1 #() 
NAND2_X1_4926_ (
  .A1({ S1698 }),
  .A2({ S1686 }),
  .ZN({ S1699 })
);
NAND4_X1 #() 
NAND4_X1_577_ (
  .A1({ S1639 }),
  .A2({ S1642 }),
  .A3({ S1655 }),
  .A4({ S1686 }),
  .ZN({ S1700 })
);
AOI21_X1 #() 
AOI21_X1_2784_ (
  .A({ S25957[916] }),
  .B1({ S1700 }),
  .B2({ S86 }),
  .ZN({ S1701 })
);
INV_X1 #() 
INV_X1_1596_ (
  .A({ S1656 }),
  .ZN({ S1702 })
);
AOI21_X1 #() 
AOI21_X1_2785_ (
  .A({ S86 }),
  .B1({ S1702 }),
  .B2({ S1658 }),
  .ZN({ S1703 })
);
AOI21_X1 #() 
AOI21_X1_2786_ (
  .A({ S1703 }),
  .B1({ S1662 }),
  .B2({ S1657 }),
  .ZN({ S1704 })
);
AOI22_X1 #() 
AOI22_X1_555_ (
  .A1({ S1704 }),
  .A2({ S25957[916] }),
  .B1({ S1699 }),
  .B2({ S1701 }),
  .ZN({ S1705 })
);
OAI21_X1 #() 
OAI21_X1_2546_ (
  .A({ S1697 }),
  .B1({ S1705 }),
  .B2({ S25957[917] }),
  .ZN({ S1706 })
);
NAND3_X1 #() 
NAND3_X1_5330_ (
  .A1({ S1649 }),
  .A2({ S25957[915] }),
  .A3({ S1686 }),
  .ZN({ S1707 })
);
NAND2_X1 #() 
NAND2_X1_4927_ (
  .A1({ S1624 }),
  .A2({ S86 }),
  .ZN({ S1708 })
);
OR2_X1 #() 
OR2_X1_66_ (
  .A1({ S1666 }),
  .A2({ S1708 }),
  .ZN({ S1709 })
);
AND2_X1 #() 
AND2_X1_301_ (
  .A1({ S1709 }),
  .A2({ S1707 }),
  .ZN({ S1710 })
);
NAND2_X1 #() 
NAND2_X1_4928_ (
  .A1({ S86 }),
  .A2({ S25957[912] }),
  .ZN({ S1711 })
);
NAND2_X1 #() 
NAND2_X1_4929_ (
  .A1({ S1698 }),
  .A2({ S1627 }),
  .ZN({ S1712 })
);
NAND3_X1 #() 
NAND3_X1_5331_ (
  .A1({ S1712 }),
  .A2({ S25957[916] }),
  .A3({ S1711 }),
  .ZN({ S1713 })
);
OAI211_X1 #() 
OAI211_X1_1713_ (
  .A({ S25957[917] }),
  .B({ S1713 }),
  .C1({ S1710 }),
  .C2({ S25957[916] }),
  .ZN({ S1714 })
);
AOI21_X1 #() 
AOI21_X1_2787_ (
  .A({ S349 }),
  .B1({ S1649 }),
  .B2({ S1631 }),
  .ZN({ S1715 })
);
NOR2_X1 #() 
NOR2_X1_1245_ (
  .A1({ S1687 }),
  .A2({ S25957[915] }),
  .ZN({ S1716 })
);
INV_X1 #() 
INV_X1_1597_ (
  .A({ S1716 }),
  .ZN({ S1717 })
);
AOI21_X1 #() 
AOI21_X1_2788_ (
  .A({ S22985 }),
  .B1({ S1650 }),
  .B2({ S25957[915] }),
  .ZN({ S1718 })
);
OAI21_X1 #() 
OAI21_X1_2547_ (
  .A({ S1718 }),
  .B1({ S1717 }),
  .B2({ S1715 }),
  .ZN({ S1719 })
);
NAND2_X1 #() 
NAND2_X1_4930_ (
  .A1({ S1649 }),
  .A2({ S25957[914] }),
  .ZN({ S1720 })
);
NOR2_X1 #() 
NOR2_X1_1246_ (
  .A1({ S1632 }),
  .A2({ S1720 }),
  .ZN({ S1721 })
);
NAND2_X1 #() 
NAND2_X1_4931_ (
  .A1({ S25957[915] }),
  .A2({ S25957[914] }),
  .ZN({ S1722 })
);
OAI21_X1 #() 
OAI21_X1_2548_ (
  .A({ S22985 }),
  .B1({ S105 }),
  .B2({ S1722 }),
  .ZN({ S1723 })
);
OAI211_X1 #() 
OAI211_X1_1714_ (
  .A({ S1719 }),
  .B({ S25608 }),
  .C1({ S1721 }),
  .C2({ S1723 }),
  .ZN({ S1724 })
);
NAND3_X1 #() 
NAND3_X1_5332_ (
  .A1({ S1724 }),
  .A2({ S1714 }),
  .A3({ S22836 }),
  .ZN({ S1725 })
);
OAI211_X1 #() 
OAI211_X1_1715_ (
  .A({ S1685 }),
  .B({ S1725 }),
  .C1({ S1706 }),
  .C2({ S22836 }),
  .ZN({ S1726 })
);
NAND2_X1 #() 
NAND2_X1_4932_ (
  .A1({ S1684 }),
  .A2({ S1726 }),
  .ZN({ S1727 })
);
NAND2_X1 #() 
NAND2_X1_4933_ (
  .A1({ S1727 }),
  .A2({ S25957[1119] }),
  .ZN({ S1728 })
);
INV_X1 #() 
INV_X1_1598_ (
  .A({ S1728 }),
  .ZN({ S1729 })
);
NAND3_X1 #() 
NAND3_X1_5333_ (
  .A1({ S1684 }),
  .A2({ S1726 }),
  .A3({ S22148 }),
  .ZN({ S1730 })
);
INV_X1 #() 
INV_X1_1599_ (
  .A({ S1730 }),
  .ZN({ S1731 })
);
NOR2_X1 #() 
NOR2_X1_1247_ (
  .A1({ S1729 }),
  .A2({ S1731 }),
  .ZN({ S25957[863] })
);
NOR2_X1 #() 
NOR2_X1_1248_ (
  .A1({ S25957[863] }),
  .A2({ S25957[1055] }),
  .ZN({ S1732 })
);
INV_X1 #() 
INV_X1_1600_ (
  .A({ S25957[863] }),
  .ZN({ S1733 })
);
NOR2_X1 #() 
NOR2_X1_1249_ (
  .A1({ S1733 }),
  .A2({ S22150 }),
  .ZN({ S1734 })
);
NOR2_X1 #() 
NOR2_X1_1250_ (
  .A1({ S1734 }),
  .A2({ S1732 }),
  .ZN({ S25957[799] })
);
XOR2_X1 #() 
XOR2_X1_79_ (
  .A({ S24901 }),
  .B({ S25957[1150] }),
  .Z({ S25957[1022] })
);
INV_X1 #() 
INV_X1_1601_ (
  .A({ S25957[1022] }),
  .ZN({ S1735 })
);
AOI21_X1 #() 
AOI21_X1_2789_ (
  .A({ S86 }),
  .B1({ S1720 }),
  .B2({ S1661 }),
  .ZN({ S1736 })
);
NAND2_X1 #() 
NAND2_X1_4934_ (
  .A1({ S86 }),
  .A2({ S1627 }),
  .ZN({ S1737 })
);
AOI22_X1 #() 
AOI22_X1_556_ (
  .A1({ S23087 }),
  .A2({ S23088 }),
  .B1({ S23260 }),
  .B2({ S23271 }),
  .ZN({ S1738 })
);
AOI21_X1 #() 
AOI21_X1_2790_ (
  .A({ S22985 }),
  .B1({ S1738 }),
  .B2({ S349 }),
  .ZN({ S1739 })
);
OAI21_X1 #() 
OAI21_X1_2549_ (
  .A({ S1739 }),
  .B1({ S25957[912] }),
  .B2({ S1737 }),
  .ZN({ S1740 })
);
OAI21_X1 #() 
OAI21_X1_2550_ (
  .A({ S22985 }),
  .B1({ S1715 }),
  .B2({ S25957[915] }),
  .ZN({ S1741 })
);
OAI21_X1 #() 
OAI21_X1_2551_ (
  .A({ S1740 }),
  .B1({ S1741 }),
  .B2({ S1736 }),
  .ZN({ S1742 })
);
INV_X1 #() 
INV_X1_1602_ (
  .A({ S1647 }),
  .ZN({ S1743 })
);
NAND4_X1 #() 
NAND4_X1_578_ (
  .A1({ S1639 }),
  .A2({ S1661 }),
  .A3({ S1655 }),
  .A4({ S86 }),
  .ZN({ S1744 })
);
OAI211_X1 #() 
OAI211_X1_1716_ (
  .A({ S25957[916] }),
  .B({ S1744 }),
  .C1({ S1743 }),
  .C2({ S86 }),
  .ZN({ S1745 })
);
INV_X1 #() 
INV_X1_1603_ (
  .A({ S1745 }),
  .ZN({ S1746 })
);
NAND2_X1 #() 
NAND2_X1_4935_ (
  .A1({ S1661 }),
  .A2({ S25957[913] }),
  .ZN({ S1747 })
);
AOI21_X1 #() 
AOI21_X1_2791_ (
  .A({ S25957[916] }),
  .B1({ S1676 }),
  .B2({ S1747 }),
  .ZN({ S1748 })
);
OAI21_X1 #() 
OAI21_X1_2552_ (
  .A({ S25957[917] }),
  .B1({ S1746 }),
  .B2({ S1748 }),
  .ZN({ S1749 })
);
OAI21_X1 #() 
OAI21_X1_2553_ (
  .A({ S1749 }),
  .B1({ S25957[917] }),
  .B2({ S1742 }),
  .ZN({ S1750 })
);
OAI211_X1 #() 
OAI211_X1_1717_ (
  .A({ S1661 }),
  .B({ S1627 }),
  .C1({ S1624 }),
  .C2({ S25957[912] }),
  .ZN({ S1751 })
);
NAND2_X1 #() 
NAND2_X1_4936_ (
  .A1({ S1751 }),
  .A2({ S25957[915] }),
  .ZN({ S1752 })
);
AOI22_X1 #() 
AOI22_X1_557_ (
  .A1({ S1752 }),
  .A2({ S22985 }),
  .B1({ S86 }),
  .B2({ S1640 }),
  .ZN({ S1753 })
);
OAI21_X1 #() 
OAI21_X1_2554_ (
  .A({ S1753 }),
  .B1({ S22985 }),
  .B2({ S1694 }),
  .ZN({ S1754 })
);
INV_X1 #() 
INV_X1_1604_ (
  .A({ S1686 }),
  .ZN({ S1755 })
);
NAND2_X1 #() 
NAND2_X1_4937_ (
  .A1({ S1655 }),
  .A2({ S25957[915] }),
  .ZN({ S1756 })
);
INV_X1 #() 
INV_X1_1605_ (
  .A({ S1640 }),
  .ZN({ S1757 })
);
OAI221_X1 #() 
OAI221_X1_145_ (
  .A({ S22985 }),
  .B1({ S1756 }),
  .B2({ S1755 }),
  .C1({ S1757 }),
  .C2({ S1708 }),
  .ZN({ S1758 })
);
NAND3_X1 #() 
NAND3_X1_5334_ (
  .A1({ S1688 }),
  .A2({ S25957[915] }),
  .A3({ S1622 }),
  .ZN({ S1759 })
);
NAND3_X1 #() 
NAND3_X1_5335_ (
  .A1({ S1663 }),
  .A2({ S1759 }),
  .A3({ S25957[916] }),
  .ZN({ S1760 })
);
NAND3_X1 #() 
NAND3_X1_5336_ (
  .A1({ S1758 }),
  .A2({ S25957[917] }),
  .A3({ S1760 }),
  .ZN({ S1761 })
);
OAI21_X1 #() 
OAI21_X1_2555_ (
  .A({ S1761 }),
  .B1({ S1754 }),
  .B2({ S25957[917] }),
  .ZN({ S1762 })
);
MUX2_X1 #() 
MUX2_X1_20_ (
  .A({ S1762 }),
  .B({ S1750 }),
  .S({ S25957[918] }),
  .Z({ S1763 })
);
NAND3_X1 #() 
NAND3_X1_5337_ (
  .A1({ S1642 }),
  .A2({ S25957[915] }),
  .A3({ S1627 }),
  .ZN({ S1764 })
);
INV_X1 #() 
INV_X1_1606_ (
  .A({ S1764 }),
  .ZN({ S1765 })
);
NAND2_X1 #() 
NAND2_X1_4938_ (
  .A1({ S1765 }),
  .A2({ S106 }),
  .ZN({ S1766 })
);
NAND2_X1 #() 
NAND2_X1_4939_ (
  .A1({ S1639 }),
  .A2({ S86 }),
  .ZN({ S1767 })
);
INV_X1 #() 
INV_X1_1607_ (
  .A({ S1767 }),
  .ZN({ S1768 })
);
AOI21_X1 #() 
AOI21_X1_2792_ (
  .A({ S1736 }),
  .B1({ S1768 }),
  .B2({ S1658 }),
  .ZN({ S1769 })
);
AOI22_X1 #() 
AOI22_X1_558_ (
  .A1({ S1769 }),
  .A2({ S25957[916] }),
  .B1({ S1701 }),
  .B2({ S1766 }),
  .ZN({ S1770 })
);
INV_X1 #() 
INV_X1_1608_ (
  .A({ S1661 }),
  .ZN({ S1771 })
);
NOR2_X1 #() 
NOR2_X1_1251_ (
  .A1({ S1674 }),
  .A2({ S1771 }),
  .ZN({ S1772 })
);
NAND2_X1 #() 
NAND2_X1_4940_ (
  .A1({ S1772 }),
  .A2({ S1639 }),
  .ZN({ S1773 })
);
OAI211_X1 #() 
OAI211_X1_1718_ (
  .A({ S1773 }),
  .B({ S25957[916] }),
  .C1({ S1626 }),
  .C2({ S25957[915] }),
  .ZN({ S1774 })
);
OAI21_X1 #() 
OAI21_X1_2556_ (
  .A({ S22985 }),
  .B1({ S1636 }),
  .B2({ S1673 }),
  .ZN({ S1775 })
);
NAND3_X1 #() 
NAND3_X1_5338_ (
  .A1({ S1774 }),
  .A2({ S25957[917] }),
  .A3({ S1775 }),
  .ZN({ S1776 })
);
OAI211_X1 #() 
OAI211_X1_1719_ (
  .A({ S25957[918] }),
  .B({ S1776 }),
  .C1({ S1770 }),
  .C2({ S25957[917] }),
  .ZN({ S1777 })
);
NAND2_X1 #() 
NAND2_X1_4941_ (
  .A1({ S1650 }),
  .A2({ S1661 }),
  .ZN({ S1778 })
);
AOI22_X1 #() 
AOI22_X1_559_ (
  .A1({ S1778 }),
  .A2({ S25957[915] }),
  .B1({ S1768 }),
  .B2({ S1658 }),
  .ZN({ S1779 })
);
NAND2_X1 #() 
NAND2_X1_4942_ (
  .A1({ S1649 }),
  .A2({ S349 }),
  .ZN({ S1780 })
);
NOR2_X1 #() 
NOR2_X1_1252_ (
  .A1({ S1780 }),
  .A2({ S25957[915] }),
  .ZN({ S1781 })
);
OAI22_X1 #() 
OAI22_X1_126_ (
  .A1({ S1779 }),
  .A2({ S25957[916] }),
  .B1({ S1677 }),
  .B2({ S1781 }),
  .ZN({ S1782 })
);
NAND2_X1 #() 
NAND2_X1_4943_ (
  .A1({ S1738 }),
  .A2({ S25957[914] }),
  .ZN({ S1783 })
);
INV_X1 #() 
INV_X1_1609_ (
  .A({ S1642 }),
  .ZN({ S1784 })
);
NAND2_X1 #() 
NAND2_X1_4944_ (
  .A1({ S1673 }),
  .A2({ S1784 }),
  .ZN({ S1785 })
);
NAND2_X1 #() 
NAND2_X1_4945_ (
  .A1({ S1785 }),
  .A2({ S1783 }),
  .ZN({ S1786 })
);
OAI21_X1 #() 
OAI21_X1_2557_ (
  .A({ S25957[916] }),
  .B1({ S1786 }),
  .B2({ S1721 }),
  .ZN({ S1787 })
);
NAND3_X1 #() 
NAND3_X1_5339_ (
  .A1({ S25921 }),
  .A2({ S25957[913] }),
  .A3({ S349 }),
  .ZN({ S1788 })
);
NAND3_X1 #() 
NAND3_X1_5340_ (
  .A1({ S1788 }),
  .A2({ S25957[915] }),
  .A3({ S1655 }),
  .ZN({ S1789 })
);
NAND4_X1 #() 
NAND4_X1_579_ (
  .A1({ S25957[913] }),
  .A2({ S25957[914] }),
  .A3({ S25919 }),
  .A4({ S25920 }),
  .ZN({ S1790 })
);
NAND2_X1 #() 
NAND2_X1_4946_ (
  .A1({ S1790 }),
  .A2({ S106 }),
  .ZN({ S1791 })
);
NAND2_X1 #() 
NAND2_X1_4947_ (
  .A1({ S1791 }),
  .A2({ S86 }),
  .ZN({ S1792 })
);
NAND3_X1 #() 
NAND3_X1_5341_ (
  .A1({ S1792 }),
  .A2({ S22985 }),
  .A3({ S1789 }),
  .ZN({ S1793 })
);
NAND3_X1 #() 
NAND3_X1_5342_ (
  .A1({ S1787 }),
  .A2({ S25957[917] }),
  .A3({ S1793 }),
  .ZN({ S1794 })
);
OAI211_X1 #() 
OAI211_X1_1720_ (
  .A({ S1794 }),
  .B({ S22836 }),
  .C1({ S1782 }),
  .C2({ S25957[917] }),
  .ZN({ S1795 })
);
AOI21_X1 #() 
AOI21_X1_2793_ (
  .A({ S1685 }),
  .B1({ S1777 }),
  .B2({ S1795 }),
  .ZN({ S1796 })
);
AOI21_X1 #() 
AOI21_X1_2794_ (
  .A({ S1796 }),
  .B1({ S1763 }),
  .B2({ S1685 }),
  .ZN({ S1797 })
);
NAND2_X1 #() 
NAND2_X1_4948_ (
  .A1({ S1797 }),
  .A2({ S1735 }),
  .ZN({ S1798 })
);
OR2_X1 #() 
OR2_X1_67_ (
  .A1({ S1797 }),
  .A2({ S1735 }),
  .ZN({ S1799 })
);
NAND2_X1 #() 
NAND2_X1_4949_ (
  .A1({ S1799 }),
  .A2({ S1798 }),
  .ZN({ S25957[894] })
);
NAND2_X1 #() 
NAND2_X1_4950_ (
  .A1({ S25957[894] }),
  .A2({ S25957[990] }),
  .ZN({ S1800 })
);
INV_X1 #() 
INV_X1_1610_ (
  .A({ S25957[990] }),
  .ZN({ S1801 })
);
INV_X1 #() 
INV_X1_1611_ (
  .A({ S25957[894] }),
  .ZN({ S1802 })
);
NAND2_X1 #() 
NAND2_X1_4951_ (
  .A1({ S1802 }),
  .A2({ S1801 }),
  .ZN({ S1803 })
);
NAND2_X1 #() 
NAND2_X1_4952_ (
  .A1({ S1803 }),
  .A2({ S1800 }),
  .ZN({ S1804 })
);
INV_X1 #() 
INV_X1_1612_ (
  .A({ S1804 }),
  .ZN({ S25957[862] })
);
NAND2_X1 #() 
NAND2_X1_4953_ (
  .A1({ S25957[862] }),
  .A2({ S22219 }),
  .ZN({ S1805 })
);
NAND2_X1 #() 
NAND2_X1_4954_ (
  .A1({ S1804 }),
  .A2({ S25957[1054] }),
  .ZN({ S1806 })
);
NAND2_X1 #() 
NAND2_X1_4955_ (
  .A1({ S1805 }),
  .A2({ S1806 }),
  .ZN({ S25957[798] })
);
INV_X1 #() 
INV_X1_1613_ (
  .A({ S24903 }),
  .ZN({ S25957[1117] })
);
NOR2_X1 #() 
NOR2_X1_1253_ (
  .A1({ S1627 }),
  .A2({ S25957[912] }),
  .ZN({ S1807 })
);
OAI21_X1 #() 
OAI21_X1_2558_ (
  .A({ S25957[915] }),
  .B1({ S1715 }),
  .B2({ S1807 }),
  .ZN({ S1808 })
);
AOI21_X1 #() 
AOI21_X1_2795_ (
  .A({ S25957[916] }),
  .B1({ S1808 }),
  .B2({ S1717 }),
  .ZN({ S1809 })
);
NAND2_X1 #() 
NAND2_X1_4956_ (
  .A1({ S1666 }),
  .A2({ S106 }),
  .ZN({ S1810 })
);
NOR2_X1 #() 
NOR2_X1_1254_ (
  .A1({ S1810 }),
  .A2({ S86 }),
  .ZN({ S1811 })
);
NAND3_X1 #() 
NAND3_X1_5343_ (
  .A1({ S1661 }),
  .A2({ S86 }),
  .A3({ S264 }),
  .ZN({ S1812 })
);
NAND2_X1 #() 
NAND2_X1_4957_ (
  .A1({ S1812 }),
  .A2({ S25957[916] }),
  .ZN({ S1813 })
);
NOR2_X1 #() 
NOR2_X1_1255_ (
  .A1({ S1811 }),
  .A2({ S1813 }),
  .ZN({ S1814 })
);
OAI21_X1 #() 
OAI21_X1_2559_ (
  .A({ S25608 }),
  .B1({ S1809 }),
  .B2({ S1814 }),
  .ZN({ S1815 })
);
NAND3_X1 #() 
NAND3_X1_5344_ (
  .A1({ S1622 }),
  .A2({ S86 }),
  .A3({ S1642 }),
  .ZN({ S1816 })
);
OAI211_X1 #() 
OAI211_X1_1721_ (
  .A({ S1816 }),
  .B({ S25957[916] }),
  .C1({ S1700 }),
  .C2({ S86 }),
  .ZN({ S1817 })
);
INV_X1 #() 
INV_X1_1614_ (
  .A({ S1631 }),
  .ZN({ S1818 })
);
NOR2_X1 #() 
NOR2_X1_1256_ (
  .A1({ S1818 }),
  .A2({ S1737 }),
  .ZN({ S1819 })
);
INV_X1 #() 
INV_X1_1615_ (
  .A({ S1819 }),
  .ZN({ S1820 })
);
NOR2_X1 #() 
NOR2_X1_1257_ (
  .A1({ S25957[916] }),
  .A2({ S1628 }),
  .ZN({ S1821 })
);
NAND2_X1 #() 
NAND2_X1_4958_ (
  .A1({ S1820 }),
  .A2({ S1821 }),
  .ZN({ S1822 })
);
NAND3_X1 #() 
NAND3_X1_5345_ (
  .A1({ S1822 }),
  .A2({ S25957[917] }),
  .A3({ S1817 }),
  .ZN({ S1823 })
);
NAND3_X1 #() 
NAND3_X1_5346_ (
  .A1({ S1815 }),
  .A2({ S22836 }),
  .A3({ S1823 }),
  .ZN({ S1824 })
);
NAND2_X1 #() 
NAND2_X1_4959_ (
  .A1({ S1627 }),
  .A2({ S25921 }),
  .ZN({ S1825 })
);
OAI21_X1 #() 
OAI21_X1_2560_ (
  .A({ S25957[916] }),
  .B1({ S1825 }),
  .B2({ S86 }),
  .ZN({ S1826 })
);
AOI21_X1 #() 
AOI21_X1_2796_ (
  .A({ S1826 }),
  .B1({ S1780 }),
  .B2({ S1633 }),
  .ZN({ S1827 })
);
OAI211_X1 #() 
OAI211_X1_1722_ (
  .A({ S1624 }),
  .B({ S25957[915] }),
  .C1({ S25921 }),
  .C2({ S264 }),
  .ZN({ S1828 })
);
NOR2_X1 #() 
NOR2_X1_1258_ (
  .A1({ S1673 }),
  .A2({ S1675 }),
  .ZN({ S1829 })
);
AOI21_X1 #() 
AOI21_X1_2797_ (
  .A({ S25957[916] }),
  .B1({ S1829 }),
  .B2({ S1828 }),
  .ZN({ S1830 })
);
OAI21_X1 #() 
OAI21_X1_2561_ (
  .A({ S25957[917] }),
  .B1({ S1827 }),
  .B2({ S1830 }),
  .ZN({ S1831 })
);
AOI22_X1 #() 
AOI22_X1_560_ (
  .A1({ S1639 }),
  .A2({ S1624 }),
  .B1({ S25921 }),
  .B2({ S25957[913] }),
  .ZN({ S1832 })
);
INV_X1 #() 
INV_X1_1616_ (
  .A({ S1832 }),
  .ZN({ S1833 })
);
NAND2_X1 #() 
NAND2_X1_4960_ (
  .A1({ S1833 }),
  .A2({ S22985 }),
  .ZN({ S1834 })
);
NAND2_X1 #() 
NAND2_X1_4961_ (
  .A1({ S1623 }),
  .A2({ S1655 }),
  .ZN({ S1835 })
);
NAND2_X1 #() 
NAND2_X1_4962_ (
  .A1({ S1835 }),
  .A2({ S86 }),
  .ZN({ S1836 })
);
NAND3_X1 #() 
NAND3_X1_5347_ (
  .A1({ S1661 }),
  .A2({ S25957[915] }),
  .A3({ S1627 }),
  .ZN({ S1837 })
);
NAND3_X1 #() 
NAND3_X1_5348_ (
  .A1({ S1836 }),
  .A2({ S25957[916] }),
  .A3({ S1837 }),
  .ZN({ S1838 })
);
OAI211_X1 #() 
OAI211_X1_1723_ (
  .A({ S1838 }),
  .B({ S25608 }),
  .C1({ S1834 }),
  .C2({ S1736 }),
  .ZN({ S1839 })
);
NAND3_X1 #() 
NAND3_X1_5349_ (
  .A1({ S1831 }),
  .A2({ S25957[918] }),
  .A3({ S1839 }),
  .ZN({ S1840 })
);
NAND3_X1 #() 
NAND3_X1_5350_ (
  .A1({ S1824 }),
  .A2({ S25957[919] }),
  .A3({ S1840 }),
  .ZN({ S1841 })
);
INV_X1 #() 
INV_X1_1617_ (
  .A({ S1788 }),
  .ZN({ S1842 })
);
OAI21_X1 #() 
OAI21_X1_2562_ (
  .A({ S1642 }),
  .B1({ S1623 }),
  .B2({ S264 }),
  .ZN({ S1843 })
);
NAND2_X1 #() 
NAND2_X1_4963_ (
  .A1({ S1843 }),
  .A2({ S25957[915] }),
  .ZN({ S1844 })
);
NAND2_X1 #() 
NAND2_X1_4964_ (
  .A1({ S1623 }),
  .A2({ S86 }),
  .ZN({ S1845 })
);
OAI21_X1 #() 
OAI21_X1_2563_ (
  .A({ S1844 }),
  .B1({ S1842 }),
  .B2({ S1845 }),
  .ZN({ S1846 })
);
NAND4_X1 #() 
NAND4_X1_580_ (
  .A1({ S1790 }),
  .A2({ S1627 }),
  .A3({ S1642 }),
  .A4({ S86 }),
  .ZN({ S1847 })
);
NAND3_X1 #() 
NAND3_X1_5351_ (
  .A1({ S1649 }),
  .A2({ S25957[915] }),
  .A3({ S349 }),
  .ZN({ S1848 })
);
AND2_X1 #() 
AND2_X1_302_ (
  .A1({ S1848 }),
  .A2({ S25957[916] }),
  .ZN({ S1849 })
);
AOI22_X1 #() 
AOI22_X1_561_ (
  .A1({ S22985 }),
  .A2({ S1846 }),
  .B1({ S1849 }),
  .B2({ S1847 }),
  .ZN({ S1850 })
);
OR2_X1 #() 
OR2_X1_68_ (
  .A1({ S1850 }),
  .A2({ S22836 }),
  .ZN({ S1851 })
);
NAND3_X1 #() 
NAND3_X1_5352_ (
  .A1({ S1633 }),
  .A2({ S1642 }),
  .A3({ S1649 }),
  .ZN({ S1852 })
);
NOR2_X1 #() 
NOR2_X1_1259_ (
  .A1({ S1832 }),
  .A2({ S1757 }),
  .ZN({ S1853 })
);
NAND2_X1 #() 
NAND2_X1_4965_ (
  .A1({ S1853 }),
  .A2({ S25957[915] }),
  .ZN({ S1854 })
);
AND2_X1 #() 
AND2_X1_303_ (
  .A1({ S1854 }),
  .A2({ S1852 }),
  .ZN({ S1855 })
);
NAND2_X1 #() 
NAND2_X1_4966_ (
  .A1({ S1660 }),
  .A2({ S86 }),
  .ZN({ S1856 })
);
OAI21_X1 #() 
OAI21_X1_2564_ (
  .A({ S1629 }),
  .B1({ S25921 }),
  .B2({ S1856 }),
  .ZN({ S1857 })
);
OAI211_X1 #() 
OAI211_X1_1724_ (
  .A({ S22836 }),
  .B({ S1857 }),
  .C1({ S1855 }),
  .C2({ S22985 }),
  .ZN({ S1858 })
);
AOI21_X1 #() 
AOI21_X1_2798_ (
  .A({ S25957[917] }),
  .B1({ S1858 }),
  .B2({ S1851 }),
  .ZN({ S1859 })
);
NAND2_X1 #() 
NAND2_X1_4967_ (
  .A1({ S1693 }),
  .A2({ S86 }),
  .ZN({ S1860 })
);
OAI21_X1 #() 
OAI21_X1_2565_ (
  .A({ S25957[915] }),
  .B1({ S1642 }),
  .B2({ S264 }),
  .ZN({ S1861 })
);
OAI21_X1 #() 
OAI21_X1_2566_ (
  .A({ S1860 }),
  .B1({ S1832 }),
  .B2({ S1861 }),
  .ZN({ S1862 })
);
NAND2_X1 #() 
NAND2_X1_4968_ (
  .A1({ S1862 }),
  .A2({ S25957[916] }),
  .ZN({ S1863 })
);
OAI21_X1 #() 
OAI21_X1_2567_ (
  .A({ S1680 }),
  .B1({ S1632 }),
  .B2({ S1771 }),
  .ZN({ S1864 })
);
OAI211_X1 #() 
OAI211_X1_1725_ (
  .A({ S1863 }),
  .B({ S25957[918] }),
  .C1({ S25957[916] }),
  .C2({ S1864 }),
  .ZN({ S1865 })
);
AND3_X1 #() 
AND3_X1_205_ (
  .A1({ S1785 }),
  .A2({ S25957[916] }),
  .A3({ S1764 }),
  .ZN({ S1866 })
);
NAND4_X1 #() 
NAND4_X1_581_ (
  .A1({ S1639 }),
  .A2({ S1661 }),
  .A3({ S86 }),
  .A4({ S25957[913] }),
  .ZN({ S1867 })
);
AOI21_X1 #() 
AOI21_X1_2799_ (
  .A({ S25957[916] }),
  .B1({ S1867 }),
  .B2({ S1676 }),
  .ZN({ S1868 })
);
OAI21_X1 #() 
OAI21_X1_2568_ (
  .A({ S22836 }),
  .B1({ S1866 }),
  .B2({ S1868 }),
  .ZN({ S1869 })
);
AOI21_X1 #() 
AOI21_X1_2800_ (
  .A({ S25608 }),
  .B1({ S1865 }),
  .B2({ S1869 }),
  .ZN({ S1870 })
);
OAI21_X1 #() 
OAI21_X1_2569_ (
  .A({ S1685 }),
  .B1({ S1859 }),
  .B2({ S1870 }),
  .ZN({ S1871 })
);
NAND2_X1 #() 
NAND2_X1_4969_ (
  .A1({ S1871 }),
  .A2({ S1841 }),
  .ZN({ S1872 })
);
NAND2_X1 #() 
NAND2_X1_4970_ (
  .A1({ S1872 }),
  .A2({ S25957[1117] }),
  .ZN({ S1873 })
);
INV_X1 #() 
INV_X1_1618_ (
  .A({ S1873 }),
  .ZN({ S1874 })
);
NOR2_X1 #() 
NOR2_X1_1260_ (
  .A1({ S1872 }),
  .A2({ S25957[1117] }),
  .ZN({ S1875 })
);
OR3_X1 #() 
OR3_X1_31_ (
  .A1({ S1874 }),
  .A2({ S1875 }),
  .A3({ S22294 }),
  .ZN({ S1876 })
);
OAI21_X1 #() 
OAI21_X1_2570_ (
  .A({ S22294 }),
  .B1({ S1874 }),
  .B2({ S1875 }),
  .ZN({ S1877 })
);
NAND2_X1 #() 
NAND2_X1_4971_ (
  .A1({ S1876 }),
  .A2({ S1877 }),
  .ZN({ S25957[797] })
);
NAND2_X1 #() 
NAND2_X1_4972_ (
  .A1({ S25062 }),
  .A2({ S25059 }),
  .ZN({ S25957[956] })
);
NAND2_X1 #() 
NAND2_X1_4973_ (
  .A1({ S1688 }),
  .A2({ S86 }),
  .ZN({ S1878 })
);
AND2_X1 #() 
AND2_X1_304_ (
  .A1({ S1849 }),
  .A2({ S1878 }),
  .ZN({ S1879 })
);
NAND3_X1 #() 
NAND3_X1_5353_ (
  .A1({ S86 }),
  .A2({ S1686 }),
  .A3({ S25921 }),
  .ZN({ S1880 })
);
AND3_X1 #() 
AND3_X1_206_ (
  .A1({ S1712 }),
  .A2({ S22985 }),
  .A3({ S1880 }),
  .ZN({ S1881 })
);
OAI21_X1 #() 
OAI21_X1_2571_ (
  .A({ S25957[917] }),
  .B1({ S1879 }),
  .B2({ S1881 }),
  .ZN({ S1882 })
);
AOI22_X1 #() 
AOI22_X1_562_ (
  .A1({ S264 }),
  .A2({ S349 }),
  .B1({ S23078 }),
  .B2({ S23086 }),
  .ZN({ S1883 })
);
NAND2_X1 #() 
NAND2_X1_4974_ (
  .A1({ S1883 }),
  .A2({ S1639 }),
  .ZN({ S1884 })
);
AOI21_X1 #() 
AOI21_X1_2801_ (
  .A({ S25957[916] }),
  .B1({ S1884 }),
  .B2({ S1707 }),
  .ZN({ S1885 })
);
OAI21_X1 #() 
OAI21_X1_2572_ (
  .A({ S25957[916] }),
  .B1({ S1819 }),
  .B2({ S1772 }),
  .ZN({ S1886 })
);
NAND2_X1 #() 
NAND2_X1_4975_ (
  .A1({ S1886 }),
  .A2({ S25608 }),
  .ZN({ S1887 })
);
OAI211_X1 #() 
OAI211_X1_1726_ (
  .A({ S1882 }),
  .B({ S25957[918] }),
  .C1({ S1885 }),
  .C2({ S1887 }),
  .ZN({ S1888 })
);
NAND2_X1 #() 
NAND2_X1_4976_ (
  .A1({ S1628 }),
  .A2({ S1623 }),
  .ZN({ S1889 })
);
NAND2_X1 #() 
NAND2_X1_4977_ (
  .A1({ S1751 }),
  .A2({ S86 }),
  .ZN({ S1890 })
);
AND2_X1 #() 
AND2_X1_305_ (
  .A1({ S1890 }),
  .A2({ S1889 }),
  .ZN({ S1891 })
);
NAND2_X1 #() 
NAND2_X1_4978_ (
  .A1({ S1650 }),
  .A2({ S86 }),
  .ZN({ S1892 })
);
NOR2_X1 #() 
NOR2_X1_1261_ (
  .A1({ S1892 }),
  .A2({ S1687 }),
  .ZN({ S1893 })
);
NOR2_X1 #() 
NOR2_X1_1262_ (
  .A1({ S1635 }),
  .A2({ S1755 }),
  .ZN({ S1894 })
);
OAI21_X1 #() 
OAI21_X1_2573_ (
  .A({ S25957[916] }),
  .B1({ S1894 }),
  .B2({ S1893 }),
  .ZN({ S1895 })
);
OAI211_X1 #() 
OAI211_X1_1727_ (
  .A({ S1895 }),
  .B({ S25608 }),
  .C1({ S25957[916] }),
  .C2({ S1891 }),
  .ZN({ S1896 })
);
NAND3_X1 #() 
NAND3_X1_5354_ (
  .A1({ S1788 }),
  .A2({ S25957[915] }),
  .A3({ S1649 }),
  .ZN({ S1897 })
);
NAND2_X1 #() 
NAND2_X1_4979_ (
  .A1({ S1642 }),
  .A2({ S25957[913] }),
  .ZN({ S1898 })
);
NAND2_X1 #() 
NAND2_X1_4980_ (
  .A1({ S1623 }),
  .A2({ S264 }),
  .ZN({ S1899 })
);
NAND2_X1 #() 
NAND2_X1_4981_ (
  .A1({ S1899 }),
  .A2({ S1898 }),
  .ZN({ S1900 })
);
AOI21_X1 #() 
AOI21_X1_2802_ (
  .A({ S22985 }),
  .B1({ S1900 }),
  .B2({ S86 }),
  .ZN({ S1901 })
);
INV_X1 #() 
INV_X1_1619_ (
  .A({ S1658 }),
  .ZN({ S1902 })
);
OAI21_X1 #() 
OAI21_X1_2574_ (
  .A({ S86 }),
  .B1({ S1902 }),
  .B2({ S1656 }),
  .ZN({ S1903 })
);
NAND2_X1 #() 
NAND2_X1_4982_ (
  .A1({ S1818 }),
  .A2({ S25957[915] }),
  .ZN({ S1904 })
);
AND3_X1 #() 
AND3_X1_207_ (
  .A1({ S1904 }),
  .A2({ S1848 }),
  .A3({ S22985 }),
  .ZN({ S1905 })
);
AOI22_X1 #() 
AOI22_X1_563_ (
  .A1({ S1903 }),
  .A2({ S1905 }),
  .B1({ S1901 }),
  .B2({ S1897 }),
  .ZN({ S1906 })
);
OAI211_X1 #() 
OAI211_X1_1728_ (
  .A({ S1896 }),
  .B({ S22836 }),
  .C1({ S25608 }),
  .C2({ S1906 }),
  .ZN({ S1907 })
);
NAND2_X1 #() 
NAND2_X1_4983_ (
  .A1({ S1907 }),
  .A2({ S1888 }),
  .ZN({ S1908 })
);
NAND2_X1 #() 
NAND2_X1_4984_ (
  .A1({ S1908 }),
  .A2({ S25957[919] }),
  .ZN({ S1909 })
);
OAI21_X1 #() 
OAI21_X1_2575_ (
  .A({ S86 }),
  .B1({ S1807 }),
  .B2({ S1625 }),
  .ZN({ S1910 })
);
NAND2_X1 #() 
NAND2_X1_4985_ (
  .A1({ S1698 }),
  .A2({ S106 }),
  .ZN({ S1911 })
);
AND2_X1 #() 
AND2_X1_306_ (
  .A1({ S1910 }),
  .A2({ S1911 }),
  .ZN({ S1912 })
);
NOR2_X1 #() 
NOR2_X1_1263_ (
  .A1({ S1912 }),
  .A2({ S25957[917] }),
  .ZN({ S1913 })
);
NOR2_X1 #() 
NOR2_X1_1264_ (
  .A1({ S1622 }),
  .A2({ S25957[915] }),
  .ZN({ S1914 })
);
NOR2_X1 #() 
NOR2_X1_1265_ (
  .A1({ S1811 }),
  .A2({ S1914 }),
  .ZN({ S1915 })
);
OAI21_X1 #() 
OAI21_X1_2576_ (
  .A({ S22985 }),
  .B1({ S1915 }),
  .B2({ S25608 }),
  .ZN({ S1916 })
);
NAND3_X1 #() 
NAND3_X1_5355_ (
  .A1({ S1694 }),
  .A2({ S25957[917] }),
  .A3({ S1836 }),
  .ZN({ S1917 })
);
NAND3_X1 #() 
NAND3_X1_5356_ (
  .A1({ S1780 }),
  .A2({ S25957[915] }),
  .A3({ S1623 }),
  .ZN({ S1918 })
);
NAND3_X1 #() 
NAND3_X1_5357_ (
  .A1({ S1820 }),
  .A2({ S25608 }),
  .A3({ S1918 }),
  .ZN({ S1919 })
);
NAND3_X1 #() 
NAND3_X1_5358_ (
  .A1({ S1919 }),
  .A2({ S1917 }),
  .A3({ S25957[916] }),
  .ZN({ S1920 })
);
OAI21_X1 #() 
OAI21_X1_2577_ (
  .A({ S1920 }),
  .B1({ S1916 }),
  .B2({ S1913 }),
  .ZN({ S1921 })
);
NAND2_X1 #() 
NAND2_X1_4986_ (
  .A1({ S1921 }),
  .A2({ S22836 }),
  .ZN({ S1922 })
);
NOR2_X1 #() 
NOR2_X1_1266_ (
  .A1({ S1625 }),
  .A2({ S1737 }),
  .ZN({ S1923 })
);
NAND2_X1 #() 
NAND2_X1_4987_ (
  .A1({ S1722 }),
  .A2({ S22985 }),
  .ZN({ S1924 })
);
AOI21_X1 #() 
AOI21_X1_2803_ (
  .A({ S1924 }),
  .B1({ S1716 }),
  .B2({ S1639 }),
  .ZN({ S1925 })
);
NOR2_X1 #() 
NOR2_X1_1267_ (
  .A1({ S1925 }),
  .A2({ S25957[917] }),
  .ZN({ S1926 })
);
OAI21_X1 #() 
OAI21_X1_2578_ (
  .A({ S1926 }),
  .B1({ S1677 }),
  .B2({ S1923 }),
  .ZN({ S1927 })
);
AOI21_X1 #() 
AOI21_X1_2804_ (
  .A({ S1835 }),
  .B1({ S1666 }),
  .B2({ S106 }),
  .ZN({ S1928 })
);
NOR2_X1 #() 
NOR2_X1_1268_ (
  .A1({ S1928 }),
  .A2({ S25957[915] }),
  .ZN({ S1929 })
);
NAND2_X1 #() 
NAND2_X1_4988_ (
  .A1({ S1844 }),
  .A2({ S22985 }),
  .ZN({ S1930 })
);
AND2_X1 #() 
AND2_X1_307_ (
  .A1({ S349 }),
  .A2({ S131 }),
  .ZN({ S1931 })
);
OAI221_X1 #() 
OAI221_X1_146_ (
  .A({ S25957[917] }),
  .B1({ S22985 }),
  .B2({ S1931 }),
  .C1({ S1929 }),
  .C2({ S1930 }),
  .ZN({ S1932 })
);
NAND3_X1 #() 
NAND3_X1_5359_ (
  .A1({ S1927 }),
  .A2({ S1932 }),
  .A3({ S25957[918] }),
  .ZN({ S1933 })
);
NAND3_X1 #() 
NAND3_X1_5360_ (
  .A1({ S1922 }),
  .A2({ S1685 }),
  .A3({ S1933 }),
  .ZN({ S1934 })
);
NAND3_X1 #() 
NAND3_X1_5361_ (
  .A1({ S1909 }),
  .A2({ S25957[1116] }),
  .A3({ S1934 }),
  .ZN({ S1935 })
);
NAND3_X1 #() 
NAND3_X1_5362_ (
  .A1({ S1907 }),
  .A2({ S25957[919] }),
  .A3({ S1888 }),
  .ZN({ S1936 })
);
AND2_X1 #() 
AND2_X1_308_ (
  .A1({ S1927 }),
  .A2({ S1932 }),
  .ZN({ S1937 })
);
OAI211_X1 #() 
OAI211_X1_1729_ (
  .A({ S22836 }),
  .B({ S1920 }),
  .C1({ S1916 }),
  .C2({ S1913 }),
  .ZN({ S1938 })
);
OAI211_X1 #() 
OAI211_X1_1730_ (
  .A({ S1685 }),
  .B({ S1938 }),
  .C1({ S1937 }),
  .C2({ S22836 }),
  .ZN({ S1939 })
);
NAND3_X1 #() 
NAND3_X1_5363_ (
  .A1({ S1939 }),
  .A2({ S1936 }),
  .A3({ S24978 }),
  .ZN({ S1940 })
);
AOI21_X1 #() 
AOI21_X1_2805_ (
  .A({ S25957[956] }),
  .B1({ S1935 }),
  .B2({ S1940 }),
  .ZN({ S1941 })
);
INV_X1 #() 
INV_X1_1620_ (
  .A({ S25957[956] }),
  .ZN({ S1942 })
);
AOI21_X1 #() 
AOI21_X1_2806_ (
  .A({ S24978 }),
  .B1({ S1939 }),
  .B2({ S1936 }),
  .ZN({ S1943 })
);
INV_X1 #() 
INV_X1_1621_ (
  .A({ S1940 }),
  .ZN({ S1944 })
);
NOR3_X1 #() 
NOR3_X1_163_ (
  .A1({ S1944 }),
  .A2({ S1943 }),
  .A3({ S1942 }),
  .ZN({ S1945 })
);
OAI21_X1 #() 
OAI21_X1_2579_ (
  .A({ S25072 }),
  .B1({ S1945 }),
  .B2({ S1941 }),
  .ZN({ S1946 })
);
OAI21_X1 #() 
OAI21_X1_2580_ (
  .A({ S1942 }),
  .B1({ S1944 }),
  .B2({ S1943 }),
  .ZN({ S1947 })
);
NAND3_X1 #() 
NAND3_X1_5364_ (
  .A1({ S1935 }),
  .A2({ S25957[956] }),
  .A3({ S1940 }),
  .ZN({ S1948 })
);
NAND3_X1 #() 
NAND3_X1_5365_ (
  .A1({ S1947 }),
  .A2({ S25957[924] }),
  .A3({ S1948 }),
  .ZN({ S1949 })
);
AND2_X1 #() 
AND2_X1_309_ (
  .A1({ S1946 }),
  .A2({ S1949 }),
  .ZN({ S25957[796] })
);
INV_X1 #() 
INV_X1_1622_ (
  .A({ S1828 }),
  .ZN({ S1950 })
);
NOR2_X1 #() 
NOR2_X1_1269_ (
  .A1({ S1767 }),
  .A2({ S1818 }),
  .ZN({ S1951 })
);
AOI22_X1 #() 
AOI22_X1_564_ (
  .A1({ S1951 }),
  .A2({ S1649 }),
  .B1({ S1950 }),
  .B2({ S1899 }),
  .ZN({ S1952 })
);
INV_X1 #() 
INV_X1_1623_ (
  .A({ S1649 }),
  .ZN({ S1953 })
);
OAI211_X1 #() 
OAI211_X1_1731_ (
  .A({ S1911 }),
  .B({ S25957[916] }),
  .C1({ S1953 }),
  .C2({ S1892 }),
  .ZN({ S1954 })
);
OAI211_X1 #() 
OAI211_X1_1732_ (
  .A({ S1954 }),
  .B({ S25957[917] }),
  .C1({ S1952 }),
  .C2({ S25957[916] }),
  .ZN({ S1955 })
);
NAND2_X1 #() 
NAND2_X1_4989_ (
  .A1({ S1853 }),
  .A2({ S86 }),
  .ZN({ S1956 })
);
AOI21_X1 #() 
AOI21_X1_2807_ (
  .A({ S22985 }),
  .B1({ S1956 }),
  .B2({ S1828 }),
  .ZN({ S1957 })
);
OAI21_X1 #() 
OAI21_X1_2581_ (
  .A({ S25608 }),
  .B1({ S1743 }),
  .B2({ S1924 }),
  .ZN({ S1958 })
);
OAI211_X1 #() 
OAI211_X1_1733_ (
  .A({ S1955 }),
  .B({ S25957[918] }),
  .C1({ S1957 }),
  .C2({ S1958 }),
  .ZN({ S1959 })
);
NOR2_X1 #() 
NOR2_X1_1270_ (
  .A1({ S1832 }),
  .A2({ S1646 }),
  .ZN({ S1960 })
);
NAND2_X1 #() 
NAND2_X1_4990_ (
  .A1({ S1960 }),
  .A2({ S25957[915] }),
  .ZN({ S1961 })
);
OAI211_X1 #() 
OAI211_X1_1734_ (
  .A({ S1961 }),
  .B({ S22985 }),
  .C1({ S1647 }),
  .C2({ S25957[915] }),
  .ZN({ S1962 })
);
OAI211_X1 #() 
OAI211_X1_1735_ (
  .A({ S25957[916] }),
  .B({ S1884 }),
  .C1({ S1902 }),
  .C2({ S86 }),
  .ZN({ S1963 })
);
NAND3_X1 #() 
NAND3_X1_5366_ (
  .A1({ S1962 }),
  .A2({ S1963 }),
  .A3({ S25608 }),
  .ZN({ S1964 })
);
NAND3_X1 #() 
NAND3_X1_5367_ (
  .A1({ S1738 }),
  .A2({ S1639 }),
  .A3({ S1661 }),
  .ZN({ S1965 })
);
OAI211_X1 #() 
OAI211_X1_1736_ (
  .A({ S22985 }),
  .B({ S1965 }),
  .C1({ S1715 }),
  .C2({ S1737 }),
  .ZN({ S1966 })
);
AOI21_X1 #() 
AOI21_X1_2808_ (
  .A({ S25957[914] }),
  .B1({ S1649 }),
  .B2({ S1631 }),
  .ZN({ S1967 })
);
INV_X1 #() 
INV_X1_1624_ (
  .A({ S1720 }),
  .ZN({ S1968 })
);
OAI21_X1 #() 
OAI21_X1_2582_ (
  .A({ S86 }),
  .B1({ S1968 }),
  .B2({ S1771 }),
  .ZN({ S1969 })
);
OAI21_X1 #() 
OAI21_X1_2583_ (
  .A({ S1969 }),
  .B1({ S1967 }),
  .B2({ S1689 }),
  .ZN({ S1970 })
);
OAI211_X1 #() 
OAI211_X1_1737_ (
  .A({ S1966 }),
  .B({ S25957[917] }),
  .C1({ S1970 }),
  .C2({ S22985 }),
  .ZN({ S1971 })
);
NAND3_X1 #() 
NAND3_X1_5368_ (
  .A1({ S1964 }),
  .A2({ S1971 }),
  .A3({ S22836 }),
  .ZN({ S1972 })
);
NAND3_X1 #() 
NAND3_X1_5369_ (
  .A1({ S1972 }),
  .A2({ S1959 }),
  .A3({ S25957[919] }),
  .ZN({ S1973 })
);
AOI21_X1 #() 
AOI21_X1_2809_ (
  .A({ S1736 }),
  .B1({ S1716 }),
  .B2({ S1657 }),
  .ZN({ S1974 })
);
NAND2_X1 #() 
NAND2_X1_4991_ (
  .A1({ S86 }),
  .A2({ S1686 }),
  .ZN({ S1975 })
);
NOR2_X1 #() 
NOR2_X1_1271_ (
  .A1({ S1953 }),
  .A2({ S1975 }),
  .ZN({ S1976 })
);
NOR2_X1 #() 
NOR2_X1_1272_ (
  .A1({ S1680 }),
  .A2({ S1660 }),
  .ZN({ S1977 })
);
OAI21_X1 #() 
OAI21_X1_2584_ (
  .A({ S22985 }),
  .B1({ S1976 }),
  .B2({ S1977 }),
  .ZN({ S1978 })
);
OAI211_X1 #() 
OAI211_X1_1738_ (
  .A({ S25957[917] }),
  .B({ S1978 }),
  .C1({ S1974 }),
  .C2({ S22985 }),
  .ZN({ S1979 })
);
NAND2_X1 #() 
NAND2_X1_4992_ (
  .A1({ S1701 }),
  .A2({ S1918 }),
  .ZN({ S1980 })
);
OAI211_X1 #() 
OAI211_X1_1739_ (
  .A({ S1623 }),
  .B({ S86 }),
  .C1({ S25921 }),
  .C2({ S264 }),
  .ZN({ S1981 })
);
OAI211_X1 #() 
OAI211_X1_1740_ (
  .A({ S1980 }),
  .B({ S25608 }),
  .C1({ S22985 }),
  .C2({ S1981 }),
  .ZN({ S1982 })
);
NAND3_X1 #() 
NAND3_X1_5370_ (
  .A1({ S1979 }),
  .A2({ S25957[918] }),
  .A3({ S1982 }),
  .ZN({ S1983 })
);
INV_X1 #() 
INV_X1_1625_ (
  .A({ S106 }),
  .ZN({ S1984 })
);
OAI211_X1 #() 
OAI211_X1_1741_ (
  .A({ S25957[916] }),
  .B({ S25957[914] }),
  .C1({ S1914 }),
  .C2({ S1984 }),
  .ZN({ S1985 })
);
NAND3_X1 #() 
NAND3_X1_5371_ (
  .A1({ S1756 }),
  .A2({ S25957[912] }),
  .A3({ S1686 }),
  .ZN({ S1986 })
);
OAI21_X1 #() 
OAI21_X1_2585_ (
  .A({ S1985 }),
  .B1({ S25957[916] }),
  .B2({ S1986 }),
  .ZN({ S1987 })
);
NAND2_X1 #() 
NAND2_X1_4993_ (
  .A1({ S1987 }),
  .A2({ S25957[917] }),
  .ZN({ S1988 })
);
OAI21_X1 #() 
OAI21_X1_2586_ (
  .A({ S25957[915] }),
  .B1({ S1967 }),
  .B2({ S1625 }),
  .ZN({ S1989 })
);
AOI21_X1 #() 
AOI21_X1_2810_ (
  .A({ S22985 }),
  .B1({ S1989 }),
  .B2({ S1860 }),
  .ZN({ S1990 })
);
INV_X1 #() 
INV_X1_1626_ (
  .A({ S1639 }),
  .ZN({ S1991 })
);
NOR2_X1 #() 
NOR2_X1_1273_ (
  .A1({ S1687 }),
  .A2({ S1991 }),
  .ZN({ S1992 })
);
AOI22_X1 #() 
AOI22_X1_565_ (
  .A1({ S1992 }),
  .A2({ S25957[915] }),
  .B1({ S1657 }),
  .B2({ S1662 }),
  .ZN({ S1993 })
);
OAI21_X1 #() 
OAI21_X1_2587_ (
  .A({ S25608 }),
  .B1({ S1993 }),
  .B2({ S25957[916] }),
  .ZN({ S1994 })
);
OAI211_X1 #() 
OAI211_X1_1742_ (
  .A({ S1988 }),
  .B({ S22836 }),
  .C1({ S1994 }),
  .C2({ S1990 }),
  .ZN({ S1995 })
);
NAND3_X1 #() 
NAND3_X1_5372_ (
  .A1({ S1995 }),
  .A2({ S1983 }),
  .A3({ S1685 }),
  .ZN({ S1996 })
);
AOI21_X1 #() 
AOI21_X1_2811_ (
  .A({ S25166 }),
  .B1({ S1973 }),
  .B2({ S1996 }),
  .ZN({ S1997 })
);
AND3_X1 #() 
AND3_X1_208_ (
  .A1({ S1973 }),
  .A2({ S25166 }),
  .A3({ S1996 }),
  .ZN({ S1998 })
);
OAI21_X1 #() 
OAI21_X1_2588_ (
  .A({ S83 }),
  .B1({ S1998 }),
  .B2({ S1997 }),
  .ZN({ S1999 })
);
NAND2_X1 #() 
NAND2_X1_4994_ (
  .A1({ S1973 }),
  .A2({ S1996 }),
  .ZN({ S2000 })
);
NAND2_X1 #() 
NAND2_X1_4995_ (
  .A1({ S2000 }),
  .A2({ S25957[1115] }),
  .ZN({ S2001 })
);
NAND3_X1 #() 
NAND3_X1_5373_ (
  .A1({ S1973 }),
  .A2({ S25166 }),
  .A3({ S1996 }),
  .ZN({ S2002 })
);
NAND3_X1 #() 
NAND3_X1_5374_ (
  .A1({ S2001 }),
  .A2({ S25957[1051] }),
  .A3({ S2002 }),
  .ZN({ S2003 })
);
AND2_X1 #() 
AND2_X1_310_ (
  .A1({ S1999 }),
  .A2({ S2003 }),
  .ZN({ S107 })
);
INV_X1 #() 
INV_X1_1627_ (
  .A({ S107 }),
  .ZN({ S25957[795] })
);
OAI21_X1 #() 
OAI21_X1_2589_ (
  .A({ S25957[915] }),
  .B1({ S1675 }),
  .B2({ S25957[913] }),
  .ZN({ S2004 })
);
NOR2_X1 #() 
NOR2_X1_1274_ (
  .A1({ S2004 }),
  .A2({ S1843 }),
  .ZN({ S2005 })
);
INV_X1 #() 
INV_X1_1628_ (
  .A({ S2005 }),
  .ZN({ S2006 })
);
NOR2_X1 #() 
NOR2_X1_1275_ (
  .A1({ S1951 }),
  .A2({ S22985 }),
  .ZN({ S2007 })
);
AOI22_X1 #() 
AOI22_X1_566_ (
  .A1({ S2006 }),
  .A2({ S2007 }),
  .B1({ S1752 }),
  .B2({ S1679 }),
  .ZN({ S2008 })
);
NAND2_X1 #() 
NAND2_X1_4996_ (
  .A1({ S1899 }),
  .A2({ S86 }),
  .ZN({ S2009 })
);
NAND3_X1 #() 
NAND3_X1_5375_ (
  .A1({ S1844 }),
  .A2({ S22985 }),
  .A3({ S2009 }),
  .ZN({ S2010 })
);
NAND4_X1 #() 
NAND4_X1_582_ (
  .A1({ S25957[916] }),
  .A2({ S1788 }),
  .A3({ S1680 }),
  .A4({ S1655 }),
  .ZN({ S2011 })
);
NAND3_X1 #() 
NAND3_X1_5376_ (
  .A1({ S2010 }),
  .A2({ S25608 }),
  .A3({ S2011 }),
  .ZN({ S2012 })
);
OAI211_X1 #() 
OAI211_X1_1743_ (
  .A({ S2012 }),
  .B({ S25957[918] }),
  .C1({ S2008 }),
  .C2({ S25608 }),
  .ZN({ S2013 })
);
OAI21_X1 #() 
OAI21_X1_2590_ (
  .A({ S25957[916] }),
  .B1({ S1902 }),
  .B2({ S86 }),
  .ZN({ S2014 })
);
NAND3_X1 #() 
NAND3_X1_5377_ (
  .A1({ S1790 }),
  .A2({ S106 }),
  .A3({ S25957[915] }),
  .ZN({ S2015 })
);
OAI21_X1 #() 
OAI21_X1_2591_ (
  .A({ S2015 }),
  .B1({ S1878 }),
  .B2({ S1757 }),
  .ZN({ S2016 })
);
NAND2_X1 #() 
NAND2_X1_4997_ (
  .A1({ S2016 }),
  .A2({ S22985 }),
  .ZN({ S2017 })
);
AOI21_X1 #() 
AOI21_X1_2812_ (
  .A({ S25957[915] }),
  .B1({ S1899 }),
  .B2({ S1790 }),
  .ZN({ S2018 })
);
OAI21_X1 #() 
OAI21_X1_2592_ (
  .A({ S2017 }),
  .B1({ S2014 }),
  .B2({ S2018 }),
  .ZN({ S2019 })
);
OAI21_X1 #() 
OAI21_X1_2593_ (
  .A({ S1911 }),
  .B1({ S1632 }),
  .B2({ S1771 }),
  .ZN({ S2020 })
);
NAND3_X1 #() 
NAND3_X1_5378_ (
  .A1({ S1852 }),
  .A2({ S1773 }),
  .A3({ S22985 }),
  .ZN({ S2021 })
);
OAI211_X1 #() 
OAI211_X1_1744_ (
  .A({ S2021 }),
  .B({ S25957[917] }),
  .C1({ S22985 }),
  .C2({ S2020 }),
  .ZN({ S2022 })
);
OAI211_X1 #() 
OAI211_X1_1745_ (
  .A({ S2022 }),
  .B({ S22836 }),
  .C1({ S25957[917] }),
  .C2({ S2019 }),
  .ZN({ S2023 })
);
NAND3_X1 #() 
NAND3_X1_5379_ (
  .A1({ S2023 }),
  .A2({ S1685 }),
  .A3({ S2013 }),
  .ZN({ S2024 })
);
NAND3_X1 #() 
NAND3_X1_5380_ (
  .A1({ S1747 }),
  .A2({ S1640 }),
  .A3({ S86 }),
  .ZN({ S2025 })
);
AND2_X1 #() 
AND2_X1_311_ (
  .A1({ S1641 }),
  .A2({ S22985 }),
  .ZN({ S2026 })
);
OAI21_X1 #() 
OAI21_X1_2594_ (
  .A({ S1910 }),
  .B1({ S1818 }),
  .B2({ S1722 }),
  .ZN({ S2027 })
);
AOI22_X1 #() 
AOI22_X1_567_ (
  .A1({ S2027 }),
  .A2({ S25957[916] }),
  .B1({ S2026 }),
  .B2({ S2025 }),
  .ZN({ S2028 })
);
OAI21_X1 #() 
OAI21_X1_2595_ (
  .A({ S1844 }),
  .B1({ S25957[915] }),
  .B2({ S1842 }),
  .ZN({ S2029 })
);
NAND4_X1 #() 
NAND4_X1_583_ (
  .A1({ S1649 }),
  .A2({ S1631 }),
  .A3({ S25957[915] }),
  .A4({ S25957[914] }),
  .ZN({ S2030 })
);
NAND2_X1 #() 
NAND2_X1_4998_ (
  .A1({ S1901 }),
  .A2({ S2030 }),
  .ZN({ S2031 })
);
OAI211_X1 #() 
OAI211_X1_1746_ (
  .A({ S2031 }),
  .B({ S25608 }),
  .C1({ S25957[916] }),
  .C2({ S2029 }),
  .ZN({ S2032 })
);
OAI211_X1 #() 
OAI211_X1_1747_ (
  .A({ S2032 }),
  .B({ S25957[918] }),
  .C1({ S2028 }),
  .C2({ S25608 }),
  .ZN({ S2033 })
);
INV_X1 #() 
INV_X1_1629_ (
  .A({ S1634 }),
  .ZN({ S2034 })
);
OAI211_X1 #() 
OAI211_X1_1748_ (
  .A({ S1689 }),
  .B({ S25957[916] }),
  .C1({ S2034 }),
  .C2({ S1643 }),
  .ZN({ S2035 })
);
NAND4_X1 #() 
NAND4_X1_584_ (
  .A1({ S1904 }),
  .A2({ S1878 }),
  .A3({ S1848 }),
  .A4({ S22985 }),
  .ZN({ S2036 })
);
NAND3_X1 #() 
NAND3_X1_5381_ (
  .A1({ S2035 }),
  .A2({ S2036 }),
  .A3({ S25957[917] }),
  .ZN({ S2037 })
);
AOI21_X1 #() 
AOI21_X1_2813_ (
  .A({ S1977 }),
  .B1({ S1778 }),
  .B2({ S86 }),
  .ZN({ S2038 })
);
OAI211_X1 #() 
OAI211_X1_1749_ (
  .A({ S25957[916] }),
  .B({ S1783 }),
  .C1({ S1810 }),
  .C2({ S25957[915] }),
  .ZN({ S2039 })
);
OAI21_X1 #() 
OAI21_X1_2596_ (
  .A({ S2039 }),
  .B1({ S2038 }),
  .B2({ S25957[916] }),
  .ZN({ S2040 })
);
NAND2_X1 #() 
NAND2_X1_4999_ (
  .A1({ S2040 }),
  .A2({ S25608 }),
  .ZN({ S2041 })
);
NAND3_X1 #() 
NAND3_X1_5382_ (
  .A1({ S2041 }),
  .A2({ S22836 }),
  .A3({ S2037 }),
  .ZN({ S2042 })
);
NAND3_X1 #() 
NAND3_X1_5383_ (
  .A1({ S2033 }),
  .A2({ S2042 }),
  .A3({ S25957[919] }),
  .ZN({ S2043 })
);
NAND3_X1 #() 
NAND3_X1_5384_ (
  .A1({ S2043 }),
  .A2({ S2024 }),
  .A3({ S25180 }),
  .ZN({ S2044 })
);
NAND2_X1 #() 
NAND2_X1_5000_ (
  .A1({ S2028 }),
  .A2({ S25957[917] }),
  .ZN({ S2045 })
);
OAI21_X1 #() 
OAI21_X1_2597_ (
  .A({ S2031 }),
  .B1({ S25957[916] }),
  .B2({ S2029 }),
  .ZN({ S2046 })
);
NAND2_X1 #() 
NAND2_X1_5001_ (
  .A1({ S2046 }),
  .A2({ S25608 }),
  .ZN({ S2047 })
);
NAND3_X1 #() 
NAND3_X1_5385_ (
  .A1({ S2047 }),
  .A2({ S2045 }),
  .A3({ S25957[918] }),
  .ZN({ S2048 })
);
NAND2_X1 #() 
NAND2_X1_5002_ (
  .A1({ S2035 }),
  .A2({ S2036 }),
  .ZN({ S2049 })
);
NAND2_X1 #() 
NAND2_X1_5003_ (
  .A1({ S2049 }),
  .A2({ S25957[917] }),
  .ZN({ S2050 })
);
OAI211_X1 #() 
OAI211_X1_1750_ (
  .A({ S2050 }),
  .B({ S22836 }),
  .C1({ S25957[917] }),
  .C2({ S2040 }),
  .ZN({ S2051 })
);
NAND3_X1 #() 
NAND3_X1_5386_ (
  .A1({ S2048 }),
  .A2({ S25957[919] }),
  .A3({ S2051 }),
  .ZN({ S2052 })
);
AND2_X1 #() 
AND2_X1_312_ (
  .A1({ S2010 }),
  .A2({ S2011 }),
  .ZN({ S2053 })
);
NAND2_X1 #() 
NAND2_X1_5004_ (
  .A1({ S2006 }),
  .A2({ S2007 }),
  .ZN({ S2054 })
);
AOI21_X1 #() 
AOI21_X1_2814_ (
  .A({ S25608 }),
  .B1({ S1752 }),
  .B2({ S1679 }),
  .ZN({ S2055 })
);
NAND2_X1 #() 
NAND2_X1_5005_ (
  .A1({ S2054 }),
  .A2({ S2055 }),
  .ZN({ S2056 })
);
OAI211_X1 #() 
OAI211_X1_1751_ (
  .A({ S2056 }),
  .B({ S25957[918] }),
  .C1({ S25957[917] }),
  .C2({ S2053 }),
  .ZN({ S2057 })
);
NAND2_X1 #() 
NAND2_X1_5006_ (
  .A1({ S1852 }),
  .A2({ S1773 }),
  .ZN({ S2058 })
);
INV_X1 #() 
INV_X1_1630_ (
  .A({ S2058 }),
  .ZN({ S2059 })
);
AOI21_X1 #() 
AOI21_X1_2815_ (
  .A({ S25608 }),
  .B1({ S2020 }),
  .B2({ S25957[916] }),
  .ZN({ S2060 })
);
OAI21_X1 #() 
OAI21_X1_2598_ (
  .A({ S2060 }),
  .B1({ S2059 }),
  .B2({ S25957[916] }),
  .ZN({ S2061 })
);
NAND2_X1 #() 
NAND2_X1_5007_ (
  .A1({ S2019 }),
  .A2({ S25608 }),
  .ZN({ S2062 })
);
NAND3_X1 #() 
NAND3_X1_5387_ (
  .A1({ S2062 }),
  .A2({ S2061 }),
  .A3({ S22836 }),
  .ZN({ S2063 })
);
NAND3_X1 #() 
NAND3_X1_5388_ (
  .A1({ S2063 }),
  .A2({ S1685 }),
  .A3({ S2057 }),
  .ZN({ S2064 })
);
NAND3_X1 #() 
NAND3_X1_5389_ (
  .A1({ S2052 }),
  .A2({ S2064 }),
  .A3({ S25957[1112] }),
  .ZN({ S2065 })
);
AOI21_X1 #() 
AOI21_X1_2816_ (
  .A({ S25957[1048] }),
  .B1({ S2065 }),
  .B2({ S2044 }),
  .ZN({ S2066 })
);
AND3_X1 #() 
AND3_X1_209_ (
  .A1({ S2065 }),
  .A2({ S2044 }),
  .A3({ S25957[1048] }),
  .ZN({ S2067 })
);
OR2_X1 #() 
OR2_X1_69_ (
  .A1({ S2067 }),
  .A2({ S2066 }),
  .ZN({ S25957[792] })
);
NOR2_X1 #() 
NOR2_X1_1276_ (
  .A1({ S22563 }),
  .A2({ S22566 }),
  .ZN({ S25957[1081] })
);
NOR2_X1 #() 
NOR2_X1_1277_ (
  .A1({ S25329 }),
  .A2({ S25311 }),
  .ZN({ S2068 })
);
XNOR2_X1 #() 
XNOR2_X1_194_ (
  .A({ S2068 }),
  .B({ S25957[1081] }),
  .ZN({ S25957[953] })
);
INV_X1 #() 
INV_X1_1631_ (
  .A({ S25957[953] }),
  .ZN({ S2069 })
);
INV_X1 #() 
INV_X1_1632_ (
  .A({ S2068 }),
  .ZN({ S25957[985] })
);
NAND2_X1 #() 
NAND2_X1_5008_ (
  .A1({ S22565 }),
  .A2({ S22564 }),
  .ZN({ S25957[1145] })
);
NAND2_X1 #() 
NAND2_X1_5009_ (
  .A1({ S25318 }),
  .A2({ S25328 }),
  .ZN({ S2070 })
);
XOR2_X1 #() 
XOR2_X1_80_ (
  .A({ S2070 }),
  .B({ S25957[1145] }),
  .Z({ S2071 })
);
NAND2_X1 #() 
NAND2_X1_5010_ (
  .A1({ S1890 }),
  .A2({ S22985 }),
  .ZN({ S2072 })
);
NAND3_X1 #() 
NAND3_X1_5390_ (
  .A1({ S1788 }),
  .A2({ S86 }),
  .A3({ S1655 }),
  .ZN({ S2073 })
);
AOI21_X1 #() 
AOI21_X1_2817_ (
  .A({ S25957[917] }),
  .B1({ S2073 }),
  .B2({ S1739 }),
  .ZN({ S2074 })
);
OAI21_X1 #() 
OAI21_X1_2599_ (
  .A({ S2074 }),
  .B1({ S2072 }),
  .B2({ S1703 }),
  .ZN({ S2075 })
);
NAND2_X1 #() 
NAND2_X1_5011_ (
  .A1({ S1661 }),
  .A2({ S25957[915] }),
  .ZN({ S2076 })
);
NOR2_X1 #() 
NOR2_X1_1278_ (
  .A1({ S1715 }),
  .A2({ S2076 }),
  .ZN({ S2077 })
);
OAI211_X1 #() 
OAI211_X1_1752_ (
  .A({ S1837 }),
  .B({ S22985 }),
  .C1({ S1953 }),
  .C2({ S1975 }),
  .ZN({ S2078 })
);
OAI211_X1 #() 
OAI211_X1_1753_ (
  .A({ S25957[917] }),
  .B({ S2078 }),
  .C1({ S2077 }),
  .C2({ S1692 }),
  .ZN({ S2079 })
);
NAND3_X1 #() 
NAND3_X1_5391_ (
  .A1({ S2075 }),
  .A2({ S22836 }),
  .A3({ S2079 }),
  .ZN({ S2080 })
);
NAND3_X1 #() 
NAND3_X1_5392_ (
  .A1({ S1708 }),
  .A2({ S1711 }),
  .A3({ S22985 }),
  .ZN({ S2081 })
);
NAND3_X1 #() 
NAND3_X1_5393_ (
  .A1({ S1828 }),
  .A2({ S1695 }),
  .A3({ S25957[916] }),
  .ZN({ S2082 })
);
OAI211_X1 #() 
OAI211_X1_1754_ (
  .A({ S25957[917] }),
  .B({ S2082 }),
  .C1({ S2005 }),
  .C2({ S2081 }),
  .ZN({ S2083 })
);
OAI211_X1 #() 
OAI211_X1_1755_ (
  .A({ S1639 }),
  .B({ S25957[915] }),
  .C1({ S25921 }),
  .C2({ S264 }),
  .ZN({ S2084 })
);
OAI211_X1 #() 
OAI211_X1_1756_ (
  .A({ S22985 }),
  .B({ S2084 }),
  .C1({ S1981 }),
  .C2({ S1807 }),
  .ZN({ S2085 })
);
NAND3_X1 #() 
NAND3_X1_5394_ (
  .A1({ S1624 }),
  .A2({ S86 }),
  .A3({ S25921 }),
  .ZN({ S2086 })
);
OAI211_X1 #() 
OAI211_X1_1757_ (
  .A({ S25957[916] }),
  .B({ S2086 }),
  .C1({ S1832 }),
  .C2({ S1861 }),
  .ZN({ S2087 })
);
NAND3_X1 #() 
NAND3_X1_5395_ (
  .A1({ S2087 }),
  .A2({ S2085 }),
  .A3({ S25608 }),
  .ZN({ S2088 })
);
NAND3_X1 #() 
NAND3_X1_5396_ (
  .A1({ S2088 }),
  .A2({ S2083 }),
  .A3({ S25957[918] }),
  .ZN({ S2089 })
);
NAND3_X1 #() 
NAND3_X1_5397_ (
  .A1({ S2080 }),
  .A2({ S25957[919] }),
  .A3({ S2089 }),
  .ZN({ S2090 })
);
NAND2_X1 #() 
NAND2_X1_5012_ (
  .A1({ S1623 }),
  .A2({ S25957[915] }),
  .ZN({ S2091 })
);
NAND2_X1 #() 
NAND2_X1_5013_ (
  .A1({ S1747 }),
  .A2({ S1640 }),
  .ZN({ S2092 })
);
NAND2_X1 #() 
NAND2_X1_5014_ (
  .A1({ S1662 }),
  .A2({ S1688 }),
  .ZN({ S2093 })
);
OAI211_X1 #() 
OAI211_X1_1758_ (
  .A({ S2093 }),
  .B({ S25957[916] }),
  .C1({ S2091 }),
  .C2({ S2092 }),
  .ZN({ S2094 })
);
NAND2_X1 #() 
NAND2_X1_5015_ (
  .A1({ S1825 }),
  .A2({ S1661 }),
  .ZN({ S2095 })
);
AOI21_X1 #() 
AOI21_X1_2818_ (
  .A({ S22836 }),
  .B1({ S1821 }),
  .B2({ S2095 }),
  .ZN({ S2096 })
);
NAND2_X1 #() 
NAND2_X1_5016_ (
  .A1({ S2094 }),
  .A2({ S2096 }),
  .ZN({ S2097 })
);
AOI21_X1 #() 
AOI21_X1_2819_ (
  .A({ S22985 }),
  .B1({ S1965 }),
  .B2({ S1880 }),
  .ZN({ S2098 })
);
OAI21_X1 #() 
OAI21_X1_2600_ (
  .A({ S22836 }),
  .B1({ S2098 }),
  .B2({ S1701 }),
  .ZN({ S2099 })
);
AOI21_X1 #() 
AOI21_X1_2820_ (
  .A({ S25608 }),
  .B1({ S2097 }),
  .B2({ S2099 }),
  .ZN({ S2100 })
);
AOI21_X1 #() 
AOI21_X1_2821_ (
  .A({ S25957[916] }),
  .B1({ S2030 }),
  .B2({ S1744 }),
  .ZN({ S2101 })
);
OAI21_X1 #() 
OAI21_X1_2601_ (
  .A({ S1784 }),
  .B1({ S25957[915] }),
  .B2({ S264 }),
  .ZN({ S2102 })
);
AOI21_X1 #() 
AOI21_X1_2822_ (
  .A({ S22985 }),
  .B1({ S25957[913] }),
  .B2({ S1675 }),
  .ZN({ S2103 })
);
AND3_X1 #() 
AND3_X1_210_ (
  .A1({ S2102 }),
  .A2({ S2103 }),
  .A3({ S1889 }),
  .ZN({ S2104 })
);
OAI21_X1 #() 
OAI21_X1_2602_ (
  .A({ S25957[918] }),
  .B1({ S2104 }),
  .B2({ S2101 }),
  .ZN({ S2105 })
);
NOR2_X1 #() 
NOR2_X1_1279_ (
  .A1({ S1737 }),
  .A2({ S1991 }),
  .ZN({ S2106 })
);
OAI21_X1 #() 
OAI21_X1_2603_ (
  .A({ S1670 }),
  .B1({ S25957[915] }),
  .B2({ S1700 }),
  .ZN({ S2107 })
);
OAI211_X1 #() 
OAI211_X1_1759_ (
  .A({ S2107 }),
  .B({ S22836 }),
  .C1({ S1677 }),
  .C2({ S2106 }),
  .ZN({ S2108 })
);
AOI21_X1 #() 
AOI21_X1_2823_ (
  .A({ S25957[917] }),
  .B1({ S2105 }),
  .B2({ S2108 }),
  .ZN({ S2109 })
);
OAI21_X1 #() 
OAI21_X1_2604_ (
  .A({ S1685 }),
  .B1({ S2109 }),
  .B2({ S2100 }),
  .ZN({ S2110 })
);
NAND3_X1 #() 
NAND3_X1_5398_ (
  .A1({ S2110 }),
  .A2({ S2071 }),
  .A3({ S2090 }),
  .ZN({ S2111 })
);
INV_X1 #() 
INV_X1_1633_ (
  .A({ S2071 }),
  .ZN({ S25957[1017] })
);
AND3_X1 #() 
AND3_X1_211_ (
  .A1({ S2080 }),
  .A2({ S25957[919] }),
  .A3({ S2089 }),
  .ZN({ S2112 })
);
INV_X1 #() 
INV_X1_1634_ (
  .A({ S2101 }),
  .ZN({ S2113 })
);
NAND3_X1 #() 
NAND3_X1_5399_ (
  .A1({ S2102 }),
  .A2({ S2103 }),
  .A3({ S1889 }),
  .ZN({ S2114 })
);
NAND3_X1 #() 
NAND3_X1_5400_ (
  .A1({ S2113 }),
  .A2({ S2114 }),
  .A3({ S25608 }),
  .ZN({ S2115 })
);
OAI21_X1 #() 
OAI21_X1_2605_ (
  .A({ S106 }),
  .B1({ S1622 }),
  .B2({ S25957[914] }),
  .ZN({ S2116 })
);
AOI22_X1 #() 
AOI22_X1_568_ (
  .A1({ S2116 }),
  .A2({ S25957[915] }),
  .B1({ S1662 }),
  .B2({ S1688 }),
  .ZN({ S2117 })
);
NAND2_X1 #() 
NAND2_X1_5017_ (
  .A1({ S2095 }),
  .A2({ S1674 }),
  .ZN({ S2118 })
);
NAND2_X1 #() 
NAND2_X1_5018_ (
  .A1({ S2118 }),
  .A2({ S22985 }),
  .ZN({ S2119 })
);
OAI211_X1 #() 
OAI211_X1_1760_ (
  .A({ S2119 }),
  .B({ S25957[917] }),
  .C1({ S2117 }),
  .C2({ S22985 }),
  .ZN({ S2120 })
);
NAND3_X1 #() 
NAND3_X1_5401_ (
  .A1({ S2120 }),
  .A2({ S2115 }),
  .A3({ S25957[918] }),
  .ZN({ S2121 })
);
NAND2_X1 #() 
NAND2_X1_5019_ (
  .A1({ S1700 }),
  .A2({ S86 }),
  .ZN({ S2122 })
);
NAND2_X1 #() 
NAND2_X1_5020_ (
  .A1({ S2122 }),
  .A2({ S22985 }),
  .ZN({ S2123 })
);
INV_X1 #() 
INV_X1_1635_ (
  .A({ S2098 }),
  .ZN({ S2124 })
);
AOI21_X1 #() 
AOI21_X1_2824_ (
  .A({ S25608 }),
  .B1({ S2124 }),
  .B2({ S2123 }),
  .ZN({ S2125 })
);
AOI21_X1 #() 
AOI21_X1_2825_ (
  .A({ S1669 }),
  .B1({ S1693 }),
  .B2({ S1768 }),
  .ZN({ S2126 })
);
OAI21_X1 #() 
OAI21_X1_2606_ (
  .A({ S25608 }),
  .B1({ S1677 }),
  .B2({ S2106 }),
  .ZN({ S2127 })
);
NOR2_X1 #() 
NOR2_X1_1280_ (
  .A1({ S2127 }),
  .A2({ S2126 }),
  .ZN({ S2128 })
);
OAI21_X1 #() 
OAI21_X1_2607_ (
  .A({ S22836 }),
  .B1({ S2125 }),
  .B2({ S2128 }),
  .ZN({ S2129 })
);
AOI21_X1 #() 
AOI21_X1_2826_ (
  .A({ S25957[919] }),
  .B1({ S2129 }),
  .B2({ S2121 }),
  .ZN({ S2130 })
);
OAI21_X1 #() 
OAI21_X1_2608_ (
  .A({ S25957[1017] }),
  .B1({ S2130 }),
  .B2({ S2112 }),
  .ZN({ S2131 })
);
NAND3_X1 #() 
NAND3_X1_5402_ (
  .A1({ S2131 }),
  .A2({ S25957[985] }),
  .A3({ S2111 }),
  .ZN({ S2132 })
);
OAI21_X1 #() 
OAI21_X1_2609_ (
  .A({ S2071 }),
  .B1({ S2130 }),
  .B2({ S2112 }),
  .ZN({ S2133 })
);
NAND3_X1 #() 
NAND3_X1_5403_ (
  .A1({ S2110 }),
  .A2({ S25957[1017] }),
  .A3({ S2090 }),
  .ZN({ S2134 })
);
NAND3_X1 #() 
NAND3_X1_5404_ (
  .A1({ S2133 }),
  .A2({ S2068 }),
  .A3({ S2134 }),
  .ZN({ S2135 })
);
AOI21_X1 #() 
AOI21_X1_2827_ (
  .A({ S2069 }),
  .B1({ S2132 }),
  .B2({ S2135 }),
  .ZN({ S2136 })
);
NAND3_X1 #() 
NAND3_X1_5405_ (
  .A1({ S2133 }),
  .A2({ S25957[985] }),
  .A3({ S2134 }),
  .ZN({ S2137 })
);
NAND3_X1 #() 
NAND3_X1_5406_ (
  .A1({ S2131 }),
  .A2({ S2068 }),
  .A3({ S2111 }),
  .ZN({ S2138 })
);
AOI21_X1 #() 
AOI21_X1_2828_ (
  .A({ S25957[953] }),
  .B1({ S2137 }),
  .B2({ S2138 }),
  .ZN({ S2139 })
);
OAI21_X1 #() 
OAI21_X1_2610_ (
  .A({ S25957[921] }),
  .B1({ S2136 }),
  .B2({ S2139 }),
  .ZN({ S2140 })
);
NAND3_X1 #() 
NAND3_X1_5407_ (
  .A1({ S2137 }),
  .A2({ S2138 }),
  .A3({ S25957[953] }),
  .ZN({ S2141 })
);
NAND3_X1 #() 
NAND3_X1_5408_ (
  .A1({ S2132 }),
  .A2({ S2135 }),
  .A3({ S2069 }),
  .ZN({ S2142 })
);
NAND3_X1 #() 
NAND3_X1_5409_ (
  .A1({ S2141 }),
  .A2({ S2142 }),
  .A3({ S1019 }),
  .ZN({ S2143 })
);
NAND2_X1 #() 
NAND2_X1_5021_ (
  .A1({ S2140 }),
  .A2({ S2143 }),
  .ZN({ S25957[793] })
);
NAND2_X1 #() 
NAND2_X1_5022_ (
  .A1({ S25400 }),
  .A2({ S25399 }),
  .ZN({ S25957[1018] })
);
XNOR2_X1 #() 
XNOR2_X1_195_ (
  .A({ S25957[1018] }),
  .B({ S22622 }),
  .ZN({ S25957[954] })
);
INV_X1 #() 
INV_X1_1636_ (
  .A({ S25957[954] }),
  .ZN({ S2144 })
);
NAND2_X1 #() 
NAND2_X1_5023_ (
  .A1({ S25397 }),
  .A2({ S25401 }),
  .ZN({ S2145 })
);
INV_X1 #() 
INV_X1_1637_ (
  .A({ S2145 }),
  .ZN({ S25957[986] })
);
NOR2_X1 #() 
NOR2_X1_1281_ (
  .A1({ S1646 }),
  .A2({ S25921 }),
  .ZN({ S2146 })
);
NAND2_X1 #() 
NAND2_X1_5024_ (
  .A1({ S2146 }),
  .A2({ S25957[915] }),
  .ZN({ S2147 })
);
OAI211_X1 #() 
OAI211_X1_1761_ (
  .A({ S2147 }),
  .B({ S25957[916] }),
  .C1({ S25957[915] }),
  .C2({ S1700 }),
  .ZN({ S2148 })
);
INV_X1 #() 
INV_X1_1638_ (
  .A({ S2148 }),
  .ZN({ S2149 })
);
NAND2_X1 #() 
NAND2_X1_5025_ (
  .A1({ S25957[915] }),
  .A2({ S25957[913] }),
  .ZN({ S2150 })
);
AOI22_X1 #() 
AOI22_X1_569_ (
  .A1({ S2150 }),
  .A2({ S25957[914] }),
  .B1({ S25921 }),
  .B2({ S25957[915] }),
  .ZN({ S2151 })
);
NAND2_X1 #() 
NAND2_X1_5026_ (
  .A1({ S106 }),
  .A2({ S22985 }),
  .ZN({ S2152 })
);
OAI21_X1 #() 
OAI21_X1_2611_ (
  .A({ S25957[917] }),
  .B1({ S2151 }),
  .B2({ S2152 }),
  .ZN({ S2153 })
);
NAND2_X1 #() 
NAND2_X1_5027_ (
  .A1({ S1738 }),
  .A2({ S1661 }),
  .ZN({ S2154 })
);
NAND3_X1 #() 
NAND3_X1_5410_ (
  .A1({ S2154 }),
  .A2({ S25957[916] }),
  .A3({ S1975 }),
  .ZN({ S2155 })
);
NAND3_X1 #() 
NAND3_X1_5411_ (
  .A1({ S1785 }),
  .A2({ S22985 }),
  .A3({ S1783 }),
  .ZN({ S2156 })
);
NAND3_X1 #() 
NAND3_X1_5412_ (
  .A1({ S2156 }),
  .A2({ S25608 }),
  .A3({ S2155 }),
  .ZN({ S2157 })
);
OAI211_X1 #() 
OAI211_X1_1762_ (
  .A({ S2157 }),
  .B({ S22836 }),
  .C1({ S2149 }),
  .C2({ S2153 }),
  .ZN({ S2158 })
);
AOI21_X1 #() 
AOI21_X1_2829_ (
  .A({ S25957[915] }),
  .B1({ S1747 }),
  .B2({ S1640 }),
  .ZN({ S2159 })
);
OAI21_X1 #() 
OAI21_X1_2612_ (
  .A({ S25957[916] }),
  .B1({ S2091 }),
  .B2({ S1755 }),
  .ZN({ S2160 })
);
NOR3_X1 #() 
NOR3_X1_164_ (
  .A1({ S1967 }),
  .A2({ S1835 }),
  .A3({ S86 }),
  .ZN({ S2161 })
);
NAND2_X1 #() 
NAND2_X1_5028_ (
  .A1({ S1708 }),
  .A2({ S22985 }),
  .ZN({ S2162 })
);
OAI221_X1 #() 
OAI221_X1_147_ (
  .A({ S25957[917] }),
  .B1({ S2159 }),
  .B2({ S2160 }),
  .C1({ S2161 }),
  .C2({ S2162 }),
  .ZN({ S2163 })
);
NOR3_X1 #() 
NOR3_X1_165_ (
  .A1({ S1968 }),
  .A2({ S1967 }),
  .A3({ S86 }),
  .ZN({ S2164 })
);
NAND2_X1 #() 
NAND2_X1_5029_ (
  .A1({ S1646 }),
  .A2({ S86 }),
  .ZN({ S2165 })
);
NAND3_X1 #() 
NAND3_X1_5413_ (
  .A1({ S1707 }),
  .A2({ S2165 }),
  .A3({ S22985 }),
  .ZN({ S2166 })
);
OAI211_X1 #() 
OAI211_X1_1763_ (
  .A({ S25608 }),
  .B({ S2166 }),
  .C1({ S2164 }),
  .C2({ S1813 }),
  .ZN({ S2167 })
);
NAND3_X1 #() 
NAND3_X1_5414_ (
  .A1({ S2163 }),
  .A2({ S2167 }),
  .A3({ S25957[918] }),
  .ZN({ S2168 })
);
NAND3_X1 #() 
NAND3_X1_5415_ (
  .A1({ S2168 }),
  .A2({ S25957[919] }),
  .A3({ S2158 }),
  .ZN({ S2169 })
);
OAI21_X1 #() 
OAI21_X1_2613_ (
  .A({ S1825 }),
  .B1({ S1883 }),
  .B2({ S1628 }),
  .ZN({ S2170 })
);
NAND2_X1 #() 
NAND2_X1_5030_ (
  .A1({ S2170 }),
  .A2({ S25957[916] }),
  .ZN({ S2171 })
);
OAI21_X1 #() 
OAI21_X1_2614_ (
  .A({ S22985 }),
  .B1({ S1975 }),
  .B2({ S25921 }),
  .ZN({ S2172 })
);
OAI211_X1 #() 
OAI211_X1_1764_ (
  .A({ S25957[917] }),
  .B({ S2171 }),
  .C1({ S1659 }),
  .C2({ S2172 }),
  .ZN({ S2173 })
);
NAND4_X1 #() 
NAND4_X1_585_ (
  .A1({ S1639 }),
  .A2({ S1642 }),
  .A3({ S1624 }),
  .A4({ S1627 }),
  .ZN({ S2174 })
);
AOI22_X1 #() 
AOI22_X1_570_ (
  .A1({ S2174 }),
  .A2({ S86 }),
  .B1({ S1698 }),
  .B2({ S1788 }),
  .ZN({ S2175 })
);
NAND3_X1 #() 
NAND3_X1_5416_ (
  .A1({ S1899 }),
  .A2({ S1898 }),
  .A3({ S86 }),
  .ZN({ S2176 })
);
NAND3_X1 #() 
NAND3_X1_5417_ (
  .A1({ S2176 }),
  .A2({ S22985 }),
  .A3({ S2154 }),
  .ZN({ S2177 })
);
OAI211_X1 #() 
OAI211_X1_1765_ (
  .A({ S2177 }),
  .B({ S25608 }),
  .C1({ S2175 }),
  .C2({ S22985 }),
  .ZN({ S2178 })
);
AND3_X1 #() 
AND3_X1_212_ (
  .A1({ S2178 }),
  .A2({ S2173 }),
  .A3({ S25957[918] }),
  .ZN({ S2179 })
);
NAND4_X1 #() 
NAND4_X1_586_ (
  .A1({ S1790 }),
  .A2({ S1627 }),
  .A3({ S1642 }),
  .A4({ S25957[915] }),
  .ZN({ S2180 })
);
NAND2_X1 #() 
NAND2_X1_5031_ (
  .A1({ S2180 }),
  .A2({ S1785 }),
  .ZN({ S2181 })
);
OAI211_X1 #() 
OAI211_X1_1766_ (
  .A({ S1623 }),
  .B({ S25957[915] }),
  .C1({ S1627 }),
  .C2({ S25957[912] }),
  .ZN({ S2182 })
);
OAI211_X1 #() 
OAI211_X1_1767_ (
  .A({ S25957[916] }),
  .B({ S2182 }),
  .C1({ S1715 }),
  .C2({ S1737 }),
  .ZN({ S2183 })
);
OAI211_X1 #() 
OAI211_X1_1768_ (
  .A({ S2183 }),
  .B({ S25957[917] }),
  .C1({ S2181 }),
  .C2({ S25957[916] }),
  .ZN({ S2184 })
);
OAI211_X1 #() 
OAI211_X1_1769_ (
  .A({ S25957[916] }),
  .B({ S2154 }),
  .C1({ S1892 }),
  .C2({ S1687 }),
  .ZN({ S2185 })
);
NAND3_X1 #() 
NAND3_X1_5418_ (
  .A1({ S1752 }),
  .A2({ S22985 }),
  .A3({ S2025 }),
  .ZN({ S2186 })
);
NAND3_X1 #() 
NAND3_X1_5419_ (
  .A1({ S2186 }),
  .A2({ S25608 }),
  .A3({ S2185 }),
  .ZN({ S2187 })
);
AOI21_X1 #() 
AOI21_X1_2830_ (
  .A({ S25957[918] }),
  .B1({ S2184 }),
  .B2({ S2187 }),
  .ZN({ S2188 })
);
OAI21_X1 #() 
OAI21_X1_2615_ (
  .A({ S1685 }),
  .B1({ S2179 }),
  .B2({ S2188 }),
  .ZN({ S2189 })
);
NAND3_X1 #() 
NAND3_X1_5420_ (
  .A1({ S2189 }),
  .A2({ S25957[1018] }),
  .A3({ S2169 }),
  .ZN({ S2190 })
);
INV_X1 #() 
INV_X1_1639_ (
  .A({ S25957[1018] }),
  .ZN({ S2191 })
);
NAND2_X1 #() 
NAND2_X1_5032_ (
  .A1({ S2181 }),
  .A2({ S22985 }),
  .ZN({ S2192 })
);
AOI21_X1 #() 
AOI21_X1_2831_ (
  .A({ S1737 }),
  .B1({ S1656 }),
  .B2({ S106 }),
  .ZN({ S2193 })
);
AOI21_X1 #() 
AOI21_X1_2832_ (
  .A({ S86 }),
  .B1({ S1825 }),
  .B2({ S1661 }),
  .ZN({ S2194 })
);
OAI21_X1 #() 
OAI21_X1_2616_ (
  .A({ S25957[916] }),
  .B1({ S2193 }),
  .B2({ S2194 }),
  .ZN({ S2195 })
);
NAND3_X1 #() 
NAND3_X1_5421_ (
  .A1({ S2192 }),
  .A2({ S2195 }),
  .A3({ S22836 }),
  .ZN({ S2196 })
);
OAI211_X1 #() 
OAI211_X1_1770_ (
  .A({ S25957[918] }),
  .B({ S2171 }),
  .C1({ S1659 }),
  .C2({ S2172 }),
  .ZN({ S2197 })
);
AOI21_X1 #() 
AOI21_X1_2833_ (
  .A({ S25957[919] }),
  .B1({ S2196 }),
  .B2({ S2197 }),
  .ZN({ S2198 })
);
NOR2_X1 #() 
NOR2_X1_1282_ (
  .A1({ S2159 }),
  .A2({ S2160 }),
  .ZN({ S2199 })
);
AOI21_X1 #() 
AOI21_X1_2834_ (
  .A({ S2162 }),
  .B1({ S1928 }),
  .B2({ S25957[915] }),
  .ZN({ S2200 })
);
OAI21_X1 #() 
OAI21_X1_2617_ (
  .A({ S25957[918] }),
  .B1({ S2200 }),
  .B2({ S2199 }),
  .ZN({ S2201 })
);
AOI22_X1 #() 
AOI22_X1_571_ (
  .A1({ S1768 }),
  .A2({ S1693 }),
  .B1({ S2146 }),
  .B2({ S25957[915] }),
  .ZN({ S2202 })
);
OAI21_X1 #() 
OAI21_X1_2618_ (
  .A({ S22985 }),
  .B1({ S2151 }),
  .B2({ S1984 }),
  .ZN({ S2203 })
);
OAI211_X1 #() 
OAI211_X1_1771_ (
  .A({ S2203 }),
  .B({ S22836 }),
  .C1({ S2202 }),
  .C2({ S22985 }),
  .ZN({ S2204 })
);
AOI21_X1 #() 
AOI21_X1_2835_ (
  .A({ S1685 }),
  .B1({ S2201 }),
  .B2({ S2204 }),
  .ZN({ S2205 })
);
OAI21_X1 #() 
OAI21_X1_2619_ (
  .A({ S25957[917] }),
  .B1({ S2205 }),
  .B2({ S2198 }),
  .ZN({ S2206 })
);
AOI21_X1 #() 
AOI21_X1_2836_ (
  .A({ S1813 }),
  .B1({ S1667 }),
  .B2({ S25957[915] }),
  .ZN({ S2207 })
);
INV_X1 #() 
INV_X1_1640_ (
  .A({ S2166 }),
  .ZN({ S2208 })
);
OAI21_X1 #() 
OAI21_X1_2620_ (
  .A({ S25957[918] }),
  .B1({ S2207 }),
  .B2({ S2208 }),
  .ZN({ S2209 })
);
NAND2_X1 #() 
NAND2_X1_5033_ (
  .A1({ S2156 }),
  .A2({ S2155 }),
  .ZN({ S2210 })
);
NAND2_X1 #() 
NAND2_X1_5034_ (
  .A1({ S2210 }),
  .A2({ S22836 }),
  .ZN({ S2211 })
);
AOI21_X1 #() 
AOI21_X1_2837_ (
  .A({ S1685 }),
  .B1({ S2209 }),
  .B2({ S2211 }),
  .ZN({ S2212 })
);
NAND2_X1 #() 
NAND2_X1_5035_ (
  .A1({ S2186 }),
  .A2({ S2185 }),
  .ZN({ S2213 })
);
NAND2_X1 #() 
NAND2_X1_5036_ (
  .A1({ S2213 }),
  .A2({ S22836 }),
  .ZN({ S2214 })
);
OAI211_X1 #() 
OAI211_X1_1772_ (
  .A({ S2177 }),
  .B({ S25957[918] }),
  .C1({ S2175 }),
  .C2({ S22985 }),
  .ZN({ S2215 })
);
AOI21_X1 #() 
AOI21_X1_2838_ (
  .A({ S25957[919] }),
  .B1({ S2214 }),
  .B2({ S2215 }),
  .ZN({ S2216 })
);
OAI21_X1 #() 
OAI21_X1_2621_ (
  .A({ S25608 }),
  .B1({ S2216 }),
  .B2({ S2212 }),
  .ZN({ S2217 })
);
NAND3_X1 #() 
NAND3_X1_5422_ (
  .A1({ S2217 }),
  .A2({ S2206 }),
  .A3({ S2191 }),
  .ZN({ S2218 })
);
NAND3_X1 #() 
NAND3_X1_5423_ (
  .A1({ S2218 }),
  .A2({ S25957[986] }),
  .A3({ S2190 }),
  .ZN({ S2219 })
);
NAND3_X1 #() 
NAND3_X1_5424_ (
  .A1({ S2189 }),
  .A2({ S2191 }),
  .A3({ S2169 }),
  .ZN({ S2220 })
);
NAND3_X1 #() 
NAND3_X1_5425_ (
  .A1({ S2217 }),
  .A2({ S2206 }),
  .A3({ S25957[1018] }),
  .ZN({ S2221 })
);
NAND3_X1 #() 
NAND3_X1_5426_ (
  .A1({ S2221 }),
  .A2({ S2145 }),
  .A3({ S2220 }),
  .ZN({ S2222 })
);
NAND3_X1 #() 
NAND3_X1_5427_ (
  .A1({ S2219 }),
  .A2({ S2222 }),
  .A3({ S2144 }),
  .ZN({ S2223 })
);
NAND3_X1 #() 
NAND3_X1_5428_ (
  .A1({ S2221 }),
  .A2({ S25957[986] }),
  .A3({ S2220 }),
  .ZN({ S2224 })
);
NAND3_X1 #() 
NAND3_X1_5429_ (
  .A1({ S2218 }),
  .A2({ S2145 }),
  .A3({ S2190 }),
  .ZN({ S2225 })
);
NAND3_X1 #() 
NAND3_X1_5430_ (
  .A1({ S2224 }),
  .A2({ S2225 }),
  .A3({ S25957[954] }),
  .ZN({ S2226 })
);
NAND3_X1 #() 
NAND3_X1_5431_ (
  .A1({ S2223 }),
  .A2({ S2226 }),
  .A3({ S25957[922] }),
  .ZN({ S2227 })
);
NAND3_X1 #() 
NAND3_X1_5432_ (
  .A1({ S2219 }),
  .A2({ S2222 }),
  .A3({ S25957[954] }),
  .ZN({ S2228 })
);
NAND3_X1 #() 
NAND3_X1_5433_ (
  .A1({ S2224 }),
  .A2({ S2225 }),
  .A3({ S2144 }),
  .ZN({ S2229 })
);
NAND3_X1 #() 
NAND3_X1_5434_ (
  .A1({ S2228 }),
  .A2({ S2229 }),
  .A3({ S1033 }),
  .ZN({ S2230 })
);
NAND2_X1 #() 
NAND2_X1_5037_ (
  .A1({ S2227 }),
  .A2({ S2230 }),
  .ZN({ S25957[794] })
);
AOI21_X1 #() 
AOI21_X1_2839_ (
  .A({ S25957[1032] }),
  .B1({ S867 }),
  .B2({ S868 }),
  .ZN({ S2231 })
);
AOI21_X1 #() 
AOI21_X1_2840_ (
  .A({ S22633 }),
  .B1({ S861 }),
  .B2({ S865 }),
  .ZN({ S2232 })
);
AOI21_X1 #() 
AOI21_X1_2841_ (
  .A({ S25957[969] }),
  .B1({ S943 }),
  .B2({ S942 }),
  .ZN({ S2233 })
);
AOI21_X1 #() 
AOI21_X1_2842_ (
  .A({ S870 }),
  .B1({ S940 }),
  .B2({ S911 }),
  .ZN({ S2234 })
);
OAI21_X1 #() 
OAI21_X1_2622_ (
  .A({ S22634 }),
  .B1({ S2233 }),
  .B2({ S2234 }),
  .ZN({ S2235 })
);
NAND3_X1 #() 
NAND3_X1_5435_ (
  .A1({ S941 }),
  .A2({ S944 }),
  .A3({ S25957[1033] }),
  .ZN({ S2236 })
);
OAI211_X1 #() 
OAI211_X1_1773_ (
  .A({ S2235 }),
  .B({ S2236 }),
  .C1({ S2232 }),
  .C2({ S2231 }),
  .ZN({ S2237 })
);
INV_X1 #() 
INV_X1_1641_ (
  .A({ S2237 }),
  .ZN({ S108 })
);
OAI211_X1 #() 
OAI211_X1_1774_ (
  .A({ S866 }),
  .B({ S869 }),
  .C1({ S946 }),
  .C2({ S945 }),
  .ZN({ S109 })
);
XOR2_X1 #() 
XOR2_X1_81_ (
  .A({ S25957[855] }),
  .B({ S25957[951] }),
  .Z({ S25957[823] })
);
INV_X1 #() 
INV_X1_1642_ (
  .A({ S25957[823] }),
  .ZN({ S2238 })
);
XNOR2_X1 #() 
XNOR2_X1_196_ (
  .A({ S22749 }),
  .B({ S25957[1143] }),
  .ZN({ S25957[1015] })
);
XOR2_X1 #() 
XOR2_X1_82_ (
  .A({ S25525 }),
  .B({ S25957[1015] }),
  .Z({ S25957[887] })
);
INV_X1 #() 
INV_X1_1643_ (
  .A({ S25957[887] }),
  .ZN({ S2239 })
);
NAND3_X1 #() 
NAND3_X1_5436_ (
  .A1({ S2237 }),
  .A2({ S109 }),
  .A3({ S25957[778] }),
  .ZN({ S2240 })
);
NAND3_X1 #() 
NAND3_X1_5437_ (
  .A1({ S1011 }),
  .A2({ S1012 }),
  .A3({ S25957[906] }),
  .ZN({ S2241 })
);
NAND3_X1 #() 
NAND3_X1_5438_ (
  .A1({ S1006 }),
  .A2({ S1009 }),
  .A3({ S25436 }),
  .ZN({ S2242 })
);
NAND2_X1 #() 
NAND2_X1_5038_ (
  .A1({ S2241 }),
  .A2({ S2242 }),
  .ZN({ S2243 })
);
OAI22_X1 #() 
OAI22_X1_127_ (
  .A1({ S2231 }),
  .A2({ S2232 }),
  .B1({ S946 }),
  .B2({ S945 }),
  .ZN({ S2244 })
);
NAND4_X1 #() 
NAND4_X1_587_ (
  .A1({ S2235 }),
  .A2({ S866 }),
  .A3({ S869 }),
  .A4({ S2236 }),
  .ZN({ S2245 })
);
NAND3_X1 #() 
NAND3_X1_5439_ (
  .A1({ S2244 }),
  .A2({ S2243 }),
  .A3({ S2245 }),
  .ZN({ S2246 })
);
AOI21_X1 #() 
AOI21_X1_2843_ (
  .A({ S101 }),
  .B1({ S2240 }),
  .B2({ S2246 }),
  .ZN({ S2247 })
);
NAND4_X1 #() 
NAND4_X1_588_ (
  .A1({ S2242 }),
  .A2({ S2235 }),
  .A3({ S2241 }),
  .A4({ S2236 }),
  .ZN({ S2248 })
);
INV_X1 #() 
INV_X1_1644_ (
  .A({ S2248 }),
  .ZN({ S2249 })
);
OAI211_X1 #() 
OAI211_X1_1775_ (
  .A({ S1010 }),
  .B({ S1013 }),
  .C1({ S2232 }),
  .C2({ S2231 }),
  .ZN({ S2250 })
);
NAND2_X1 #() 
NAND2_X1_5039_ (
  .A1({ S2250 }),
  .A2({ S101 }),
  .ZN({ S2251 })
);
NOR2_X1 #() 
NOR2_X1_1283_ (
  .A1({ S2251 }),
  .A2({ S2249 }),
  .ZN({ S2252 })
);
OAI21_X1 #() 
OAI21_X1_2623_ (
  .A({ S25957[780] }),
  .B1({ S2247 }),
  .B2({ S2252 }),
  .ZN({ S2253 })
);
OAI21_X1 #() 
OAI21_X1_2624_ (
  .A({ S25416 }),
  .B1({ S706 }),
  .B2({ S709 }),
  .ZN({ S2254 })
);
NAND3_X1 #() 
NAND3_X1_5440_ (
  .A1({ S711 }),
  .A2({ S712 }),
  .A3({ S25957[908] }),
  .ZN({ S2255 })
);
NAND2_X1 #() 
NAND2_X1_5040_ (
  .A1({ S2254 }),
  .A2({ S2255 }),
  .ZN({ S2256 })
);
NAND3_X1 #() 
NAND3_X1_5441_ (
  .A1({ S25957[777] }),
  .A2({ S2243 }),
  .A3({ S25957[776] }),
  .ZN({ S2257 })
);
NAND2_X1 #() 
NAND2_X1_5041_ (
  .A1({ S2235 }),
  .A2({ S2236 }),
  .ZN({ S2258 })
);
NAND2_X1 #() 
NAND2_X1_5042_ (
  .A1({ S2250 }),
  .A2({ S2258 }),
  .ZN({ S2259 })
);
NAND2_X1 #() 
NAND2_X1_5043_ (
  .A1({ S2259 }),
  .A2({ S2257 }),
  .ZN({ S2260 })
);
INV_X1 #() 
INV_X1_1645_ (
  .A({ S2260 }),
  .ZN({ S2261 })
);
NAND4_X1 #() 
NAND4_X1_589_ (
  .A1({ S2241 }),
  .A2({ S2242 }),
  .A3({ S866 }),
  .A4({ S869 }),
  .ZN({ S2262 })
);
NAND2_X1 #() 
NAND2_X1_5044_ (
  .A1({ S2262 }),
  .A2({ S101 }),
  .ZN({ S2263 })
);
AOI22_X1 #() 
AOI22_X1_572_ (
  .A1({ S2242 }),
  .A2({ S2241 }),
  .B1({ S2235 }),
  .B2({ S2236 }),
  .ZN({ S2264 })
);
NAND2_X1 #() 
NAND2_X1_5045_ (
  .A1({ S2264 }),
  .A2({ S25957[779] }),
  .ZN({ S2265 })
);
OAI211_X1 #() 
OAI211_X1_1776_ (
  .A({ S2256 }),
  .B({ S2265 }),
  .C1({ S2261 }),
  .C2({ S2263 }),
  .ZN({ S2266 })
);
AOI21_X1 #() 
AOI21_X1_2844_ (
  .A({ S25957[781] }),
  .B1({ S2266 }),
  .B2({ S2253 }),
  .ZN({ S2267 })
);
INV_X1 #() 
INV_X1_1646_ (
  .A({ S25957[782] }),
  .ZN({ S2268 })
);
AOI22_X1 #() 
AOI22_X1_573_ (
  .A1({ S1010 }),
  .A2({ S1013 }),
  .B1({ S869 }),
  .B2({ S866 }),
  .ZN({ S2269 })
);
NAND2_X1 #() 
NAND2_X1_5046_ (
  .A1({ S101 }),
  .A2({ S25957[777] }),
  .ZN({ S2270 })
);
OAI21_X1 #() 
OAI21_X1_2625_ (
  .A({ S25957[779] }),
  .B1({ S2269 }),
  .B2({ S2258 }),
  .ZN({ S2271 })
);
OAI211_X1 #() 
OAI211_X1_1777_ (
  .A({ S2271 }),
  .B({ S25957[780] }),
  .C1({ S2269 }),
  .C2({ S2270 }),
  .ZN({ S2272 })
);
NAND4_X1 #() 
NAND4_X1_590_ (
  .A1({ S1010 }),
  .A2({ S1013 }),
  .A3({ S866 }),
  .A4({ S869 }),
  .ZN({ S2273 })
);
OAI21_X1 #() 
OAI21_X1_2626_ (
  .A({ S101 }),
  .B1({ S2273 }),
  .B2({ S25957[777] }),
  .ZN({ S2274 })
);
NOR2_X1 #() 
NOR2_X1_1284_ (
  .A1({ S2237 }),
  .A2({ S101 }),
  .ZN({ S2275 })
);
INV_X1 #() 
INV_X1_1647_ (
  .A({ S2275 }),
  .ZN({ S2276 })
);
NAND3_X1 #() 
NAND3_X1_5442_ (
  .A1({ S2276 }),
  .A2({ S2256 }),
  .A3({ S2274 }),
  .ZN({ S2277 })
);
NAND3_X1 #() 
NAND3_X1_5443_ (
  .A1({ S2277 }),
  .A2({ S2272 }),
  .A3({ S25957[781] }),
  .ZN({ S2278 })
);
NAND2_X1 #() 
NAND2_X1_5047_ (
  .A1({ S2278 }),
  .A2({ S2268 }),
  .ZN({ S2279 })
);
AOI22_X1 #() 
AOI22_X1_574_ (
  .A1({ S2235 }),
  .A2({ S2236 }),
  .B1({ S869 }),
  .B2({ S866 }),
  .ZN({ S2280 })
);
NAND2_X1 #() 
NAND2_X1_5048_ (
  .A1({ S109 }),
  .A2({ S2243 }),
  .ZN({ S2281 })
);
NOR2_X1 #() 
NOR2_X1_1285_ (
  .A1({ S2231 }),
  .A2({ S2232 }),
  .ZN({ S2282 })
);
NAND3_X1 #() 
NAND3_X1_5444_ (
  .A1({ S2282 }),
  .A2({ S2258 }),
  .A3({ S25957[778] }),
  .ZN({ S2283 })
);
AOI22_X1 #() 
AOI22_X1_575_ (
  .A1({ S2281 }),
  .A2({ S2283 }),
  .B1({ S2280 }),
  .B2({ S25957[779] }),
  .ZN({ S2284 })
);
OAI211_X1 #() 
OAI211_X1_1778_ (
  .A({ S2241 }),
  .B({ S2242 }),
  .C1({ S946 }),
  .C2({ S945 }),
  .ZN({ S2285 })
);
NAND3_X1 #() 
NAND3_X1_5445_ (
  .A1({ S2237 }),
  .A2({ S2285 }),
  .A3({ S25957[779] }),
  .ZN({ S2286 })
);
NAND2_X1 #() 
NAND2_X1_5049_ (
  .A1({ S2245 }),
  .A2({ S101 }),
  .ZN({ S2287 })
);
NAND3_X1 #() 
NAND3_X1_5446_ (
  .A1({ S2286 }),
  .A2({ S25957[780] }),
  .A3({ S2287 }),
  .ZN({ S2288 })
);
OAI21_X1 #() 
OAI21_X1_2627_ (
  .A({ S2288 }),
  .B1({ S2284 }),
  .B2({ S25957[780] }),
  .ZN({ S2289 })
);
NAND3_X1 #() 
NAND3_X1_5447_ (
  .A1({ S2282 }),
  .A2({ S25957[777] }),
  .A3({ S25957[778] }),
  .ZN({ S2290 })
);
NOR2_X1 #() 
NOR2_X1_1286_ (
  .A1({ S25957[780] }),
  .A2({ S101 }),
  .ZN({ S2291 })
);
NAND3_X1 #() 
NAND3_X1_5448_ (
  .A1({ S2291 }),
  .A2({ S2244 }),
  .A3({ S2290 }),
  .ZN({ S2292 })
);
NOR2_X1 #() 
NOR2_X1_1287_ (
  .A1({ S25957[780] }),
  .A2({ S25957[779] }),
  .ZN({ S2293 })
);
NAND3_X1 #() 
NAND3_X1_5449_ (
  .A1({ S2293 }),
  .A2({ S2257 }),
  .A3({ S2283 }),
  .ZN({ S2294 })
);
NAND2_X1 #() 
NAND2_X1_5050_ (
  .A1({ S2292 }),
  .A2({ S2294 }),
  .ZN({ S2295 })
);
NAND3_X1 #() 
NAND3_X1_5450_ (
  .A1({ S2243 }),
  .A2({ S2258 }),
  .A3({ S25957[776] }),
  .ZN({ S2296 })
);
INV_X1 #() 
INV_X1_1648_ (
  .A({ S2296 }),
  .ZN({ S2297 })
);
NAND2_X1 #() 
NAND2_X1_5051_ (
  .A1({ S2273 }),
  .A2({ S101 }),
  .ZN({ S2298 })
);
NAND2_X1 #() 
NAND2_X1_5052_ (
  .A1({ S2262 }),
  .A2({ S25957[779] }),
  .ZN({ S2299 })
);
OAI22_X1 #() 
OAI22_X1_128_ (
  .A1({ S2297 }),
  .A2({ S2299 }),
  .B1({ S2298 }),
  .B2({ S2258 }),
  .ZN({ S2300 })
);
OAI21_X1 #() 
OAI21_X1_2628_ (
  .A({ S25957[781] }),
  .B1({ S2300 }),
  .B2({ S2256 }),
  .ZN({ S2301 })
);
OAI221_X1 #() 
OAI221_X1_148_ (
  .A({ S25957[782] }),
  .B1({ S2289 }),
  .B2({ S25957[781] }),
  .C1({ S2301 }),
  .C2({ S2295 }),
  .ZN({ S2302 })
);
OAI21_X1 #() 
OAI21_X1_2629_ (
  .A({ S2302 }),
  .B1({ S2279 }),
  .B2({ S2267 }),
  .ZN({ S2303 })
);
NAND2_X1 #() 
NAND2_X1_5053_ (
  .A1({ S2303 }),
  .A2({ S25957[783] }),
  .ZN({ S2304 })
);
INV_X1 #() 
INV_X1_1649_ (
  .A({ S25957[783] }),
  .ZN({ S2305 })
);
NAND2_X1 #() 
NAND2_X1_5054_ (
  .A1({ S2256 }),
  .A2({ S25957[779] }),
  .ZN({ S2306 })
);
NOR2_X1 #() 
NOR2_X1_1288_ (
  .A1({ S2250 }),
  .A2({ S2258 }),
  .ZN({ S2307 })
);
OAI21_X1 #() 
OAI21_X1_2630_ (
  .A({ S25957[779] }),
  .B1({ S2262 }),
  .B2({ S25957[777] }),
  .ZN({ S2308 })
);
INV_X1 #() 
INV_X1_1650_ (
  .A({ S2298 }),
  .ZN({ S2309 })
);
AOI21_X1 #() 
AOI21_X1_2845_ (
  .A({ S2256 }),
  .B1({ S2309 }),
  .B2({ S2290 }),
  .ZN({ S2310 })
);
OAI21_X1 #() 
OAI21_X1_2631_ (
  .A({ S2310 }),
  .B1({ S2307 }),
  .B2({ S2308 }),
  .ZN({ S2311 })
);
NAND2_X1 #() 
NAND2_X1_5055_ (
  .A1({ S2244 }),
  .A2({ S2243 }),
  .ZN({ S2312 })
);
NAND2_X1 #() 
NAND2_X1_5056_ (
  .A1({ S2312 }),
  .A2({ S2285 }),
  .ZN({ S2313 })
);
INV_X1 #() 
INV_X1_1651_ (
  .A({ S2313 }),
  .ZN({ S2314 })
);
INV_X1 #() 
INV_X1_1652_ (
  .A({ S25957[781] }),
  .ZN({ S2315 })
);
NAND2_X1 #() 
NAND2_X1_5057_ (
  .A1({ S2237 }),
  .A2({ S25957[778] }),
  .ZN({ S2316 })
);
INV_X1 #() 
INV_X1_1653_ (
  .A({ S2316 }),
  .ZN({ S2317 })
);
AOI21_X1 #() 
AOI21_X1_2846_ (
  .A({ S2315 }),
  .B1({ S2317 }),
  .B2({ S2293 }),
  .ZN({ S2318 })
);
OAI211_X1 #() 
OAI211_X1_1779_ (
  .A({ S2311 }),
  .B({ S2318 }),
  .C1({ S2306 }),
  .C2({ S2314 }),
  .ZN({ S2319 })
);
NAND4_X1 #() 
NAND4_X1_591_ (
  .A1({ S1013 }),
  .A2({ S2235 }),
  .A3({ S1010 }),
  .A4({ S2236 }),
  .ZN({ S2320 })
);
NOR2_X1 #() 
NOR2_X1_1289_ (
  .A1({ S2269 }),
  .A2({ S101 }),
  .ZN({ S2321 })
);
NAND2_X1 #() 
NAND2_X1_5058_ (
  .A1({ S2321 }),
  .A2({ S2320 }),
  .ZN({ S2322 })
);
NAND3_X1 #() 
NAND3_X1_5451_ (
  .A1({ S2285 }),
  .A2({ S2320 }),
  .A3({ S25957[776] }),
  .ZN({ S2323 })
);
AOI21_X1 #() 
AOI21_X1_2847_ (
  .A({ S25957[780] }),
  .B1({ S2323 }),
  .B2({ S101 }),
  .ZN({ S2324 })
);
AOI21_X1 #() 
AOI21_X1_2848_ (
  .A({ S101 }),
  .B1({ S2246 }),
  .B2({ S2316 }),
  .ZN({ S2325 })
);
NAND3_X1 #() 
NAND3_X1_5452_ (
  .A1({ S2244 }),
  .A2({ S25957[778] }),
  .A3({ S2245 }),
  .ZN({ S2326 })
);
AOI21_X1 #() 
AOI21_X1_2849_ (
  .A({ S25957[779] }),
  .B1({ S2326 }),
  .B2({ S2273 }),
  .ZN({ S2327 })
);
NOR3_X1 #() 
NOR3_X1_166_ (
  .A1({ S2327 }),
  .A2({ S2325 }),
  .A3({ S2256 }),
  .ZN({ S2328 })
);
AOI21_X1 #() 
AOI21_X1_2850_ (
  .A({ S2328 }),
  .B1({ S2324 }),
  .B2({ S2322 }),
  .ZN({ S2329 })
);
OAI21_X1 #() 
OAI21_X1_2632_ (
  .A({ S2319 }),
  .B1({ S2329 }),
  .B2({ S25957[781] }),
  .ZN({ S2330 })
);
NAND2_X1 #() 
NAND2_X1_5059_ (
  .A1({ S2237 }),
  .A2({ S2243 }),
  .ZN({ S2331 })
);
INV_X1 #() 
INV_X1_1654_ (
  .A({ S2331 }),
  .ZN({ S2332 })
);
NAND2_X1 #() 
NAND2_X1_5060_ (
  .A1({ S2248 }),
  .A2({ S101 }),
  .ZN({ S2333 })
);
NOR2_X1 #() 
NOR2_X1_1290_ (
  .A1({ S2280 }),
  .A2({ S101 }),
  .ZN({ S2334 })
);
NAND2_X1 #() 
NAND2_X1_5061_ (
  .A1({ S2334 }),
  .A2({ S2320 }),
  .ZN({ S2335 })
);
OAI21_X1 #() 
OAI21_X1_2633_ (
  .A({ S2335 }),
  .B1({ S2332 }),
  .B2({ S2333 }),
  .ZN({ S2336 })
);
NAND2_X1 #() 
NAND2_X1_5062_ (
  .A1({ S101 }),
  .A2({ S25957[776] }),
  .ZN({ S2337 })
);
NAND2_X1 #() 
NAND2_X1_5063_ (
  .A1({ S2243 }),
  .A2({ S2258 }),
  .ZN({ S2338 })
);
NAND2_X1 #() 
NAND2_X1_5064_ (
  .A1({ S2321 }),
  .A2({ S2338 }),
  .ZN({ S2339 })
);
AND3_X1 #() 
AND3_X1_213_ (
  .A1({ S2339 }),
  .A2({ S2337 }),
  .A3({ S25957[780] }),
  .ZN({ S2340 })
);
AOI211_X1 #() 
AOI211_X1_87_ (
  .A({ S2315 }),
  .B({ S2340 }),
  .C1({ S2256 }),
  .C2({ S2336 }),
  .ZN({ S2341 })
);
AOI21_X1 #() 
AOI21_X1_2851_ (
  .A({ S2243 }),
  .B1({ S2244 }),
  .B2({ S2245 }),
  .ZN({ S2342 })
);
NAND2_X1 #() 
NAND2_X1_5065_ (
  .A1({ S2257 }),
  .A2({ S101 }),
  .ZN({ S2343 })
);
NOR2_X1 #() 
NOR2_X1_1291_ (
  .A1({ S2343 }),
  .A2({ S2342 }),
  .ZN({ S2344 })
);
NAND4_X1 #() 
NAND4_X1_592_ (
  .A1({ S2244 }),
  .A2({ S2245 }),
  .A3({ S101 }),
  .A4({ S25957[778] }),
  .ZN({ S2345 })
);
OAI211_X1 #() 
OAI211_X1_1780_ (
  .A({ S2345 }),
  .B({ S2256 }),
  .C1({ S101 }),
  .C2({ S2316 }),
  .ZN({ S2346 })
);
INV_X1 #() 
INV_X1_1655_ (
  .A({ S2290 }),
  .ZN({ S2347 })
);
OAI21_X1 #() 
OAI21_X1_2634_ (
  .A({ S25957[780] }),
  .B1({ S2347 }),
  .B2({ S101 }),
  .ZN({ S2348 })
);
OAI211_X1 #() 
OAI211_X1_1781_ (
  .A({ S2315 }),
  .B({ S2346 }),
  .C1({ S2348 }),
  .C2({ S2344 }),
  .ZN({ S2349 })
);
NAND2_X1 #() 
NAND2_X1_5066_ (
  .A1({ S2349 }),
  .A2({ S2268 }),
  .ZN({ S2350 })
);
OAI221_X1 #() 
OAI221_X1_149_ (
  .A({ S2305 }),
  .B1({ S2330 }),
  .B2({ S2268 }),
  .C1({ S2350 }),
  .C2({ S2341 }),
  .ZN({ S2351 })
);
NAND2_X1 #() 
NAND2_X1_5067_ (
  .A1({ S2351 }),
  .A2({ S2304 }),
  .ZN({ S2352 })
);
NAND2_X1 #() 
NAND2_X1_5068_ (
  .A1({ S2352 }),
  .A2({ S2239 }),
  .ZN({ S2353 })
);
NAND3_X1 #() 
NAND3_X1_5453_ (
  .A1({ S2351 }),
  .A2({ S25957[887] }),
  .A3({ S2304 }),
  .ZN({ S2354 })
);
NAND2_X1 #() 
NAND2_X1_5069_ (
  .A1({ S2353 }),
  .A2({ S2354 }),
  .ZN({ S25957[759] })
);
NAND2_X1 #() 
NAND2_X1_5070_ (
  .A1({ S25957[759] }),
  .A2({ S25527 }),
  .ZN({ S2355 })
);
INV_X1 #() 
INV_X1_1656_ (
  .A({ S25957[759] }),
  .ZN({ S2356 })
);
NAND2_X1 #() 
NAND2_X1_5071_ (
  .A1({ S2356 }),
  .A2({ S25957[855] }),
  .ZN({ S2357 })
);
NAND2_X1 #() 
NAND2_X1_5072_ (
  .A1({ S2357 }),
  .A2({ S2355 }),
  .ZN({ S25957[727] })
);
NAND2_X1 #() 
NAND2_X1_5073_ (
  .A1({ S25957[727] }),
  .A2({ S2238 }),
  .ZN({ S2358 })
);
NAND3_X1 #() 
NAND3_X1_5454_ (
  .A1({ S2357 }),
  .A2({ S25957[823] }),
  .A3({ S2355 }),
  .ZN({ S2359 })
);
NAND3_X1 #() 
NAND3_X1_5455_ (
  .A1({ S2358 }),
  .A2({ S2359 }),
  .A3({ S25957[791] }),
  .ZN({ S2360 })
);
INV_X1 #() 
INV_X1_1657_ (
  .A({ S25957[791] }),
  .ZN({ S2361 })
);
NAND2_X1 #() 
NAND2_X1_5074_ (
  .A1({ S2358 }),
  .A2({ S2359 }),
  .ZN({ S25957[695] })
);
NAND2_X1 #() 
NAND2_X1_5075_ (
  .A1({ S25957[695] }),
  .A2({ S2361 }),
  .ZN({ S2362 })
);
NAND2_X1 #() 
NAND2_X1_5076_ (
  .A1({ S2362 }),
  .A2({ S2360 }),
  .ZN({ S25957[663] })
);
NAND2_X1 #() 
NAND2_X1_5077_ (
  .A1({ S22830 }),
  .A2({ S22829 }),
  .ZN({ S2363 })
);
INV_X1 #() 
INV_X1_1658_ (
  .A({ S2363 }),
  .ZN({ S25957[950] })
);
NAND2_X1 #() 
NAND2_X1_5078_ (
  .A1({ S22825 }),
  .A2({ S22796 }),
  .ZN({ S2364 })
);
XNOR2_X1 #() 
XNOR2_X1_197_ (
  .A({ S2364 }),
  .B({ S25957[1142] }),
  .ZN({ S25957[1014] })
);
XOR2_X1 #() 
XOR2_X1_83_ (
  .A({ S25602 }),
  .B({ S25957[1014] }),
  .Z({ S2365 })
);
INV_X1 #() 
INV_X1_1659_ (
  .A({ S2365 }),
  .ZN({ S25957[886] })
);
NAND2_X1 #() 
NAND2_X1_5079_ (
  .A1({ S2338 }),
  .A2({ S2282 }),
  .ZN({ S2366 })
);
INV_X1 #() 
INV_X1_1660_ (
  .A({ S2320 }),
  .ZN({ S2367 })
);
NAND2_X1 #() 
NAND2_X1_5080_ (
  .A1({ S2367 }),
  .A2({ S25957[779] }),
  .ZN({ S2368 })
);
OAI211_X1 #() 
OAI211_X1_1782_ (
  .A({ S2368 }),
  .B({ S25957[780] }),
  .C1({ S2366 }),
  .C2({ S25957[779] }),
  .ZN({ S2369 })
);
NAND3_X1 #() 
NAND3_X1_5456_ (
  .A1({ S2250 }),
  .A2({ S2248 }),
  .A3({ S2262 }),
  .ZN({ S2370 })
);
NAND2_X1 #() 
NAND2_X1_5081_ (
  .A1({ S2370 }),
  .A2({ S25957[779] }),
  .ZN({ S2371 })
);
OAI21_X1 #() 
OAI21_X1_2635_ (
  .A({ S2371 }),
  .B1({ S25957[779] }),
  .B2({ S2342 }),
  .ZN({ S2372 })
);
OAI21_X1 #() 
OAI21_X1_2636_ (
  .A({ S2369 }),
  .B1({ S2372 }),
  .B2({ S25957[780] }),
  .ZN({ S2373 })
);
OAI211_X1 #() 
OAI211_X1_1783_ (
  .A({ S2241 }),
  .B({ S2242 }),
  .C1({ S2232 }),
  .C2({ S2231 }),
  .ZN({ S2374 })
);
AOI21_X1 #() 
AOI21_X1_2852_ (
  .A({ S101 }),
  .B1({ S2374 }),
  .B2({ S2245 }),
  .ZN({ S2375 })
);
INV_X1 #() 
INV_X1_1661_ (
  .A({ S2250 }),
  .ZN({ S2376 })
);
NOR2_X1 #() 
NOR2_X1_1292_ (
  .A1({ S2376 }),
  .A2({ S2270 }),
  .ZN({ S2377 })
);
OR3_X1 #() 
OR3_X1_32_ (
  .A1({ S2377 }),
  .A2({ S2375 }),
  .A3({ S25957[780] }),
  .ZN({ S2378 })
);
NAND3_X1 #() 
NAND3_X1_5457_ (
  .A1({ S2285 }),
  .A2({ S2262 }),
  .A3({ S101 }),
  .ZN({ S2379 })
);
NOR2_X1 #() 
NOR2_X1_1293_ (
  .A1({ S2379 }),
  .A2({ S2376 }),
  .ZN({ S2380 })
);
OAI21_X1 #() 
OAI21_X1_2637_ (
  .A({ S25957[780] }),
  .B1({ S2380 }),
  .B2({ S2375 }),
  .ZN({ S2381 })
);
NAND3_X1 #() 
NAND3_X1_5458_ (
  .A1({ S2378 }),
  .A2({ S25957[781] }),
  .A3({ S2381 }),
  .ZN({ S2382 })
);
OAI21_X1 #() 
OAI21_X1_2638_ (
  .A({ S2382 }),
  .B1({ S2373 }),
  .B2({ S25957[781] }),
  .ZN({ S2383 })
);
INV_X1 #() 
INV_X1_1662_ (
  .A({ S2285 }),
  .ZN({ S2384 })
);
NOR2_X1 #() 
NOR2_X1_1294_ (
  .A1({ S2384 }),
  .A2({ S2367 }),
  .ZN({ S2385 })
);
INV_X1 #() 
INV_X1_1663_ (
  .A({ S2385 }),
  .ZN({ S2386 })
);
NAND3_X1 #() 
NAND3_X1_5459_ (
  .A1({ S2296 }),
  .A2({ S101 }),
  .A3({ S2248 }),
  .ZN({ S2387 })
);
OAI21_X1 #() 
OAI21_X1_2639_ (
  .A({ S2387 }),
  .B1({ S2386 }),
  .B2({ S101 }),
  .ZN({ S2388 })
);
NAND2_X1 #() 
NAND2_X1_5082_ (
  .A1({ S2283 }),
  .A2({ S2237 }),
  .ZN({ S2389 })
);
OAI211_X1 #() 
OAI211_X1_1784_ (
  .A({ S25957[780] }),
  .B({ S2251 }),
  .C1({ S2389 }),
  .C2({ S101 }),
  .ZN({ S2390 })
);
OAI211_X1 #() 
OAI211_X1_1785_ (
  .A({ S25957[781] }),
  .B({ S2390 }),
  .C1({ S2388 }),
  .C2({ S25957[780] }),
  .ZN({ S2391 })
);
NAND2_X1 #() 
NAND2_X1_5083_ (
  .A1({ S2313 }),
  .A2({ S25957[779] }),
  .ZN({ S2392 })
);
NAND2_X1 #() 
NAND2_X1_5084_ (
  .A1({ S2264 }),
  .A2({ S101 }),
  .ZN({ S2393 })
);
OAI21_X1 #() 
OAI21_X1_2640_ (
  .A({ S2392 }),
  .B1({ S2282 }),
  .B2({ S2393 }),
  .ZN({ S2394 })
);
NAND2_X1 #() 
NAND2_X1_5085_ (
  .A1({ S2245 }),
  .A2({ S2243 }),
  .ZN({ S2395 })
);
NAND2_X1 #() 
NAND2_X1_5086_ (
  .A1({ S2290 }),
  .A2({ S2395 }),
  .ZN({ S2396 })
);
AOI22_X1 #() 
AOI22_X1_576_ (
  .A1({ S2394 }),
  .A2({ S25957[780] }),
  .B1({ S2396 }),
  .B2({ S2291 }),
  .ZN({ S2397 })
);
OAI211_X1 #() 
OAI211_X1_1786_ (
  .A({ S2391 }),
  .B({ S2268 }),
  .C1({ S2397 }),
  .C2({ S25957[781] }),
  .ZN({ S2398 })
);
OAI211_X1 #() 
OAI211_X1_1787_ (
  .A({ S2398 }),
  .B({ S2305 }),
  .C1({ S2268 }),
  .C2({ S2383 }),
  .ZN({ S2399 })
);
NAND4_X1 #() 
NAND4_X1_593_ (
  .A1({ S2237 }),
  .A2({ S109 }),
  .A3({ S101 }),
  .A4({ S2243 }),
  .ZN({ S2400 })
);
NAND2_X1 #() 
NAND2_X1_5087_ (
  .A1({ S2269 }),
  .A2({ S101 }),
  .ZN({ S2401 })
);
NAND2_X1 #() 
NAND2_X1_5088_ (
  .A1({ S2400 }),
  .A2({ S2401 }),
  .ZN({ S2402 })
);
NAND2_X1 #() 
NAND2_X1_5089_ (
  .A1({ S2371 }),
  .A2({ S25957[780] }),
  .ZN({ S2403 })
);
NAND2_X1 #() 
NAND2_X1_5090_ (
  .A1({ S2249 }),
  .A2({ S25957[779] }),
  .ZN({ S2404 })
);
NAND3_X1 #() 
NAND3_X1_5460_ (
  .A1({ S2338 }),
  .A2({ S25957[779] }),
  .A3({ S25957[776] }),
  .ZN({ S2405 })
);
NAND3_X1 #() 
NAND3_X1_5461_ (
  .A1({ S2324 }),
  .A2({ S2404 }),
  .A3({ S2405 }),
  .ZN({ S2406 })
);
OAI21_X1 #() 
OAI21_X1_2641_ (
  .A({ S2406 }),
  .B1({ S2402 }),
  .B2({ S2403 }),
  .ZN({ S2407 })
);
NAND2_X1 #() 
NAND2_X1_5091_ (
  .A1({ S2244 }),
  .A2({ S25957[778] }),
  .ZN({ S2408 })
);
NAND2_X1 #() 
NAND2_X1_5092_ (
  .A1({ S2408 }),
  .A2({ S2281 }),
  .ZN({ S2409 })
);
NAND2_X1 #() 
NAND2_X1_5093_ (
  .A1({ S2409 }),
  .A2({ S25957[779] }),
  .ZN({ S2410 })
);
NAND3_X1 #() 
NAND3_X1_5462_ (
  .A1({ S2374 }),
  .A2({ S2248 }),
  .A3({ S101 }),
  .ZN({ S2411 })
);
AOI21_X1 #() 
AOI21_X1_2853_ (
  .A({ S2256 }),
  .B1({ S2410 }),
  .B2({ S2411 }),
  .ZN({ S2412 })
);
AOI21_X1 #() 
AOI21_X1_2854_ (
  .A({ S25957[780] }),
  .B1({ S2286 }),
  .B2({ S2270 }),
  .ZN({ S2413 })
);
OAI21_X1 #() 
OAI21_X1_2642_ (
  .A({ S25957[781] }),
  .B1({ S2412 }),
  .B2({ S2413 }),
  .ZN({ S2414 })
);
OAI21_X1 #() 
OAI21_X1_2643_ (
  .A({ S2414 }),
  .B1({ S2407 }),
  .B2({ S25957[781] }),
  .ZN({ S2415 })
);
NAND2_X1 #() 
NAND2_X1_5094_ (
  .A1({ S2273 }),
  .A2({ S25957[777] }),
  .ZN({ S2416 })
);
NAND2_X1 #() 
NAND2_X1_5095_ (
  .A1({ S2416 }),
  .A2({ S2338 }),
  .ZN({ S2417 })
);
NAND2_X1 #() 
NAND2_X1_5096_ (
  .A1({ S2417 }),
  .A2({ S25957[779] }),
  .ZN({ S2418 })
);
NAND3_X1 #() 
NAND3_X1_5463_ (
  .A1({ S2240 }),
  .A2({ S101 }),
  .A3({ S2281 }),
  .ZN({ S2419 })
);
AND2_X1 #() 
AND2_X1_313_ (
  .A1({ S2418 }),
  .A2({ S2419 }),
  .ZN({ S2420 })
);
OAI22_X1 #() 
OAI22_X1_129_ (
  .A1({ S2270 }),
  .A2({ S2273 }),
  .B1({ S2248 }),
  .B2({ S101 }),
  .ZN({ S2421 })
);
INV_X1 #() 
INV_X1_1664_ (
  .A({ S2421 }),
  .ZN({ S2422 })
);
NAND3_X1 #() 
NAND3_X1_5464_ (
  .A1({ S2422 }),
  .A2({ S25957[780] }),
  .A3({ S2345 }),
  .ZN({ S2423 })
);
OAI211_X1 #() 
OAI211_X1_1788_ (
  .A({ S25957[781] }),
  .B({ S2423 }),
  .C1({ S2420 }),
  .C2({ S25957[780] }),
  .ZN({ S2424 })
);
NAND2_X1 #() 
NAND2_X1_5097_ (
  .A1({ S25957[779] }),
  .A2({ S2258 }),
  .ZN({ S2425 })
);
NAND2_X1 #() 
NAND2_X1_5098_ (
  .A1({ S2269 }),
  .A2({ S25957[779] }),
  .ZN({ S2426 })
);
NAND2_X1 #() 
NAND2_X1_5099_ (
  .A1({ S2426 }),
  .A2({ S2425 }),
  .ZN({ S2427 })
);
NOR2_X1 #() 
NOR2_X1_1295_ (
  .A1({ S2312 }),
  .A2({ S25957[779] }),
  .ZN({ S2428 })
);
OAI21_X1 #() 
OAI21_X1_2644_ (
  .A({ S25957[780] }),
  .B1({ S2428 }),
  .B2({ S2427 }),
  .ZN({ S2429 })
);
OAI21_X1 #() 
OAI21_X1_2645_ (
  .A({ S2250 }),
  .B1({ S2248 }),
  .B2({ S25957[776] }),
  .ZN({ S2430 })
);
NAND2_X1 #() 
NAND2_X1_5100_ (
  .A1({ S2430 }),
  .A2({ S25957[779] }),
  .ZN({ S2431 })
);
NAND3_X1 #() 
NAND3_X1_5465_ (
  .A1({ S2431 }),
  .A2({ S2400 }),
  .A3({ S2401 }),
  .ZN({ S2432 })
);
OAI211_X1 #() 
OAI211_X1_1789_ (
  .A({ S2429 }),
  .B({ S2315 }),
  .C1({ S25957[780] }),
  .C2({ S2432 }),
  .ZN({ S2433 })
);
NAND3_X1 #() 
NAND3_X1_5466_ (
  .A1({ S2424 }),
  .A2({ S2268 }),
  .A3({ S2433 }),
  .ZN({ S2434 })
);
OAI211_X1 #() 
OAI211_X1_1790_ (
  .A({ S25957[783] }),
  .B({ S2434 }),
  .C1({ S2415 }),
  .C2({ S2268 }),
  .ZN({ S2435 })
);
NAND3_X1 #() 
NAND3_X1_5467_ (
  .A1({ S2399 }),
  .A2({ S2435 }),
  .A3({ S25957[886] }),
  .ZN({ S2436 })
);
NAND2_X1 #() 
NAND2_X1_5101_ (
  .A1({ S2399 }),
  .A2({ S2435 }),
  .ZN({ S2437 })
);
NAND2_X1 #() 
NAND2_X1_5102_ (
  .A1({ S2437 }),
  .A2({ S2365 }),
  .ZN({ S2438 })
);
NAND2_X1 #() 
NAND2_X1_5103_ (
  .A1({ S2438 }),
  .A2({ S2436 }),
  .ZN({ S2439 })
);
NAND2_X1 #() 
NAND2_X1_5104_ (
  .A1({ S2439 }),
  .A2({ S25957[950] }),
  .ZN({ S2440 })
);
INV_X1 #() 
INV_X1_1665_ (
  .A({ S2439 }),
  .ZN({ S25957[758] })
);
NAND2_X1 #() 
NAND2_X1_5105_ (
  .A1({ S25957[758] }),
  .A2({ S2363 }),
  .ZN({ S2441 })
);
NAND3_X1 #() 
NAND3_X1_5468_ (
  .A1({ S2441 }),
  .A2({ S25607 }),
  .A3({ S2440 }),
  .ZN({ S2442 })
);
NAND2_X1 #() 
NAND2_X1_5106_ (
  .A1({ S2441 }),
  .A2({ S2440 }),
  .ZN({ S25957[694] })
);
NAND2_X1 #() 
NAND2_X1_5107_ (
  .A1({ S25957[694] }),
  .A2({ S25957[790] }),
  .ZN({ S2443 })
);
NAND2_X1 #() 
NAND2_X1_5108_ (
  .A1({ S2443 }),
  .A2({ S2442 }),
  .ZN({ S2444 })
);
INV_X1 #() 
INV_X1_1666_ (
  .A({ S2444 }),
  .ZN({ S25957[662] })
);
NAND2_X1 #() 
NAND2_X1_5109_ (
  .A1({ S22919 }),
  .A2({ S22918 }),
  .ZN({ S2445 })
);
NAND2_X1 #() 
NAND2_X1_5110_ (
  .A1({ S2320 }),
  .A2({ S2273 }),
  .ZN({ S2446 })
);
NOR2_X1 #() 
NOR2_X1_1296_ (
  .A1({ S2446 }),
  .A2({ S2287 }),
  .ZN({ S2447 })
);
OAI21_X1 #() 
OAI21_X1_2646_ (
  .A({ S25957[780] }),
  .B1({ S2366 }),
  .B2({ S101 }),
  .ZN({ S2448 })
);
AOI21_X1 #() 
AOI21_X1_2855_ (
  .A({ S25957[779] }),
  .B1({ S2374 }),
  .B2({ S2258 }),
  .ZN({ S2449 })
);
NAND2_X1 #() 
NAND2_X1_5111_ (
  .A1({ S2245 }),
  .A2({ S25957[778] }),
  .ZN({ S2450 })
);
NAND2_X1 #() 
NAND2_X1_5112_ (
  .A1({ S2331 }),
  .A2({ S2450 }),
  .ZN({ S2451 })
);
AOI21_X1 #() 
AOI21_X1_2856_ (
  .A({ S2449 }),
  .B1({ S2451 }),
  .B2({ S25957[779] }),
  .ZN({ S2452 })
);
OAI221_X1 #() 
OAI221_X1_150_ (
  .A({ S25957[781] }),
  .B1({ S2447 }),
  .B2({ S2448 }),
  .C1({ S2452 }),
  .C2({ S25957[780] }),
  .ZN({ S2453 })
);
NAND3_X1 #() 
NAND3_X1_5469_ (
  .A1({ S2245 }),
  .A2({ S25957[779] }),
  .A3({ S2243 }),
  .ZN({ S2454 })
);
NAND2_X1 #() 
NAND2_X1_5113_ (
  .A1({ S2450 }),
  .A2({ S101 }),
  .ZN({ S2455 })
);
NAND3_X1 #() 
NAND3_X1_5470_ (
  .A1({ S2455 }),
  .A2({ S25957[780] }),
  .A3({ S2454 }),
  .ZN({ S2456 })
);
AND2_X1 #() 
AND2_X1_314_ (
  .A1({ S2371 }),
  .A2({ S2345 }),
  .ZN({ S2457 })
);
OAI211_X1 #() 
OAI211_X1_1791_ (
  .A({ S2315 }),
  .B({ S2456 }),
  .C1({ S2457 }),
  .C2({ S25957[780] }),
  .ZN({ S2458 })
);
NAND3_X1 #() 
NAND3_X1_5471_ (
  .A1({ S2453 }),
  .A2({ S25957[782] }),
  .A3({ S2458 }),
  .ZN({ S2459 })
);
NAND3_X1 #() 
NAND3_X1_5472_ (
  .A1({ S2237 }),
  .A2({ S101 }),
  .A3({ S2273 }),
  .ZN({ S2460 })
);
OAI211_X1 #() 
OAI211_X1_1792_ (
  .A({ S2460 }),
  .B({ S25957[780] }),
  .C1({ S2323 }),
  .C2({ S101 }),
  .ZN({ S2461 })
);
NAND3_X1 #() 
NAND3_X1_5473_ (
  .A1({ S2338 }),
  .A2({ S101 }),
  .A3({ S2245 }),
  .ZN({ S2462 })
);
NOR2_X1 #() 
NOR2_X1_1297_ (
  .A1({ S101 }),
  .A2({ S25957[777] }),
  .ZN({ S2463 })
);
NOR2_X1 #() 
NOR2_X1_1298_ (
  .A1({ S2463 }),
  .A2({ S25957[780] }),
  .ZN({ S2464 })
);
AOI21_X1 #() 
AOI21_X1_2857_ (
  .A({ S2315 }),
  .B1({ S2462 }),
  .B2({ S2464 }),
  .ZN({ S2465 })
);
INV_X1 #() 
INV_X1_1667_ (
  .A({ S2273 }),
  .ZN({ S2466 })
);
NAND2_X1 #() 
NAND2_X1_5114_ (
  .A1({ S2466 }),
  .A2({ S2258 }),
  .ZN({ S2467 })
);
AND2_X1 #() 
AND2_X1_315_ (
  .A1({ S2467 }),
  .A2({ S2240 }),
  .ZN({ S2468 })
);
OAI211_X1 #() 
OAI211_X1_1793_ (
  .A({ S2256 }),
  .B({ S2343 }),
  .C1({ S2468 }),
  .C2({ S101 }),
  .ZN({ S2469 })
);
INV_X1 #() 
INV_X1_1668_ (
  .A({ S109 }),
  .ZN({ S2470 })
);
NOR2_X1 #() 
NOR2_X1_1299_ (
  .A1({ S2331 }),
  .A2({ S2470 }),
  .ZN({ S2471 })
);
NAND2_X1 #() 
NAND2_X1_5115_ (
  .A1({ S2471 }),
  .A2({ S25957[779] }),
  .ZN({ S2472 })
);
NAND2_X1 #() 
NAND2_X1_5116_ (
  .A1({ S109 }),
  .A2({ S2285 }),
  .ZN({ S2473 })
);
NAND2_X1 #() 
NAND2_X1_5117_ (
  .A1({ S2473 }),
  .A2({ S101 }),
  .ZN({ S2474 })
);
NAND2_X1 #() 
NAND2_X1_5118_ (
  .A1({ S2472 }),
  .A2({ S2474 }),
  .ZN({ S2475 })
);
AOI21_X1 #() 
AOI21_X1_2858_ (
  .A({ S25957[781] }),
  .B1({ S2475 }),
  .B2({ S25957[780] }),
  .ZN({ S2476 })
);
AOI22_X1 #() 
AOI22_X1_577_ (
  .A1({ S2476 }),
  .A2({ S2469 }),
  .B1({ S2465 }),
  .B2({ S2461 }),
  .ZN({ S2477 })
);
OAI21_X1 #() 
OAI21_X1_2647_ (
  .A({ S2459 }),
  .B1({ S2477 }),
  .B2({ S25957[782] }),
  .ZN({ S2478 })
);
NAND2_X1 #() 
NAND2_X1_5119_ (
  .A1({ S2478 }),
  .A2({ S25957[783] }),
  .ZN({ S2479 })
);
NAND2_X1 #() 
NAND2_X1_5120_ (
  .A1({ S2446 }),
  .A2({ S25957[779] }),
  .ZN({ S2480 })
);
NAND2_X1 #() 
NAND2_X1_5121_ (
  .A1({ S2316 }),
  .A2({ S2257 }),
  .ZN({ S2481 })
);
NAND2_X1 #() 
NAND2_X1_5122_ (
  .A1({ S2481 }),
  .A2({ S101 }),
  .ZN({ S2482 })
);
NAND3_X1 #() 
NAND3_X1_5474_ (
  .A1({ S2482 }),
  .A2({ S25957[780] }),
  .A3({ S2480 }),
  .ZN({ S2483 })
);
NAND4_X1 #() 
NAND4_X1_594_ (
  .A1({ S2250 }),
  .A2({ S2285 }),
  .A3({ S2262 }),
  .A4({ S25957[779] }),
  .ZN({ S2484 })
);
NAND2_X1 #() 
NAND2_X1_5123_ (
  .A1({ S2484 }),
  .A2({ S2269 }),
  .ZN({ S2485 })
);
INV_X1 #() 
INV_X1_1669_ (
  .A({ S2485 }),
  .ZN({ S2486 })
);
NOR2_X1 #() 
NOR2_X1_1300_ (
  .A1({ S2245 }),
  .A2({ S25957[778] }),
  .ZN({ S2487 })
);
NAND2_X1 #() 
NAND2_X1_5124_ (
  .A1({ S2256 }),
  .A2({ S101 }),
  .ZN({ S2488 })
);
OAI22_X1 #() 
OAI22_X1_130_ (
  .A1({ S2484 }),
  .A2({ S25957[780] }),
  .B1({ S2488 }),
  .B2({ S2487 }),
  .ZN({ S2489 })
);
INV_X1 #() 
INV_X1_1670_ (
  .A({ S2489 }),
  .ZN({ S2490 })
);
OAI21_X1 #() 
OAI21_X1_2648_ (
  .A({ S2483 }),
  .B1({ S2486 }),
  .B2({ S2490 }),
  .ZN({ S2491 })
);
NAND4_X1 #() 
NAND4_X1_595_ (
  .A1({ S788 }),
  .A2({ S791 }),
  .A3({ S866 }),
  .A4({ S869 }),
  .ZN({ S2492 })
);
NAND3_X1 #() 
NAND3_X1_5475_ (
  .A1({ S2250 }),
  .A2({ S101 }),
  .A3({ S2245 }),
  .ZN({ S2493 })
);
AND2_X1 #() 
AND2_X1_316_ (
  .A1({ S2493 }),
  .A2({ S2492 }),
  .ZN({ S2494 })
);
NAND3_X1 #() 
NAND3_X1_5476_ (
  .A1({ S2282 }),
  .A2({ S25957[777] }),
  .A3({ S2243 }),
  .ZN({ S2495 })
);
NAND3_X1 #() 
NAND3_X1_5477_ (
  .A1({ S2326 }),
  .A2({ S25957[779] }),
  .A3({ S2495 }),
  .ZN({ S2496 })
);
OAI211_X1 #() 
OAI211_X1_1794_ (
  .A({ S2496 }),
  .B({ S25957[780] }),
  .C1({ S25957[779] }),
  .C2({ S2313 }),
  .ZN({ S2497 })
);
OAI211_X1 #() 
OAI211_X1_1795_ (
  .A({ S2497 }),
  .B({ S25957[781] }),
  .C1({ S25957[780] }),
  .C2({ S2494 }),
  .ZN({ S2498 })
);
OAI211_X1 #() 
OAI211_X1_1796_ (
  .A({ S2498 }),
  .B({ S25957[782] }),
  .C1({ S2491 }),
  .C2({ S25957[781] }),
  .ZN({ S2499 })
);
NOR2_X1 #() 
NOR2_X1_1301_ (
  .A1({ S2248 }),
  .A2({ S25957[779] }),
  .ZN({ S2500 })
);
OAI211_X1 #() 
OAI211_X1_1797_ (
  .A({ S2256 }),
  .B({ S25957[776] }),
  .C1({ S2500 }),
  .C2({ S2463 }),
  .ZN({ S2501 })
);
AOI21_X1 #() 
AOI21_X1_2859_ (
  .A({ S101 }),
  .B1({ S2240 }),
  .B2({ S2312 }),
  .ZN({ S2502 })
);
AOI21_X1 #() 
AOI21_X1_2860_ (
  .A({ S25957[779] }),
  .B1({ S2283 }),
  .B2({ S2237 }),
  .ZN({ S2503 })
);
OR2_X1 #() 
OR2_X1_70_ (
  .A1({ S2503 }),
  .A2({ S2256 }),
  .ZN({ S2504 })
);
OAI21_X1 #() 
OAI21_X1_2649_ (
  .A({ S2501 }),
  .B1({ S2504 }),
  .B2({ S2502 }),
  .ZN({ S2505 })
);
NAND4_X1 #() 
NAND4_X1_596_ (
  .A1({ S788 }),
  .A2({ S2241 }),
  .A3({ S2242 }),
  .A4({ S791 }),
  .ZN({ S2506 })
);
INV_X1 #() 
INV_X1_1671_ (
  .A({ S2506 }),
  .ZN({ S2507 })
);
OAI211_X1 #() 
OAI211_X1_1798_ (
  .A({ S2256 }),
  .B({ S2262 }),
  .C1({ S2377 }),
  .C2({ S2507 }),
  .ZN({ S2508 })
);
NAND2_X1 #() 
NAND2_X1_5125_ (
  .A1({ S2487 }),
  .A2({ S101 }),
  .ZN({ S2509 })
);
NAND4_X1 #() 
NAND4_X1_597_ (
  .A1({ S2276 }),
  .A2({ S2509 }),
  .A3({ S25957[780] }),
  .A4({ S2506 }),
  .ZN({ S2510 })
);
AOI21_X1 #() 
AOI21_X1_2861_ (
  .A({ S2315 }),
  .B1({ S2508 }),
  .B2({ S2510 }),
  .ZN({ S2511 })
);
AOI21_X1 #() 
AOI21_X1_2862_ (
  .A({ S2511 }),
  .B1({ S2505 }),
  .B2({ S2315 }),
  .ZN({ S2512 })
);
OAI21_X1 #() 
OAI21_X1_2650_ (
  .A({ S2499 }),
  .B1({ S2512 }),
  .B2({ S25957[782] }),
  .ZN({ S2513 })
);
NAND2_X1 #() 
NAND2_X1_5126_ (
  .A1({ S2513 }),
  .A2({ S2305 }),
  .ZN({ S2514 })
);
NAND2_X1 #() 
NAND2_X1_5127_ (
  .A1({ S2479 }),
  .A2({ S2514 }),
  .ZN({ S2515 })
);
NAND2_X1 #() 
NAND2_X1_5128_ (
  .A1({ S2515 }),
  .A2({ S25957[885] }),
  .ZN({ S2516 })
);
NAND3_X1 #() 
NAND3_X1_5478_ (
  .A1({ S2479 }),
  .A2({ S2514 }),
  .A3({ S25666 }),
  .ZN({ S2517 })
);
AOI21_X1 #() 
AOI21_X1_2863_ (
  .A({ S2445 }),
  .B1({ S2516 }),
  .B2({ S2517 }),
  .ZN({ S2518 })
);
NAND3_X1 #() 
NAND3_X1_5479_ (
  .A1({ S2516 }),
  .A2({ S2445 }),
  .A3({ S2517 }),
  .ZN({ S2519 })
);
INV_X1 #() 
INV_X1_1672_ (
  .A({ S2519 }),
  .ZN({ S2520 })
);
OAI21_X1 #() 
OAI21_X1_2651_ (
  .A({ S25673 }),
  .B1({ S2520 }),
  .B2({ S2518 }),
  .ZN({ S2521 })
);
INV_X1 #() 
INV_X1_1673_ (
  .A({ S2518 }),
  .ZN({ S2522 })
);
NAND3_X1 #() 
NAND3_X1_5480_ (
  .A1({ S2522 }),
  .A2({ S25957[789] }),
  .A3({ S2519 }),
  .ZN({ S2523 })
);
AND2_X1 #() 
AND2_X1_317_ (
  .A1({ S2521 }),
  .A2({ S2523 }),
  .ZN({ S25957[661] })
);
NOR2_X1 #() 
NOR2_X1_1302_ (
  .A1({ S25741 }),
  .A2({ S25745 }),
  .ZN({ S25957[852] })
);
XNOR2_X1 #() 
XNOR2_X1_198_ (
  .A({ S25957[852] }),
  .B({ S25676 }),
  .ZN({ S25957[820] })
);
NAND2_X1 #() 
NAND2_X1_5129_ (
  .A1({ S25746 }),
  .A2({ S25749 }),
  .ZN({ S2524 })
);
NAND2_X1 #() 
NAND2_X1_5130_ (
  .A1({ S25744 }),
  .A2({ S25743 }),
  .ZN({ S25957[884] })
);
INV_X1 #() 
INV_X1_1674_ (
  .A({ S25957[884] }),
  .ZN({ S2525 })
);
NAND3_X1 #() 
NAND3_X1_5481_ (
  .A1({ S2320 }),
  .A2({ S101 }),
  .A3({ S2282 }),
  .ZN({ S2526 })
);
AND2_X1 #() 
AND2_X1_318_ (
  .A1({ S2339 }),
  .A2({ S2526 }),
  .ZN({ S2527 })
);
OAI21_X1 #() 
OAI21_X1_2652_ (
  .A({ S101 }),
  .B1({ S2262 }),
  .B2({ S25957[777] }),
  .ZN({ S2528 })
);
NAND2_X1 #() 
NAND2_X1_5131_ (
  .A1({ S2480 }),
  .A2({ S2528 }),
  .ZN({ S2529 })
);
NAND2_X1 #() 
NAND2_X1_5132_ (
  .A1({ S2529 }),
  .A2({ S25957[780] }),
  .ZN({ S2530 })
);
OAI211_X1 #() 
OAI211_X1_1799_ (
  .A({ S2530 }),
  .B({ S25957[781] }),
  .C1({ S2527 }),
  .C2({ S25957[780] }),
  .ZN({ S2531 })
);
OAI21_X1 #() 
OAI21_X1_2653_ (
  .A({ S2462 }),
  .B1({ S2376 }),
  .B2({ S2425 }),
  .ZN({ S2532 })
);
NAND2_X1 #() 
NAND2_X1_5133_ (
  .A1({ S2532 }),
  .A2({ S25957[780] }),
  .ZN({ S2533 })
);
INV_X1 #() 
INV_X1_1675_ (
  .A({ S2335 }),
  .ZN({ S2534 })
);
NAND3_X1 #() 
NAND3_X1_5482_ (
  .A1({ S2338 }),
  .A2({ S101 }),
  .A3({ S2262 }),
  .ZN({ S2535 })
);
INV_X1 #() 
INV_X1_1676_ (
  .A({ S2535 }),
  .ZN({ S2536 })
);
OAI21_X1 #() 
OAI21_X1_2654_ (
  .A({ S2256 }),
  .B1({ S2534 }),
  .B2({ S2536 }),
  .ZN({ S2537 })
);
NAND3_X1 #() 
NAND3_X1_5483_ (
  .A1({ S2537 }),
  .A2({ S2533 }),
  .A3({ S2315 }),
  .ZN({ S2538 })
);
AND2_X1 #() 
AND2_X1_319_ (
  .A1({ S2538 }),
  .A2({ S2531 }),
  .ZN({ S2539 })
);
OAI221_X1 #() 
OAI221_X1_151_ (
  .A({ S2256 }),
  .B1({ S2425 }),
  .B2({ S2269 }),
  .C1({ S2455 }),
  .C2({ S2487 }),
  .ZN({ S2540 })
);
AOI21_X1 #() 
AOI21_X1_2864_ (
  .A({ S25957[779] }),
  .B1({ S2331 }),
  .B2({ S2450 }),
  .ZN({ S2541 })
);
INV_X1 #() 
INV_X1_1677_ (
  .A({ S2541 }),
  .ZN({ S2542 })
);
AOI21_X1 #() 
AOI21_X1_2865_ (
  .A({ S2256 }),
  .B1({ S2385 }),
  .B2({ S2321 }),
  .ZN({ S2543 })
);
NAND2_X1 #() 
NAND2_X1_5134_ (
  .A1({ S2543 }),
  .A2({ S2542 }),
  .ZN({ S2544 })
);
NAND2_X1 #() 
NAND2_X1_5135_ (
  .A1({ S2544 }),
  .A2({ S2540 }),
  .ZN({ S2545 })
);
NAND4_X1 #() 
NAND4_X1_598_ (
  .A1({ S2257 }),
  .A2({ S2262 }),
  .A3({ S109 }),
  .A4({ S2285 }),
  .ZN({ S2546 })
);
NAND3_X1 #() 
NAND3_X1_5484_ (
  .A1({ S2291 }),
  .A2({ S2312 }),
  .A3({ S2290 }),
  .ZN({ S2547 })
);
OAI21_X1 #() 
OAI21_X1_2655_ (
  .A({ S2547 }),
  .B1({ S2546 }),
  .B2({ S2488 }),
  .ZN({ S2548 })
);
AOI21_X1 #() 
AOI21_X1_2866_ (
  .A({ S25957[779] }),
  .B1({ S2408 }),
  .B2({ S2395 }),
  .ZN({ S2549 })
);
NAND2_X1 #() 
NAND2_X1_5136_ (
  .A1({ S2244 }),
  .A2({ S25957[779] }),
  .ZN({ S2550 })
);
OAI21_X1 #() 
OAI21_X1_2656_ (
  .A({ S25957[780] }),
  .B1({ S2550 }),
  .B2({ S2487 }),
  .ZN({ S2551 })
);
OAI21_X1 #() 
OAI21_X1_2657_ (
  .A({ S25957[781] }),
  .B1({ S2551 }),
  .B2({ S2549 }),
  .ZN({ S2552 })
);
OAI221_X1 #() 
OAI221_X1_152_ (
  .A({ S2268 }),
  .B1({ S2548 }),
  .B2({ S2552 }),
  .C1({ S2545 }),
  .C2({ S25957[781] }),
  .ZN({ S2553 })
);
OAI211_X1 #() 
OAI211_X1_1800_ (
  .A({ S2553 }),
  .B({ S25957[783] }),
  .C1({ S2268 }),
  .C2({ S2539 }),
  .ZN({ S2554 })
);
NOR2_X1 #() 
NOR2_X1_1303_ (
  .A1({ S2507 }),
  .A2({ S25957[780] }),
  .ZN({ S2555 })
);
OAI21_X1 #() 
OAI21_X1_2658_ (
  .A({ S2555 }),
  .B1({ S2307 }),
  .B2({ S2263 }),
  .ZN({ S2556 })
);
OAI211_X1 #() 
OAI211_X1_1801_ (
  .A({ S2271 }),
  .B({ S25957[780] }),
  .C1({ S2411 }),
  .C2({ S2264 }),
  .ZN({ S2557 })
);
NAND3_X1 #() 
NAND3_X1_5485_ (
  .A1({ S2556 }),
  .A2({ S2557 }),
  .A3({ S2315 }),
  .ZN({ S2558 })
);
AOI21_X1 #() 
AOI21_X1_2867_ (
  .A({ S2243 }),
  .B1({ S2282 }),
  .B2({ S25957[777] }),
  .ZN({ S2559 })
);
OAI21_X1 #() 
OAI21_X1_2659_ (
  .A({ S101 }),
  .B1({ S2471 }),
  .B2({ S2559 }),
  .ZN({ S2560 })
);
NAND2_X1 #() 
NAND2_X1_5137_ (
  .A1({ S2484 }),
  .A2({ S2256 }),
  .ZN({ S2561 })
);
INV_X1 #() 
INV_X1_1678_ (
  .A({ S2561 }),
  .ZN({ S2562 })
);
NAND2_X1 #() 
NAND2_X1_5138_ (
  .A1({ S2560 }),
  .A2({ S2562 }),
  .ZN({ S2563 })
);
INV_X1 #() 
INV_X1_1679_ (
  .A({ S132 }),
  .ZN({ S2564 })
);
OAI21_X1 #() 
OAI21_X1_2660_ (
  .A({ S25957[780] }),
  .B1({ S2564 }),
  .B2({ S25957[778] }),
  .ZN({ S2565 })
);
NAND3_X1 #() 
NAND3_X1_5486_ (
  .A1({ S2563 }),
  .A2({ S25957[781] }),
  .A3({ S2565 }),
  .ZN({ S2566 })
);
NAND2_X1 #() 
NAND2_X1_5139_ (
  .A1({ S2566 }),
  .A2({ S2558 }),
  .ZN({ S2567 })
);
NAND3_X1 #() 
NAND3_X1_5487_ (
  .A1({ S2392 }),
  .A2({ S25957[780] }),
  .A3({ S2455 }),
  .ZN({ S2568 })
);
OAI21_X1 #() 
OAI21_X1_2661_ (
  .A({ S2472 }),
  .B1({ S2258 }),
  .B2({ S2337 }),
  .ZN({ S2569 })
);
OAI21_X1 #() 
OAI21_X1_2662_ (
  .A({ S2568 }),
  .B1({ S2569 }),
  .B2({ S25957[780] }),
  .ZN({ S2570 })
);
NAND3_X1 #() 
NAND3_X1_5488_ (
  .A1({ S2374 }),
  .A2({ S109 }),
  .A3({ S25957[779] }),
  .ZN({ S2571 })
);
NAND3_X1 #() 
NAND3_X1_5489_ (
  .A1({ S2281 }),
  .A2({ S2283 }),
  .A3({ S101 }),
  .ZN({ S2572 })
);
AOI21_X1 #() 
AOI21_X1_2868_ (
  .A({ S25957[780] }),
  .B1({ S2572 }),
  .B2({ S2571 }),
  .ZN({ S2573 })
);
NAND4_X1 #() 
NAND4_X1_599_ (
  .A1({ S2374 }),
  .A2({ S2320 }),
  .A3({ S2273 }),
  .A4({ S25957[779] }),
  .ZN({ S2574 })
);
AND3_X1 #() 
AND3_X1_214_ (
  .A1({ S2574 }),
  .A2({ S2462 }),
  .A3({ S25957[780] }),
  .ZN({ S2575 })
);
OAI21_X1 #() 
OAI21_X1_2663_ (
  .A({ S2315 }),
  .B1({ S2573 }),
  .B2({ S2575 }),
  .ZN({ S2576 })
);
OAI211_X1 #() 
OAI211_X1_1802_ (
  .A({ S2268 }),
  .B({ S2576 }),
  .C1({ S2570 }),
  .C2({ S2315 }),
  .ZN({ S2577 })
);
OAI211_X1 #() 
OAI211_X1_1803_ (
  .A({ S2577 }),
  .B({ S2305 }),
  .C1({ S2268 }),
  .C2({ S2567 }),
  .ZN({ S2578 })
);
NAND3_X1 #() 
NAND3_X1_5490_ (
  .A1({ S2578 }),
  .A2({ S2554 }),
  .A3({ S2525 }),
  .ZN({ S2579 })
);
NAND2_X1 #() 
NAND2_X1_5140_ (
  .A1({ S2567 }),
  .A2({ S25957[782] }),
  .ZN({ S2580 })
);
NAND2_X1 #() 
NAND2_X1_5141_ (
  .A1({ S2570 }),
  .A2({ S25957[781] }),
  .ZN({ S2581 })
);
OR3_X1 #() 
OR3_X1_33_ (
  .A1({ S2573 }),
  .A2({ S2575 }),
  .A3({ S25957[781] }),
  .ZN({ S2582 })
);
NAND3_X1 #() 
NAND3_X1_5491_ (
  .A1({ S2581 }),
  .A2({ S2582 }),
  .A3({ S2268 }),
  .ZN({ S2583 })
);
NAND3_X1 #() 
NAND3_X1_5492_ (
  .A1({ S2583 }),
  .A2({ S2580 }),
  .A3({ S2305 }),
  .ZN({ S2584 })
);
INV_X1 #() 
INV_X1_1680_ (
  .A({ S2545 }),
  .ZN({ S2585 })
);
NOR2_X1 #() 
NOR2_X1_1304_ (
  .A1({ S2552 }),
  .A2({ S2548 }),
  .ZN({ S2586 })
);
AOI21_X1 #() 
AOI21_X1_2869_ (
  .A({ S2586 }),
  .B1({ S2585 }),
  .B2({ S2315 }),
  .ZN({ S2587 })
);
NAND3_X1 #() 
NAND3_X1_5493_ (
  .A1({ S2538 }),
  .A2({ S2531 }),
  .A3({ S25957[782] }),
  .ZN({ S2588 })
);
OAI211_X1 #() 
OAI211_X1_1804_ (
  .A({ S25957[783] }),
  .B({ S2588 }),
  .C1({ S2587 }),
  .C2({ S25957[782] }),
  .ZN({ S2589 })
);
NAND3_X1 #() 
NAND3_X1_5494_ (
  .A1({ S2584 }),
  .A2({ S2589 }),
  .A3({ S25957[884] }),
  .ZN({ S2590 })
);
AOI21_X1 #() 
AOI21_X1_2870_ (
  .A({ S25957[948] }),
  .B1({ S2590 }),
  .B2({ S2579 }),
  .ZN({ S2591 })
);
NAND3_X1 #() 
NAND3_X1_5495_ (
  .A1({ S2578 }),
  .A2({ S2554 }),
  .A3({ S25957[884] }),
  .ZN({ S2592 })
);
NAND3_X1 #() 
NAND3_X1_5496_ (
  .A1({ S2584 }),
  .A2({ S2589 }),
  .A3({ S2525 }),
  .ZN({ S2593 })
);
AOI21_X1 #() 
AOI21_X1_2871_ (
  .A({ S25676 }),
  .B1({ S2593 }),
  .B2({ S2592 }),
  .ZN({ S2594 })
);
OAI21_X1 #() 
OAI21_X1_2664_ (
  .A({ S2524 }),
  .B1({ S2591 }),
  .B2({ S2594 }),
  .ZN({ S2595 })
);
NAND3_X1 #() 
NAND3_X1_5497_ (
  .A1({ S2593 }),
  .A2({ S2592 }),
  .A3({ S25676 }),
  .ZN({ S2596 })
);
NAND3_X1 #() 
NAND3_X1_5498_ (
  .A1({ S2590 }),
  .A2({ S2579 }),
  .A3({ S25957[948] }),
  .ZN({ S2597 })
);
NAND3_X1 #() 
NAND3_X1_5499_ (
  .A1({ S2596 }),
  .A2({ S2597 }),
  .A3({ S25957[788] }),
  .ZN({ S2598 })
);
NAND2_X1 #() 
NAND2_X1_5142_ (
  .A1({ S2595 }),
  .A2({ S2598 }),
  .ZN({ S25957[660] })
);
NOR2_X1 #() 
NOR2_X1_1305_ (
  .A1({ S25827 }),
  .A2({ S25826 }),
  .ZN({ S25957[819] })
);
NOR2_X1 #() 
NOR2_X1_1306_ (
  .A1({ S23076 }),
  .A2({ S23075 }),
  .ZN({ S25957[979] })
);
INV_X1 #() 
INV_X1_1681_ (
  .A({ S25957[979] }),
  .ZN({ S2599 })
);
NAND3_X1 #() 
NAND3_X1_5500_ (
  .A1({ S2244 }),
  .A2({ S2320 }),
  .A3({ S101 }),
  .ZN({ S2600 })
);
OAI211_X1 #() 
OAI211_X1_1805_ (
  .A({ S2600 }),
  .B({ S2256 }),
  .C1({ S2249 }),
  .C2({ S2492 }),
  .ZN({ S2601 })
);
OAI211_X1 #() 
OAI211_X1_1806_ (
  .A({ S25957[781] }),
  .B({ S2601 }),
  .C1({ S2403 }),
  .C2({ S2344 }),
  .ZN({ S2602 })
);
NAND4_X1 #() 
NAND4_X1_600_ (
  .A1({ S2285 }),
  .A2({ S2320 }),
  .A3({ S101 }),
  .A4({ S25957[776] }),
  .ZN({ S2603 })
);
OAI211_X1 #() 
OAI211_X1_1807_ (
  .A({ S2603 }),
  .B({ S2256 }),
  .C1({ S2297 }),
  .C2({ S2299 }),
  .ZN({ S2604 })
);
NAND3_X1 #() 
NAND3_X1_5501_ (
  .A1({ S2237 }),
  .A2({ S2374 }),
  .A3({ S101 }),
  .ZN({ S2605 })
);
INV_X1 #() 
INV_X1_1682_ (
  .A({ S2605 }),
  .ZN({ S2606 })
);
OAI211_X1 #() 
OAI211_X1_1808_ (
  .A({ S2604 }),
  .B({ S2315 }),
  .C1({ S2256 }),
  .C2({ S2606 }),
  .ZN({ S2607 })
);
NAND2_X1 #() 
NAND2_X1_5143_ (
  .A1({ S2602 }),
  .A2({ S2607 }),
  .ZN({ S2608 })
);
NAND2_X1 #() 
NAND2_X1_5144_ (
  .A1({ S2608 }),
  .A2({ S25957[782] }),
  .ZN({ S2609 })
);
INV_X1 #() 
INV_X1_1683_ (
  .A({ S2326 }),
  .ZN({ S2610 })
);
OAI211_X1 #() 
OAI211_X1_1809_ (
  .A({ S25957[780] }),
  .B({ S2308 }),
  .C1({ S2610 }),
  .C2({ S25957[779] }),
  .ZN({ S2611 })
);
OAI221_X1 #() 
OAI221_X1_153_ (
  .A({ S2256 }),
  .B1({ S2280 }),
  .B2({ S2269 }),
  .C1({ S2384 }),
  .C2({ S101 }),
  .ZN({ S2612 })
);
AND3_X1 #() 
AND3_X1_215_ (
  .A1({ S2611 }),
  .A2({ S25957[781] }),
  .A3({ S2612 }),
  .ZN({ S2613 })
);
NAND4_X1 #() 
NAND4_X1_601_ (
  .A1({ S2374 }),
  .A2({ S2244 }),
  .A3({ S2245 }),
  .A4({ S25957[779] }),
  .ZN({ S2614 })
);
NAND3_X1 #() 
NAND3_X1_5502_ (
  .A1({ S2387 }),
  .A2({ S2614 }),
  .A3({ S25957[780] }),
  .ZN({ S2615 })
);
AOI21_X1 #() 
AOI21_X1_2872_ (
  .A({ S101 }),
  .B1({ S2331 }),
  .B2({ S2374 }),
  .ZN({ S2616 })
);
OAI21_X1 #() 
OAI21_X1_2665_ (
  .A({ S2256 }),
  .B1({ S2327 }),
  .B2({ S2616 }),
  .ZN({ S2617 })
);
AOI21_X1 #() 
AOI21_X1_2873_ (
  .A({ S25957[781] }),
  .B1({ S2617 }),
  .B2({ S2615 }),
  .ZN({ S2618 })
);
OAI21_X1 #() 
OAI21_X1_2666_ (
  .A({ S2268 }),
  .B1({ S2618 }),
  .B2({ S2613 }),
  .ZN({ S2619 })
);
NAND3_X1 #() 
NAND3_X1_5503_ (
  .A1({ S2619 }),
  .A2({ S2609 }),
  .A3({ S2305 }),
  .ZN({ S2620 })
);
NAND2_X1 #() 
NAND2_X1_5145_ (
  .A1({ S2416 }),
  .A2({ S25957[779] }),
  .ZN({ S2621 })
);
NAND3_X1 #() 
NAND3_X1_5504_ (
  .A1({ S2326 }),
  .A2({ S101 }),
  .A3({ S2296 }),
  .ZN({ S2622 })
);
AND2_X1 #() 
AND2_X1_320_ (
  .A1({ S2622 }),
  .A2({ S2621 }),
  .ZN({ S2623 })
);
NAND2_X1 #() 
NAND2_X1_5146_ (
  .A1({ S2374 }),
  .A2({ S2245 }),
  .ZN({ S2624 })
);
NAND2_X1 #() 
NAND2_X1_5147_ (
  .A1({ S2555 }),
  .A2({ S2624 }),
  .ZN({ S2625 })
);
OAI211_X1 #() 
OAI211_X1_1810_ (
  .A({ S2315 }),
  .B({ S2625 }),
  .C1({ S2623 }),
  .C2({ S2256 }),
  .ZN({ S2626 })
);
NAND2_X1 #() 
NAND2_X1_5148_ (
  .A1({ S2338 }),
  .A2({ S25957[779] }),
  .ZN({ S2627 })
);
NOR2_X1 #() 
NOR2_X1_1307_ (
  .A1({ S2370 }),
  .A2({ S2627 }),
  .ZN({ S2628 })
);
NAND2_X1 #() 
NAND2_X1_5149_ (
  .A1({ S2269 }),
  .A2({ S25957[777] }),
  .ZN({ S2629 })
);
AOI21_X1 #() 
AOI21_X1_2874_ (
  .A({ S25957[779] }),
  .B1({ S2246 }),
  .B2({ S2629 }),
  .ZN({ S2630 })
);
OAI21_X1 #() 
OAI21_X1_2667_ (
  .A({ S2256 }),
  .B1({ S2630 }),
  .B2({ S2628 }),
  .ZN({ S2631 })
);
NAND3_X1 #() 
NAND3_X1_5505_ (
  .A1({ S2290 }),
  .A2({ S101 }),
  .A3({ S2244 }),
  .ZN({ S2632 })
);
NAND3_X1 #() 
NAND3_X1_5506_ (
  .A1({ S2632 }),
  .A2({ S25957[780] }),
  .A3({ S2571 }),
  .ZN({ S2633 })
);
NAND3_X1 #() 
NAND3_X1_5507_ (
  .A1({ S2631 }),
  .A2({ S25957[781] }),
  .A3({ S2633 }),
  .ZN({ S2634 })
);
NAND3_X1 #() 
NAND3_X1_5508_ (
  .A1({ S2626 }),
  .A2({ S2634 }),
  .A3({ S25957[782] }),
  .ZN({ S2635 })
);
AOI21_X1 #() 
AOI21_X1_2875_ (
  .A({ S2256 }),
  .B1({ S2370 }),
  .B2({ S101 }),
  .ZN({ S2636 })
);
OAI21_X1 #() 
OAI21_X1_2668_ (
  .A({ S2636 }),
  .B1({ S2471 }),
  .B2({ S2308 }),
  .ZN({ S2637 })
);
NAND4_X1 #() 
NAND4_X1_602_ (
  .A1({ S2250 }),
  .A2({ S2262 }),
  .A3({ S25957[779] }),
  .A4({ S25957[777] }),
  .ZN({ S2638 })
);
NAND3_X1 #() 
NAND3_X1_5509_ (
  .A1({ S2240 }),
  .A2({ S101 }),
  .A3({ S2338 }),
  .ZN({ S2639 })
);
NAND3_X1 #() 
NAND3_X1_5510_ (
  .A1({ S2639 }),
  .A2({ S2256 }),
  .A3({ S2638 }),
  .ZN({ S2640 })
);
NAND3_X1 #() 
NAND3_X1_5511_ (
  .A1({ S2637 }),
  .A2({ S25957[781] }),
  .A3({ S2640 }),
  .ZN({ S2641 })
);
OAI221_X1 #() 
OAI221_X1_154_ (
  .A({ S2256 }),
  .B1({ S25957[779] }),
  .B2({ S2624 }),
  .C1({ S2610 }),
  .C2({ S2627 }),
  .ZN({ S2642 })
);
AOI21_X1 #() 
AOI21_X1_2876_ (
  .A({ S25957[778] }),
  .B1({ S2237 }),
  .B2({ S109 }),
  .ZN({ S2643 })
);
OAI211_X1 #() 
OAI211_X1_1811_ (
  .A({ S25957[780] }),
  .B({ S2535 }),
  .C1({ S2643 }),
  .C2({ S101 }),
  .ZN({ S2644 })
);
NAND3_X1 #() 
NAND3_X1_5512_ (
  .A1({ S2642 }),
  .A2({ S2315 }),
  .A3({ S2644 }),
  .ZN({ S2645 })
);
NAND3_X1 #() 
NAND3_X1_5513_ (
  .A1({ S2645 }),
  .A2({ S2641 }),
  .A3({ S2268 }),
  .ZN({ S2646 })
);
NAND3_X1 #() 
NAND3_X1_5514_ (
  .A1({ S2635 }),
  .A2({ S25957[783] }),
  .A3({ S2646 }),
  .ZN({ S2647 })
);
NAND3_X1 #() 
NAND3_X1_5515_ (
  .A1({ S2620 }),
  .A2({ S2647 }),
  .A3({ S2599 }),
  .ZN({ S2648 })
);
NAND2_X1 #() 
NAND2_X1_5150_ (
  .A1({ S2635 }),
  .A2({ S2646 }),
  .ZN({ S2649 })
);
NAND2_X1 #() 
NAND2_X1_5151_ (
  .A1({ S2649 }),
  .A2({ S25957[783] }),
  .ZN({ S2650 })
);
AND2_X1 #() 
AND2_X1_321_ (
  .A1({ S2617 }),
  .A2({ S2615 }),
  .ZN({ S2651 })
);
NAND3_X1 #() 
NAND3_X1_5516_ (
  .A1({ S2611 }),
  .A2({ S25957[781] }),
  .A3({ S2612 }),
  .ZN({ S2652 })
);
OAI211_X1 #() 
OAI211_X1_1812_ (
  .A({ S2268 }),
  .B({ S2652 }),
  .C1({ S2651 }),
  .C2({ S25957[781] }),
  .ZN({ S2653 })
);
NAND3_X1 #() 
NAND3_X1_5517_ (
  .A1({ S2602 }),
  .A2({ S2607 }),
  .A3({ S25957[782] }),
  .ZN({ S2654 })
);
NAND3_X1 #() 
NAND3_X1_5518_ (
  .A1({ S2653 }),
  .A2({ S2305 }),
  .A3({ S2654 }),
  .ZN({ S2655 })
);
NAND3_X1 #() 
NAND3_X1_5519_ (
  .A1({ S2650 }),
  .A2({ S2655 }),
  .A3({ S25957[979] }),
  .ZN({ S2656 })
);
NAND3_X1 #() 
NAND3_X1_5520_ (
  .A1({ S2656 }),
  .A2({ S25957[819] }),
  .A3({ S2648 }),
  .ZN({ S2657 })
);
INV_X1 #() 
INV_X1_1684_ (
  .A({ S25957[819] }),
  .ZN({ S2658 })
);
AND3_X1 #() 
AND3_X1_216_ (
  .A1({ S2620 }),
  .A2({ S2599 }),
  .A3({ S2647 }),
  .ZN({ S2659 })
);
AOI21_X1 #() 
AOI21_X1_2877_ (
  .A({ S2599 }),
  .B1({ S2620 }),
  .B2({ S2647 }),
  .ZN({ S2660 })
);
OAI21_X1 #() 
OAI21_X1_2669_ (
  .A({ S2658 }),
  .B1({ S2659 }),
  .B2({ S2660 }),
  .ZN({ S2661 })
);
NAND3_X1 #() 
NAND3_X1_5521_ (
  .A1({ S2661 }),
  .A2({ S25957[787] }),
  .A3({ S2657 }),
  .ZN({ S2662 })
);
OAI21_X1 #() 
OAI21_X1_2670_ (
  .A({ S25957[819] }),
  .B1({ S2659 }),
  .B2({ S2660 }),
  .ZN({ S2663 })
);
NAND3_X1 #() 
NAND3_X1_5522_ (
  .A1({ S2656 }),
  .A2({ S2658 }),
  .A3({ S2648 }),
  .ZN({ S2664 })
);
NAND3_X1 #() 
NAND3_X1_5523_ (
  .A1({ S2663 }),
  .A2({ S98 }),
  .A3({ S2664 }),
  .ZN({ S2665 })
);
NAND2_X1 #() 
NAND2_X1_5152_ (
  .A1({ S2662 }),
  .A2({ S2665 }),
  .ZN({ S110 })
);
AND2_X1 #() 
AND2_X1_322_ (
  .A1({ S2665 }),
  .A2({ S2662 }),
  .ZN({ S25957[659] })
);
NOR2_X1 #() 
NOR2_X1_1308_ (
  .A1({ S23140 }),
  .A2({ S23141 }),
  .ZN({ S25957[1008] })
);
NAND2_X1 #() 
NAND2_X1_5153_ (
  .A1({ S25859 }),
  .A2({ S25881 }),
  .ZN({ S2666 })
);
XOR2_X1 #() 
XOR2_X1_84_ (
  .A({ S2666 }),
  .B({ S25957[1008] }),
  .Z({ S2667 })
);
INV_X1 #() 
INV_X1_1685_ (
  .A({ S2667 }),
  .ZN({ S25957[880] })
);
AOI21_X1 #() 
AOI21_X1_2878_ (
  .A({ S101 }),
  .B1({ S2290 }),
  .B2({ S2395 }),
  .ZN({ S2668 })
);
AOI21_X1 #() 
AOI21_X1_2879_ (
  .A({ S101 }),
  .B1({ S2240 }),
  .B2({ S2257 }),
  .ZN({ S2669 })
);
NAND3_X1 #() 
NAND3_X1_5524_ (
  .A1({ S2262 }),
  .A2({ S2245 }),
  .A3({ S101 }),
  .ZN({ S2670 })
);
NAND2_X1 #() 
NAND2_X1_5154_ (
  .A1({ S2670 }),
  .A2({ S25957[780] }),
  .ZN({ S2671 })
);
NAND2_X1 #() 
NAND2_X1_5155_ (
  .A1({ S2298 }),
  .A2({ S2256 }),
  .ZN({ S2672 })
);
OAI22_X1 #() 
OAI22_X1_131_ (
  .A1({ S2669 }),
  .A2({ S2671 }),
  .B1({ S2668 }),
  .B2({ S2672 }),
  .ZN({ S2673 })
);
AOI21_X1 #() 
AOI21_X1_2880_ (
  .A({ S25957[776] }),
  .B1({ S2320 }),
  .B2({ S101 }),
  .ZN({ S2674 })
);
OAI21_X1 #() 
OAI21_X1_2671_ (
  .A({ S25957[780] }),
  .B1({ S2674 }),
  .B2({ S2384 }),
  .ZN({ S2675 })
);
AOI22_X1 #() 
AOI22_X1_578_ (
  .A1({ S2506 }),
  .A2({ S2492 }),
  .B1({ S2237 }),
  .B2({ S25957[778] }),
  .ZN({ S2676 })
);
OAI21_X1 #() 
OAI21_X1_2672_ (
  .A({ S2256 }),
  .B1({ S2676 }),
  .B2({ S2449 }),
  .ZN({ S2677 })
);
NAND3_X1 #() 
NAND3_X1_5525_ (
  .A1({ S2677 }),
  .A2({ S2315 }),
  .A3({ S2675 }),
  .ZN({ S2678 })
);
OAI211_X1 #() 
OAI211_X1_1813_ (
  .A({ S2678 }),
  .B({ S25957[782] }),
  .C1({ S2315 }),
  .C2({ S2673 }),
  .ZN({ S2679 })
);
AOI21_X1 #() 
AOI21_X1_2881_ (
  .A({ S25957[778] }),
  .B1({ S2282 }),
  .B2({ S25957[777] }),
  .ZN({ S2680 })
);
AOI21_X1 #() 
AOI21_X1_2882_ (
  .A({ S101 }),
  .B1({ S2680 }),
  .B2({ S2244 }),
  .ZN({ S2681 })
);
AOI21_X1 #() 
AOI21_X1_2883_ (
  .A({ S25957[779] }),
  .B1({ S2326 }),
  .B2({ S2338 }),
  .ZN({ S2682 })
);
OAI21_X1 #() 
OAI21_X1_2673_ (
  .A({ S25957[780] }),
  .B1({ S2682 }),
  .B2({ S2681 }),
  .ZN({ S2683 })
);
AOI21_X1 #() 
AOI21_X1_2884_ (
  .A({ S101 }),
  .B1({ S2282 }),
  .B2({ S2258 }),
  .ZN({ S2684 })
);
NAND2_X1 #() 
NAND2_X1_5156_ (
  .A1({ S2684 }),
  .A2({ S2629 }),
  .ZN({ S2685 })
);
OAI211_X1 #() 
OAI211_X1_1814_ (
  .A({ S2685 }),
  .B({ S2256 }),
  .C1({ S2297 }),
  .C2({ S2528 }),
  .ZN({ S2686 })
);
NAND3_X1 #() 
NAND3_X1_5526_ (
  .A1({ S2683 }),
  .A2({ S2315 }),
  .A3({ S2686 }),
  .ZN({ S2687 })
);
OAI21_X1 #() 
OAI21_X1_2674_ (
  .A({ S2256 }),
  .B1({ S2259 }),
  .B2({ S2299 }),
  .ZN({ S2688 })
);
NAND3_X1 #() 
NAND3_X1_5527_ (
  .A1({ S2493 }),
  .A2({ S2571 }),
  .A3({ S25957[780] }),
  .ZN({ S2689 })
);
OAI21_X1 #() 
OAI21_X1_2675_ (
  .A({ S2689 }),
  .B1({ S2688 }),
  .B2({ S2503 }),
  .ZN({ S2690 })
);
AOI21_X1 #() 
AOI21_X1_2885_ (
  .A({ S25957[782] }),
  .B1({ S2690 }),
  .B2({ S25957[781] }),
  .ZN({ S2691 })
);
NAND2_X1 #() 
NAND2_X1_5157_ (
  .A1({ S2691 }),
  .A2({ S2687 }),
  .ZN({ S2692 })
);
NAND3_X1 #() 
NAND3_X1_5528_ (
  .A1({ S2692 }),
  .A2({ S2679 }),
  .A3({ S2305 }),
  .ZN({ S2693 })
);
NAND4_X1 #() 
NAND4_X1_603_ (
  .A1({ S2244 }),
  .A2({ S2245 }),
  .A3({ S25957[779] }),
  .A4({ S25957[778] }),
  .ZN({ S2694 })
);
INV_X1 #() 
INV_X1_1686_ (
  .A({ S2694 }),
  .ZN({ S2695 })
);
OAI21_X1 #() 
OAI21_X1_2676_ (
  .A({ S25957[780] }),
  .B1({ S2549 }),
  .B2({ S2695 }),
  .ZN({ S2696 })
);
AOI21_X1 #() 
AOI21_X1_2886_ (
  .A({ S25957[781] }),
  .B1({ S2696 }),
  .B2({ S2490 }),
  .ZN({ S2697 })
);
OAI211_X1 #() 
OAI211_X1_1815_ (
  .A({ S2256 }),
  .B({ S2574 }),
  .C1({ S2343 }),
  .C2({ S2473 }),
  .ZN({ S2698 })
);
NAND2_X1 #() 
NAND2_X1_5158_ (
  .A1({ S2507 }),
  .A2({ S2245 }),
  .ZN({ S2699 })
);
NAND3_X1 #() 
NAND3_X1_5529_ (
  .A1({ S2572 }),
  .A2({ S2699 }),
  .A3({ S25957[780] }),
  .ZN({ S2700 })
);
AND3_X1 #() 
AND3_X1_217_ (
  .A1({ S2700 }),
  .A2({ S2698 }),
  .A3({ S25957[781] }),
  .ZN({ S2701 })
);
OAI21_X1 #() 
OAI21_X1_2677_ (
  .A({ S25957[782] }),
  .B1({ S2697 }),
  .B2({ S2701 }),
  .ZN({ S2702 })
);
OAI21_X1 #() 
OAI21_X1_2678_ (
  .A({ S2528 }),
  .B1({ S2550 }),
  .B2({ S2559 }),
  .ZN({ S2703 })
);
NAND2_X1 #() 
NAND2_X1_5159_ (
  .A1({ S2703 }),
  .A2({ S2256 }),
  .ZN({ S2704 })
);
NAND2_X1 #() 
NAND2_X1_5160_ (
  .A1({ S2605 }),
  .A2({ S2308 }),
  .ZN({ S2705 })
);
AOI21_X1 #() 
AOI21_X1_2887_ (
  .A({ S25957[776] }),
  .B1({ S25957[777] }),
  .B2({ S25957[778] }),
  .ZN({ S2706 })
);
AOI21_X1 #() 
AOI21_X1_2888_ (
  .A({ S2256 }),
  .B1({ S2706 }),
  .B2({ S101 }),
  .ZN({ S2707 })
);
NAND2_X1 #() 
NAND2_X1_5161_ (
  .A1({ S2705 }),
  .A2({ S2707 }),
  .ZN({ S2708 })
);
NAND3_X1 #() 
NAND3_X1_5530_ (
  .A1({ S2704 }),
  .A2({ S25957[781] }),
  .A3({ S2708 }),
  .ZN({ S2709 })
);
NAND3_X1 #() 
NAND3_X1_5531_ (
  .A1({ S2404 }),
  .A2({ S2400 }),
  .A3({ S25957[780] }),
  .ZN({ S2710 })
);
INV_X1 #() 
INV_X1_1687_ (
  .A({ S2492 }),
  .ZN({ S2711 })
);
AOI22_X1 #() 
AOI22_X1_579_ (
  .A1({ S2430 }),
  .A2({ S101 }),
  .B1({ S2248 }),
  .B2({ S2711 }),
  .ZN({ S2712 })
);
OAI211_X1 #() 
OAI211_X1_1816_ (
  .A({ S2315 }),
  .B({ S2710 }),
  .C1({ S2712 }),
  .C2({ S25957[780] }),
  .ZN({ S2713 })
);
NAND3_X1 #() 
NAND3_X1_5532_ (
  .A1({ S2709 }),
  .A2({ S2713 }),
  .A3({ S2268 }),
  .ZN({ S2714 })
);
NAND3_X1 #() 
NAND3_X1_5533_ (
  .A1({ S2702 }),
  .A2({ S25957[783] }),
  .A3({ S2714 }),
  .ZN({ S2715 })
);
NAND3_X1 #() 
NAND3_X1_5534_ (
  .A1({ S2715 }),
  .A2({ S25957[880] }),
  .A3({ S2693 }),
  .ZN({ S2716 })
);
AOI22_X1 #() 
AOI22_X1_580_ (
  .A1({ S2258 }),
  .A2({ S25957[776] }),
  .B1({ S1010 }),
  .B2({ S1013 }),
  .ZN({ S2717 })
);
OAI21_X1 #() 
OAI21_X1_2679_ (
  .A({ S101 }),
  .B1({ S2680 }),
  .B2({ S2717 }),
  .ZN({ S2718 })
);
AOI21_X1 #() 
AOI21_X1_2889_ (
  .A({ S2256 }),
  .B1({ S2718 }),
  .B2({ S2694 }),
  .ZN({ S2719 })
);
OAI21_X1 #() 
OAI21_X1_2680_ (
  .A({ S2315 }),
  .B1({ S2719 }),
  .B2({ S2489 }),
  .ZN({ S2720 })
);
NAND3_X1 #() 
NAND3_X1_5535_ (
  .A1({ S2700 }),
  .A2({ S2698 }),
  .A3({ S25957[781] }),
  .ZN({ S2721 })
);
AOI21_X1 #() 
AOI21_X1_2890_ (
  .A({ S2268 }),
  .B1({ S2720 }),
  .B2({ S2721 }),
  .ZN({ S2722 })
);
AND3_X1 #() 
AND3_X1_218_ (
  .A1({ S2709 }),
  .A2({ S2713 }),
  .A3({ S2268 }),
  .ZN({ S2723 })
);
OAI21_X1 #() 
OAI21_X1_2681_ (
  .A({ S25957[783] }),
  .B1({ S2722 }),
  .B2({ S2723 }),
  .ZN({ S2724 })
);
NAND2_X1 #() 
NAND2_X1_5162_ (
  .A1({ S2240 }),
  .A2({ S2257 }),
  .ZN({ S2725 })
);
AOI21_X1 #() 
AOI21_X1_2891_ (
  .A({ S2671 }),
  .B1({ S2725 }),
  .B2({ S25957[779] }),
  .ZN({ S2726 })
);
NOR2_X1 #() 
NOR2_X1_1309_ (
  .A1({ S2668 }),
  .A2({ S2672 }),
  .ZN({ S2727 })
);
OAI21_X1 #() 
OAI21_X1_2682_ (
  .A({ S25957[781] }),
  .B1({ S2726 }),
  .B2({ S2727 }),
  .ZN({ S2728 })
);
NOR2_X1 #() 
NOR2_X1_1310_ (
  .A1({ S2711 }),
  .A2({ S2256 }),
  .ZN({ S2729 })
);
AOI21_X1 #() 
AOI21_X1_2892_ (
  .A({ S25957[781] }),
  .B1({ S2729 }),
  .B2({ S2417 }),
  .ZN({ S2730 })
);
OAI21_X1 #() 
OAI21_X1_2683_ (
  .A({ S2730 }),
  .B1({ S2561 }),
  .B2({ S2449 }),
  .ZN({ S2731 })
);
AOI21_X1 #() 
AOI21_X1_2893_ (
  .A({ S2268 }),
  .B1({ S2728 }),
  .B2({ S2731 }),
  .ZN({ S2732 })
);
NAND2_X1 #() 
NAND2_X1_5163_ (
  .A1({ S2263 }),
  .A2({ S2270 }),
  .ZN({ S2733 })
);
AOI22_X1 #() 
AOI22_X1_581_ (
  .A1({ S2733 }),
  .A2({ S2296 }),
  .B1({ S2684 }),
  .B2({ S2629 }),
  .ZN({ S2734 })
);
AOI21_X1 #() 
AOI21_X1_2894_ (
  .A({ S2256 }),
  .B1({ S2264 }),
  .B2({ S101 }),
  .ZN({ S2735 })
);
OAI211_X1 #() 
OAI211_X1_1817_ (
  .A({ S2735 }),
  .B({ S2345 }),
  .C1({ S2643 }),
  .C2({ S101 }),
  .ZN({ S2736 })
);
OAI211_X1 #() 
OAI211_X1_1818_ (
  .A({ S2736 }),
  .B({ S2315 }),
  .C1({ S2734 }),
  .C2({ S25957[780] }),
  .ZN({ S2737 })
);
OAI211_X1 #() 
OAI211_X1_1819_ (
  .A({ S2689 }),
  .B({ S25957[781] }),
  .C1({ S2688 }),
  .C2({ S2503 }),
  .ZN({ S2738 })
);
AOI21_X1 #() 
AOI21_X1_2895_ (
  .A({ S25957[782] }),
  .B1({ S2737 }),
  .B2({ S2738 }),
  .ZN({ S2739 })
);
OAI21_X1 #() 
OAI21_X1_2684_ (
  .A({ S2305 }),
  .B1({ S2732 }),
  .B2({ S2739 }),
  .ZN({ S2740 })
);
NAND3_X1 #() 
NAND3_X1_5536_ (
  .A1({ S2724 }),
  .A2({ S2740 }),
  .A3({ S2667 }),
  .ZN({ S2741 })
);
NAND3_X1 #() 
NAND3_X1_5537_ (
  .A1({ S2741 }),
  .A2({ S2716 }),
  .A3({ S25957[944] }),
  .ZN({ S2742 })
);
NAND3_X1 #() 
NAND3_X1_5538_ (
  .A1({ S2715 }),
  .A2({ S2667 }),
  .A3({ S2693 }),
  .ZN({ S2743 })
);
NAND3_X1 #() 
NAND3_X1_5539_ (
  .A1({ S2724 }),
  .A2({ S2740 }),
  .A3({ S25957[880] }),
  .ZN({ S2744 })
);
NAND3_X1 #() 
NAND3_X1_5540_ (
  .A1({ S2744 }),
  .A2({ S2743 }),
  .A3({ S25834 }),
  .ZN({ S2745 })
);
NAND3_X1 #() 
NAND3_X1_5541_ (
  .A1({ S2742 }),
  .A2({ S2745 }),
  .A3({ S25957[784] }),
  .ZN({ S2746 })
);
NAND3_X1 #() 
NAND3_X1_5542_ (
  .A1({ S25917 }),
  .A2({ S25921 }),
  .A3({ S25914 }),
  .ZN({ S2747 })
);
NAND3_X1 #() 
NAND3_X1_5543_ (
  .A1({ S25922 }),
  .A2({ S25957[912] }),
  .A3({ S25923 }),
  .ZN({ S2748 })
);
NAND2_X1 #() 
NAND2_X1_5164_ (
  .A1({ S2747 }),
  .A2({ S2748 }),
  .ZN({ S2749 })
);
NAND3_X1 #() 
NAND3_X1_5544_ (
  .A1({ S2744 }),
  .A2({ S2743 }),
  .A3({ S25957[944] }),
  .ZN({ S2750 })
);
NAND3_X1 #() 
NAND3_X1_5545_ (
  .A1({ S2741 }),
  .A2({ S2716 }),
  .A3({ S25834 }),
  .ZN({ S2751 })
);
NAND3_X1 #() 
NAND3_X1_5546_ (
  .A1({ S2750 }),
  .A2({ S2751 }),
  .A3({ S2749 }),
  .ZN({ S2752 })
);
NAND2_X1 #() 
NAND2_X1_5165_ (
  .A1({ S2746 }),
  .A2({ S2752 }),
  .ZN({ S25957[656] })
);
NOR2_X1 #() 
NOR2_X1_1311_ (
  .A1({ S259 }),
  .A2({ S258 }),
  .ZN({ S2753 })
);
INV_X1 #() 
INV_X1_1688_ (
  .A({ S2753 }),
  .ZN({ S25957[849] })
);
NAND2_X1 #() 
NAND2_X1_5166_ (
  .A1({ S23269 }),
  .A2({ S23268 }),
  .ZN({ S25957[1009] })
);
NAND2_X1 #() 
NAND2_X1_5167_ (
  .A1({ S255 }),
  .A2({ S250 }),
  .ZN({ S2754 })
);
XOR2_X1 #() 
XOR2_X1_85_ (
  .A({ S2754 }),
  .B({ S25957[1009] }),
  .Z({ S2755 })
);
NAND2_X1 #() 
NAND2_X1_5168_ (
  .A1({ S2323 }),
  .A2({ S101 }),
  .ZN({ S2756 })
);
NAND2_X1 #() 
NAND2_X1_5169_ (
  .A1({ S2756 }),
  .A2({ S2256 }),
  .ZN({ S2757 })
);
AND2_X1 #() 
AND2_X1_323_ (
  .A1({ S2638 }),
  .A2({ S2526 }),
  .ZN({ S2758 })
);
OAI211_X1 #() 
OAI211_X1_1820_ (
  .A({ S2757 }),
  .B({ S25957[781] }),
  .C1({ S2758 }),
  .C2({ S2256 }),
  .ZN({ S2759 })
);
NAND3_X1 #() 
NAND3_X1_5547_ (
  .A1({ S2535 }),
  .A2({ S2271 }),
  .A3({ S25957[780] }),
  .ZN({ S2760 })
);
NAND3_X1 #() 
NAND3_X1_5548_ (
  .A1({ S2603 }),
  .A2({ S2256 }),
  .A3({ S2265 }),
  .ZN({ S2761 })
);
NAND2_X1 #() 
NAND2_X1_5170_ (
  .A1({ S2760 }),
  .A2({ S2761 }),
  .ZN({ S2762 })
);
NAND2_X1 #() 
NAND2_X1_5171_ (
  .A1({ S2762 }),
  .A2({ S2315 }),
  .ZN({ S2763 })
);
NAND3_X1 #() 
NAND3_X1_5549_ (
  .A1({ S2763 }),
  .A2({ S2759 }),
  .A3({ S2268 }),
  .ZN({ S2764 })
);
OAI211_X1 #() 
OAI211_X1_1821_ (
  .A({ S2614 }),
  .B({ S25957[780] }),
  .C1({ S2376 }),
  .C2({ S2528 }),
  .ZN({ S2765 })
);
AOI21_X1 #() 
AOI21_X1_2896_ (
  .A({ S2269 }),
  .B1({ S2466 }),
  .B2({ S2258 }),
  .ZN({ S2766 })
);
AOI21_X1 #() 
AOI21_X1_2897_ (
  .A({ S2315 }),
  .B1({ S2766 }),
  .B2({ S2464 }),
  .ZN({ S2767 })
);
OAI211_X1 #() 
OAI211_X1_1822_ (
  .A({ S2694 }),
  .B({ S2256 }),
  .C1({ S2379 }),
  .C2({ S2376 }),
  .ZN({ S2768 })
);
OAI21_X1 #() 
OAI21_X1_2685_ (
  .A({ S25957[779] }),
  .B1({ S2342 }),
  .B2({ S2307 }),
  .ZN({ S2769 })
);
NAND2_X1 #() 
NAND2_X1_5172_ (
  .A1({ S2298 }),
  .A2({ S2270 }),
  .ZN({ S2770 })
);
AOI21_X1 #() 
AOI21_X1_2898_ (
  .A({ S2256 }),
  .B1({ S2770 }),
  .B2({ S2629 }),
  .ZN({ S2771 })
);
AOI21_X1 #() 
AOI21_X1_2899_ (
  .A({ S25957[781] }),
  .B1({ S2771 }),
  .B2({ S2769 }),
  .ZN({ S2772 })
);
AOI22_X1 #() 
AOI22_X1_582_ (
  .A1({ S2772 }),
  .A2({ S2768 }),
  .B1({ S2767 }),
  .B2({ S2765 }),
  .ZN({ S2773 })
);
OAI211_X1 #() 
OAI211_X1_1823_ (
  .A({ S2305 }),
  .B({ S2764 }),
  .C1({ S2773 }),
  .C2({ S2268 }),
  .ZN({ S2774 })
);
NAND2_X1 #() 
NAND2_X1_5173_ (
  .A1({ S2496 }),
  .A2({ S2707 }),
  .ZN({ S2775 })
);
NAND3_X1 #() 
NAND3_X1_5550_ (
  .A1({ S2237 }),
  .A2({ S25957[779] }),
  .A3({ S2262 }),
  .ZN({ S2776 })
);
INV_X1 #() 
INV_X1_1689_ (
  .A({ S2262 }),
  .ZN({ S2777 })
);
AOI21_X1 #() 
AOI21_X1_2900_ (
  .A({ S25957[780] }),
  .B1({ S2777 }),
  .B2({ S101 }),
  .ZN({ S2778 })
);
NAND3_X1 #() 
NAND3_X1_5551_ (
  .A1({ S2778 }),
  .A2({ S2400 }),
  .A3({ S2776 }),
  .ZN({ S2779 })
);
NAND3_X1 #() 
NAND3_X1_5552_ (
  .A1({ S2775 }),
  .A2({ S2779 }),
  .A3({ S2315 }),
  .ZN({ S2780 })
);
NAND3_X1 #() 
NAND3_X1_5553_ (
  .A1({ S2333 }),
  .A2({ S2256 }),
  .A3({ S2337 }),
  .ZN({ S2781 })
);
NAND3_X1 #() 
NAND3_X1_5554_ (
  .A1({ S2621 }),
  .A2({ S25957[780] }),
  .A3({ S2379 }),
  .ZN({ S2782 })
);
OAI211_X1 #() 
OAI211_X1_1824_ (
  .A({ S2782 }),
  .B({ S25957[781] }),
  .C1({ S2669 }),
  .C2({ S2781 }),
  .ZN({ S2783 })
);
NAND2_X1 #() 
NAND2_X1_5174_ (
  .A1({ S2780 }),
  .A2({ S2783 }),
  .ZN({ S2784 })
);
NAND2_X1 #() 
NAND2_X1_5175_ (
  .A1({ S2784 }),
  .A2({ S25957[782] }),
  .ZN({ S2785 })
);
NAND2_X1 #() 
NAND2_X1_5176_ (
  .A1({ S2326 }),
  .A2({ S2273 }),
  .ZN({ S2786 })
);
AOI22_X1 #() 
AOI22_X1_583_ (
  .A1({ S2786 }),
  .A2({ S25957[779] }),
  .B1({ S2309 }),
  .B2({ S2290 }),
  .ZN({ S2787 })
);
OAI211_X1 #() 
OAI211_X1_1825_ (
  .A({ S2454 }),
  .B({ S2256 }),
  .C1({ S2333 }),
  .C2({ S2470 }),
  .ZN({ S2788 })
);
OAI211_X1 #() 
OAI211_X1_1826_ (
  .A({ S25957[781] }),
  .B({ S2788 }),
  .C1({ S2787 }),
  .C2({ S2256 }),
  .ZN({ S2789 })
);
AOI21_X1 #() 
AOI21_X1_2901_ (
  .A({ S25957[779] }),
  .B1({ S25957[778] }),
  .B2({ S2245 }),
  .ZN({ S2790 })
);
AOI22_X1 #() 
AOI22_X1_584_ (
  .A1({ S2546 }),
  .A2({ S25957[779] }),
  .B1({ S2790 }),
  .B2({ S2495 }),
  .ZN({ S2791 })
);
OAI211_X1 #() 
OAI211_X1_1827_ (
  .A({ S2285 }),
  .B({ S101 }),
  .C1({ S2245 }),
  .C2({ S25957[778] }),
  .ZN({ S2792 })
);
NAND2_X1 #() 
NAND2_X1_5177_ (
  .A1({ S2368 }),
  .A2({ S2792 }),
  .ZN({ S2793 })
);
NAND2_X1 #() 
NAND2_X1_5178_ (
  .A1({ S2793 }),
  .A2({ S25957[780] }),
  .ZN({ S2794 })
);
OAI211_X1 #() 
OAI211_X1_1828_ (
  .A({ S2315 }),
  .B({ S2794 }),
  .C1({ S2791 }),
  .C2({ S25957[780] }),
  .ZN({ S2795 })
);
NAND3_X1 #() 
NAND3_X1_5555_ (
  .A1({ S2789 }),
  .A2({ S2795 }),
  .A3({ S2268 }),
  .ZN({ S2796 })
);
NAND3_X1 #() 
NAND3_X1_5556_ (
  .A1({ S2796 }),
  .A2({ S2785 }),
  .A3({ S25957[783] }),
  .ZN({ S2797 })
);
NAND3_X1 #() 
NAND3_X1_5557_ (
  .A1({ S2797 }),
  .A2({ S2774 }),
  .A3({ S2755 }),
  .ZN({ S2798 })
);
INV_X1 #() 
INV_X1_1690_ (
  .A({ S2755 }),
  .ZN({ S25957[881] })
);
OAI21_X1 #() 
OAI21_X1_2686_ (
  .A({ S2256 }),
  .B1({ S2455 }),
  .B2({ S2487 }),
  .ZN({ S2799 })
);
OAI22_X1 #() 
OAI22_X1_132_ (
  .A1({ S2799 }),
  .A2({ S2325 }),
  .B1({ S2793 }),
  .B2({ S2256 }),
  .ZN({ S2800 })
);
AOI21_X1 #() 
AOI21_X1_2902_ (
  .A({ S25957[782] }),
  .B1({ S2800 }),
  .B2({ S2315 }),
  .ZN({ S2801 })
);
AOI22_X1 #() 
AOI22_X1_585_ (
  .A1({ S2801 }),
  .A2({ S2789 }),
  .B1({ S2784 }),
  .B2({ S25957[782] }),
  .ZN({ S2802 })
);
NAND3_X1 #() 
NAND3_X1_5558_ (
  .A1({ S2760 }),
  .A2({ S2761 }),
  .A3({ S2315 }),
  .ZN({ S2803 })
);
AOI21_X1 #() 
AOI21_X1_2903_ (
  .A({ S2256 }),
  .B1({ S2638 }),
  .B2({ S2526 }),
  .ZN({ S2804 })
);
OAI21_X1 #() 
OAI21_X1_2687_ (
  .A({ S25957[781] }),
  .B1({ S2804 }),
  .B2({ S2324 }),
  .ZN({ S2805 })
);
AOI21_X1 #() 
AOI21_X1_2904_ (
  .A({ S25957[782] }),
  .B1({ S2805 }),
  .B2({ S2803 }),
  .ZN({ S2806 })
);
NAND2_X1 #() 
NAND2_X1_5179_ (
  .A1({ S2767 }),
  .A2({ S2765 }),
  .ZN({ S2807 })
);
INV_X1 #() 
INV_X1_1691_ (
  .A({ S2629 }),
  .ZN({ S2808 })
);
OAI21_X1 #() 
OAI21_X1_2688_ (
  .A({ S25957[780] }),
  .B1({ S2808 }),
  .B2({ S2274 }),
  .ZN({ S2809 })
);
OAI211_X1 #() 
OAI211_X1_1829_ (
  .A({ S2768 }),
  .B({ S2315 }),
  .C1({ S2809 }),
  .C2({ S2669 }),
  .ZN({ S2810 })
);
AOI21_X1 #() 
AOI21_X1_2905_ (
  .A({ S2268 }),
  .B1({ S2810 }),
  .B2({ S2807 }),
  .ZN({ S2811 })
);
OAI21_X1 #() 
OAI21_X1_2689_ (
  .A({ S2305 }),
  .B1({ S2811 }),
  .B2({ S2806 }),
  .ZN({ S2812 })
);
OAI211_X1 #() 
OAI211_X1_1830_ (
  .A({ S2812 }),
  .B({ S25957[881] }),
  .C1({ S2802 }),
  .C2({ S2305 }),
  .ZN({ S2813 })
);
NAND3_X1 #() 
NAND3_X1_5559_ (
  .A1({ S2813 }),
  .A2({ S2798 }),
  .A3({ S25957[849] }),
  .ZN({ S2814 })
);
NAND3_X1 #() 
NAND3_X1_5560_ (
  .A1({ S2797 }),
  .A2({ S2774 }),
  .A3({ S25957[881] }),
  .ZN({ S2815 })
);
OAI211_X1 #() 
OAI211_X1_1831_ (
  .A({ S2812 }),
  .B({ S2755 }),
  .C1({ S2802 }),
  .C2({ S2305 }),
  .ZN({ S2816 })
);
NAND3_X1 #() 
NAND3_X1_5561_ (
  .A1({ S2816 }),
  .A2({ S2815 }),
  .A3({ S2753 }),
  .ZN({ S2817 })
);
AOI21_X1 #() 
AOI21_X1_2906_ (
  .A({ S25957[913] }),
  .B1({ S2814 }),
  .B2({ S2817 }),
  .ZN({ S2818 })
);
AND3_X1 #() 
AND3_X1_219_ (
  .A1({ S2817 }),
  .A2({ S2814 }),
  .A3({ S25957[913] }),
  .ZN({ S2819 })
);
NOR2_X1 #() 
NOR2_X1_1312_ (
  .A1({ S2819 }),
  .A2({ S2818 }),
  .ZN({ S25957[657] })
);
NOR2_X1 #() 
NOR2_X1_1313_ (
  .A1({ S345 }),
  .A2({ S346 }),
  .ZN({ S25957[978] })
);
NAND2_X1 #() 
NAND2_X1_5180_ (
  .A1({ S2250 }),
  .A2({ S25957[777] }),
  .ZN({ S2820 })
);
NAND4_X1 #() 
NAND4_X1_604_ (
  .A1({ S2820 }),
  .A2({ S2262 }),
  .A3({ S25957[779] }),
  .A4({ S2296 }),
  .ZN({ S2821 })
);
AOI22_X1 #() 
AOI22_X1_586_ (
  .A1({ S2334 }),
  .A2({ S2320 }),
  .B1({ S2264 }),
  .B2({ S101 }),
  .ZN({ S2822 })
);
AOI21_X1 #() 
AOI21_X1_2907_ (
  .A({ S2256 }),
  .B1({ S2473 }),
  .B2({ S101 }),
  .ZN({ S2823 })
);
AOI22_X1 #() 
AOI22_X1_587_ (
  .A1({ S2822 }),
  .A2({ S2256 }),
  .B1({ S2821 }),
  .B2({ S2823 }),
  .ZN({ S2824 })
);
OAI211_X1 #() 
OAI211_X1_1832_ (
  .A({ S25957[779] }),
  .B({ S2450 }),
  .C1({ S2331 }),
  .C2({ S2470 }),
  .ZN({ S2825 })
);
NAND3_X1 #() 
NAND3_X1_5562_ (
  .A1({ S2825 }),
  .A2({ S2256 }),
  .A3({ S2333 }),
  .ZN({ S2826 })
);
NAND3_X1 #() 
NAND3_X1_5563_ (
  .A1({ S2259 }),
  .A2({ S101 }),
  .A3({ S2257 }),
  .ZN({ S2827 })
);
AOI21_X1 #() 
AOI21_X1_2908_ (
  .A({ S2256 }),
  .B1({ S2321 }),
  .B2({ S2320 }),
  .ZN({ S2828 })
);
AOI21_X1 #() 
AOI21_X1_2909_ (
  .A({ S2315 }),
  .B1({ S2828 }),
  .B2({ S2827 }),
  .ZN({ S2829 })
);
AOI22_X1 #() 
AOI22_X1_588_ (
  .A1({ S2824 }),
  .A2({ S2315 }),
  .B1({ S2829 }),
  .B2({ S2826 }),
  .ZN({ S2830 })
);
NAND2_X1 #() 
NAND2_X1_5181_ (
  .A1({ S2367 }),
  .A2({ S101 }),
  .ZN({ S2831 })
);
NAND2_X1 #() 
NAND2_X1_5182_ (
  .A1({ S2820 }),
  .A2({ S25957[779] }),
  .ZN({ S2832 })
);
NAND3_X1 #() 
NAND3_X1_5564_ (
  .A1({ S2832 }),
  .A2({ S25957[780] }),
  .A3({ S2831 }),
  .ZN({ S2833 })
);
OAI211_X1 #() 
OAI211_X1_1833_ (
  .A({ S2833 }),
  .B({ S2315 }),
  .C1({ S25957[780] }),
  .C2({ S2422 }),
  .ZN({ S2834 })
);
NAND4_X1 #() 
NAND4_X1_605_ (
  .A1({ S2694 }),
  .A2({ S2411 }),
  .A3({ S2454 }),
  .A4({ S2256 }),
  .ZN({ S2835 })
);
NAND3_X1 #() 
NAND3_X1_5565_ (
  .A1({ S2405 }),
  .A2({ S2603 }),
  .A3({ S25957[780] }),
  .ZN({ S2836 })
);
NAND2_X1 #() 
NAND2_X1_5183_ (
  .A1({ S2835 }),
  .A2({ S2836 }),
  .ZN({ S2837 })
);
NAND2_X1 #() 
NAND2_X1_5184_ (
  .A1({ S2837 }),
  .A2({ S25957[781] }),
  .ZN({ S2838 })
);
NAND3_X1 #() 
NAND3_X1_5566_ (
  .A1({ S2838 }),
  .A2({ S2834 }),
  .A3({ S2268 }),
  .ZN({ S2839 })
);
OAI211_X1 #() 
OAI211_X1_1834_ (
  .A({ S2839 }),
  .B({ S25957[783] }),
  .C1({ S2830 }),
  .C2({ S2268 }),
  .ZN({ S2840 })
);
INV_X1 #() 
INV_X1_1692_ (
  .A({ S2500 }),
  .ZN({ S2841 })
);
NAND2_X1 #() 
NAND2_X1_5185_ (
  .A1({ S2321 }),
  .A2({ S2495 }),
  .ZN({ S2842 })
);
NAND4_X1 #() 
NAND4_X1_606_ (
  .A1({ S2842 }),
  .A2({ S2841 }),
  .A3({ S2605 }),
  .A4({ S25957[780] }),
  .ZN({ S2843 })
);
NAND3_X1 #() 
NAND3_X1_5567_ (
  .A1({ S2718 }),
  .A2({ S2256 }),
  .A3({ S2832 }),
  .ZN({ S2844 })
);
NAND2_X1 #() 
NAND2_X1_5186_ (
  .A1({ S2844 }),
  .A2({ S2843 }),
  .ZN({ S2845 })
);
NAND2_X1 #() 
NAND2_X1_5187_ (
  .A1({ S2845 }),
  .A2({ S2315 }),
  .ZN({ S2846 })
);
NAND3_X1 #() 
NAND3_X1_5568_ (
  .A1({ S2338 }),
  .A2({ S25957[779] }),
  .A3({ S2244 }),
  .ZN({ S2847 })
);
AOI21_X1 #() 
AOI21_X1_2910_ (
  .A({ S2256 }),
  .B1({ S2847 }),
  .B2({ S2605 }),
  .ZN({ S2848 })
);
INV_X1 #() 
INV_X1_1693_ (
  .A({ S2848 }),
  .ZN({ S2849 })
);
OAI21_X1 #() 
OAI21_X1_2690_ (
  .A({ S2256 }),
  .B1({ S2446 }),
  .B2({ S2263 }),
  .ZN({ S2850 })
);
OAI211_X1 #() 
OAI211_X1_1835_ (
  .A({ S2849 }),
  .B({ S25957[781] }),
  .C1({ S2247 }),
  .C2({ S2850 }),
  .ZN({ S2851 })
);
NAND3_X1 #() 
NAND3_X1_5569_ (
  .A1({ S2846 }),
  .A2({ S25957[782] }),
  .A3({ S2851 }),
  .ZN({ S2852 })
);
AOI21_X1 #() 
AOI21_X1_2911_ (
  .A({ S25957[781] }),
  .B1({ S2396 }),
  .B2({ S2291 }),
  .ZN({ S2853 })
);
AOI21_X1 #() 
AOI21_X1_2912_ (
  .A({ S101 }),
  .B1({ S2248 }),
  .B2({ S2245 }),
  .ZN({ S2854 })
);
OAI21_X1 #() 
OAI21_X1_2691_ (
  .A({ S25957[780] }),
  .B1({ S2541 }),
  .B2({ S2854 }),
  .ZN({ S2855 })
);
NAND2_X1 #() 
NAND2_X1_5188_ (
  .A1({ S2260 }),
  .A2({ S2293 }),
  .ZN({ S2856 })
);
NAND3_X1 #() 
NAND3_X1_5570_ (
  .A1({ S2855 }),
  .A2({ S2853 }),
  .A3({ S2856 }),
  .ZN({ S2857 })
);
NAND2_X1 #() 
NAND2_X1_5189_ (
  .A1({ S2467 }),
  .A2({ S2321 }),
  .ZN({ S2858 })
);
AOI21_X1 #() 
AOI21_X1_2913_ (
  .A({ S2256 }),
  .B1({ S2639 }),
  .B2({ S2858 }),
  .ZN({ S2859 })
);
NOR2_X1 #() 
NOR2_X1_1314_ (
  .A1({ S2270 }),
  .A2({ S2273 }),
  .ZN({ S2860 })
);
AOI21_X1 #() 
AOI21_X1_2914_ (
  .A({ S2860 }),
  .B1({ S2481 }),
  .B2({ S25957[779] }),
  .ZN({ S2861 })
);
OAI21_X1 #() 
OAI21_X1_2692_ (
  .A({ S25957[781] }),
  .B1({ S2861 }),
  .B2({ S25957[780] }),
  .ZN({ S2862 })
);
OAI211_X1 #() 
OAI211_X1_1836_ (
  .A({ S2857 }),
  .B({ S2268 }),
  .C1({ S2862 }),
  .C2({ S2859 }),
  .ZN({ S2863 })
);
NAND3_X1 #() 
NAND3_X1_5571_ (
  .A1({ S2852 }),
  .A2({ S2863 }),
  .A3({ S2305 }),
  .ZN({ S2864 })
);
AOI21_X1 #() 
AOI21_X1_2915_ (
  .A({ S25957[978] }),
  .B1({ S2864 }),
  .B2({ S2840 }),
  .ZN({ S2865 })
);
INV_X1 #() 
INV_X1_1694_ (
  .A({ S25957[978] }),
  .ZN({ S2866 })
);
NAND2_X1 #() 
NAND2_X1_5190_ (
  .A1({ S2821 }),
  .A2({ S2823 }),
  .ZN({ S2867 })
);
NAND2_X1 #() 
NAND2_X1_5191_ (
  .A1({ S2822 }),
  .A2({ S2256 }),
  .ZN({ S2868 })
);
NAND3_X1 #() 
NAND3_X1_5572_ (
  .A1({ S2868 }),
  .A2({ S2315 }),
  .A3({ S2867 }),
  .ZN({ S2869 })
);
NAND2_X1 #() 
NAND2_X1_5192_ (
  .A1({ S2829 }),
  .A2({ S2826 }),
  .ZN({ S2870 })
);
NAND3_X1 #() 
NAND3_X1_5573_ (
  .A1({ S2870 }),
  .A2({ S2869 }),
  .A3({ S25957[782] }),
  .ZN({ S2871 })
);
NAND2_X1 #() 
NAND2_X1_5193_ (
  .A1({ S2838 }),
  .A2({ S2834 }),
  .ZN({ S2872 })
);
NAND2_X1 #() 
NAND2_X1_5194_ (
  .A1({ S2872 }),
  .A2({ S2268 }),
  .ZN({ S2873 })
);
NAND3_X1 #() 
NAND3_X1_5574_ (
  .A1({ S2873 }),
  .A2({ S2871 }),
  .A3({ S25957[783] }),
  .ZN({ S2874 })
);
NOR2_X1 #() 
NOR2_X1_1315_ (
  .A1({ S2247 }),
  .A2({ S2850 }),
  .ZN({ S2875 })
);
OAI21_X1 #() 
OAI21_X1_2693_ (
  .A({ S25957[781] }),
  .B1({ S2875 }),
  .B2({ S2848 }),
  .ZN({ S2876 })
);
NAND3_X1 #() 
NAND3_X1_5575_ (
  .A1({ S2844 }),
  .A2({ S2843 }),
  .A3({ S2315 }),
  .ZN({ S2877 })
);
NAND3_X1 #() 
NAND3_X1_5576_ (
  .A1({ S2876 }),
  .A2({ S25957[782] }),
  .A3({ S2877 }),
  .ZN({ S2878 })
);
AND2_X1 #() 
AND2_X1_324_ (
  .A1({ S2853 }),
  .A2({ S2856 }),
  .ZN({ S2879 })
);
INV_X1 #() 
INV_X1_1695_ (
  .A({ S2859 }),
  .ZN({ S2880 })
);
NAND3_X1 #() 
NAND3_X1_5577_ (
  .A1({ S2331 }),
  .A2({ S2629 }),
  .A3({ S25957[779] }),
  .ZN({ S2881 })
);
NAND2_X1 #() 
NAND2_X1_5195_ (
  .A1({ S2881 }),
  .A2({ S2509 }),
  .ZN({ S2882 })
);
AOI21_X1 #() 
AOI21_X1_2916_ (
  .A({ S2315 }),
  .B1({ S2882 }),
  .B2({ S2256 }),
  .ZN({ S2883 })
);
AOI22_X1 #() 
AOI22_X1_589_ (
  .A1({ S2880 }),
  .A2({ S2883 }),
  .B1({ S2879 }),
  .B2({ S2855 }),
  .ZN({ S2884 })
);
OAI211_X1 #() 
OAI211_X1_1837_ (
  .A({ S2878 }),
  .B({ S2305 }),
  .C1({ S2884 }),
  .C2({ S25957[782] }),
  .ZN({ S2885 })
);
AOI21_X1 #() 
AOI21_X1_2917_ (
  .A({ S2866 }),
  .B1({ S2885 }),
  .B2({ S2874 }),
  .ZN({ S2886 })
);
OAI21_X1 #() 
OAI21_X1_2694_ (
  .A({ S349 }),
  .B1({ S2886 }),
  .B2({ S2865 }),
  .ZN({ S2887 })
);
NAND3_X1 #() 
NAND3_X1_5578_ (
  .A1({ S2885 }),
  .A2({ S2866 }),
  .A3({ S2874 }),
  .ZN({ S2888 })
);
NAND3_X1 #() 
NAND3_X1_5579_ (
  .A1({ S2864 }),
  .A2({ S2840 }),
  .A3({ S25957[978] }),
  .ZN({ S2889 })
);
NAND3_X1 #() 
NAND3_X1_5580_ (
  .A1({ S2888 }),
  .A2({ S2889 }),
  .A3({ S25957[914] }),
  .ZN({ S2890 })
);
NAND2_X1 #() 
NAND2_X1_5196_ (
  .A1({ S2887 }),
  .A2({ S2890 }),
  .ZN({ S25957[658] })
);
NAND3_X1 #() 
NAND3_X1_5581_ (
  .A1({ S1559 }),
  .A2({ S1558 }),
  .A3({ S25957[897] }),
  .ZN({ S2891 })
);
NAND3_X1 #() 
NAND3_X1_5582_ (
  .A1({ S1551 }),
  .A2({ S1556 }),
  .A3({ S490 }),
  .ZN({ S2892 })
);
NAND3_X1 #() 
NAND3_X1_5583_ (
  .A1({ S25957[768] }),
  .A2({ S2891 }),
  .A3({ S2892 }),
  .ZN({ S2893 })
);
INV_X1 #() 
INV_X1_1696_ (
  .A({ S2893 }),
  .ZN({ S111 })
);
AOI21_X1 #() 
AOI21_X1_2918_ (
  .A({ S24456 }),
  .B1({ S1507 }),
  .B2({ S1487 }),
  .ZN({ S2894 })
);
AOI21_X1 #() 
AOI21_X1_2919_ (
  .A({ S25957[1088] }),
  .B1({ S1439 }),
  .B2({ S1462 }),
  .ZN({ S2895 })
);
OAI21_X1 #() 
OAI21_X1_2695_ (
  .A({ S23360 }),
  .B1({ S2894 }),
  .B2({ S2895 }),
  .ZN({ S2896 })
);
NAND3_X1 #() 
NAND3_X1_5584_ (
  .A1({ S1508 }),
  .A2({ S1463 }),
  .A3({ S25957[1024] }),
  .ZN({ S2897 })
);
NAND2_X1 #() 
NAND2_X1_5197_ (
  .A1({ S2896 }),
  .A2({ S2897 }),
  .ZN({ S2898 })
);
NAND3_X1 #() 
NAND3_X1_5585_ (
  .A1({ S2898 }),
  .A2({ S1557 }),
  .A3({ S1560 }),
  .ZN({ S112 })
);
XNOR2_X1 #() 
XNOR2_X1_199_ (
  .A({ S23473 }),
  .B({ S25957[1135] }),
  .ZN({ S25957[1007] })
);
XNOR2_X1 #() 
XNOR2_X1_200_ (
  .A({ S469 }),
  .B({ S25957[1007] }),
  .ZN({ S25957[879] })
);
INV_X1 #() 
INV_X1_1697_ (
  .A({ S25957[879] }),
  .ZN({ S2899 })
);
INV_X1 #() 
INV_X1_1698_ (
  .A({ S25957[774] }),
  .ZN({ S2900 })
);
AND2_X1 #() 
AND2_X1_325_ (
  .A1({ S1341 }),
  .A2({ S1343 }),
  .ZN({ S2901 })
);
NAND2_X1 #() 
NAND2_X1_5198_ (
  .A1({ S2891 }),
  .A2({ S2892 }),
  .ZN({ S2902 })
);
AOI21_X1 #() 
AOI21_X1_2920_ (
  .A({ S25957[898] }),
  .B1({ S1619 }),
  .B2({ S1620 }),
  .ZN({ S2903 })
);
AND3_X1 #() 
AND3_X1_220_ (
  .A1({ S1620 }),
  .A2({ S1619 }),
  .A3({ S25957[898] }),
  .ZN({ S2904 })
);
OAI21_X1 #() 
OAI21_X1_2696_ (
  .A({ S2902 }),
  .B1({ S2904 }),
  .B2({ S2903 }),
  .ZN({ S2905 })
);
NAND2_X1 #() 
NAND2_X1_5199_ (
  .A1({ S2905 }),
  .A2({ S25957[771] }),
  .ZN({ S2906 })
);
NOR2_X1 #() 
NOR2_X1_1316_ (
  .A1({ S2906 }),
  .A2({ S111 }),
  .ZN({ S2907 })
);
AOI21_X1 #() 
AOI21_X1_2921_ (
  .A({ S25957[771] }),
  .B1({ S25957[769] }),
  .B2({ S2898 }),
  .ZN({ S2908 })
);
NOR3_X1 #() 
NOR3_X1_167_ (
  .A1({ S2907 }),
  .A2({ S2908 }),
  .A3({ S2901 }),
  .ZN({ S2909 })
);
OAI21_X1 #() 
OAI21_X1_2697_ (
  .A({ S2898 }),
  .B1({ S2904 }),
  .B2({ S2903 }),
  .ZN({ S2910 })
);
NOR2_X1 #() 
NOR2_X1_1317_ (
  .A1({ S2904 }),
  .A2({ S2903 }),
  .ZN({ S2911 })
);
NAND3_X1 #() 
NAND3_X1_5586_ (
  .A1({ S25957[768] }),
  .A2({ S1557 }),
  .A3({ S1560 }),
  .ZN({ S2912 })
);
INV_X1 #() 
INV_X1_1699_ (
  .A({ S2912 }),
  .ZN({ S2913 })
);
NAND2_X1 #() 
NAND2_X1_5200_ (
  .A1({ S2911 }),
  .A2({ S2913 }),
  .ZN({ S2914 })
);
NAND3_X1 #() 
NAND3_X1_5587_ (
  .A1({ S2914 }),
  .A2({ S25957[771] }),
  .A3({ S2910 }),
  .ZN({ S2915 })
);
NAND3_X1 #() 
NAND3_X1_5588_ (
  .A1({ S1618 }),
  .A2({ S2898 }),
  .A3({ S1621 }),
  .ZN({ S2916 })
);
NOR2_X1 #() 
NOR2_X1_1318_ (
  .A1({ S25957[771] }),
  .A2({ S2902 }),
  .ZN({ S2917 })
);
NAND2_X1 #() 
NAND2_X1_5201_ (
  .A1({ S2917 }),
  .A2({ S2916 }),
  .ZN({ S2918 })
);
AOI21_X1 #() 
AOI21_X1_2922_ (
  .A({ S2901 }),
  .B1({ S2915 }),
  .B2({ S2918 }),
  .ZN({ S2919 })
);
OAI211_X1 #() 
OAI211_X1_1838_ (
  .A({ S2898 }),
  .B({ S2902 }),
  .C1({ S2904 }),
  .C2({ S2903 }),
  .ZN({ S2920 })
);
NAND4_X1 #() 
NAND4_X1_607_ (
  .A1({ S1618 }),
  .A2({ S25957[769] }),
  .A3({ S25957[768] }),
  .A4({ S1621 }),
  .ZN({ S2921 })
);
NAND3_X1 #() 
NAND3_X1_5589_ (
  .A1({ S2920 }),
  .A2({ S2921 }),
  .A3({ S104 }),
  .ZN({ S2922 })
);
OAI211_X1 #() 
OAI211_X1_1839_ (
  .A({ S2898 }),
  .B({ S25957[769] }),
  .C1({ S2904 }),
  .C2({ S2903 }),
  .ZN({ S2923 })
);
NAND3_X1 #() 
NAND3_X1_5590_ (
  .A1({ S2923 }),
  .A2({ S25957[771] }),
  .A3({ S2912 }),
  .ZN({ S2924 })
);
AND3_X1 #() 
AND3_X1_221_ (
  .A1({ S2922 }),
  .A2({ S2924 }),
  .A3({ S2901 }),
  .ZN({ S2925 })
);
OAI21_X1 #() 
OAI21_X1_2698_ (
  .A({ S25957[773] }),
  .B1({ S2925 }),
  .B2({ S2919 }),
  .ZN({ S2926 })
);
INV_X1 #() 
INV_X1_1700_ (
  .A({ S25957[773] }),
  .ZN({ S2927 })
);
NAND3_X1 #() 
NAND3_X1_5591_ (
  .A1({ S112 }),
  .A2({ S1618 }),
  .A3({ S1621 }),
  .ZN({ S2928 })
);
AOI21_X1 #() 
AOI21_X1_2923_ (
  .A({ S104 }),
  .B1({ S2891 }),
  .B2({ S2892 }),
  .ZN({ S2929 })
);
AOI22_X1 #() 
AOI22_X1_590_ (
  .A1({ S2920 }),
  .A2({ S2928 }),
  .B1({ S25957[768] }),
  .B2({ S2929 }),
  .ZN({ S2930 })
);
OAI21_X1 #() 
OAI21_X1_2699_ (
  .A({ S2927 }),
  .B1({ S2930 }),
  .B2({ S25957[772] }),
  .ZN({ S2931 })
);
OAI21_X1 #() 
OAI21_X1_2700_ (
  .A({ S2926 }),
  .B1({ S2909 }),
  .B2({ S2931 }),
  .ZN({ S2932 })
);
OAI21_X1 #() 
OAI21_X1_2701_ (
  .A({ S25957[769] }),
  .B1({ S2904 }),
  .B2({ S2903 }),
  .ZN({ S2933 })
);
INV_X1 #() 
INV_X1_1701_ (
  .A({ S2933 }),
  .ZN({ S2934 })
);
NAND4_X1 #() 
NAND4_X1_608_ (
  .A1({ S2893 }),
  .A2({ S112 }),
  .A3({ S1618 }),
  .A4({ S1621 }),
  .ZN({ S2935 })
);
NAND3_X1 #() 
NAND3_X1_5592_ (
  .A1({ S2898 }),
  .A2({ S2891 }),
  .A3({ S2892 }),
  .ZN({ S2936 })
);
OAI211_X1 #() 
OAI211_X1_1840_ (
  .A({ S2912 }),
  .B({ S2936 }),
  .C1({ S2904 }),
  .C2({ S2903 }),
  .ZN({ S2937 })
);
NAND3_X1 #() 
NAND3_X1_5593_ (
  .A1({ S2937 }),
  .A2({ S2935 }),
  .A3({ S25957[771] }),
  .ZN({ S2938 })
);
NAND3_X1 #() 
NAND3_X1_5594_ (
  .A1({ S1618 }),
  .A2({ S25957[768] }),
  .A3({ S1621 }),
  .ZN({ S2939 })
);
NAND2_X1 #() 
NAND2_X1_5202_ (
  .A1({ S2939 }),
  .A2({ S104 }),
  .ZN({ S2940 })
);
OAI21_X1 #() 
OAI21_X1_2702_ (
  .A({ S2938 }),
  .B1({ S2934 }),
  .B2({ S2940 }),
  .ZN({ S2941 })
);
NAND2_X1 #() 
NAND2_X1_5203_ (
  .A1({ S2941 }),
  .A2({ S25957[772] }),
  .ZN({ S2942 })
);
NAND2_X1 #() 
NAND2_X1_5204_ (
  .A1({ S2910 }),
  .A2({ S104 }),
  .ZN({ S2943 })
);
NAND2_X1 #() 
NAND2_X1_5205_ (
  .A1({ S2935 }),
  .A2({ S2933 }),
  .ZN({ S2944 })
);
AOI21_X1 #() 
AOI21_X1_2924_ (
  .A({ S25957[772] }),
  .B1({ S2911 }),
  .B2({ S2929 }),
  .ZN({ S2945 })
);
OAI21_X1 #() 
OAI21_X1_2703_ (
  .A({ S2945 }),
  .B1({ S2944 }),
  .B2({ S2943 }),
  .ZN({ S2946 })
);
AOI21_X1 #() 
AOI21_X1_2925_ (
  .A({ S25957[773] }),
  .B1({ S2942 }),
  .B2({ S2946 }),
  .ZN({ S2947 })
);
OAI21_X1 #() 
OAI21_X1_2704_ (
  .A({ S25957[768] }),
  .B1({ S2904 }),
  .B2({ S2903 }),
  .ZN({ S2948 })
);
INV_X1 #() 
INV_X1_1702_ (
  .A({ S2948 }),
  .ZN({ S2949 })
);
INV_X1 #() 
INV_X1_1703_ (
  .A({ S2917 }),
  .ZN({ S2950 })
);
NAND3_X1 #() 
NAND3_X1_5595_ (
  .A1({ S25957[770] }),
  .A2({ S25957[771] }),
  .A3({ S25957[768] }),
  .ZN({ S2951 })
);
INV_X1 #() 
INV_X1_1704_ (
  .A({ S2929 }),
  .ZN({ S2952 })
);
AND3_X1 #() 
AND3_X1_222_ (
  .A1({ S2951 }),
  .A2({ S25957[772] }),
  .A3({ S2952 }),
  .ZN({ S2953 })
);
OAI21_X1 #() 
OAI21_X1_2705_ (
  .A({ S2953 }),
  .B1({ S2949 }),
  .B2({ S2950 }),
  .ZN({ S2954 })
);
NAND4_X1 #() 
NAND4_X1_609_ (
  .A1({ S1618 }),
  .A2({ S2902 }),
  .A3({ S2898 }),
  .A4({ S1621 }),
  .ZN({ S2955 })
);
NAND2_X1 #() 
NAND2_X1_5206_ (
  .A1({ S2955 }),
  .A2({ S104 }),
  .ZN({ S2956 })
);
NAND3_X1 #() 
NAND3_X1_5596_ (
  .A1({ S2956 }),
  .A2({ S2901 }),
  .A3({ S2893 }),
  .ZN({ S2957 })
);
NAND3_X1 #() 
NAND3_X1_5597_ (
  .A1({ S2954 }),
  .A2({ S25957[773] }),
  .A3({ S2957 }),
  .ZN({ S2958 })
);
NAND2_X1 #() 
NAND2_X1_5207_ (
  .A1({ S2958 }),
  .A2({ S2900 }),
  .ZN({ S2959 })
);
OAI22_X1 #() 
OAI22_X1_133_ (
  .A1({ S2932 }),
  .A2({ S2900 }),
  .B1({ S2947 }),
  .B2({ S2959 }),
  .ZN({ S2960 })
);
NAND2_X1 #() 
NAND2_X1_5208_ (
  .A1({ S2960 }),
  .A2({ S25957[775] }),
  .ZN({ S2961 })
);
XNOR2_X1 #() 
XNOR2_X1_201_ (
  .A({ S1141 }),
  .B({ S24137 }),
  .ZN({ S2962 })
);
NAND2_X1 #() 
NAND2_X1_5209_ (
  .A1({ S2914 }),
  .A2({ S2933 }),
  .ZN({ S2963 })
);
NAND2_X1 #() 
NAND2_X1_5210_ (
  .A1({ S2963 }),
  .A2({ S25957[771] }),
  .ZN({ S2964 })
);
OAI21_X1 #() 
OAI21_X1_2706_ (
  .A({ S2893 }),
  .B1({ S2904 }),
  .B2({ S2903 }),
  .ZN({ S2965 })
);
NAND2_X1 #() 
NAND2_X1_5211_ (
  .A1({ S2965 }),
  .A2({ S104 }),
  .ZN({ S2966 })
);
NAND3_X1 #() 
NAND3_X1_5598_ (
  .A1({ S2964 }),
  .A2({ S2901 }),
  .A3({ S2966 }),
  .ZN({ S2967 })
);
NAND2_X1 #() 
NAND2_X1_5212_ (
  .A1({ S2916 }),
  .A2({ S2912 }),
  .ZN({ S2968 })
);
AOI21_X1 #() 
AOI21_X1_2926_ (
  .A({ S2936 }),
  .B1({ S1621 }),
  .B2({ S1618 }),
  .ZN({ S2969 })
);
NAND2_X1 #() 
NAND2_X1_5213_ (
  .A1({ S2916 }),
  .A2({ S104 }),
  .ZN({ S2970 })
);
NOR2_X1 #() 
NOR2_X1_1319_ (
  .A1({ S2970 }),
  .A2({ S2969 }),
  .ZN({ S2971 })
);
NAND3_X1 #() 
NAND3_X1_5599_ (
  .A1({ S25957[770] }),
  .A2({ S25957[771] }),
  .A3({ S25957[769] }),
  .ZN({ S2972 })
);
NAND2_X1 #() 
NAND2_X1_5214_ (
  .A1({ S2972 }),
  .A2({ S25957[772] }),
  .ZN({ S2973 })
);
AOI211_X1 #() 
AOI211_X1_88_ (
  .A({ S2973 }),
  .B({ S2971 }),
  .C1({ S2968 }),
  .C2({ S25957[771] }),
  .ZN({ S2974 })
);
NOR2_X1 #() 
NOR2_X1_1320_ (
  .A1({ S2974 }),
  .A2({ S2927 }),
  .ZN({ S2975 })
);
NAND3_X1 #() 
NAND3_X1_5600_ (
  .A1({ S1618 }),
  .A2({ S25957[769] }),
  .A3({ S1621 }),
  .ZN({ S2976 })
);
NAND3_X1 #() 
NAND3_X1_5601_ (
  .A1({ S2948 }),
  .A2({ S2976 }),
  .A3({ S25957[771] }),
  .ZN({ S2977 })
);
NAND3_X1 #() 
NAND3_X1_5602_ (
  .A1({ S2912 }),
  .A2({ S1618 }),
  .A3({ S1621 }),
  .ZN({ S2978 })
);
NAND2_X1 #() 
NAND2_X1_5215_ (
  .A1({ S2965 }),
  .A2({ S2978 }),
  .ZN({ S2979 })
);
AOI21_X1 #() 
AOI21_X1_2927_ (
  .A({ S25957[772] }),
  .B1({ S2979 }),
  .B2({ S104 }),
  .ZN({ S2980 })
);
NAND4_X1 #() 
NAND4_X1_610_ (
  .A1({ S2912 }),
  .A2({ S2936 }),
  .A3({ S1618 }),
  .A4({ S1621 }),
  .ZN({ S2981 })
);
AOI21_X1 #() 
AOI21_X1_2928_ (
  .A({ S104 }),
  .B1({ S2981 }),
  .B2({ S2965 }),
  .ZN({ S2982 })
);
AOI21_X1 #() 
AOI21_X1_2929_ (
  .A({ S25957[771] }),
  .B1({ S2937 }),
  .B2({ S2916 }),
  .ZN({ S2983 })
);
NOR3_X1 #() 
NOR3_X1_168_ (
  .A1({ S2983 }),
  .A2({ S2982 }),
  .A3({ S2901 }),
  .ZN({ S2984 })
);
AOI21_X1 #() 
AOI21_X1_2930_ (
  .A({ S2984 }),
  .B1({ S2980 }),
  .B2({ S2977 }),
  .ZN({ S2985 })
);
INV_X1 #() 
INV_X1_1705_ (
  .A({ S2985 }),
  .ZN({ S2986 })
);
AOI22_X1 #() 
AOI22_X1_591_ (
  .A1({ S2986 }),
  .A2({ S2927 }),
  .B1({ S2967 }),
  .B2({ S2975 }),
  .ZN({ S2987 })
);
NAND2_X1 #() 
NAND2_X1_5216_ (
  .A1({ S2910 }),
  .A2({ S25957[771] }),
  .ZN({ S2988 })
);
NAND2_X1 #() 
NAND2_X1_5217_ (
  .A1({ S2921 }),
  .A2({ S104 }),
  .ZN({ S2989 })
);
INV_X1 #() 
INV_X1_1706_ (
  .A({ S2989 }),
  .ZN({ S2990 })
);
OAI211_X1 #() 
OAI211_X1_1841_ (
  .A({ S2893 }),
  .B({ S112 }),
  .C1({ S2904 }),
  .C2({ S2903 }),
  .ZN({ S2991 })
);
AOI21_X1 #() 
AOI21_X1_2931_ (
  .A({ S2901 }),
  .B1({ S2990 }),
  .B2({ S2991 }),
  .ZN({ S2992 })
);
NAND3_X1 #() 
NAND3_X1_5603_ (
  .A1({ S2992 }),
  .A2({ S2988 }),
  .A3({ S2952 }),
  .ZN({ S2993 })
);
AOI22_X1 #() 
AOI22_X1_592_ (
  .A1({ S1618 }),
  .A2({ S1621 }),
  .B1({ S25957[769] }),
  .B2({ S2898 }),
  .ZN({ S2994 })
);
AOI21_X1 #() 
AOI21_X1_2932_ (
  .A({ S25957[771] }),
  .B1({ S2902 }),
  .B2({ S25957[768] }),
  .ZN({ S2995 })
);
NAND2_X1 #() 
NAND2_X1_5218_ (
  .A1({ S2994 }),
  .A2({ S2995 }),
  .ZN({ S2996 })
);
OAI211_X1 #() 
OAI211_X1_1842_ (
  .A({ S2996 }),
  .B({ S2901 }),
  .C1({ S104 }),
  .C2({ S2965 }),
  .ZN({ S2997 })
);
NAND3_X1 #() 
NAND3_X1_5604_ (
  .A1({ S2993 }),
  .A2({ S2927 }),
  .A3({ S2997 }),
  .ZN({ S2998 })
);
NAND3_X1 #() 
NAND3_X1_5605_ (
  .A1({ S2893 }),
  .A2({ S1618 }),
  .A3({ S1621 }),
  .ZN({ S2999 })
);
INV_X1 #() 
INV_X1_1707_ (
  .A({ S2999 }),
  .ZN({ S3000 })
);
AOI21_X1 #() 
AOI21_X1_2933_ (
  .A({ S25957[771] }),
  .B1({ S25957[770] }),
  .B2({ S25957[769] }),
  .ZN({ S3001 })
);
INV_X1 #() 
INV_X1_1708_ (
  .A({ S3001 }),
  .ZN({ S3002 })
);
NAND3_X1 #() 
NAND3_X1_5606_ (
  .A1({ S2976 }),
  .A2({ S25957[771] }),
  .A3({ S2912 }),
  .ZN({ S3003 })
);
OAI211_X1 #() 
OAI211_X1_1843_ (
  .A({ S2901 }),
  .B({ S3003 }),
  .C1({ S3002 }),
  .C2({ S3000 }),
  .ZN({ S3004 })
);
NAND2_X1 #() 
NAND2_X1_5219_ (
  .A1({ S104 }),
  .A2({ S25957[768] }),
  .ZN({ S3005 })
);
NAND3_X1 #() 
NAND3_X1_5607_ (
  .A1({ S1618 }),
  .A2({ S2902 }),
  .A3({ S1621 }),
  .ZN({ S3006 })
);
NAND3_X1 #() 
NAND3_X1_5608_ (
  .A1({ S2948 }),
  .A2({ S3006 }),
  .A3({ S25957[771] }),
  .ZN({ S3007 })
);
AND2_X1 #() 
AND2_X1_326_ (
  .A1({ S3007 }),
  .A2({ S3005 }),
  .ZN({ S3008 })
);
OAI21_X1 #() 
OAI21_X1_2707_ (
  .A({ S3004 }),
  .B1({ S2901 }),
  .B2({ S3008 }),
  .ZN({ S3009 })
);
AOI21_X1 #() 
AOI21_X1_2934_ (
  .A({ S25957[774] }),
  .B1({ S3009 }),
  .B2({ S25957[773] }),
  .ZN({ S3010 })
);
AOI22_X1 #() 
AOI22_X1_593_ (
  .A1({ S2987 }),
  .A2({ S25957[774] }),
  .B1({ S2998 }),
  .B2({ S3010 }),
  .ZN({ S3011 })
);
NAND2_X1 #() 
NAND2_X1_5220_ (
  .A1({ S3011 }),
  .A2({ S2962 }),
  .ZN({ S3012 })
);
NAND2_X1 #() 
NAND2_X1_5221_ (
  .A1({ S3012 }),
  .A2({ S2961 }),
  .ZN({ S3013 })
);
NAND2_X1 #() 
NAND2_X1_5222_ (
  .A1({ S3013 }),
  .A2({ S2899 }),
  .ZN({ S3014 })
);
NAND3_X1 #() 
NAND3_X1_5609_ (
  .A1({ S3012 }),
  .A2({ S25957[879] }),
  .A3({ S2961 }),
  .ZN({ S3015 })
);
NAND2_X1 #() 
NAND2_X1_5223_ (
  .A1({ S3014 }),
  .A2({ S3015 }),
  .ZN({ S25957[751] })
);
NAND2_X1 #() 
NAND2_X1_5224_ (
  .A1({ S25957[751] }),
  .A2({ S474 }),
  .ZN({ S3016 })
);
NAND3_X1 #() 
NAND3_X1_5610_ (
  .A1({ S3014 }),
  .A2({ S25957[847] }),
  .A3({ S3015 }),
  .ZN({ S3017 })
);
NAND2_X1 #() 
NAND2_X1_5225_ (
  .A1({ S3016 }),
  .A2({ S3017 }),
  .ZN({ S25957[719] })
);
NAND2_X1 #() 
NAND2_X1_5226_ (
  .A1({ S25957[719] }),
  .A2({ S25957[911] }),
  .ZN({ S3018 })
);
NAND3_X1 #() 
NAND3_X1_5611_ (
  .A1({ S3016 }),
  .A2({ S3017 }),
  .A3({ S25568 }),
  .ZN({ S3019 })
);
NAND2_X1 #() 
NAND2_X1_5227_ (
  .A1({ S3018 }),
  .A2({ S3019 }),
  .ZN({ S3020 })
);
INV_X1 #() 
INV_X1_1709_ (
  .A({ S3020 }),
  .ZN({ S25957[655] })
);
INV_X1 #() 
INV_X1_1710_ (
  .A({ S2939 }),
  .ZN({ S3021 })
);
NOR2_X1 #() 
NOR2_X1_1321_ (
  .A1({ S2911 }),
  .A2({ S2913 }),
  .ZN({ S3022 })
);
OAI21_X1 #() 
OAI21_X1_2708_ (
  .A({ S25957[771] }),
  .B1({ S3022 }),
  .B2({ S3021 }),
  .ZN({ S3023 })
);
INV_X1 #() 
INV_X1_1711_ (
  .A({ S2935 }),
  .ZN({ S3024 })
);
OAI21_X1 #() 
OAI21_X1_2709_ (
  .A({ S104 }),
  .B1({ S3024 }),
  .B2({ S2949 }),
  .ZN({ S3025 })
);
AND2_X1 #() 
AND2_X1_327_ (
  .A1({ S3025 }),
  .A2({ S3023 }),
  .ZN({ S3026 })
);
INV_X1 #() 
INV_X1_1712_ (
  .A({ S3005 }),
  .ZN({ S3027 })
);
NAND3_X1 #() 
NAND3_X1_5612_ (
  .A1({ S2905 }),
  .A2({ S2976 }),
  .A3({ S3027 }),
  .ZN({ S3028 })
);
INV_X1 #() 
INV_X1_1713_ (
  .A({ S3028 }),
  .ZN({ S3029 })
);
AOI21_X1 #() 
AOI21_X1_2935_ (
  .A({ S25957[768] }),
  .B1({ S1618 }),
  .B2({ S1621 }),
  .ZN({ S3030 })
);
NAND2_X1 #() 
NAND2_X1_5228_ (
  .A1({ S3030 }),
  .A2({ S2929 }),
  .ZN({ S3031 })
);
OAI211_X1 #() 
OAI211_X1_1844_ (
  .A({ S3031 }),
  .B({ S2901 }),
  .C1({ S104 }),
  .C2({ S2999 }),
  .ZN({ S3032 })
);
OAI221_X1 #() 
OAI221_X1_155_ (
  .A({ S2927 }),
  .B1({ S3029 }),
  .B2({ S3032 }),
  .C1({ S3026 }),
  .C2({ S2901 }),
  .ZN({ S3033 })
);
OAI21_X1 #() 
OAI21_X1_2710_ (
  .A({ S112 }),
  .B1({ S2904 }),
  .B2({ S2903 }),
  .ZN({ S3034 })
);
NAND4_X1 #() 
NAND4_X1_611_ (
  .A1({ S2910 }),
  .A2({ S2939 }),
  .A3({ S25957[771] }),
  .A4({ S2902 }),
  .ZN({ S3035 })
);
OAI21_X1 #() 
OAI21_X1_2711_ (
  .A({ S3035 }),
  .B1({ S25957[771] }),
  .B2({ S3034 }),
  .ZN({ S3036 })
);
NOR2_X1 #() 
NOR2_X1_1322_ (
  .A1({ S2907 }),
  .A2({ S2917 }),
  .ZN({ S3037 })
);
MUX2_X1 #() 
MUX2_X1_21_ (
  .A({ S3036 }),
  .B({ S3037 }),
  .S({ S2901 }),
  .Z({ S3038 })
);
AOI21_X1 #() 
AOI21_X1_2936_ (
  .A({ S2900 }),
  .B1({ S3038 }),
  .B2({ S25957[773] }),
  .ZN({ S3039 })
);
NAND4_X1 #() 
NAND4_X1_612_ (
  .A1({ S2921 }),
  .A2({ S2933 }),
  .A3({ S3006 }),
  .A4({ S25957[771] }),
  .ZN({ S3040 })
);
OAI211_X1 #() 
OAI211_X1_1845_ (
  .A({ S25957[768] }),
  .B({ S25957[769] }),
  .C1({ S2904 }),
  .C2({ S2903 }),
  .ZN({ S3041 })
);
NAND3_X1 #() 
NAND3_X1_5613_ (
  .A1({ S3041 }),
  .A2({ S104 }),
  .A3({ S112 }),
  .ZN({ S3042 })
);
NAND3_X1 #() 
NAND3_X1_5614_ (
  .A1({ S3040 }),
  .A2({ S2901 }),
  .A3({ S3042 }),
  .ZN({ S3043 })
);
NAND4_X1 #() 
NAND4_X1_613_ (
  .A1({ S1618 }),
  .A2({ S25957[769] }),
  .A3({ S2898 }),
  .A4({ S1621 }),
  .ZN({ S3044 })
);
AOI21_X1 #() 
AOI21_X1_2937_ (
  .A({ S25957[771] }),
  .B1({ S2937 }),
  .B2({ S3044 }),
  .ZN({ S3045 })
);
OAI211_X1 #() 
OAI211_X1_1846_ (
  .A({ S3043 }),
  .B({ S25957[773] }),
  .C1({ S2973 }),
  .C2({ S3045 }),
  .ZN({ S3046 })
);
OAI21_X1 #() 
OAI21_X1_2712_ (
  .A({ S2936 }),
  .B1({ S2904 }),
  .B2({ S2903 }),
  .ZN({ S3047 })
);
NAND3_X1 #() 
NAND3_X1_5615_ (
  .A1({ S3047 }),
  .A2({ S25957[771] }),
  .A3({ S2916 }),
  .ZN({ S3048 })
);
AOI21_X1 #() 
AOI21_X1_2938_ (
  .A({ S25957[772] }),
  .B1({ S3025 }),
  .B2({ S3048 }),
  .ZN({ S3049 })
);
INV_X1 #() 
INV_X1_1714_ (
  .A({ S2978 }),
  .ZN({ S3050 })
);
NAND2_X1 #() 
NAND2_X1_5229_ (
  .A1({ S3050 }),
  .A2({ S104 }),
  .ZN({ S3051 })
);
AOI21_X1 #() 
AOI21_X1_2939_ (
  .A({ S3049 }),
  .B1({ S2953 }),
  .B2({ S3051 }),
  .ZN({ S3052 })
);
OAI21_X1 #() 
OAI21_X1_2713_ (
  .A({ S3046 }),
  .B1({ S3052 }),
  .B2({ S25957[773] }),
  .ZN({ S3053 })
);
AOI22_X1 #() 
AOI22_X1_594_ (
  .A1({ S3053 }),
  .A2({ S2900 }),
  .B1({ S3039 }),
  .B2({ S3033 }),
  .ZN({ S3054 })
);
INV_X1 #() 
INV_X1_1715_ (
  .A({ S2940 }),
  .ZN({ S3055 })
);
NAND2_X1 #() 
NAND2_X1_5230_ (
  .A1({ S2948 }),
  .A2({ S2936 }),
  .ZN({ S3056 })
);
AOI22_X1 #() 
AOI22_X1_595_ (
  .A1({ S3055 }),
  .A2({ S2965 }),
  .B1({ S3056 }),
  .B2({ S25957[771] }),
  .ZN({ S3057 })
);
NAND2_X1 #() 
NAND2_X1_5231_ (
  .A1({ S2939 }),
  .A2({ S112 }),
  .ZN({ S3058 })
);
NOR2_X1 #() 
NOR2_X1_1323_ (
  .A1({ S25957[771] }),
  .A2({ S25957[769] }),
  .ZN({ S3059 })
);
OAI21_X1 #() 
OAI21_X1_2714_ (
  .A({ S2901 }),
  .B1({ S3058 }),
  .B2({ S3059 }),
  .ZN({ S3060 })
);
OAI211_X1 #() 
OAI211_X1_1847_ (
  .A({ S3060 }),
  .B({ S25957[773] }),
  .C1({ S3057 }),
  .C2({ S2901 }),
  .ZN({ S3061 })
);
NAND2_X1 #() 
NAND2_X1_5232_ (
  .A1({ S2991 }),
  .A2({ S104 }),
  .ZN({ S3062 })
);
NAND3_X1 #() 
NAND3_X1_5616_ (
  .A1({ S3023 }),
  .A2({ S2901 }),
  .A3({ S3062 }),
  .ZN({ S3063 })
);
NAND2_X1 #() 
NAND2_X1_5233_ (
  .A1({ S2910 }),
  .A2({ S2936 }),
  .ZN({ S3064 })
);
NAND2_X1 #() 
NAND2_X1_5234_ (
  .A1({ S3064 }),
  .A2({ S104 }),
  .ZN({ S3065 })
);
NAND4_X1 #() 
NAND4_X1_614_ (
  .A1({ S25957[771] }),
  .A2({ S1618 }),
  .A3({ S25957[769] }),
  .A4({ S1621 }),
  .ZN({ S3066 })
);
NAND3_X1 #() 
NAND3_X1_5617_ (
  .A1({ S3065 }),
  .A2({ S25957[772] }),
  .A3({ S3066 }),
  .ZN({ S3067 })
);
NAND3_X1 #() 
NAND3_X1_5618_ (
  .A1({ S3063 }),
  .A2({ S2927 }),
  .A3({ S3067 }),
  .ZN({ S3068 })
);
AOI21_X1 #() 
AOI21_X1_2940_ (
  .A({ S2900 }),
  .B1({ S3068 }),
  .B2({ S3061 }),
  .ZN({ S3069 })
);
INV_X1 #() 
INV_X1_1716_ (
  .A({ S2976 }),
  .ZN({ S3070 })
);
NAND2_X1 #() 
NAND2_X1_5235_ (
  .A1({ S3001 }),
  .A2({ S2914 }),
  .ZN({ S3071 })
);
OAI21_X1 #() 
OAI21_X1_2715_ (
  .A({ S3071 }),
  .B1({ S3070 }),
  .B2({ S2906 }),
  .ZN({ S3072 })
);
NAND3_X1 #() 
NAND3_X1_5619_ (
  .A1({ S2920 }),
  .A2({ S25957[771] }),
  .A3({ S2893 }),
  .ZN({ S3073 })
);
NAND3_X1 #() 
NAND3_X1_5620_ (
  .A1({ S3073 }),
  .A2({ S25957[772] }),
  .A3({ S2940 }),
  .ZN({ S3074 })
);
OAI211_X1 #() 
OAI211_X1_1848_ (
  .A({ S25957[773] }),
  .B({ S3074 }),
  .C1({ S3072 }),
  .C2({ S25957[772] }),
  .ZN({ S3075 })
);
AND4_X1 #() 
AND4_X1_12_ (
  .A1({ S25957[772] }),
  .A2({ S2964 }),
  .A3({ S2950 }),
  .A4({ S2940 }),
  .ZN({ S3076 })
);
NAND3_X1 #() 
NAND3_X1_5621_ (
  .A1({ S2936 }),
  .A2({ S1618 }),
  .A3({ S1621 }),
  .ZN({ S3077 })
);
NAND2_X1 #() 
NAND2_X1_5236_ (
  .A1({ S2923 }),
  .A2({ S3077 }),
  .ZN({ S3078 })
);
NAND3_X1 #() 
NAND3_X1_5622_ (
  .A1({ S3078 }),
  .A2({ S2901 }),
  .A3({ S25957[771] }),
  .ZN({ S3079 })
);
INV_X1 #() 
INV_X1_1717_ (
  .A({ S3079 }),
  .ZN({ S3080 })
);
OAI21_X1 #() 
OAI21_X1_2716_ (
  .A({ S2927 }),
  .B1({ S3076 }),
  .B2({ S3080 }),
  .ZN({ S3081 })
);
NAND2_X1 #() 
NAND2_X1_5237_ (
  .A1({ S3081 }),
  .A2({ S3075 }),
  .ZN({ S3082 })
);
AOI21_X1 #() 
AOI21_X1_2941_ (
  .A({ S3069 }),
  .B1({ S2900 }),
  .B2({ S3082 }),
  .ZN({ S3083 })
);
MUX2_X1 #() 
MUX2_X1_22_ (
  .A({ S3083 }),
  .B({ S3054 }),
  .S({ S25957[775] }),
  .Z({ S3084 })
);
XNOR2_X1 #() 
XNOR2_X1_202_ (
  .A({ S3084 }),
  .B({ S20130 }),
  .ZN({ S25957[654] })
);
INV_X1 #() 
INV_X1_1718_ (
  .A({ S633 }),
  .ZN({ S25957[845] })
);
NOR2_X1 #() 
NOR2_X1_1324_ (
  .A1({ S23621 }),
  .A2({ S23620 }),
  .ZN({ S3085 })
);
XOR2_X1 #() 
XOR2_X1_86_ (
  .A({ S3085 }),
  .B({ S25957[1133] }),
  .Z({ S25957[1005] })
);
AND2_X1 #() 
AND2_X1_328_ (
  .A1({ S629 }),
  .A2({ S591 }),
  .ZN({ S3086 })
);
XNOR2_X1 #() 
XNOR2_X1_203_ (
  .A({ S3086 }),
  .B({ S25957[1005] }),
  .ZN({ S25957[877] })
);
NAND2_X1 #() 
NAND2_X1_5238_ (
  .A1({ S2908 }),
  .A2({ S2939 }),
  .ZN({ S3087 })
);
OAI21_X1 #() 
OAI21_X1_2717_ (
  .A({ S3087 }),
  .B1({ S104 }),
  .B2({ S25957[768] }),
  .ZN({ S3088 })
);
NAND2_X1 #() 
NAND2_X1_5239_ (
  .A1({ S3088 }),
  .A2({ S25957[773] }),
  .ZN({ S3089 })
);
NAND3_X1 #() 
NAND3_X1_5623_ (
  .A1({ S2965 }),
  .A2({ S25957[771] }),
  .A3({ S2939 }),
  .ZN({ S3090 })
);
INV_X1 #() 
INV_X1_1719_ (
  .A({ S3090 }),
  .ZN({ S3091 })
);
AOI21_X1 #() 
AOI21_X1_2942_ (
  .A({ S25957[771] }),
  .B1({ S3077 }),
  .B2({ S2910 }),
  .ZN({ S3092 })
);
OAI21_X1 #() 
OAI21_X1_2718_ (
  .A({ S2927 }),
  .B1({ S3091 }),
  .B2({ S3092 }),
  .ZN({ S3093 })
);
AOI21_X1 #() 
AOI21_X1_2943_ (
  .A({ S25957[772] }),
  .B1({ S3093 }),
  .B2({ S3089 }),
  .ZN({ S3094 })
);
NAND2_X1 #() 
NAND2_X1_5240_ (
  .A1({ S3050 }),
  .A2({ S25957[771] }),
  .ZN({ S3095 })
);
NAND3_X1 #() 
NAND3_X1_5624_ (
  .A1({ S3041 }),
  .A2({ S2999 }),
  .A3({ S104 }),
  .ZN({ S3096 })
);
NAND3_X1 #() 
NAND3_X1_5625_ (
  .A1({ S3095 }),
  .A2({ S2927 }),
  .A3({ S3096 }),
  .ZN({ S3097 })
);
INV_X1 #() 
INV_X1_1720_ (
  .A({ S2963 }),
  .ZN({ S3098 })
);
NAND3_X1 #() 
NAND3_X1_5626_ (
  .A1({ S2937 }),
  .A2({ S25957[771] }),
  .A3({ S3044 }),
  .ZN({ S3099 })
);
OAI211_X1 #() 
OAI211_X1_1849_ (
  .A({ S3099 }),
  .B({ S25957[773] }),
  .C1({ S25957[771] }),
  .C2({ S3098 }),
  .ZN({ S3100 })
);
AOI21_X1 #() 
AOI21_X1_2944_ (
  .A({ S2901 }),
  .B1({ S3100 }),
  .B2({ S3097 }),
  .ZN({ S3101 })
);
OAI21_X1 #() 
OAI21_X1_2719_ (
  .A({ S25957[774] }),
  .B1({ S3101 }),
  .B2({ S3094 }),
  .ZN({ S3102 })
);
NAND2_X1 #() 
NAND2_X1_5241_ (
  .A1({ S3044 }),
  .A2({ S104 }),
  .ZN({ S3103 })
);
OAI211_X1 #() 
OAI211_X1_1850_ (
  .A({ S3103 }),
  .B({ S25957[772] }),
  .C1({ S104 }),
  .C2({ S2999 }),
  .ZN({ S3104 })
);
NAND2_X1 #() 
NAND2_X1_5242_ (
  .A1({ S2939 }),
  .A2({ S25957[769] }),
  .ZN({ S3105 })
);
OAI211_X1 #() 
OAI211_X1_1851_ (
  .A({ S2951 }),
  .B({ S2901 }),
  .C1({ S2943 }),
  .C2({ S3105 }),
  .ZN({ S3106 })
);
AND3_X1 #() 
AND3_X1_223_ (
  .A1({ S3106 }),
  .A2({ S3104 }),
  .A3({ S25957[773] }),
  .ZN({ S3107 })
);
NAND3_X1 #() 
NAND3_X1_5627_ (
  .A1({ S2914 }),
  .A2({ S2937 }),
  .A3({ S25957[771] }),
  .ZN({ S3108 })
);
NAND3_X1 #() 
NAND3_X1_5628_ (
  .A1({ S2908 }),
  .A2({ S2916 }),
  .A3({ S2912 }),
  .ZN({ S3109 })
);
NAND3_X1 #() 
NAND3_X1_5629_ (
  .A1({ S3108 }),
  .A2({ S25957[772] }),
  .A3({ S3109 }),
  .ZN({ S3110 })
);
OAI22_X1 #() 
OAI22_X1_134_ (
  .A1({ S2898 }),
  .A2({ S2952 }),
  .B1({ S3041 }),
  .B2({ S25957[771] }),
  .ZN({ S3111 })
);
NAND2_X1 #() 
NAND2_X1_5243_ (
  .A1({ S3111 }),
  .A2({ S2901 }),
  .ZN({ S3112 })
);
AOI21_X1 #() 
AOI21_X1_2945_ (
  .A({ S25957[773] }),
  .B1({ S3110 }),
  .B2({ S3112 }),
  .ZN({ S3113 })
);
OAI21_X1 #() 
OAI21_X1_2720_ (
  .A({ S2900 }),
  .B1({ S3107 }),
  .B2({ S3113 }),
  .ZN({ S3114 })
);
AND2_X1 #() 
AND2_X1_329_ (
  .A1({ S3102 }),
  .A2({ S3114 }),
  .ZN({ S3115 })
);
NOR2_X1 #() 
NOR2_X1_1325_ (
  .A1({ S3115 }),
  .A2({ S25957[775] }),
  .ZN({ S3116 })
);
NAND3_X1 #() 
NAND3_X1_5630_ (
  .A1({ S3023 }),
  .A2({ S2901 }),
  .A3({ S2996 }),
  .ZN({ S3117 })
);
NAND2_X1 #() 
NAND2_X1_5244_ (
  .A1({ S3077 }),
  .A2({ S25957[771] }),
  .ZN({ S3118 })
);
NAND2_X1 #() 
NAND2_X1_5245_ (
  .A1({ S2994 }),
  .A2({ S104 }),
  .ZN({ S3119 })
);
NAND3_X1 #() 
NAND3_X1_5631_ (
  .A1({ S3119 }),
  .A2({ S25957[772] }),
  .A3({ S3118 }),
  .ZN({ S3120 })
);
NAND3_X1 #() 
NAND3_X1_5632_ (
  .A1({ S3117 }),
  .A2({ S2927 }),
  .A3({ S3120 }),
  .ZN({ S3121 })
);
OAI21_X1 #() 
OAI21_X1_2721_ (
  .A({ S25957[771] }),
  .B1({ S3000 }),
  .B2({ S2994 }),
  .ZN({ S3122 })
);
AOI22_X1 #() 
AOI22_X1_596_ (
  .A1({ S25957[770] }),
  .A2({ S3027 }),
  .B1({ S25957[769] }),
  .B2({ S104 }),
  .ZN({ S3123 })
);
NAND3_X1 #() 
NAND3_X1_5633_ (
  .A1({ S3122 }),
  .A2({ S2901 }),
  .A3({ S3123 }),
  .ZN({ S3124 })
);
OAI21_X1 #() 
OAI21_X1_2722_ (
  .A({ S104 }),
  .B1({ S3050 }),
  .B2({ S2969 }),
  .ZN({ S3125 })
);
OAI211_X1 #() 
OAI211_X1_1852_ (
  .A({ S3125 }),
  .B({ S25957[772] }),
  .C1({ S104 }),
  .C2({ S3064 }),
  .ZN({ S3126 })
);
NAND3_X1 #() 
NAND3_X1_5634_ (
  .A1({ S3126 }),
  .A2({ S25957[773] }),
  .A3({ S3124 }),
  .ZN({ S3127 })
);
NAND3_X1 #() 
NAND3_X1_5635_ (
  .A1({ S3127 }),
  .A2({ S3121 }),
  .A3({ S25957[774] }),
  .ZN({ S3128 })
);
AND2_X1 #() 
AND2_X1_330_ (
  .A1({ S2991 }),
  .A2({ S2955 }),
  .ZN({ S3129 })
);
OAI21_X1 #() 
OAI21_X1_2723_ (
  .A({ S2989 }),
  .B1({ S3129 }),
  .B2({ S104 }),
  .ZN({ S3130 })
);
NAND2_X1 #() 
NAND2_X1_5246_ (
  .A1({ S3024 }),
  .A2({ S25957[771] }),
  .ZN({ S3131 })
);
AOI21_X1 #() 
AOI21_X1_2946_ (
  .A({ S2901 }),
  .B1({ S2939 }),
  .B2({ S3059 }),
  .ZN({ S3132 })
);
AOI22_X1 #() 
AOI22_X1_597_ (
  .A1({ S3130 }),
  .A2({ S2901 }),
  .B1({ S3131 }),
  .B2({ S3132 }),
  .ZN({ S3133 })
);
OAI21_X1 #() 
OAI21_X1_2724_ (
  .A({ S104 }),
  .B1({ S3030 }),
  .B2({ S2913 }),
  .ZN({ S3134 })
);
OAI211_X1 #() 
OAI211_X1_1853_ (
  .A({ S3134 }),
  .B({ S25957[772] }),
  .C1({ S2979 }),
  .C2({ S104 }),
  .ZN({ S3135 })
);
NAND2_X1 #() 
NAND2_X1_5247_ (
  .A1({ S2908 }),
  .A2({ S3006 }),
  .ZN({ S3136 })
);
NAND3_X1 #() 
NAND3_X1_5636_ (
  .A1({ S3136 }),
  .A2({ S2901 }),
  .A3({ S2952 }),
  .ZN({ S3137 })
);
NAND3_X1 #() 
NAND3_X1_5637_ (
  .A1({ S3135 }),
  .A2({ S25957[773] }),
  .A3({ S3137 }),
  .ZN({ S3138 })
);
OAI211_X1 #() 
OAI211_X1_1854_ (
  .A({ S2900 }),
  .B({ S3138 }),
  .C1({ S3133 }),
  .C2({ S25957[773] }),
  .ZN({ S3139 })
);
NAND3_X1 #() 
NAND3_X1_5638_ (
  .A1({ S3139 }),
  .A2({ S25957[775] }),
  .A3({ S3128 }),
  .ZN({ S3140 })
);
INV_X1 #() 
INV_X1_1721_ (
  .A({ S3140 }),
  .ZN({ S3141 })
);
OAI21_X1 #() 
OAI21_X1_2725_ (
  .A({ S25957[877] }),
  .B1({ S3116 }),
  .B2({ S3141 }),
  .ZN({ S3142 })
);
INV_X1 #() 
INV_X1_1722_ (
  .A({ S25957[877] }),
  .ZN({ S3143 })
);
OAI211_X1 #() 
OAI211_X1_1855_ (
  .A({ S3140 }),
  .B({ S3143 }),
  .C1({ S3115 }),
  .C2({ S25957[775] }),
  .ZN({ S3144 })
);
NAND2_X1 #() 
NAND2_X1_5248_ (
  .A1({ S3142 }),
  .A2({ S3144 }),
  .ZN({ S25957[749] })
);
NAND2_X1 #() 
NAND2_X1_5249_ (
  .A1({ S25957[749] }),
  .A2({ S25957[845] }),
  .ZN({ S3145 })
);
NAND3_X1 #() 
NAND3_X1_5639_ (
  .A1({ S3142 }),
  .A2({ S633 }),
  .A3({ S3144 }),
  .ZN({ S3146 })
);
NAND3_X1 #() 
NAND3_X1_5640_ (
  .A1({ S3145 }),
  .A2({ S3146 }),
  .A3({ S25957[909] }),
  .ZN({ S3147 })
);
NAND3_X1 #() 
NAND3_X1_5641_ (
  .A1({ S3142 }),
  .A2({ S25957[845] }),
  .A3({ S3144 }),
  .ZN({ S3148 })
);
OAI21_X1 #() 
OAI21_X1_2726_ (
  .A({ S3143 }),
  .B1({ S3116 }),
  .B2({ S3141 }),
  .ZN({ S3149 })
);
OAI211_X1 #() 
OAI211_X1_1856_ (
  .A({ S3140 }),
  .B({ S25957[877] }),
  .C1({ S3115 }),
  .C2({ S25957[775] }),
  .ZN({ S3150 })
);
NAND3_X1 #() 
NAND3_X1_5642_ (
  .A1({ S3149 }),
  .A2({ S633 }),
  .A3({ S3150 }),
  .ZN({ S3151 })
);
NAND3_X1 #() 
NAND3_X1_5643_ (
  .A1({ S3148 }),
  .A2({ S3151 }),
  .A3({ S25484 }),
  .ZN({ S3152 })
);
AND2_X1 #() 
AND2_X1_331_ (
  .A1({ S3147 }),
  .A2({ S3152 }),
  .ZN({ S25957[653] })
);
NOR2_X1 #() 
NOR2_X1_1326_ (
  .A1({ S706 }),
  .A2({ S709 }),
  .ZN({ S25957[812] })
);
NOR2_X1 #() 
NOR2_X1_1327_ (
  .A1({ S23709 }),
  .A2({ S23712 }),
  .ZN({ S25957[972] })
);
INV_X1 #() 
INV_X1_1723_ (
  .A({ S2921 }),
  .ZN({ S3153 })
);
AOI21_X1 #() 
AOI21_X1_2947_ (
  .A({ S25957[772] }),
  .B1({ S25957[770] }),
  .B2({ S25957[771] }),
  .ZN({ S3154 })
);
OAI21_X1 #() 
OAI21_X1_2727_ (
  .A({ S3154 }),
  .B1({ S2943 }),
  .B2({ S3153 }),
  .ZN({ S3155 })
);
OAI221_X1 #() 
OAI221_X1_156_ (
  .A({ S2953 }),
  .B1({ S25957[770] }),
  .B2({ S2950 }),
  .C1({ S25957[771] }),
  .C2({ S2920 }),
  .ZN({ S3156 })
);
NAND3_X1 #() 
NAND3_X1_5644_ (
  .A1({ S3156 }),
  .A2({ S2927 }),
  .A3({ S3155 }),
  .ZN({ S3157 })
);
AND2_X1 #() 
AND2_X1_332_ (
  .A1({ S2911 }),
  .A2({ S133 }),
  .ZN({ S3158 })
);
AOI21_X1 #() 
AOI21_X1_2948_ (
  .A({ S25957[771] }),
  .B1({ S2935 }),
  .B2({ S3047 }),
  .ZN({ S3159 })
);
NAND2_X1 #() 
NAND2_X1_5250_ (
  .A1({ S3090 }),
  .A2({ S2901 }),
  .ZN({ S3160 })
);
OAI221_X1 #() 
OAI221_X1_157_ (
  .A({ S25957[773] }),
  .B1({ S3158 }),
  .B2({ S2901 }),
  .C1({ S3160 }),
  .C2({ S3159 }),
  .ZN({ S3161 })
);
NAND3_X1 #() 
NAND3_X1_5645_ (
  .A1({ S3157 }),
  .A2({ S2962 }),
  .A3({ S3161 }),
  .ZN({ S3162 })
);
NAND2_X1 #() 
NAND2_X1_5251_ (
  .A1({ S112 }),
  .A2({ S104 }),
  .ZN({ S3163 })
);
AND2_X1 #() 
AND2_X1_333_ (
  .A1({ S2978 }),
  .A2({ S3163 }),
  .ZN({ S3164 })
);
NAND2_X1 #() 
NAND2_X1_5252_ (
  .A1({ S3164 }),
  .A2({ S25957[772] }),
  .ZN({ S3165 })
);
NAND3_X1 #() 
NAND3_X1_5646_ (
  .A1({ S2976 }),
  .A2({ S104 }),
  .A3({ S2898 }),
  .ZN({ S3166 })
);
NAND3_X1 #() 
NAND3_X1_5647_ (
  .A1({ S3007 }),
  .A2({ S3166 }),
  .A3({ S2901 }),
  .ZN({ S3167 })
);
NAND3_X1 #() 
NAND3_X1_5648_ (
  .A1({ S3165 }),
  .A2({ S3167 }),
  .A3({ S25957[773] }),
  .ZN({ S3168 })
);
NAND3_X1 #() 
NAND3_X1_5649_ (
  .A1({ S2910 }),
  .A2({ S3006 }),
  .A3({ S104 }),
  .ZN({ S3169 })
);
NAND3_X1 #() 
NAND3_X1_5650_ (
  .A1({ S3169 }),
  .A2({ S3003 }),
  .A3({ S2901 }),
  .ZN({ S3170 })
);
OAI21_X1 #() 
OAI21_X1_2728_ (
  .A({ S3136 }),
  .B1({ S3021 }),
  .B2({ S2952 }),
  .ZN({ S3171 })
);
OAI211_X1 #() 
OAI211_X1_1857_ (
  .A({ S3170 }),
  .B({ S2927 }),
  .C1({ S3171 }),
  .C2({ S2901 }),
  .ZN({ S3172 })
);
NAND3_X1 #() 
NAND3_X1_5651_ (
  .A1({ S25957[775] }),
  .A2({ S3168 }),
  .A3({ S3172 }),
  .ZN({ S3173 })
);
NAND2_X1 #() 
NAND2_X1_5253_ (
  .A1({ S3162 }),
  .A2({ S3173 }),
  .ZN({ S3174 })
);
NAND2_X1 #() 
NAND2_X1_5254_ (
  .A1({ S3174 }),
  .A2({ S25957[774] }),
  .ZN({ S3175 })
);
AOI21_X1 #() 
AOI21_X1_2949_ (
  .A({ S25957[771] }),
  .B1({ S2981 }),
  .B2({ S2965 }),
  .ZN({ S3176 })
);
NAND2_X1 #() 
NAND2_X1_5255_ (
  .A1({ S2969 }),
  .A2({ S25957[771] }),
  .ZN({ S3177 })
);
NAND3_X1 #() 
NAND3_X1_5652_ (
  .A1({ S3095 }),
  .A2({ S2901 }),
  .A3({ S3177 }),
  .ZN({ S3178 })
);
NAND2_X1 #() 
NAND2_X1_5256_ (
  .A1({ S2981 }),
  .A2({ S25957[771] }),
  .ZN({ S3179 })
);
NAND4_X1 #() 
NAND4_X1_615_ (
  .A1({ S2910 }),
  .A2({ S3006 }),
  .A3({ S104 }),
  .A4({ S2893 }),
  .ZN({ S3180 })
);
OAI21_X1 #() 
OAI21_X1_2729_ (
  .A({ S3180 }),
  .B1({ S3179 }),
  .B2({ S3022 }),
  .ZN({ S3181 })
);
NAND2_X1 #() 
NAND2_X1_5257_ (
  .A1({ S3181 }),
  .A2({ S25957[772] }),
  .ZN({ S3182 })
);
OAI211_X1 #() 
OAI211_X1_1858_ (
  .A({ S3182 }),
  .B({ S25957[773] }),
  .C1({ S3176 }),
  .C2({ S3178 }),
  .ZN({ S3183 })
);
NOR2_X1 #() 
NOR2_X1_1328_ (
  .A1({ S2949 }),
  .A2({ S2952 }),
  .ZN({ S3184 })
);
OAI21_X1 #() 
OAI21_X1_2730_ (
  .A({ S2901 }),
  .B1({ S3103 }),
  .B2({ S2994 }),
  .ZN({ S3185 })
);
NAND3_X1 #() 
NAND3_X1_5653_ (
  .A1({ S2923 }),
  .A2({ S2921 }),
  .A3({ S104 }),
  .ZN({ S3186 })
);
NAND3_X1 #() 
NAND3_X1_5654_ (
  .A1({ S3047 }),
  .A2({ S25957[771] }),
  .A3({ S2976 }),
  .ZN({ S3187 })
);
NAND3_X1 #() 
NAND3_X1_5655_ (
  .A1({ S3186 }),
  .A2({ S3187 }),
  .A3({ S25957[772] }),
  .ZN({ S3188 })
);
OAI211_X1 #() 
OAI211_X1_1859_ (
  .A({ S3188 }),
  .B({ S2927 }),
  .C1({ S3185 }),
  .C2({ S3184 }),
  .ZN({ S3189 })
);
NAND3_X1 #() 
NAND3_X1_5656_ (
  .A1({ S3183 }),
  .A2({ S25957[775] }),
  .A3({ S3189 }),
  .ZN({ S3190 })
);
AND3_X1 #() 
AND3_X1_224_ (
  .A1({ S2964 }),
  .A2({ S25957[772] }),
  .A3({ S3119 }),
  .ZN({ S3191 })
);
NAND2_X1 #() 
NAND2_X1_5258_ (
  .A1({ S3027 }),
  .A2({ S25957[769] }),
  .ZN({ S3192 })
);
AOI21_X1 #() 
AOI21_X1_2950_ (
  .A({ S25957[772] }),
  .B1({ S3131 }),
  .B2({ S3192 }),
  .ZN({ S3193 })
);
OAI21_X1 #() 
OAI21_X1_2731_ (
  .A({ S25957[773] }),
  .B1({ S3191 }),
  .B2({ S3193 }),
  .ZN({ S3194 })
);
NAND3_X1 #() 
NAND3_X1_5657_ (
  .A1({ S2978 }),
  .A2({ S2948 }),
  .A3({ S25957[771] }),
  .ZN({ S3195 })
);
AOI21_X1 #() 
AOI21_X1_2951_ (
  .A({ S2901 }),
  .B1({ S3195 }),
  .B2({ S3136 }),
  .ZN({ S3196 })
);
NAND3_X1 #() 
NAND3_X1_5658_ (
  .A1({ S2948 }),
  .A2({ S25957[771] }),
  .A3({ S112 }),
  .ZN({ S3197 })
);
NAND3_X1 #() 
NAND3_X1_5659_ (
  .A1({ S2920 }),
  .A2({ S2928 }),
  .A3({ S104 }),
  .ZN({ S3198 })
);
NAND3_X1 #() 
NAND3_X1_5660_ (
  .A1({ S3198 }),
  .A2({ S2901 }),
  .A3({ S3197 }),
  .ZN({ S3199 })
);
NAND2_X1 #() 
NAND2_X1_5259_ (
  .A1({ S3199 }),
  .A2({ S2927 }),
  .ZN({ S3200 })
);
OAI211_X1 #() 
OAI211_X1_1860_ (
  .A({ S3194 }),
  .B({ S2962 }),
  .C1({ S3196 }),
  .C2({ S3200 }),
  .ZN({ S3201 })
);
NAND2_X1 #() 
NAND2_X1_5260_ (
  .A1({ S3201 }),
  .A2({ S3190 }),
  .ZN({ S3202 })
);
NAND2_X1 #() 
NAND2_X1_5261_ (
  .A1({ S3202 }),
  .A2({ S2900 }),
  .ZN({ S3203 })
);
AOI21_X1 #() 
AOI21_X1_2952_ (
  .A({ S25957[972] }),
  .B1({ S3203 }),
  .B2({ S3175 }),
  .ZN({ S3204 })
);
NAND3_X1 #() 
NAND3_X1_5661_ (
  .A1({ S3203 }),
  .A2({ S25957[972] }),
  .A3({ S3175 }),
  .ZN({ S3205 })
);
INV_X1 #() 
INV_X1_1724_ (
  .A({ S3205 }),
  .ZN({ S3206 })
);
OAI21_X1 #() 
OAI21_X1_2732_ (
  .A({ S25416 }),
  .B1({ S3206 }),
  .B2({ S3204 }),
  .ZN({ S3207 })
);
INV_X1 #() 
INV_X1_1725_ (
  .A({ S3204 }),
  .ZN({ S3208 })
);
NAND3_X1 #() 
NAND3_X1_5662_ (
  .A1({ S3208 }),
  .A2({ S25957[908] }),
  .A3({ S3205 }),
  .ZN({ S3209 })
);
NAND2_X1 #() 
NAND2_X1_5262_ (
  .A1({ S3207 }),
  .A2({ S3209 }),
  .ZN({ S25957[652] })
);
NAND2_X1 #() 
NAND2_X1_5263_ (
  .A1({ S23784 }),
  .A2({ S23770 }),
  .ZN({ S25957[971] })
);
INV_X1 #() 
INV_X1_1726_ (
  .A({ S25957[971] }),
  .ZN({ S3210 })
);
NAND3_X1 #() 
NAND3_X1_5663_ (
  .A1({ S2933 }),
  .A2({ S25957[771] }),
  .A3({ S2893 }),
  .ZN({ S3211 })
);
NAND3_X1 #() 
NAND3_X1_5664_ (
  .A1({ S2914 }),
  .A2({ S2937 }),
  .A3({ S104 }),
  .ZN({ S3212 })
);
AOI21_X1 #() 
AOI21_X1_2953_ (
  .A({ S2901 }),
  .B1({ S3212 }),
  .B2({ S3211 }),
  .ZN({ S3213 })
);
AOI21_X1 #() 
AOI21_X1_2954_ (
  .A({ S3213 }),
  .B1({ S3154 }),
  .B2({ S3056 }),
  .ZN({ S3214 })
);
NAND2_X1 #() 
NAND2_X1_5264_ (
  .A1({ S3214 }),
  .A2({ S2927 }),
  .ZN({ S3215 })
);
NAND3_X1 #() 
NAND3_X1_5665_ (
  .A1({ S2968 }),
  .A2({ S25957[771] }),
  .A3({ S3006 }),
  .ZN({ S3216 })
);
NAND3_X1 #() 
NAND3_X1_5666_ (
  .A1({ S2995 }),
  .A2({ S2910 }),
  .A3({ S2936 }),
  .ZN({ S3217 })
);
AOI21_X1 #() 
AOI21_X1_2955_ (
  .A({ S25957[772] }),
  .B1({ S3216 }),
  .B2({ S3217 }),
  .ZN({ S3218 })
);
AOI21_X1 #() 
AOI21_X1_2956_ (
  .A({ S2901 }),
  .B1({ S2995 }),
  .B2({ S2923 }),
  .ZN({ S3219 })
);
AND2_X1 #() 
AND2_X1_334_ (
  .A1({ S3219 }),
  .A2({ S3197 }),
  .ZN({ S3220 })
);
NOR2_X1 #() 
NOR2_X1_1329_ (
  .A1({ S3218 }),
  .A2({ S3220 }),
  .ZN({ S3221 })
);
AOI21_X1 #() 
AOI21_X1_2957_ (
  .A({ S2900 }),
  .B1({ S3221 }),
  .B2({ S25957[773] }),
  .ZN({ S3222 })
);
NAND2_X1 #() 
NAND2_X1_5265_ (
  .A1({ S3222 }),
  .A2({ S3215 }),
  .ZN({ S3223 })
);
NAND4_X1 #() 
NAND4_X1_616_ (
  .A1({ S2910 }),
  .A2({ S2939 }),
  .A3({ S25957[771] }),
  .A4({ S25957[769] }),
  .ZN({ S3224 })
);
NAND3_X1 #() 
NAND3_X1_5667_ (
  .A1({ S2991 }),
  .A2({ S104 }),
  .A3({ S3006 }),
  .ZN({ S3225 })
);
NAND2_X1 #() 
NAND2_X1_5266_ (
  .A1({ S3225 }),
  .A2({ S3224 }),
  .ZN({ S3226 })
);
NAND2_X1 #() 
NAND2_X1_5267_ (
  .A1({ S3226 }),
  .A2({ S2901 }),
  .ZN({ S3227 })
);
AND2_X1 #() 
AND2_X1_335_ (
  .A1({ S2935 }),
  .A2({ S2920 }),
  .ZN({ S3228 })
);
OAI211_X1 #() 
OAI211_X1_1861_ (
  .A({ S104 }),
  .B({ S2939 }),
  .C1({ S2911 }),
  .C2({ S2913 }),
  .ZN({ S3229 })
);
OAI211_X1 #() 
OAI211_X1_1862_ (
  .A({ S25957[772] }),
  .B({ S3229 }),
  .C1({ S3228 }),
  .C2({ S104 }),
  .ZN({ S3230 })
);
AND2_X1 #() 
AND2_X1_336_ (
  .A1({ S3227 }),
  .A2({ S3230 }),
  .ZN({ S3231 })
);
AOI21_X1 #() 
AOI21_X1_2958_ (
  .A({ S25957[768] }),
  .B1({ S2891 }),
  .B2({ S2892 }),
  .ZN({ S3232 })
);
NAND4_X1 #() 
NAND4_X1_617_ (
  .A1({ S25957[770] }),
  .A2({ S25957[771] }),
  .A3({ S2912 }),
  .A4({ S2936 }),
  .ZN({ S3233 })
);
OAI221_X1 #() 
OAI221_X1_158_ (
  .A({ S3233 }),
  .B1({ S104 }),
  .B2({ S3006 }),
  .C1({ S2940 }),
  .C2({ S3232 }),
  .ZN({ S3234 })
);
NAND2_X1 #() 
NAND2_X1_5268_ (
  .A1({ S3234 }),
  .A2({ S2901 }),
  .ZN({ S3235 })
);
NAND3_X1 #() 
NAND3_X1_5668_ (
  .A1({ S3179 }),
  .A2({ S3169 }),
  .A3({ S25957[772] }),
  .ZN({ S3236 })
);
NAND3_X1 #() 
NAND3_X1_5669_ (
  .A1({ S3235 }),
  .A2({ S2927 }),
  .A3({ S3236 }),
  .ZN({ S3237 })
);
OAI211_X1 #() 
OAI211_X1_1863_ (
  .A({ S3237 }),
  .B({ S2900 }),
  .C1({ S3231 }),
  .C2({ S2927 }),
  .ZN({ S3238 })
);
NAND3_X1 #() 
NAND3_X1_5670_ (
  .A1({ S3223 }),
  .A2({ S3238 }),
  .A3({ S25957[775] }),
  .ZN({ S3239 })
);
AOI21_X1 #() 
AOI21_X1_2959_ (
  .A({ S25957[771] }),
  .B1({ S3006 }),
  .B2({ S25957[768] }),
  .ZN({ S3240 })
);
NAND3_X1 #() 
NAND3_X1_5671_ (
  .A1({ S2915 }),
  .A2({ S2901 }),
  .A3({ S3028 }),
  .ZN({ S3241 })
);
OAI21_X1 #() 
OAI21_X1_2733_ (
  .A({ S3241 }),
  .B1({ S2901 }),
  .B2({ S3240 }),
  .ZN({ S3242 })
);
NAND2_X1 #() 
NAND2_X1_5269_ (
  .A1({ S3242 }),
  .A2({ S2927 }),
  .ZN({ S3243 })
);
NAND3_X1 #() 
NAND3_X1_5672_ (
  .A1({ S2933 }),
  .A2({ S25957[771] }),
  .A3({ S2898 }),
  .ZN({ S3244 })
);
AOI21_X1 #() 
AOI21_X1_2960_ (
  .A({ S25957[772] }),
  .B1({ S2995 }),
  .B2({ S2976 }),
  .ZN({ S3245 })
);
AOI22_X1 #() 
AOI22_X1_598_ (
  .A1({ S2992 }),
  .A2({ S3023 }),
  .B1({ S3245 }),
  .B2({ S3244 }),
  .ZN({ S3246 })
);
OAI211_X1 #() 
OAI211_X1_1864_ (
  .A({ S3243 }),
  .B({ S25957[774] }),
  .C1({ S3246 }),
  .C2({ S2927 }),
  .ZN({ S3247 })
);
NAND3_X1 #() 
NAND3_X1_5673_ (
  .A1({ S2935 }),
  .A2({ S25957[771] }),
  .A3({ S3034 }),
  .ZN({ S3248 })
);
NAND3_X1 #() 
NAND3_X1_5674_ (
  .A1({ S3071 }),
  .A2({ S25957[772] }),
  .A3({ S3248 }),
  .ZN({ S3249 })
);
AOI21_X1 #() 
AOI21_X1_2961_ (
  .A({ S104 }),
  .B1({ S2999 }),
  .B2({ S2948 }),
  .ZN({ S3250 })
);
OAI21_X1 #() 
OAI21_X1_2734_ (
  .A({ S2901 }),
  .B1({ S2983 }),
  .B2({ S3250 }),
  .ZN({ S3251 })
);
NAND3_X1 #() 
NAND3_X1_5675_ (
  .A1({ S3251 }),
  .A2({ S3249 }),
  .A3({ S2927 }),
  .ZN({ S3252 })
);
NAND3_X1 #() 
NAND3_X1_5676_ (
  .A1({ S2996 }),
  .A2({ S25957[772] }),
  .A3({ S3031 }),
  .ZN({ S3253 })
);
NAND3_X1 #() 
NAND3_X1_5677_ (
  .A1({ S2906 }),
  .A2({ S2910 }),
  .A3({ S2978 }),
  .ZN({ S3254 })
);
NAND2_X1 #() 
NAND2_X1_5270_ (
  .A1({ S3254 }),
  .A2({ S2901 }),
  .ZN({ S3255 })
);
NAND3_X1 #() 
NAND3_X1_5678_ (
  .A1({ S3255 }),
  .A2({ S25957[773] }),
  .A3({ S3253 }),
  .ZN({ S3256 })
);
NAND3_X1 #() 
NAND3_X1_5679_ (
  .A1({ S3252 }),
  .A2({ S2900 }),
  .A3({ S3256 }),
  .ZN({ S3257 })
);
NAND3_X1 #() 
NAND3_X1_5680_ (
  .A1({ S3247 }),
  .A2({ S2962 }),
  .A3({ S3257 }),
  .ZN({ S3258 })
);
AOI21_X1 #() 
AOI21_X1_2962_ (
  .A({ S3210 }),
  .B1({ S3239 }),
  .B2({ S3258 }),
  .ZN({ S3259 })
);
OAI21_X1 #() 
OAI21_X1_2735_ (
  .A({ S25957[773] }),
  .B1({ S3218 }),
  .B2({ S3220 }),
  .ZN({ S3260 })
);
OAI211_X1 #() 
OAI211_X1_1865_ (
  .A({ S25957[774] }),
  .B({ S3260 }),
  .C1({ S3214 }),
  .C2({ S25957[773] }),
  .ZN({ S3261 })
);
AND2_X1 #() 
AND2_X1_337_ (
  .A1({ S3235 }),
  .A2({ S3236 }),
  .ZN({ S3262 })
);
NAND3_X1 #() 
NAND3_X1_5681_ (
  .A1({ S3227 }),
  .A2({ S3230 }),
  .A3({ S25957[773] }),
  .ZN({ S3263 })
);
OAI211_X1 #() 
OAI211_X1_1866_ (
  .A({ S3263 }),
  .B({ S2900 }),
  .C1({ S3262 }),
  .C2({ S25957[773] }),
  .ZN({ S3264 })
);
NAND3_X1 #() 
NAND3_X1_5682_ (
  .A1({ S3264 }),
  .A2({ S25957[775] }),
  .A3({ S3261 }),
  .ZN({ S3265 })
);
NAND2_X1 #() 
NAND2_X1_5271_ (
  .A1({ S3246 }),
  .A2({ S25957[773] }),
  .ZN({ S3266 })
);
OAI211_X1 #() 
OAI211_X1_1867_ (
  .A({ S3241 }),
  .B({ S2927 }),
  .C1({ S2901 }),
  .C2({ S3240 }),
  .ZN({ S3267 })
);
NAND3_X1 #() 
NAND3_X1_5683_ (
  .A1({ S3266 }),
  .A2({ S25957[774] }),
  .A3({ S3267 }),
  .ZN({ S3268 })
);
AND2_X1 #() 
AND2_X1_338_ (
  .A1({ S3252 }),
  .A2({ S3256 }),
  .ZN({ S3269 })
);
OAI211_X1 #() 
OAI211_X1_1868_ (
  .A({ S3268 }),
  .B({ S2962 }),
  .C1({ S25957[774] }),
  .C2({ S3269 }),
  .ZN({ S3270 })
);
AOI21_X1 #() 
AOI21_X1_2963_ (
  .A({ S25957[971] }),
  .B1({ S3270 }),
  .B2({ S3265 }),
  .ZN({ S3271 })
);
OAI21_X1 #() 
OAI21_X1_2736_ (
  .A({ S89 }),
  .B1({ S3271 }),
  .B2({ S3259 }),
  .ZN({ S3272 })
);
NAND3_X1 #() 
NAND3_X1_5684_ (
  .A1({ S3270 }),
  .A2({ S3265 }),
  .A3({ S25957[971] }),
  .ZN({ S3273 })
);
NAND3_X1 #() 
NAND3_X1_5685_ (
  .A1({ S3239 }),
  .A2({ S3258 }),
  .A3({ S3210 }),
  .ZN({ S3274 })
);
NAND3_X1 #() 
NAND3_X1_5686_ (
  .A1({ S3273 }),
  .A2({ S3274 }),
  .A3({ S25957[907] }),
  .ZN({ S3275 })
);
NAND2_X1 #() 
NAND2_X1_5272_ (
  .A1({ S3272 }),
  .A2({ S3275 }),
  .ZN({ S113 })
);
AND2_X1 #() 
AND2_X1_339_ (
  .A1({ S3272 }),
  .A2({ S3275 }),
  .ZN({ S25957[651] })
);
NOR2_X1 #() 
NOR2_X1_1330_ (
  .A1({ S16516 }),
  .A2({ S16560 }),
  .ZN({ S25957[1192] })
);
NAND2_X1 #() 
NAND2_X1_5273_ (
  .A1({ S21258 }),
  .A2({ S21261 }),
  .ZN({ S25957[1096] })
);
XOR2_X1 #() 
XOR2_X1_87_ (
  .A({ S25957[1096] }),
  .B({ S25957[1192] }),
  .Z({ S25957[1064] })
);
INV_X1 #() 
INV_X1_1727_ (
  .A({ S25957[1064] }),
  .ZN({ S3276 })
);
XNOR2_X1 #() 
XNOR2_X1_204_ (
  .A({ S25957[968] }),
  .B({ S3276 }),
  .ZN({ S25957[936] })
);
INV_X1 #() 
INV_X1_1728_ (
  .A({ S25957[936] }),
  .ZN({ S3277 })
);
NAND2_X1 #() 
NAND2_X1_5274_ (
  .A1({ S860 }),
  .A2({ S840 }),
  .ZN({ S3278 })
);
NAND3_X1 #() 
NAND3_X1_5687_ (
  .A1({ S2939 }),
  .A2({ S25957[771] }),
  .A3({ S2893 }),
  .ZN({ S3279 })
);
NAND4_X1 #() 
NAND4_X1_618_ (
  .A1({ S2921 }),
  .A2({ S2933 }),
  .A3({ S3006 }),
  .A4({ S104 }),
  .ZN({ S3280 })
);
NAND3_X1 #() 
NAND3_X1_5688_ (
  .A1({ S3280 }),
  .A2({ S25957[772] }),
  .A3({ S3279 }),
  .ZN({ S3281 })
);
NAND3_X1 #() 
NAND3_X1_5689_ (
  .A1({ S3090 }),
  .A2({ S3123 }),
  .A3({ S2901 }),
  .ZN({ S3282 })
);
NAND2_X1 #() 
NAND2_X1_5275_ (
  .A1({ S3281 }),
  .A2({ S3282 }),
  .ZN({ S3283 })
);
NAND2_X1 #() 
NAND2_X1_5276_ (
  .A1({ S3283 }),
  .A2({ S2927 }),
  .ZN({ S3284 })
);
OAI21_X1 #() 
OAI21_X1_2737_ (
  .A({ S25957[771] }),
  .B1({ S2904 }),
  .B2({ S2903 }),
  .ZN({ S3285 })
);
OAI21_X1 #() 
OAI21_X1_2738_ (
  .A({ S2901 }),
  .B1({ S3285 }),
  .B2({ S2936 }),
  .ZN({ S3286 })
);
NAND4_X1 #() 
NAND4_X1_619_ (
  .A1({ S2936 }),
  .A2({ S1618 }),
  .A3({ S25957[771] }),
  .A4({ S1621 }),
  .ZN({ S3287 })
);
NAND2_X1 #() 
NAND2_X1_5277_ (
  .A1({ S2970 }),
  .A2({ S3287 }),
  .ZN({ S3288 })
);
AOI21_X1 #() 
AOI21_X1_2964_ (
  .A({ S104 }),
  .B1({ S2991 }),
  .B2({ S2921 }),
  .ZN({ S3289 })
);
NAND2_X1 #() 
NAND2_X1_5278_ (
  .A1({ S2936 }),
  .A2({ S104 }),
  .ZN({ S3290 })
);
OAI21_X1 #() 
OAI21_X1_2739_ (
  .A({ S25957[772] }),
  .B1({ S3030 }),
  .B2({ S3290 }),
  .ZN({ S3291 })
);
OAI221_X1 #() 
OAI221_X1_159_ (
  .A({ S25957[773] }),
  .B1({ S3288 }),
  .B2({ S3286 }),
  .C1({ S3289 }),
  .C2({ S3291 }),
  .ZN({ S3292 })
);
NAND3_X1 #() 
NAND3_X1_5690_ (
  .A1({ S3284 }),
  .A2({ S25957[774] }),
  .A3({ S3292 }),
  .ZN({ S3293 })
);
NAND3_X1 #() 
NAND3_X1_5691_ (
  .A1({ S2991 }),
  .A2({ S25957[771] }),
  .A3({ S2928 }),
  .ZN({ S3294 })
);
NAND3_X1 #() 
NAND3_X1_5692_ (
  .A1({ S2978 }),
  .A2({ S3034 }),
  .A3({ S104 }),
  .ZN({ S3295 })
);
NAND3_X1 #() 
NAND3_X1_5693_ (
  .A1({ S3294 }),
  .A2({ S2901 }),
  .A3({ S3295 }),
  .ZN({ S3296 })
);
AOI21_X1 #() 
AOI21_X1_2965_ (
  .A({ S2901 }),
  .B1({ S2911 }),
  .B2({ S3059 }),
  .ZN({ S3297 })
);
NAND3_X1 #() 
NAND3_X1_5694_ (
  .A1({ S3297 }),
  .A2({ S2996 }),
  .A3({ S3179 }),
  .ZN({ S3298 })
);
NAND3_X1 #() 
NAND3_X1_5695_ (
  .A1({ S3296 }),
  .A2({ S3298 }),
  .A3({ S2927 }),
  .ZN({ S3299 })
);
NAND3_X1 #() 
NAND3_X1_5696_ (
  .A1({ S3109 }),
  .A2({ S3035 }),
  .A3({ S2901 }),
  .ZN({ S3300 })
);
NAND3_X1 #() 
NAND3_X1_5697_ (
  .A1({ S3087 }),
  .A2({ S3197 }),
  .A3({ S25957[772] }),
  .ZN({ S3301 })
);
NAND3_X1 #() 
NAND3_X1_5698_ (
  .A1({ S3300 }),
  .A2({ S25957[773] }),
  .A3({ S3301 }),
  .ZN({ S3302 })
);
NAND2_X1 #() 
NAND2_X1_5279_ (
  .A1({ S3299 }),
  .A2({ S3302 }),
  .ZN({ S3303 })
);
NAND2_X1 #() 
NAND2_X1_5280_ (
  .A1({ S3303 }),
  .A2({ S2900 }),
  .ZN({ S3304 })
);
NAND3_X1 #() 
NAND3_X1_5699_ (
  .A1({ S3304 }),
  .A2({ S3293 }),
  .A3({ S2962 }),
  .ZN({ S3305 })
);
NAND3_X1 #() 
NAND3_X1_5700_ (
  .A1({ S3090 }),
  .A2({ S2901 }),
  .A3({ S3103 }),
  .ZN({ S3306 })
);
NAND2_X1 #() 
NAND2_X1_5281_ (
  .A1({ S2937 }),
  .A2({ S25957[771] }),
  .ZN({ S3307 })
);
NAND2_X1 #() 
NAND2_X1_5282_ (
  .A1({ S3307 }),
  .A2({ S3180 }),
  .ZN({ S3308 })
);
AOI21_X1 #() 
AOI21_X1_2966_ (
  .A({ S25957[773] }),
  .B1({ S3308 }),
  .B2({ S25957[772] }),
  .ZN({ S3309 })
);
NAND2_X1 #() 
NAND2_X1_5283_ (
  .A1({ S2944 }),
  .A2({ S104 }),
  .ZN({ S3310 })
);
NAND3_X1 #() 
NAND3_X1_5701_ (
  .A1({ S3310 }),
  .A2({ S2901 }),
  .A3({ S3195 }),
  .ZN({ S3311 })
);
AOI21_X1 #() 
AOI21_X1_2967_ (
  .A({ S2901 }),
  .B1({ S2994 }),
  .B2({ S25957[771] }),
  .ZN({ S3312 })
);
AOI21_X1 #() 
AOI21_X1_2968_ (
  .A({ S2927 }),
  .B1({ S3312 }),
  .B2({ S3198 }),
  .ZN({ S3313 })
);
AOI22_X1 #() 
AOI22_X1_599_ (
  .A1({ S3309 }),
  .A2({ S3306 }),
  .B1({ S3311 }),
  .B2({ S3313 }),
  .ZN({ S3314 })
);
AOI21_X1 #() 
AOI21_X1_2969_ (
  .A({ S104 }),
  .B1({ S25957[770] }),
  .B2({ S3232 }),
  .ZN({ S3315 })
);
NAND3_X1 #() 
NAND3_X1_5702_ (
  .A1({ S2933 }),
  .A2({ S104 }),
  .A3({ S2898 }),
  .ZN({ S3316 })
);
OAI211_X1 #() 
OAI211_X1_1869_ (
  .A({ S25957[772] }),
  .B({ S3316 }),
  .C1({ S3240 }),
  .C2({ S3315 }),
  .ZN({ S3317 })
);
OAI211_X1 #() 
OAI211_X1_1870_ (
  .A({ S2978 }),
  .B({ S3163 }),
  .C1({ S3285 }),
  .C2({ S2936 }),
  .ZN({ S3318 })
);
NAND2_X1 #() 
NAND2_X1_5284_ (
  .A1({ S3318 }),
  .A2({ S2901 }),
  .ZN({ S3319 })
);
NAND3_X1 #() 
NAND3_X1_5703_ (
  .A1({ S3317 }),
  .A2({ S25957[773] }),
  .A3({ S3319 }),
  .ZN({ S3320 })
);
OAI211_X1 #() 
OAI211_X1_1871_ (
  .A({ S2972 }),
  .B({ S25957[772] }),
  .C1({ S2935 }),
  .C2({ S25957[771] }),
  .ZN({ S3321 })
);
AOI21_X1 #() 
AOI21_X1_2970_ (
  .A({ S104 }),
  .B1({ S2916 }),
  .B2({ S112 }),
  .ZN({ S3322 })
);
AOI21_X1 #() 
AOI21_X1_2971_ (
  .A({ S25957[771] }),
  .B1({ S2923 }),
  .B2({ S2939 }),
  .ZN({ S3323 })
);
OAI21_X1 #() 
OAI21_X1_2740_ (
  .A({ S2901 }),
  .B1({ S3323 }),
  .B2({ S3322 }),
  .ZN({ S3324 })
);
NAND3_X1 #() 
NAND3_X1_5704_ (
  .A1({ S3324 }),
  .A2({ S2927 }),
  .A3({ S3321 }),
  .ZN({ S3325 })
);
NAND3_X1 #() 
NAND3_X1_5705_ (
  .A1({ S3325 }),
  .A2({ S3320 }),
  .A3({ S2900 }),
  .ZN({ S3326 })
);
OAI211_X1 #() 
OAI211_X1_1872_ (
  .A({ S25957[775] }),
  .B({ S3326 }),
  .C1({ S3314 }),
  .C2({ S2900 }),
  .ZN({ S3327 })
);
NAND3_X1 #() 
NAND3_X1_5706_ (
  .A1({ S3305 }),
  .A2({ S3327 }),
  .A3({ S3278 }),
  .ZN({ S3328 })
);
INV_X1 #() 
INV_X1_1729_ (
  .A({ S3278 }),
  .ZN({ S25957[872] })
);
AOI21_X1 #() 
AOI21_X1_2972_ (
  .A({ S25957[771] }),
  .B1({ S2911 }),
  .B2({ S2902 }),
  .ZN({ S3329 })
);
AOI22_X1 #() 
AOI22_X1_600_ (
  .A1({ S3329 }),
  .A2({ S2968 }),
  .B1({ S25957[771] }),
  .B2({ S2937 }),
  .ZN({ S3330 })
);
OAI211_X1 #() 
OAI211_X1_1873_ (
  .A({ S2927 }),
  .B({ S3306 }),
  .C1({ S3330 }),
  .C2({ S2901 }),
  .ZN({ S3331 })
);
AOI21_X1 #() 
AOI21_X1_2973_ (
  .A({ S25957[771] }),
  .B1({ S2935 }),
  .B2({ S2933 }),
  .ZN({ S3332 })
);
NAND2_X1 #() 
NAND2_X1_5285_ (
  .A1({ S3195 }),
  .A2({ S2901 }),
  .ZN({ S3333 })
);
NAND3_X1 #() 
NAND3_X1_5707_ (
  .A1({ S25957[770] }),
  .A2({ S25957[771] }),
  .A3({ S2936 }),
  .ZN({ S3334 })
);
NAND3_X1 #() 
NAND3_X1_5708_ (
  .A1({ S3198 }),
  .A2({ S25957[772] }),
  .A3({ S3334 }),
  .ZN({ S3335 })
);
OAI211_X1 #() 
OAI211_X1_1874_ (
  .A({ S3335 }),
  .B({ S25957[773] }),
  .C1({ S3332 }),
  .C2({ S3333 }),
  .ZN({ S3336 })
);
AOI21_X1 #() 
AOI21_X1_2974_ (
  .A({ S2900 }),
  .B1({ S3331 }),
  .B2({ S3336 }),
  .ZN({ S3337 })
);
AND3_X1 #() 
AND3_X1_225_ (
  .A1({ S3325 }),
  .A2({ S3320 }),
  .A3({ S2900 }),
  .ZN({ S3338 })
);
OAI21_X1 #() 
OAI21_X1_2741_ (
  .A({ S25957[775] }),
  .B1({ S3338 }),
  .B2({ S3337 }),
  .ZN({ S3339 })
);
OAI22_X1 #() 
OAI22_X1_135_ (
  .A1({ S3289 }),
  .A2({ S3291 }),
  .B1({ S3288 }),
  .B2({ S3286 }),
  .ZN({ S3340 })
);
NAND2_X1 #() 
NAND2_X1_5286_ (
  .A1({ S3340 }),
  .A2({ S25957[773] }),
  .ZN({ S3341 })
);
NAND3_X1 #() 
NAND3_X1_5709_ (
  .A1({ S3281 }),
  .A2({ S3282 }),
  .A3({ S2927 }),
  .ZN({ S3342 })
);
AOI21_X1 #() 
AOI21_X1_2975_ (
  .A({ S2900 }),
  .B1({ S3341 }),
  .B2({ S3342 }),
  .ZN({ S3343 })
);
AOI21_X1 #() 
AOI21_X1_2976_ (
  .A({ S25957[774] }),
  .B1({ S3299 }),
  .B2({ S3302 }),
  .ZN({ S3344 })
);
OAI21_X1 #() 
OAI21_X1_2742_ (
  .A({ S2962 }),
  .B1({ S3343 }),
  .B2({ S3344 }),
  .ZN({ S3345 })
);
NAND3_X1 #() 
NAND3_X1_5710_ (
  .A1({ S3339 }),
  .A2({ S3345 }),
  .A3({ S25957[872] }),
  .ZN({ S3346 })
);
AOI21_X1 #() 
AOI21_X1_2977_ (
  .A({ S3277 }),
  .B1({ S3346 }),
  .B2({ S3328 }),
  .ZN({ S3347 })
);
NAND3_X1 #() 
NAND3_X1_5711_ (
  .A1({ S3339 }),
  .A2({ S3345 }),
  .A3({ S3278 }),
  .ZN({ S3348 })
);
NAND3_X1 #() 
NAND3_X1_5712_ (
  .A1({ S3305 }),
  .A2({ S3327 }),
  .A3({ S25957[872] }),
  .ZN({ S3349 })
);
AOI21_X1 #() 
AOI21_X1_2978_ (
  .A({ S25957[936] }),
  .B1({ S3348 }),
  .B2({ S3349 }),
  .ZN({ S3350 })
);
OAI21_X1 #() 
OAI21_X1_2743_ (
  .A({ S2282 }),
  .B1({ S3347 }),
  .B2({ S3350 }),
  .ZN({ S3351 })
);
NAND3_X1 #() 
NAND3_X1_5713_ (
  .A1({ S3348 }),
  .A2({ S3349 }),
  .A3({ S25957[936] }),
  .ZN({ S3352 })
);
NAND3_X1 #() 
NAND3_X1_5714_ (
  .A1({ S3346 }),
  .A2({ S3328 }),
  .A3({ S3277 }),
  .ZN({ S3353 })
);
NAND3_X1 #() 
NAND3_X1_5715_ (
  .A1({ S3352 }),
  .A2({ S3353 }),
  .A3({ S25957[776] }),
  .ZN({ S3354 })
);
NAND2_X1 #() 
NAND2_X1_5287_ (
  .A1({ S3351 }),
  .A2({ S3354 }),
  .ZN({ S25957[648] })
);
NAND2_X1 #() 
NAND2_X1_5288_ (
  .A1({ S23923 }),
  .A2({ S23924 }),
  .ZN({ S25957[937] })
);
NOR2_X1 #() 
NOR2_X1_1331_ (
  .A1({ S2233 }),
  .A2({ S2234 }),
  .ZN({ S25957[841] })
);
XOR2_X1 #() 
XOR2_X1_88_ (
  .A({ S25957[841] }),
  .B({ S25957[937] }),
  .Z({ S25957[809] })
);
INV_X1 #() 
INV_X1_1730_ (
  .A({ S25957[809] }),
  .ZN({ S3355 })
);
INV_X1 #() 
INV_X1_1731_ (
  .A({ S25957[841] }),
  .ZN({ S3356 })
);
NAND2_X1 #() 
NAND2_X1_5289_ (
  .A1({ S940 }),
  .A2({ S911 }),
  .ZN({ S25957[873] })
);
INV_X1 #() 
INV_X1_1732_ (
  .A({ S25957[873] }),
  .ZN({ S3357 })
);
NAND3_X1 #() 
NAND3_X1_5716_ (
  .A1({ S2920 }),
  .A2({ S104 }),
  .A3({ S2939 }),
  .ZN({ S3358 })
);
NAND3_X1 #() 
NAND3_X1_5717_ (
  .A1({ S3248 }),
  .A2({ S3358 }),
  .A3({ S25957[772] }),
  .ZN({ S3359 })
);
NAND3_X1 #() 
NAND3_X1_5718_ (
  .A1({ S2910 }),
  .A2({ S2939 }),
  .A3({ S2936 }),
  .ZN({ S3360 })
);
NOR2_X1 #() 
NOR2_X1_1332_ (
  .A1({ S2929 }),
  .A2({ S25957[772] }),
  .ZN({ S3361 })
);
AOI21_X1 #() 
AOI21_X1_2979_ (
  .A({ S2927 }),
  .B1({ S3360 }),
  .B2({ S3361 }),
  .ZN({ S3362 })
);
NAND2_X1 #() 
NAND2_X1_5290_ (
  .A1({ S3362 }),
  .A2({ S3359 }),
  .ZN({ S3363 })
);
AOI22_X1 #() 
AOI22_X1_601_ (
  .A1({ S1618 }),
  .A2({ S1621 }),
  .B1({ S25957[769] }),
  .B2({ S25957[768] }),
  .ZN({ S3364 })
);
OAI211_X1 #() 
OAI211_X1_1875_ (
  .A({ S3233 }),
  .B({ S2901 }),
  .C1({ S2940 }),
  .C2({ S3364 }),
  .ZN({ S3365 })
);
NAND3_X1 #() 
NAND3_X1_5719_ (
  .A1({ S3041 }),
  .A2({ S2955 }),
  .A3({ S104 }),
  .ZN({ S3366 })
);
NAND2_X1 #() 
NAND2_X1_5291_ (
  .A1({ S3366 }),
  .A2({ S25957[772] }),
  .ZN({ S3367 })
);
OAI211_X1 #() 
OAI211_X1_1876_ (
  .A({ S3365 }),
  .B({ S2927 }),
  .C1({ S3367 }),
  .C2({ S3289 }),
  .ZN({ S3368 })
);
NAND3_X1 #() 
NAND3_X1_5720_ (
  .A1({ S3368 }),
  .A2({ S3363 }),
  .A3({ S25957[774] }),
  .ZN({ S3369 })
);
AOI21_X1 #() 
AOI21_X1_2980_ (
  .A({ S2901 }),
  .B1({ S3224 }),
  .B2({ S3166 }),
  .ZN({ S3370 })
);
OAI21_X1 #() 
OAI21_X1_2744_ (
  .A({ S25957[773] }),
  .B1({ S3370 }),
  .B2({ S2980 }),
  .ZN({ S3371 })
);
NAND4_X1 #() 
NAND4_X1_620_ (
  .A1({ S3169 }),
  .A2({ S2952 }),
  .A3({ S2951 }),
  .A4({ S25957[772] }),
  .ZN({ S3372 })
);
AOI21_X1 #() 
AOI21_X1_2981_ (
  .A({ S25957[773] }),
  .B1({ S3028 }),
  .B2({ S2945 }),
  .ZN({ S3373 })
);
AOI21_X1 #() 
AOI21_X1_2982_ (
  .A({ S25957[774] }),
  .B1({ S3373 }),
  .B2({ S3372 }),
  .ZN({ S3374 })
);
NAND2_X1 #() 
NAND2_X1_5292_ (
  .A1({ S3371 }),
  .A2({ S3374 }),
  .ZN({ S3375 })
);
NAND3_X1 #() 
NAND3_X1_5721_ (
  .A1({ S3369 }),
  .A2({ S3375 }),
  .A3({ S2962 }),
  .ZN({ S3376 })
);
NAND3_X1 #() 
NAND3_X1_5722_ (
  .A1({ S3099 }),
  .A2({ S25957[772] }),
  .A3({ S3316 }),
  .ZN({ S3377 })
);
NAND3_X1 #() 
NAND3_X1_5723_ (
  .A1({ S2910 }),
  .A2({ S25957[771] }),
  .A3({ S2893 }),
  .ZN({ S3378 })
);
NAND2_X1 #() 
NAND2_X1_5293_ (
  .A1({ S2948 }),
  .A2({ S2893 }),
  .ZN({ S3379 })
);
OAI211_X1 #() 
OAI211_X1_1877_ (
  .A({ S2901 }),
  .B({ S3378 }),
  .C1({ S2956 }),
  .C2({ S3379 }),
  .ZN({ S3380 })
);
NAND3_X1 #() 
NAND3_X1_5724_ (
  .A1({ S3377 }),
  .A2({ S3380 }),
  .A3({ S2927 }),
  .ZN({ S3381 })
);
OAI21_X1 #() 
OAI21_X1_2745_ (
  .A({ S2901 }),
  .B1({ S2969 }),
  .B2({ S25957[771] }),
  .ZN({ S3382 })
);
NAND3_X1 #() 
NAND3_X1_5725_ (
  .A1({ S3211 }),
  .A2({ S2966 }),
  .A3({ S25957[772] }),
  .ZN({ S3383 })
);
OAI211_X1 #() 
OAI211_X1_1878_ (
  .A({ S3383 }),
  .B({ S25957[773] }),
  .C1({ S3289 }),
  .C2({ S3382 }),
  .ZN({ S3384 })
);
NAND3_X1 #() 
NAND3_X1_5726_ (
  .A1({ S3381 }),
  .A2({ S3384 }),
  .A3({ S25957[774] }),
  .ZN({ S3385 })
);
AOI21_X1 #() 
AOI21_X1_2983_ (
  .A({ S104 }),
  .B1({ S2937 }),
  .B2({ S2916 }),
  .ZN({ S3386 })
);
OAI21_X1 #() 
OAI21_X1_2746_ (
  .A({ S25957[772] }),
  .B1({ S2970 }),
  .B2({ S2969 }),
  .ZN({ S3387 })
);
NAND2_X1 #() 
NAND2_X1_5294_ (
  .A1({ S2995 }),
  .A2({ S2976 }),
  .ZN({ S3388 })
);
NAND3_X1 #() 
NAND3_X1_5727_ (
  .A1({ S3388 }),
  .A2({ S3118 }),
  .A3({ S2901 }),
  .ZN({ S3389 })
);
OAI211_X1 #() 
OAI211_X1_1879_ (
  .A({ S3389 }),
  .B({ S25957[773] }),
  .C1({ S3387 }),
  .C2({ S3386 }),
  .ZN({ S3390 })
);
NAND3_X1 #() 
NAND3_X1_5728_ (
  .A1({ S3044 }),
  .A2({ S2905 }),
  .A3({ S104 }),
  .ZN({ S3391 })
);
NAND3_X1 #() 
NAND3_X1_5729_ (
  .A1({ S3391 }),
  .A2({ S25957[772] }),
  .A3({ S3066 }),
  .ZN({ S3392 })
);
OAI211_X1 #() 
OAI211_X1_1880_ (
  .A({ S3392 }),
  .B({ S2927 }),
  .C1({ S3185 }),
  .C2({ S2982 }),
  .ZN({ S3393 })
);
NAND3_X1 #() 
NAND3_X1_5730_ (
  .A1({ S3393 }),
  .A2({ S3390 }),
  .A3({ S2900 }),
  .ZN({ S3394 })
);
NAND3_X1 #() 
NAND3_X1_5731_ (
  .A1({ S3385 }),
  .A2({ S3394 }),
  .A3({ S25957[775] }),
  .ZN({ S3395 })
);
NAND3_X1 #() 
NAND3_X1_5732_ (
  .A1({ S3395 }),
  .A2({ S3376 }),
  .A3({ S3357 }),
  .ZN({ S3396 })
);
NAND2_X1 #() 
NAND2_X1_5295_ (
  .A1({ S3395 }),
  .A2({ S3376 }),
  .ZN({ S3397 })
);
NAND2_X1 #() 
NAND2_X1_5296_ (
  .A1({ S3397 }),
  .A2({ S25957[873] }),
  .ZN({ S3398 })
);
NAND3_X1 #() 
NAND3_X1_5733_ (
  .A1({ S3398 }),
  .A2({ S3356 }),
  .A3({ S3396 }),
  .ZN({ S3399 })
);
NAND3_X1 #() 
NAND3_X1_5734_ (
  .A1({ S3395 }),
  .A2({ S3376 }),
  .A3({ S25957[873] }),
  .ZN({ S3400 })
);
NAND2_X1 #() 
NAND2_X1_5297_ (
  .A1({ S3397 }),
  .A2({ S3357 }),
  .ZN({ S3401 })
);
NAND3_X1 #() 
NAND3_X1_5735_ (
  .A1({ S3401 }),
  .A2({ S25957[841] }),
  .A3({ S3400 }),
  .ZN({ S3402 })
);
NAND3_X1 #() 
NAND3_X1_5736_ (
  .A1({ S3399 }),
  .A2({ S3402 }),
  .A3({ S3355 }),
  .ZN({ S3403 })
);
AOI21_X1 #() 
AOI21_X1_2984_ (
  .A({ S25957[841] }),
  .B1({ S3401 }),
  .B2({ S3400 }),
  .ZN({ S3404 })
);
AOI21_X1 #() 
AOI21_X1_2985_ (
  .A({ S3356 }),
  .B1({ S3398 }),
  .B2({ S3396 }),
  .ZN({ S3405 })
);
OAI21_X1 #() 
OAI21_X1_2747_ (
  .A({ S25957[809] }),
  .B1({ S3404 }),
  .B2({ S3405 }),
  .ZN({ S3406 })
);
NAND3_X1 #() 
NAND3_X1_5737_ (
  .A1({ S3406 }),
  .A2({ S25957[777] }),
  .A3({ S3403 }),
  .ZN({ S3407 })
);
OAI21_X1 #() 
OAI21_X1_2748_ (
  .A({ S3355 }),
  .B1({ S3404 }),
  .B2({ S3405 }),
  .ZN({ S3408 })
);
NAND3_X1 #() 
NAND3_X1_5738_ (
  .A1({ S3399 }),
  .A2({ S3402 }),
  .A3({ S25957[809] }),
  .ZN({ S3409 })
);
NAND3_X1 #() 
NAND3_X1_5739_ (
  .A1({ S3408 }),
  .A2({ S2258 }),
  .A3({ S3409 }),
  .ZN({ S3410 })
);
NAND2_X1 #() 
NAND2_X1_5298_ (
  .A1({ S3407 }),
  .A2({ S3410 }),
  .ZN({ S25957[649] })
);
NAND2_X1 #() 
NAND2_X1_5299_ (
  .A1({ S1011 }),
  .A2({ S1012 }),
  .ZN({ S3411 })
);
INV_X1 #() 
INV_X1_1733_ (
  .A({ S3411 }),
  .ZN({ S25957[810] })
);
NOR2_X1 #() 
NOR2_X1_1333_ (
  .A1({ S24007 }),
  .A2({ S24008 }),
  .ZN({ S25957[970] })
);
INV_X1 #() 
INV_X1_1734_ (
  .A({ S25957[970] }),
  .ZN({ S3412 })
);
NAND3_X1 #() 
NAND3_X1_5740_ (
  .A1({ S2935 }),
  .A2({ S25957[771] }),
  .A3({ S3047 }),
  .ZN({ S3413 })
);
AND3_X1 #() 
AND3_X1_226_ (
  .A1({ S3002 }),
  .A2({ S3413 }),
  .A3({ S2901 }),
  .ZN({ S3414 })
);
NAND2_X1 #() 
NAND2_X1_5300_ (
  .A1({ S2977 }),
  .A2({ S25957[772] }),
  .ZN({ S3415 })
);
OAI21_X1 #() 
OAI21_X1_2749_ (
  .A({ S25957[773] }),
  .B1({ S3415 }),
  .B2({ S3332 }),
  .ZN({ S3416 })
);
OAI21_X1 #() 
OAI21_X1_2750_ (
  .A({ S3132 }),
  .B1({ S2944 }),
  .B2({ S2988 }),
  .ZN({ S3417 })
);
AOI21_X1 #() 
AOI21_X1_2986_ (
  .A({ S25957[772] }),
  .B1({ S3059 }),
  .B2({ S2911 }),
  .ZN({ S3418 })
);
AOI21_X1 #() 
AOI21_X1_2987_ (
  .A({ S25957[773] }),
  .B1({ S3418 }),
  .B2({ S3003 }),
  .ZN({ S3419 })
);
NAND2_X1 #() 
NAND2_X1_5301_ (
  .A1({ S3417 }),
  .A2({ S3419 }),
  .ZN({ S3420 })
);
OAI211_X1 #() 
OAI211_X1_1881_ (
  .A({ S3420 }),
  .B({ S25957[774] }),
  .C1({ S3416 }),
  .C2({ S3414 }),
  .ZN({ S3421 })
);
NAND2_X1 #() 
NAND2_X1_5302_ (
  .A1({ S3034 }),
  .A2({ S104 }),
  .ZN({ S3422 })
);
OAI211_X1 #() 
OAI211_X1_1882_ (
  .A({ S25957[771] }),
  .B({ S2936 }),
  .C1({ S2911 }),
  .C2({ S2912 }),
  .ZN({ S3423 })
);
AOI21_X1 #() 
AOI21_X1_2988_ (
  .A({ S25957[772] }),
  .B1({ S3423 }),
  .B2({ S3422 }),
  .ZN({ S3424 })
);
NAND3_X1 #() 
NAND3_X1_5741_ (
  .A1({ S3006 }),
  .A2({ S25957[771] }),
  .A3({ S25957[768] }),
  .ZN({ S3425 })
);
AOI21_X1 #() 
AOI21_X1_2989_ (
  .A({ S2901 }),
  .B1({ S3028 }),
  .B2({ S3425 }),
  .ZN({ S3426 })
);
OAI21_X1 #() 
OAI21_X1_2751_ (
  .A({ S25957[773] }),
  .B1({ S3424 }),
  .B2({ S3426 }),
  .ZN({ S3427 })
);
NAND3_X1 #() 
NAND3_X1_5742_ (
  .A1({ S2939 }),
  .A2({ S25957[771] }),
  .A3({ S25957[769] }),
  .ZN({ S3428 })
);
OAI211_X1 #() 
OAI211_X1_1883_ (
  .A({ S3428 }),
  .B({ S25957[772] }),
  .C1({ S3070 }),
  .C2({ S25957[771] }),
  .ZN({ S3429 })
);
NOR3_X1 #() 
NOR3_X1_169_ (
  .A1({ S2904 }),
  .A2({ S2903 }),
  .A3({ S25957[768] }),
  .ZN({ S3430 })
);
AOI21_X1 #() 
AOI21_X1_2990_ (
  .A({ S25957[772] }),
  .B1({ S3430 }),
  .B2({ S2917 }),
  .ZN({ S3431 })
);
NAND2_X1 #() 
NAND2_X1_5303_ (
  .A1({ S3431 }),
  .A2({ S2972 }),
  .ZN({ S3432 })
);
NAND3_X1 #() 
NAND3_X1_5743_ (
  .A1({ S3432 }),
  .A2({ S3429 }),
  .A3({ S2927 }),
  .ZN({ S3433 })
);
NAND3_X1 #() 
NAND3_X1_5744_ (
  .A1({ S3427 }),
  .A2({ S2900 }),
  .A3({ S3433 }),
  .ZN({ S3434 })
);
NAND3_X1 #() 
NAND3_X1_5745_ (
  .A1({ S3434 }),
  .A2({ S3421 }),
  .A3({ S25957[775] }),
  .ZN({ S3435 })
);
NAND3_X1 #() 
NAND3_X1_5746_ (
  .A1({ S3077 }),
  .A2({ S2910 }),
  .A3({ S25957[771] }),
  .ZN({ S3436 })
);
NAND2_X1 #() 
NAND2_X1_5304_ (
  .A1({ S2999 }),
  .A2({ S104 }),
  .ZN({ S3437 })
);
OAI211_X1 #() 
OAI211_X1_1884_ (
  .A({ S3436 }),
  .B({ S25957[772] }),
  .C1({ S3437 }),
  .C2({ S3022 }),
  .ZN({ S3438 })
);
NAND3_X1 #() 
NAND3_X1_5747_ (
  .A1({ S3180 }),
  .A2({ S2901 }),
  .A3({ S3428 }),
  .ZN({ S3439 })
);
NAND3_X1 #() 
NAND3_X1_5748_ (
  .A1({ S3438 }),
  .A2({ S2927 }),
  .A3({ S3439 }),
  .ZN({ S3440 })
);
AND3_X1 #() 
AND3_X1_227_ (
  .A1({ S3006 }),
  .A2({ S2912 }),
  .A3({ S25957[771] }),
  .ZN({ S3441 })
);
OAI21_X1 #() 
OAI21_X1_2752_ (
  .A({ S25957[772] }),
  .B1({ S3441 }),
  .B2({ S3240 }),
  .ZN({ S3442 })
);
AOI21_X1 #() 
AOI21_X1_2991_ (
  .A({ S25957[772] }),
  .B1({ S2976 }),
  .B2({ S3027 }),
  .ZN({ S3443 })
);
NAND2_X1 #() 
NAND2_X1_5305_ (
  .A1({ S2938 }),
  .A2({ S3443 }),
  .ZN({ S3444 })
);
NAND3_X1 #() 
NAND3_X1_5749_ (
  .A1({ S3442 }),
  .A2({ S25957[773] }),
  .A3({ S3444 }),
  .ZN({ S3445 })
);
AND3_X1 #() 
AND3_X1_228_ (
  .A1({ S3445 }),
  .A2({ S3440 }),
  .A3({ S25957[774] }),
  .ZN({ S3446 })
);
NAND3_X1 #() 
NAND3_X1_5750_ (
  .A1({ S2955 }),
  .A2({ S2948 }),
  .A3({ S25957[771] }),
  .ZN({ S3447 })
);
NAND3_X1 #() 
NAND3_X1_5751_ (
  .A1({ S3225 }),
  .A2({ S3447 }),
  .A3({ S25957[772] }),
  .ZN({ S3448 })
);
NAND3_X1 #() 
NAND3_X1_5752_ (
  .A1({ S3041 }),
  .A2({ S2999 }),
  .A3({ S25957[771] }),
  .ZN({ S3449 })
);
AOI21_X1 #() 
AOI21_X1_2992_ (
  .A({ S2927 }),
  .B1({ S3431 }),
  .B2({ S3449 }),
  .ZN({ S3450 })
);
NAND2_X1 #() 
NAND2_X1_5306_ (
  .A1({ S3450 }),
  .A2({ S3448 }),
  .ZN({ S3451 })
);
AOI21_X1 #() 
AOI21_X1_2993_ (
  .A({ S2901 }),
  .B1({ S3186 }),
  .B2({ S3428 }),
  .ZN({ S3452 })
);
NAND2_X1 #() 
NAND2_X1_5307_ (
  .A1({ S2912 }),
  .A2({ S2936 }),
  .ZN({ S3453 })
);
AOI21_X1 #() 
AOI21_X1_2994_ (
  .A({ S25957[772] }),
  .B1({ S3453 }),
  .B2({ S2911 }),
  .ZN({ S3454 })
);
NAND2_X1 #() 
NAND2_X1_5308_ (
  .A1({ S3454 }),
  .A2({ S3001 }),
  .ZN({ S3455 })
);
NAND2_X1 #() 
NAND2_X1_5309_ (
  .A1({ S3079 }),
  .A2({ S3455 }),
  .ZN({ S3456 })
);
OAI21_X1 #() 
OAI21_X1_2753_ (
  .A({ S2927 }),
  .B1({ S3456 }),
  .B2({ S3452 }),
  .ZN({ S3457 })
);
AOI21_X1 #() 
AOI21_X1_2995_ (
  .A({ S25957[774] }),
  .B1({ S3457 }),
  .B2({ S3451 }),
  .ZN({ S3458 })
);
OAI21_X1 #() 
OAI21_X1_2754_ (
  .A({ S2962 }),
  .B1({ S3458 }),
  .B2({ S3446 }),
  .ZN({ S3459 })
);
AOI21_X1 #() 
AOI21_X1_2996_ (
  .A({ S3412 }),
  .B1({ S3459 }),
  .B2({ S3435 }),
  .ZN({ S3460 })
);
AND3_X1 #() 
AND3_X1_229_ (
  .A1({ S3434 }),
  .A2({ S3421 }),
  .A3({ S25957[775] }),
  .ZN({ S3461 })
);
NAND3_X1 #() 
NAND3_X1_5753_ (
  .A1({ S3445 }),
  .A2({ S3440 }),
  .A3({ S25957[774] }),
  .ZN({ S3462 })
);
AND2_X1 #() 
AND2_X1_340_ (
  .A1({ S3450 }),
  .A2({ S3448 }),
  .ZN({ S3463 })
);
AOI21_X1 #() 
AOI21_X1_2997_ (
  .A({ S25957[771] }),
  .B1({ S2999 }),
  .B2({ S3047 }),
  .ZN({ S3464 })
);
AOI21_X1 #() 
AOI21_X1_2998_ (
  .A({ S104 }),
  .B1({ S2933 }),
  .B2({ S2936 }),
  .ZN({ S3465 })
);
OAI21_X1 #() 
OAI21_X1_2755_ (
  .A({ S25957[772] }),
  .B1({ S3464 }),
  .B2({ S3465 }),
  .ZN({ S3466 })
);
OAI21_X1 #() 
OAI21_X1_2756_ (
  .A({ S3287 }),
  .B1({ S3285 }),
  .B2({ S2936 }),
  .ZN({ S3467 })
);
AOI22_X1 #() 
AOI22_X1_602_ (
  .A1({ S3467 }),
  .A2({ S2901 }),
  .B1({ S3454 }),
  .B2({ S3001 }),
  .ZN({ S3468 })
);
AOI21_X1 #() 
AOI21_X1_2999_ (
  .A({ S25957[773] }),
  .B1({ S3468 }),
  .B2({ S3466 }),
  .ZN({ S3469 })
);
OAI21_X1 #() 
OAI21_X1_2757_ (
  .A({ S2900 }),
  .B1({ S3469 }),
  .B2({ S3463 }),
  .ZN({ S3470 })
);
AOI21_X1 #() 
AOI21_X1_3000_ (
  .A({ S25957[775] }),
  .B1({ S3470 }),
  .B2({ S3462 }),
  .ZN({ S3471 })
);
NOR3_X1 #() 
NOR3_X1_170_ (
  .A1({ S3471 }),
  .A2({ S3461 }),
  .A3({ S25957[970] }),
  .ZN({ S3472 })
);
OAI21_X1 #() 
OAI21_X1_2758_ (
  .A({ S25957[810] }),
  .B1({ S3472 }),
  .B2({ S3460 }),
  .ZN({ S3473 })
);
OAI21_X1 #() 
OAI21_X1_2759_ (
  .A({ S25957[970] }),
  .B1({ S3471 }),
  .B2({ S3461 }),
  .ZN({ S3474 })
);
NAND3_X1 #() 
NAND3_X1_5754_ (
  .A1({ S3459 }),
  .A2({ S3412 }),
  .A3({ S3435 }),
  .ZN({ S3475 })
);
NAND3_X1 #() 
NAND3_X1_5755_ (
  .A1({ S3474 }),
  .A2({ S3411 }),
  .A3({ S3475 }),
  .ZN({ S3476 })
);
NAND3_X1 #() 
NAND3_X1_5756_ (
  .A1({ S3473 }),
  .A2({ S2243 }),
  .A3({ S3476 }),
  .ZN({ S3477 })
);
OAI21_X1 #() 
OAI21_X1_2760_ (
  .A({ S3411 }),
  .B1({ S3472 }),
  .B2({ S3460 }),
  .ZN({ S3478 })
);
NAND3_X1 #() 
NAND3_X1_5757_ (
  .A1({ S3474 }),
  .A2({ S25957[810] }),
  .A3({ S3475 }),
  .ZN({ S3479 })
);
NAND3_X1 #() 
NAND3_X1_5758_ (
  .A1({ S3478 }),
  .A2({ S25957[778] }),
  .A3({ S3479 }),
  .ZN({ S3480 })
);
NAND2_X1 #() 
NAND2_X1_5310_ (
  .A1({ S3477 }),
  .A2({ S3480 }),
  .ZN({ S25957[650] })
);
NOR2_X1 #() 
NOR2_X1_1334_ (
  .A1({ S2067 }),
  .A2({ S2066 }),
  .ZN({ S3481 })
);
AOI21_X1 #() 
AOI21_X1_3001_ (
  .A({ S3481 }),
  .B1({ S2140 }),
  .B2({ S2143 }),
  .ZN({ S114 })
);
NAND3_X1 #() 
NAND3_X1_5759_ (
  .A1({ S2140 }),
  .A2({ S3481 }),
  .A3({ S2143 }),
  .ZN({ S115 })
);
INV_X1 #() 
INV_X1_1735_ (
  .A({ S1141 }),
  .ZN({ S25957[807] })
);
XNOR2_X1 #() 
XNOR2_X1_205_ (
  .A({ S24131 }),
  .B({ S25957[1223] }),
  .ZN({ S25957[967] })
);
XNOR2_X1 #() 
XNOR2_X1_206_ (
  .A({ S1137 }),
  .B({ S25957[967] }),
  .ZN({ S25957[839] })
);
INV_X1 #() 
INV_X1_1736_ (
  .A({ S1137 }),
  .ZN({ S25957[871] })
);
INV_X1 #() 
INV_X1_1737_ (
  .A({ S25957[797] }),
  .ZN({ S3482 })
);
NAND2_X1 #() 
NAND2_X1_5311_ (
  .A1({ S1946 }),
  .A2({ S1949 }),
  .ZN({ S3483 })
);
NAND3_X1 #() 
NAND3_X1_5760_ (
  .A1({ S2140 }),
  .A2({ S25957[792] }),
  .A3({ S2143 }),
  .ZN({ S3484 })
);
INV_X1 #() 
INV_X1_1738_ (
  .A({ S3484 }),
  .ZN({ S3485 })
);
NAND3_X1 #() 
NAND3_X1_5761_ (
  .A1({ S2228 }),
  .A2({ S2229 }),
  .A3({ S25957[922] }),
  .ZN({ S3486 })
);
NAND3_X1 #() 
NAND3_X1_5762_ (
  .A1({ S2223 }),
  .A2({ S2226 }),
  .A3({ S1033 }),
  .ZN({ S3487 })
);
NAND2_X1 #() 
NAND2_X1_5312_ (
  .A1({ S3486 }),
  .A2({ S3487 }),
  .ZN({ S3488 })
);
NAND3_X1 #() 
NAND3_X1_5763_ (
  .A1({ S2141 }),
  .A2({ S2142 }),
  .A3({ S25957[921] }),
  .ZN({ S3489 })
);
OAI21_X1 #() 
OAI21_X1_2761_ (
  .A({ S1019 }),
  .B1({ S2136 }),
  .B2({ S2139 }),
  .ZN({ S3490 })
);
NAND3_X1 #() 
NAND3_X1_5764_ (
  .A1({ S3490 }),
  .A2({ S3481 }),
  .A3({ S3489 }),
  .ZN({ S3491 })
);
NOR2_X1 #() 
NOR2_X1_1335_ (
  .A1({ S3491 }),
  .A2({ S3488 }),
  .ZN({ S3492 })
);
OAI21_X1 #() 
OAI21_X1_2762_ (
  .A({ S25957[795] }),
  .B1({ S3492 }),
  .B2({ S3485 }),
  .ZN({ S3493 })
);
AOI22_X1 #() 
AOI22_X1_603_ (
  .A1({ S3490 }),
  .A2({ S3489 }),
  .B1({ S3486 }),
  .B2({ S3487 }),
  .ZN({ S3494 })
);
NAND3_X1 #() 
NAND3_X1_5765_ (
  .A1({ S25957[792] }),
  .A2({ S3486 }),
  .A3({ S3487 }),
  .ZN({ S3495 })
);
NAND2_X1 #() 
NAND2_X1_5313_ (
  .A1({ S3491 }),
  .A2({ S3495 }),
  .ZN({ S3496 })
);
NOR2_X1 #() 
NOR2_X1_1336_ (
  .A1({ S3496 }),
  .A2({ S3494 }),
  .ZN({ S3497 })
);
NAND2_X1 #() 
NAND2_X1_5314_ (
  .A1({ S3497 }),
  .A2({ S107 }),
  .ZN({ S3498 })
);
NAND3_X1 #() 
NAND3_X1_5766_ (
  .A1({ S3498 }),
  .A2({ S3483 }),
  .A3({ S3493 }),
  .ZN({ S3499 })
);
NAND3_X1 #() 
NAND3_X1_5767_ (
  .A1({ S3484 }),
  .A2({ S25957[795] }),
  .A3({ S3488 }),
  .ZN({ S3500 })
);
NAND2_X1 #() 
NAND2_X1_5315_ (
  .A1({ S3500 }),
  .A2({ S25957[796] }),
  .ZN({ S3501 })
);
NAND3_X1 #() 
NAND3_X1_5768_ (
  .A1({ S2227 }),
  .A2({ S2230 }),
  .A3({ S3481 }),
  .ZN({ S3502 })
);
INV_X1 #() 
INV_X1_1739_ (
  .A({ S3502 }),
  .ZN({ S3503 })
);
NAND3_X1 #() 
NAND3_X1_5769_ (
  .A1({ S3490 }),
  .A2({ S107 }),
  .A3({ S3489 }),
  .ZN({ S3504 })
);
AOI21_X1 #() 
AOI21_X1_3002_ (
  .A({ S3481 }),
  .B1({ S2227 }),
  .B2({ S2230 }),
  .ZN({ S3505 })
);
NAND2_X1 #() 
NAND2_X1_5316_ (
  .A1({ S3505 }),
  .A2({ S25957[795] }),
  .ZN({ S3506 })
);
OAI21_X1 #() 
OAI21_X1_2763_ (
  .A({ S3506 }),
  .B1({ S3503 }),
  .B2({ S3504 }),
  .ZN({ S3507 })
);
OAI21_X1 #() 
OAI21_X1_2764_ (
  .A({ S3499 }),
  .B1({ S3501 }),
  .B2({ S3507 }),
  .ZN({ S3508 })
);
NAND4_X1 #() 
NAND4_X1_621_ (
  .A1({ S2140 }),
  .A2({ S2143 }),
  .A3({ S3486 }),
  .A4({ S3487 }),
  .ZN({ S3509 })
);
INV_X1 #() 
INV_X1_1740_ (
  .A({ S3509 }),
  .ZN({ S3510 })
);
NAND3_X1 #() 
NAND3_X1_5770_ (
  .A1({ S3490 }),
  .A2({ S25957[792] }),
  .A3({ S3489 }),
  .ZN({ S3511 })
);
NAND2_X1 #() 
NAND2_X1_5317_ (
  .A1({ S3511 }),
  .A2({ S25957[795] }),
  .ZN({ S3512 })
);
NOR2_X1 #() 
NOR2_X1_1337_ (
  .A1({ S3512 }),
  .A2({ S3510 }),
  .ZN({ S3513 })
);
AOI21_X1 #() 
AOI21_X1_3003_ (
  .A({ S3513 }),
  .B1({ S3491 }),
  .B2({ S107 }),
  .ZN({ S3514 })
);
NAND2_X1 #() 
NAND2_X1_5318_ (
  .A1({ S3514 }),
  .A2({ S25957[796] }),
  .ZN({ S3515 })
);
NAND4_X1 #() 
NAND4_X1_622_ (
  .A1({ S2140 }),
  .A2({ S2143 }),
  .A3({ S2227 }),
  .A4({ S2230 }),
  .ZN({ S3516 })
);
NAND4_X1 #() 
NAND4_X1_623_ (
  .A1({ S3490 }),
  .A2({ S3489 }),
  .A3({ S3486 }),
  .A4({ S3487 }),
  .ZN({ S3517 })
);
OAI211_X1 #() 
OAI211_X1_1885_ (
  .A({ S3517 }),
  .B({ S3495 }),
  .C1({ S3516 }),
  .C2({ S25957[792] }),
  .ZN({ S3518 })
);
NOR2_X1 #() 
NOR2_X1_1338_ (
  .A1({ S3484 }),
  .A2({ S107 }),
  .ZN({ S3519 })
);
OAI21_X1 #() 
OAI21_X1_2765_ (
  .A({ S3483 }),
  .B1({ S3518 }),
  .B2({ S3519 }),
  .ZN({ S3520 })
);
NAND3_X1 #() 
NAND3_X1_5771_ (
  .A1({ S3515 }),
  .A2({ S3482 }),
  .A3({ S3520 }),
  .ZN({ S3521 })
);
OAI211_X1 #() 
OAI211_X1_1886_ (
  .A({ S3521 }),
  .B({ S25957[798] }),
  .C1({ S3508 }),
  .C2({ S3482 }),
  .ZN({ S3522 })
);
INV_X1 #() 
INV_X1_1741_ (
  .A({ S25957[798] }),
  .ZN({ S3523 })
);
AOI21_X1 #() 
AOI21_X1_3004_ (
  .A({ S25957[792] }),
  .B1({ S3490 }),
  .B2({ S3489 }),
  .ZN({ S3524 })
);
NAND2_X1 #() 
NAND2_X1_5319_ (
  .A1({ S3524 }),
  .A2({ S3488 }),
  .ZN({ S3525 })
);
AND2_X1 #() 
AND2_X1_341_ (
  .A1({ S3525 }),
  .A2({ S3512 }),
  .ZN({ S3526 })
);
NAND2_X1 #() 
NAND2_X1_5320_ (
  .A1({ S3490 }),
  .A2({ S3489 }),
  .ZN({ S3527 })
);
NAND2_X1 #() 
NAND2_X1_5321_ (
  .A1({ S3527 }),
  .A2({ S25957[795] }),
  .ZN({ S3528 })
);
AND3_X1 #() 
AND3_X1_230_ (
  .A1({ S3506 }),
  .A2({ S3528 }),
  .A3({ S25957[796] }),
  .ZN({ S3529 })
);
OAI21_X1 #() 
OAI21_X1_2766_ (
  .A({ S3529 }),
  .B1({ S3505 }),
  .B2({ S3504 }),
  .ZN({ S3530 })
);
OAI21_X1 #() 
OAI21_X1_2767_ (
  .A({ S3530 }),
  .B1({ S25957[796] }),
  .B2({ S3526 }),
  .ZN({ S3531 })
);
INV_X1 #() 
INV_X1_1742_ (
  .A({ S3517 }),
  .ZN({ S3532 })
);
AOI21_X1 #() 
AOI21_X1_3005_ (
  .A({ S3488 }),
  .B1({ S3484 }),
  .B2({ S3491 }),
  .ZN({ S3533 })
);
AOI21_X1 #() 
AOI21_X1_3006_ (
  .A({ S25957[794] }),
  .B1({ S3511 }),
  .B2({ S115 }),
  .ZN({ S3534 })
);
OAI21_X1 #() 
OAI21_X1_2768_ (
  .A({ S25957[795] }),
  .B1({ S3533 }),
  .B2({ S3534 }),
  .ZN({ S3535 })
);
NAND3_X1 #() 
NAND3_X1_5772_ (
  .A1({ S25957[792] }),
  .A2({ S2227 }),
  .A3({ S2230 }),
  .ZN({ S3536 })
);
NAND2_X1 #() 
NAND2_X1_5322_ (
  .A1({ S3536 }),
  .A2({ S107 }),
  .ZN({ S3537 })
);
OAI21_X1 #() 
OAI21_X1_2769_ (
  .A({ S3535 }),
  .B1({ S3532 }),
  .B2({ S3537 }),
  .ZN({ S3538 })
);
NAND3_X1 #() 
NAND3_X1_5773_ (
  .A1({ S3511 }),
  .A2({ S115 }),
  .A3({ S3488 }),
  .ZN({ S3539 })
);
AOI21_X1 #() 
AOI21_X1_3007_ (
  .A({ S25957[795] }),
  .B1({ S3539 }),
  .B2({ S3517 }),
  .ZN({ S3540 })
);
NOR2_X1 #() 
NOR2_X1_1339_ (
  .A1({ S3516 }),
  .A2({ S107 }),
  .ZN({ S3541 })
);
AOI21_X1 #() 
AOI21_X1_3008_ (
  .A({ S25957[792] }),
  .B1({ S2227 }),
  .B2({ S2230 }),
  .ZN({ S3542 })
);
NOR2_X1 #() 
NOR2_X1_1340_ (
  .A1({ S3542 }),
  .A2({ S25957[795] }),
  .ZN({ S3543 })
);
OAI21_X1 #() 
OAI21_X1_2770_ (
  .A({ S3483 }),
  .B1({ S3541 }),
  .B2({ S3543 }),
  .ZN({ S3544 })
);
OAI221_X1 #() 
OAI221_X1_160_ (
  .A({ S3482 }),
  .B1({ S3540 }),
  .B2({ S3544 }),
  .C1({ S3538 }),
  .C2({ S3483 }),
  .ZN({ S3545 })
);
OAI211_X1 #() 
OAI211_X1_1887_ (
  .A({ S3545 }),
  .B({ S3523 }),
  .C1({ S3482 }),
  .C2({ S3531 }),
  .ZN({ S3546 })
);
NAND3_X1 #() 
NAND3_X1_5774_ (
  .A1({ S3546 }),
  .A2({ S25957[799] }),
  .A3({ S3522 }),
  .ZN({ S3547 })
);
INV_X1 #() 
INV_X1_1743_ (
  .A({ S3547 }),
  .ZN({ S3548 })
);
NOR2_X1 #() 
NOR2_X1_1341_ (
  .A1({ S3497 }),
  .A2({ S107 }),
  .ZN({ S3549 })
);
NAND2_X1 #() 
NAND2_X1_5323_ (
  .A1({ S3502 }),
  .A2({ S107 }),
  .ZN({ S3550 })
);
OAI21_X1 #() 
OAI21_X1_2771_ (
  .A({ S25957[796] }),
  .B1({ S3492 }),
  .B2({ S3550 }),
  .ZN({ S3551 })
);
NAND2_X1 #() 
NAND2_X1_5324_ (
  .A1({ S3484 }),
  .A2({ S3488 }),
  .ZN({ S3552 })
);
AOI21_X1 #() 
AOI21_X1_3009_ (
  .A({ S107 }),
  .B1({ S3527 }),
  .B2({ S25957[794] }),
  .ZN({ S3553 })
);
NAND2_X1 #() 
NAND2_X1_5325_ (
  .A1({ S3553 }),
  .A2({ S3552 }),
  .ZN({ S3554 })
);
NAND3_X1 #() 
NAND3_X1_5775_ (
  .A1({ S3486 }),
  .A2({ S3487 }),
  .A3({ S3481 }),
  .ZN({ S3555 })
);
NAND3_X1 #() 
NAND3_X1_5776_ (
  .A1({ S3509 }),
  .A2({ S107 }),
  .A3({ S3555 }),
  .ZN({ S3556 })
);
NAND3_X1 #() 
NAND3_X1_5777_ (
  .A1({ S3554 }),
  .A2({ S3483 }),
  .A3({ S3556 }),
  .ZN({ S3557 })
);
OAI211_X1 #() 
OAI211_X1_1888_ (
  .A({ S25957[797] }),
  .B({ S3557 }),
  .C1({ S3549 }),
  .C2({ S3551 }),
  .ZN({ S3558 })
);
NAND4_X1 #() 
NAND4_X1_624_ (
  .A1({ S3490 }),
  .A2({ S3489 }),
  .A3({ S2227 }),
  .A4({ S2230 }),
  .ZN({ S3559 })
);
NOR2_X1 #() 
NOR2_X1_1342_ (
  .A1({ S3505 }),
  .A2({ S107 }),
  .ZN({ S3560 })
);
NAND2_X1 #() 
NAND2_X1_5326_ (
  .A1({ S3560 }),
  .A2({ S3559 }),
  .ZN({ S3561 })
);
NAND4_X1 #() 
NAND4_X1_625_ (
  .A1({ S3559 }),
  .A2({ S3509 }),
  .A3({ S3502 }),
  .A4({ S3555 }),
  .ZN({ S3562 })
);
AOI21_X1 #() 
AOI21_X1_3010_ (
  .A({ S25957[796] }),
  .B1({ S3562 }),
  .B2({ S107 }),
  .ZN({ S3563 })
);
NAND3_X1 #() 
NAND3_X1_5778_ (
  .A1({ S3511 }),
  .A2({ S115 }),
  .A3({ S25957[794] }),
  .ZN({ S3564 })
);
AOI21_X1 #() 
AOI21_X1_3011_ (
  .A({ S25957[795] }),
  .B1({ S3488 }),
  .B2({ S25957[792] }),
  .ZN({ S3565 })
);
NAND2_X1 #() 
NAND2_X1_5327_ (
  .A1({ S3564 }),
  .A2({ S3565 }),
  .ZN({ S3566 })
);
NAND2_X1 #() 
NAND2_X1_5328_ (
  .A1({ S3511 }),
  .A2({ S25957[794] }),
  .ZN({ S3567 })
);
NAND3_X1 #() 
NAND3_X1_5779_ (
  .A1({ S3484 }),
  .A2({ S3491 }),
  .A3({ S3488 }),
  .ZN({ S3568 })
);
AOI21_X1 #() 
AOI21_X1_3012_ (
  .A({ S107 }),
  .B1({ S3568 }),
  .B2({ S3567 }),
  .ZN({ S3569 })
);
NOR2_X1 #() 
NOR2_X1_1343_ (
  .A1({ S3569 }),
  .A2({ S3483 }),
  .ZN({ S3570 })
);
AOI22_X1 #() 
AOI22_X1_604_ (
  .A1({ S3570 }),
  .A2({ S3566 }),
  .B1({ S3563 }),
  .B2({ S3561 }),
  .ZN({ S3571 })
);
OAI211_X1 #() 
OAI211_X1_1889_ (
  .A({ S25957[798] }),
  .B({ S3558 }),
  .C1({ S3571 }),
  .C2({ S25957[797] }),
  .ZN({ S3572 })
);
NAND2_X1 #() 
NAND2_X1_5329_ (
  .A1({ S3560 }),
  .A2({ S3516 }),
  .ZN({ S3573 })
);
OAI21_X1 #() 
OAI21_X1_2772_ (
  .A({ S3573 }),
  .B1({ S25957[795] }),
  .B2({ S3481 }),
  .ZN({ S3574 })
);
NAND2_X1 #() 
NAND2_X1_5330_ (
  .A1({ S3511 }),
  .A2({ S3488 }),
  .ZN({ S3575 })
);
INV_X1 #() 
INV_X1_1744_ (
  .A({ S3575 }),
  .ZN({ S3576 })
);
NAND2_X1 #() 
NAND2_X1_5331_ (
  .A1({ S3517 }),
  .A2({ S107 }),
  .ZN({ S3577 })
);
NAND3_X1 #() 
NAND3_X1_5780_ (
  .A1({ S3559 }),
  .A2({ S25957[795] }),
  .A3({ S3484 }),
  .ZN({ S3578 })
);
OAI21_X1 #() 
OAI21_X1_2773_ (
  .A({ S3578 }),
  .B1({ S3576 }),
  .B2({ S3577 }),
  .ZN({ S3579 })
);
NAND2_X1 #() 
NAND2_X1_5332_ (
  .A1({ S3579 }),
  .A2({ S3483 }),
  .ZN({ S3580 })
);
OAI211_X1 #() 
OAI211_X1_1890_ (
  .A({ S3580 }),
  .B({ S25957[797] }),
  .C1({ S3483 }),
  .C2({ S3574 }),
  .ZN({ S3581 })
);
NOR2_X1 #() 
NOR2_X1_1344_ (
  .A1({ S3511 }),
  .A2({ S25957[794] }),
  .ZN({ S3582 })
);
NAND2_X1 #() 
NAND2_X1_5333_ (
  .A1({ S3564 }),
  .A2({ S107 }),
  .ZN({ S3583 })
);
OAI221_X1 #() 
OAI221_X1_161_ (
  .A({ S25957[796] }),
  .B1({ S3492 }),
  .B2({ S107 }),
  .C1({ S3583 }),
  .C2({ S3582 }),
  .ZN({ S3584 })
);
NAND4_X1 #() 
NAND4_X1_626_ (
  .A1({ S3484 }),
  .A2({ S3491 }),
  .A3({ S107 }),
  .A4({ S25957[794] }),
  .ZN({ S3585 })
);
AOI21_X1 #() 
AOI21_X1_3013_ (
  .A({ S107 }),
  .B1({ S2227 }),
  .B2({ S2230 }),
  .ZN({ S3586 })
);
NAND2_X1 #() 
NAND2_X1_5334_ (
  .A1({ S3586 }),
  .A2({ S3511 }),
  .ZN({ S3587 })
);
NAND3_X1 #() 
NAND3_X1_5781_ (
  .A1({ S3585 }),
  .A2({ S3483 }),
  .A3({ S3587 }),
  .ZN({ S3588 })
);
NAND3_X1 #() 
NAND3_X1_5782_ (
  .A1({ S3584 }),
  .A2({ S3482 }),
  .A3({ S3588 }),
  .ZN({ S3589 })
);
NAND3_X1 #() 
NAND3_X1_5783_ (
  .A1({ S3589 }),
  .A2({ S3581 }),
  .A3({ S3523 }),
  .ZN({ S3590 })
);
AOI21_X1 #() 
AOI21_X1_3014_ (
  .A({ S25957[799] }),
  .B1({ S3572 }),
  .B2({ S3590 }),
  .ZN({ S3591 })
);
OR3_X1 #() 
OR3_X1_34_ (
  .A1({ S3548 }),
  .A2({ S3591 }),
  .A3({ S25957[871] }),
  .ZN({ S3592 })
);
OAI21_X1 #() 
OAI21_X1_2774_ (
  .A({ S25957[871] }),
  .B1({ S3548 }),
  .B2({ S3591 }),
  .ZN({ S3593 })
);
NAND2_X1 #() 
NAND2_X1_5335_ (
  .A1({ S3592 }),
  .A2({ S3593 }),
  .ZN({ S25957[743] })
);
NAND2_X1 #() 
NAND2_X1_5336_ (
  .A1({ S25957[743] }),
  .A2({ S25957[839] }),
  .ZN({ S3594 })
);
INV_X1 #() 
INV_X1_1745_ (
  .A({ S25957[839] }),
  .ZN({ S3595 })
);
NAND3_X1 #() 
NAND3_X1_5784_ (
  .A1({ S3592 }),
  .A2({ S3595 }),
  .A3({ S3593 }),
  .ZN({ S3596 })
);
NAND3_X1 #() 
NAND3_X1_5785_ (
  .A1({ S3594 }),
  .A2({ S25957[807] }),
  .A3({ S3596 }),
  .ZN({ S3597 })
);
NAND2_X1 #() 
NAND2_X1_5337_ (
  .A1({ S25957[743] }),
  .A2({ S3595 }),
  .ZN({ S3598 })
);
NAND3_X1 #() 
NAND3_X1_5786_ (
  .A1({ S3592 }),
  .A2({ S25957[839] }),
  .A3({ S3593 }),
  .ZN({ S3599 })
);
NAND3_X1 #() 
NAND3_X1_5787_ (
  .A1({ S3598 }),
  .A2({ S1141 }),
  .A3({ S3599 }),
  .ZN({ S3600 })
);
NAND3_X1 #() 
NAND3_X1_5788_ (
  .A1({ S3597 }),
  .A2({ S3600 }),
  .A3({ S2962 }),
  .ZN({ S3601 })
);
NAND3_X1 #() 
NAND3_X1_5789_ (
  .A1({ S3594 }),
  .A2({ S1141 }),
  .A3({ S3596 }),
  .ZN({ S3602 })
);
NAND3_X1 #() 
NAND3_X1_5790_ (
  .A1({ S3598 }),
  .A2({ S25957[807] }),
  .A3({ S3599 }),
  .ZN({ S3603 })
);
NAND3_X1 #() 
NAND3_X1_5791_ (
  .A1({ S3602 }),
  .A2({ S3603 }),
  .A3({ S25957[775] }),
  .ZN({ S3604 })
);
NAND2_X1 #() 
NAND2_X1_5338_ (
  .A1({ S3601 }),
  .A2({ S3604 }),
  .ZN({ S25957[647] })
);
INV_X1 #() 
INV_X1_1746_ (
  .A({ S1214 }),
  .ZN({ S3605 })
);
INV_X1 #() 
INV_X1_1747_ (
  .A({ S1218 }),
  .ZN({ S3606 })
);
NOR2_X1 #() 
NOR2_X1_1345_ (
  .A1({ S3606 }),
  .A2({ S3605 }),
  .ZN({ S25957[806] })
);
NAND2_X1 #() 
NAND2_X1_5339_ (
  .A1({ S3511 }),
  .A2({ S115 }),
  .ZN({ S3607 })
);
INV_X1 #() 
INV_X1_1748_ (
  .A({ S3607 }),
  .ZN({ S3608 })
);
NAND2_X1 #() 
NAND2_X1_5340_ (
  .A1({ S3559 }),
  .A2({ S107 }),
  .ZN({ S3609 })
);
NAND3_X1 #() 
NAND3_X1_5792_ (
  .A1({ S25957[793] }),
  .A2({ S3481 }),
  .A3({ S3488 }),
  .ZN({ S3610 })
);
NAND2_X1 #() 
NAND2_X1_5341_ (
  .A1({ S3610 }),
  .A2({ S25957[795] }),
  .ZN({ S3611 })
);
OAI221_X1 #() 
OAI221_X1_162_ (
  .A({ S3483 }),
  .B1({ S3608 }),
  .B2({ S3609 }),
  .C1({ S3611 }),
  .C2({ S3510 }),
  .ZN({ S3612 })
);
NAND2_X1 #() 
NAND2_X1_5342_ (
  .A1({ S3586 }),
  .A2({ S25957[793] }),
  .ZN({ S3613 })
);
INV_X1 #() 
INV_X1_1749_ (
  .A({ S3504 }),
  .ZN({ S3614 })
);
NAND2_X1 #() 
NAND2_X1_5343_ (
  .A1({ S3614 }),
  .A2({ S3503 }),
  .ZN({ S3615 })
);
NAND3_X1 #() 
NAND3_X1_5793_ (
  .A1({ S3615 }),
  .A2({ S3585 }),
  .A3({ S3613 }),
  .ZN({ S3616 })
);
AOI21_X1 #() 
AOI21_X1_3015_ (
  .A({ S3482 }),
  .B1({ S3616 }),
  .B2({ S25957[796] }),
  .ZN({ S3617 })
);
AOI21_X1 #() 
AOI21_X1_3016_ (
  .A({ S25957[794] }),
  .B1({ S3484 }),
  .B2({ S3491 }),
  .ZN({ S3618 })
);
NOR2_X1 #() 
NOR2_X1_1346_ (
  .A1({ S3495 }),
  .A2({ S25957[795] }),
  .ZN({ S3619 })
);
AOI21_X1 #() 
AOI21_X1_3017_ (
  .A({ S3619 }),
  .B1({ S3618 }),
  .B2({ S107 }),
  .ZN({ S3620 })
);
NAND2_X1 #() 
NAND2_X1_5344_ (
  .A1({ S3517 }),
  .A2({ S3481 }),
  .ZN({ S3621 })
);
NAND3_X1 #() 
NAND3_X1_5794_ (
  .A1({ S3621 }),
  .A2({ S25957[795] }),
  .A3({ S3495 }),
  .ZN({ S3622 })
);
AOI21_X1 #() 
AOI21_X1_3018_ (
  .A({ S25957[796] }),
  .B1({ S3620 }),
  .B2({ S3622 }),
  .ZN({ S3623 })
);
NAND2_X1 #() 
NAND2_X1_5345_ (
  .A1({ S3559 }),
  .A2({ S3502 }),
  .ZN({ S3624 })
);
NAND2_X1 #() 
NAND2_X1_5346_ (
  .A1({ S3624 }),
  .A2({ S107 }),
  .ZN({ S3625 })
);
AOI21_X1 #() 
AOI21_X1_3019_ (
  .A({ S3623 }),
  .B1({ S3529 }),
  .B2({ S3625 }),
  .ZN({ S3626 })
);
AOI22_X1 #() 
AOI22_X1_605_ (
  .A1({ S3626 }),
  .A2({ S3482 }),
  .B1({ S3612 }),
  .B2({ S3617 }),
  .ZN({ S3627 })
);
AOI21_X1 #() 
AOI21_X1_3020_ (
  .A({ S107 }),
  .B1({ S3511 }),
  .B2({ S3488 }),
  .ZN({ S3628 })
);
NAND2_X1 #() 
NAND2_X1_5347_ (
  .A1({ S3628 }),
  .A2({ S115 }),
  .ZN({ S3629 })
);
NAND2_X1 #() 
NAND2_X1_5348_ (
  .A1({ S3484 }),
  .A2({ S25957[794] }),
  .ZN({ S3630 })
);
AOI21_X1 #() 
AOI21_X1_3021_ (
  .A({ S107 }),
  .B1({ S3630 }),
  .B2({ S3536 }),
  .ZN({ S3631 })
);
NOR2_X1 #() 
NOR2_X1_1347_ (
  .A1({ S3631 }),
  .A2({ S3483 }),
  .ZN({ S3632 })
);
AOI22_X1 #() 
AOI22_X1_606_ (
  .A1({ S3632 }),
  .A2({ S3620 }),
  .B1({ S3563 }),
  .B2({ S3629 }),
  .ZN({ S3633 })
);
NAND2_X1 #() 
NAND2_X1_5349_ (
  .A1({ S115 }),
  .A2({ S25957[794] }),
  .ZN({ S3634 })
);
NAND4_X1 #() 
NAND4_X1_627_ (
  .A1({ S3536 }),
  .A2({ S3555 }),
  .A3({ S3527 }),
  .A4({ S25957[795] }),
  .ZN({ S3635 })
);
OAI211_X1 #() 
OAI211_X1_1891_ (
  .A({ S3635 }),
  .B({ S25957[796] }),
  .C1({ S25957[795] }),
  .C2({ S3634 }),
  .ZN({ S3636 })
);
OAI21_X1 #() 
OAI21_X1_2775_ (
  .A({ S3483 }),
  .B1({ S3513 }),
  .B2({ S3614 }),
  .ZN({ S3637 })
);
NAND3_X1 #() 
NAND3_X1_5795_ (
  .A1({ S3637 }),
  .A2({ S25957[797] }),
  .A3({ S3636 }),
  .ZN({ S3638 })
);
OAI21_X1 #() 
OAI21_X1_2776_ (
  .A({ S3638 }),
  .B1({ S3633 }),
  .B2({ S25957[797] }),
  .ZN({ S3639 })
);
NAND2_X1 #() 
NAND2_X1_5350_ (
  .A1({ S3639 }),
  .A2({ S25957[798] }),
  .ZN({ S3640 })
);
OAI211_X1 #() 
OAI211_X1_1892_ (
  .A({ S3640 }),
  .B({ S25957[799] }),
  .C1({ S25957[798] }),
  .C2({ S3627 }),
  .ZN({ S3641 })
);
INV_X1 #() 
INV_X1_1750_ (
  .A({ S25957[799] }),
  .ZN({ S3642 })
);
NOR2_X1 #() 
NOR2_X1_1348_ (
  .A1({ S3565 }),
  .A2({ S3483 }),
  .ZN({ S3643 })
);
AND3_X1 #() 
AND3_X1_231_ (
  .A1({ S3554 }),
  .A2({ S3643 }),
  .A3({ S3504 }),
  .ZN({ S3644 })
);
NAND2_X1 #() 
NAND2_X1_5351_ (
  .A1({ S3516 }),
  .A2({ S3536 }),
  .ZN({ S3645 })
);
OAI21_X1 #() 
OAI21_X1_2777_ (
  .A({ S25957[795] }),
  .B1({ S3492 }),
  .B2({ S3645 }),
  .ZN({ S3646 })
);
NOR2_X1 #() 
NOR2_X1_1349_ (
  .A1({ S3646 }),
  .A2({ S25957[796] }),
  .ZN({ S3647 })
);
OAI21_X1 #() 
OAI21_X1_2778_ (
  .A({ S3482 }),
  .B1({ S3647 }),
  .B2({ S3644 }),
  .ZN({ S3648 })
);
INV_X1 #() 
INV_X1_1751_ (
  .A({ S3559 }),
  .ZN({ S3649 })
);
INV_X1 #() 
INV_X1_1752_ (
  .A({ S3553 }),
  .ZN({ S3650 })
);
OAI211_X1 #() 
OAI211_X1_1893_ (
  .A({ S3517 }),
  .B({ S107 }),
  .C1({ S3484 }),
  .C2({ S25957[794] }),
  .ZN({ S3651 })
);
OAI21_X1 #() 
OAI21_X1_2779_ (
  .A({ S3651 }),
  .B1({ S3650 }),
  .B2({ S3649 }),
  .ZN({ S3652 })
);
NAND2_X1 #() 
NAND2_X1_5352_ (
  .A1({ S3524 }),
  .A2({ S25957[794] }),
  .ZN({ S3653 })
);
NAND3_X1 #() 
NAND3_X1_5796_ (
  .A1({ S3653 }),
  .A2({ S25957[795] }),
  .A3({ S3511 }),
  .ZN({ S3654 })
);
AOI21_X1 #() 
AOI21_X1_3022_ (
  .A({ S3482 }),
  .B1({ S3654 }),
  .B2({ S3643 }),
  .ZN({ S3655 })
);
OAI21_X1 #() 
OAI21_X1_2780_ (
  .A({ S3655 }),
  .B1({ S25957[796] }),
  .B2({ S3652 }),
  .ZN({ S3656 })
);
NAND3_X1 #() 
NAND3_X1_5797_ (
  .A1({ S3648 }),
  .A2({ S3523 }),
  .A3({ S3656 }),
  .ZN({ S3657 })
);
NAND3_X1 #() 
NAND3_X1_5798_ (
  .A1({ S3517 }),
  .A2({ S3555 }),
  .A3({ S3536 }),
  .ZN({ S3658 })
);
NAND2_X1 #() 
NAND2_X1_5353_ (
  .A1({ S3658 }),
  .A2({ S25957[795] }),
  .ZN({ S3659 })
);
NAND3_X1 #() 
NAND3_X1_5799_ (
  .A1({ S3659 }),
  .A2({ S3583 }),
  .A3({ S3483 }),
  .ZN({ S3660 })
);
NAND2_X1 #() 
NAND2_X1_5354_ (
  .A1({ S3649 }),
  .A2({ S25957[795] }),
  .ZN({ S3661 })
);
NAND3_X1 #() 
NAND3_X1_5800_ (
  .A1({ S3516 }),
  .A2({ S107 }),
  .A3({ S3481 }),
  .ZN({ S3662 })
);
NAND3_X1 #() 
NAND3_X1_5801_ (
  .A1({ S3661 }),
  .A2({ S25957[796] }),
  .A3({ S3662 }),
  .ZN({ S3663 })
);
NAND3_X1 #() 
NAND3_X1_5802_ (
  .A1({ S3660 }),
  .A2({ S3482 }),
  .A3({ S3663 }),
  .ZN({ S3664 })
);
AOI21_X1 #() 
AOI21_X1_3023_ (
  .A({ S3481 }),
  .B1({ S3486 }),
  .B2({ S3487 }),
  .ZN({ S3665 })
);
OAI21_X1 #() 
OAI21_X1_2781_ (
  .A({ S3506 }),
  .B1({ S3527 }),
  .B2({ S3665 }),
  .ZN({ S3666 })
);
AOI21_X1 #() 
AOI21_X1_3024_ (
  .A({ S107 }),
  .B1({ S3491 }),
  .B2({ S3495 }),
  .ZN({ S3667 })
);
NAND4_X1 #() 
NAND4_X1_628_ (
  .A1({ S3509 }),
  .A2({ S107 }),
  .A3({ S3555 }),
  .A4({ S3536 }),
  .ZN({ S3668 })
);
INV_X1 #() 
INV_X1_1753_ (
  .A({ S3668 }),
  .ZN({ S3669 })
);
OAI21_X1 #() 
OAI21_X1_2782_ (
  .A({ S25957[796] }),
  .B1({ S3669 }),
  .B2({ S3667 }),
  .ZN({ S3670 })
);
OAI211_X1 #() 
OAI211_X1_1894_ (
  .A({ S3670 }),
  .B({ S25957[797] }),
  .C1({ S25957[796] }),
  .C2({ S3666 }),
  .ZN({ S3671 })
);
NAND3_X1 #() 
NAND3_X1_5803_ (
  .A1({ S3671 }),
  .A2({ S25957[798] }),
  .A3({ S3664 }),
  .ZN({ S3672 })
);
NAND3_X1 #() 
NAND3_X1_5804_ (
  .A1({ S3657 }),
  .A2({ S3672 }),
  .A3({ S3642 }),
  .ZN({ S3673 })
);
NAND3_X1 #() 
NAND3_X1_5805_ (
  .A1({ S3641 }),
  .A2({ S24211 }),
  .A3({ S3673 }),
  .ZN({ S3674 })
);
NAND2_X1 #() 
NAND2_X1_5355_ (
  .A1({ S3641 }),
  .A2({ S3673 }),
  .ZN({ S3675 })
);
NAND2_X1 #() 
NAND2_X1_5356_ (
  .A1({ S3675 }),
  .A2({ S25957[966] }),
  .ZN({ S3676 })
);
NAND2_X1 #() 
NAND2_X1_5357_ (
  .A1({ S3676 }),
  .A2({ S3674 }),
  .ZN({ S25957[710] })
);
NAND2_X1 #() 
NAND2_X1_5358_ (
  .A1({ S25957[710] }),
  .A2({ S25957[806] }),
  .ZN({ S3677 })
);
INV_X1 #() 
INV_X1_1754_ (
  .A({ S3677 }),
  .ZN({ S3678 })
);
NOR2_X1 #() 
NOR2_X1_1350_ (
  .A1({ S25957[710] }),
  .A2({ S25957[806] }),
  .ZN({ S3679 })
);
NOR2_X1 #() 
NOR2_X1_1351_ (
  .A1({ S3678 }),
  .A2({ S3679 }),
  .ZN({ S25957[678] })
);
NOR2_X1 #() 
NOR2_X1_1352_ (
  .A1({ S25957[678] }),
  .A2({ S25957[774] }),
  .ZN({ S3680 })
);
NOR3_X1 #() 
NOR3_X1_171_ (
  .A1({ S3678 }),
  .A2({ S3679 }),
  .A3({ S2900 }),
  .ZN({ S3681 })
);
NOR2_X1 #() 
NOR2_X1_1353_ (
  .A1({ S3680 }),
  .A2({ S3681 }),
  .ZN({ S25957[646] })
);
NOR2_X1 #() 
NOR2_X1_1354_ (
  .A1({ S1284 }),
  .A2({ S1281 }),
  .ZN({ S3682 })
);
INV_X1 #() 
INV_X1_1755_ (
  .A({ S3682 }),
  .ZN({ S25957[837] })
);
NAND2_X1 #() 
NAND2_X1_5359_ (
  .A1({ S24288 }),
  .A2({ S24286 }),
  .ZN({ S3683 })
);
XNOR2_X1 #() 
XNOR2_X1_207_ (
  .A({ S3683 }),
  .B({ S25957[1125] }),
  .ZN({ S25957[997] })
);
XOR2_X1 #() 
XOR2_X1_89_ (
  .A({ S1279 }),
  .B({ S25957[997] }),
  .Z({ S25957[869] })
);
NAND3_X1 #() 
NAND3_X1_5806_ (
  .A1({ S3516 }),
  .A2({ S25957[795] }),
  .A3({ S3481 }),
  .ZN({ S3684 })
);
NAND3_X1 #() 
NAND3_X1_5807_ (
  .A1({ S3552 }),
  .A2({ S107 }),
  .A3({ S3491 }),
  .ZN({ S3685 })
);
NAND3_X1 #() 
NAND3_X1_5808_ (
  .A1({ S3685 }),
  .A2({ S25957[796] }),
  .A3({ S3684 }),
  .ZN({ S3686 })
);
NAND2_X1 #() 
NAND2_X1_5360_ (
  .A1({ S3491 }),
  .A2({ S25957[794] }),
  .ZN({ S3687 })
);
NAND2_X1 #() 
NAND2_X1_5361_ (
  .A1({ S3575 }),
  .A2({ S3687 }),
  .ZN({ S3688 })
);
OAI21_X1 #() 
OAI21_X1_2783_ (
  .A({ S3504 }),
  .B1({ S3495 }),
  .B2({ S25957[795] }),
  .ZN({ S3689 })
);
AOI21_X1 #() 
AOI21_X1_3025_ (
  .A({ S3689 }),
  .B1({ S3688 }),
  .B2({ S25957[795] }),
  .ZN({ S3690 })
);
OAI211_X1 #() 
OAI211_X1_1895_ (
  .A({ S3686 }),
  .B({ S25957[797] }),
  .C1({ S3690 }),
  .C2({ S25957[796] }),
  .ZN({ S3691 })
);
NAND3_X1 #() 
NAND3_X1_5809_ (
  .A1({ S25957[793] }),
  .A2({ S25957[795] }),
  .A3({ S3481 }),
  .ZN({ S3692 })
);
AOI21_X1 #() 
AOI21_X1_3026_ (
  .A({ S3483 }),
  .B1({ S3687 }),
  .B2({ S3692 }),
  .ZN({ S3693 })
);
AOI21_X1 #() 
AOI21_X1_3027_ (
  .A({ S25957[796] }),
  .B1({ S3659 }),
  .B2({ S3585 }),
  .ZN({ S3694 })
);
OR3_X1 #() 
OR3_X1_35_ (
  .A1({ S3694 }),
  .A2({ S3693 }),
  .A3({ S25957[797] }),
  .ZN({ S3695 })
);
NAND3_X1 #() 
NAND3_X1_5810_ (
  .A1({ S3695 }),
  .A2({ S3691 }),
  .A3({ S25957[798] }),
  .ZN({ S3696 })
);
OAI211_X1 #() 
OAI211_X1_1896_ (
  .A({ S3484 }),
  .B({ S3555 }),
  .C1({ S3488 }),
  .C2({ S107 }),
  .ZN({ S3697 })
);
AOI21_X1 #() 
AOI21_X1_3028_ (
  .A({ S3483 }),
  .B1({ S3697 }),
  .B2({ S3587 }),
  .ZN({ S3698 })
);
NAND3_X1 #() 
NAND3_X1_5811_ (
  .A1({ S3516 }),
  .A2({ S107 }),
  .A3({ S3491 }),
  .ZN({ S3699 })
);
AND2_X1 #() 
AND2_X1_342_ (
  .A1({ S3528 }),
  .A2({ S3483 }),
  .ZN({ S3700 })
);
AOI211_X1 #() 
AOI211_X1_89_ (
  .A({ S3482 }),
  .B({ S3698 }),
  .C1({ S3699 }),
  .C2({ S3700 }),
  .ZN({ S3701 })
);
NAND2_X1 #() 
NAND2_X1_5362_ (
  .A1({ S3618 }),
  .A2({ S25957[795] }),
  .ZN({ S3702 })
);
NAND2_X1 #() 
NAND2_X1_5363_ (
  .A1({ S3565 }),
  .A2({ S3527 }),
  .ZN({ S3703 })
);
NAND3_X1 #() 
NAND3_X1_5812_ (
  .A1({ S3702 }),
  .A2({ S25957[796] }),
  .A3({ S3703 }),
  .ZN({ S3704 })
);
NAND2_X1 #() 
NAND2_X1_5364_ (
  .A1({ S114 }),
  .A2({ S3488 }),
  .ZN({ S3705 })
);
NAND3_X1 #() 
NAND3_X1_5813_ (
  .A1({ S3564 }),
  .A2({ S3525 }),
  .A3({ S25957[795] }),
  .ZN({ S3706 })
);
OAI211_X1 #() 
OAI211_X1_1897_ (
  .A({ S3706 }),
  .B({ S3483 }),
  .C1({ S25957[795] }),
  .C2({ S3705 }),
  .ZN({ S3707 })
);
AOI21_X1 #() 
AOI21_X1_3029_ (
  .A({ S25957[797] }),
  .B1({ S3707 }),
  .B2({ S3704 }),
  .ZN({ S3708 })
);
OAI21_X1 #() 
OAI21_X1_2784_ (
  .A({ S3523 }),
  .B1({ S3701 }),
  .B2({ S3708 }),
  .ZN({ S3709 })
);
NAND3_X1 #() 
NAND3_X1_5814_ (
  .A1({ S3709 }),
  .A2({ S3696 }),
  .A3({ S25957[799] }),
  .ZN({ S3710 })
);
NAND4_X1 #() 
NAND4_X1_629_ (
  .A1({ S3484 }),
  .A2({ S3491 }),
  .A3({ S107 }),
  .A4({ S3502 }),
  .ZN({ S3711 })
);
NAND3_X1 #() 
NAND3_X1_5815_ (
  .A1({ S3484 }),
  .A2({ S3491 }),
  .A3({ S25957[794] }),
  .ZN({ S3712 })
);
OAI21_X1 #() 
OAI21_X1_2785_ (
  .A({ S3712 }),
  .B1({ S25957[794] }),
  .B2({ S3484 }),
  .ZN({ S3713 })
);
OAI21_X1 #() 
OAI21_X1_2786_ (
  .A({ S3711 }),
  .B1({ S3713 }),
  .B2({ S107 }),
  .ZN({ S3714 })
);
NAND4_X1 #() 
NAND4_X1_630_ (
  .A1({ S3490 }),
  .A2({ S3489 }),
  .A3({ S25957[792] }),
  .A4({ S107 }),
  .ZN({ S3715 })
);
NOR2_X1 #() 
NOR2_X1_1355_ (
  .A1({ S3715 }),
  .A2({ S3488 }),
  .ZN({ S3716 })
);
OAI21_X1 #() 
OAI21_X1_2787_ (
  .A({ S3483 }),
  .B1({ S3716 }),
  .B2({ S3519 }),
  .ZN({ S3717 })
);
OAI211_X1 #() 
OAI211_X1_1898_ (
  .A({ S3482 }),
  .B({ S3717 }),
  .C1({ S3714 }),
  .C2({ S3483 }),
  .ZN({ S3718 })
);
NAND2_X1 #() 
NAND2_X1_5365_ (
  .A1({ S3488 }),
  .A2({ S107 }),
  .ZN({ S3719 })
);
AOI21_X1 #() 
AOI21_X1_3030_ (
  .A({ S25957[796] }),
  .B1({ S3719 }),
  .B2({ S3495 }),
  .ZN({ S3720 })
);
NAND2_X1 #() 
NAND2_X1_5366_ (
  .A1({ S3666 }),
  .A2({ S3720 }),
  .ZN({ S3721 })
);
NAND3_X1 #() 
NAND3_X1_5816_ (
  .A1({ S3516 }),
  .A2({ S25957[795] }),
  .A3({ S3502 }),
  .ZN({ S3722 })
);
NAND3_X1 #() 
NAND3_X1_5817_ (
  .A1({ S3615 }),
  .A2({ S25957[796] }),
  .A3({ S3722 }),
  .ZN({ S3723 })
);
NAND3_X1 #() 
NAND3_X1_5818_ (
  .A1({ S3721 }),
  .A2({ S25957[797] }),
  .A3({ S3723 }),
  .ZN({ S3724 })
);
NAND3_X1 #() 
NAND3_X1_5819_ (
  .A1({ S3718 }),
  .A2({ S3523 }),
  .A3({ S3724 }),
  .ZN({ S3725 })
);
NAND2_X1 #() 
NAND2_X1_5367_ (
  .A1({ S3509 }),
  .A2({ S3555 }),
  .ZN({ S3726 })
);
NAND2_X1 #() 
NAND2_X1_5368_ (
  .A1({ S3536 }),
  .A2({ S25957[795] }),
  .ZN({ S3727 })
);
OAI21_X1 #() 
OAI21_X1_2788_ (
  .A({ S107 }),
  .B1({ S3491 }),
  .B2({ S25957[794] }),
  .ZN({ S3728 })
);
OAI21_X1 #() 
OAI21_X1_2789_ (
  .A({ S3728 }),
  .B1({ S3726 }),
  .B2({ S3727 }),
  .ZN({ S3729 })
);
NAND2_X1 #() 
NAND2_X1_5369_ (
  .A1({ S3729 }),
  .A2({ S3483 }),
  .ZN({ S3730 })
);
AOI21_X1 #() 
AOI21_X1_3031_ (
  .A({ S107 }),
  .B1({ S3488 }),
  .B2({ S25957[792] }),
  .ZN({ S3731 })
);
NAND2_X1 #() 
NAND2_X1_5370_ (
  .A1({ S3567 }),
  .A2({ S3731 }),
  .ZN({ S3732 })
);
NAND2_X1 #() 
NAND2_X1_5371_ (
  .A1({ S3732 }),
  .A2({ S3505 }),
  .ZN({ S3733 })
);
INV_X1 #() 
INV_X1_1756_ (
  .A({ S3733 }),
  .ZN({ S3734 })
);
AOI21_X1 #() 
AOI21_X1_3032_ (
  .A({ S25957[795] }),
  .B1({ S3705 }),
  .B2({ S3567 }),
  .ZN({ S3735 })
);
OAI22_X1 #() 
OAI22_X1_136_ (
  .A1({ S3734 }),
  .A2({ S3730 }),
  .B1({ S3501 }),
  .B2({ S3735 }),
  .ZN({ S3736 })
);
AOI21_X1 #() 
AOI21_X1_3033_ (
  .A({ S3619 }),
  .B1({ S3504 }),
  .B2({ S3481 }),
  .ZN({ S3737 })
);
AOI21_X1 #() 
AOI21_X1_3034_ (
  .A({ S3488 }),
  .B1({ S3511 }),
  .B2({ S115 }),
  .ZN({ S3738 })
);
NAND3_X1 #() 
NAND3_X1_5820_ (
  .A1({ S3552 }),
  .A2({ S107 }),
  .A3({ S3509 }),
  .ZN({ S3739 })
);
OAI211_X1 #() 
OAI211_X1_1899_ (
  .A({ S3739 }),
  .B({ S25957[796] }),
  .C1({ S3611 }),
  .C2({ S3738 }),
  .ZN({ S3740 })
);
OAI211_X1 #() 
OAI211_X1_1900_ (
  .A({ S3740 }),
  .B({ S25957[797] }),
  .C1({ S25957[796] }),
  .C2({ S3737 }),
  .ZN({ S3741 })
);
OAI211_X1 #() 
OAI211_X1_1901_ (
  .A({ S25957[798] }),
  .B({ S3741 }),
  .C1({ S3736 }),
  .C2({ S25957[797] }),
  .ZN({ S3742 })
);
NAND3_X1 #() 
NAND3_X1_5821_ (
  .A1({ S3742 }),
  .A2({ S3725 }),
  .A3({ S3642 }),
  .ZN({ S3743 })
);
NAND3_X1 #() 
NAND3_X1_5822_ (
  .A1({ S3710 }),
  .A2({ S3743 }),
  .A3({ S25957[869] }),
  .ZN({ S3744 })
);
INV_X1 #() 
INV_X1_1757_ (
  .A({ S25957[869] }),
  .ZN({ S3745 })
);
NAND2_X1 #() 
NAND2_X1_5372_ (
  .A1({ S3710 }),
  .A2({ S3743 }),
  .ZN({ S3746 })
);
NAND2_X1 #() 
NAND2_X1_5373_ (
  .A1({ S3746 }),
  .A2({ S3745 }),
  .ZN({ S3747 })
);
NAND2_X1 #() 
NAND2_X1_5374_ (
  .A1({ S3747 }),
  .A2({ S3744 }),
  .ZN({ S25957[741] })
);
INV_X1 #() 
INV_X1_1758_ (
  .A({ S25957[741] }),
  .ZN({ S3748 })
);
NAND2_X1 #() 
NAND2_X1_5375_ (
  .A1({ S3748 }),
  .A2({ S25957[837] }),
  .ZN({ S3749 })
);
NAND2_X1 #() 
NAND2_X1_5376_ (
  .A1({ S25957[741] }),
  .A2({ S3682 }),
  .ZN({ S3750 })
);
NAND3_X1 #() 
NAND3_X1_5823_ (
  .A1({ S3749 }),
  .A2({ S3750 }),
  .A3({ S354 }),
  .ZN({ S3751 })
);
NAND2_X1 #() 
NAND2_X1_5377_ (
  .A1({ S25957[741] }),
  .A2({ S25957[837] }),
  .ZN({ S3752 })
);
NAND2_X1 #() 
NAND2_X1_5378_ (
  .A1({ S3748 }),
  .A2({ S3682 }),
  .ZN({ S3753 })
);
NAND3_X1 #() 
NAND3_X1_5824_ (
  .A1({ S3753 }),
  .A2({ S25957[901] }),
  .A3({ S3752 }),
  .ZN({ S3754 })
);
AND2_X1 #() 
AND2_X1_343_ (
  .A1({ S3751 }),
  .A2({ S3754 }),
  .ZN({ S25957[645] })
);
NOR2_X1 #() 
NOR2_X1_1356_ (
  .A1({ S1339 }),
  .A2({ S1340 }),
  .ZN({ S25957[836] })
);
XOR2_X1 #() 
XOR2_X1_90_ (
  .A({ S25957[836] }),
  .B({ S25957[932] }),
  .Z({ S25957[804] })
);
INV_X1 #() 
INV_X1_1759_ (
  .A({ S25957[804] }),
  .ZN({ S3755 })
);
INV_X1 #() 
INV_X1_1760_ (
  .A({ S25957[836] }),
  .ZN({ S3756 })
);
NOR2_X1 #() 
NOR2_X1_1357_ (
  .A1({ S24355 }),
  .A2({ S24356 }),
  .ZN({ S25957[996] })
);
NAND2_X1 #() 
NAND2_X1_5379_ (
  .A1({ S1310 }),
  .A2({ S1337 }),
  .ZN({ S3757 })
);
XOR2_X1 #() 
XOR2_X1_91_ (
  .A({ S3757 }),
  .B({ S25957[996] }),
  .Z({ S3758 })
);
NOR2_X1 #() 
NOR2_X1_1358_ (
  .A1({ S3528 }),
  .A2({ S3665 }),
  .ZN({ S3759 })
);
NAND3_X1 #() 
NAND3_X1_5825_ (
  .A1({ S3516 }),
  .A2({ S107 }),
  .A3({ S3555 }),
  .ZN({ S3760 })
);
NAND3_X1 #() 
NAND3_X1_5826_ (
  .A1({ S3578 }),
  .A2({ S3760 }),
  .A3({ S3483 }),
  .ZN({ S3761 })
);
NAND2_X1 #() 
NAND2_X1_5380_ (
  .A1({ S3699 }),
  .A2({ S25957[796] }),
  .ZN({ S3762 })
);
OAI211_X1 #() 
OAI211_X1_1902_ (
  .A({ S3761 }),
  .B({ S3482 }),
  .C1({ S3759 }),
  .C2({ S3762 }),
  .ZN({ S3763 })
);
NAND3_X1 #() 
NAND3_X1_5827_ (
  .A1({ S3559 }),
  .A2({ S107 }),
  .A3({ S3481 }),
  .ZN({ S3764 })
);
NAND3_X1 #() 
NAND3_X1_5828_ (
  .A1({ S3573 }),
  .A2({ S3483 }),
  .A3({ S3764 }),
  .ZN({ S3765 })
);
OAI21_X1 #() 
OAI21_X1_2790_ (
  .A({ S107 }),
  .B1({ S3555 }),
  .B2({ S25957[793] }),
  .ZN({ S3766 })
);
AOI21_X1 #() 
AOI21_X1_3035_ (
  .A({ S3483 }),
  .B1({ S3488 }),
  .B2({ S3484 }),
  .ZN({ S3767 })
);
AOI21_X1 #() 
AOI21_X1_3036_ (
  .A({ S3482 }),
  .B1({ S3767 }),
  .B2({ S3766 }),
  .ZN({ S3768 })
);
NAND2_X1 #() 
NAND2_X1_5381_ (
  .A1({ S3765 }),
  .A2({ S3768 }),
  .ZN({ S3769 })
);
NAND2_X1 #() 
NAND2_X1_5382_ (
  .A1({ S3763 }),
  .A2({ S3769 }),
  .ZN({ S3770 })
);
NAND2_X1 #() 
NAND2_X1_5383_ (
  .A1({ S3770 }),
  .A2({ S25957[798] }),
  .ZN({ S3771 })
);
NAND3_X1 #() 
NAND3_X1_5829_ (
  .A1({ S25957[793] }),
  .A2({ S3481 }),
  .A3({ S25957[794] }),
  .ZN({ S3772 })
);
NAND3_X1 #() 
NAND3_X1_5830_ (
  .A1({ S3705 }),
  .A2({ S3772 }),
  .A3({ S107 }),
  .ZN({ S3773 })
);
NAND3_X1 #() 
NAND3_X1_5831_ (
  .A1({ S3687 }),
  .A2({ S25957[795] }),
  .A3({ S3559 }),
  .ZN({ S3774 })
);
NAND3_X1 #() 
NAND3_X1_5832_ (
  .A1({ S3773 }),
  .A2({ S3774 }),
  .A3({ S25957[796] }),
  .ZN({ S3775 })
);
OAI21_X1 #() 
OAI21_X1_2791_ (
  .A({ S107 }),
  .B1({ S3492 }),
  .B2({ S3645 }),
  .ZN({ S3776 })
);
AOI21_X1 #() 
AOI21_X1_3037_ (
  .A({ S25957[796] }),
  .B1({ S3560 }),
  .B2({ S3527 }),
  .ZN({ S3777 })
);
NAND2_X1 #() 
NAND2_X1_5384_ (
  .A1({ S3776 }),
  .A2({ S3777 }),
  .ZN({ S3778 })
);
AOI21_X1 #() 
AOI21_X1_3038_ (
  .A({ S25957[797] }),
  .B1({ S3778 }),
  .B2({ S3775 }),
  .ZN({ S3779 })
);
OAI21_X1 #() 
OAI21_X1_2792_ (
  .A({ S107 }),
  .B1({ S3534 }),
  .B2({ S3726 }),
  .ZN({ S3780 })
);
AND3_X1 #() 
AND3_X1_232_ (
  .A1({ S3500 }),
  .A2({ S3483 }),
  .A3({ S3692 }),
  .ZN({ S3781 })
);
OAI211_X1 #() 
OAI211_X1_1903_ (
  .A({ S3527 }),
  .B({ S25957[792] }),
  .C1({ S25957[794] }),
  .C2({ S25957[795] }),
  .ZN({ S3782 })
);
NAND2_X1 #() 
NAND2_X1_5385_ (
  .A1({ S3782 }),
  .A2({ S3610 }),
  .ZN({ S3783 })
);
AOI22_X1 #() 
AOI22_X1_607_ (
  .A1({ S3780 }),
  .A2({ S3781 }),
  .B1({ S25957[796] }),
  .B2({ S3783 }),
  .ZN({ S3784 })
);
OAI21_X1 #() 
OAI21_X1_2793_ (
  .A({ S3523 }),
  .B1({ S3784 }),
  .B2({ S3482 }),
  .ZN({ S3785 })
);
OAI211_X1 #() 
OAI211_X1_1904_ (
  .A({ S3771 }),
  .B({ S25957[799] }),
  .C1({ S3785 }),
  .C2({ S3779 }),
  .ZN({ S3786 })
);
AOI22_X1 #() 
AOI22_X1_608_ (
  .A1({ S3518 }),
  .A2({ S107 }),
  .B1({ S115 }),
  .B2({ S3560 }),
  .ZN({ S3787 })
);
NAND4_X1 #() 
NAND4_X1_631_ (
  .A1({ S3559 }),
  .A2({ S3495 }),
  .A3({ S25957[795] }),
  .A4({ S3502 }),
  .ZN({ S3788 })
);
NAND3_X1 #() 
NAND3_X1_5833_ (
  .A1({ S3788 }),
  .A2({ S25957[796] }),
  .A3({ S3699 }),
  .ZN({ S3789 })
);
OAI211_X1 #() 
OAI211_X1_1905_ (
  .A({ S3482 }),
  .B({ S3789 }),
  .C1({ S3787 }),
  .C2({ S25957[796] }),
  .ZN({ S3790 })
);
AOI22_X1 #() 
AOI22_X1_609_ (
  .A1({ S3618 }),
  .A2({ S25957[795] }),
  .B1({ S25957[792] }),
  .B2({ S3614 }),
  .ZN({ S3791 })
);
NAND2_X1 #() 
NAND2_X1_5386_ (
  .A1({ S3509 }),
  .A2({ S3495 }),
  .ZN({ S3792 })
);
NAND2_X1 #() 
NAND2_X1_5387_ (
  .A1({ S3792 }),
  .A2({ S107 }),
  .ZN({ S3793 })
);
NAND3_X1 #() 
NAND3_X1_5834_ (
  .A1({ S3554 }),
  .A2({ S3793 }),
  .A3({ S25957[796] }),
  .ZN({ S3794 })
);
OAI211_X1 #() 
OAI211_X1_1906_ (
  .A({ S3794 }),
  .B({ S25957[797] }),
  .C1({ S3791 }),
  .C2({ S25957[796] }),
  .ZN({ S3795 })
);
NAND3_X1 #() 
NAND3_X1_5835_ (
  .A1({ S3790 }),
  .A2({ S3795 }),
  .A3({ S3523 }),
  .ZN({ S3796 })
);
OAI21_X1 #() 
OAI21_X1_2794_ (
  .A({ S25957[795] }),
  .B1({ S3505 }),
  .B2({ S3527 }),
  .ZN({ S3797 })
);
NAND3_X1 #() 
NAND3_X1_5836_ (
  .A1({ S3517 }),
  .A2({ S107 }),
  .A3({ S3495 }),
  .ZN({ S3798 })
);
OAI211_X1 #() 
OAI211_X1_1907_ (
  .A({ S25957[796] }),
  .B({ S3797 }),
  .C1({ S3798 }),
  .C2({ S3494 }),
  .ZN({ S3799 })
);
OAI211_X1 #() 
OAI211_X1_1908_ (
  .A({ S107 }),
  .B({ S3555 }),
  .C1({ S3511 }),
  .C2({ S25957[794] }),
  .ZN({ S3800 })
);
NOR2_X1 #() 
NOR2_X1_1359_ (
  .A1({ S25957[796] }),
  .A2({ S3586 }),
  .ZN({ S3801 })
);
AOI21_X1 #() 
AOI21_X1_3039_ (
  .A({ S25957[797] }),
  .B1({ S3801 }),
  .B2({ S3800 }),
  .ZN({ S3802 })
);
NAND2_X1 #() 
NAND2_X1_5388_ (
  .A1({ S3802 }),
  .A2({ S3799 }),
  .ZN({ S3803 })
);
INV_X1 #() 
INV_X1_1761_ (
  .A({ S3803 }),
  .ZN({ S3804 })
);
OAI21_X1 #() 
OAI21_X1_2795_ (
  .A({ S107 }),
  .B1({ S3491 }),
  .B2({ S3488 }),
  .ZN({ S3805 })
);
NOR2_X1 #() 
NOR2_X1_1360_ (
  .A1({ S3534 }),
  .A2({ S3805 }),
  .ZN({ S3806 })
);
INV_X1 #() 
INV_X1_1762_ (
  .A({ S3806 }),
  .ZN({ S3807 })
);
AOI21_X1 #() 
AOI21_X1_3040_ (
  .A({ S25957[796] }),
  .B1({ S3567 }),
  .B2({ S3731 }),
  .ZN({ S3808 })
);
AND2_X1 #() 
AND2_X1_344_ (
  .A1({ S3488 }),
  .A2({ S134 }),
  .ZN({ S3809 })
);
OAI21_X1 #() 
OAI21_X1_2796_ (
  .A({ S25957[797] }),
  .B1({ S3809 }),
  .B2({ S3483 }),
  .ZN({ S3810 })
);
AOI21_X1 #() 
AOI21_X1_3041_ (
  .A({ S3810 }),
  .B1({ S3807 }),
  .B2({ S3808 }),
  .ZN({ S3811 })
);
OAI21_X1 #() 
OAI21_X1_2797_ (
  .A({ S25957[798] }),
  .B1({ S3811 }),
  .B2({ S3804 }),
  .ZN({ S3812 })
);
NAND3_X1 #() 
NAND3_X1_5837_ (
  .A1({ S3812 }),
  .A2({ S3796 }),
  .A3({ S3642 }),
  .ZN({ S3813 })
);
NAND3_X1 #() 
NAND3_X1_5838_ (
  .A1({ S3786 }),
  .A2({ S3813 }),
  .A3({ S3758 }),
  .ZN({ S3814 })
);
INV_X1 #() 
INV_X1_1763_ (
  .A({ S3758 }),
  .ZN({ S25957[868] })
);
AOI21_X1 #() 
AOI21_X1_3042_ (
  .A({ S3523 }),
  .B1({ S3763 }),
  .B2({ S3769 }),
  .ZN({ S3815 })
);
NAND2_X1 #() 
NAND2_X1_5389_ (
  .A1({ S3780 }),
  .A2({ S3781 }),
  .ZN({ S3816 })
);
AOI21_X1 #() 
AOI21_X1_3043_ (
  .A({ S3482 }),
  .B1({ S3783 }),
  .B2({ S25957[796] }),
  .ZN({ S3817 })
);
NAND2_X1 #() 
NAND2_X1_5390_ (
  .A1({ S3816 }),
  .A2({ S3817 }),
  .ZN({ S3818 })
);
NAND3_X1 #() 
NAND3_X1_5839_ (
  .A1({ S3778 }),
  .A2({ S3775 }),
  .A3({ S3482 }),
  .ZN({ S3819 })
);
AOI21_X1 #() 
AOI21_X1_3044_ (
  .A({ S25957[798] }),
  .B1({ S3819 }),
  .B2({ S3818 }),
  .ZN({ S3820 })
);
OAI21_X1 #() 
OAI21_X1_2798_ (
  .A({ S25957[799] }),
  .B1({ S3820 }),
  .B2({ S3815 }),
  .ZN({ S3821 })
);
NAND3_X1 #() 
NAND3_X1_5840_ (
  .A1({ S115 }),
  .A2({ S3495 }),
  .A3({ S25957[795] }),
  .ZN({ S3822 })
);
NAND2_X1 #() 
NAND2_X1_5391_ (
  .A1({ S115 }),
  .A2({ S3488 }),
  .ZN({ S3823 })
);
NAND3_X1 #() 
NAND3_X1_5841_ (
  .A1({ S3653 }),
  .A2({ S3823 }),
  .A3({ S107 }),
  .ZN({ S3824 })
);
AOI21_X1 #() 
AOI21_X1_3045_ (
  .A({ S25957[796] }),
  .B1({ S3824 }),
  .B2({ S3822 }),
  .ZN({ S3825 })
);
INV_X1 #() 
INV_X1_1764_ (
  .A({ S3789 }),
  .ZN({ S3826 })
);
OAI21_X1 #() 
OAI21_X1_2799_ (
  .A({ S3482 }),
  .B1({ S3825 }),
  .B2({ S3826 }),
  .ZN({ S3827 })
);
AOI22_X1 #() 
AOI22_X1_610_ (
  .A1({ S3552 }),
  .A2({ S3553 }),
  .B1({ S3792 }),
  .B2({ S107 }),
  .ZN({ S3828 })
);
AND2_X1 #() 
AND2_X1_345_ (
  .A1({ S3715 }),
  .A2({ S3483 }),
  .ZN({ S3829 })
);
AOI21_X1 #() 
AOI21_X1_3046_ (
  .A({ S3482 }),
  .B1({ S3702 }),
  .B2({ S3829 }),
  .ZN({ S3830 })
);
OAI21_X1 #() 
OAI21_X1_2800_ (
  .A({ S3830 }),
  .B1({ S3483 }),
  .B2({ S3828 }),
  .ZN({ S3831 })
);
AOI21_X1 #() 
AOI21_X1_3047_ (
  .A({ S25957[798] }),
  .B1({ S3831 }),
  .B2({ S3827 }),
  .ZN({ S3832 })
);
OAI21_X1 #() 
OAI21_X1_2801_ (
  .A({ S3483 }),
  .B1({ S3726 }),
  .B2({ S3727 }),
  .ZN({ S3833 })
);
OAI221_X1 #() 
OAI221_X1_163_ (
  .A({ S25957[797] }),
  .B1({ S3483 }),
  .B2({ S3809 }),
  .C1({ S3806 }),
  .C2({ S3833 }),
  .ZN({ S3834 })
);
AOI21_X1 #() 
AOI21_X1_3048_ (
  .A({ S3523 }),
  .B1({ S3834 }),
  .B2({ S3803 }),
  .ZN({ S3835 })
);
OAI21_X1 #() 
OAI21_X1_2802_ (
  .A({ S3642 }),
  .B1({ S3832 }),
  .B2({ S3835 }),
  .ZN({ S3836 })
);
NAND3_X1 #() 
NAND3_X1_5842_ (
  .A1({ S3836 }),
  .A2({ S25957[868] }),
  .A3({ S3821 }),
  .ZN({ S3837 })
);
NAND3_X1 #() 
NAND3_X1_5843_ (
  .A1({ S3837 }),
  .A2({ S3756 }),
  .A3({ S3814 }),
  .ZN({ S3838 })
);
NAND3_X1 #() 
NAND3_X1_5844_ (
  .A1({ S3786 }),
  .A2({ S3813 }),
  .A3({ S25957[868] }),
  .ZN({ S3839 })
);
NAND3_X1 #() 
NAND3_X1_5845_ (
  .A1({ S3836 }),
  .A2({ S3758 }),
  .A3({ S3821 }),
  .ZN({ S3840 })
);
NAND3_X1 #() 
NAND3_X1_5846_ (
  .A1({ S3840 }),
  .A2({ S25957[836] }),
  .A3({ S3839 }),
  .ZN({ S3841 })
);
NAND3_X1 #() 
NAND3_X1_5847_ (
  .A1({ S3838 }),
  .A2({ S3841 }),
  .A3({ S3755 }),
  .ZN({ S3842 })
);
NAND3_X1 #() 
NAND3_X1_5848_ (
  .A1({ S3837 }),
  .A2({ S25957[836] }),
  .A3({ S3814 }),
  .ZN({ S3843 })
);
NAND3_X1 #() 
NAND3_X1_5849_ (
  .A1({ S3840 }),
  .A2({ S3756 }),
  .A3({ S3839 }),
  .ZN({ S3844 })
);
NAND3_X1 #() 
NAND3_X1_5850_ (
  .A1({ S3843 }),
  .A2({ S3844 }),
  .A3({ S25957[804] }),
  .ZN({ S3845 })
);
NAND3_X1 #() 
NAND3_X1_5851_ (
  .A1({ S3842 }),
  .A2({ S3845 }),
  .A3({ S25957[772] }),
  .ZN({ S3846 })
);
NAND3_X1 #() 
NAND3_X1_5852_ (
  .A1({ S3843 }),
  .A2({ S3844 }),
  .A3({ S3755 }),
  .ZN({ S3847 })
);
NAND3_X1 #() 
NAND3_X1_5853_ (
  .A1({ S3838 }),
  .A2({ S3841 }),
  .A3({ S25957[804] }),
  .ZN({ S3848 })
);
NAND3_X1 #() 
NAND3_X1_5854_ (
  .A1({ S3847 }),
  .A2({ S3848 }),
  .A3({ S2901 }),
  .ZN({ S3849 })
);
AND2_X1 #() 
AND2_X1_346_ (
  .A1({ S3849 }),
  .A2({ S3846 }),
  .ZN({ S25957[644] })
);
NAND2_X1 #() 
NAND2_X1_5392_ (
  .A1({ S24440 }),
  .A2({ S24443 }),
  .ZN({ S25957[931] })
);
NOR2_X1 #() 
NOR2_X1_1361_ (
  .A1({ S1417 }),
  .A2({ S1395 }),
  .ZN({ S25957[835] })
);
XOR2_X1 #() 
XOR2_X1_92_ (
  .A({ S25957[835] }),
  .B({ S25957[931] }),
  .Z({ S25957[803] })
);
NOR2_X1 #() 
NOR2_X1_1362_ (
  .A1({ S24450 }),
  .A2({ S24451 }),
  .ZN({ S25957[963] })
);
INV_X1 #() 
INV_X1_1765_ (
  .A({ S25957[963] }),
  .ZN({ S3850 })
);
NAND2_X1 #() 
NAND2_X1_5393_ (
  .A1({ S3537 }),
  .A2({ S3504 }),
  .ZN({ S3851 })
);
AOI21_X1 #() 
AOI21_X1_3049_ (
  .A({ S107 }),
  .B1({ S3502 }),
  .B2({ S25957[793] }),
  .ZN({ S3852 })
);
AOI21_X1 #() 
AOI21_X1_3050_ (
  .A({ S3852 }),
  .B1({ S3851 }),
  .B2({ S3712 }),
  .ZN({ S3853 })
);
NAND2_X1 #() 
NAND2_X1_5394_ (
  .A1({ S3801 }),
  .A2({ S3496 }),
  .ZN({ S3854 })
);
OAI211_X1 #() 
OAI211_X1_1909_ (
  .A({ S3482 }),
  .B({ S3854 }),
  .C1({ S3853 }),
  .C2({ S3483 }),
  .ZN({ S3855 })
);
OAI211_X1 #() 
OAI211_X1_1910_ (
  .A({ S25957[796] }),
  .B({ S3822 }),
  .C1({ S3805 }),
  .C2({ S3485 }),
  .ZN({ S3856 })
);
AOI22_X1 #() 
AOI22_X1_611_ (
  .A1({ S3667 }),
  .A2({ S3517 }),
  .B1({ S3543 }),
  .B2({ S3607 }),
  .ZN({ S3857 })
);
OAI211_X1 #() 
OAI211_X1_1911_ (
  .A({ S25957[797] }),
  .B({ S3856 }),
  .C1({ S3857 }),
  .C2({ S25957[796] }),
  .ZN({ S3858 })
);
NAND3_X1 #() 
NAND3_X1_5855_ (
  .A1({ S3858 }),
  .A2({ S3855 }),
  .A3({ S25957[798] }),
  .ZN({ S3859 })
);
NAND2_X1 #() 
NAND2_X1_5395_ (
  .A1({ S3658 }),
  .A2({ S107 }),
  .ZN({ S3860 })
);
NAND3_X1 #() 
NAND3_X1_5856_ (
  .A1({ S3539 }),
  .A2({ S3653 }),
  .A3({ S25957[795] }),
  .ZN({ S3861 })
);
NAND3_X1 #() 
NAND3_X1_5857_ (
  .A1({ S3861 }),
  .A2({ S3860 }),
  .A3({ S25957[796] }),
  .ZN({ S3862 })
);
NAND3_X1 #() 
NAND3_X1_5858_ (
  .A1({ S3564 }),
  .A2({ S107 }),
  .A3({ S3516 }),
  .ZN({ S3863 })
);
AOI21_X1 #() 
AOI21_X1_3051_ (
  .A({ S107 }),
  .B1({ S25957[794] }),
  .B2({ S3481 }),
  .ZN({ S3864 })
);
NOR2_X1 #() 
NOR2_X1_1363_ (
  .A1({ S3665 }),
  .A2({ S3527 }),
  .ZN({ S3865 })
);
AOI21_X1 #() 
AOI21_X1_3052_ (
  .A({ S25957[796] }),
  .B1({ S3865 }),
  .B2({ S3864 }),
  .ZN({ S3866 })
);
NAND2_X1 #() 
NAND2_X1_5396_ (
  .A1({ S3866 }),
  .A2({ S3863 }),
  .ZN({ S3867 })
);
AOI21_X1 #() 
AOI21_X1_3053_ (
  .A({ S3482 }),
  .B1({ S3862 }),
  .B2({ S3867 }),
  .ZN({ S3868 })
);
NAND2_X1 #() 
NAND2_X1_5397_ (
  .A1({ S3559 }),
  .A2({ S25957[795] }),
  .ZN({ S3869 })
);
NAND3_X1 #() 
NAND3_X1_5859_ (
  .A1({ S115 }),
  .A2({ S3536 }),
  .A3({ S107 }),
  .ZN({ S3870 })
);
OAI211_X1 #() 
OAI211_X1_1912_ (
  .A({ S3483 }),
  .B({ S3870 }),
  .C1({ S3533 }),
  .C2({ S3869 }),
  .ZN({ S3871 })
);
NAND4_X1 #() 
NAND4_X1_632_ (
  .A1({ S3484 }),
  .A2({ S3491 }),
  .A3({ S25957[795] }),
  .A4({ S3488 }),
  .ZN({ S3872 })
);
OAI21_X1 #() 
OAI21_X1_2803_ (
  .A({ S107 }),
  .B1({ S3494 }),
  .B2({ S3542 }),
  .ZN({ S3873 })
);
NAND3_X1 #() 
NAND3_X1_5860_ (
  .A1({ S3873 }),
  .A2({ S25957[796] }),
  .A3({ S3872 }),
  .ZN({ S3874 })
);
AND3_X1 #() 
AND3_X1_233_ (
  .A1({ S3871 }),
  .A2({ S3874 }),
  .A3({ S3482 }),
  .ZN({ S3875 })
);
OAI21_X1 #() 
OAI21_X1_2804_ (
  .A({ S3523 }),
  .B1({ S3868 }),
  .B2({ S3875 }),
  .ZN({ S3876 })
);
NAND3_X1 #() 
NAND3_X1_5861_ (
  .A1({ S3876 }),
  .A2({ S25957[799] }),
  .A3({ S3859 }),
  .ZN({ S3877 })
);
OAI211_X1 #() 
OAI211_X1_1913_ (
  .A({ S3659 }),
  .B({ S25957[796] }),
  .C1({ S3583 }),
  .C2({ S3582 }),
  .ZN({ S3878 })
);
NAND3_X1 #() 
NAND3_X1_5862_ (
  .A1({ S3511 }),
  .A2({ S3495 }),
  .A3({ S107 }),
  .ZN({ S3879 })
);
NOR2_X1 #() 
NOR2_X1_1364_ (
  .A1({ S3879 }),
  .A2({ S3483 }),
  .ZN({ S3880 })
);
INV_X1 #() 
INV_X1_1766_ (
  .A({ S3880 }),
  .ZN({ S3881 })
);
NAND3_X1 #() 
NAND3_X1_5863_ (
  .A1({ S3559 }),
  .A2({ S3502 }),
  .A3({ S3495 }),
  .ZN({ S3882 })
);
NAND2_X1 #() 
NAND2_X1_5398_ (
  .A1({ S3719 }),
  .A2({ S3715 }),
  .ZN({ S3883 })
);
AOI22_X1 #() 
AOI22_X1_612_ (
  .A1({ S3883 }),
  .A2({ S3552 }),
  .B1({ S3882 }),
  .B2({ S25957[795] }),
  .ZN({ S3884 })
);
OAI21_X1 #() 
OAI21_X1_2805_ (
  .A({ S3881 }),
  .B1({ S3884 }),
  .B2({ S25957[796] }),
  .ZN({ S3885 })
);
NAND3_X1 #() 
NAND3_X1_5864_ (
  .A1({ S3559 }),
  .A2({ S107 }),
  .A3({ S3484 }),
  .ZN({ S3886 })
);
NAND2_X1 #() 
NAND2_X1_5399_ (
  .A1({ S115 }),
  .A2({ S3502 }),
  .ZN({ S3887 })
);
AOI21_X1 #() 
AOI21_X1_3054_ (
  .A({ S25957[796] }),
  .B1({ S3887 }),
  .B2({ S25957[795] }),
  .ZN({ S3888 })
);
AOI21_X1 #() 
AOI21_X1_3055_ (
  .A({ S3482 }),
  .B1({ S3888 }),
  .B2({ S3886 }),
  .ZN({ S3889 })
);
AOI22_X1 #() 
AOI22_X1_613_ (
  .A1({ S3885 }),
  .A2({ S3482 }),
  .B1({ S3889 }),
  .B2({ S3878 }),
  .ZN({ S3890 })
);
AOI21_X1 #() 
AOI21_X1_3056_ (
  .A({ S3524 }),
  .B1({ S114 }),
  .B2({ S3488 }),
  .ZN({ S3891 })
);
OAI211_X1 #() 
OAI211_X1_1914_ (
  .A({ S25957[796] }),
  .B({ S3651 }),
  .C1({ S3891 }),
  .C2({ S107 }),
  .ZN({ S3892 })
);
NAND2_X1 #() 
NAND2_X1_5400_ (
  .A1({ S3575 }),
  .A2({ S3495 }),
  .ZN({ S3893 })
);
AOI22_X1 #() 
AOI22_X1_614_ (
  .A1({ S3893 }),
  .A2({ S25957[795] }),
  .B1({ S3564 }),
  .B2({ S3565 }),
  .ZN({ S3894 })
);
OAI211_X1 #() 
OAI211_X1_1915_ (
  .A({ S3892 }),
  .B({ S3482 }),
  .C1({ S3894 }),
  .C2({ S25957[796] }),
  .ZN({ S3895 })
);
NAND3_X1 #() 
NAND3_X1_5865_ (
  .A1({ S3524 }),
  .A2({ S25957[795] }),
  .A3({ S25957[794] }),
  .ZN({ S3896 })
);
NAND3_X1 #() 
NAND3_X1_5866_ (
  .A1({ S3585 }),
  .A2({ S3896 }),
  .A3({ S25957[796] }),
  .ZN({ S3897 })
);
NAND2_X1 #() 
NAND2_X1_5401_ (
  .A1({ S3559 }),
  .A2({ S25957[792] }),
  .ZN({ S3898 })
);
OAI21_X1 #() 
OAI21_X1_2806_ (
  .A({ S3483 }),
  .B1({ S3553 }),
  .B2({ S3898 }),
  .ZN({ S3899 })
);
NAND3_X1 #() 
NAND3_X1_5867_ (
  .A1({ S3899 }),
  .A2({ S3897 }),
  .A3({ S25957[797] }),
  .ZN({ S3900 })
);
NAND3_X1 #() 
NAND3_X1_5868_ (
  .A1({ S3895 }),
  .A2({ S3523 }),
  .A3({ S3900 }),
  .ZN({ S3901 })
);
OAI211_X1 #() 
OAI211_X1_1916_ (
  .A({ S3642 }),
  .B({ S3901 }),
  .C1({ S3890 }),
  .C2({ S3523 }),
  .ZN({ S3902 })
);
NAND3_X1 #() 
NAND3_X1_5869_ (
  .A1({ S3902 }),
  .A2({ S3877 }),
  .A3({ S3850 }),
  .ZN({ S3903 })
);
NAND2_X1 #() 
NAND2_X1_5402_ (
  .A1({ S3876 }),
  .A2({ S3859 }),
  .ZN({ S3904 })
);
NAND2_X1 #() 
NAND2_X1_5403_ (
  .A1({ S3904 }),
  .A2({ S25957[799] }),
  .ZN({ S3905 })
);
NAND2_X1 #() 
NAND2_X1_5404_ (
  .A1({ S3878 }),
  .A2({ S3889 }),
  .ZN({ S3906 })
);
NAND2_X1 #() 
NAND2_X1_5405_ (
  .A1({ S3882 }),
  .A2({ S25957[795] }),
  .ZN({ S3907 })
);
NAND2_X1 #() 
NAND2_X1_5406_ (
  .A1({ S3883 }),
  .A2({ S3552 }),
  .ZN({ S3908 })
);
AOI21_X1 #() 
AOI21_X1_3057_ (
  .A({ S25957[796] }),
  .B1({ S3908 }),
  .B2({ S3907 }),
  .ZN({ S3909 })
);
OAI21_X1 #() 
OAI21_X1_2807_ (
  .A({ S3482 }),
  .B1({ S3909 }),
  .B2({ S3880 }),
  .ZN({ S3910 })
);
AOI21_X1 #() 
AOI21_X1_3058_ (
  .A({ S3523 }),
  .B1({ S3910 }),
  .B2({ S3906 }),
  .ZN({ S3911 })
);
OAI211_X1 #() 
OAI211_X1_1917_ (
  .A({ S25957[795] }),
  .B({ S115 }),
  .C1({ S3511 }),
  .C2({ S25957[794] }),
  .ZN({ S3912 })
);
AOI21_X1 #() 
AOI21_X1_3059_ (
  .A({ S3483 }),
  .B1({ S3739 }),
  .B2({ S3912 }),
  .ZN({ S3913 })
);
NAND3_X1 #() 
NAND3_X1_5870_ (
  .A1({ S3705 }),
  .A2({ S25957[795] }),
  .A3({ S3555 }),
  .ZN({ S3914 })
);
AOI21_X1 #() 
AOI21_X1_3060_ (
  .A({ S25957[796] }),
  .B1({ S3914 }),
  .B2({ S3566 }),
  .ZN({ S3915 })
);
NOR3_X1 #() 
NOR3_X1_172_ (
  .A1({ S3915 }),
  .A2({ S3913 }),
  .A3({ S25957[797] }),
  .ZN({ S3916 })
);
NAND2_X1 #() 
NAND2_X1_5407_ (
  .A1({ S3900 }),
  .A2({ S3523 }),
  .ZN({ S3917 })
);
NOR2_X1 #() 
NOR2_X1_1365_ (
  .A1({ S3916 }),
  .A2({ S3917 }),
  .ZN({ S3918 })
);
OAI21_X1 #() 
OAI21_X1_2808_ (
  .A({ S3642 }),
  .B1({ S3911 }),
  .B2({ S3918 }),
  .ZN({ S3919 })
);
NAND3_X1 #() 
NAND3_X1_5871_ (
  .A1({ S3905 }),
  .A2({ S3919 }),
  .A3({ S25957[963] }),
  .ZN({ S3920 })
);
AOI21_X1 #() 
AOI21_X1_3061_ (
  .A({ S25957[803] }),
  .B1({ S3920 }),
  .B2({ S3903 }),
  .ZN({ S3921 })
);
INV_X1 #() 
INV_X1_1767_ (
  .A({ S25957[803] }),
  .ZN({ S3922 })
);
AND3_X1 #() 
AND3_X1_234_ (
  .A1({ S3902 }),
  .A2({ S3877 }),
  .A3({ S3850 }),
  .ZN({ S3923 })
);
AOI21_X1 #() 
AOI21_X1_3062_ (
  .A({ S3850 }),
  .B1({ S3902 }),
  .B2({ S3877 }),
  .ZN({ S3924 })
);
NOR3_X1 #() 
NOR3_X1_173_ (
  .A1({ S3923 }),
  .A2({ S3924 }),
  .A3({ S3922 }),
  .ZN({ S3925 })
);
OAI21_X1 #() 
OAI21_X1_2809_ (
  .A({ S104 }),
  .B1({ S3925 }),
  .B2({ S3921 }),
  .ZN({ S3926 })
);
OAI21_X1 #() 
OAI21_X1_2810_ (
  .A({ S3922 }),
  .B1({ S3923 }),
  .B2({ S3924 }),
  .ZN({ S3927 })
);
NAND3_X1 #() 
NAND3_X1_5872_ (
  .A1({ S3920 }),
  .A2({ S25957[803] }),
  .A3({ S3903 }),
  .ZN({ S3928 })
);
NAND3_X1 #() 
NAND3_X1_5873_ (
  .A1({ S3927 }),
  .A2({ S3928 }),
  .A3({ S25957[771] }),
  .ZN({ S3929 })
);
NAND2_X1 #() 
NAND2_X1_5408_ (
  .A1({ S3926 }),
  .A2({ S3929 }),
  .ZN({ S0 })
);
OAI21_X1 #() 
OAI21_X1_2811_ (
  .A({ S25957[771] }),
  .B1({ S3925 }),
  .B2({ S3921 }),
  .ZN({ S3930 })
);
NAND3_X1 #() 
NAND3_X1_5874_ (
  .A1({ S3927 }),
  .A2({ S3928 }),
  .A3({ S104 }),
  .ZN({ S3931 })
);
NAND2_X1 #() 
NAND2_X1_5409_ (
  .A1({ S3930 }),
  .A2({ S3931 }),
  .ZN({ S25957[643] })
);
NOR2_X1 #() 
NOR2_X1_1366_ (
  .A1({ S2894 }),
  .A2({ S2895 }),
  .ZN({ S25957[832] })
);
NAND2_X1 #() 
NAND2_X1_5410_ (
  .A1({ S24556 }),
  .A2({ S24555 }),
  .ZN({ S25957[992] })
);
NAND2_X1 #() 
NAND2_X1_5411_ (
  .A1({ S1439 }),
  .A2({ S1462 }),
  .ZN({ S3932 })
);
XOR2_X1 #() 
XOR2_X1_93_ (
  .A({ S3932 }),
  .B({ S25957[992] }),
  .Z({ S3933 })
);
INV_X1 #() 
INV_X1_1768_ (
  .A({ S3933 }),
  .ZN({ S25957[864] })
);
NAND3_X1 #() 
NAND3_X1_5875_ (
  .A1({ S3568 }),
  .A2({ S107 }),
  .A3({ S3509 }),
  .ZN({ S3934 })
);
NAND3_X1 #() 
NAND3_X1_5876_ (
  .A1({ S3934 }),
  .A2({ S3483 }),
  .A3({ S3788 }),
  .ZN({ S3935 })
);
NAND2_X1 #() 
NAND2_X1_5412_ (
  .A1({ S3792 }),
  .A2({ S25957[795] }),
  .ZN({ S3936 })
);
NAND3_X1 #() 
NAND3_X1_5877_ (
  .A1({ S3824 }),
  .A2({ S25957[796] }),
  .A3({ S3936 }),
  .ZN({ S3937 })
);
NAND3_X1 #() 
NAND3_X1_5878_ (
  .A1({ S3935 }),
  .A2({ S3937 }),
  .A3({ S25957[797] }),
  .ZN({ S3938 })
);
AOI21_X1 #() 
AOI21_X1_3063_ (
  .A({ S25957[796] }),
  .B1({ S3732 }),
  .B2({ S3728 }),
  .ZN({ S3939 })
);
NAND3_X1 #() 
NAND3_X1_5879_ (
  .A1({ S3517 }),
  .A2({ S115 }),
  .A3({ S3536 }),
  .ZN({ S3940 })
);
NAND2_X1 #() 
NAND2_X1_5413_ (
  .A1({ S3940 }),
  .A2({ S107 }),
  .ZN({ S3941 })
);
NAND3_X1 #() 
NAND3_X1_5880_ (
  .A1({ S3586 }),
  .A2({ S3484 }),
  .A3({ S3491 }),
  .ZN({ S3942 })
);
AOI21_X1 #() 
AOI21_X1_3064_ (
  .A({ S3483 }),
  .B1({ S3941 }),
  .B2({ S3942 }),
  .ZN({ S3943 })
);
OAI21_X1 #() 
OAI21_X1_2812_ (
  .A({ S3482 }),
  .B1({ S3943 }),
  .B2({ S3939 }),
  .ZN({ S3944 })
);
NAND3_X1 #() 
NAND3_X1_5881_ (
  .A1({ S3944 }),
  .A2({ S25957[798] }),
  .A3({ S3938 }),
  .ZN({ S3945 })
);
NOR2_X1 #() 
NOR2_X1_1367_ (
  .A1({ S115 }),
  .A2({ S3488 }),
  .ZN({ S3946 })
);
OAI22_X1 #() 
OAI22_X1_137_ (
  .A1({ S3879 }),
  .A2({ S3887 }),
  .B1({ S3946 }),
  .B2({ S107 }),
  .ZN({ S3947 })
);
NAND4_X1 #() 
NAND4_X1_633_ (
  .A1({ S3766 }),
  .A2({ S3500 }),
  .A3({ S3692 }),
  .A4({ S3483 }),
  .ZN({ S3948 })
);
OAI211_X1 #() 
OAI211_X1_1918_ (
  .A({ S25957[797] }),
  .B({ S3948 }),
  .C1({ S3947 }),
  .C2({ S3483 }),
  .ZN({ S3949 })
);
NAND3_X1 #() 
NAND3_X1_5882_ (
  .A1({ S3517 }),
  .A2({ S25957[795] }),
  .A3({ S3481 }),
  .ZN({ S3950 })
);
NAND4_X1 #() 
NAND4_X1_634_ (
  .A1({ S115 }),
  .A2({ S3495 }),
  .A3({ S3502 }),
  .A4({ S107 }),
  .ZN({ S3951 })
);
NAND2_X1 #() 
NAND2_X1_5414_ (
  .A1({ S3951 }),
  .A2({ S3950 }),
  .ZN({ S3952 })
);
OAI21_X1 #() 
OAI21_X1_2813_ (
  .A({ S3613 }),
  .B1({ S3607 }),
  .B2({ S3719 }),
  .ZN({ S3953 })
);
NAND2_X1 #() 
NAND2_X1_5415_ (
  .A1({ S3953 }),
  .A2({ S25957[796] }),
  .ZN({ S3954 })
);
OAI211_X1 #() 
OAI211_X1_1919_ (
  .A({ S3954 }),
  .B({ S3482 }),
  .C1({ S25957[796] }),
  .C2({ S3952 }),
  .ZN({ S3955 })
);
NAND3_X1 #() 
NAND3_X1_5883_ (
  .A1({ S3955 }),
  .A2({ S3949 }),
  .A3({ S3523 }),
  .ZN({ S3956 })
);
NAND3_X1 #() 
NAND3_X1_5884_ (
  .A1({ S3945 }),
  .A2({ S3956 }),
  .A3({ S25957[799] }),
  .ZN({ S3957 })
);
NAND2_X1 #() 
NAND2_X1_5416_ (
  .A1({ S3494 }),
  .A2({ S107 }),
  .ZN({ S3958 })
);
OAI211_X1 #() 
OAI211_X1_1920_ (
  .A({ S3958 }),
  .B({ S3585 }),
  .C1({ S3534 }),
  .C2({ S107 }),
  .ZN({ S3959 })
);
NAND2_X1 #() 
NAND2_X1_5417_ (
  .A1({ S3959 }),
  .A2({ S25957[796] }),
  .ZN({ S3960 })
);
NOR2_X1 #() 
NOR2_X1_1368_ (
  .A1({ S3484 }),
  .A2({ S25957[794] }),
  .ZN({ S3961 })
);
NAND2_X1 #() 
NAND2_X1_5418_ (
  .A1({ S114 }),
  .A2({ S25957[794] }),
  .ZN({ S3962 })
);
NAND3_X1 #() 
NAND3_X1_5885_ (
  .A1({ S3962 }),
  .A2({ S25957[795] }),
  .A3({ S115 }),
  .ZN({ S3963 })
);
OAI211_X1 #() 
OAI211_X1_1921_ (
  .A({ S3963 }),
  .B({ S3483 }),
  .C1({ S3961 }),
  .C2({ S3766 }),
  .ZN({ S3964 })
);
NAND3_X1 #() 
NAND3_X1_5886_ (
  .A1({ S3960 }),
  .A2({ S3482 }),
  .A3({ S3964 }),
  .ZN({ S3965 })
);
NAND2_X1 #() 
NAND2_X1_5419_ (
  .A1({ S3491 }),
  .A2({ S3488 }),
  .ZN({ S3966 })
);
NAND3_X1 #() 
NAND3_X1_5887_ (
  .A1({ S3772 }),
  .A2({ S3966 }),
  .A3({ S25957[795] }),
  .ZN({ S3967 })
);
NAND2_X1 #() 
NAND2_X1_5420_ (
  .A1({ S3503 }),
  .A2({ S107 }),
  .ZN({ S3968 })
);
NAND3_X1 #() 
NAND3_X1_5888_ (
  .A1({ S3967 }),
  .A2({ S3483 }),
  .A3({ S3968 }),
  .ZN({ S3969 })
);
NAND3_X1 #() 
NAND3_X1_5889_ (
  .A1({ S3564 }),
  .A2({ S3705 }),
  .A3({ S25957[795] }),
  .ZN({ S3970 })
);
NAND3_X1 #() 
NAND3_X1_5890_ (
  .A1({ S3970 }),
  .A2({ S25957[796] }),
  .A3({ S3662 }),
  .ZN({ S3971 })
);
NAND3_X1 #() 
NAND3_X1_5891_ (
  .A1({ S3971 }),
  .A2({ S25957[797] }),
  .A3({ S3969 }),
  .ZN({ S3972 })
);
AOI21_X1 #() 
AOI21_X1_3065_ (
  .A({ S25957[792] }),
  .B1({ S3559 }),
  .B2({ S107 }),
  .ZN({ S3973 })
);
NAND2_X1 #() 
NAND2_X1_5421_ (
  .A1({ S25957[796] }),
  .A2({ S3509 }),
  .ZN({ S3974 })
);
OAI221_X1 #() 
OAI221_X1_164_ (
  .A({ S3482 }),
  .B1({ S3973 }),
  .B2({ S3974 }),
  .C1({ S3833 }),
  .C2({ S3689 }),
  .ZN({ S3975 })
);
NAND2_X1 #() 
NAND2_X1_5422_ (
  .A1({ S3972 }),
  .A2({ S3975 }),
  .ZN({ S3976 })
);
INV_X1 #() 
INV_X1_1769_ (
  .A({ S3491 }),
  .ZN({ S3977 })
);
OAI211_X1 #() 
OAI211_X1_1922_ (
  .A({ S3822 }),
  .B({ S25957[796] }),
  .C1({ S3977 }),
  .C2({ S3537 }),
  .ZN({ S3978 })
);
NAND3_X1 #() 
NAND3_X1_5892_ (
  .A1({ S3711 }),
  .A2({ S3635 }),
  .A3({ S3483 }),
  .ZN({ S3979 })
);
NAND2_X1 #() 
NAND2_X1_5423_ (
  .A1({ S3979 }),
  .A2({ S3978 }),
  .ZN({ S3980 })
);
AOI21_X1 #() 
AOI21_X1_3066_ (
  .A({ S25957[798] }),
  .B1({ S3980 }),
  .B2({ S25957[797] }),
  .ZN({ S3981 })
);
AOI22_X1 #() 
AOI22_X1_615_ (
  .A1({ S3976 }),
  .A2({ S25957[798] }),
  .B1({ S3965 }),
  .B2({ S3981 }),
  .ZN({ S3982 })
);
OAI211_X1 #() 
OAI211_X1_1923_ (
  .A({ S3957 }),
  .B({ S25957[864] }),
  .C1({ S3982 }),
  .C2({ S25957[799] }),
  .ZN({ S3983 })
);
NAND2_X1 #() 
NAND2_X1_5424_ (
  .A1({ S3665 }),
  .A2({ S107 }),
  .ZN({ S3984 })
);
NAND3_X1 #() 
NAND3_X1_5893_ (
  .A1({ S3886 }),
  .A2({ S3942 }),
  .A3({ S3984 }),
  .ZN({ S3985 })
);
NAND2_X1 #() 
NAND2_X1_5425_ (
  .A1({ S3985 }),
  .A2({ S25957[796] }),
  .ZN({ S3986 })
);
NAND3_X1 #() 
NAND3_X1_5894_ (
  .A1({ S3986 }),
  .A2({ S3730 }),
  .A3({ S3482 }),
  .ZN({ S3987 })
);
AOI21_X1 #() 
AOI21_X1_3067_ (
  .A({ S25957[796] }),
  .B1({ S3934 }),
  .B2({ S3788 }),
  .ZN({ S3988 })
);
AOI21_X1 #() 
AOI21_X1_3068_ (
  .A({ S107 }),
  .B1({ S3509 }),
  .B2({ S3495 }),
  .ZN({ S3989 })
);
AOI21_X1 #() 
AOI21_X1_3069_ (
  .A({ S3989 }),
  .B1({ S3518 }),
  .B2({ S107 }),
  .ZN({ S3990 })
);
OAI21_X1 #() 
OAI21_X1_2814_ (
  .A({ S25957[797] }),
  .B1({ S3990 }),
  .B2({ S3483 }),
  .ZN({ S3991 })
);
OAI211_X1 #() 
OAI211_X1_1924_ (
  .A({ S3987 }),
  .B({ S25957[798] }),
  .C1({ S3991 }),
  .C2({ S3988 }),
  .ZN({ S3992 })
);
NAND2_X1 #() 
NAND2_X1_5426_ (
  .A1({ S3952 }),
  .A2({ S3483 }),
  .ZN({ S3993 })
);
OAI211_X1 #() 
OAI211_X1_1925_ (
  .A({ S3993 }),
  .B({ S3482 }),
  .C1({ S3483 }),
  .C2({ S3953 }),
  .ZN({ S3994 })
);
NAND2_X1 #() 
NAND2_X1_5427_ (
  .A1({ S3947 }),
  .A2({ S25957[796] }),
  .ZN({ S3995 })
);
NAND3_X1 #() 
NAND3_X1_5895_ (
  .A1({ S3766 }),
  .A2({ S3500 }),
  .A3({ S3692 }),
  .ZN({ S3996 })
);
AOI21_X1 #() 
AOI21_X1_3070_ (
  .A({ S3482 }),
  .B1({ S3996 }),
  .B2({ S3483 }),
  .ZN({ S3997 })
);
NAND2_X1 #() 
NAND2_X1_5428_ (
  .A1({ S3997 }),
  .A2({ S3995 }),
  .ZN({ S3998 })
);
NAND3_X1 #() 
NAND3_X1_5896_ (
  .A1({ S3994 }),
  .A2({ S3998 }),
  .A3({ S3523 }),
  .ZN({ S3999 })
);
AOI21_X1 #() 
AOI21_X1_3071_ (
  .A({ S3642 }),
  .B1({ S3992 }),
  .B2({ S3999 }),
  .ZN({ S4000 })
);
AOI21_X1 #() 
AOI21_X1_3072_ (
  .A({ S107 }),
  .B1({ S3772 }),
  .B2({ S3966 }),
  .ZN({ S4001 })
);
NAND3_X1 #() 
NAND3_X1_5897_ (
  .A1({ S3491 }),
  .A2({ S3555 }),
  .A3({ S107 }),
  .ZN({ S4002 })
);
OAI211_X1 #() 
OAI211_X1_1926_ (
  .A({ S25957[796] }),
  .B({ S4002 }),
  .C1({ S3738 }),
  .C2({ S3722 }),
  .ZN({ S4003 })
);
NAND2_X1 #() 
NAND2_X1_5429_ (
  .A1({ S3550 }),
  .A2({ S3483 }),
  .ZN({ S4004 })
);
OAI211_X1 #() 
OAI211_X1_1927_ (
  .A({ S4003 }),
  .B({ S25957[797] }),
  .C1({ S4001 }),
  .C2({ S4004 }),
  .ZN({ S4005 })
);
OAI21_X1 #() 
OAI21_X1_2815_ (
  .A({ S25957[796] }),
  .B1({ S3973 }),
  .B2({ S3510 }),
  .ZN({ S4006 })
);
AOI21_X1 #() 
AOI21_X1_3073_ (
  .A({ S3689 }),
  .B1({ S3731 }),
  .B2({ S3567 }),
  .ZN({ S4007 })
);
OAI211_X1 #() 
OAI211_X1_1928_ (
  .A({ S4006 }),
  .B({ S3482 }),
  .C1({ S4007 }),
  .C2({ S25957[796] }),
  .ZN({ S4008 })
);
NAND3_X1 #() 
NAND3_X1_5898_ (
  .A1({ S4005 }),
  .A2({ S25957[798] }),
  .A3({ S4008 }),
  .ZN({ S4009 })
);
NAND2_X1 #() 
NAND2_X1_5430_ (
  .A1({ S3965 }),
  .A2({ S3981 }),
  .ZN({ S4010 })
);
AOI21_X1 #() 
AOI21_X1_3074_ (
  .A({ S25957[799] }),
  .B1({ S4010 }),
  .B2({ S4009 }),
  .ZN({ S4011 })
);
OAI21_X1 #() 
OAI21_X1_2816_ (
  .A({ S3933 }),
  .B1({ S4000 }),
  .B2({ S4011 }),
  .ZN({ S4012 })
);
NAND3_X1 #() 
NAND3_X1_5899_ (
  .A1({ S4012 }),
  .A2({ S25957[832] }),
  .A3({ S3983 }),
  .ZN({ S4013 })
);
INV_X1 #() 
INV_X1_1770_ (
  .A({ S25957[832] }),
  .ZN({ S4014 })
);
OAI211_X1 #() 
OAI211_X1_1929_ (
  .A({ S3957 }),
  .B({ S3933 }),
  .C1({ S3982 }),
  .C2({ S25957[799] }),
  .ZN({ S4015 })
);
OAI21_X1 #() 
OAI21_X1_2817_ (
  .A({ S25957[864] }),
  .B1({ S4000 }),
  .B2({ S4011 }),
  .ZN({ S4016 })
);
NAND3_X1 #() 
NAND3_X1_5900_ (
  .A1({ S4016 }),
  .A2({ S4014 }),
  .A3({ S4015 }),
  .ZN({ S4017 })
);
NAND3_X1 #() 
NAND3_X1_5901_ (
  .A1({ S4013 }),
  .A2({ S4017 }),
  .A3({ S499 }),
  .ZN({ S4018 })
);
NAND3_X1 #() 
NAND3_X1_5902_ (
  .A1({ S4012 }),
  .A2({ S4014 }),
  .A3({ S3983 }),
  .ZN({ S4019 })
);
NAND3_X1 #() 
NAND3_X1_5903_ (
  .A1({ S4016 }),
  .A2({ S25957[832] }),
  .A3({ S4015 }),
  .ZN({ S4020 })
);
NAND3_X1 #() 
NAND3_X1_5904_ (
  .A1({ S4019 }),
  .A2({ S4020 }),
  .A3({ S25957[896] }),
  .ZN({ S4021 })
);
NAND2_X1 #() 
NAND2_X1_5431_ (
  .A1({ S4018 }),
  .A2({ S4021 }),
  .ZN({ S25957[640] })
);
NOR2_X1 #() 
NOR2_X1_1369_ (
  .A1({ S3891 }),
  .A2({ S107 }),
  .ZN({ S4022 })
);
NAND4_X1 #() 
NAND4_X1_635_ (
  .A1({ S3525 }),
  .A2({ S3528 }),
  .A3({ S3495 }),
  .A4({ S3483 }),
  .ZN({ S4023 })
);
OAI21_X1 #() 
OAI21_X1_2818_ (
  .A({ S25957[796] }),
  .B1({ S3946 }),
  .B2({ S3537 }),
  .ZN({ S4024 })
);
OAI211_X1 #() 
OAI211_X1_1930_ (
  .A({ S4023 }),
  .B({ S25957[797] }),
  .C1({ S4022 }),
  .C2({ S4024 }),
  .ZN({ S4025 })
);
AOI21_X1 #() 
AOI21_X1_3075_ (
  .A({ S25957[796] }),
  .B1({ S3668 }),
  .B2({ S3942 }),
  .ZN({ S4026 })
);
OAI211_X1 #() 
OAI211_X1_1931_ (
  .A({ S3527 }),
  .B({ S3488 }),
  .C1({ S3481 }),
  .C2({ S25957[795] }),
  .ZN({ S4027 })
);
AOI21_X1 #() 
AOI21_X1_3076_ (
  .A({ S3483 }),
  .B1({ S114 }),
  .B2({ S25957[794] }),
  .ZN({ S4028 })
);
AND3_X1 #() 
AND3_X1_235_ (
  .A1({ S4028 }),
  .A2({ S4027 }),
  .A3({ S3950 }),
  .ZN({ S4029 })
);
OAI21_X1 #() 
OAI21_X1_2819_ (
  .A({ S3482 }),
  .B1({ S4029 }),
  .B2({ S4026 }),
  .ZN({ S4030 })
);
AOI21_X1 #() 
AOI21_X1_3077_ (
  .A({ S3523 }),
  .B1({ S4030 }),
  .B2({ S4025 }),
  .ZN({ S4031 })
);
NAND4_X1 #() 
NAND4_X1_636_ (
  .A1({ S3536 }),
  .A2({ S3555 }),
  .A3({ S25957[793] }),
  .A4({ S25957[795] }),
  .ZN({ S4032 })
);
AOI21_X1 #() 
AOI21_X1_3078_ (
  .A({ S3483 }),
  .B1({ S4032 }),
  .B2({ S3764 }),
  .ZN({ S4033 })
);
OAI21_X1 #() 
OAI21_X1_2820_ (
  .A({ S25957[797] }),
  .B1({ S3563 }),
  .B2({ S4033 }),
  .ZN({ S4034 })
);
AOI21_X1 #() 
AOI21_X1_3079_ (
  .A({ S25957[796] }),
  .B1({ S3494 }),
  .B2({ S25957[795] }),
  .ZN({ S4035 })
);
NAND2_X1 #() 
NAND2_X1_5432_ (
  .A1({ S3908 }),
  .A2({ S4035 }),
  .ZN({ S4036 })
);
NAND3_X1 #() 
NAND3_X1_5905_ (
  .A1({ S3797 }),
  .A2({ S3760 }),
  .A3({ S25957[796] }),
  .ZN({ S4037 })
);
NAND3_X1 #() 
NAND3_X1_5906_ (
  .A1({ S4036 }),
  .A2({ S3482 }),
  .A3({ S4037 }),
  .ZN({ S4038 })
);
AOI21_X1 #() 
AOI21_X1_3080_ (
  .A({ S25957[798] }),
  .B1({ S4034 }),
  .B2({ S4038 }),
  .ZN({ S4039 })
);
OAI21_X1 #() 
OAI21_X1_2821_ (
  .A({ S3642 }),
  .B1({ S4031 }),
  .B2({ S4039 }),
  .ZN({ S4040 })
);
OAI211_X1 #() 
OAI211_X1_1932_ (
  .A({ S3556 }),
  .B({ S25957[796] }),
  .C1({ S3532 }),
  .C2({ S3512 }),
  .ZN({ S4041 })
);
OAI211_X1 #() 
OAI211_X1_1933_ (
  .A({ S3483 }),
  .B({ S3805 }),
  .C1({ S3738 }),
  .C2({ S3722 }),
  .ZN({ S4042 })
);
NAND3_X1 #() 
NAND3_X1_5907_ (
  .A1({ S4042 }),
  .A2({ S4041 }),
  .A3({ S25957[797] }),
  .ZN({ S4043 })
);
NOR2_X1 #() 
NOR2_X1_1370_ (
  .A1({ S115 }),
  .A2({ S25957[794] }),
  .ZN({ S4044 })
);
NAND3_X1 #() 
NAND3_X1_5908_ (
  .A1({ S3511 }),
  .A2({ S3555 }),
  .A3({ S25957[795] }),
  .ZN({ S4045 })
);
OAI211_X1 #() 
OAI211_X1_1934_ (
  .A({ S3483 }),
  .B({ S4045 }),
  .C1({ S3879 }),
  .C2({ S4044 }),
  .ZN({ S4046 })
);
NAND2_X1 #() 
NAND2_X1_5433_ (
  .A1({ S3887 }),
  .A2({ S107 }),
  .ZN({ S4047 })
);
OAI211_X1 #() 
OAI211_X1_1935_ (
  .A({ S4047 }),
  .B({ S25957[796] }),
  .C1({ S3611 }),
  .C2({ S3738 }),
  .ZN({ S4048 })
);
NAND3_X1 #() 
NAND3_X1_5909_ (
  .A1({ S4048 }),
  .A2({ S3482 }),
  .A3({ S4046 }),
  .ZN({ S4049 })
);
NAND3_X1 #() 
NAND3_X1_5910_ (
  .A1({ S4049 }),
  .A2({ S4043 }),
  .A3({ S25957[798] }),
  .ZN({ S4050 })
);
OAI211_X1 #() 
OAI211_X1_1936_ (
  .A({ S3886 }),
  .B({ S3483 }),
  .C1({ S3645 }),
  .C2({ S107 }),
  .ZN({ S4051 })
);
AOI21_X1 #() 
AOI21_X1_3081_ (
  .A({ S107 }),
  .B1({ S3962 }),
  .B2({ S3621 }),
  .ZN({ S4052 })
);
OAI211_X1 #() 
OAI211_X1_1937_ (
  .A({ S4051 }),
  .B({ S25957[797] }),
  .C1({ S4052 }),
  .C2({ S3551 }),
  .ZN({ S4053 })
);
NAND3_X1 #() 
NAND3_X1_5911_ (
  .A1({ S3615 }),
  .A2({ S3509 }),
  .A3({ S3869 }),
  .ZN({ S4054 })
);
NAND2_X1 #() 
NAND2_X1_5434_ (
  .A1({ S4054 }),
  .A2({ S25957[796] }),
  .ZN({ S4055 })
);
NAND2_X1 #() 
NAND2_X1_5435_ (
  .A1({ S3776 }),
  .A2({ S3483 }),
  .ZN({ S4056 })
);
OAI211_X1 #() 
OAI211_X1_1938_ (
  .A({ S3482 }),
  .B({ S4055 }),
  .C1({ S4056 }),
  .C2({ S3569 }),
  .ZN({ S4057 })
);
NAND3_X1 #() 
NAND3_X1_5912_ (
  .A1({ S4057 }),
  .A2({ S3523 }),
  .A3({ S4053 }),
  .ZN({ S4058 })
);
NAND3_X1 #() 
NAND3_X1_5913_ (
  .A1({ S4058 }),
  .A2({ S25957[799] }),
  .A3({ S4050 }),
  .ZN({ S4059 })
);
AND3_X1 #() 
AND3_X1_236_ (
  .A1({ S4059 }),
  .A2({ S4040 }),
  .A3({ S25957[961] }),
  .ZN({ S4060 })
);
AOI21_X1 #() 
AOI21_X1_3082_ (
  .A({ S25957[961] }),
  .B1({ S4059 }),
  .B2({ S4040 }),
  .ZN({ S4061 })
);
OAI21_X1 #() 
OAI21_X1_2822_ (
  .A({ S25957[897] }),
  .B1({ S4060 }),
  .B2({ S4061 }),
  .ZN({ S4062 })
);
NAND3_X1 #() 
NAND3_X1_5914_ (
  .A1({ S4059 }),
  .A2({ S4040 }),
  .A3({ S25957[961] }),
  .ZN({ S4063 })
);
AND3_X1 #() 
AND3_X1_237_ (
  .A1({ S4034 }),
  .A2({ S4038 }),
  .A3({ S3642 }),
  .ZN({ S4064 })
);
OAI21_X1 #() 
OAI21_X1_2823_ (
  .A({ S4051 }),
  .B1({ S4052 }),
  .B2({ S3551 }),
  .ZN({ S4065 })
);
NAND2_X1 #() 
NAND2_X1_5436_ (
  .A1({ S4065 }),
  .A2({ S25957[797] }),
  .ZN({ S4066 })
);
NAND4_X1 #() 
NAND4_X1_637_ (
  .A1({ S3615 }),
  .A2({ S3869 }),
  .A3({ S3509 }),
  .A4({ S25957[796] }),
  .ZN({ S4067 })
);
AOI21_X1 #() 
AOI21_X1_3083_ (
  .A({ S25957[795] }),
  .B1({ S3772 }),
  .B2({ S3966 }),
  .ZN({ S4068 })
);
OAI21_X1 #() 
OAI21_X1_2824_ (
  .A({ S3483 }),
  .B1({ S3569 }),
  .B2({ S4068 }),
  .ZN({ S4069 })
);
NAND3_X1 #() 
NAND3_X1_5915_ (
  .A1({ S4069 }),
  .A2({ S3482 }),
  .A3({ S4067 }),
  .ZN({ S4070 })
);
AOI21_X1 #() 
AOI21_X1_3084_ (
  .A({ S3642 }),
  .B1({ S4070 }),
  .B2({ S4066 }),
  .ZN({ S4071 })
);
OAI21_X1 #() 
OAI21_X1_2825_ (
  .A({ S3523 }),
  .B1({ S4071 }),
  .B2({ S4064 }),
  .ZN({ S4072 })
);
NAND3_X1 #() 
NAND3_X1_5916_ (
  .A1({ S4049 }),
  .A2({ S4043 }),
  .A3({ S25957[799] }),
  .ZN({ S4073 })
);
NAND3_X1 #() 
NAND3_X1_5917_ (
  .A1({ S4030 }),
  .A2({ S4025 }),
  .A3({ S3642 }),
  .ZN({ S4074 })
);
NAND2_X1 #() 
NAND2_X1_5437_ (
  .A1({ S4074 }),
  .A2({ S4073 }),
  .ZN({ S4075 })
);
NAND2_X1 #() 
NAND2_X1_5438_ (
  .A1({ S4075 }),
  .A2({ S25957[798] }),
  .ZN({ S4076 })
);
NAND4_X1 #() 
NAND4_X1_638_ (
  .A1({ S4072 }),
  .A2({ S4076 }),
  .A3({ S24631 }),
  .A4({ S24634 }),
  .ZN({ S4077 })
);
NAND3_X1 #() 
NAND3_X1_5918_ (
  .A1({ S4077 }),
  .A2({ S490 }),
  .A3({ S4063 }),
  .ZN({ S4078 })
);
NAND2_X1 #() 
NAND2_X1_5439_ (
  .A1({ S4062 }),
  .A2({ S4078 }),
  .ZN({ S25957[641] })
);
NOR2_X1 #() 
NOR2_X1_1371_ (
  .A1({ S355 }),
  .A2({ S356 }),
  .ZN({ S25957[962] })
);
AOI21_X1 #() 
AOI21_X1_3085_ (
  .A({ S3482 }),
  .B1({ S3543 }),
  .B2({ S3552 }),
  .ZN({ S4079 })
);
NAND2_X1 #() 
NAND2_X1_5440_ (
  .A1({ S3535 }),
  .A2({ S4079 }),
  .ZN({ S4080 })
);
OAI21_X1 #() 
OAI21_X1_2826_ (
  .A({ S25957[795] }),
  .B1({ S3665 }),
  .B2({ S3527 }),
  .ZN({ S4081 })
);
NAND3_X1 #() 
NAND3_X1_5919_ (
  .A1({ S4081 }),
  .A2({ S3886 }),
  .A3({ S3984 }),
  .ZN({ S4082 })
);
NAND2_X1 #() 
NAND2_X1_5441_ (
  .A1({ S4082 }),
  .A2({ S3482 }),
  .ZN({ S4083 })
);
AOI21_X1 #() 
AOI21_X1_3086_ (
  .A({ S25957[796] }),
  .B1({ S4080 }),
  .B2({ S4083 }),
  .ZN({ S4084 })
);
INV_X1 #() 
INV_X1_1771_ (
  .A({ S3879 }),
  .ZN({ S4085 })
);
NAND2_X1 #() 
NAND2_X1_5442_ (
  .A1({ S3495 }),
  .A2({ S25957[795] }),
  .ZN({ S4086 })
);
NOR2_X1 #() 
NOR2_X1_1372_ (
  .A1({ S3491 }),
  .A2({ S25957[794] }),
  .ZN({ S4087 })
);
NAND3_X1 #() 
NAND3_X1_5920_ (
  .A1({ S25957[793] }),
  .A2({ S107 }),
  .A3({ S25957[794] }),
  .ZN({ S4088 })
);
OAI21_X1 #() 
OAI21_X1_2827_ (
  .A({ S4088 }),
  .B1({ S4087 }),
  .B2({ S4086 }),
  .ZN({ S4089 })
);
AOI21_X1 #() 
AOI21_X1_3087_ (
  .A({ S4085 }),
  .B1({ S4089 }),
  .B2({ S3482 }),
  .ZN({ S4090 })
);
AND4_X1 #() 
AND4_X1_13_ (
  .A1({ S25957[797] }),
  .A2({ S25957[796] }),
  .A3({ S25957[795] }),
  .A4({ S3484 }),
  .ZN({ S4091 })
);
AOI21_X1 #() 
AOI21_X1_3088_ (
  .A({ S25957[799] }),
  .B1({ S4091 }),
  .B2({ S3516 }),
  .ZN({ S4092 })
);
OAI21_X1 #() 
OAI21_X1_2828_ (
  .A({ S4092 }),
  .B1({ S4090 }),
  .B2({ S3483 }),
  .ZN({ S4093 })
);
NOR2_X1 #() 
NOR2_X1_1373_ (
  .A1({ S4084 }),
  .A2({ S4093 }),
  .ZN({ S4094 })
);
NAND2_X1 #() 
NAND2_X1_5443_ (
  .A1({ S3703 }),
  .A2({ S25957[796] }),
  .ZN({ S4095 })
);
AND3_X1 #() 
AND3_X1_238_ (
  .A1({ S3539 }),
  .A2({ S25957[795] }),
  .A3({ S3630 }),
  .ZN({ S4096 })
);
NAND3_X1 #() 
NAND3_X1_5921_ (
  .A1({ S3958 }),
  .A2({ S3578 }),
  .A3({ S3483 }),
  .ZN({ S4097 })
);
OAI21_X1 #() 
OAI21_X1_2829_ (
  .A({ S4097 }),
  .B1({ S4096 }),
  .B2({ S4095 }),
  .ZN({ S4098 })
);
NAND2_X1 #() 
NAND2_X1_5444_ (
  .A1({ S4098 }),
  .A2({ S3482 }),
  .ZN({ S4099 })
);
NOR2_X1 #() 
NOR2_X1_1374_ (
  .A1({ S3649 }),
  .A2({ S4086 }),
  .ZN({ S4100 })
);
OAI21_X1 #() 
OAI21_X1_2830_ (
  .A({ S25957[796] }),
  .B1({ S3540 }),
  .B2({ S4100 }),
  .ZN({ S4101 })
);
AOI21_X1 #() 
AOI21_X1_3089_ (
  .A({ S107 }),
  .B1({ S3491 }),
  .B2({ S25957[794] }),
  .ZN({ S4102 })
);
NAND2_X1 #() 
NAND2_X1_5445_ (
  .A1({ S4102 }),
  .A2({ S3539 }),
  .ZN({ S4103 })
);
NAND2_X1 #() 
NAND2_X1_5446_ (
  .A1({ S4103 }),
  .A2({ S3577 }),
  .ZN({ S4104 })
);
NAND2_X1 #() 
NAND2_X1_5447_ (
  .A1({ S4104 }),
  .A2({ S3483 }),
  .ZN({ S4105 })
);
NAND3_X1 #() 
NAND3_X1_5922_ (
  .A1({ S4105 }),
  .A2({ S4101 }),
  .A3({ S25957[797] }),
  .ZN({ S4106 })
);
AOI21_X1 #() 
AOI21_X1_3090_ (
  .A({ S3642 }),
  .B1({ S4106 }),
  .B2({ S4099 }),
  .ZN({ S4107 })
);
OAI21_X1 #() 
OAI21_X1_2831_ (
  .A({ S25957[798] }),
  .B1({ S4107 }),
  .B2({ S4094 }),
  .ZN({ S4108 })
);
NAND3_X1 #() 
NAND3_X1_5923_ (
  .A1({ S3516 }),
  .A2({ S25957[795] }),
  .A3({ S25957[792] }),
  .ZN({ S4109 })
);
OAI211_X1 #() 
OAI211_X1_1939_ (
  .A({ S25957[796] }),
  .B({ S4109 }),
  .C1({ S3556 }),
  .C2({ S3624 }),
  .ZN({ S4110 })
);
OAI211_X1 #() 
OAI211_X1_1940_ (
  .A({ S25957[795] }),
  .B({ S3491 }),
  .C1({ S3484 }),
  .C2({ S3488 }),
  .ZN({ S4111 })
);
NAND3_X1 #() 
NAND3_X1_5924_ (
  .A1({ S4111 }),
  .A2({ S3798 }),
  .A3({ S3483 }),
  .ZN({ S4112 })
);
NAND3_X1 #() 
NAND3_X1_5925_ (
  .A1({ S4110 }),
  .A2({ S25957[797] }),
  .A3({ S4112 }),
  .ZN({ S4113 })
);
NAND3_X1 #() 
NAND3_X1_5926_ (
  .A1({ S3615 }),
  .A2({ S3483 }),
  .A3({ S3613 }),
  .ZN({ S4114 })
);
NAND3_X1 #() 
NAND3_X1_5927_ (
  .A1({ S3536 }),
  .A2({ S25957[793] }),
  .A3({ S25957[795] }),
  .ZN({ S4115 })
);
NAND3_X1 #() 
NAND3_X1_5928_ (
  .A1({ S3609 }),
  .A2({ S4115 }),
  .A3({ S25957[796] }),
  .ZN({ S4116 })
);
NAND3_X1 #() 
NAND3_X1_5929_ (
  .A1({ S4114 }),
  .A2({ S4116 }),
  .A3({ S3482 }),
  .ZN({ S4117 })
);
AND3_X1 #() 
AND3_X1_239_ (
  .A1({ S4113 }),
  .A2({ S25957[799] }),
  .A3({ S4117 }),
  .ZN({ S4118 })
);
NAND3_X1 #() 
NAND3_X1_5930_ (
  .A1({ S3934 }),
  .A2({ S3482 }),
  .A3({ S3967 }),
  .ZN({ S4119 })
);
AOI22_X1 #() 
AOI22_X1_616_ (
  .A1({ S3628 }),
  .A2({ S3962 }),
  .B1({ S3614 }),
  .B2({ S3503 }),
  .ZN({ S4120 })
);
OAI211_X1 #() 
OAI211_X1_1941_ (
  .A({ S4119 }),
  .B({ S3483 }),
  .C1({ S3482 }),
  .C2({ S4120 }),
  .ZN({ S4121 })
);
NAND3_X1 #() 
NAND3_X1_5931_ (
  .A1({ S3525 }),
  .A2({ S25957[795] }),
  .A3({ S3495 }),
  .ZN({ S4122 })
);
NAND2_X1 #() 
NAND2_X1_5448_ (
  .A1({ S3863 }),
  .A2({ S4122 }),
  .ZN({ S4123 })
);
NAND2_X1 #() 
NAND2_X1_5449_ (
  .A1({ S4123 }),
  .A2({ S25957[797] }),
  .ZN({ S4124 })
);
OAI21_X1 #() 
OAI21_X1_2832_ (
  .A({ S4115 }),
  .B1({ S3805 }),
  .B2({ S3582 }),
  .ZN({ S4125 })
);
AOI21_X1 #() 
AOI21_X1_3091_ (
  .A({ S3483 }),
  .B1({ S4125 }),
  .B2({ S3482 }),
  .ZN({ S4126 })
);
NAND2_X1 #() 
NAND2_X1_5450_ (
  .A1({ S4124 }),
  .A2({ S4126 }),
  .ZN({ S4127 })
);
AOI21_X1 #() 
AOI21_X1_3092_ (
  .A({ S25957[799] }),
  .B1({ S4127 }),
  .B2({ S4121 }),
  .ZN({ S4128 })
);
OAI21_X1 #() 
OAI21_X1_2833_ (
  .A({ S3523 }),
  .B1({ S4128 }),
  .B2({ S4118 }),
  .ZN({ S4129 })
);
AOI21_X1 #() 
AOI21_X1_3093_ (
  .A({ S25957[962] }),
  .B1({ S4108 }),
  .B2({ S4129 }),
  .ZN({ S4130 })
);
INV_X1 #() 
INV_X1_1772_ (
  .A({ S25957[962] }),
  .ZN({ S4131 })
);
AOI21_X1 #() 
AOI21_X1_3094_ (
  .A({ S3483 }),
  .B1({ S3934 }),
  .B2({ S3561 }),
  .ZN({ S4132 })
);
AOI21_X1 #() 
AOI21_X1_3095_ (
  .A({ S25957[796] }),
  .B1({ S4103 }),
  .B2({ S3577 }),
  .ZN({ S4133 })
);
OAI21_X1 #() 
OAI21_X1_2834_ (
  .A({ S25957[797] }),
  .B1({ S4132 }),
  .B2({ S4133 }),
  .ZN({ S4134 })
);
OAI211_X1 #() 
OAI211_X1_1942_ (
  .A({ S3482 }),
  .B({ S4097 }),
  .C1({ S4096 }),
  .C2({ S4095 }),
  .ZN({ S4135 })
);
AOI21_X1 #() 
AOI21_X1_3096_ (
  .A({ S3523 }),
  .B1({ S4134 }),
  .B2({ S4135 }),
  .ZN({ S4136 })
);
AOI21_X1 #() 
AOI21_X1_3097_ (
  .A({ S25957[798] }),
  .B1({ S4113 }),
  .B2({ S4117 }),
  .ZN({ S4137 })
);
OAI21_X1 #() 
OAI21_X1_2835_ (
  .A({ S25957[799] }),
  .B1({ S4136 }),
  .B2({ S4137 }),
  .ZN({ S4138 })
);
AOI21_X1 #() 
AOI21_X1_3098_ (
  .A({ S3483 }),
  .B1({ S3773 }),
  .B2({ S4115 }),
  .ZN({ S4139 })
);
NAND3_X1 #() 
NAND3_X1_5932_ (
  .A1({ S3539 }),
  .A2({ S107 }),
  .A3({ S3517 }),
  .ZN({ S4140 })
);
AOI21_X1 #() 
AOI21_X1_3099_ (
  .A({ S25957[796] }),
  .B1({ S3646 }),
  .B2({ S4140 }),
  .ZN({ S4141 })
);
OAI21_X1 #() 
OAI21_X1_2836_ (
  .A({ S3482 }),
  .B1({ S4141 }),
  .B2({ S4139 }),
  .ZN({ S4142 })
);
NAND3_X1 #() 
NAND3_X1_5933_ (
  .A1({ S3863 }),
  .A2({ S4122 }),
  .A3({ S25957[796] }),
  .ZN({ S4143 })
);
AOI21_X1 #() 
AOI21_X1_3100_ (
  .A({ S3482 }),
  .B1({ S4120 }),
  .B2({ S3483 }),
  .ZN({ S4144 })
);
AOI21_X1 #() 
AOI21_X1_3101_ (
  .A({ S25957[798] }),
  .B1({ S4144 }),
  .B2({ S4143 }),
  .ZN({ S4145 })
);
NAND2_X1 #() 
NAND2_X1_5451_ (
  .A1({ S4145 }),
  .A2({ S4142 }),
  .ZN({ S4146 })
);
OAI21_X1 #() 
OAI21_X1_2837_ (
  .A({ S25957[795] }),
  .B1({ S3542 }),
  .B2({ S25957[793] }),
  .ZN({ S4147 })
);
AOI21_X1 #() 
AOI21_X1_3102_ (
  .A({ S3483 }),
  .B1({ S4147 }),
  .B2({ S3879 }),
  .ZN({ S4148 })
);
AOI21_X1 #() 
AOI21_X1_3103_ (
  .A({ S25957[796] }),
  .B1({ S3543 }),
  .B2({ S3552 }),
  .ZN({ S4149 })
);
AOI21_X1 #() 
AOI21_X1_3104_ (
  .A({ S4148 }),
  .B1({ S3535 }),
  .B2({ S4149 }),
  .ZN({ S4150 })
);
NAND3_X1 #() 
NAND3_X1_5934_ (
  .A1({ S3941 }),
  .A2({ S3483 }),
  .A3({ S4081 }),
  .ZN({ S4151 })
);
NAND2_X1 #() 
NAND2_X1_5452_ (
  .A1({ S3560 }),
  .A2({ S3610 }),
  .ZN({ S4152 })
);
NAND3_X1 #() 
NAND3_X1_5935_ (
  .A1({ S3516 }),
  .A2({ S3517 }),
  .A3({ S25957[792] }),
  .ZN({ S4153 })
);
NAND2_X1 #() 
NAND2_X1_5453_ (
  .A1({ S4153 }),
  .A2({ S107 }),
  .ZN({ S4154 })
);
NAND3_X1 #() 
NAND3_X1_5936_ (
  .A1({ S4154 }),
  .A2({ S25957[796] }),
  .A3({ S4152 }),
  .ZN({ S4155 })
);
NAND3_X1 #() 
NAND3_X1_5937_ (
  .A1({ S4155 }),
  .A2({ S4151 }),
  .A3({ S3482 }),
  .ZN({ S4156 })
);
OAI211_X1 #() 
OAI211_X1_1943_ (
  .A({ S4156 }),
  .B({ S25957[798] }),
  .C1({ S4150 }),
  .C2({ S3482 }),
  .ZN({ S4157 })
);
NAND3_X1 #() 
NAND3_X1_5938_ (
  .A1({ S4146 }),
  .A2({ S3642 }),
  .A3({ S4157 }),
  .ZN({ S4158 })
);
AOI21_X1 #() 
AOI21_X1_3105_ (
  .A({ S4131 }),
  .B1({ S4138 }),
  .B2({ S4158 }),
  .ZN({ S4159 })
);
OAI21_X1 #() 
OAI21_X1_2838_ (
  .A({ S359 }),
  .B1({ S4130 }),
  .B2({ S4159 }),
  .ZN({ S4160 })
);
NAND3_X1 #() 
NAND3_X1_5939_ (
  .A1({ S4138 }),
  .A2({ S4131 }),
  .A3({ S4158 }),
  .ZN({ S4161 })
);
NAND3_X1 #() 
NAND3_X1_5940_ (
  .A1({ S4108 }),
  .A2({ S4129 }),
  .A3({ S25957[962] }),
  .ZN({ S4162 })
);
NAND3_X1 #() 
NAND3_X1_5941_ (
  .A1({ S4162 }),
  .A2({ S4161 }),
  .A3({ S25957[898] }),
  .ZN({ S4163 })
);
NAND2_X1 #() 
NAND2_X1_5454_ (
  .A1({ S4160 }),
  .A2({ S4163 }),
  .ZN({ S25957[642] })
);
OAI21_X1 #() 
OAI21_X1_2839_ (
  .A({ S264 }),
  .B1({ S260 }),
  .B2({ S257 }),
  .ZN({ S4164 })
);
NAND3_X1 #() 
NAND3_X1_5942_ (
  .A1({ S265 }),
  .A2({ S25957[913] }),
  .A3({ S266 }),
  .ZN({ S4165 })
);
NAND3_X1 #() 
NAND3_X1_5943_ (
  .A1({ S25957[784] }),
  .A2({ S4164 }),
  .A3({ S4165 }),
  .ZN({ S4166 })
);
INV_X1 #() 
INV_X1_1773_ (
  .A({ S4166 }),
  .ZN({ S1 })
);
NAND3_X1 #() 
NAND3_X1_5944_ (
  .A1({ S2749 }),
  .A2({ S261 }),
  .A3({ S267 }),
  .ZN({ S2 })
);
XNOR2_X1 #() 
XNOR2_X1_208_ (
  .A({ S24826 }),
  .B({ S25957[1151] }),
  .ZN({ S25957[1023] })
);
XNOR2_X1 #() 
XNOR2_X1_209_ (
  .A({ S1727 }),
  .B({ S25957[1023] }),
  .ZN({ S4167 })
);
INV_X1 #() 
INV_X1_1774_ (
  .A({ S4167 }),
  .ZN({ S25957[895] })
);
AOI21_X1 #() 
AOI21_X1_3106_ (
  .A({ S349 }),
  .B1({ S350 }),
  .B2({ S351 }),
  .ZN({ S4168 })
);
AND3_X1 #() 
AND3_X1_240_ (
  .A1({ S351 }),
  .A2({ S350 }),
  .A3({ S349 }),
  .ZN({ S4169 })
);
NOR2_X1 #() 
NOR2_X1_1375_ (
  .A1({ S4169 }),
  .A2({ S4168 }),
  .ZN({ S4170 })
);
NAND4_X1 #() 
NAND4_X1_639_ (
  .A1({ S4170 }),
  .A2({ S267 }),
  .A3({ S261 }),
  .A4({ S25957[784] }),
  .ZN({ S4171 })
);
AOI21_X1 #() 
AOI21_X1_3107_ (
  .A({ S98 }),
  .B1({ S2749 }),
  .B2({ S25957[786] }),
  .ZN({ S4172 })
);
NAND2_X1 #() 
NAND2_X1_5455_ (
  .A1({ S4172 }),
  .A2({ S4171 }),
  .ZN({ S4173 })
);
NAND4_X1 #() 
NAND4_X1_640_ (
  .A1({ S344 }),
  .A2({ S25918 }),
  .A3({ S25924 }),
  .A4({ S352 }),
  .ZN({ S4174 })
);
NAND3_X1 #() 
NAND3_X1_5945_ (
  .A1({ S25957[785] }),
  .A2({ S4174 }),
  .A3({ S98 }),
  .ZN({ S4175 })
);
AND2_X1 #() 
AND2_X1_347_ (
  .A1({ S4175 }),
  .A2({ S25957[788] }),
  .ZN({ S4176 })
);
NAND3_X1 #() 
NAND3_X1_5946_ (
  .A1({ S2749 }),
  .A2({ S4164 }),
  .A3({ S4165 }),
  .ZN({ S4177 })
);
NAND3_X1 #() 
NAND3_X1_5947_ (
  .A1({ S25957[784] }),
  .A2({ S261 }),
  .A3({ S267 }),
  .ZN({ S4178 })
);
AOI21_X1 #() 
AOI21_X1_3108_ (
  .A({ S4170 }),
  .B1({ S4177 }),
  .B2({ S4178 }),
  .ZN({ S4179 })
);
NAND4_X1 #() 
NAND4_X1_641_ (
  .A1({ S344 }),
  .A2({ S2747 }),
  .A3({ S2748 }),
  .A4({ S352 }),
  .ZN({ S4180 })
);
NOR2_X1 #() 
NOR2_X1_1376_ (
  .A1({ S25957[785] }),
  .A2({ S4180 }),
  .ZN({ S4181 })
);
OAI21_X1 #() 
OAI21_X1_2840_ (
  .A({ S25957[787] }),
  .B1({ S4179 }),
  .B2({ S4181 }),
  .ZN({ S4182 })
);
NAND3_X1 #() 
NAND3_X1_5948_ (
  .A1({ S25957[786] }),
  .A2({ S4164 }),
  .A3({ S4165 }),
  .ZN({ S4183 })
);
NAND2_X1 #() 
NAND2_X1_5456_ (
  .A1({ S4183 }),
  .A2({ S98 }),
  .ZN({ S4184 })
);
NAND2_X1 #() 
NAND2_X1_5457_ (
  .A1({ S4184 }),
  .A2({ S2524 }),
  .ZN({ S4185 })
);
OAI211_X1 #() 
OAI211_X1_1944_ (
  .A({ S25918 }),
  .B({ S25924 }),
  .C1({ S4169 }),
  .C2({ S4168 }),
  .ZN({ S4186 })
);
NAND3_X1 #() 
NAND3_X1_5949_ (
  .A1({ S2524 }),
  .A2({ S4166 }),
  .A3({ S4186 }),
  .ZN({ S4187 })
);
NAND2_X1 #() 
NAND2_X1_5458_ (
  .A1({ S4185 }),
  .A2({ S4187 }),
  .ZN({ S4188 })
);
AOI22_X1 #() 
AOI22_X1_617_ (
  .A1({ S4182 }),
  .A2({ S4188 }),
  .B1({ S4176 }),
  .B2({ S4173 }),
  .ZN({ S4189 })
);
NAND4_X1 #() 
NAND4_X1_642_ (
  .A1({ S4164 }),
  .A2({ S4165 }),
  .A3({ S344 }),
  .A4({ S352 }),
  .ZN({ S4190 })
);
NAND2_X1 #() 
NAND2_X1_5459_ (
  .A1({ S4190 }),
  .A2({ S25957[787] }),
  .ZN({ S4191 })
);
NAND4_X1 #() 
NAND4_X1_643_ (
  .A1({ S25957[786] }),
  .A2({ S2749 }),
  .A3({ S261 }),
  .A4({ S267 }),
  .ZN({ S4192 })
);
INV_X1 #() 
INV_X1_1775_ (
  .A({ S4192 }),
  .ZN({ S4193 })
);
NAND2_X1 #() 
NAND2_X1_5460_ (
  .A1({ S2 }),
  .A2({ S4170 }),
  .ZN({ S4194 })
);
NAND3_X1 #() 
NAND3_X1_5950_ (
  .A1({ S4194 }),
  .A2({ S98 }),
  .A3({ S4192 }),
  .ZN({ S4195 })
);
OAI211_X1 #() 
OAI211_X1_1945_ (
  .A({ S4195 }),
  .B({ S2524 }),
  .C1({ S4191 }),
  .C2({ S4193 }),
  .ZN({ S4196 })
);
NAND3_X1 #() 
NAND3_X1_5951_ (
  .A1({ S25957[786] }),
  .A2({ S261 }),
  .A3({ S267 }),
  .ZN({ S4197 })
);
NAND3_X1 #() 
NAND3_X1_5952_ (
  .A1({ S4197 }),
  .A2({ S4166 }),
  .A3({ S25957[787] }),
  .ZN({ S4198 })
);
NAND2_X1 #() 
NAND2_X1_5461_ (
  .A1({ S4177 }),
  .A2({ S98 }),
  .ZN({ S4199 })
);
AND2_X1 #() 
AND2_X1_348_ (
  .A1({ S4198 }),
  .A2({ S4199 }),
  .ZN({ S4200 })
);
OAI211_X1 #() 
OAI211_X1_1946_ (
  .A({ S4196 }),
  .B({ S25673 }),
  .C1({ S2524 }),
  .C2({ S4200 }),
  .ZN({ S4201 })
);
OAI211_X1 #() 
OAI211_X1_1947_ (
  .A({ S4201 }),
  .B({ S25957[790] }),
  .C1({ S4189 }),
  .C2({ S25673 }),
  .ZN({ S4202 })
);
NAND3_X1 #() 
NAND3_X1_5953_ (
  .A1({ S4166 }),
  .A2({ S2 }),
  .A3({ S25957[786] }),
  .ZN({ S4203 })
);
NAND3_X1 #() 
NAND3_X1_5954_ (
  .A1({ S4177 }),
  .A2({ S4178 }),
  .A3({ S4170 }),
  .ZN({ S4204 })
);
AOI21_X1 #() 
AOI21_X1_3109_ (
  .A({ S98 }),
  .B1({ S4203 }),
  .B2({ S4204 }),
  .ZN({ S4205 })
);
AOI22_X1 #() 
AOI22_X1_618_ (
  .A1({ S261 }),
  .A2({ S267 }),
  .B1({ S352 }),
  .B2({ S344 }),
  .ZN({ S4206 })
);
NAND2_X1 #() 
NAND2_X1_5462_ (
  .A1({ S4180 }),
  .A2({ S98 }),
  .ZN({ S4207 })
);
NOR2_X1 #() 
NOR2_X1_1377_ (
  .A1({ S4207 }),
  .A2({ S4206 }),
  .ZN({ S4208 })
);
OAI21_X1 #() 
OAI21_X1_2841_ (
  .A({ S25957[788] }),
  .B1({ S4205 }),
  .B2({ S4208 }),
  .ZN({ S4209 })
);
AOI22_X1 #() 
AOI22_X1_619_ (
  .A1({ S25957[786] }),
  .A2({ S2749 }),
  .B1({ S25833 }),
  .B2({ S25828 }),
  .ZN({ S4210 })
);
NAND2_X1 #() 
NAND2_X1_5463_ (
  .A1({ S25957[785] }),
  .A2({ S4180 }),
  .ZN({ S4211 })
);
NAND3_X1 #() 
NAND3_X1_5955_ (
  .A1({ S4171 }),
  .A2({ S4211 }),
  .A3({ S4210 }),
  .ZN({ S4212 })
);
NAND4_X1 #() 
NAND4_X1_644_ (
  .A1({ S261 }),
  .A2({ S267 }),
  .A3({ S344 }),
  .A4({ S352 }),
  .ZN({ S4213 })
);
INV_X1 #() 
INV_X1_1776_ (
  .A({ S4213 }),
  .ZN({ S4214 })
);
AOI21_X1 #() 
AOI21_X1_3110_ (
  .A({ S25957[788] }),
  .B1({ S4214 }),
  .B2({ S25957[787] }),
  .ZN({ S4215 })
);
NAND2_X1 #() 
NAND2_X1_5464_ (
  .A1({ S4215 }),
  .A2({ S4212 }),
  .ZN({ S4216 })
);
AOI21_X1 #() 
AOI21_X1_3111_ (
  .A({ S25957[789] }),
  .B1({ S4209 }),
  .B2({ S4216 }),
  .ZN({ S4217 })
);
OAI211_X1 #() 
OAI211_X1_1948_ (
  .A({ S2747 }),
  .B({ S2748 }),
  .C1({ S4169 }),
  .C2({ S4168 }),
  .ZN({ S4218 })
);
NAND2_X1 #() 
NAND2_X1_5465_ (
  .A1({ S25957[785] }),
  .A2({ S98 }),
  .ZN({ S4219 })
);
INV_X1 #() 
INV_X1_1777_ (
  .A({ S4219 }),
  .ZN({ S4220 })
);
INV_X1 #() 
INV_X1_1778_ (
  .A({ S4218 }),
  .ZN({ S4221 })
);
NAND2_X1 #() 
NAND2_X1_5466_ (
  .A1({ S4221 }),
  .A2({ S25957[787] }),
  .ZN({ S4222 })
);
NAND4_X1 #() 
NAND4_X1_645_ (
  .A1({ S261 }),
  .A2({ S267 }),
  .A3({ S25828 }),
  .A4({ S25833 }),
  .ZN({ S4223 })
);
INV_X1 #() 
INV_X1_1779_ (
  .A({ S4223 }),
  .ZN({ S4224 })
);
NOR2_X1 #() 
NOR2_X1_1378_ (
  .A1({ S4224 }),
  .A2({ S2524 }),
  .ZN({ S4225 })
);
NAND2_X1 #() 
NAND2_X1_5467_ (
  .A1({ S4225 }),
  .A2({ S4222 }),
  .ZN({ S4226 })
);
AOI21_X1 #() 
AOI21_X1_3112_ (
  .A({ S4226 }),
  .B1({ S4220 }),
  .B2({ S4218 }),
  .ZN({ S4227 })
);
NAND4_X1 #() 
NAND4_X1_646_ (
  .A1({ S4170 }),
  .A2({ S267 }),
  .A3({ S261 }),
  .A4({ S2749 }),
  .ZN({ S4228 })
);
NAND2_X1 #() 
NAND2_X1_5468_ (
  .A1({ S4228 }),
  .A2({ S98 }),
  .ZN({ S4229 })
);
AOI21_X1 #() 
AOI21_X1_3113_ (
  .A({ S25957[788] }),
  .B1({ S1 }),
  .B2({ S25957[787] }),
  .ZN({ S4230 })
);
AOI211_X1 #() 
AOI211_X1_90_ (
  .A({ S25673 }),
  .B({ S4227 }),
  .C1({ S4229 }),
  .C2({ S4230 }),
  .ZN({ S4231 })
);
OAI21_X1 #() 
OAI21_X1_2842_ (
  .A({ S25607 }),
  .B1({ S4231 }),
  .B2({ S4217 }),
  .ZN({ S4232 })
);
AOI21_X1 #() 
AOI21_X1_3114_ (
  .A({ S2361 }),
  .B1({ S4232 }),
  .B2({ S4202 }),
  .ZN({ S4233 })
);
INV_X1 #() 
INV_X1_1780_ (
  .A({ S4190 }),
  .ZN({ S4234 })
);
NAND2_X1 #() 
NAND2_X1_5469_ (
  .A1({ S25957[787] }),
  .A2({ S4218 }),
  .ZN({ S4235 })
);
NAND4_X1 #() 
NAND4_X1_647_ (
  .A1({ S4197 }),
  .A2({ S4190 }),
  .A3({ S4174 }),
  .A4({ S4186 }),
  .ZN({ S4236 })
);
AOI21_X1 #() 
AOI21_X1_3115_ (
  .A({ S25957[788] }),
  .B1({ S4236 }),
  .B2({ S98 }),
  .ZN({ S4237 })
);
OAI21_X1 #() 
OAI21_X1_2843_ (
  .A({ S4237 }),
  .B1({ S4234 }),
  .B2({ S4235 }),
  .ZN({ S4238 })
);
NAND2_X1 #() 
NAND2_X1_5470_ (
  .A1({ S4166 }),
  .A2({ S25957[786] }),
  .ZN({ S4239 })
);
AOI21_X1 #() 
AOI21_X1_3116_ (
  .A({ S98 }),
  .B1({ S4204 }),
  .B2({ S4239 }),
  .ZN({ S4240 })
);
INV_X1 #() 
INV_X1_1781_ (
  .A({ S4207 }),
  .ZN({ S4241 })
);
NAND2_X1 #() 
NAND2_X1_5471_ (
  .A1({ S4203 }),
  .A2({ S4241 }),
  .ZN({ S4242 })
);
NAND2_X1 #() 
NAND2_X1_5472_ (
  .A1({ S4242 }),
  .A2({ S25957[788] }),
  .ZN({ S4243 })
);
OAI21_X1 #() 
OAI21_X1_2844_ (
  .A({ S4238 }),
  .B1({ S4240 }),
  .B2({ S4243 }),
  .ZN({ S4244 })
);
NAND2_X1 #() 
NAND2_X1_5473_ (
  .A1({ S4244 }),
  .A2({ S25673 }),
  .ZN({ S4245 })
);
AOI21_X1 #() 
AOI21_X1_3117_ (
  .A({ S2524 }),
  .B1({ S4206 }),
  .B2({ S25957[787] }),
  .ZN({ S4246 })
);
INV_X1 #() 
INV_X1_1782_ (
  .A({ S4246 }),
  .ZN({ S4247 })
);
NAND2_X1 #() 
NAND2_X1_5474_ (
  .A1({ S4174 }),
  .A2({ S98 }),
  .ZN({ S4248 })
);
NAND2_X1 #() 
NAND2_X1_5475_ (
  .A1({ S4164 }),
  .A2({ S4165 }),
  .ZN({ S4249 })
);
NOR2_X1 #() 
NOR2_X1_1379_ (
  .A1({ S4186 }),
  .A2({ S4249 }),
  .ZN({ S4250 })
);
NOR2_X1 #() 
NOR2_X1_1380_ (
  .A1({ S4250 }),
  .A2({ S4248 }),
  .ZN({ S4251 })
);
AOI211_X1 #() 
AOI211_X1_91_ (
  .A({ S4251 }),
  .B({ S4247 }),
  .C1({ S4172 }),
  .C2({ S4166 }),
  .ZN({ S4252 })
);
NAND2_X1 #() 
NAND2_X1_5476_ (
  .A1({ S4197 }),
  .A2({ S4186 }),
  .ZN({ S4253 })
);
NAND2_X1 #() 
NAND2_X1_5477_ (
  .A1({ S4178 }),
  .A2({ S4170 }),
  .ZN({ S4254 })
);
AOI21_X1 #() 
AOI21_X1_3118_ (
  .A({ S98 }),
  .B1({ S4254 }),
  .B2({ S4197 }),
  .ZN({ S4255 })
);
AOI21_X1 #() 
AOI21_X1_3119_ (
  .A({ S4255 }),
  .B1({ S4253 }),
  .B2({ S98 }),
  .ZN({ S4256 })
);
OAI21_X1 #() 
OAI21_X1_2845_ (
  .A({ S25957[789] }),
  .B1({ S4256 }),
  .B2({ S25957[788] }),
  .ZN({ S4257 })
);
OAI211_X1 #() 
OAI211_X1_1949_ (
  .A({ S4245 }),
  .B({ S25957[790] }),
  .C1({ S4257 }),
  .C2({ S4252 }),
  .ZN({ S4258 })
);
AOI22_X1 #() 
AOI22_X1_620_ (
  .A1({ S25828 }),
  .A2({ S25833 }),
  .B1({ S25924 }),
  .B2({ S25918 }),
  .ZN({ S4259 })
);
NOR2_X1 #() 
NOR2_X1_1381_ (
  .A1({ S4214 }),
  .A2({ S4235 }),
  .ZN({ S4260 })
);
NOR3_X1 #() 
NOR3_X1_174_ (
  .A1({ S4260 }),
  .A2({ S4259 }),
  .A3({ S2524 }),
  .ZN({ S4261 })
);
NAND2_X1 #() 
NAND2_X1_5478_ (
  .A1({ S4166 }),
  .A2({ S4170 }),
  .ZN({ S4262 })
);
INV_X1 #() 
INV_X1_1783_ (
  .A({ S4262 }),
  .ZN({ S4263 })
);
NAND3_X1 #() 
NAND3_X1_5956_ (
  .A1({ S4190 }),
  .A2({ S4178 }),
  .A3({ S25957[787] }),
  .ZN({ S4264 })
);
OAI21_X1 #() 
OAI21_X1_2846_ (
  .A({ S4264 }),
  .B1({ S4263 }),
  .B2({ S4184 }),
  .ZN({ S4265 })
);
AOI21_X1 #() 
AOI21_X1_3120_ (
  .A({ S4261 }),
  .B1({ S2524 }),
  .B2({ S4265 }),
  .ZN({ S4266 })
);
OAI21_X1 #() 
OAI21_X1_2847_ (
  .A({ S98 }),
  .B1({ S4249 }),
  .B2({ S4180 }),
  .ZN({ S4267 })
);
OAI21_X1 #() 
OAI21_X1_2848_ (
  .A({ S25957[788] }),
  .B1({ S4179 }),
  .B2({ S4267 }),
  .ZN({ S4268 })
);
NOR3_X1 #() 
NOR3_X1_175_ (
  .A1({ S4268 }),
  .A2({ S4172 }),
  .A3({ S4224 }),
  .ZN({ S4269 })
);
NAND4_X1 #() 
NAND4_X1_648_ (
  .A1({ S4177 }),
  .A2({ S4178 }),
  .A3({ S98 }),
  .A4({ S25957[786] }),
  .ZN({ S4270 })
);
INV_X1 #() 
INV_X1_1784_ (
  .A({ S4270 }),
  .ZN({ S4271 })
);
AOI211_X1 #() 
AOI211_X1_92_ (
  .A({ S25957[788] }),
  .B({ S4271 }),
  .C1({ S25957[787] }),
  .C2({ S4253 }),
  .ZN({ S4272 })
);
OAI21_X1 #() 
OAI21_X1_2849_ (
  .A({ S25673 }),
  .B1({ S4272 }),
  .B2({ S4269 }),
  .ZN({ S4273 })
);
OAI21_X1 #() 
OAI21_X1_2850_ (
  .A({ S4273 }),
  .B1({ S25673 }),
  .B2({ S4266 }),
  .ZN({ S4274 })
);
NAND2_X1 #() 
NAND2_X1_5479_ (
  .A1({ S4274 }),
  .A2({ S25607 }),
  .ZN({ S4275 })
);
AOI21_X1 #() 
AOI21_X1_3121_ (
  .A({ S25957[791] }),
  .B1({ S4275 }),
  .B2({ S4258 }),
  .ZN({ S4276 })
);
OR3_X1 #() 
OR3_X1_36_ (
  .A1({ S4276 }),
  .A2({ S4233 }),
  .A3({ S25957[895] }),
  .ZN({ S4277 })
);
OAI21_X1 #() 
OAI21_X1_2851_ (
  .A({ S25957[895] }),
  .B1({ S4233 }),
  .B2({ S4276 }),
  .ZN({ S4278 })
);
NAND2_X1 #() 
NAND2_X1_5480_ (
  .A1({ S4277 }),
  .A2({ S4278 }),
  .ZN({ S25957[767] })
);
NAND2_X1 #() 
NAND2_X1_5481_ (
  .A1({ S25957[767] }),
  .A2({ S25957[863] }),
  .ZN({ S4279 })
);
NAND3_X1 #() 
NAND3_X1_5957_ (
  .A1({ S4277 }),
  .A2({ S1733 }),
  .A3({ S4278 }),
  .ZN({ S4280 })
);
NAND2_X1 #() 
NAND2_X1_5482_ (
  .A1({ S4279 }),
  .A2({ S4280 }),
  .ZN({ S4281 })
);
INV_X1 #() 
INV_X1_1785_ (
  .A({ S4281 }),
  .ZN({ S25957[735] })
);
NAND2_X1 #() 
NAND2_X1_5483_ (
  .A1({ S25957[735] }),
  .A2({ S25957[927] }),
  .ZN({ S4282 })
);
NAND2_X1 #() 
NAND2_X1_5484_ (
  .A1({ S4281 }),
  .A2({ S24835 }),
  .ZN({ S4283 })
);
NAND2_X1 #() 
NAND2_X1_5485_ (
  .A1({ S4282 }),
  .A2({ S4283 }),
  .ZN({ S4284 })
);
INV_X1 #() 
INV_X1_1786_ (
  .A({ S4284 }),
  .ZN({ S25957[671] })
);
XOR2_X1 #() 
XOR2_X1_94_ (
  .A({ S25957[990] }),
  .B({ S25957[1086] }),
  .Z({ S25957[958] })
);
AOI22_X1 #() 
AOI22_X1_621_ (
  .A1({ S344 }),
  .A2({ S352 }),
  .B1({ S2748 }),
  .B2({ S2747 }),
  .ZN({ S4285 })
);
AOI21_X1 #() 
AOI21_X1_3122_ (
  .A({ S98 }),
  .B1({ S4285 }),
  .B2({ S4249 }),
  .ZN({ S4286 })
);
NAND2_X1 #() 
NAND2_X1_5486_ (
  .A1({ S4286 }),
  .A2({ S4166 }),
  .ZN({ S4287 })
);
NAND3_X1 #() 
NAND3_X1_5958_ (
  .A1({ S4287 }),
  .A2({ S25957[788] }),
  .A3({ S4207 }),
  .ZN({ S4288 })
);
INV_X1 #() 
INV_X1_1787_ (
  .A({ S4197 }),
  .ZN({ S4289 })
);
OAI22_X1 #() 
OAI22_X1_138_ (
  .A1({ S4184 }),
  .A2({ S4181 }),
  .B1({ S4191 }),
  .B2({ S4289 }),
  .ZN({ S4290 })
);
OAI21_X1 #() 
OAI21_X1_2852_ (
  .A({ S4288 }),
  .B1({ S4290 }),
  .B2({ S25957[788] }),
  .ZN({ S4291 })
);
AOI21_X1 #() 
AOI21_X1_3123_ (
  .A({ S4255 }),
  .B1({ S4259 }),
  .B2({ S4214 }),
  .ZN({ S4292 })
);
NAND4_X1 #() 
NAND4_X1_649_ (
  .A1({ S25957[786] }),
  .A2({ S2749 }),
  .A3({ S4164 }),
  .A4({ S4165 }),
  .ZN({ S4293 })
);
NAND3_X1 #() 
NAND3_X1_5959_ (
  .A1({ S4293 }),
  .A2({ S4213 }),
  .A3({ S4180 }),
  .ZN({ S4294 })
);
AOI21_X1 #() 
AOI21_X1_3124_ (
  .A({ S25957[788] }),
  .B1({ S4294 }),
  .B2({ S25957[787] }),
  .ZN({ S4295 })
);
AOI21_X1 #() 
AOI21_X1_3125_ (
  .A({ S4295 }),
  .B1({ S4292 }),
  .B2({ S25957[788] }),
  .ZN({ S4296 })
);
NAND2_X1 #() 
NAND2_X1_5487_ (
  .A1({ S4296 }),
  .A2({ S25673 }),
  .ZN({ S4297 })
);
OAI211_X1 #() 
OAI211_X1_1950_ (
  .A({ S4297 }),
  .B({ S25607 }),
  .C1({ S25673 }),
  .C2({ S4291 }),
  .ZN({ S4298 })
);
NAND3_X1 #() 
NAND3_X1_5960_ (
  .A1({ S25957[787] }),
  .A2({ S25957[785] }),
  .A3({ S4170 }),
  .ZN({ S4299 })
);
NAND2_X1 #() 
NAND2_X1_5488_ (
  .A1({ S4213 }),
  .A2({ S98 }),
  .ZN({ S4300 })
);
OAI21_X1 #() 
OAI21_X1_2853_ (
  .A({ S4299 }),
  .B1({ S4300 }),
  .B2({ S25957[784] }),
  .ZN({ S4301 })
);
OAI211_X1 #() 
OAI211_X1_1951_ (
  .A({ S4186 }),
  .B({ S4180 }),
  .C1({ S4249 }),
  .C2({ S4170 }),
  .ZN({ S4302 })
);
AOI21_X1 #() 
AOI21_X1_3126_ (
  .A({ S25957[788] }),
  .B1({ S4302 }),
  .B2({ S25957[787] }),
  .ZN({ S4303 })
);
OAI21_X1 #() 
OAI21_X1_2854_ (
  .A({ S4303 }),
  .B1({ S25957[787] }),
  .B2({ S4179 }),
  .ZN({ S4304 })
);
OAI21_X1 #() 
OAI21_X1_2855_ (
  .A({ S4304 }),
  .B1({ S2524 }),
  .B2({ S4301 }),
  .ZN({ S4305 })
);
NAND3_X1 #() 
NAND3_X1_5961_ (
  .A1({ S4210 }),
  .A2({ S4197 }),
  .A3({ S4180 }),
  .ZN({ S4306 })
);
NAND2_X1 #() 
NAND2_X1_5489_ (
  .A1({ S4177 }),
  .A2({ S4218 }),
  .ZN({ S4307 })
);
NAND2_X1 #() 
NAND2_X1_5490_ (
  .A1({ S4307 }),
  .A2({ S25957[787] }),
  .ZN({ S4308 })
);
NAND3_X1 #() 
NAND3_X1_5962_ (
  .A1({ S4308 }),
  .A2({ S4306 }),
  .A3({ S25957[788] }),
  .ZN({ S4309 })
);
AOI21_X1 #() 
AOI21_X1_3127_ (
  .A({ S25957[788] }),
  .B1({ S4222 }),
  .B2({ S4211 }),
  .ZN({ S4310 })
);
NOR2_X1 #() 
NOR2_X1_1382_ (
  .A1({ S4310 }),
  .A2({ S25673 }),
  .ZN({ S4311 })
);
AOI22_X1 #() 
AOI22_X1_622_ (
  .A1({ S4305 }),
  .A2({ S25673 }),
  .B1({ S4309 }),
  .B2({ S4311 }),
  .ZN({ S4312 })
);
OAI21_X1 #() 
OAI21_X1_2856_ (
  .A({ S4298 }),
  .B1({ S25607 }),
  .B2({ S4312 }),
  .ZN({ S4313 })
);
NOR2_X1 #() 
NOR2_X1_1383_ (
  .A1({ S4220 }),
  .A2({ S25957[788] }),
  .ZN({ S4314 })
);
NAND2_X1 #() 
NAND2_X1_5491_ (
  .A1({ S4302 }),
  .A2({ S25957[787] }),
  .ZN({ S4315 })
);
NAND3_X1 #() 
NAND3_X1_5963_ (
  .A1({ S4183 }),
  .A2({ S98 }),
  .A3({ S4218 }),
  .ZN({ S4316 })
);
AND3_X1 #() 
AND3_X1_241_ (
  .A1({ S4315 }),
  .A2({ S4316 }),
  .A3({ S4299 }),
  .ZN({ S4317 })
);
AOI22_X1 #() 
AOI22_X1_623_ (
  .A1({ S4317 }),
  .A2({ S25957[788] }),
  .B1({ S4198 }),
  .B2({ S4314 }),
  .ZN({ S4318 })
);
NAND2_X1 #() 
NAND2_X1_5492_ (
  .A1({ S4204 }),
  .A2({ S4210 }),
  .ZN({ S4319 })
);
AND2_X1 #() 
AND2_X1_349_ (
  .A1({ S4319 }),
  .A2({ S4315 }),
  .ZN({ S4320 })
);
NAND3_X1 #() 
NAND3_X1_5964_ (
  .A1({ S4197 }),
  .A2({ S4190 }),
  .A3({ S4259 }),
  .ZN({ S4321 })
);
OAI21_X1 #() 
OAI21_X1_2857_ (
  .A({ S25957[787] }),
  .B1({ S4263 }),
  .B2({ S4193 }),
  .ZN({ S4322 })
);
NAND3_X1 #() 
NAND3_X1_5965_ (
  .A1({ S4322 }),
  .A2({ S2524 }),
  .A3({ S4321 }),
  .ZN({ S4323 })
);
OAI211_X1 #() 
OAI211_X1_1952_ (
  .A({ S4323 }),
  .B({ S25673 }),
  .C1({ S2524 }),
  .C2({ S4320 }),
  .ZN({ S4324 })
);
OAI21_X1 #() 
OAI21_X1_2858_ (
  .A({ S4324 }),
  .B1({ S25673 }),
  .B2({ S4318 }),
  .ZN({ S4325 })
);
NAND2_X1 #() 
NAND2_X1_5493_ (
  .A1({ S4325 }),
  .A2({ S25957[790] }),
  .ZN({ S4326 })
);
NAND2_X1 #() 
NAND2_X1_5494_ (
  .A1({ S4177 }),
  .A2({ S4178 }),
  .ZN({ S4327 })
);
NAND2_X1 #() 
NAND2_X1_5495_ (
  .A1({ S4206 }),
  .A2({ S25957[787] }),
  .ZN({ S4328 })
);
NAND2_X1 #() 
NAND2_X1_5496_ (
  .A1({ S4213 }),
  .A2({ S4180 }),
  .ZN({ S4329 })
);
NAND2_X1 #() 
NAND2_X1_5497_ (
  .A1({ S4329 }),
  .A2({ S25957[787] }),
  .ZN({ S4330 })
);
OAI211_X1 #() 
OAI211_X1_1953_ (
  .A({ S4330 }),
  .B({ S4328 }),
  .C1({ S4207 }),
  .C2({ S4327 }),
  .ZN({ S4331 })
);
NAND4_X1 #() 
NAND4_X1_650_ (
  .A1({ S4170 }),
  .A2({ S4165 }),
  .A3({ S4164 }),
  .A4({ S2749 }),
  .ZN({ S4332 })
);
OAI21_X1 #() 
OAI21_X1_2859_ (
  .A({ S4328 }),
  .B1({ S25957[787] }),
  .B2({ S4332 }),
  .ZN({ S4333 })
);
OAI21_X1 #() 
OAI21_X1_2860_ (
  .A({ S25957[788] }),
  .B1({ S4333 }),
  .B2({ S4271 }),
  .ZN({ S4334 })
);
OAI21_X1 #() 
OAI21_X1_2861_ (
  .A({ S4334 }),
  .B1({ S25957[788] }),
  .B2({ S4331 }),
  .ZN({ S4335 })
);
AOI21_X1 #() 
AOI21_X1_3128_ (
  .A({ S98 }),
  .B1({ S4293 }),
  .B2({ S4180 }),
  .ZN({ S4336 })
);
AOI21_X1 #() 
AOI21_X1_3129_ (
  .A({ S4336 }),
  .B1({ S4210 }),
  .B2({ S4204 }),
  .ZN({ S4337 })
);
NOR2_X1 #() 
NOR2_X1_1384_ (
  .A1({ S4254 }),
  .A2({ S25957[787] }),
  .ZN({ S4338 })
);
OAI221_X1 #() 
OAI221_X1_165_ (
  .A({ S25673 }),
  .B1({ S4226 }),
  .B2({ S4338 }),
  .C1({ S4337 }),
  .C2({ S25957[788] }),
  .ZN({ S4339 })
);
OAI21_X1 #() 
OAI21_X1_2862_ (
  .A({ S4339 }),
  .B1({ S25673 }),
  .B2({ S4335 }),
  .ZN({ S4340 })
);
INV_X1 #() 
INV_X1_1788_ (
  .A({ S4340 }),
  .ZN({ S4341 })
);
OAI21_X1 #() 
OAI21_X1_2863_ (
  .A({ S4326 }),
  .B1({ S25957[790] }),
  .B2({ S4341 }),
  .ZN({ S4342 })
);
OR2_X1 #() 
OR2_X1_71_ (
  .A1({ S4342 }),
  .A2({ S2361 }),
  .ZN({ S4343 })
);
OAI211_X1 #() 
OAI211_X1_1954_ (
  .A({ S4343 }),
  .B({ S1802 }),
  .C1({ S4313 }),
  .C2({ S25957[791] }),
  .ZN({ S4344 })
);
NAND2_X1 #() 
NAND2_X1_5498_ (
  .A1({ S4342 }),
  .A2({ S25957[791] }),
  .ZN({ S4345 })
);
NAND2_X1 #() 
NAND2_X1_5499_ (
  .A1({ S4313 }),
  .A2({ S2361 }),
  .ZN({ S4346 })
);
NAND3_X1 #() 
NAND3_X1_5966_ (
  .A1({ S4345 }),
  .A2({ S4346 }),
  .A3({ S25957[894] }),
  .ZN({ S4347 })
);
AOI21_X1 #() 
AOI21_X1_3130_ (
  .A({ S25957[958] }),
  .B1({ S4344 }),
  .B2({ S4347 }),
  .ZN({ S4348 })
);
NAND3_X1 #() 
NAND3_X1_5967_ (
  .A1({ S4344 }),
  .A2({ S4347 }),
  .A3({ S25957[958] }),
  .ZN({ S4349 })
);
INV_X1 #() 
INV_X1_1789_ (
  .A({ S4349 }),
  .ZN({ S4350 })
);
OAI21_X1 #() 
OAI21_X1_2864_ (
  .A({ S25957[798] }),
  .B1({ S4350 }),
  .B2({ S4348 }),
  .ZN({ S4351 })
);
INV_X1 #() 
INV_X1_1790_ (
  .A({ S4348 }),
  .ZN({ S4352 })
);
NAND3_X1 #() 
NAND3_X1_5968_ (
  .A1({ S4352 }),
  .A2({ S3523 }),
  .A3({ S4349 }),
  .ZN({ S4353 })
);
NAND2_X1 #() 
NAND2_X1_5500_ (
  .A1({ S4351 }),
  .A2({ S4353 }),
  .ZN({ S4354 })
);
INV_X1 #() 
INV_X1_1791_ (
  .A({ S4354 }),
  .ZN({ S25957[670] })
);
NOR2_X1 #() 
NOR2_X1_1385_ (
  .A1({ S1874 }),
  .A2({ S1875 }),
  .ZN({ S4355 })
);
INV_X1 #() 
INV_X1_1792_ (
  .A({ S4355 }),
  .ZN({ S25957[861] })
);
NAND2_X1 #() 
NAND2_X1_5501_ (
  .A1({ S24933 }),
  .A2({ S24965 }),
  .ZN({ S4356 })
);
XOR2_X1 #() 
XOR2_X1_95_ (
  .A({ S4356 }),
  .B({ S25957[1149] }),
  .Z({ S25957[1021] })
);
XNOR2_X1 #() 
XNOR2_X1_210_ (
  .A({ S1872 }),
  .B({ S25957[1021] }),
  .ZN({ S25957[893] })
);
AOI21_X1 #() 
AOI21_X1_3131_ (
  .A({ S4170 }),
  .B1({ S25957[785] }),
  .B2({ S2749 }),
  .ZN({ S4357 })
);
AOI21_X1 #() 
AOI21_X1_3132_ (
  .A({ S98 }),
  .B1({ S4357 }),
  .B2({ S4178 }),
  .ZN({ S4358 })
);
INV_X1 #() 
INV_X1_1793_ (
  .A({ S4180 }),
  .ZN({ S4359 })
);
AOI21_X1 #() 
AOI21_X1_3133_ (
  .A({ S25957[787] }),
  .B1({ S4359 }),
  .B2({ S25957[785] }),
  .ZN({ S4360 })
);
AOI21_X1 #() 
AOI21_X1_3134_ (
  .A({ S4360 }),
  .B1({ S4358 }),
  .B2({ S4194 }),
  .ZN({ S4361 })
);
NAND3_X1 #() 
NAND3_X1_5969_ (
  .A1({ S4166 }),
  .A2({ S2 }),
  .A3({ S4170 }),
  .ZN({ S4362 })
);
NOR2_X1 #() 
NOR2_X1_1386_ (
  .A1({ S4362 }),
  .A2({ S98 }),
  .ZN({ S4363 })
);
OAI21_X1 #() 
OAI21_X1_2865_ (
  .A({ S25957[788] }),
  .B1({ S4207 }),
  .B2({ S25957[785] }),
  .ZN({ S4364 })
);
OAI22_X1 #() 
OAI22_X1_139_ (
  .A1({ S4361 }),
  .A2({ S25957[788] }),
  .B1({ S4363 }),
  .B2({ S4364 }),
  .ZN({ S4365 })
);
NAND2_X1 #() 
NAND2_X1_5502_ (
  .A1({ S4365 }),
  .A2({ S25673 }),
  .ZN({ S4366 })
);
AOI21_X1 #() 
AOI21_X1_3135_ (
  .A({ S2749 }),
  .B1({ S4164 }),
  .B2({ S4165 }),
  .ZN({ S4367 })
);
OAI21_X1 #() 
OAI21_X1_2866_ (
  .A({ S98 }),
  .B1({ S4367 }),
  .B2({ S4285 }),
  .ZN({ S4368 })
);
OAI211_X1 #() 
OAI211_X1_1955_ (
  .A({ S4368 }),
  .B({ S25957[788] }),
  .C1({ S4236 }),
  .C2({ S98 }),
  .ZN({ S4369 })
);
NAND2_X1 #() 
NAND2_X1_5503_ (
  .A1({ S4197 }),
  .A2({ S4166 }),
  .ZN({ S4370 })
);
NAND2_X1 #() 
NAND2_X1_5504_ (
  .A1({ S4370 }),
  .A2({ S98 }),
  .ZN({ S4371 })
);
NAND3_X1 #() 
NAND3_X1_5970_ (
  .A1({ S4371 }),
  .A2({ S2524 }),
  .A3({ S4223 }),
  .ZN({ S4372 })
);
NAND3_X1 #() 
NAND3_X1_5971_ (
  .A1({ S4369 }),
  .A2({ S4372 }),
  .A3({ S25957[789] }),
  .ZN({ S4373 })
);
AOI21_X1 #() 
AOI21_X1_3136_ (
  .A({ S25957[790] }),
  .B1({ S4366 }),
  .B2({ S4373 }),
  .ZN({ S4374 })
);
OAI21_X1 #() 
OAI21_X1_2867_ (
  .A({ S25957[788] }),
  .B1({ S4357 }),
  .B2({ S25957[787] }),
  .ZN({ S4375 })
);
AOI21_X1 #() 
AOI21_X1_3137_ (
  .A({ S4375 }),
  .B1({ S4329 }),
  .B2({ S25957[787] }),
  .ZN({ S4376 })
);
AOI21_X1 #() 
AOI21_X1_3138_ (
  .A({ S25957[788] }),
  .B1({ S4315 }),
  .B2({ S4270 }),
  .ZN({ S4377 })
);
OAI21_X1 #() 
OAI21_X1_2868_ (
  .A({ S25673 }),
  .B1({ S4376 }),
  .B2({ S4377 }),
  .ZN({ S4378 })
);
NAND2_X1 #() 
NAND2_X1_5505_ (
  .A1({ S4177 }),
  .A2({ S25957[786] }),
  .ZN({ S4379 })
);
AOI21_X1 #() 
AOI21_X1_3139_ (
  .A({ S98 }),
  .B1({ S4379 }),
  .B2({ S4262 }),
  .ZN({ S4380 })
);
AOI22_X1 #() 
AOI22_X1_624_ (
  .A1({ S25957[786] }),
  .A2({ S25957[784] }),
  .B1({ S4164 }),
  .B2({ S4165 }),
  .ZN({ S4381 })
);
OAI21_X1 #() 
OAI21_X1_2869_ (
  .A({ S2524 }),
  .B1({ S4381 }),
  .B2({ S25957[787] }),
  .ZN({ S4382 })
);
NAND2_X1 #() 
NAND2_X1_5506_ (
  .A1({ S4190 }),
  .A2({ S4174 }),
  .ZN({ S4383 })
);
NAND4_X1 #() 
NAND4_X1_651_ (
  .A1({ S25828 }),
  .A2({ S25833 }),
  .A3({ S25918 }),
  .A4({ S25924 }),
  .ZN({ S4384 })
);
NAND2_X1 #() 
NAND2_X1_5507_ (
  .A1({ S4293 }),
  .A2({ S98 }),
  .ZN({ S4385 })
);
OAI22_X1 #() 
OAI22_X1_140_ (
  .A1({ S4385 }),
  .A2({ S4383 }),
  .B1({ S4384 }),
  .B2({ S4214 }),
  .ZN({ S4386 })
);
AOI21_X1 #() 
AOI21_X1_3140_ (
  .A({ S25673 }),
  .B1({ S4386 }),
  .B2({ S25957[788] }),
  .ZN({ S4387 })
);
OAI21_X1 #() 
OAI21_X1_2870_ (
  .A({ S4387 }),
  .B1({ S4380 }),
  .B2({ S4382 }),
  .ZN({ S4388 })
);
AOI21_X1 #() 
AOI21_X1_3141_ (
  .A({ S25607 }),
  .B1({ S4388 }),
  .B2({ S4378 }),
  .ZN({ S4389 })
);
OAI21_X1 #() 
OAI21_X1_2871_ (
  .A({ S25957[791] }),
  .B1({ S4374 }),
  .B2({ S4389 }),
  .ZN({ S4390 })
);
OAI21_X1 #() 
OAI21_X1_2872_ (
  .A({ S4384 }),
  .B1({ S4199 }),
  .B2({ S4359 }),
  .ZN({ S4391 })
);
NAND2_X1 #() 
NAND2_X1_5508_ (
  .A1({ S4391 }),
  .A2({ S2524 }),
  .ZN({ S4392 })
);
NAND3_X1 #() 
NAND3_X1_5972_ (
  .A1({ S4177 }),
  .A2({ S4178 }),
  .A3({ S25957[786] }),
  .ZN({ S4393 })
);
NAND3_X1 #() 
NAND3_X1_5973_ (
  .A1({ S4393 }),
  .A2({ S25957[787] }),
  .A3({ S4332 }),
  .ZN({ S4394 })
);
NAND3_X1 #() 
NAND3_X1_5974_ (
  .A1({ S4254 }),
  .A2({ S98 }),
  .A3({ S4197 }),
  .ZN({ S4395 })
);
NAND3_X1 #() 
NAND3_X1_5975_ (
  .A1({ S4394 }),
  .A2({ S25957[788] }),
  .A3({ S4395 }),
  .ZN({ S4396 })
);
NAND3_X1 #() 
NAND3_X1_5976_ (
  .A1({ S4396 }),
  .A2({ S4392 }),
  .A3({ S25957[789] }),
  .ZN({ S4397 })
);
NAND3_X1 #() 
NAND3_X1_5977_ (
  .A1({ S4178 }),
  .A2({ S25957[787] }),
  .A3({ S4170 }),
  .ZN({ S4398 })
);
NAND4_X1 #() 
NAND4_X1_652_ (
  .A1({ S25957[786] }),
  .A2({ S25957[784] }),
  .A3({ S4164 }),
  .A4({ S4165 }),
  .ZN({ S4399 })
);
NAND3_X1 #() 
NAND3_X1_5978_ (
  .A1({ S4262 }),
  .A2({ S98 }),
  .A3({ S4399 }),
  .ZN({ S4400 })
);
NAND3_X1 #() 
NAND3_X1_5979_ (
  .A1({ S4400 }),
  .A2({ S25957[788] }),
  .A3({ S4398 }),
  .ZN({ S4401 })
);
INV_X1 #() 
INV_X1_1794_ (
  .A({ S4332 }),
  .ZN({ S4402 })
);
NOR2_X1 #() 
NOR2_X1_1387_ (
  .A1({ S4402 }),
  .A2({ S4221 }),
  .ZN({ S4403 })
);
NAND2_X1 #() 
NAND2_X1_5509_ (
  .A1({ S25957[787] }),
  .A2({ S4180 }),
  .ZN({ S4404 })
);
NOR2_X1 #() 
NOR2_X1_1388_ (
  .A1({ S4253 }),
  .A2({ S4404 }),
  .ZN({ S4405 })
);
AOI21_X1 #() 
AOI21_X1_3142_ (
  .A({ S4405 }),
  .B1({ S4403 }),
  .B2({ S98 }),
  .ZN({ S4406 })
);
OAI211_X1 #() 
OAI211_X1_1956_ (
  .A({ S25673 }),
  .B({ S4401 }),
  .C1({ S4406 }),
  .C2({ S25957[788] }),
  .ZN({ S4407 })
);
NAND3_X1 #() 
NAND3_X1_5980_ (
  .A1({ S4407 }),
  .A2({ S25957[790] }),
  .A3({ S4397 }),
  .ZN({ S4408 })
);
OAI21_X1 #() 
OAI21_X1_2873_ (
  .A({ S98 }),
  .B1({ S4249 }),
  .B2({ S4174 }),
  .ZN({ S4409 })
);
OAI21_X1 #() 
OAI21_X1_2874_ (
  .A({ S4409 }),
  .B1({ S4262 }),
  .B2({ S98 }),
  .ZN({ S4410 })
);
NAND2_X1 #() 
NAND2_X1_5510_ (
  .A1({ S4410 }),
  .A2({ S25957[788] }),
  .ZN({ S4411 })
);
NAND2_X1 #() 
NAND2_X1_5511_ (
  .A1({ S4186 }),
  .A2({ S98 }),
  .ZN({ S4412 })
);
NAND2_X1 #() 
NAND2_X1_5512_ (
  .A1({ S4222 }),
  .A2({ S4412 }),
  .ZN({ S4413 })
);
NAND2_X1 #() 
NAND2_X1_5513_ (
  .A1({ S4310 }),
  .A2({ S4413 }),
  .ZN({ S4414 })
);
AOI21_X1 #() 
AOI21_X1_3143_ (
  .A({ S25673 }),
  .B1({ S4414 }),
  .B2({ S4411 }),
  .ZN({ S4415 })
);
AOI211_X1 #() 
AOI211_X1_93_ (
  .A({ S98 }),
  .B({ S4181 }),
  .C1({ S4357 }),
  .C2({ S4178 }),
  .ZN({ S4416 })
);
NAND4_X1 #() 
NAND4_X1_653_ (
  .A1({ S4178 }),
  .A2({ S4177 }),
  .A3({ S4174 }),
  .A4({ S98 }),
  .ZN({ S4417 })
);
NAND2_X1 #() 
NAND2_X1_5514_ (
  .A1({ S4417 }),
  .A2({ S25957[788] }),
  .ZN({ S4418 })
);
NOR3_X1 #() 
NOR3_X1_176_ (
  .A1({ S4234 }),
  .A2({ S25957[788] }),
  .A3({ S2749 }),
  .ZN({ S4419 })
);
OAI21_X1 #() 
OAI21_X1_2875_ (
  .A({ S4419 }),
  .B1({ S4220 }),
  .B2({ S4224 }),
  .ZN({ S4420 })
);
OAI21_X1 #() 
OAI21_X1_2876_ (
  .A({ S4420 }),
  .B1({ S4416 }),
  .B2({ S4418 }),
  .ZN({ S4421 })
);
AOI21_X1 #() 
AOI21_X1_3144_ (
  .A({ S4415 }),
  .B1({ S25673 }),
  .B2({ S4421 }),
  .ZN({ S4422 })
);
OAI21_X1 #() 
OAI21_X1_2877_ (
  .A({ S4408 }),
  .B1({ S4422 }),
  .B2({ S25957[790] }),
  .ZN({ S4423 })
);
NAND2_X1 #() 
NAND2_X1_5515_ (
  .A1({ S4423 }),
  .A2({ S2361 }),
  .ZN({ S4424 })
);
NAND2_X1 #() 
NAND2_X1_5516_ (
  .A1({ S4390 }),
  .A2({ S4424 }),
  .ZN({ S4425 })
);
NAND2_X1 #() 
NAND2_X1_5517_ (
  .A1({ S4425 }),
  .A2({ S25957[893] }),
  .ZN({ S4426 })
);
INV_X1 #() 
INV_X1_1795_ (
  .A({ S25957[893] }),
  .ZN({ S4427 })
);
NAND3_X1 #() 
NAND3_X1_5981_ (
  .A1({ S4390 }),
  .A2({ S4424 }),
  .A3({ S4427 }),
  .ZN({ S4428 })
);
NAND3_X1 #() 
NAND3_X1_5982_ (
  .A1({ S4426 }),
  .A2({ S4428 }),
  .A3({ S25957[861] }),
  .ZN({ S4429 })
);
NAND2_X1 #() 
NAND2_X1_5518_ (
  .A1({ S4425 }),
  .A2({ S4427 }),
  .ZN({ S4430 })
);
NAND3_X1 #() 
NAND3_X1_5983_ (
  .A1({ S4390 }),
  .A2({ S4424 }),
  .A3({ S25957[893] }),
  .ZN({ S4431 })
);
NAND3_X1 #() 
NAND3_X1_5984_ (
  .A1({ S4430 }),
  .A2({ S4431 }),
  .A3({ S4355 }),
  .ZN({ S4432 })
);
NAND3_X1 #() 
NAND3_X1_5985_ (
  .A1({ S4429 }),
  .A2({ S4432 }),
  .A3({ S25957[925] }),
  .ZN({ S4433 })
);
NAND3_X1 #() 
NAND3_X1_5986_ (
  .A1({ S4430 }),
  .A2({ S4431 }),
  .A3({ S25957[861] }),
  .ZN({ S4434 })
);
NAND3_X1 #() 
NAND3_X1_5987_ (
  .A1({ S4426 }),
  .A2({ S4428 }),
  .A3({ S4355 }),
  .ZN({ S4435 })
);
NAND3_X1 #() 
NAND3_X1_5988_ (
  .A1({ S4434 }),
  .A2({ S4435 }),
  .A3({ S1084 }),
  .ZN({ S4436 })
);
NAND2_X1 #() 
NAND2_X1_5519_ (
  .A1({ S4433 }),
  .A2({ S4436 }),
  .ZN({ S25957[669] })
);
NOR2_X1 #() 
NOR2_X1_1389_ (
  .A1({ S1945 }),
  .A2({ S1941 }),
  .ZN({ S25957[828] })
);
NOR2_X1 #() 
NOR2_X1_1390_ (
  .A1({ S1944 }),
  .A2({ S1943 }),
  .ZN({ S25957[860] })
);
NAND2_X1 #() 
NAND2_X1_5520_ (
  .A1({ S25069 }),
  .A2({ S25068 }),
  .ZN({ S25957[1020] })
);
NAND2_X1 #() 
NAND2_X1_5521_ (
  .A1({ S1909 }),
  .A2({ S1934 }),
  .ZN({ S4437 })
);
XOR2_X1 #() 
XOR2_X1_96_ (
  .A({ S4437 }),
  .B({ S25957[1020] }),
  .Z({ S4438 })
);
INV_X1 #() 
INV_X1_1796_ (
  .A({ S4438 }),
  .ZN({ S25957[892] })
);
NAND2_X1 #() 
NAND2_X1_5522_ (
  .A1({ S4362 }),
  .A2({ S4379 }),
  .ZN({ S4439 })
);
AOI21_X1 #() 
AOI21_X1_3145_ (
  .A({ S4405 }),
  .B1({ S98 }),
  .B2({ S4439 }),
  .ZN({ S4440 })
);
AND2_X1 #() 
AND2_X1_350_ (
  .A1({ S4170 }),
  .A2({ S135 }),
  .ZN({ S4441 })
);
AOI21_X1 #() 
AOI21_X1_3146_ (
  .A({ S25673 }),
  .B1({ S25957[788] }),
  .B2({ S4441 }),
  .ZN({ S4442 })
);
OAI21_X1 #() 
OAI21_X1_2878_ (
  .A({ S4442 }),
  .B1({ S4440 }),
  .B2({ S25957[788] }),
  .ZN({ S4443 })
);
AOI21_X1 #() 
AOI21_X1_3147_ (
  .A({ S25957[787] }),
  .B1({ S4192 }),
  .B2({ S4190 }),
  .ZN({ S4444 })
);
NOR2_X1 #() 
NOR2_X1_1391_ (
  .A1({ S4226 }),
  .A2({ S4444 }),
  .ZN({ S4445 })
);
OAI211_X1 #() 
OAI211_X1_1957_ (
  .A({ S25828 }),
  .B({ S25833 }),
  .C1({ S4169 }),
  .C2({ S4168 }),
  .ZN({ S4446 })
);
INV_X1 #() 
INV_X1_1797_ (
  .A({ S4446 }),
  .ZN({ S4447 })
);
AOI211_X1 #() 
AOI211_X1_94_ (
  .A({ S4447 }),
  .B({ S25957[788] }),
  .C1({ S4360 }),
  .C2({ S4186 }),
  .ZN({ S4448 })
);
OAI21_X1 #() 
OAI21_X1_2879_ (
  .A({ S25673 }),
  .B1({ S4445 }),
  .B2({ S4448 }),
  .ZN({ S4449 })
);
NAND3_X1 #() 
NAND3_X1_5989_ (
  .A1({ S4449 }),
  .A2({ S4443 }),
  .A3({ S25957[790] }),
  .ZN({ S4450 })
);
NAND2_X1 #() 
NAND2_X1_5523_ (
  .A1({ S4259 }),
  .A2({ S25957[785] }),
  .ZN({ S4451 })
);
NAND2_X1 #() 
NAND2_X1_5524_ (
  .A1({ S4451 }),
  .A2({ S2524 }),
  .ZN({ S4452 })
);
OAI22_X1 #() 
OAI22_X1_141_ (
  .A1({ S4375 }),
  .A2({ S4255 }),
  .B1({ S4363 }),
  .B2({ S4452 }),
  .ZN({ S4453 })
);
NAND2_X1 #() 
NAND2_X1_5525_ (
  .A1({ S4453 }),
  .A2({ S25957[789] }),
  .ZN({ S4454 })
);
AOI21_X1 #() 
AOI21_X1_3148_ (
  .A({ S98 }),
  .B1({ S25957[784] }),
  .B2({ S25957[786] }),
  .ZN({ S4455 })
);
OAI21_X1 #() 
OAI21_X1_2880_ (
  .A({ S98 }),
  .B1({ S4186 }),
  .B2({ S25957[785] }),
  .ZN({ S4456 })
);
INV_X1 #() 
INV_X1_1798_ (
  .A({ S4456 }),
  .ZN({ S4457 })
);
AOI22_X1 #() 
AOI22_X1_625_ (
  .A1({ S4457 }),
  .A2({ S4194 }),
  .B1({ S4455 }),
  .B2({ S2 }),
  .ZN({ S4458 })
);
NAND2_X1 #() 
NAND2_X1_5526_ (
  .A1({ S4254 }),
  .A2({ S4455 }),
  .ZN({ S4459 })
);
NAND3_X1 #() 
NAND3_X1_5990_ (
  .A1({ S4371 }),
  .A2({ S4459 }),
  .A3({ S25957[788] }),
  .ZN({ S4460 })
);
OAI211_X1 #() 
OAI211_X1_1958_ (
  .A({ S25673 }),
  .B({ S4460 }),
  .C1({ S4458 }),
  .C2({ S25957[788] }),
  .ZN({ S4461 })
);
NAND3_X1 #() 
NAND3_X1_5991_ (
  .A1({ S4454 }),
  .A2({ S4461 }),
  .A3({ S25607 }),
  .ZN({ S4462 })
);
NAND2_X1 #() 
NAND2_X1_5527_ (
  .A1({ S4450 }),
  .A2({ S4462 }),
  .ZN({ S4463 })
);
NAND2_X1 #() 
NAND2_X1_5528_ (
  .A1({ S4463 }),
  .A2({ S2361 }),
  .ZN({ S4464 })
);
NAND3_X1 #() 
NAND3_X1_5992_ (
  .A1({ S4456 }),
  .A2({ S4398 }),
  .A3({ S25957[788] }),
  .ZN({ S4465 })
);
NAND3_X1 #() 
NAND3_X1_5993_ (
  .A1({ S4190 }),
  .A2({ S98 }),
  .A3({ S2749 }),
  .ZN({ S4466 })
);
NOR2_X1 #() 
NOR2_X1_1392_ (
  .A1({ S4260 }),
  .A2({ S25957[788] }),
  .ZN({ S4467 })
);
AOI21_X1 #() 
AOI21_X1_3149_ (
  .A({ S25673 }),
  .B1({ S4467 }),
  .B2({ S4466 }),
  .ZN({ S4468 })
);
NAND2_X1 #() 
NAND2_X1_5529_ (
  .A1({ S4468 }),
  .A2({ S4465 }),
  .ZN({ S4469 })
);
OAI211_X1 #() 
OAI211_X1_1959_ (
  .A({ S4371 }),
  .B({ S25957[788] }),
  .C1({ S4223 }),
  .C2({ S4359 }),
  .ZN({ S4470 })
);
NAND2_X1 #() 
NAND2_X1_5530_ (
  .A1({ S4210 }),
  .A2({ S4213 }),
  .ZN({ S4471 })
);
NAND3_X1 #() 
NAND3_X1_5994_ (
  .A1({ S4471 }),
  .A2({ S4264 }),
  .A3({ S2524 }),
  .ZN({ S4472 })
);
NAND3_X1 #() 
NAND3_X1_5995_ (
  .A1({ S4470 }),
  .A2({ S25673 }),
  .A3({ S4472 }),
  .ZN({ S4473 })
);
NAND3_X1 #() 
NAND3_X1_5996_ (
  .A1({ S4469 }),
  .A2({ S25957[790] }),
  .A3({ S4473 }),
  .ZN({ S4474 })
);
AOI21_X1 #() 
AOI21_X1_3150_ (
  .A({ S25957[787] }),
  .B1({ S4204 }),
  .B2({ S4239 }),
  .ZN({ S4475 })
);
NAND3_X1 #() 
NAND3_X1_5997_ (
  .A1({ S4285 }),
  .A2({ S25957[787] }),
  .A3({ S25957[785] }),
  .ZN({ S4476 })
);
NAND2_X1 #() 
NAND2_X1_5531_ (
  .A1({ S4398 }),
  .A2({ S4476 }),
  .ZN({ S4477 })
);
OAI21_X1 #() 
OAI21_X1_2881_ (
  .A({ S2524 }),
  .B1({ S4475 }),
  .B2({ S4477 }),
  .ZN({ S4478 })
);
NAND2_X1 #() 
NAND2_X1_5532_ (
  .A1({ S4327 }),
  .A2({ S4172 }),
  .ZN({ S4479 })
);
NAND4_X1 #() 
NAND4_X1_654_ (
  .A1({ S4213 }),
  .A2({ S4166 }),
  .A3({ S98 }),
  .A4({ S4186 }),
  .ZN({ S4480 })
);
NAND3_X1 #() 
NAND3_X1_5998_ (
  .A1({ S4479 }),
  .A2({ S25957[788] }),
  .A3({ S4480 }),
  .ZN({ S4481 })
);
AOI21_X1 #() 
AOI21_X1_3151_ (
  .A({ S25673 }),
  .B1({ S4478 }),
  .B2({ S4481 }),
  .ZN({ S4482 })
);
OAI221_X1 #() 
OAI221_X1_166_ (
  .A({ S2524 }),
  .B1({ S4223 }),
  .B2({ S4221 }),
  .C1({ S4409 }),
  .C2({ S4357 }),
  .ZN({ S4483 })
);
NAND3_X1 #() 
NAND3_X1_5999_ (
  .A1({ S4455 }),
  .A2({ S4197 }),
  .A3({ S4190 }),
  .ZN({ S4484 })
);
OAI211_X1 #() 
OAI211_X1_1960_ (
  .A({ S4484 }),
  .B({ S25957[788] }),
  .C1({ S4250 }),
  .C2({ S4267 }),
  .ZN({ S4485 })
);
NAND3_X1 #() 
NAND3_X1_6000_ (
  .A1({ S4485 }),
  .A2({ S4483 }),
  .A3({ S25673 }),
  .ZN({ S4486 })
);
NAND2_X1 #() 
NAND2_X1_5533_ (
  .A1({ S4486 }),
  .A2({ S25607 }),
  .ZN({ S4487 })
);
OAI211_X1 #() 
OAI211_X1_1961_ (
  .A({ S4474 }),
  .B({ S25957[791] }),
  .C1({ S4482 }),
  .C2({ S4487 }),
  .ZN({ S4488 })
);
NAND3_X1 #() 
NAND3_X1_6001_ (
  .A1({ S4464 }),
  .A2({ S4488 }),
  .A3({ S25957[892] }),
  .ZN({ S4489 })
);
OAI21_X1 #() 
OAI21_X1_2882_ (
  .A({ S4474 }),
  .B1({ S4482 }),
  .B2({ S4487 }),
  .ZN({ S4490 })
);
NAND2_X1 #() 
NAND2_X1_5534_ (
  .A1({ S4490 }),
  .A2({ S25957[791] }),
  .ZN({ S4491 })
);
NAND3_X1 #() 
NAND3_X1_6002_ (
  .A1({ S4450 }),
  .A2({ S4462 }),
  .A3({ S2361 }),
  .ZN({ S4492 })
);
NAND3_X1 #() 
NAND3_X1_6003_ (
  .A1({ S4491 }),
  .A2({ S4492 }),
  .A3({ S4438 }),
  .ZN({ S4493 })
);
NAND2_X1 #() 
NAND2_X1_5535_ (
  .A1({ S4493 }),
  .A2({ S4489 }),
  .ZN({ S25957[764] })
);
NAND2_X1 #() 
NAND2_X1_5536_ (
  .A1({ S25957[764] }),
  .A2({ S25957[860] }),
  .ZN({ S4494 })
);
INV_X1 #() 
INV_X1_1799_ (
  .A({ S25957[860] }),
  .ZN({ S4495 })
);
NAND3_X1 #() 
NAND3_X1_6004_ (
  .A1({ S4493 }),
  .A2({ S4489 }),
  .A3({ S4495 }),
  .ZN({ S4496 })
);
NAND3_X1 #() 
NAND3_X1_6005_ (
  .A1({ S4494 }),
  .A2({ S4496 }),
  .A3({ S25072 }),
  .ZN({ S4497 })
);
NAND3_X1 #() 
NAND3_X1_6006_ (
  .A1({ S4464 }),
  .A2({ S4488 }),
  .A3({ S4438 }),
  .ZN({ S4498 })
);
NAND3_X1 #() 
NAND3_X1_6007_ (
  .A1({ S4491 }),
  .A2({ S4492 }),
  .A3({ S25957[892] }),
  .ZN({ S4499 })
);
NAND3_X1 #() 
NAND3_X1_6008_ (
  .A1({ S4499 }),
  .A2({ S4498 }),
  .A3({ S4495 }),
  .ZN({ S4500 })
);
NAND3_X1 #() 
NAND3_X1_6009_ (
  .A1({ S4493 }),
  .A2({ S4489 }),
  .A3({ S25957[860] }),
  .ZN({ S4501 })
);
NAND3_X1 #() 
NAND3_X1_6010_ (
  .A1({ S4500 }),
  .A2({ S4501 }),
  .A3({ S25957[924] }),
  .ZN({ S4502 })
);
NAND2_X1 #() 
NAND2_X1_5537_ (
  .A1({ S4497 }),
  .A2({ S4502 }),
  .ZN({ S25957[668] })
);
NAND2_X1 #() 
NAND2_X1_5538_ (
  .A1({ S25175 }),
  .A2({ S25172 }),
  .ZN({ S4503 })
);
NAND2_X1 #() 
NAND2_X1_5539_ (
  .A1({ S25163 }),
  .A2({ S25162 }),
  .ZN({ S25957[1019] })
);
XOR2_X1 #() 
XOR2_X1_97_ (
  .A({ S2000 }),
  .B({ S25957[1019] }),
  .Z({ S4504 })
);
INV_X1 #() 
INV_X1_1800_ (
  .A({ S4504 }),
  .ZN({ S25957[891] })
);
NAND2_X1 #() 
NAND2_X1_5540_ (
  .A1({ S4302 }),
  .A2({ S98 }),
  .ZN({ S4505 })
);
AOI21_X1 #() 
AOI21_X1_3152_ (
  .A({ S2524 }),
  .B1({ S4362 }),
  .B2({ S4286 }),
  .ZN({ S4506 })
);
NAND3_X1 #() 
NAND3_X1_6011_ (
  .A1({ S4203 }),
  .A2({ S98 }),
  .A3({ S4213 }),
  .ZN({ S4507 })
);
AOI22_X1 #() 
AOI22_X1_626_ (
  .A1({ S4170 }),
  .A2({ S25957[784] }),
  .B1({ S261 }),
  .B2({ S267 }),
  .ZN({ S4508 })
);
AOI21_X1 #() 
AOI21_X1_3153_ (
  .A({ S25957[788] }),
  .B1({ S4172 }),
  .B2({ S4508 }),
  .ZN({ S4509 })
);
AOI22_X1 #() 
AOI22_X1_627_ (
  .A1({ S4506 }),
  .A2({ S4505 }),
  .B1({ S4507 }),
  .B2({ S4509 }),
  .ZN({ S4510 })
);
NAND2_X1 #() 
NAND2_X1_5541_ (
  .A1({ S4307 }),
  .A2({ S98 }),
  .ZN({ S4511 })
);
INV_X1 #() 
INV_X1_1801_ (
  .A({ S4399 }),
  .ZN({ S4512 })
);
OAI21_X1 #() 
OAI21_X1_2883_ (
  .A({ S25957[787] }),
  .B1({ S4512 }),
  .B2({ S4381 }),
  .ZN({ S4513 })
);
NAND3_X1 #() 
NAND3_X1_6012_ (
  .A1({ S4513 }),
  .A2({ S4511 }),
  .A3({ S2524 }),
  .ZN({ S4514 })
);
NAND3_X1 #() 
NAND3_X1_6013_ (
  .A1({ S4190 }),
  .A2({ S98 }),
  .A3({ S4218 }),
  .ZN({ S4515 })
);
OAI211_X1 #() 
OAI211_X1_1962_ (
  .A({ S25957[788] }),
  .B({ S4515 }),
  .C1({ S4204 }),
  .C2({ S98 }),
  .ZN({ S4516 })
);
NAND3_X1 #() 
NAND3_X1_6014_ (
  .A1({ S4514 }),
  .A2({ S25673 }),
  .A3({ S4516 }),
  .ZN({ S4517 })
);
OAI211_X1 #() 
OAI211_X1_1963_ (
  .A({ S4517 }),
  .B({ S25607 }),
  .C1({ S4510 }),
  .C2({ S25673 }),
  .ZN({ S4518 })
);
NAND3_X1 #() 
NAND3_X1_6015_ (
  .A1({ S4183 }),
  .A2({ S4166 }),
  .A3({ S25957[787] }),
  .ZN({ S4519 })
);
NAND3_X1 #() 
NAND3_X1_6016_ (
  .A1({ S4393 }),
  .A2({ S98 }),
  .A3({ S4171 }),
  .ZN({ S4520 })
);
AOI21_X1 #() 
AOI21_X1_3154_ (
  .A({ S2524 }),
  .B1({ S4520 }),
  .B2({ S4519 }),
  .ZN({ S4521 })
);
NAND3_X1 #() 
NAND3_X1_6017_ (
  .A1({ S4307 }),
  .A2({ S2524 }),
  .A3({ S4446 }),
  .ZN({ S4522 })
);
NAND2_X1 #() 
NAND2_X1_5542_ (
  .A1({ S4522 }),
  .A2({ S25673 }),
  .ZN({ S4523 })
);
NAND4_X1 #() 
NAND4_X1_655_ (
  .A1({ S4213 }),
  .A2({ S4166 }),
  .A3({ S25957[787] }),
  .A4({ S4186 }),
  .ZN({ S4524 })
);
NAND3_X1 #() 
NAND3_X1_6018_ (
  .A1({ S4210 }),
  .A2({ S4177 }),
  .A3({ S4178 }),
  .ZN({ S4525 })
);
AOI21_X1 #() 
AOI21_X1_3155_ (
  .A({ S25957[788] }),
  .B1({ S4525 }),
  .B2({ S4524 }),
  .ZN({ S4526 })
);
NAND3_X1 #() 
NAND3_X1_6019_ (
  .A1({ S4293 }),
  .A2({ S98 }),
  .A3({ S4178 }),
  .ZN({ S4527 })
);
INV_X1 #() 
INV_X1_1802_ (
  .A({ S4527 }),
  .ZN({ S4528 })
);
AOI21_X1 #() 
AOI21_X1_3156_ (
  .A({ S25957[784] }),
  .B1({ S4164 }),
  .B2({ S4165 }),
  .ZN({ S4529 })
);
OAI21_X1 #() 
OAI21_X1_2884_ (
  .A({ S25957[788] }),
  .B1({ S4235 }),
  .B2({ S4529 }),
  .ZN({ S4530 })
);
OAI21_X1 #() 
OAI21_X1_2885_ (
  .A({ S25957[789] }),
  .B1({ S4528 }),
  .B2({ S4530 }),
  .ZN({ S4531 })
);
OAI22_X1 #() 
OAI22_X1_142_ (
  .A1({ S4521 }),
  .A2({ S4523 }),
  .B1({ S4531 }),
  .B2({ S4526 }),
  .ZN({ S4532 })
);
NAND2_X1 #() 
NAND2_X1_5543_ (
  .A1({ S4532 }),
  .A2({ S25957[790] }),
  .ZN({ S4533 })
);
NAND3_X1 #() 
NAND3_X1_6020_ (
  .A1({ S4533 }),
  .A2({ S4518 }),
  .A3({ S25957[791] }),
  .ZN({ S4534 })
);
AOI21_X1 #() 
AOI21_X1_3157_ (
  .A({ S98 }),
  .B1({ S4367 }),
  .B2({ S25957[786] }),
  .ZN({ S4535 })
);
AOI21_X1 #() 
AOI21_X1_3158_ (
  .A({ S25957[787] }),
  .B1({ S4190 }),
  .B2({ S25957[784] }),
  .ZN({ S4536 })
);
OAI21_X1 #() 
OAI21_X1_2886_ (
  .A({ S2524 }),
  .B1({ S4535 }),
  .B2({ S4536 }),
  .ZN({ S4537 })
);
OAI211_X1 #() 
OAI211_X1_1964_ (
  .A({ S4270 }),
  .B({ S25957[788] }),
  .C1({ S98 }),
  .C2({ S4192 }),
  .ZN({ S4538 })
);
NAND2_X1 #() 
NAND2_X1_5544_ (
  .A1({ S4537 }),
  .A2({ S4538 }),
  .ZN({ S4539 })
);
NAND2_X1 #() 
NAND2_X1_5545_ (
  .A1({ S4539 }),
  .A2({ S25957[789] }),
  .ZN({ S4540 })
);
NAND4_X1 #() 
NAND4_X1_656_ (
  .A1({ S4177 }),
  .A2({ S4178 }),
  .A3({ S25957[787] }),
  .A4({ S4218 }),
  .ZN({ S4541 })
);
OAI21_X1 #() 
OAI21_X1_2887_ (
  .A({ S4541 }),
  .B1({ S4181 }),
  .B2({ S4184 }),
  .ZN({ S4542 })
);
NAND2_X1 #() 
NAND2_X1_5546_ (
  .A1({ S4542 }),
  .A2({ S25957[788] }),
  .ZN({ S4543 })
);
NAND3_X1 #() 
NAND3_X1_6021_ (
  .A1({ S25957[785] }),
  .A2({ S25957[784] }),
  .A3({ S4170 }),
  .ZN({ S4544 })
);
AOI22_X1 #() 
AOI22_X1_628_ (
  .A1({ S4203 }),
  .A2({ S4241 }),
  .B1({ S4172 }),
  .B2({ S4544 }),
  .ZN({ S4545 })
);
NAND2_X1 #() 
NAND2_X1_5547_ (
  .A1({ S4545 }),
  .A2({ S2524 }),
  .ZN({ S4546 })
);
NAND3_X1 #() 
NAND3_X1_6022_ (
  .A1({ S4546 }),
  .A2({ S4543 }),
  .A3({ S25673 }),
  .ZN({ S4547 })
);
NAND3_X1 #() 
NAND3_X1_6023_ (
  .A1({ S4540 }),
  .A2({ S4547 }),
  .A3({ S25607 }),
  .ZN({ S4548 })
);
INV_X1 #() 
INV_X1_1803_ (
  .A({ S4315 }),
  .ZN({ S4549 })
);
NOR2_X1 #() 
NOR2_X1_1393_ (
  .A1({ S4268 }),
  .A2({ S4549 }),
  .ZN({ S4550 })
);
NAND3_X1 #() 
NAND3_X1_6024_ (
  .A1({ S4183 }),
  .A2({ S25957[787] }),
  .A3({ S2749 }),
  .ZN({ S4551 })
);
NAND3_X1 #() 
NAND3_X1_6025_ (
  .A1({ S4190 }),
  .A2({ S4178 }),
  .A3({ S98 }),
  .ZN({ S4552 })
);
NAND2_X1 #() 
NAND2_X1_5548_ (
  .A1({ S4551 }),
  .A2({ S4552 }),
  .ZN({ S4553 })
);
OAI21_X1 #() 
OAI21_X1_2888_ (
  .A({ S25957[789] }),
  .B1({ S4553 }),
  .B2({ S25957[788] }),
  .ZN({ S4554 })
);
NAND3_X1 #() 
NAND3_X1_6026_ (
  .A1({ S4166 }),
  .A2({ S98 }),
  .A3({ S4218 }),
  .ZN({ S4555 })
);
NAND2_X1 #() 
NAND2_X1_5549_ (
  .A1({ S4555 }),
  .A2({ S25957[788] }),
  .ZN({ S4556 })
);
NAND2_X1 #() 
NAND2_X1_5550_ (
  .A1({ S4173 }),
  .A2({ S4321 }),
  .ZN({ S4557 })
);
OAI211_X1 #() 
OAI211_X1_1965_ (
  .A({ S25673 }),
  .B({ S4556 }),
  .C1({ S4557 }),
  .C2({ S25957[788] }),
  .ZN({ S4558 })
);
OAI211_X1 #() 
OAI211_X1_1966_ (
  .A({ S4558 }),
  .B({ S25957[790] }),
  .C1({ S4550 }),
  .C2({ S4554 }),
  .ZN({ S4559 })
);
NAND3_X1 #() 
NAND3_X1_6027_ (
  .A1({ S4548 }),
  .A2({ S2361 }),
  .A3({ S4559 }),
  .ZN({ S4560 })
);
NAND3_X1 #() 
NAND3_X1_6028_ (
  .A1({ S4534 }),
  .A2({ S4560 }),
  .A3({ S25957[891] }),
  .ZN({ S4561 })
);
NOR2_X1 #() 
NOR2_X1_1394_ (
  .A1({ S4529 }),
  .A2({ S4207 }),
  .ZN({ S4562 })
);
NAND2_X1 #() 
NAND2_X1_5551_ (
  .A1({ S4218 }),
  .A2({ S4249 }),
  .ZN({ S4563 })
);
AOI21_X1 #() 
AOI21_X1_3159_ (
  .A({ S98 }),
  .B1({ S4563 }),
  .B2({ S4399 }),
  .ZN({ S4564 })
);
OAI21_X1 #() 
OAI21_X1_2889_ (
  .A({ S2524 }),
  .B1({ S4564 }),
  .B2({ S4562 }),
  .ZN({ S4565 })
);
NAND2_X1 #() 
NAND2_X1_5552_ (
  .A1({ S4204 }),
  .A2({ S25957[787] }),
  .ZN({ S4566 })
);
AOI21_X1 #() 
AOI21_X1_3160_ (
  .A({ S2524 }),
  .B1({ S4210 }),
  .B2({ S4213 }),
  .ZN({ S4567 })
);
AOI21_X1 #() 
AOI21_X1_3161_ (
  .A({ S25957[789] }),
  .B1({ S4566 }),
  .B2({ S4567 }),
  .ZN({ S4568 })
);
NAND2_X1 #() 
NAND2_X1_5553_ (
  .A1({ S4568 }),
  .A2({ S4565 }),
  .ZN({ S4569 })
);
NAND2_X1 #() 
NAND2_X1_5554_ (
  .A1({ S4506 }),
  .A2({ S4505 }),
  .ZN({ S4570 })
);
AOI21_X1 #() 
AOI21_X1_3162_ (
  .A({ S25673 }),
  .B1({ S4507 }),
  .B2({ S4509 }),
  .ZN({ S4571 })
);
NAND2_X1 #() 
NAND2_X1_5555_ (
  .A1({ S4571 }),
  .A2({ S4570 }),
  .ZN({ S4572 })
);
NAND3_X1 #() 
NAND3_X1_6029_ (
  .A1({ S4572 }),
  .A2({ S25607 }),
  .A3({ S4569 }),
  .ZN({ S4573 })
);
OAI211_X1 #() 
OAI211_X1_1967_ (
  .A({ S4573 }),
  .B({ S25957[791] }),
  .C1({ S25607 }),
  .C2({ S4532 }),
  .ZN({ S4574 })
);
AOI21_X1 #() 
AOI21_X1_3163_ (
  .A({ S25957[787] }),
  .B1({ S4213 }),
  .B2({ S25957[784] }),
  .ZN({ S4575 })
);
NAND2_X1 #() 
NAND2_X1_5556_ (
  .A1({ S4575 }),
  .A2({ S25957[788] }),
  .ZN({ S4576 })
);
NAND2_X1 #() 
NAND2_X1_5557_ (
  .A1({ S4557 }),
  .A2({ S2524 }),
  .ZN({ S4577 })
);
NAND3_X1 #() 
NAND3_X1_6030_ (
  .A1({ S4577 }),
  .A2({ S25673 }),
  .A3({ S4576 }),
  .ZN({ S4578 })
);
AOI22_X1 #() 
AOI22_X1_629_ (
  .A1({ S4360 }),
  .A2({ S4203 }),
  .B1({ S4302 }),
  .B2({ S25957[787] }),
  .ZN({ S4579 })
);
NAND2_X1 #() 
NAND2_X1_5558_ (
  .A1({ S4553 }),
  .A2({ S2524 }),
  .ZN({ S4580 })
);
OAI211_X1 #() 
OAI211_X1_1968_ (
  .A({ S4580 }),
  .B({ S25957[789] }),
  .C1({ S4579 }),
  .C2({ S2524 }),
  .ZN({ S4581 })
);
NAND3_X1 #() 
NAND3_X1_6031_ (
  .A1({ S4581 }),
  .A2({ S4578 }),
  .A3({ S25957[790] }),
  .ZN({ S4582 })
);
OAI211_X1 #() 
OAI211_X1_1969_ (
  .A({ S4541 }),
  .B({ S25957[788] }),
  .C1({ S4181 }),
  .C2({ S4184 }),
  .ZN({ S4583 })
);
OAI211_X1 #() 
OAI211_X1_1970_ (
  .A({ S4583 }),
  .B({ S25673 }),
  .C1({ S4545 }),
  .C2({ S25957[788] }),
  .ZN({ S4584 })
);
NAND3_X1 #() 
NAND3_X1_6032_ (
  .A1({ S4537 }),
  .A2({ S4538 }),
  .A3({ S25957[789] }),
  .ZN({ S4585 })
);
NAND3_X1 #() 
NAND3_X1_6033_ (
  .A1({ S4584 }),
  .A2({ S25607 }),
  .A3({ S4585 }),
  .ZN({ S4586 })
);
NAND3_X1 #() 
NAND3_X1_6034_ (
  .A1({ S4582 }),
  .A2({ S2361 }),
  .A3({ S4586 }),
  .ZN({ S4587 })
);
NAND3_X1 #() 
NAND3_X1_6035_ (
  .A1({ S4574 }),
  .A2({ S4587 }),
  .A3({ S4504 }),
  .ZN({ S4588 })
);
NAND3_X1 #() 
NAND3_X1_6036_ (
  .A1({ S4561 }),
  .A2({ S4588 }),
  .A3({ S4503 }),
  .ZN({ S4589 })
);
INV_X1 #() 
INV_X1_1804_ (
  .A({ S4503 }),
  .ZN({ S25957[955] })
);
NAND3_X1 #() 
NAND3_X1_6037_ (
  .A1({ S4574 }),
  .A2({ S4587 }),
  .A3({ S25957[891] }),
  .ZN({ S4590 })
);
NAND3_X1 #() 
NAND3_X1_6038_ (
  .A1({ S4534 }),
  .A2({ S4560 }),
  .A3({ S4504 }),
  .ZN({ S4591 })
);
NAND3_X1 #() 
NAND3_X1_6039_ (
  .A1({ S4591 }),
  .A2({ S4590 }),
  .A3({ S25957[955] }),
  .ZN({ S4592 })
);
NAND3_X1 #() 
NAND3_X1_6040_ (
  .A1({ S4589 }),
  .A2({ S4592 }),
  .A3({ S25957[795] }),
  .ZN({ S4593 })
);
NAND3_X1 #() 
NAND3_X1_6041_ (
  .A1({ S4561 }),
  .A2({ S4588 }),
  .A3({ S25957[955] }),
  .ZN({ S4594 })
);
NAND3_X1 #() 
NAND3_X1_6042_ (
  .A1({ S4591 }),
  .A2({ S4590 }),
  .A3({ S4503 }),
  .ZN({ S4595 })
);
NAND3_X1 #() 
NAND3_X1_6043_ (
  .A1({ S4594 }),
  .A2({ S4595 }),
  .A3({ S107 }),
  .ZN({ S4596 })
);
AND2_X1 #() 
AND2_X1_351_ (
  .A1({ S4596 }),
  .A2({ S4593 }),
  .ZN({ S3 })
);
NAND2_X1 #() 
NAND2_X1_5559_ (
  .A1({ S4593 }),
  .A2({ S4596 }),
  .ZN({ S25957[667] })
);
NAND2_X1 #() 
NAND2_X1_5560_ (
  .A1({ S25259 }),
  .A2({ S25262 }),
  .ZN({ S4597 })
);
NAND2_X1 #() 
NAND2_X1_5561_ (
  .A1({ S22515 }),
  .A2({ S22516 }),
  .ZN({ S25957[1144] })
);
NAND2_X1 #() 
NAND2_X1_5562_ (
  .A1({ S25239 }),
  .A2({ S25257 }),
  .ZN({ S4598 })
);
XNOR2_X1 #() 
XNOR2_X1_211_ (
  .A({ S4598 }),
  .B({ S25957[1144] }),
  .ZN({ S25957[1016] })
);
NAND2_X1 #() 
NAND2_X1_5563_ (
  .A1({ S2043 }),
  .A2({ S2024 }),
  .ZN({ S4599 })
);
XNOR2_X1 #() 
XNOR2_X1_212_ (
  .A({ S4599 }),
  .B({ S25957[1016] }),
  .ZN({ S25957[888] })
);
INV_X1 #() 
INV_X1_1805_ (
  .A({ S25957[888] }),
  .ZN({ S4600 })
);
NAND3_X1 #() 
NAND3_X1_6044_ (
  .A1({ S4456 }),
  .A2({ S4398 }),
  .A3({ S4476 }),
  .ZN({ S4601 })
);
NAND2_X1 #() 
NAND2_X1_5564_ (
  .A1({ S4601 }),
  .A2({ S2524 }),
  .ZN({ S4602 })
);
NAND3_X1 #() 
NAND3_X1_6045_ (
  .A1({ S4183 }),
  .A2({ S98 }),
  .A3({ S2749 }),
  .ZN({ S4603 })
);
OAI211_X1 #() 
OAI211_X1_1971_ (
  .A({ S25957[788] }),
  .B({ S4603 }),
  .C1({ S4575 }),
  .C2({ S4286 }),
  .ZN({ S4604 })
);
AND3_X1 #() 
AND3_X1_242_ (
  .A1({ S4602 }),
  .A2({ S25607 }),
  .A3({ S4604 }),
  .ZN({ S4605 })
);
OAI21_X1 #() 
OAI21_X1_2890_ (
  .A({ S98 }),
  .B1({ S4181 }),
  .B2({ S4508 }),
  .ZN({ S4606 })
);
NAND3_X1 #() 
NAND3_X1_6046_ (
  .A1({ S4606 }),
  .A2({ S2524 }),
  .A3({ S4459 }),
  .ZN({ S4607 })
);
AOI21_X1 #() 
AOI21_X1_3164_ (
  .A({ S2524 }),
  .B1({ S4447 }),
  .B2({ S4177 }),
  .ZN({ S4608 })
);
NAND2_X1 #() 
NAND2_X1_5565_ (
  .A1({ S4195 }),
  .A2({ S4608 }),
  .ZN({ S4609 })
);
AOI21_X1 #() 
AOI21_X1_3165_ (
  .A({ S25607 }),
  .B1({ S4607 }),
  .B2({ S4609 }),
  .ZN({ S4610 })
);
OAI21_X1 #() 
OAI21_X1_2891_ (
  .A({ S25957[789] }),
  .B1({ S4605 }),
  .B2({ S4610 }),
  .ZN({ S4611 })
);
NAND4_X1 #() 
NAND4_X1_657_ (
  .A1({ S2 }),
  .A2({ S98 }),
  .A3({ S4218 }),
  .A4({ S4174 }),
  .ZN({ S4612 })
);
AOI21_X1 #() 
AOI21_X1_3166_ (
  .A({ S25957[788] }),
  .B1({ S4612 }),
  .B2({ S4551 }),
  .ZN({ S4613 })
);
NAND4_X1 #() 
NAND4_X1_658_ (
  .A1({ S4166 }),
  .A2({ S2 }),
  .A3({ S98 }),
  .A4({ S4170 }),
  .ZN({ S4614 })
);
NAND2_X1 #() 
NAND2_X1_5566_ (
  .A1({ S4246 }),
  .A2({ S4614 }),
  .ZN({ S4615 })
);
NAND2_X1 #() 
NAND2_X1_5567_ (
  .A1({ S4615 }),
  .A2({ S25607 }),
  .ZN({ S4616 })
);
NAND3_X1 #() 
NAND3_X1_6047_ (
  .A1({ S4213 }),
  .A2({ S4166 }),
  .A3({ S4186 }),
  .ZN({ S4617 })
);
NAND2_X1 #() 
NAND2_X1_5568_ (
  .A1({ S4617 }),
  .A2({ S98 }),
  .ZN({ S4618 })
);
NAND3_X1 #() 
NAND3_X1_6048_ (
  .A1({ S4447 }),
  .A2({ S4177 }),
  .A3({ S4178 }),
  .ZN({ S4619 })
);
AOI21_X1 #() 
AOI21_X1_3167_ (
  .A({ S2524 }),
  .B1({ S4618 }),
  .B2({ S4619 }),
  .ZN({ S4620 })
);
NAND2_X1 #() 
NAND2_X1_5569_ (
  .A1({ S4446 }),
  .A2({ S4384 }),
  .ZN({ S4621 })
);
AOI22_X1 #() 
AOI22_X1_630_ (
  .A1({ S4239 }),
  .A2({ S4621 }),
  .B1({ S4332 }),
  .B2({ S98 }),
  .ZN({ S4622 })
);
OAI21_X1 #() 
OAI21_X1_2892_ (
  .A({ S25957[790] }),
  .B1({ S4622 }),
  .B2({ S25957[788] }),
  .ZN({ S4623 })
);
OAI22_X1 #() 
OAI22_X1_143_ (
  .A1({ S4623 }),
  .A2({ S4620 }),
  .B1({ S4616 }),
  .B2({ S4613 }),
  .ZN({ S4624 })
);
NAND2_X1 #() 
NAND2_X1_5570_ (
  .A1({ S4624 }),
  .A2({ S25673 }),
  .ZN({ S4625 })
);
NAND3_X1 #() 
NAND3_X1_6049_ (
  .A1({ S4611 }),
  .A2({ S25957[791] }),
  .A3({ S4625 }),
  .ZN({ S4626 })
);
NAND3_X1 #() 
NAND3_X1_6050_ (
  .A1({ S4393 }),
  .A2({ S25957[787] }),
  .A3({ S4262 }),
  .ZN({ S4627 })
);
NAND2_X1 #() 
NAND2_X1_5571_ (
  .A1({ S4213 }),
  .A2({ S2749 }),
  .ZN({ S4628 })
);
AOI21_X1 #() 
AOI21_X1_3168_ (
  .A({ S2524 }),
  .B1({ S4628 }),
  .B2({ S98 }),
  .ZN({ S4629 })
);
AOI22_X1 #() 
AOI22_X1_631_ (
  .A1({ S4295 }),
  .A2({ S4248 }),
  .B1({ S4627 }),
  .B2({ S4629 }),
  .ZN({ S4630 })
);
NAND4_X1 #() 
NAND4_X1_659_ (
  .A1({ S25957[788] }),
  .A2({ S4332 }),
  .A3({ S4197 }),
  .A4({ S4384 }),
  .ZN({ S4631 })
);
OAI211_X1 #() 
OAI211_X1_1972_ (
  .A({ S25673 }),
  .B({ S4631 }),
  .C1({ S4405 }),
  .C2({ S4382 }),
  .ZN({ S4632 })
);
OAI211_X1 #() 
OAI211_X1_1973_ (
  .A({ S25957[790] }),
  .B({ S4632 }),
  .C1({ S4630 }),
  .C2({ S25673 }),
  .ZN({ S4633 })
);
NAND2_X1 #() 
NAND2_X1_5572_ (
  .A1({ S4417 }),
  .A2({ S4191 }),
  .ZN({ S4634 })
);
OAI22_X1 #() 
OAI22_X1_144_ (
  .A1({ S4199 }),
  .A2({ S4359 }),
  .B1({ S4235 }),
  .B2({ S4529 }),
  .ZN({ S4635 })
);
AOI22_X1 #() 
AOI22_X1_632_ (
  .A1({ S4634 }),
  .A2({ S4303 }),
  .B1({ S4635 }),
  .B2({ S25957[788] }),
  .ZN({ S4636 })
);
AOI21_X1 #() 
AOI21_X1_3169_ (
  .A({ S25957[787] }),
  .B1({ S4563 }),
  .B2({ S4399 }),
  .ZN({ S4637 })
);
AOI22_X1 #() 
AOI22_X1_633_ (
  .A1({ S4213 }),
  .A2({ S4180 }),
  .B1({ S4249 }),
  .B2({ S25957[784] }),
  .ZN({ S4638 })
);
OAI21_X1 #() 
OAI21_X1_2893_ (
  .A({ S25957[788] }),
  .B1({ S4638 }),
  .B2({ S98 }),
  .ZN({ S4639 })
);
NAND4_X1 #() 
NAND4_X1_660_ (
  .A1({ S4177 }),
  .A2({ S4178 }),
  .A3({ S25957[787] }),
  .A4({ S4180 }),
  .ZN({ S4640 })
);
OAI211_X1 #() 
OAI211_X1_1974_ (
  .A({ S4640 }),
  .B({ S2524 }),
  .C1({ S4316 }),
  .C2({ S4383 }),
  .ZN({ S4641 })
);
OAI211_X1 #() 
OAI211_X1_1975_ (
  .A({ S4641 }),
  .B({ S25673 }),
  .C1({ S4639 }),
  .C2({ S4637 }),
  .ZN({ S4642 })
);
OAI211_X1 #() 
OAI211_X1_1976_ (
  .A({ S4642 }),
  .B({ S25607 }),
  .C1({ S4636 }),
  .C2({ S25673 }),
  .ZN({ S4643 })
);
NAND3_X1 #() 
NAND3_X1_6051_ (
  .A1({ S4643 }),
  .A2({ S4633 }),
  .A3({ S2361 }),
  .ZN({ S4644 })
);
NAND3_X1 #() 
NAND3_X1_6052_ (
  .A1({ S4626 }),
  .A2({ S4600 }),
  .A3({ S4644 }),
  .ZN({ S4645 })
);
AOI21_X1 #() 
AOI21_X1_3170_ (
  .A({ S25673 }),
  .B1({ S4195 }),
  .B2({ S4608 }),
  .ZN({ S4646 })
);
NAND2_X1 #() 
NAND2_X1_5573_ (
  .A1({ S4480 }),
  .A2({ S25957[788] }),
  .ZN({ S4647 })
);
OAI22_X1 #() 
OAI22_X1_145_ (
  .A1({ S4358 }),
  .A2({ S4647 }),
  .B1({ S4622 }),
  .B2({ S25957[788] }),
  .ZN({ S4648 })
);
AOI22_X1 #() 
AOI22_X1_634_ (
  .A1({ S4648 }),
  .A2({ S25673 }),
  .B1({ S4607 }),
  .B2({ S4646 }),
  .ZN({ S4649 })
);
AND2_X1 #() 
AND2_X1_352_ (
  .A1({ S4612 }),
  .A2({ S4551 }),
  .ZN({ S4650 })
);
OAI211_X1 #() 
OAI211_X1_1977_ (
  .A({ S25673 }),
  .B({ S4615 }),
  .C1({ S4650 }),
  .C2({ S25957[788] }),
  .ZN({ S4651 })
);
NAND3_X1 #() 
NAND3_X1_6053_ (
  .A1({ S4602 }),
  .A2({ S25957[789] }),
  .A3({ S4604 }),
  .ZN({ S4652 })
);
NAND3_X1 #() 
NAND3_X1_6054_ (
  .A1({ S4652 }),
  .A2({ S4651 }),
  .A3({ S25607 }),
  .ZN({ S4653 })
);
OAI211_X1 #() 
OAI211_X1_1978_ (
  .A({ S4653 }),
  .B({ S25957[791] }),
  .C1({ S4649 }),
  .C2({ S25607 }),
  .ZN({ S4654 })
);
NAND2_X1 #() 
NAND2_X1_5574_ (
  .A1({ S4627 }),
  .A2({ S4629 }),
  .ZN({ S4655 })
);
NAND4_X1 #() 
NAND4_X1_661_ (
  .A1({ S4330 }),
  .A2({ S4476 }),
  .A3({ S4248 }),
  .A4({ S2524 }),
  .ZN({ S4656 })
);
AOI21_X1 #() 
AOI21_X1_3171_ (
  .A({ S25673 }),
  .B1({ S4655 }),
  .B2({ S4656 }),
  .ZN({ S4657 })
);
INV_X1 #() 
INV_X1_1806_ (
  .A({ S4632 }),
  .ZN({ S4658 })
);
OAI21_X1 #() 
OAI21_X1_2894_ (
  .A({ S25957[790] }),
  .B1({ S4657 }),
  .B2({ S4658 }),
  .ZN({ S4659 })
);
NAND2_X1 #() 
NAND2_X1_5575_ (
  .A1({ S4303 }),
  .A2({ S4634 }),
  .ZN({ S4660 })
);
NAND2_X1 #() 
NAND2_X1_5576_ (
  .A1({ S4635 }),
  .A2({ S25957[788] }),
  .ZN({ S4661 })
);
AOI21_X1 #() 
AOI21_X1_3172_ (
  .A({ S25673 }),
  .B1({ S4660 }),
  .B2({ S4661 }),
  .ZN({ S4662 })
);
AOI21_X1 #() 
AOI21_X1_3173_ (
  .A({ S98 }),
  .B1({ S4329 }),
  .B2({ S4178 }),
  .ZN({ S4663 })
);
OAI21_X1 #() 
OAI21_X1_2895_ (
  .A({ S25957[788] }),
  .B1({ S4663 }),
  .B2({ S4637 }),
  .ZN({ S4664 })
);
AOI21_X1 #() 
AOI21_X1_3174_ (
  .A({ S25957[787] }),
  .B1({ S4171 }),
  .B2({ S4192 }),
  .ZN({ S4665 })
);
INV_X1 #() 
INV_X1_1807_ (
  .A({ S4640 }),
  .ZN({ S4666 })
);
OAI21_X1 #() 
OAI21_X1_2896_ (
  .A({ S2524 }),
  .B1({ S4666 }),
  .B2({ S4665 }),
  .ZN({ S4667 })
);
AOI21_X1 #() 
AOI21_X1_3175_ (
  .A({ S25957[789] }),
  .B1({ S4664 }),
  .B2({ S4667 }),
  .ZN({ S4668 })
);
OAI21_X1 #() 
OAI21_X1_2897_ (
  .A({ S25607 }),
  .B1({ S4668 }),
  .B2({ S4662 }),
  .ZN({ S4669 })
);
NAND3_X1 #() 
NAND3_X1_6055_ (
  .A1({ S4669 }),
  .A2({ S2361 }),
  .A3({ S4659 }),
  .ZN({ S4670 })
);
NAND3_X1 #() 
NAND3_X1_6056_ (
  .A1({ S4670 }),
  .A2({ S25957[888] }),
  .A3({ S4654 }),
  .ZN({ S4671 })
);
AOI21_X1 #() 
AOI21_X1_3176_ (
  .A({ S4597 }),
  .B1({ S4671 }),
  .B2({ S4645 }),
  .ZN({ S4672 })
);
INV_X1 #() 
INV_X1_1808_ (
  .A({ S4597 }),
  .ZN({ S25957[952] })
);
NAND3_X1 #() 
NAND3_X1_6057_ (
  .A1({ S4626 }),
  .A2({ S25957[888] }),
  .A3({ S4644 }),
  .ZN({ S4673 })
);
NAND3_X1 #() 
NAND3_X1_6058_ (
  .A1({ S4670 }),
  .A2({ S4600 }),
  .A3({ S4654 }),
  .ZN({ S4674 })
);
AOI21_X1 #() 
AOI21_X1_3177_ (
  .A({ S25957[952] }),
  .B1({ S4674 }),
  .B2({ S4673 }),
  .ZN({ S4675 })
);
OAI21_X1 #() 
OAI21_X1_2898_ (
  .A({ S25957[792] }),
  .B1({ S4672 }),
  .B2({ S4675 }),
  .ZN({ S4676 })
);
NAND3_X1 #() 
NAND3_X1_6059_ (
  .A1({ S4674 }),
  .A2({ S4673 }),
  .A3({ S25957[952] }),
  .ZN({ S4677 })
);
NAND3_X1 #() 
NAND3_X1_6060_ (
  .A1({ S4671 }),
  .A2({ S4645 }),
  .A3({ S4597 }),
  .ZN({ S4678 })
);
NAND3_X1 #() 
NAND3_X1_6061_ (
  .A1({ S4677 }),
  .A2({ S4678 }),
  .A3({ S3481 }),
  .ZN({ S4679 })
);
NAND2_X1 #() 
NAND2_X1_5577_ (
  .A1({ S4676 }),
  .A2({ S4679 }),
  .ZN({ S25957[664] })
);
NOR2_X1 #() 
NOR2_X1_1395_ (
  .A1({ S2136 }),
  .A2({ S2139 }),
  .ZN({ S25957[825] })
);
NAND2_X1 #() 
NAND2_X1_5578_ (
  .A1({ S2137 }),
  .A2({ S2138 }),
  .ZN({ S4680 })
);
INV_X1 #() 
INV_X1_1809_ (
  .A({ S4680 }),
  .ZN({ S25957[857] })
);
NAND2_X1 #() 
NAND2_X1_5579_ (
  .A1({ S2131 }),
  .A2({ S2111 }),
  .ZN({ S25957[889] })
);
INV_X1 #() 
INV_X1_1810_ (
  .A({ S25957[889] }),
  .ZN({ S4681 })
);
OAI211_X1 #() 
OAI211_X1_1979_ (
  .A({ S4519 }),
  .B({ S25957[788] }),
  .C1({ S4289 }),
  .C2({ S4412 }),
  .ZN({ S4682 })
);
NAND3_X1 #() 
NAND3_X1_6062_ (
  .A1({ S4627 }),
  .A2({ S2524 }),
  .A3({ S4385 }),
  .ZN({ S4683 })
);
NAND3_X1 #() 
NAND3_X1_6063_ (
  .A1({ S4683 }),
  .A2({ S25957[789] }),
  .A3({ S4682 }),
  .ZN({ S4684 })
);
AOI21_X1 #() 
AOI21_X1_3178_ (
  .A({ S25957[784] }),
  .B1({ S25957[785] }),
  .B2({ S25957[786] }),
  .ZN({ S4685 })
);
AOI21_X1 #() 
AOI21_X1_3179_ (
  .A({ S2524 }),
  .B1({ S4685 }),
  .B2({ S98 }),
  .ZN({ S4686 })
);
NAND2_X1 #() 
NAND2_X1_5580_ (
  .A1({ S4394 }),
  .A2({ S4686 }),
  .ZN({ S4687 })
);
NAND4_X1 #() 
NAND4_X1_662_ (
  .A1({ S4228 }),
  .A2({ S4218 }),
  .A3({ S4166 }),
  .A4({ S98 }),
  .ZN({ S4688 })
);
AOI21_X1 #() 
AOI21_X1_3180_ (
  .A({ S25957[788] }),
  .B1({ S4172 }),
  .B2({ S4166 }),
  .ZN({ S4689 })
);
AOI21_X1 #() 
AOI21_X1_3181_ (
  .A({ S25957[789] }),
  .B1({ S4689 }),
  .B2({ S4688 }),
  .ZN({ S4690 })
);
AOI21_X1 #() 
AOI21_X1_3182_ (
  .A({ S25607 }),
  .B1({ S4690 }),
  .B2({ S4687 }),
  .ZN({ S4691 })
);
NAND2_X1 #() 
NAND2_X1_5581_ (
  .A1({ S4691 }),
  .A2({ S4684 }),
  .ZN({ S4692 })
);
OAI21_X1 #() 
OAI21_X1_2899_ (
  .A({ S2524 }),
  .B1({ S4409 }),
  .B2({ S4357 }),
  .ZN({ S4693 })
);
NAND3_X1 #() 
NAND3_X1_6064_ (
  .A1({ S4249 }),
  .A2({ S98 }),
  .A3({ S4170 }),
  .ZN({ S4694 })
);
NAND4_X1 #() 
NAND4_X1_663_ (
  .A1({ S4299 }),
  .A2({ S4175 }),
  .A3({ S4694 }),
  .A4({ S25957[788] }),
  .ZN({ S4695 })
);
OAI211_X1 #() 
OAI211_X1_1980_ (
  .A({ S25673 }),
  .B({ S4695 }),
  .C1({ S4240 }),
  .C2({ S4693 }),
  .ZN({ S4696 })
);
NOR2_X1 #() 
NOR2_X1_1396_ (
  .A1({ S4179 }),
  .A2({ S4404 }),
  .ZN({ S4697 })
);
OAI21_X1 #() 
OAI21_X1_2900_ (
  .A({ S25957[788] }),
  .B1({ S4250 }),
  .B2({ S4248 }),
  .ZN({ S4698 })
);
NAND3_X1 #() 
NAND3_X1_6065_ (
  .A1({ S4213 }),
  .A2({ S25957[787] }),
  .A3({ S4180 }),
  .ZN({ S4699 })
);
NAND3_X1 #() 
NAND3_X1_6066_ (
  .A1({ S4552 }),
  .A2({ S4699 }),
  .A3({ S2524 }),
  .ZN({ S4700 })
);
OAI211_X1 #() 
OAI211_X1_1981_ (
  .A({ S25957[789] }),
  .B({ S4700 }),
  .C1({ S4697 }),
  .C2({ S4698 }),
  .ZN({ S4701 })
);
NAND3_X1 #() 
NAND3_X1_6067_ (
  .A1({ S4696 }),
  .A2({ S4701 }),
  .A3({ S25607 }),
  .ZN({ S4702 })
);
NAND3_X1 #() 
NAND3_X1_6068_ (
  .A1({ S4692 }),
  .A2({ S25957[791] }),
  .A3({ S4702 }),
  .ZN({ S4703 })
);
AOI21_X1 #() 
AOI21_X1_3183_ (
  .A({ S98 }),
  .B1({ S4203 }),
  .B2({ S4544 }),
  .ZN({ S4704 })
);
NAND3_X1 #() 
NAND3_X1_6069_ (
  .A1({ S4228 }),
  .A2({ S4399 }),
  .A3({ S98 }),
  .ZN({ S4705 })
);
NAND2_X1 #() 
NAND2_X1_5582_ (
  .A1({ S4705 }),
  .A2({ S25957[788] }),
  .ZN({ S4706 })
);
NAND3_X1 #() 
NAND3_X1_6070_ (
  .A1({ S4306 }),
  .A2({ S4619 }),
  .A3({ S2524 }),
  .ZN({ S4707 })
);
OAI211_X1 #() 
OAI211_X1_1982_ (
  .A({ S4707 }),
  .B({ S25673 }),
  .C1({ S4704 }),
  .C2({ S4706 }),
  .ZN({ S4708 })
);
OAI211_X1 #() 
OAI211_X1_1983_ (
  .A({ S4541 }),
  .B({ S25957[788] }),
  .C1({ S4207 }),
  .C2({ S4193 }),
  .ZN({ S4709 })
);
AND3_X1 #() 
AND3_X1_243_ (
  .A1({ S4223 }),
  .A2({ S2524 }),
  .A3({ S4218 }),
  .ZN({ S4710 })
);
AOI21_X1 #() 
AOI21_X1_3184_ (
  .A({ S25673 }),
  .B1({ S4710 }),
  .B2({ S4228 }),
  .ZN({ S4711 })
);
AOI21_X1 #() 
AOI21_X1_3185_ (
  .A({ S25607 }),
  .B1({ S4711 }),
  .B2({ S4709 }),
  .ZN({ S4712 })
);
NAND2_X1 #() 
NAND2_X1_5583_ (
  .A1({ S4712 }),
  .A2({ S4708 }),
  .ZN({ S4713 })
);
NAND4_X1 #() 
NAND4_X1_664_ (
  .A1({ S25957[787] }),
  .A2({ S4186 }),
  .A3({ S25957[785] }),
  .A4({ S4180 }),
  .ZN({ S4714 })
);
AOI21_X1 #() 
AOI21_X1_3186_ (
  .A({ S2524 }),
  .B1({ S4714 }),
  .B2({ S4466 }),
  .ZN({ S4715 })
);
OAI21_X1 #() 
OAI21_X1_2901_ (
  .A({ S25957[789] }),
  .B1({ S4237 }),
  .B2({ S4715 }),
  .ZN({ S4716 })
);
NAND2_X1 #() 
NAND2_X1_5584_ (
  .A1({ S4215 }),
  .A2({ S4321 }),
  .ZN({ S4717 })
);
NAND3_X1 #() 
NAND3_X1_6071_ (
  .A1({ S4225 }),
  .A2({ S4471 }),
  .A3({ S4222 }),
  .ZN({ S4718 })
);
NAND3_X1 #() 
NAND3_X1_6072_ (
  .A1({ S4717 }),
  .A2({ S4718 }),
  .A3({ S25673 }),
  .ZN({ S4719 })
);
NAND3_X1 #() 
NAND3_X1_6073_ (
  .A1({ S4716 }),
  .A2({ S4719 }),
  .A3({ S25607 }),
  .ZN({ S4720 })
);
NAND3_X1 #() 
NAND3_X1_6074_ (
  .A1({ S4720 }),
  .A2({ S4713 }),
  .A3({ S2361 }),
  .ZN({ S4721 })
);
NAND3_X1 #() 
NAND3_X1_6075_ (
  .A1({ S4703 }),
  .A2({ S4721 }),
  .A3({ S4681 }),
  .ZN({ S4722 })
);
NAND2_X1 #() 
NAND2_X1_5585_ (
  .A1({ S4703 }),
  .A2({ S4721 }),
  .ZN({ S4723 })
);
NAND2_X1 #() 
NAND2_X1_5586_ (
  .A1({ S4723 }),
  .A2({ S25957[889] }),
  .ZN({ S4724 })
);
NAND3_X1 #() 
NAND3_X1_6076_ (
  .A1({ S4724 }),
  .A2({ S25957[857] }),
  .A3({ S4722 }),
  .ZN({ S4725 })
);
NAND2_X1 #() 
NAND2_X1_5587_ (
  .A1({ S4723 }),
  .A2({ S4681 }),
  .ZN({ S4726 })
);
NAND3_X1 #() 
NAND3_X1_6077_ (
  .A1({ S4703 }),
  .A2({ S4721 }),
  .A3({ S25957[889] }),
  .ZN({ S4727 })
);
NAND3_X1 #() 
NAND3_X1_6078_ (
  .A1({ S4726 }),
  .A2({ S4680 }),
  .A3({ S4727 }),
  .ZN({ S4728 })
);
NAND3_X1 #() 
NAND3_X1_6079_ (
  .A1({ S4725 }),
  .A2({ S4728 }),
  .A3({ S25957[825] }),
  .ZN({ S4729 })
);
INV_X1 #() 
INV_X1_1811_ (
  .A({ S25957[825] }),
  .ZN({ S4730 })
);
NAND3_X1 #() 
NAND3_X1_6080_ (
  .A1({ S4726 }),
  .A2({ S25957[857] }),
  .A3({ S4727 }),
  .ZN({ S4731 })
);
NAND3_X1 #() 
NAND3_X1_6081_ (
  .A1({ S4724 }),
  .A2({ S4680 }),
  .A3({ S4722 }),
  .ZN({ S4732 })
);
NAND3_X1 #() 
NAND3_X1_6082_ (
  .A1({ S4731 }),
  .A2({ S4732 }),
  .A3({ S4730 }),
  .ZN({ S4733 })
);
NAND3_X1 #() 
NAND3_X1_6083_ (
  .A1({ S4729 }),
  .A2({ S4733 }),
  .A3({ S25957[793] }),
  .ZN({ S4734 })
);
NAND3_X1 #() 
NAND3_X1_6084_ (
  .A1({ S4731 }),
  .A2({ S4732 }),
  .A3({ S25957[825] }),
  .ZN({ S4735 })
);
NAND3_X1 #() 
NAND3_X1_6085_ (
  .A1({ S4725 }),
  .A2({ S4728 }),
  .A3({ S4730 }),
  .ZN({ S4736 })
);
NAND3_X1 #() 
NAND3_X1_6086_ (
  .A1({ S4735 }),
  .A2({ S4736 }),
  .A3({ S3527 }),
  .ZN({ S4737 })
);
NAND2_X1 #() 
NAND2_X1_5588_ (
  .A1({ S4734 }),
  .A2({ S4737 }),
  .ZN({ S25957[665] })
);
OAI211_X1 #() 
OAI211_X1_1984_ (
  .A({ S25957[787] }),
  .B({ S4177 }),
  .C1({ S4178 }),
  .C2({ S4170 }),
  .ZN({ S4738 })
);
AOI21_X1 #() 
AOI21_X1_3187_ (
  .A({ S25957[788] }),
  .B1({ S4738 }),
  .B2({ S4316 }),
  .ZN({ S4739 })
);
NAND3_X1 #() 
NAND3_X1_6087_ (
  .A1({ S4213 }),
  .A2({ S25957[787] }),
  .A3({ S25957[784] }),
  .ZN({ S4740 })
);
AOI21_X1 #() 
AOI21_X1_3188_ (
  .A({ S2524 }),
  .B1({ S4321 }),
  .B2({ S4740 }),
  .ZN({ S4741 })
);
OAI21_X1 #() 
OAI21_X1_2902_ (
  .A({ S25957[789] }),
  .B1({ S4739 }),
  .B2({ S4741 }),
  .ZN({ S4742 })
);
NAND2_X1 #() 
NAND2_X1_5589_ (
  .A1({ S4190 }),
  .A2({ S98 }),
  .ZN({ S4743 })
);
NAND3_X1 #() 
NAND3_X1_6088_ (
  .A1({ S25957[787] }),
  .A2({ S25957[785] }),
  .A3({ S4180 }),
  .ZN({ S4744 })
);
NAND3_X1 #() 
NAND3_X1_6089_ (
  .A1({ S4743 }),
  .A2({ S4744 }),
  .A3({ S25957[788] }),
  .ZN({ S4745 })
);
OAI211_X1 #() 
OAI211_X1_1985_ (
  .A({ S25673 }),
  .B({ S4745 }),
  .C1({ S4333 }),
  .C2({ S25957[788] }),
  .ZN({ S4746 })
);
NAND3_X1 #() 
NAND3_X1_6090_ (
  .A1({ S4742 }),
  .A2({ S25607 }),
  .A3({ S4746 }),
  .ZN({ S4747 })
);
AOI21_X1 #() 
AOI21_X1_3189_ (
  .A({ S4357 }),
  .B1({ S4170 }),
  .B2({ S4327 }),
  .ZN({ S4748 })
);
AOI21_X1 #() 
AOI21_X1_3190_ (
  .A({ S4185 }),
  .B1({ S4748 }),
  .B2({ S25957[787] }),
  .ZN({ S4749 })
);
AOI21_X1 #() 
AOI21_X1_3191_ (
  .A({ S25957[787] }),
  .B1({ S4171 }),
  .B2({ S4211 }),
  .ZN({ S4750 })
);
OAI21_X1 #() 
OAI21_X1_2903_ (
  .A({ S25957[788] }),
  .B1({ S4234 }),
  .B2({ S4235 }),
  .ZN({ S4751 })
);
OAI21_X1 #() 
OAI21_X1_2904_ (
  .A({ S25957[789] }),
  .B1({ S4751 }),
  .B2({ S4750 }),
  .ZN({ S4752 })
);
AND3_X1 #() 
AND3_X1_244_ (
  .A1({ S4172 }),
  .A2({ S4211 }),
  .A3({ S4171 }),
  .ZN({ S4753 })
);
NAND3_X1 #() 
NAND3_X1_6091_ (
  .A1({ S4264 }),
  .A2({ S2524 }),
  .A3({ S4694 }),
  .ZN({ S4754 })
);
OAI211_X1 #() 
OAI211_X1_1986_ (
  .A({ S25673 }),
  .B({ S4754 }),
  .C1({ S4753 }),
  .C2({ S4364 }),
  .ZN({ S4755 })
);
OAI211_X1 #() 
OAI211_X1_1987_ (
  .A({ S4755 }),
  .B({ S25957[790] }),
  .C1({ S4749 }),
  .C2({ S4752 }),
  .ZN({ S4756 })
);
NAND3_X1 #() 
NAND3_X1_6092_ (
  .A1({ S4756 }),
  .A2({ S4747 }),
  .A3({ S25957[791] }),
  .ZN({ S4757 })
);
NAND3_X1 #() 
NAND3_X1_6093_ (
  .A1({ S4213 }),
  .A2({ S4178 }),
  .A3({ S25957[787] }),
  .ZN({ S4758 })
);
NAND2_X1 #() 
NAND2_X1_5590_ (
  .A1({ S4758 }),
  .A2({ S4555 }),
  .ZN({ S4759 })
);
NAND2_X1 #() 
NAND2_X1_5591_ (
  .A1({ S4759 }),
  .A2({ S25957[788] }),
  .ZN({ S4760 })
);
OAI21_X1 #() 
OAI21_X1_2905_ (
  .A({ S2524 }),
  .B1({ S4743 }),
  .B2({ S2749 }),
  .ZN({ S4761 })
);
OAI211_X1 #() 
OAI211_X1_1988_ (
  .A({ S4760 }),
  .B({ S25957[789] }),
  .C1({ S4205 }),
  .C2({ S4761 }),
  .ZN({ S4762 })
);
NAND4_X1 #() 
NAND4_X1_665_ (
  .A1({ S4213 }),
  .A2({ S25957[787] }),
  .A3({ S4180 }),
  .A4({ S4186 }),
  .ZN({ S4763 })
);
OAI21_X1 #() 
OAI21_X1_2906_ (
  .A({ S4259 }),
  .B1({ S4289 }),
  .B2({ S4234 }),
  .ZN({ S4764 })
);
NAND3_X1 #() 
NAND3_X1_6094_ (
  .A1({ S4764 }),
  .A2({ S25957[788] }),
  .A3({ S4763 }),
  .ZN({ S4765 })
);
NAND3_X1 #() 
NAND3_X1_6095_ (
  .A1({ S4480 }),
  .A2({ S2524 }),
  .A3({ S4744 }),
  .ZN({ S4766 })
);
NAND3_X1 #() 
NAND3_X1_6096_ (
  .A1({ S4765 }),
  .A2({ S25673 }),
  .A3({ S4766 }),
  .ZN({ S4767 })
);
NAND3_X1 #() 
NAND3_X1_6097_ (
  .A1({ S4767 }),
  .A2({ S4762 }),
  .A3({ S25957[790] }),
  .ZN({ S4768 })
);
NOR2_X1 #() 
NOR2_X1_1397_ (
  .A1({ S4179 }),
  .A2({ S4300 }),
  .ZN({ S4769 })
);
NOR2_X1 #() 
NOR2_X1_1398_ (
  .A1({ S25957[785] }),
  .A2({ S4174 }),
  .ZN({ S4770 })
);
OAI21_X1 #() 
OAI21_X1_2907_ (
  .A({ S25957[788] }),
  .B1({ S4770 }),
  .B2({ S4235 }),
  .ZN({ S4771 })
);
AOI21_X1 #() 
AOI21_X1_3192_ (
  .A({ S98 }),
  .B1({ S4239 }),
  .B2({ S4544 }),
  .ZN({ S4772 })
);
OAI21_X1 #() 
OAI21_X1_2908_ (
  .A({ S2524 }),
  .B1({ S4219 }),
  .B2({ S4174 }),
  .ZN({ S4773 })
);
OAI22_X1 #() 
OAI22_X1_146_ (
  .A1({ S4769 }),
  .A2({ S4771 }),
  .B1({ S4772 }),
  .B2({ S4773 }),
  .ZN({ S4774 })
);
NAND2_X1 #() 
NAND2_X1_5592_ (
  .A1({ S4774 }),
  .A2({ S25957[789] }),
  .ZN({ S4775 })
);
OAI21_X1 #() 
OAI21_X1_2909_ (
  .A({ S4744 }),
  .B1({ S4267 }),
  .B2({ S4250 }),
  .ZN({ S4776 })
);
NAND2_X1 #() 
NAND2_X1_5593_ (
  .A1({ S4776 }),
  .A2({ S25957[788] }),
  .ZN({ S4777 })
);
NAND4_X1 #() 
NAND4_X1_666_ (
  .A1({ S4293 }),
  .A2({ S4180 }),
  .A3({ S4213 }),
  .A4({ S25957[787] }),
  .ZN({ S4778 })
);
NAND3_X1 #() 
NAND3_X1_6098_ (
  .A1({ S4606 }),
  .A2({ S2524 }),
  .A3({ S4778 }),
  .ZN({ S4779 })
);
NAND3_X1 #() 
NAND3_X1_6099_ (
  .A1({ S4779 }),
  .A2({ S4777 }),
  .A3({ S25673 }),
  .ZN({ S4780 })
);
NAND3_X1 #() 
NAND3_X1_6100_ (
  .A1({ S4775 }),
  .A2({ S25607 }),
  .A3({ S4780 }),
  .ZN({ S4781 })
);
NAND2_X1 #() 
NAND2_X1_5594_ (
  .A1({ S4781 }),
  .A2({ S4768 }),
  .ZN({ S4782 })
);
NAND2_X1 #() 
NAND2_X1_5595_ (
  .A1({ S4782 }),
  .A2({ S2361 }),
  .ZN({ S4783 })
);
AOI21_X1 #() 
AOI21_X1_3193_ (
  .A({ S2145 }),
  .B1({ S4783 }),
  .B2({ S4757 }),
  .ZN({ S4784 })
);
AND3_X1 #() 
AND3_X1_245_ (
  .A1({ S4756 }),
  .A2({ S4747 }),
  .A3({ S25957[791] }),
  .ZN({ S4785 })
);
AOI21_X1 #() 
AOI21_X1_3194_ (
  .A({ S25957[791] }),
  .B1({ S4781 }),
  .B2({ S4768 }),
  .ZN({ S4786 })
);
NOR3_X1 #() 
NOR3_X1_177_ (
  .A1({ S4786 }),
  .A2({ S4785 }),
  .A3({ S25957[986] }),
  .ZN({ S4787 })
);
OAI21_X1 #() 
OAI21_X1_2910_ (
  .A({ S1033 }),
  .B1({ S4784 }),
  .B2({ S4787 }),
  .ZN({ S4788 })
);
OAI21_X1 #() 
OAI21_X1_2911_ (
  .A({ S25957[986] }),
  .B1({ S4786 }),
  .B2({ S4785 }),
  .ZN({ S4789 })
);
NAND3_X1 #() 
NAND3_X1_6101_ (
  .A1({ S4783 }),
  .A2({ S2145 }),
  .A3({ S4757 }),
  .ZN({ S4790 })
);
NAND3_X1 #() 
NAND3_X1_6102_ (
  .A1({ S4790 }),
  .A2({ S25957[922] }),
  .A3({ S4789 }),
  .ZN({ S4791 })
);
NAND2_X1 #() 
NAND2_X1_5596_ (
  .A1({ S4788 }),
  .A2({ S4791 }),
  .ZN({ S25957[666] })
);
AOI21_X1 #() 
AOI21_X1_3195_ (
  .A({ S25957[776] }),
  .B1({ S3352 }),
  .B2({ S3353 }),
  .ZN({ S4792 })
);
AND3_X1 #() 
AND3_X1_246_ (
  .A1({ S3353 }),
  .A2({ S3352 }),
  .A3({ S25957[776] }),
  .ZN({ S4793 })
);
NOR2_X1 #() 
NOR2_X1_1399_ (
  .A1({ S4793 }),
  .A2({ S4792 }),
  .ZN({ S4794 })
);
AOI21_X1 #() 
AOI21_X1_3196_ (
  .A({ S4794 }),
  .B1({ S3407 }),
  .B2({ S3410 }),
  .ZN({ S4 })
);
NAND3_X1 #() 
NAND3_X1_6103_ (
  .A1({ S3407 }),
  .A2({ S3410 }),
  .A3({ S4794 }),
  .ZN({ S5 })
);
NAND3_X1 #() 
NAND3_X1_6104_ (
  .A1({ S2358 }),
  .A2({ S2359 }),
  .A3({ S2361 }),
  .ZN({ S4795 })
);
NAND2_X1 #() 
NAND2_X1_5597_ (
  .A1({ S25957[695] }),
  .A2({ S25957[791] }),
  .ZN({ S4796 })
);
NAND2_X1 #() 
NAND2_X1_5598_ (
  .A1({ S4796 }),
  .A2({ S4795 }),
  .ZN({ S4797 })
);
NAND2_X1 #() 
NAND2_X1_5599_ (
  .A1({ S3147 }),
  .A2({ S3152 }),
  .ZN({ S4798 })
);
NAND2_X1 #() 
NAND2_X1_5600_ (
  .A1({ S25957[650] }),
  .A2({ S25957[648] }),
  .ZN({ S4799 })
);
NAND2_X1 #() 
NAND2_X1_5601_ (
  .A1({ S25957[649] }),
  .A2({ S113 }),
  .ZN({ S4800 })
);
INV_X1 #() 
INV_X1_1812_ (
  .A({ S4800 }),
  .ZN({ S4801 })
);
NAND2_X1 #() 
NAND2_X1_5602_ (
  .A1({ S4801 }),
  .A2({ S4799 }),
  .ZN({ S4802 })
);
INV_X1 #() 
INV_X1_1813_ (
  .A({ S25957[652] }),
  .ZN({ S4803 })
);
AOI21_X1 #() 
AOI21_X1_3197_ (
  .A({ S113 }),
  .B1({ S25957[649] }),
  .B2({ S4799 }),
  .ZN({ S4804 })
);
NOR2_X1 #() 
NOR2_X1_1400_ (
  .A1({ S4804 }),
  .A2({ S4803 }),
  .ZN({ S4805 })
);
AND2_X1 #() 
AND2_X1_353_ (
  .A1({ S3410 }),
  .A2({ S3407 }),
  .ZN({ S4806 })
);
NOR2_X1 #() 
NOR2_X1_1401_ (
  .A1({ S25957[650] }),
  .A2({ S25957[648] }),
  .ZN({ S4807 })
);
NAND2_X1 #() 
NAND2_X1_5603_ (
  .A1({ S4806 }),
  .A2({ S4807 }),
  .ZN({ S4808 })
);
AOI211_X1 #() 
AOI211_X1_95_ (
  .A({ S4 }),
  .B({ S25957[652] }),
  .C1({ S4808 }),
  .C2({ S113 }),
  .ZN({ S4809 })
);
AOI211_X1 #() 
AOI211_X1_96_ (
  .A({ S4798 }),
  .B({ S4809 }),
  .C1({ S4802 }),
  .C2({ S4805 }),
  .ZN({ S4810 })
);
NAND3_X1 #() 
NAND3_X1_6105_ (
  .A1({ S3407 }),
  .A2({ S3410 }),
  .A3({ S25957[648] }),
  .ZN({ S4811 })
);
NAND4_X1 #() 
NAND4_X1_667_ (
  .A1({ S3407 }),
  .A2({ S3410 }),
  .A3({ S3477 }),
  .A4({ S3480 }),
  .ZN({ S4812 })
);
NAND3_X1 #() 
NAND3_X1_6106_ (
  .A1({ S4794 }),
  .A2({ S3477 }),
  .A3({ S3480 }),
  .ZN({ S4813 })
);
NAND2_X1 #() 
NAND2_X1_5604_ (
  .A1({ S4812 }),
  .A2({ S4813 }),
  .ZN({ S4814 })
);
AOI22_X1 #() 
AOI22_X1_635_ (
  .A1({ S4814 }),
  .A2({ S5 }),
  .B1({ S25957[650] }),
  .B2({ S4811 }),
  .ZN({ S4815 })
);
AND2_X1 #() 
AND2_X1_354_ (
  .A1({ S3480 }),
  .A2({ S3477 }),
  .ZN({ S4816 })
);
AOI21_X1 #() 
AOI21_X1_3198_ (
  .A({ S113 }),
  .B1({ S4806 }),
  .B2({ S4816 }),
  .ZN({ S4817 })
);
NOR2_X1 #() 
NOR2_X1_1402_ (
  .A1({ S4817 }),
  .A2({ S25957[652] }),
  .ZN({ S4818 })
);
OAI21_X1 #() 
OAI21_X1_2912_ (
  .A({ S4818 }),
  .B1({ S4815 }),
  .B2({ S25957[651] }),
  .ZN({ S4819 })
);
INV_X1 #() 
INV_X1_1814_ (
  .A({ S4819 }),
  .ZN({ S4820 })
);
AOI21_X1 #() 
AOI21_X1_3199_ (
  .A({ S2258 }),
  .B1({ S3408 }),
  .B2({ S3409 }),
  .ZN({ S4821 })
);
AOI21_X1 #() 
AOI21_X1_3200_ (
  .A({ S25957[777] }),
  .B1({ S3406 }),
  .B2({ S3403 }),
  .ZN({ S4822 })
);
OAI21_X1 #() 
OAI21_X1_2913_ (
  .A({ S25957[650] }),
  .B1({ S4821 }),
  .B2({ S4822 }),
  .ZN({ S4823 })
);
AOI21_X1 #() 
AOI21_X1_3201_ (
  .A({ S25957[651] }),
  .B1({ S4816 }),
  .B2({ S25957[648] }),
  .ZN({ S4824 })
);
OAI21_X1 #() 
OAI21_X1_2914_ (
  .A({ S25957[648] }),
  .B1({ S4821 }),
  .B2({ S4822 }),
  .ZN({ S4825 })
);
NAND3_X1 #() 
NAND3_X1_6107_ (
  .A1({ S4825 }),
  .A2({ S4816 }),
  .A3({ S5 }),
  .ZN({ S4826 })
);
NAND3_X1 #() 
NAND3_X1_6108_ (
  .A1({ S25957[650] }),
  .A2({ S3407 }),
  .A3({ S3410 }),
  .ZN({ S4827 })
);
NAND2_X1 #() 
NAND2_X1_5605_ (
  .A1({ S4827 }),
  .A2({ S4799 }),
  .ZN({ S4828 })
);
AOI21_X1 #() 
AOI21_X1_3202_ (
  .A({ S113 }),
  .B1({ S4828 }),
  .B2({ S4811 }),
  .ZN({ S4829 })
);
AOI22_X1 #() 
AOI22_X1_636_ (
  .A1({ S4829 }),
  .A2({ S4826 }),
  .B1({ S4824 }),
  .B2({ S4823 }),
  .ZN({ S4830 })
);
AOI211_X1 #() 
AOI211_X1_97_ (
  .A({ S25957[653] }),
  .B({ S4820 }),
  .C1({ S25957[652] }),
  .C2({ S4830 }),
  .ZN({ S4831 })
);
OR2_X1 #() 
OR2_X1_72_ (
  .A1({ S4831 }),
  .A2({ S4810 }),
  .ZN({ S4832 })
);
AOI21_X1 #() 
AOI21_X1_3203_ (
  .A({ S25957[648] }),
  .B1({ S3407 }),
  .B2({ S3410 }),
  .ZN({ S4833 })
);
AOI21_X1 #() 
AOI21_X1_3204_ (
  .A({ S113 }),
  .B1({ S25957[649] }),
  .B2({ S25957[648] }),
  .ZN({ S4834 })
);
NAND2_X1 #() 
NAND2_X1_5606_ (
  .A1({ S4834 }),
  .A2({ S4827 }),
  .ZN({ S4835 })
);
OAI21_X1 #() 
OAI21_X1_2915_ (
  .A({ S4835 }),
  .B1({ S25957[651] }),
  .B2({ S4833 }),
  .ZN({ S4836 })
);
NOR2_X1 #() 
NOR2_X1_1403_ (
  .A1({ S25957[649] }),
  .A2({ S113 }),
  .ZN({ S4837 })
);
NAND2_X1 #() 
NAND2_X1_5607_ (
  .A1({ S4837 }),
  .A2({ S25957[648] }),
  .ZN({ S4838 })
);
NAND4_X1 #() 
NAND4_X1_668_ (
  .A1({ S4838 }),
  .A2({ S4823 }),
  .A3({ S4799 }),
  .A4({ S4808 }),
  .ZN({ S4839 })
);
NAND2_X1 #() 
NAND2_X1_5608_ (
  .A1({ S4839 }),
  .A2({ S4803 }),
  .ZN({ S4840 })
);
OAI211_X1 #() 
OAI211_X1_1989_ (
  .A({ S4840 }),
  .B({ S4798 }),
  .C1({ S4803 }),
  .C2({ S4836 }),
  .ZN({ S4841 })
);
NAND2_X1 #() 
NAND2_X1_5609_ (
  .A1({ S4811 }),
  .A2({ S4816 }),
  .ZN({ S4842 })
);
NOR2_X1 #() 
NOR2_X1_1404_ (
  .A1({ S4842 }),
  .A2({ S113 }),
  .ZN({ S4843 })
);
AOI21_X1 #() 
AOI21_X1_3205_ (
  .A({ S25957[651] }),
  .B1({ S4816 }),
  .B2({ S4794 }),
  .ZN({ S4844 })
);
INV_X1 #() 
INV_X1_1815_ (
  .A({ S4844 }),
  .ZN({ S4845 })
);
AOI21_X1 #() 
AOI21_X1_3206_ (
  .A({ S113 }),
  .B1({ S3477 }),
  .B2({ S3480 }),
  .ZN({ S4846 })
);
NAND2_X1 #() 
NAND2_X1_5610_ (
  .A1({ S4846 }),
  .A2({ S25957[648] }),
  .ZN({ S4847 })
);
OAI21_X1 #() 
OAI21_X1_2916_ (
  .A({ S4847 }),
  .B1({ S4845 }),
  .B2({ S4806 }),
  .ZN({ S4848 })
);
NOR3_X1 #() 
NOR3_X1_178_ (
  .A1({ S4848 }),
  .A2({ S4843 }),
  .A3({ S4803 }),
  .ZN({ S4849 })
);
NAND4_X1 #() 
NAND4_X1_669_ (
  .A1({ S25957[650] }),
  .A2({ S3410 }),
  .A3({ S3407 }),
  .A4({ S4794 }),
  .ZN({ S4850 })
);
OAI211_X1 #() 
OAI211_X1_1990_ (
  .A({ S3477 }),
  .B({ S3480 }),
  .C1({ S4793 }),
  .C2({ S4792 }),
  .ZN({ S4851 })
);
INV_X1 #() 
INV_X1_1816_ (
  .A({ S4851 }),
  .ZN({ S4852 })
);
NAND2_X1 #() 
NAND2_X1_5611_ (
  .A1({ S4852 }),
  .A2({ S25957[649] }),
  .ZN({ S4853 })
);
NAND2_X1 #() 
NAND2_X1_5612_ (
  .A1({ S4853 }),
  .A2({ S4850 }),
  .ZN({ S4854 })
);
NAND2_X1 #() 
NAND2_X1_5613_ (
  .A1({ S4803 }),
  .A2({ S113 }),
  .ZN({ S4855 })
);
OAI211_X1 #() 
OAI211_X1_1991_ (
  .A({ S4794 }),
  .B({ S25957[650] }),
  .C1({ S4821 }),
  .C2({ S4822 }),
  .ZN({ S4856 })
);
NOR2_X1 #() 
NOR2_X1_1405_ (
  .A1({ S25957[652] }),
  .A2({ S113 }),
  .ZN({ S4857 })
);
NAND3_X1 #() 
NAND3_X1_6109_ (
  .A1({ S4856 }),
  .A2({ S4857 }),
  .A3({ S4811 }),
  .ZN({ S4858 })
);
OAI211_X1 #() 
OAI211_X1_1992_ (
  .A({ S4858 }),
  .B({ S25957[653] }),
  .C1({ S4854 }),
  .C2({ S4855 }),
  .ZN({ S4859 })
);
OAI211_X1 #() 
OAI211_X1_1993_ (
  .A({ S4841 }),
  .B({ S25957[654] }),
  .C1({ S4849 }),
  .C2({ S4859 }),
  .ZN({ S4860 })
);
OAI211_X1 #() 
OAI211_X1_1994_ (
  .A({ S25957[655] }),
  .B({ S4860 }),
  .C1({ S4832 }),
  .C2({ S25957[654] }),
  .ZN({ S4861 })
);
INV_X1 #() 
INV_X1_1817_ (
  .A({ S25957[654] }),
  .ZN({ S4862 })
);
AOI21_X1 #() 
AOI21_X1_3207_ (
  .A({ S25957[650] }),
  .B1({ S3410 }),
  .B2({ S3407 }),
  .ZN({ S4863 })
);
AOI21_X1 #() 
AOI21_X1_3208_ (
  .A({ S113 }),
  .B1({ S25957[650] }),
  .B2({ S25957[648] }),
  .ZN({ S4864 })
);
INV_X1 #() 
INV_X1_1818_ (
  .A({ S4864 }),
  .ZN({ S4865 })
);
NOR2_X1 #() 
NOR2_X1_1406_ (
  .A1({ S4865 }),
  .A2({ S4863 }),
  .ZN({ S4866 })
);
NOR2_X1 #() 
NOR2_X1_1407_ (
  .A1({ S4806 }),
  .A2({ S4799 }),
  .ZN({ S4867 })
);
OAI21_X1 #() 
OAI21_X1_2917_ (
  .A({ S113 }),
  .B1({ S25957[649] }),
  .B2({ S4851 }),
  .ZN({ S4868 })
);
OAI21_X1 #() 
OAI21_X1_2918_ (
  .A({ S4803 }),
  .B1({ S4867 }),
  .B2({ S4868 }),
  .ZN({ S4869 })
);
AOI21_X1 #() 
AOI21_X1_3209_ (
  .A({ S4816 }),
  .B1({ S4825 }),
  .B2({ S5 }),
  .ZN({ S4870 })
);
OAI21_X1 #() 
OAI21_X1_2919_ (
  .A({ S113 }),
  .B1({ S4870 }),
  .B2({ S4807 }),
  .ZN({ S4871 })
);
NAND2_X1 #() 
NAND2_X1_5614_ (
  .A1({ S4825 }),
  .A2({ S25957[650] }),
  .ZN({ S4872 })
);
OAI21_X1 #() 
OAI21_X1_2920_ (
  .A({ S4794 }),
  .B1({ S4821 }),
  .B2({ S4822 }),
  .ZN({ S4873 })
);
NAND3_X1 #() 
NAND3_X1_6110_ (
  .A1({ S4873 }),
  .A2({ S4816 }),
  .A3({ S4811 }),
  .ZN({ S4874 })
);
AOI21_X1 #() 
AOI21_X1_3210_ (
  .A({ S113 }),
  .B1({ S4874 }),
  .B2({ S4872 }),
  .ZN({ S4875 })
);
INV_X1 #() 
INV_X1_1819_ (
  .A({ S4875 }),
  .ZN({ S4876 })
);
NAND3_X1 #() 
NAND3_X1_6111_ (
  .A1({ S4876 }),
  .A2({ S25957[652] }),
  .A3({ S4871 }),
  .ZN({ S4877 })
);
OAI21_X1 #() 
OAI21_X1_2921_ (
  .A({ S4877 }),
  .B1({ S4866 }),
  .B2({ S4869 }),
  .ZN({ S4878 })
);
INV_X1 #() 
INV_X1_1820_ (
  .A({ S4878 }),
  .ZN({ S4879 })
);
NOR2_X1 #() 
NOR2_X1_1408_ (
  .A1({ S4854 }),
  .A2({ S113 }),
  .ZN({ S4880 })
);
INV_X1 #() 
INV_X1_1821_ (
  .A({ S4856 }),
  .ZN({ S4881 })
);
OAI21_X1 #() 
OAI21_X1_2922_ (
  .A({ S25957[652] }),
  .B1({ S4881 }),
  .B2({ S4845 }),
  .ZN({ S4882 })
);
NAND2_X1 #() 
NAND2_X1_5615_ (
  .A1({ S4806 }),
  .A2({ S4852 }),
  .ZN({ S4883 })
);
NAND2_X1 #() 
NAND2_X1_5616_ (
  .A1({ S4883 }),
  .A2({ S4823 }),
  .ZN({ S4884 })
);
NAND2_X1 #() 
NAND2_X1_5617_ (
  .A1({ S4884 }),
  .A2({ S25957[651] }),
  .ZN({ S4885 })
);
INV_X1 #() 
INV_X1_1822_ (
  .A({ S4885 }),
  .ZN({ S4886 })
);
NAND2_X1 #() 
NAND2_X1_5618_ (
  .A1({ S25957[650] }),
  .A2({ S4794 }),
  .ZN({ S4887 })
);
NAND2_X1 #() 
NAND2_X1_5619_ (
  .A1({ S4827 }),
  .A2({ S4887 }),
  .ZN({ S4888 })
);
OAI21_X1 #() 
OAI21_X1_2923_ (
  .A({ S4803 }),
  .B1({ S4888 }),
  .B2({ S25957[651] }),
  .ZN({ S4889 })
);
OAI221_X1 #() 
OAI221_X1_167_ (
  .A({ S25957[653] }),
  .B1({ S4880 }),
  .B2({ S4882 }),
  .C1({ S4886 }),
  .C2({ S4889 }),
  .ZN({ S4890 })
);
OAI21_X1 #() 
OAI21_X1_2924_ (
  .A({ S4890 }),
  .B1({ S4879 }),
  .B2({ S25957[653] }),
  .ZN({ S4891 })
);
NAND2_X1 #() 
NAND2_X1_5620_ (
  .A1({ S4888 }),
  .A2({ S5 }),
  .ZN({ S4892 })
);
AOI21_X1 #() 
AOI21_X1_3211_ (
  .A({ S25957[651] }),
  .B1({ S4852 }),
  .B2({ S25957[649] }),
  .ZN({ S4893 })
);
NAND2_X1 #() 
NAND2_X1_5621_ (
  .A1({ S4892 }),
  .A2({ S4893 }),
  .ZN({ S4894 })
);
OAI21_X1 #() 
OAI21_X1_2925_ (
  .A({ S4894 }),
  .B1({ S113 }),
  .B2({ S4881 }),
  .ZN({ S4895 })
);
NAND2_X1 #() 
NAND2_X1_5622_ (
  .A1({ S4828 }),
  .A2({ S4811 }),
  .ZN({ S4896 })
);
NOR2_X1 #() 
NOR2_X1_1409_ (
  .A1({ S4896 }),
  .A2({ S25957[651] }),
  .ZN({ S4897 })
);
NAND2_X1 #() 
NAND2_X1_5623_ (
  .A1({ S25957[650] }),
  .A2({ S25957[651] }),
  .ZN({ S4898 })
);
NOR2_X1 #() 
NOR2_X1_1410_ (
  .A1({ S4 }),
  .A2({ S4898 }),
  .ZN({ S4899 })
);
OR3_X1 #() 
OR3_X1_37_ (
  .A1({ S4897 }),
  .A2({ S4899 }),
  .A3({ S25957[652] }),
  .ZN({ S4900 })
);
OAI21_X1 #() 
OAI21_X1_2926_ (
  .A({ S4900 }),
  .B1({ S4895 }),
  .B2({ S4803 }),
  .ZN({ S4901 })
);
NOR2_X1 #() 
NOR2_X1_1411_ (
  .A1({ S4794 }),
  .A2({ S25957[651] }),
  .ZN({ S4902 })
);
INV_X1 #() 
INV_X1_1823_ (
  .A({ S4812 }),
  .ZN({ S4903 })
);
NOR2_X1 #() 
NOR2_X1_1412_ (
  .A1({ S4903 }),
  .A2({ S4865 }),
  .ZN({ S4904 })
);
OAI21_X1 #() 
OAI21_X1_2927_ (
  .A({ S25957[652] }),
  .B1({ S4904 }),
  .B2({ S4902 }),
  .ZN({ S4905 })
);
NAND2_X1 #() 
NAND2_X1_5624_ (
  .A1({ S4823 }),
  .A2({ S113 }),
  .ZN({ S4906 })
);
NOR2_X1 #() 
NOR2_X1_1413_ (
  .A1({ S4906 }),
  .A2({ S4814 }),
  .ZN({ S4907 })
);
OAI21_X1 #() 
OAI21_X1_2928_ (
  .A({ S4816 }),
  .B1({ S4821 }),
  .B2({ S4822 }),
  .ZN({ S4908 })
);
NAND3_X1 #() 
NAND3_X1_6112_ (
  .A1({ S4908 }),
  .A2({ S25957[651] }),
  .A3({ S4811 }),
  .ZN({ S4909 })
);
NAND2_X1 #() 
NAND2_X1_5625_ (
  .A1({ S4909 }),
  .A2({ S4803 }),
  .ZN({ S4910 })
);
OAI21_X1 #() 
OAI21_X1_2929_ (
  .A({ S4905 }),
  .B1({ S4907 }),
  .B2({ S4910 }),
  .ZN({ S4911 })
);
AOI21_X1 #() 
AOI21_X1_3212_ (
  .A({ S25957[654] }),
  .B1({ S4911 }),
  .B2({ S25957[653] }),
  .ZN({ S4912 })
);
OAI21_X1 #() 
OAI21_X1_2930_ (
  .A({ S4912 }),
  .B1({ S25957[653] }),
  .B2({ S4901 }),
  .ZN({ S4913 })
);
OAI21_X1 #() 
OAI21_X1_2931_ (
  .A({ S4913 }),
  .B1({ S4891 }),
  .B2({ S4862 }),
  .ZN({ S4914 })
);
NAND2_X1 #() 
NAND2_X1_5626_ (
  .A1({ S4914 }),
  .A2({ S3020 }),
  .ZN({ S4915 })
);
NAND3_X1 #() 
NAND3_X1_6113_ (
  .A1({ S4861 }),
  .A2({ S4915 }),
  .A3({ S2356 }),
  .ZN({ S4916 })
);
NAND2_X1 #() 
NAND2_X1_5627_ (
  .A1({ S4861 }),
  .A2({ S4915 }),
  .ZN({ S4917 })
);
NAND2_X1 #() 
NAND2_X1_5628_ (
  .A1({ S4917 }),
  .A2({ S25957[759] }),
  .ZN({ S4918 })
);
NAND2_X1 #() 
NAND2_X1_5629_ (
  .A1({ S4918 }),
  .A2({ S4916 }),
  .ZN({ S25957[631] })
);
NOR2_X1 #() 
NOR2_X1_1414_ (
  .A1({ S25957[631] }),
  .A2({ S25957[823] }),
  .ZN({ S4919 })
);
INV_X1 #() 
INV_X1_1824_ (
  .A({ S25957[631] }),
  .ZN({ S4920 })
);
NOR2_X1 #() 
NOR2_X1_1415_ (
  .A1({ S4920 }),
  .A2({ S2238 }),
  .ZN({ S4921 })
);
OAI21_X1 #() 
OAI21_X1_2932_ (
  .A({ S4797 }),
  .B1({ S4921 }),
  .B2({ S4919 }),
  .ZN({ S4922 })
);
NOR2_X1 #() 
NOR2_X1_1416_ (
  .A1({ S4921 }),
  .A2({ S4919 }),
  .ZN({ S25957[567] })
);
NAND2_X1 #() 
NAND2_X1_5630_ (
  .A1({ S25957[567] }),
  .A2({ S25957[663] }),
  .ZN({ S4923 })
);
NAND2_X1 #() 
NAND2_X1_5631_ (
  .A1({ S4923 }),
  .A2({ S4922 }),
  .ZN({ S4924 })
);
INV_X1 #() 
INV_X1_1825_ (
  .A({ S4924 }),
  .ZN({ S25957[535] })
);
XNOR2_X1 #() 
XNOR2_X1_213_ (
  .A({ S25957[854] }),
  .B({ S2363 }),
  .ZN({ S25957[822] })
);
INV_X1 #() 
INV_X1_1826_ (
  .A({ S4869 }),
  .ZN({ S4925 })
);
AOI21_X1 #() 
AOI21_X1_3213_ (
  .A({ S25957[651] }),
  .B1({ S25957[650] }),
  .B2({ S4794 }),
  .ZN({ S4926 })
);
NAND2_X1 #() 
NAND2_X1_5632_ (
  .A1({ S4874 }),
  .A2({ S4926 }),
  .ZN({ S4927 })
);
NAND4_X1 #() 
NAND4_X1_670_ (
  .A1({ S25957[650] }),
  .A2({ S3410 }),
  .A3({ S3407 }),
  .A4({ S25957[648] }),
  .ZN({ S4928 })
);
NAND3_X1 #() 
NAND3_X1_6114_ (
  .A1({ S4928 }),
  .A2({ S25957[651] }),
  .A3({ S4813 }),
  .ZN({ S4929 })
);
AND2_X1 #() 
AND2_X1_355_ (
  .A1({ S4929 }),
  .A2({ S25957[652] }),
  .ZN({ S4930 })
);
INV_X1 #() 
INV_X1_1827_ (
  .A({ S5 }),
  .ZN({ S4931 })
);
NAND3_X1 #() 
NAND3_X1_6115_ (
  .A1({ S4812 }),
  .A2({ S25957[651] }),
  .A3({ S4813 }),
  .ZN({ S4932 })
);
OR2_X1 #() 
OR2_X1_73_ (
  .A1({ S4932 }),
  .A2({ S4931 }),
  .ZN({ S4933 })
);
AOI22_X1 #() 
AOI22_X1_637_ (
  .A1({ S4925 }),
  .A2({ S4933 }),
  .B1({ S4930 }),
  .B2({ S4927 }),
  .ZN({ S4934 })
);
NAND3_X1 #() 
NAND3_X1_6116_ (
  .A1({ S5 }),
  .A2({ S113 }),
  .A3({ S25957[650] }),
  .ZN({ S4935 })
);
NAND4_X1 #() 
NAND4_X1_671_ (
  .A1({ S4806 }),
  .A2({ S25957[651] }),
  .A3({ S4887 }),
  .A4({ S4851 }),
  .ZN({ S4936 })
);
AOI21_X1 #() 
AOI21_X1_3214_ (
  .A({ S4803 }),
  .B1({ S4935 }),
  .B2({ S4936 }),
  .ZN({ S4937 })
);
NOR2_X1 #() 
NOR2_X1_1417_ (
  .A1({ S4801 }),
  .A2({ S25957[652] }),
  .ZN({ S4938 })
);
AOI211_X1 #() 
AOI211_X1_98_ (
  .A({ S4798 }),
  .B({ S4937 }),
  .C1({ S4835 }),
  .C2({ S4938 }),
  .ZN({ S4939 })
);
AOI21_X1 #() 
AOI21_X1_3215_ (
  .A({ S4939 }),
  .B1({ S4934 }),
  .B2({ S4798 }),
  .ZN({ S4940 })
);
INV_X1 #() 
INV_X1_1828_ (
  .A({ S4897 }),
  .ZN({ S4941 })
);
OAI22_X1 #() 
OAI22_X1_147_ (
  .A1({ S4800 }),
  .A2({ S4813 }),
  .B1({ S4806 }),
  .B2({ S4898 }),
  .ZN({ S4942 })
);
INV_X1 #() 
INV_X1_1829_ (
  .A({ S4942 }),
  .ZN({ S4943 })
);
AOI21_X1 #() 
AOI21_X1_3216_ (
  .A({ S4803 }),
  .B1({ S4941 }),
  .B2({ S4943 }),
  .ZN({ S4944 })
);
NAND4_X1 #() 
NAND4_X1_672_ (
  .A1({ S4857 }),
  .A2({ S4823 }),
  .A3({ S4851 }),
  .A4({ S4812 }),
  .ZN({ S4945 })
);
NAND3_X1 #() 
NAND3_X1_6117_ (
  .A1({ S25957[649] }),
  .A2({ S25957[648] }),
  .A3({ S25957[650] }),
  .ZN({ S4946 })
);
NAND2_X1 #() 
NAND2_X1_5633_ (
  .A1({ S4946 }),
  .A2({ S5 }),
  .ZN({ S4947 })
);
OAI211_X1 #() 
OAI211_X1_1995_ (
  .A({ S4945 }),
  .B({ S25957[653] }),
  .C1({ S4947 }),
  .C2({ S4855 }),
  .ZN({ S4948 })
);
OAI21_X1 #() 
OAI21_X1_2933_ (
  .A({ S4805 }),
  .B1({ S25957[651] }),
  .B2({ S4842 }),
  .ZN({ S4949 })
);
NAND2_X1 #() 
NAND2_X1_5634_ (
  .A1({ S4856 }),
  .A2({ S4851 }),
  .ZN({ S4950 })
);
AOI22_X1 #() 
AOI22_X1_638_ (
  .A1({ S4950 }),
  .A2({ S25957[651] }),
  .B1({ S4874 }),
  .B2({ S4926 }),
  .ZN({ S4951 })
);
OAI21_X1 #() 
OAI21_X1_2934_ (
  .A({ S4949 }),
  .B1({ S4951 }),
  .B2({ S25957[652] }),
  .ZN({ S4952 })
);
OAI221_X1 #() 
OAI221_X1_168_ (
  .A({ S4862 }),
  .B1({ S4944 }),
  .B2({ S4948 }),
  .C1({ S4952 }),
  .C2({ S25957[653] }),
  .ZN({ S4953 })
);
OAI211_X1 #() 
OAI211_X1_1996_ (
  .A({ S4953 }),
  .B({ S25957[655] }),
  .C1({ S4940 }),
  .C2({ S4862 }),
  .ZN({ S4954 })
);
NAND2_X1 #() 
NAND2_X1_5635_ (
  .A1({ S4856 }),
  .A2({ S4928 }),
  .ZN({ S4955 })
);
NOR2_X1 #() 
NOR2_X1_1418_ (
  .A1({ S4955 }),
  .A2({ S25957[651] }),
  .ZN({ S4956 })
);
NAND2_X1 #() 
NAND2_X1_5636_ (
  .A1({ S4929 }),
  .A2({ S4803 }),
  .ZN({ S4957 })
);
NAND3_X1 #() 
NAND3_X1_6118_ (
  .A1({ S4812 }),
  .A2({ S113 }),
  .A3({ S4794 }),
  .ZN({ S4958 })
);
AOI21_X1 #() 
AOI21_X1_3217_ (
  .A({ S4803 }),
  .B1({ S4863 }),
  .B2({ S25957[651] }),
  .ZN({ S4959 })
);
AOI21_X1 #() 
AOI21_X1_3218_ (
  .A({ S25957[653] }),
  .B1({ S4959 }),
  .B2({ S4958 }),
  .ZN({ S4960 })
);
OAI21_X1 #() 
OAI21_X1_2935_ (
  .A({ S4960 }),
  .B1({ S4956 }),
  .B2({ S4957 }),
  .ZN({ S4961 })
);
NAND2_X1 #() 
NAND2_X1_5637_ (
  .A1({ S4873 }),
  .A2({ S4799 }),
  .ZN({ S4962 })
);
NAND2_X1 #() 
NAND2_X1_5638_ (
  .A1({ S4825 }),
  .A2({ S4813 }),
  .ZN({ S4963 })
);
AOI22_X1 #() 
AOI22_X1_639_ (
  .A1({ S4963 }),
  .A2({ S4824 }),
  .B1({ S4962 }),
  .B2({ S25957[651] }),
  .ZN({ S4964 })
);
AOI21_X1 #() 
AOI21_X1_3219_ (
  .A({ S25957[652] }),
  .B1({ S25957[649] }),
  .B2({ S4851 }),
  .ZN({ S4965 })
);
AOI21_X1 #() 
AOI21_X1_3220_ (
  .A({ S4798 }),
  .B1({ S4965 }),
  .B2({ S4847 }),
  .ZN({ S4966 })
);
OAI21_X1 #() 
OAI21_X1_2936_ (
  .A({ S4966 }),
  .B1({ S4964 }),
  .B2({ S4803 }),
  .ZN({ S4967 })
);
NAND2_X1 #() 
NAND2_X1_5639_ (
  .A1({ S4967 }),
  .A2({ S4961 }),
  .ZN({ S4968 })
);
NAND2_X1 #() 
NAND2_X1_5640_ (
  .A1({ S4968 }),
  .A2({ S25957[654] }),
  .ZN({ S4969 })
);
NAND2_X1 #() 
NAND2_X1_5641_ (
  .A1({ S4823 }),
  .A2({ S4812 }),
  .ZN({ S4970 })
);
AOI21_X1 #() 
AOI21_X1_3221_ (
  .A({ S4816 }),
  .B1({ S3410 }),
  .B2({ S3407 }),
  .ZN({ S4971 })
);
NOR2_X1 #() 
NOR2_X1_1419_ (
  .A1({ S4868 }),
  .A2({ S4971 }),
  .ZN({ S4972 })
);
AOI21_X1 #() 
AOI21_X1_3222_ (
  .A({ S4972 }),
  .B1({ S4970 }),
  .B2({ S25957[651] }),
  .ZN({ S4973 })
);
AOI21_X1 #() 
AOI21_X1_3223_ (
  .A({ S25957[648] }),
  .B1({ S3477 }),
  .B2({ S3480 }),
  .ZN({ S4974 })
);
AOI21_X1 #() 
AOI21_X1_3224_ (
  .A({ S113 }),
  .B1({ S4806 }),
  .B2({ S4974 }),
  .ZN({ S4975 })
);
AOI211_X1 #() 
AOI211_X1_99_ (
  .A({ S4824 }),
  .B({ S4803 }),
  .C1({ S4975 }),
  .C2({ S4825 }),
  .ZN({ S4976 })
);
AOI21_X1 #() 
AOI21_X1_3225_ (
  .A({ S4976 }),
  .B1({ S4973 }),
  .B2({ S4803 }),
  .ZN({ S4977 })
);
NAND3_X1 #() 
NAND3_X1_6119_ (
  .A1({ S4856 }),
  .A2({ S4812 }),
  .A3({ S4851 }),
  .ZN({ S4978 })
);
NAND2_X1 #() 
NAND2_X1_5642_ (
  .A1({ S4978 }),
  .A2({ S4857 }),
  .ZN({ S4979 })
);
NAND3_X1 #() 
NAND3_X1_6120_ (
  .A1({ S4885 }),
  .A2({ S25957[652] }),
  .A3({ S4868 }),
  .ZN({ S4980 })
);
NAND3_X1 #() 
NAND3_X1_6121_ (
  .A1({ S4980 }),
  .A2({ S4798 }),
  .A3({ S4979 }),
  .ZN({ S4981 })
);
OAI211_X1 #() 
OAI211_X1_1997_ (
  .A({ S4862 }),
  .B({ S4981 }),
  .C1({ S4977 }),
  .C2({ S4798 }),
  .ZN({ S4982 })
);
NAND3_X1 #() 
NAND3_X1_6122_ (
  .A1({ S4982 }),
  .A2({ S3020 }),
  .A3({ S4969 }),
  .ZN({ S4983 })
);
NAND3_X1 #() 
NAND3_X1_6123_ (
  .A1({ S4954 }),
  .A2({ S25957[758] }),
  .A3({ S4983 }),
  .ZN({ S4984 })
);
NAND2_X1 #() 
NAND2_X1_5643_ (
  .A1({ S4982 }),
  .A2({ S4969 }),
  .ZN({ S4985 })
);
NAND2_X1 #() 
NAND2_X1_5644_ (
  .A1({ S4985 }),
  .A2({ S3020 }),
  .ZN({ S4986 })
);
OAI21_X1 #() 
OAI21_X1_2937_ (
  .A({ S4953 }),
  .B1({ S4940 }),
  .B2({ S4862 }),
  .ZN({ S4987 })
);
NAND2_X1 #() 
NAND2_X1_5645_ (
  .A1({ S4987 }),
  .A2({ S25957[655] }),
  .ZN({ S4988 })
);
NAND3_X1 #() 
NAND3_X1_6124_ (
  .A1({ S4988 }),
  .A2({ S2439 }),
  .A3({ S4986 }),
  .ZN({ S4989 })
);
NAND2_X1 #() 
NAND2_X1_5646_ (
  .A1({ S4989 }),
  .A2({ S4984 }),
  .ZN({ S25957[630] })
);
NAND2_X1 #() 
NAND2_X1_5647_ (
  .A1({ S25957[630] }),
  .A2({ S25957[822] }),
  .ZN({ S4990 })
);
INV_X1 #() 
INV_X1_1830_ (
  .A({ S4990 }),
  .ZN({ S4991 })
);
NOR2_X1 #() 
NOR2_X1_1420_ (
  .A1({ S25957[630] }),
  .A2({ S25957[822] }),
  .ZN({ S4992 })
);
OAI21_X1 #() 
OAI21_X1_2938_ (
  .A({ S25957[662] }),
  .B1({ S4991 }),
  .B2({ S4992 }),
  .ZN({ S4993 })
);
NOR2_X1 #() 
NOR2_X1_1421_ (
  .A1({ S4991 }),
  .A2({ S4992 }),
  .ZN({ S25957[566] })
);
NAND2_X1 #() 
NAND2_X1_5648_ (
  .A1({ S25957[566] }),
  .A2({ S2444 }),
  .ZN({ S4994 })
);
NAND2_X1 #() 
NAND2_X1_5649_ (
  .A1({ S4994 }),
  .A2({ S4993 }),
  .ZN({ S25957[534] })
);
NAND2_X1 #() 
NAND2_X1_5650_ (
  .A1({ S2521 }),
  .A2({ S2523 }),
  .ZN({ S4995 })
);
NOR2_X1 #() 
NOR2_X1_1422_ (
  .A1({ S2520 }),
  .A2({ S2518 }),
  .ZN({ S25957[693] })
);
XNOR2_X1 #() 
XNOR2_X1_214_ (
  .A({ S25662 }),
  .B({ S22837 }),
  .ZN({ S25957[853] })
);
INV_X1 #() 
INV_X1_1831_ (
  .A({ S25957[853] }),
  .ZN({ S4996 })
);
NAND4_X1 #() 
NAND4_X1_673_ (
  .A1({ S4812 }),
  .A2({ S4827 }),
  .A3({ S4813 }),
  .A4({ S4799 }),
  .ZN({ S4997 })
);
AND2_X1 #() 
AND2_X1_356_ (
  .A1({ S4997 }),
  .A2({ S4857 }),
  .ZN({ S4998 })
);
NAND3_X1 #() 
NAND3_X1_6125_ (
  .A1({ S4842 }),
  .A2({ S4856 }),
  .A3({ S113 }),
  .ZN({ S4999 })
);
AOI21_X1 #() 
AOI21_X1_3226_ (
  .A({ S4803 }),
  .B1({ S4817 }),
  .B2({ S4794 }),
  .ZN({ S5000 })
);
NAND4_X1 #() 
NAND4_X1_674_ (
  .A1({ S4812 }),
  .A2({ S4803 }),
  .A3({ S5 }),
  .A4({ S113 }),
  .ZN({ S5001 })
);
NAND2_X1 #() 
NAND2_X1_5651_ (
  .A1({ S5001 }),
  .A2({ S25957[653] }),
  .ZN({ S5002 })
);
AOI211_X1 #() 
AOI211_X1_100_ (
  .A({ S5002 }),
  .B({ S4998 }),
  .C1({ S5000 }),
  .C2({ S4999 }),
  .ZN({ S5003 })
);
NAND3_X1 #() 
NAND3_X1_6126_ (
  .A1({ S4812 }),
  .A2({ S25957[651] }),
  .A3({ S4851 }),
  .ZN({ S5004 })
);
AOI21_X1 #() 
AOI21_X1_3227_ (
  .A({ S4803 }),
  .B1({ S4828 }),
  .B2({ S113 }),
  .ZN({ S5005 })
);
NAND2_X1 #() 
NAND2_X1_5652_ (
  .A1({ S5005 }),
  .A2({ S5004 }),
  .ZN({ S5006 })
);
OAI21_X1 #() 
OAI21_X1_2939_ (
  .A({ S5006 }),
  .B1({ S4897 }),
  .B2({ S4957 }),
  .ZN({ S5007 })
);
AOI21_X1 #() 
AOI21_X1_3228_ (
  .A({ S5003 }),
  .B1({ S4798 }),
  .B2({ S5007 }),
  .ZN({ S5008 })
);
NOR2_X1 #() 
NOR2_X1_1423_ (
  .A1({ S5008 }),
  .A2({ S3020 }),
  .ZN({ S5009 })
);
NAND2_X1 #() 
NAND2_X1_5653_ (
  .A1({ S4807 }),
  .A2({ S25957[649] }),
  .ZN({ S5010 })
);
AOI21_X1 #() 
AOI21_X1_3229_ (
  .A({ S113 }),
  .B1({ S4896 }),
  .B2({ S5010 }),
  .ZN({ S5011 })
);
OAI21_X1 #() 
OAI21_X1_2940_ (
  .A({ S25957[652] }),
  .B1({ S5011 }),
  .B2({ S4972 }),
  .ZN({ S5012 })
);
NOR2_X1 #() 
NOR2_X1_1424_ (
  .A1({ S25957[648] }),
  .A2({ S113 }),
  .ZN({ S5013 })
);
NAND2_X1 #() 
NAND2_X1_5654_ (
  .A1({ S4824 }),
  .A2({ S4873 }),
  .ZN({ S5014 })
);
INV_X1 #() 
INV_X1_1832_ (
  .A({ S5014 }),
  .ZN({ S5015 })
);
OAI21_X1 #() 
OAI21_X1_2941_ (
  .A({ S4803 }),
  .B1({ S5015 }),
  .B2({ S5013 }),
  .ZN({ S5016 })
);
NAND3_X1 #() 
NAND3_X1_6127_ (
  .A1({ S5012 }),
  .A2({ S25957[653] }),
  .A3({ S5016 }),
  .ZN({ S5017 })
);
NOR2_X1 #() 
NOR2_X1_1425_ (
  .A1({ S4843 }),
  .A2({ S4803 }),
  .ZN({ S5018 })
);
NAND2_X1 #() 
NAND2_X1_5655_ (
  .A1({ S4946 }),
  .A2({ S113 }),
  .ZN({ S5019 })
);
OAI21_X1 #() 
OAI21_X1_2942_ (
  .A({ S5018 }),
  .B1({ S4814 }),
  .B2({ S5019 }),
  .ZN({ S5020 })
);
NAND3_X1 #() 
NAND3_X1_6128_ (
  .A1({ S4812 }),
  .A2({ S4887 }),
  .A3({ S4851 }),
  .ZN({ S5021 })
);
NAND3_X1 #() 
NAND3_X1_6129_ (
  .A1({ S5021 }),
  .A2({ S4803 }),
  .A3({ S113 }),
  .ZN({ S5022 })
);
AOI21_X1 #() 
AOI21_X1_3230_ (
  .A({ S113 }),
  .B1({ S4816 }),
  .B2({ S25957[648] }),
  .ZN({ S5023 })
);
NAND4_X1 #() 
NAND4_X1_675_ (
  .A1({ S5023 }),
  .A2({ S4811 }),
  .A3({ S4887 }),
  .A4({ S4803 }),
  .ZN({ S5024 })
);
NAND4_X1 #() 
NAND4_X1_676_ (
  .A1({ S5020 }),
  .A2({ S4798 }),
  .A3({ S5022 }),
  .A4({ S5024 }),
  .ZN({ S5025 })
);
AOI21_X1 #() 
AOI21_X1_3231_ (
  .A({ S25957[655] }),
  .B1({ S5017 }),
  .B2({ S5025 }),
  .ZN({ S5026 })
);
OAI21_X1 #() 
OAI21_X1_2943_ (
  .A({ S25957[654] }),
  .B1({ S5009 }),
  .B2({ S5026 }),
  .ZN({ S5027 })
);
NAND2_X1 #() 
NAND2_X1_5656_ (
  .A1({ S4963 }),
  .A2({ S4898 }),
  .ZN({ S5028 })
);
OAI211_X1 #() 
OAI211_X1_1998_ (
  .A({ S5028 }),
  .B({ S25957[652] }),
  .C1({ S113 }),
  .C2({ S4872 }),
  .ZN({ S5029 })
);
AOI21_X1 #() 
AOI21_X1_3232_ (
  .A({ S25957[651] }),
  .B1({ S4825 }),
  .B2({ S4827 }),
  .ZN({ S5030 })
);
OAI21_X1 #() 
OAI21_X1_2944_ (
  .A({ S4803 }),
  .B1({ S5030 }),
  .B2({ S4837 }),
  .ZN({ S5031 })
);
NAND3_X1 #() 
NAND3_X1_6130_ (
  .A1({ S5029 }),
  .A2({ S25957[653] }),
  .A3({ S5031 }),
  .ZN({ S5032 })
);
AOI21_X1 #() 
AOI21_X1_3233_ (
  .A({ S25957[650] }),
  .B1({ S4873 }),
  .B2({ S4811 }),
  .ZN({ S5033 })
);
NAND2_X1 #() 
NAND2_X1_5657_ (
  .A1({ S5033 }),
  .A2({ S25957[651] }),
  .ZN({ S5034 })
);
NAND2_X1 #() 
NAND2_X1_5658_ (
  .A1({ S4824 }),
  .A2({ S4806 }),
  .ZN({ S5035 })
);
AOI21_X1 #() 
AOI21_X1_3234_ (
  .A({ S4803 }),
  .B1({ S5034 }),
  .B2({ S5035 }),
  .ZN({ S5036 })
);
NAND3_X1 #() 
NAND3_X1_6131_ (
  .A1({ S4892 }),
  .A2({ S4808 }),
  .A3({ S4857 }),
  .ZN({ S5037 })
);
OAI21_X1 #() 
OAI21_X1_2945_ (
  .A({ S5037 }),
  .B1({ S4853 }),
  .B2({ S4855 }),
  .ZN({ S5038 })
);
OAI21_X1 #() 
OAI21_X1_2946_ (
  .A({ S4798 }),
  .B1({ S5038 }),
  .B2({ S5036 }),
  .ZN({ S5039 })
);
AOI21_X1 #() 
AOI21_X1_3235_ (
  .A({ S3020 }),
  .B1({ S5039 }),
  .B2({ S5032 }),
  .ZN({ S5040 })
);
AOI21_X1 #() 
AOI21_X1_3236_ (
  .A({ S25957[651] }),
  .B1({ S4807 }),
  .B2({ S25957[649] }),
  .ZN({ S5041 })
);
AOI21_X1 #() 
AOI21_X1_3237_ (
  .A({ S5041 }),
  .B1({ S4814 }),
  .B2({ S25957[651] }),
  .ZN({ S5042 })
);
NAND2_X1 #() 
NAND2_X1_5659_ (
  .A1({ S4887 }),
  .A2({ S113 }),
  .ZN({ S5043 })
);
NAND2_X1 #() 
NAND2_X1_5660_ (
  .A1({ S25957[649] }),
  .A2({ S4851 }),
  .ZN({ S5044 })
);
OAI21_X1 #() 
OAI21_X1_2947_ (
  .A({ S4847 }),
  .B1({ S5044 }),
  .B2({ S5043 }),
  .ZN({ S5045 })
);
NAND2_X1 #() 
NAND2_X1_5661_ (
  .A1({ S5045 }),
  .A2({ S4803 }),
  .ZN({ S5046 })
);
OAI211_X1 #() 
OAI211_X1_1999_ (
  .A({ S5046 }),
  .B({ S25957[653] }),
  .C1({ S5042 }),
  .C2({ S4803 }),
  .ZN({ S5047 })
);
NAND3_X1 #() 
NAND3_X1_6132_ (
  .A1({ S4896 }),
  .A2({ S25957[651] }),
  .A3({ S4883 }),
  .ZN({ S5048 })
);
NAND3_X1 #() 
NAND3_X1_6133_ (
  .A1({ S4844 }),
  .A2({ S4873 }),
  .A3({ S4811 }),
  .ZN({ S5049 })
);
NAND3_X1 #() 
NAND3_X1_6134_ (
  .A1({ S5048 }),
  .A2({ S25957[652] }),
  .A3({ S5049 }),
  .ZN({ S5050 })
);
AOI22_X1 #() 
AOI22_X1_640_ (
  .A1({ S4837 }),
  .A2({ S25957[648] }),
  .B1({ S4971 }),
  .B2({ S4902 }),
  .ZN({ S5051 })
);
OAI211_X1 #() 
OAI211_X1_2000_ (
  .A({ S5050 }),
  .B({ S4798 }),
  .C1({ S25957[652] }),
  .C2({ S5051 }),
  .ZN({ S5052 })
);
AOI21_X1 #() 
AOI21_X1_3238_ (
  .A({ S25957[655] }),
  .B1({ S5052 }),
  .B2({ S5047 }),
  .ZN({ S5053 })
);
OAI21_X1 #() 
OAI21_X1_2948_ (
  .A({ S4862 }),
  .B1({ S5040 }),
  .B2({ S5053 }),
  .ZN({ S5054 })
);
NAND3_X1 #() 
NAND3_X1_6135_ (
  .A1({ S5027 }),
  .A2({ S5054 }),
  .A3({ S4996 }),
  .ZN({ S5055 })
);
INV_X1 #() 
INV_X1_1833_ (
  .A({ S5055 }),
  .ZN({ S5056 })
);
AOI21_X1 #() 
AOI21_X1_3239_ (
  .A({ S4996 }),
  .B1({ S5027 }),
  .B2({ S5054 }),
  .ZN({ S5057 })
);
OAI21_X1 #() 
OAI21_X1_2949_ (
  .A({ S25957[693] }),
  .B1({ S5056 }),
  .B2({ S5057 }),
  .ZN({ S5058 })
);
INV_X1 #() 
INV_X1_1834_ (
  .A({ S25957[693] }),
  .ZN({ S5059 })
);
NAND2_X1 #() 
NAND2_X1_5662_ (
  .A1({ S5027 }),
  .A2({ S5054 }),
  .ZN({ S5060 })
);
NAND2_X1 #() 
NAND2_X1_5663_ (
  .A1({ S5060 }),
  .A2({ S25957[853] }),
  .ZN({ S5061 })
);
NAND3_X1 #() 
NAND3_X1_6136_ (
  .A1({ S5061 }),
  .A2({ S5059 }),
  .A3({ S5055 }),
  .ZN({ S5062 })
);
NAND3_X1 #() 
NAND3_X1_6137_ (
  .A1({ S5058 }),
  .A2({ S5062 }),
  .A3({ S4995 }),
  .ZN({ S5063 })
);
NAND3_X1 #() 
NAND3_X1_6138_ (
  .A1({ S5061 }),
  .A2({ S25957[693] }),
  .A3({ S5055 }),
  .ZN({ S5064 })
);
OAI21_X1 #() 
OAI21_X1_2950_ (
  .A({ S5059 }),
  .B1({ S5056 }),
  .B2({ S5057 }),
  .ZN({ S5065 })
);
NAND3_X1 #() 
NAND3_X1_6139_ (
  .A1({ S5065 }),
  .A2({ S5064 }),
  .A3({ S25957[661] }),
  .ZN({ S5066 })
);
AND2_X1 #() 
AND2_X1_357_ (
  .A1({ S5066 }),
  .A2({ S5063 }),
  .ZN({ S25957[533] })
);
NAND2_X1 #() 
NAND2_X1_5664_ (
  .A1({ S2596 }),
  .A2({ S2597 }),
  .ZN({ S25957[692] })
);
INV_X1 #() 
INV_X1_1835_ (
  .A({ S25957[852] }),
  .ZN({ S5067 })
);
INV_X1 #() 
INV_X1_1836_ (
  .A({ S4997 }),
  .ZN({ S5068 })
);
NAND2_X1 #() 
NAND2_X1_5665_ (
  .A1({ S4970 }),
  .A2({ S4834 }),
  .ZN({ S5069 })
);
OAI21_X1 #() 
OAI21_X1_2951_ (
  .A({ S5069 }),
  .B1({ S5068 }),
  .B2({ S25957[651] }),
  .ZN({ S5070 })
);
NAND3_X1 #() 
NAND3_X1_6140_ (
  .A1({ S5041 }),
  .A2({ S4827 }),
  .A3({ S4799 }),
  .ZN({ S5071 })
);
AOI21_X1 #() 
AOI21_X1_3240_ (
  .A({ S25957[652] }),
  .B1({ S4837 }),
  .B2({ S4799 }),
  .ZN({ S5072 })
);
AOI21_X1 #() 
AOI21_X1_3241_ (
  .A({ S25957[653] }),
  .B1({ S5071 }),
  .B2({ S5072 }),
  .ZN({ S5073 })
);
OAI21_X1 #() 
OAI21_X1_2952_ (
  .A({ S5073 }),
  .B1({ S5070 }),
  .B2({ S4803 }),
  .ZN({ S5074 })
);
NAND2_X1 #() 
NAND2_X1_5666_ (
  .A1({ S4874 }),
  .A2({ S4872 }),
  .ZN({ S5075 })
);
NOR2_X1 #() 
NOR2_X1_1426_ (
  .A1({ S25957[650] }),
  .A2({ S25957[651] }),
  .ZN({ S5076 })
);
OAI21_X1 #() 
OAI21_X1_2953_ (
  .A({ S5010 }),
  .B1({ S4811 }),
  .B2({ S5076 }),
  .ZN({ S5077 })
);
AOI21_X1 #() 
AOI21_X1_3242_ (
  .A({ S4798 }),
  .B1({ S5077 }),
  .B2({ S25957[652] }),
  .ZN({ S5078 })
);
NAND3_X1 #() 
NAND3_X1_6141_ (
  .A1({ S4842 }),
  .A2({ S4856 }),
  .A3({ S4857 }),
  .ZN({ S5079 })
);
OAI211_X1 #() 
OAI211_X1_2001_ (
  .A({ S5078 }),
  .B({ S5079 }),
  .C1({ S5075 }),
  .C2({ S4855 }),
  .ZN({ S5080 })
);
NAND3_X1 #() 
NAND3_X1_6142_ (
  .A1({ S5074 }),
  .A2({ S5080 }),
  .A3({ S4862 }),
  .ZN({ S5081 })
);
NAND2_X1 #() 
NAND2_X1_5667_ (
  .A1({ S4926 }),
  .A2({ S4812 }),
  .ZN({ S5082 })
);
INV_X1 #() 
INV_X1_1837_ (
  .A({ S5082 }),
  .ZN({ S5083 })
);
NAND2_X1 #() 
NAND2_X1_5668_ (
  .A1({ S5023 }),
  .A2({ S4806 }),
  .ZN({ S5084 })
);
INV_X1 #() 
INV_X1_1838_ (
  .A({ S5030 }),
  .ZN({ S5085 })
);
NAND3_X1 #() 
NAND3_X1_6143_ (
  .A1({ S5085 }),
  .A2({ S25957[652] }),
  .A3({ S5084 }),
  .ZN({ S5086 })
);
OAI211_X1 #() 
OAI211_X1_2002_ (
  .A({ S5086 }),
  .B({ S4798 }),
  .C1({ S4910 }),
  .C2({ S5083 }),
  .ZN({ S5087 })
);
AOI21_X1 #() 
AOI21_X1_3243_ (
  .A({ S25957[651] }),
  .B1({ S25957[649] }),
  .B2({ S4816 }),
  .ZN({ S5088 })
);
NAND2_X1 #() 
NAND2_X1_5669_ (
  .A1({ S5088 }),
  .A2({ S4794 }),
  .ZN({ S5089 })
);
INV_X1 #() 
INV_X1_1839_ (
  .A({ S5089 }),
  .ZN({ S5090 })
);
NOR3_X1 #() 
NOR3_X1_179_ (
  .A1({ S5090 }),
  .A2({ S4904 }),
  .A3({ S25957[652] }),
  .ZN({ S5091 })
);
NAND3_X1 #() 
NAND3_X1_6144_ (
  .A1({ S5018 }),
  .A2({ S4800 }),
  .A3({ S5043 }),
  .ZN({ S5092 })
);
NAND2_X1 #() 
NAND2_X1_5670_ (
  .A1({ S5092 }),
  .A2({ S25957[653] }),
  .ZN({ S5093 })
);
OAI211_X1 #() 
OAI211_X1_2003_ (
  .A({ S25957[654] }),
  .B({ S5087 }),
  .C1({ S5093 }),
  .C2({ S5091 }),
  .ZN({ S5094 })
);
NAND3_X1 #() 
NAND3_X1_6145_ (
  .A1({ S5094 }),
  .A2({ S25957[655] }),
  .A3({ S5081 }),
  .ZN({ S5095 })
);
INV_X1 #() 
INV_X1_1840_ (
  .A({ S4850 }),
  .ZN({ S5096 })
);
OAI21_X1 #() 
OAI21_X1_2954_ (
  .A({ S113 }),
  .B1({ S5096 }),
  .B2({ S4863 }),
  .ZN({ S5097 })
);
NAND2_X1 #() 
NAND2_X1_5671_ (
  .A1({ S5097 }),
  .A2({ S4805 }),
  .ZN({ S5098 })
);
NAND2_X1 #() 
NAND2_X1_5672_ (
  .A1({ S4893 }),
  .A2({ S4887 }),
  .ZN({ S5099 })
);
NOR2_X1 #() 
NOR2_X1_1427_ (
  .A1({ S4846 }),
  .A2({ S25957[652] }),
  .ZN({ S5100 })
);
NAND2_X1 #() 
NAND2_X1_5673_ (
  .A1({ S5099 }),
  .A2({ S5100 }),
  .ZN({ S5101 })
);
NAND3_X1 #() 
NAND3_X1_6146_ (
  .A1({ S5098 }),
  .A2({ S5101 }),
  .A3({ S4798 }),
  .ZN({ S5102 })
);
NAND3_X1 #() 
NAND3_X1_6147_ (
  .A1({ S5023 }),
  .A2({ S4887 }),
  .A3({ S4811 }),
  .ZN({ S5103 })
);
OAI21_X1 #() 
OAI21_X1_2955_ (
  .A({ S113 }),
  .B1({ S5033 }),
  .B2({ S4828 }),
  .ZN({ S5104 })
);
NAND3_X1 #() 
NAND3_X1_6148_ (
  .A1({ S5104 }),
  .A2({ S4803 }),
  .A3({ S5103 }),
  .ZN({ S5105 })
);
NAND2_X1 #() 
NAND2_X1_5674_ (
  .A1({ S4816 }),
  .A2({ S136 }),
  .ZN({ S5106 })
);
AOI21_X1 #() 
AOI21_X1_3244_ (
  .A({ S4798 }),
  .B1({ S25957[652] }),
  .B2({ S5106 }),
  .ZN({ S5107 })
);
NAND2_X1 #() 
NAND2_X1_5675_ (
  .A1({ S5105 }),
  .A2({ S5107 }),
  .ZN({ S5108 })
);
AOI21_X1 #() 
AOI21_X1_3245_ (
  .A({ S4862 }),
  .B1({ S5108 }),
  .B2({ S5102 }),
  .ZN({ S5109 })
);
NAND2_X1 #() 
NAND2_X1_5676_ (
  .A1({ S5 }),
  .A2({ S4816 }),
  .ZN({ S5110 })
);
NAND3_X1 #() 
NAND3_X1_6149_ (
  .A1({ S5110 }),
  .A2({ S113 }),
  .A3({ S4850 }),
  .ZN({ S5111 })
);
OAI21_X1 #() 
OAI21_X1_2956_ (
  .A({ S5111 }),
  .B1({ S4931 }),
  .B2({ S4865 }),
  .ZN({ S5112 })
);
NAND3_X1 #() 
NAND3_X1_6150_ (
  .A1({ S5112 }),
  .A2({ S3207 }),
  .A3({ S3209 }),
  .ZN({ S5113 })
);
NAND2_X1 #() 
NAND2_X1_5677_ (
  .A1({ S4842 }),
  .A2({ S4864 }),
  .ZN({ S5114 })
);
NAND3_X1 #() 
NAND3_X1_6151_ (
  .A1({ S5085 }),
  .A2({ S25957[652] }),
  .A3({ S5114 }),
  .ZN({ S5115 })
);
NAND3_X1 #() 
NAND3_X1_6152_ (
  .A1({ S5113 }),
  .A2({ S4798 }),
  .A3({ S5115 }),
  .ZN({ S5116 })
);
OAI21_X1 #() 
OAI21_X1_2957_ (
  .A({ S5034 }),
  .B1({ S25957[651] }),
  .B2({ S4825 }),
  .ZN({ S5117 })
);
AOI22_X1 #() 
AOI22_X1_641_ (
  .A1({ S5117 }),
  .A2({ S4803 }),
  .B1({ S4885 }),
  .B2({ S5005 }),
  .ZN({ S5118 })
);
AOI21_X1 #() 
AOI21_X1_3246_ (
  .A({ S25957[654] }),
  .B1({ S5118 }),
  .B2({ S25957[653] }),
  .ZN({ S5119 })
);
AOI21_X1 #() 
AOI21_X1_3247_ (
  .A({ S5109 }),
  .B1({ S5119 }),
  .B2({ S5116 }),
  .ZN({ S5120 })
);
OAI211_X1 #() 
OAI211_X1_2004_ (
  .A({ S5095 }),
  .B({ S5067 }),
  .C1({ S5120 }),
  .C2({ S25957[655] }),
  .ZN({ S5121 })
);
OAI21_X1 #() 
OAI21_X1_2958_ (
  .A({ S5095 }),
  .B1({ S5120 }),
  .B2({ S25957[655] }),
  .ZN({ S5122 })
);
NAND2_X1 #() 
NAND2_X1_5678_ (
  .A1({ S5122 }),
  .A2({ S25957[852] }),
  .ZN({ S5123 })
);
NAND3_X1 #() 
NAND3_X1_6153_ (
  .A1({ S5123 }),
  .A2({ S2524 }),
  .A3({ S5121 }),
  .ZN({ S5124 })
);
NAND2_X1 #() 
NAND2_X1_5679_ (
  .A1({ S5122 }),
  .A2({ S5067 }),
  .ZN({ S5125 })
);
OAI211_X1 #() 
OAI211_X1_2005_ (
  .A({ S5095 }),
  .B({ S25957[852] }),
  .C1({ S5120 }),
  .C2({ S25957[655] }),
  .ZN({ S5126 })
);
NAND3_X1 #() 
NAND3_X1_6154_ (
  .A1({ S5125 }),
  .A2({ S25957[788] }),
  .A3({ S5126 }),
  .ZN({ S5127 })
);
NAND2_X1 #() 
NAND2_X1_5680_ (
  .A1({ S5124 }),
  .A2({ S5127 }),
  .ZN({ S5128 })
);
INV_X1 #() 
INV_X1_1841_ (
  .A({ S5128 }),
  .ZN({ S25957[532] })
);
NAND2_X1 #() 
NAND2_X1_5681_ (
  .A1({ S2661 }),
  .A2({ S2657 }),
  .ZN({ S5129 })
);
INV_X1 #() 
INV_X1_1842_ (
  .A({ S5129 }),
  .ZN({ S25957[691] })
);
NOR2_X1 #() 
NOR2_X1_1428_ (
  .A1({ S25829 }),
  .A2({ S25830 }),
  .ZN({ S5130 })
);
NAND2_X1 #() 
NAND2_X1_5682_ (
  .A1({ S4928 }),
  .A2({ S4813 }),
  .ZN({ S5131 })
);
NAND2_X1 #() 
NAND2_X1_5683_ (
  .A1({ S4817 }),
  .A2({ S5131 }),
  .ZN({ S5132 })
);
NOR2_X1 #() 
NOR2_X1_1429_ (
  .A1({ S4833 }),
  .A2({ S25957[651] }),
  .ZN({ S5133 })
);
NAND2_X1 #() 
NAND2_X1_5684_ (
  .A1({ S4963 }),
  .A2({ S5133 }),
  .ZN({ S5134 })
);
AOI21_X1 #() 
AOI21_X1_3248_ (
  .A({ S25957[652] }),
  .B1({ S5132 }),
  .B2({ S5134 }),
  .ZN({ S5135 })
);
AOI21_X1 #() 
AOI21_X1_3249_ (
  .A({ S4803 }),
  .B1({ S4864 }),
  .B2({ S5 }),
  .ZN({ S5136 })
);
NAND3_X1 #() 
NAND3_X1_6155_ (
  .A1({ S4856 }),
  .A2({ S113 }),
  .A3({ S4811 }),
  .ZN({ S5137 })
);
NAND2_X1 #() 
NAND2_X1_5685_ (
  .A1({ S5137 }),
  .A2({ S5136 }),
  .ZN({ S5138 })
);
NAND2_X1 #() 
NAND2_X1_5686_ (
  .A1({ S5138 }),
  .A2({ S25957[653] }),
  .ZN({ S5139 })
);
NOR2_X1 #() 
NOR2_X1_1430_ (
  .A1({ S5135 }),
  .A2({ S5139 }),
  .ZN({ S5140 })
);
NAND2_X1 #() 
NAND2_X1_5687_ (
  .A1({ S4834 }),
  .A2({ S4823 }),
  .ZN({ S5141 })
);
NAND3_X1 #() 
NAND3_X1_6156_ (
  .A1({ S4896 }),
  .A2({ S113 }),
  .A3({ S4883 }),
  .ZN({ S5142 })
);
NAND2_X1 #() 
NAND2_X1_5688_ (
  .A1({ S5142 }),
  .A2({ S5141 }),
  .ZN({ S5143 })
);
NAND2_X1 #() 
NAND2_X1_5689_ (
  .A1({ S4962 }),
  .A2({ S5100 }),
  .ZN({ S5144 })
);
NAND2_X1 #() 
NAND2_X1_5690_ (
  .A1({ S5144 }),
  .A2({ S4798 }),
  .ZN({ S5145 })
);
AOI21_X1 #() 
AOI21_X1_3250_ (
  .A({ S5145 }),
  .B1({ S5143 }),
  .B2({ S25957[652] }),
  .ZN({ S5146 })
);
OAI21_X1 #() 
OAI21_X1_2959_ (
  .A({ S25957[654] }),
  .B1({ S5146 }),
  .B2({ S5140 }),
  .ZN({ S5147 })
);
NAND4_X1 #() 
NAND4_X1_677_ (
  .A1({ S4856 }),
  .A2({ S4928 }),
  .A3({ S113 }),
  .A4({ S4812 }),
  .ZN({ S5148 })
);
NAND4_X1 #() 
NAND4_X1_678_ (
  .A1({ S25957[649] }),
  .A2({ S4887 }),
  .A3({ S25957[651] }),
  .A4({ S4851 }),
  .ZN({ S5149 })
);
INV_X1 #() 
INV_X1_1843_ (
  .A({ S5149 }),
  .ZN({ S5150 })
);
NOR2_X1 #() 
NOR2_X1_1431_ (
  .A1({ S5150 }),
  .A2({ S25957[652] }),
  .ZN({ S5151 })
);
NAND2_X1 #() 
NAND2_X1_5691_ (
  .A1({ S4826 }),
  .A2({ S4975 }),
  .ZN({ S5152 })
);
AOI21_X1 #() 
AOI21_X1_3251_ (
  .A({ S4803 }),
  .B1({ S4844 }),
  .B2({ S4928 }),
  .ZN({ S5153 })
);
AOI22_X1 #() 
AOI22_X1_642_ (
  .A1({ S5151 }),
  .A2({ S5148 }),
  .B1({ S5152 }),
  .B2({ S5153 }),
  .ZN({ S5154 })
);
OAI21_X1 #() 
OAI21_X1_2960_ (
  .A({ S113 }),
  .B1({ S4903 }),
  .B2({ S4974 }),
  .ZN({ S5155 })
);
OAI211_X1 #() 
OAI211_X1_2006_ (
  .A({ S5155 }),
  .B({ S25957[652] }),
  .C1({ S113 }),
  .C2({ S4874 }),
  .ZN({ S5156 })
);
NAND2_X1 #() 
NAND2_X1_5692_ (
  .A1({ S4824 }),
  .A2({ S5 }),
  .ZN({ S5157 })
);
NAND2_X1 #() 
NAND2_X1_5693_ (
  .A1({ S4908 }),
  .A2({ S25957[651] }),
  .ZN({ S5158 })
);
OAI211_X1 #() 
OAI211_X1_2007_ (
  .A({ S4803 }),
  .B({ S5157 }),
  .C1({ S4955 }),
  .C2({ S5158 }),
  .ZN({ S5159 })
);
NAND3_X1 #() 
NAND3_X1_6157_ (
  .A1({ S5156 }),
  .A2({ S5159 }),
  .A3({ S4798 }),
  .ZN({ S5160 })
);
OAI211_X1 #() 
OAI211_X1_2008_ (
  .A({ S5160 }),
  .B({ S4862 }),
  .C1({ S5154 }),
  .C2({ S4798 }),
  .ZN({ S5161 })
);
NAND3_X1 #() 
NAND3_X1_6158_ (
  .A1({ S5147 }),
  .A2({ S5161 }),
  .A3({ S25957[655] }),
  .ZN({ S5162 })
);
AOI21_X1 #() 
AOI21_X1_3252_ (
  .A({ S25957[651] }),
  .B1({ S25957[650] }),
  .B2({ S25957[648] }),
  .ZN({ S5163 })
);
INV_X1 #() 
INV_X1_1844_ (
  .A({ S5163 }),
  .ZN({ S5164 })
);
OAI21_X1 #() 
OAI21_X1_2961_ (
  .A({ S25957[652] }),
  .B1({ S5164 }),
  .B2({ S4 }),
  .ZN({ S5165 })
);
AND3_X1 #() 
AND3_X1_247_ (
  .A1({ S4908 }),
  .A2({ S4827 }),
  .A3({ S4902 }),
  .ZN({ S5166 })
);
OAI211_X1 #() 
OAI211_X1_2009_ (
  .A({ S4803 }),
  .B({ S4847 }),
  .C1({ S4842 }),
  .C2({ S113 }),
  .ZN({ S5167 })
);
OAI21_X1 #() 
OAI21_X1_2962_ (
  .A({ S5165 }),
  .B1({ S5167 }),
  .B2({ S5166 }),
  .ZN({ S5168 })
);
NAND2_X1 #() 
NAND2_X1_5694_ (
  .A1({ S4930 }),
  .A2({ S4894 }),
  .ZN({ S5169 })
);
NAND2_X1 #() 
NAND2_X1_5695_ (
  .A1({ S5088 }),
  .A2({ S4811 }),
  .ZN({ S5170 })
);
AOI21_X1 #() 
AOI21_X1_3253_ (
  .A({ S25957[652] }),
  .B1({ S4823 }),
  .B2({ S5013 }),
  .ZN({ S5171 })
);
AOI21_X1 #() 
AOI21_X1_3254_ (
  .A({ S4798 }),
  .B1({ S5170 }),
  .B2({ S5171 }),
  .ZN({ S5172 })
);
NAND2_X1 #() 
NAND2_X1_5696_ (
  .A1({ S5169 }),
  .A2({ S5172 }),
  .ZN({ S5173 })
);
OAI211_X1 #() 
OAI211_X1_2010_ (
  .A({ S5173 }),
  .B({ S25957[654] }),
  .C1({ S25957[653] }),
  .C2({ S5168 }),
  .ZN({ S5174 })
);
NAND2_X1 #() 
NAND2_X1_5697_ (
  .A1({ S4850 }),
  .A2({ S25957[651] }),
  .ZN({ S5175 })
);
OAI211_X1 #() 
OAI211_X1_2011_ (
  .A({ S25957[652] }),
  .B({ S5175 }),
  .C1({ S4870 }),
  .C2({ S25957[651] }),
  .ZN({ S5176 })
);
AND2_X1 #() 
AND2_X1_358_ (
  .A1({ S4928 }),
  .A2({ S25957[651] }),
  .ZN({ S5177 })
);
AOI21_X1 #() 
AOI21_X1_3255_ (
  .A({ S25957[651] }),
  .B1({ S4908 }),
  .B2({ S25957[648] }),
  .ZN({ S5178 })
);
OR2_X1 #() 
OR2_X1_74_ (
  .A1({ S5178 }),
  .A2({ S5177 }),
  .ZN({ S5179 })
);
OAI211_X1 #() 
OAI211_X1_2012_ (
  .A({ S5176 }),
  .B({ S25957[653] }),
  .C1({ S5179 }),
  .C2({ S25957[652] }),
  .ZN({ S5180 })
);
NAND3_X1 #() 
NAND3_X1_6159_ (
  .A1({ S4873 }),
  .A2({ S4811 }),
  .A3({ S4864 }),
  .ZN({ S5181 })
);
INV_X1 #() 
INV_X1_1845_ (
  .A({ S5181 }),
  .ZN({ S5182 })
);
OAI21_X1 #() 
OAI21_X1_2963_ (
  .A({ S25957[652] }),
  .B1({ S5182 }),
  .B2({ S4972 }),
  .ZN({ S5183 })
);
AOI21_X1 #() 
AOI21_X1_3256_ (
  .A({ S4807 }),
  .B1({ S4828 }),
  .B2({ S4811 }),
  .ZN({ S5184 })
);
NAND3_X1 #() 
NAND3_X1_6160_ (
  .A1({ S4853 }),
  .A2({ S25957[651] }),
  .A3({ S4887 }),
  .ZN({ S5185 })
);
OAI211_X1 #() 
OAI211_X1_2013_ (
  .A({ S4803 }),
  .B({ S5185 }),
  .C1({ S5184 }),
  .C2({ S25957[651] }),
  .ZN({ S5186 })
);
NAND3_X1 #() 
NAND3_X1_6161_ (
  .A1({ S5186 }),
  .A2({ S5183 }),
  .A3({ S4798 }),
  .ZN({ S5187 })
);
NAND3_X1 #() 
NAND3_X1_6162_ (
  .A1({ S5180 }),
  .A2({ S5187 }),
  .A3({ S4862 }),
  .ZN({ S5188 })
);
NAND3_X1 #() 
NAND3_X1_6163_ (
  .A1({ S5188 }),
  .A2({ S5174 }),
  .A3({ S3020 }),
  .ZN({ S5189 })
);
NAND3_X1 #() 
NAND3_X1_6164_ (
  .A1({ S5162 }),
  .A2({ S5130 }),
  .A3({ S5189 }),
  .ZN({ S5190 })
);
INV_X1 #() 
INV_X1_1846_ (
  .A({ S5130 }),
  .ZN({ S25957[851] })
);
AOI21_X1 #() 
AOI21_X1_3257_ (
  .A({ S4803 }),
  .B1({ S5142 }),
  .B2({ S5141 }),
  .ZN({ S5191 })
);
OAI21_X1 #() 
OAI21_X1_2964_ (
  .A({ S25957[654] }),
  .B1({ S5191 }),
  .B2({ S5145 }),
  .ZN({ S5192 })
);
NAND3_X1 #() 
NAND3_X1_6165_ (
  .A1({ S5148 }),
  .A2({ S4803 }),
  .A3({ S5149 }),
  .ZN({ S5193 })
);
NAND2_X1 #() 
NAND2_X1_5698_ (
  .A1({ S5152 }),
  .A2({ S5153 }),
  .ZN({ S5194 })
);
NAND3_X1 #() 
NAND3_X1_6166_ (
  .A1({ S5194 }),
  .A2({ S25957[653] }),
  .A3({ S5193 }),
  .ZN({ S5195 })
);
OAI21_X1 #() 
OAI21_X1_2965_ (
  .A({ S5157 }),
  .B1({ S4955 }),
  .B2({ S5158 }),
  .ZN({ S5196 })
);
NAND2_X1 #() 
NAND2_X1_5699_ (
  .A1({ S5196 }),
  .A2({ S4803 }),
  .ZN({ S5197 })
);
OAI21_X1 #() 
OAI21_X1_2966_ (
  .A({ S25957[651] }),
  .B1({ S4842 }),
  .B2({ S4833 }),
  .ZN({ S5198 })
);
AOI21_X1 #() 
AOI21_X1_3258_ (
  .A({ S4803 }),
  .B1({ S4926 }),
  .B2({ S4812 }),
  .ZN({ S5199 })
);
AOI21_X1 #() 
AOI21_X1_3259_ (
  .A({ S25957[653] }),
  .B1({ S5198 }),
  .B2({ S5199 }),
  .ZN({ S5200 })
);
NAND2_X1 #() 
NAND2_X1_5700_ (
  .A1({ S5197 }),
  .A2({ S5200 }),
  .ZN({ S5201 })
);
NAND3_X1 #() 
NAND3_X1_6167_ (
  .A1({ S5201 }),
  .A2({ S5195 }),
  .A3({ S4862 }),
  .ZN({ S5202 })
);
OAI211_X1 #() 
OAI211_X1_2014_ (
  .A({ S5202 }),
  .B({ S25957[655] }),
  .C1({ S5192 }),
  .C2({ S5140 }),
  .ZN({ S5203 })
);
AOI22_X1 #() 
AOI22_X1_643_ (
  .A1({ S4930 }),
  .A2({ S4894 }),
  .B1({ S5170 }),
  .B2({ S5171 }),
  .ZN({ S5204 })
);
NAND2_X1 #() 
NAND2_X1_5701_ (
  .A1({ S5168 }),
  .A2({ S4798 }),
  .ZN({ S5205 })
);
OAI211_X1 #() 
OAI211_X1_2015_ (
  .A({ S5205 }),
  .B({ S25957[654] }),
  .C1({ S5204 }),
  .C2({ S4798 }),
  .ZN({ S5206 })
);
AOI21_X1 #() 
AOI21_X1_3260_ (
  .A({ S4975 }),
  .B1({ S4896 }),
  .B2({ S113 }),
  .ZN({ S5207 })
);
OAI21_X1 #() 
OAI21_X1_2967_ (
  .A({ S4803 }),
  .B1({ S5178 }),
  .B2({ S5177 }),
  .ZN({ S5208 })
);
OAI211_X1 #() 
OAI211_X1_2016_ (
  .A({ S5208 }),
  .B({ S25957[653] }),
  .C1({ S5207 }),
  .C2({ S4803 }),
  .ZN({ S5209 })
);
AOI21_X1 #() 
AOI21_X1_3261_ (
  .A({ S25957[652] }),
  .B1({ S4871 }),
  .B2({ S5185 }),
  .ZN({ S5210 })
);
OAI21_X1 #() 
OAI21_X1_2968_ (
  .A({ S25957[652] }),
  .B1({ S4868 }),
  .B2({ S4971 }),
  .ZN({ S5211 })
);
OAI21_X1 #() 
OAI21_X1_2969_ (
  .A({ S4798 }),
  .B1({ S5211 }),
  .B2({ S5182 }),
  .ZN({ S5212 })
);
OAI211_X1 #() 
OAI211_X1_2017_ (
  .A({ S5209 }),
  .B({ S4862 }),
  .C1({ S5210 }),
  .C2({ S5212 }),
  .ZN({ S5213 })
);
NAND3_X1 #() 
NAND3_X1_6168_ (
  .A1({ S5213 }),
  .A2({ S5206 }),
  .A3({ S3020 }),
  .ZN({ S5214 })
);
NAND3_X1 #() 
NAND3_X1_6169_ (
  .A1({ S5214 }),
  .A2({ S5203 }),
  .A3({ S25957[851] }),
  .ZN({ S5215 })
);
NAND3_X1 #() 
NAND3_X1_6170_ (
  .A1({ S5190 }),
  .A2({ S5215 }),
  .A3({ S25957[691] }),
  .ZN({ S5216 })
);
AOI21_X1 #() 
AOI21_X1_3262_ (
  .A({ S25957[851] }),
  .B1({ S5214 }),
  .B2({ S5203 }),
  .ZN({ S5217 })
);
AOI21_X1 #() 
AOI21_X1_3263_ (
  .A({ S5130 }),
  .B1({ S5162 }),
  .B2({ S5189 }),
  .ZN({ S5218 })
);
OAI21_X1 #() 
OAI21_X1_2970_ (
  .A({ S5129 }),
  .B1({ S5218 }),
  .B2({ S5217 }),
  .ZN({ S5219 })
);
NAND3_X1 #() 
NAND3_X1_6171_ (
  .A1({ S5219 }),
  .A2({ S110 }),
  .A3({ S5216 }),
  .ZN({ S5220 })
);
OAI21_X1 #() 
OAI21_X1_2971_ (
  .A({ S25957[691] }),
  .B1({ S5218 }),
  .B2({ S5217 }),
  .ZN({ S5221 })
);
NAND3_X1 #() 
NAND3_X1_6172_ (
  .A1({ S5190 }),
  .A2({ S5215 }),
  .A3({ S5129 }),
  .ZN({ S5222 })
);
NAND3_X1 #() 
NAND3_X1_6173_ (
  .A1({ S5221 }),
  .A2({ S25957[659] }),
  .A3({ S5222 }),
  .ZN({ S5223 })
);
NAND2_X1 #() 
NAND2_X1_5702_ (
  .A1({ S5220 }),
  .A2({ S5223 }),
  .ZN({ S6 })
);
NAND3_X1 #() 
NAND3_X1_6174_ (
  .A1({ S5219 }),
  .A2({ S25957[659] }),
  .A3({ S5216 }),
  .ZN({ S5224 })
);
NAND3_X1 #() 
NAND3_X1_6175_ (
  .A1({ S5221 }),
  .A2({ S110 }),
  .A3({ S5222 }),
  .ZN({ S5225 })
);
NAND2_X1 #() 
NAND2_X1_5703_ (
  .A1({ S5224 }),
  .A2({ S5225 }),
  .ZN({ S25957[531] })
);
NAND2_X1 #() 
NAND2_X1_5704_ (
  .A1({ S25917 }),
  .A2({ S25914 }),
  .ZN({ S25957[816] })
);
INV_X1 #() 
INV_X1_1847_ (
  .A({ S25957[816] }),
  .ZN({ S5226 })
);
NAND2_X1 #() 
NAND2_X1_5705_ (
  .A1({ S2741 }),
  .A2({ S2716 }),
  .ZN({ S25957[752] })
);
NAND4_X1 #() 
NAND4_X1_679_ (
  .A1({ S4853 }),
  .A2({ S4856 }),
  .A3({ S25957[651] }),
  .A4({ S4928 }),
  .ZN({ S5227 })
);
AOI21_X1 #() 
AOI21_X1_3264_ (
  .A({ S4803 }),
  .B1({ S5227 }),
  .B2({ S4958 }),
  .ZN({ S5228 })
);
INV_X1 #() 
INV_X1_1848_ (
  .A({ S4857 }),
  .ZN({ S5229 })
);
NAND3_X1 #() 
NAND3_X1_6176_ (
  .A1({ S4803 }),
  .A2({ S113 }),
  .A3({ S4807 }),
  .ZN({ S5230 })
);
OAI211_X1 #() 
OAI211_X1_2018_ (
  .A({ S25957[653] }),
  .B({ S5230 }),
  .C1({ S4978 }),
  .C2({ S5229 }),
  .ZN({ S5231 })
);
OAI21_X1 #() 
OAI21_X1_2972_ (
  .A({ S25957[648] }),
  .B1({ S25957[649] }),
  .B2({ S4816 }),
  .ZN({ S5232 })
);
NAND2_X1 #() 
NAND2_X1_5706_ (
  .A1({ S5232 }),
  .A2({ S25957[651] }),
  .ZN({ S5233 })
);
NAND4_X1 #() 
NAND4_X1_680_ (
  .A1({ S4823 }),
  .A2({ S4851 }),
  .A3({ S4812 }),
  .A4({ S113 }),
  .ZN({ S5234 })
);
AOI21_X1 #() 
AOI21_X1_3265_ (
  .A({ S4803 }),
  .B1({ S5233 }),
  .B2({ S5234 }),
  .ZN({ S5235 })
);
NAND3_X1 #() 
NAND3_X1_6177_ (
  .A1({ S5024 }),
  .A2({ S4798 }),
  .A3({ S5001 }),
  .ZN({ S5236 })
);
OAI22_X1 #() 
OAI22_X1_148_ (
  .A1({ S5228 }),
  .A2({ S5231 }),
  .B1({ S5235 }),
  .B2({ S5236 }),
  .ZN({ S5237 })
);
NAND2_X1 #() 
NAND2_X1_5707_ (
  .A1({ S5237 }),
  .A2({ S25957[654] }),
  .ZN({ S5238 })
);
NAND4_X1 #() 
NAND4_X1_681_ (
  .A1({ S4908 }),
  .A2({ S4873 }),
  .A3({ S4811 }),
  .A4({ S25957[651] }),
  .ZN({ S5239 })
);
OAI211_X1 #() 
OAI211_X1_2019_ (
  .A({ S4806 }),
  .B({ S113 }),
  .C1({ S4974 }),
  .C2({ S4852 }),
  .ZN({ S5240 })
);
NAND3_X1 #() 
NAND3_X1_6178_ (
  .A1({ S5239 }),
  .A2({ S5240 }),
  .A3({ S4803 }),
  .ZN({ S5241 })
);
NAND4_X1 #() 
NAND4_X1_682_ (
  .A1({ S4856 }),
  .A2({ S4908 }),
  .A3({ S113 }),
  .A4({ S4928 }),
  .ZN({ S5242 })
);
NAND3_X1 #() 
NAND3_X1_6179_ (
  .A1({ S5198 }),
  .A2({ S5242 }),
  .A3({ S25957[652] }),
  .ZN({ S5243 })
);
NAND3_X1 #() 
NAND3_X1_6180_ (
  .A1({ S5243 }),
  .A2({ S4798 }),
  .A3({ S5241 }),
  .ZN({ S5244 })
);
NAND3_X1 #() 
NAND3_X1_6181_ (
  .A1({ S5049 }),
  .A2({ S4803 }),
  .A3({ S4936 }),
  .ZN({ S5245 })
);
AOI21_X1 #() 
AOI21_X1_3266_ (
  .A({ S4798 }),
  .B1({ S5136 }),
  .B2({ S5014 }),
  .ZN({ S5246 })
);
AOI21_X1 #() 
AOI21_X1_3267_ (
  .A({ S25957[654] }),
  .B1({ S5246 }),
  .B2({ S5245 }),
  .ZN({ S5247 })
);
AOI21_X1 #() 
AOI21_X1_3268_ (
  .A({ S25957[655] }),
  .B1({ S5244 }),
  .B2({ S5247 }),
  .ZN({ S5248 })
);
NAND2_X1 #() 
NAND2_X1_5708_ (
  .A1({ S5238 }),
  .A2({ S5248 }),
  .ZN({ S5249 })
);
NAND2_X1 #() 
NAND2_X1_5709_ (
  .A1({ S5010 }),
  .A2({ S113 }),
  .ZN({ S5250 })
);
NAND3_X1 #() 
NAND3_X1_6182_ (
  .A1({ S5103 }),
  .A2({ S5250 }),
  .A3({ S4803 }),
  .ZN({ S5251 })
);
AOI22_X1 #() 
AOI22_X1_644_ (
  .A1({ S4844 }),
  .A2({ S4928 }),
  .B1({ S4806 }),
  .B2({ S5076 }),
  .ZN({ S5252 })
);
NAND3_X1 #() 
NAND3_X1_6183_ (
  .A1({ S4873 }),
  .A2({ S4811 }),
  .A3({ S4846 }),
  .ZN({ S5253 })
);
NAND3_X1 #() 
NAND3_X1_6184_ (
  .A1({ S5252 }),
  .A2({ S25957[652] }),
  .A3({ S5253 }),
  .ZN({ S5254 })
);
NAND3_X1 #() 
NAND3_X1_6185_ (
  .A1({ S5254 }),
  .A2({ S4798 }),
  .A3({ S5251 }),
  .ZN({ S5255 })
);
AOI21_X1 #() 
AOI21_X1_3269_ (
  .A({ S4803 }),
  .B1({ S4873 }),
  .B2({ S4846 }),
  .ZN({ S5256 })
);
NAND2_X1 #() 
NAND2_X1_5710_ (
  .A1({ S5111 }),
  .A2({ S5256 }),
  .ZN({ S5257 })
);
AOI21_X1 #() 
AOI21_X1_3270_ (
  .A({ S25957[651] }),
  .B1({ S4826 }),
  .B2({ S4823 }),
  .ZN({ S5258 })
);
NAND2_X1 #() 
NAND2_X1_5711_ (
  .A1({ S5114 }),
  .A2({ S4803 }),
  .ZN({ S5259 })
);
OAI211_X1 #() 
OAI211_X1_2020_ (
  .A({ S5257 }),
  .B({ S25957[653] }),
  .C1({ S5258 }),
  .C2({ S5259 }),
  .ZN({ S5260 })
);
NAND3_X1 #() 
NAND3_X1_6186_ (
  .A1({ S5260 }),
  .A2({ S5255 }),
  .A3({ S25957[654] }),
  .ZN({ S5261 })
);
NAND3_X1 #() 
NAND3_X1_6187_ (
  .A1({ S4825 }),
  .A2({ S5 }),
  .A3({ S5076 }),
  .ZN({ S5262 })
);
NAND2_X1 #() 
NAND2_X1_5712_ (
  .A1({ S4823 }),
  .A2({ S5013 }),
  .ZN({ S5263 })
);
NAND4_X1 #() 
NAND4_X1_683_ (
  .A1({ S5 }),
  .A2({ S4813 }),
  .A3({ S113 }),
  .A4({ S4799 }),
  .ZN({ S5264 })
);
NAND2_X1 #() 
NAND2_X1_5713_ (
  .A1({ S5263 }),
  .A2({ S5264 }),
  .ZN({ S5265 })
);
AOI21_X1 #() 
AOI21_X1_3271_ (
  .A({ S4803 }),
  .B1({ S4846 }),
  .B2({ S25957[649] }),
  .ZN({ S5266 })
);
AOI22_X1 #() 
AOI22_X1_645_ (
  .A1({ S5265 }),
  .A2({ S4803 }),
  .B1({ S5266 }),
  .B2({ S5262 }),
  .ZN({ S5267 })
);
NAND4_X1 #() 
NAND4_X1_684_ (
  .A1({ S4883 }),
  .A2({ S4887 }),
  .A3({ S113 }),
  .A4({ S25957[652] }),
  .ZN({ S5268 })
);
AOI21_X1 #() 
AOI21_X1_3272_ (
  .A({ S4798 }),
  .B1({ S5229 }),
  .B2({ S5096 }),
  .ZN({ S5269 })
);
NAND3_X1 #() 
NAND3_X1_6188_ (
  .A1({ S5269 }),
  .A2({ S5268 }),
  .A3({ S5079 }),
  .ZN({ S5270 })
);
OAI211_X1 #() 
OAI211_X1_2021_ (
  .A({ S4862 }),
  .B({ S5270 }),
  .C1({ S5267 }),
  .C2({ S25957[653] }),
  .ZN({ S5271 })
);
NAND3_X1 #() 
NAND3_X1_6189_ (
  .A1({ S5261 }),
  .A2({ S5271 }),
  .A3({ S25957[655] }),
  .ZN({ S5272 })
);
NAND3_X1 #() 
NAND3_X1_6190_ (
  .A1({ S5249 }),
  .A2({ S5272 }),
  .A3({ S25957[752] }),
  .ZN({ S5273 })
);
INV_X1 #() 
INV_X1_1849_ (
  .A({ S25957[752] }),
  .ZN({ S5274 })
);
NAND2_X1 #() 
NAND2_X1_5714_ (
  .A1({ S5249 }),
  .A2({ S5272 }),
  .ZN({ S5275 })
);
NAND2_X1 #() 
NAND2_X1_5715_ (
  .A1({ S5275 }),
  .A2({ S5274 }),
  .ZN({ S5276 })
);
NAND3_X1 #() 
NAND3_X1_6191_ (
  .A1({ S5276 }),
  .A2({ S5226 }),
  .A3({ S5273 }),
  .ZN({ S5277 })
);
NAND3_X1 #() 
NAND3_X1_6192_ (
  .A1({ S5249 }),
  .A2({ S5272 }),
  .A3({ S5274 }),
  .ZN({ S5278 })
);
NAND2_X1 #() 
NAND2_X1_5716_ (
  .A1({ S5275 }),
  .A2({ S25957[752] }),
  .ZN({ S5279 })
);
NAND3_X1 #() 
NAND3_X1_6193_ (
  .A1({ S5279 }),
  .A2({ S25957[816] }),
  .A3({ S5278 }),
  .ZN({ S5280 })
);
NAND3_X1 #() 
NAND3_X1_6194_ (
  .A1({ S5277 }),
  .A2({ S5280 }),
  .A3({ S25957[656] }),
  .ZN({ S5281 })
);
AND2_X1 #() 
AND2_X1_359_ (
  .A1({ S2752 }),
  .A2({ S2746 }),
  .ZN({ S5282 })
);
AOI21_X1 #() 
AOI21_X1_3273_ (
  .A({ S25957[816] }),
  .B1({ S5279 }),
  .B2({ S5278 }),
  .ZN({ S5283 })
);
AOI21_X1 #() 
AOI21_X1_3274_ (
  .A({ S5226 }),
  .B1({ S5276 }),
  .B2({ S5273 }),
  .ZN({ S5284 })
);
OAI21_X1 #() 
OAI21_X1_2973_ (
  .A({ S5282 }),
  .B1({ S5283 }),
  .B2({ S5284 }),
  .ZN({ S5285 })
);
NAND2_X1 #() 
NAND2_X1_5717_ (
  .A1({ S5285 }),
  .A2({ S5281 }),
  .ZN({ S25957[528] })
);
NOR2_X1 #() 
NOR2_X1_1432_ (
  .A1({ S260 }),
  .A2({ S257 }),
  .ZN({ S25957[817] })
);
INV_X1 #() 
INV_X1_1850_ (
  .A({ S25957[817] }),
  .ZN({ S5286 })
);
NAND2_X1 #() 
NAND2_X1_5718_ (
  .A1({ S2816 }),
  .A2({ S2815 }),
  .ZN({ S25957[753] })
);
INV_X1 #() 
INV_X1_1851_ (
  .A({ S25957[753] }),
  .ZN({ S5287 })
);
NAND2_X1 #() 
NAND2_X1_5719_ (
  .A1({ S4824 }),
  .A2({ S4850 }),
  .ZN({ S5288 })
);
NAND2_X1 #() 
NAND2_X1_5720_ (
  .A1({ S5181 }),
  .A2({ S5288 }),
  .ZN({ S5289 })
);
NOR2_X1 #() 
NOR2_X1_1433_ (
  .A1({ S5289 }),
  .A2({ S4803 }),
  .ZN({ S5290 })
);
OAI21_X1 #() 
OAI21_X1_2974_ (
  .A({ S4803 }),
  .B1({ S25957[649] }),
  .B2({ S113 }),
  .ZN({ S5291 })
);
NAND2_X1 #() 
NAND2_X1_5721_ (
  .A1({ S4808 }),
  .A2({ S4799 }),
  .ZN({ S5292 })
);
OAI21_X1 #() 
OAI21_X1_2975_ (
  .A({ S25957[653] }),
  .B1({ S5292 }),
  .B2({ S5291 }),
  .ZN({ S5293 })
);
NOR2_X1 #() 
NOR2_X1_1434_ (
  .A1({ S5290 }),
  .A2({ S5293 }),
  .ZN({ S5294 })
);
NAND3_X1 #() 
NAND3_X1_6195_ (
  .A1({ S4853 }),
  .A2({ S4856 }),
  .A3({ S4928 }),
  .ZN({ S5295 })
);
AOI21_X1 #() 
AOI21_X1_3275_ (
  .A({ S4803 }),
  .B1({ S5295 }),
  .B2({ S25957[651] }),
  .ZN({ S5296 })
);
NAND3_X1 #() 
NAND3_X1_6196_ (
  .A1({ S4808 }),
  .A2({ S113 }),
  .A3({ S4946 }),
  .ZN({ S5297 })
);
AOI21_X1 #() 
AOI21_X1_3276_ (
  .A({ S4898 }),
  .B1({ S4825 }),
  .B2({ S5 }),
  .ZN({ S5298 })
);
NAND4_X1 #() 
NAND4_X1_685_ (
  .A1({ S4811 }),
  .A2({ S4851 }),
  .A3({ S4887 }),
  .A4({ S113 }),
  .ZN({ S5299 })
);
NAND2_X1 #() 
NAND2_X1_5722_ (
  .A1({ S5299 }),
  .A2({ S4803 }),
  .ZN({ S5300 })
);
OAI21_X1 #() 
OAI21_X1_2976_ (
  .A({ S4798 }),
  .B1({ S5300 }),
  .B2({ S5298 }),
  .ZN({ S5301 })
);
AOI21_X1 #() 
AOI21_X1_3277_ (
  .A({ S5301 }),
  .B1({ S5297 }),
  .B2({ S5296 }),
  .ZN({ S5302 })
);
OAI21_X1 #() 
OAI21_X1_2977_ (
  .A({ S25957[654] }),
  .B1({ S5302 }),
  .B2({ S5294 }),
  .ZN({ S5303 })
);
AOI21_X1 #() 
AOI21_X1_3278_ (
  .A({ S4803 }),
  .B1({ S5089 }),
  .B2({ S5149 }),
  .ZN({ S5304 })
);
INV_X1 #() 
INV_X1_1852_ (
  .A({ S5304 }),
  .ZN({ S5305 })
);
NAND3_X1 #() 
NAND3_X1_6197_ (
  .A1({ S5305 }),
  .A2({ S25957[653] }),
  .A3({ S4869 }),
  .ZN({ S5306 })
);
OAI21_X1 #() 
OAI21_X1_2978_ (
  .A({ S25957[652] }),
  .B1({ S5083 }),
  .B2({ S4804 }),
  .ZN({ S5307 })
);
OAI211_X1 #() 
OAI211_X1_2022_ (
  .A({ S5307 }),
  .B({ S4798 }),
  .C1({ S4869 }),
  .C2({ S4817 }),
  .ZN({ S5308 })
);
NAND3_X1 #() 
NAND3_X1_6198_ (
  .A1({ S5306 }),
  .A2({ S5308 }),
  .A3({ S4862 }),
  .ZN({ S5309 })
);
AOI21_X1 #() 
AOI21_X1_3279_ (
  .A({ S25957[655] }),
  .B1({ S5303 }),
  .B2({ S5309 }),
  .ZN({ S5310 })
);
NAND2_X1 #() 
NAND2_X1_5723_ (
  .A1({ S4874 }),
  .A2({ S5163 }),
  .ZN({ S5311 })
);
AOI21_X1 #() 
AOI21_X1_3280_ (
  .A({ S25957[652] }),
  .B1({ S4834 }),
  .B2({ S4887 }),
  .ZN({ S5312 })
);
NAND2_X1 #() 
NAND2_X1_5724_ (
  .A1({ S5311 }),
  .A2({ S5312 }),
  .ZN({ S5313 })
);
NAND2_X1 #() 
NAND2_X1_5725_ (
  .A1({ S5010 }),
  .A2({ S25957[651] }),
  .ZN({ S5314 })
);
NAND3_X1 #() 
NAND3_X1_6199_ (
  .A1({ S4823 }),
  .A2({ S113 }),
  .A3({ S4794 }),
  .ZN({ S5315 })
);
OAI211_X1 #() 
OAI211_X1_2023_ (
  .A({ S25957[652] }),
  .B({ S5315 }),
  .C1({ S4870 }),
  .C2({ S5314 }),
  .ZN({ S5316 })
);
NAND3_X1 #() 
NAND3_X1_6200_ (
  .A1({ S5316 }),
  .A2({ S5313 }),
  .A3({ S4798 }),
  .ZN({ S5317 })
);
AOI21_X1 #() 
AOI21_X1_3281_ (
  .A({ S113 }),
  .B1({ S4892 }),
  .B2({ S4853 }),
  .ZN({ S5318 })
);
OAI21_X1 #() 
OAI21_X1_2979_ (
  .A({ S4803 }),
  .B1({ S4881 }),
  .B2({ S25957[651] }),
  .ZN({ S5319 })
);
AOI21_X1 #() 
AOI21_X1_3282_ (
  .A({ S4803 }),
  .B1({ S4926 }),
  .B2({ S4827 }),
  .ZN({ S5320 })
);
AOI21_X1 #() 
AOI21_X1_3283_ (
  .A({ S4798 }),
  .B1({ S5141 }),
  .B2({ S5320 }),
  .ZN({ S5321 })
);
OAI21_X1 #() 
OAI21_X1_2980_ (
  .A({ S5321 }),
  .B1({ S5318 }),
  .B2({ S5319 }),
  .ZN({ S5322 })
);
NAND3_X1 #() 
NAND3_X1_6201_ (
  .A1({ S5317 }),
  .A2({ S5322 }),
  .A3({ S25957[654] }),
  .ZN({ S5323 })
);
AOI21_X1 #() 
AOI21_X1_3284_ (
  .A({ S113 }),
  .B1({ S4896 }),
  .B2({ S4813 }),
  .ZN({ S5324 })
);
NAND3_X1 #() 
NAND3_X1_6202_ (
  .A1({ S5170 }),
  .A2({ S4803 }),
  .A3({ S5004 }),
  .ZN({ S5325 })
);
OAI211_X1 #() 
OAI211_X1_2024_ (
  .A({ S25957[653] }),
  .B({ S5325 }),
  .C1({ S5324 }),
  .C2({ S4882 }),
  .ZN({ S5326 })
);
NAND2_X1 #() 
NAND2_X1_5726_ (
  .A1({ S5071 }),
  .A2({ S4803 }),
  .ZN({ S5327 })
);
NAND3_X1 #() 
NAND3_X1_6203_ (
  .A1({ S5010 }),
  .A2({ S113 }),
  .A3({ S4827 }),
  .ZN({ S5328 })
);
AOI21_X1 #() 
AOI21_X1_3285_ (
  .A({ S25957[653] }),
  .B1({ S5328 }),
  .B2({ S4959 }),
  .ZN({ S5329 })
);
OAI21_X1 #() 
OAI21_X1_2981_ (
  .A({ S5329 }),
  .B1({ S5327 }),
  .B2({ S4875 }),
  .ZN({ S5330 })
);
NAND3_X1 #() 
NAND3_X1_6204_ (
  .A1({ S5326 }),
  .A2({ S5330 }),
  .A3({ S4862 }),
  .ZN({ S5331 })
);
AND3_X1 #() 
AND3_X1_248_ (
  .A1({ S5331 }),
  .A2({ S5323 }),
  .A3({ S25957[655] }),
  .ZN({ S5332 })
);
OAI21_X1 #() 
OAI21_X1_2982_ (
  .A({ S5287 }),
  .B1({ S5310 }),
  .B2({ S5332 }),
  .ZN({ S5333 })
);
OAI221_X1 #() 
OAI221_X1_169_ (
  .A({ S25957[653] }),
  .B1({ S5292 }),
  .B2({ S5291 }),
  .C1({ S5289 }),
  .C2({ S4803 }),
  .ZN({ S5334 })
);
AOI22_X1 #() 
AOI22_X1_646_ (
  .A1({ S4888 }),
  .A2({ S5 }),
  .B1({ S25957[648] }),
  .B2({ S4863 }),
  .ZN({ S5335 })
);
OAI211_X1 #() 
OAI211_X1_2025_ (
  .A({ S25957[652] }),
  .B({ S5297 }),
  .C1({ S5335 }),
  .C2({ S113 }),
  .ZN({ S5336 })
);
AOI21_X1 #() 
AOI21_X1_3286_ (
  .A({ S25957[652] }),
  .B1({ S4963 }),
  .B2({ S4824 }),
  .ZN({ S5337 })
);
AOI21_X1 #() 
AOI21_X1_3287_ (
  .A({ S25957[653] }),
  .B1({ S5337 }),
  .B2({ S5253 }),
  .ZN({ S5338 })
);
NAND2_X1 #() 
NAND2_X1_5727_ (
  .A1({ S5338 }),
  .A2({ S5336 }),
  .ZN({ S5339 })
);
AOI21_X1 #() 
AOI21_X1_3288_ (
  .A({ S4862 }),
  .B1({ S5339 }),
  .B2({ S5334 }),
  .ZN({ S5340 })
);
INV_X1 #() 
INV_X1_1853_ (
  .A({ S4804 }),
  .ZN({ S5341 })
);
AOI21_X1 #() 
AOI21_X1_3289_ (
  .A({ S4803 }),
  .B1({ S5341 }),
  .B2({ S5082 }),
  .ZN({ S5342 })
);
NOR2_X1 #() 
NOR2_X1_1435_ (
  .A1({ S4869 }),
  .A2({ S4817 }),
  .ZN({ S5343 })
);
OAI21_X1 #() 
OAI21_X1_2983_ (
  .A({ S4798 }),
  .B1({ S5343 }),
  .B2({ S5342 }),
  .ZN({ S5344 })
);
OAI21_X1 #() 
OAI21_X1_2984_ (
  .A({ S25957[653] }),
  .B1({ S4925 }),
  .B2({ S5304 }),
  .ZN({ S5345 })
);
AOI21_X1 #() 
AOI21_X1_3290_ (
  .A({ S25957[654] }),
  .B1({ S5344 }),
  .B2({ S5345 }),
  .ZN({ S5346 })
);
OAI21_X1 #() 
OAI21_X1_2985_ (
  .A({ S3020 }),
  .B1({ S5346 }),
  .B2({ S5340 }),
  .ZN({ S5347 })
);
NAND3_X1 #() 
NAND3_X1_6205_ (
  .A1({ S5331 }),
  .A2({ S5323 }),
  .A3({ S25957[655] }),
  .ZN({ S5348 })
);
NAND3_X1 #() 
NAND3_X1_6206_ (
  .A1({ S5347 }),
  .A2({ S25957[753] }),
  .A3({ S5348 }),
  .ZN({ S5349 })
);
NAND3_X1 #() 
NAND3_X1_6207_ (
  .A1({ S5333 }),
  .A2({ S5349 }),
  .A3({ S5286 }),
  .ZN({ S5350 })
);
NAND3_X1 #() 
NAND3_X1_6208_ (
  .A1({ S5347 }),
  .A2({ S5287 }),
  .A3({ S5348 }),
  .ZN({ S5351 })
);
OAI21_X1 #() 
OAI21_X1_2986_ (
  .A({ S25957[753] }),
  .B1({ S5310 }),
  .B2({ S5332 }),
  .ZN({ S5352 })
);
NAND3_X1 #() 
NAND3_X1_6209_ (
  .A1({ S5352 }),
  .A2({ S5351 }),
  .A3({ S25957[817] }),
  .ZN({ S5353 })
);
NAND3_X1 #() 
NAND3_X1_6210_ (
  .A1({ S5350 }),
  .A2({ S5353 }),
  .A3({ S25957[657] }),
  .ZN({ S5354 })
);
AOI21_X1 #() 
AOI21_X1_3291_ (
  .A({ S2753 }),
  .B1({ S2816 }),
  .B2({ S2815 }),
  .ZN({ S5355 })
);
AOI21_X1 #() 
AOI21_X1_3292_ (
  .A({ S25957[849] }),
  .B1({ S2813 }),
  .B2({ S2798 }),
  .ZN({ S5356 })
);
OAI21_X1 #() 
OAI21_X1_2987_ (
  .A({ S264 }),
  .B1({ S5355 }),
  .B2({ S5356 }),
  .ZN({ S5357 })
);
NAND3_X1 #() 
NAND3_X1_6211_ (
  .A1({ S2814 }),
  .A2({ S2817 }),
  .A3({ S25957[913] }),
  .ZN({ S5358 })
);
NAND2_X1 #() 
NAND2_X1_5728_ (
  .A1({ S5357 }),
  .A2({ S5358 }),
  .ZN({ S5359 })
);
AOI21_X1 #() 
AOI21_X1_3293_ (
  .A({ S25957[817] }),
  .B1({ S5352 }),
  .B2({ S5351 }),
  .ZN({ S5360 })
);
AOI21_X1 #() 
AOI21_X1_3294_ (
  .A({ S5286 }),
  .B1({ S5333 }),
  .B2({ S5349 }),
  .ZN({ S5361 })
);
OAI21_X1 #() 
OAI21_X1_2988_ (
  .A({ S5359 }),
  .B1({ S5360 }),
  .B2({ S5361 }),
  .ZN({ S5362 })
);
NAND2_X1 #() 
NAND2_X1_5729_ (
  .A1({ S5362 }),
  .A2({ S5354 }),
  .ZN({ S25957[529] })
);
NOR2_X1 #() 
NOR2_X1_1436_ (
  .A1({ S340 }),
  .A2({ S343 }),
  .ZN({ S25957[818] })
);
INV_X1 #() 
INV_X1_1854_ (
  .A({ S25957[818] }),
  .ZN({ S5363 })
);
NAND2_X1 #() 
NAND2_X1_5730_ (
  .A1({ S315 }),
  .A2({ S339 }),
  .ZN({ S25957[882] })
);
NAND2_X1 #() 
NAND2_X1_5731_ (
  .A1({ S2885 }),
  .A2({ S2874 }),
  .ZN({ S5364 })
);
OR2_X1 #() 
OR2_X1_75_ (
  .A1({ S5364 }),
  .A2({ S25957[882] }),
  .ZN({ S5365 })
);
NAND2_X1 #() 
NAND2_X1_5732_ (
  .A1({ S5364 }),
  .A2({ S25957[882] }),
  .ZN({ S5366 })
);
NAND2_X1 #() 
NAND2_X1_5733_ (
  .A1({ S5365 }),
  .A2({ S5366 }),
  .ZN({ S25957[754] })
);
NAND3_X1 #() 
NAND3_X1_6212_ (
  .A1({ S4827 }),
  .A2({ S25957[651] }),
  .A3({ S4799 }),
  .ZN({ S5367 })
);
OAI211_X1 #() 
OAI211_X1_2026_ (
  .A({ S4906 }),
  .B({ S4803 }),
  .C1({ S5033 }),
  .C2({ S5367 }),
  .ZN({ S5368 })
);
INV_X1 #() 
INV_X1_1855_ (
  .A({ S4866 }),
  .ZN({ S5369 })
);
AOI21_X1 #() 
AOI21_X1_3295_ (
  .A({ S4971 }),
  .B1({ S4814 }),
  .B2({ S5 }),
  .ZN({ S5370 })
);
OAI211_X1 #() 
OAI211_X1_2027_ (
  .A({ S5369 }),
  .B({ S25957[652] }),
  .C1({ S5370 }),
  .C2({ S25957[651] }),
  .ZN({ S5371 })
);
NAND3_X1 #() 
NAND3_X1_6213_ (
  .A1({ S5371 }),
  .A2({ S25957[653] }),
  .A3({ S5368 }),
  .ZN({ S5372 })
);
NAND2_X1 #() 
NAND2_X1_5734_ (
  .A1({ S4806 }),
  .A2({ S5076 }),
  .ZN({ S5373 })
);
NAND3_X1 #() 
NAND3_X1_6214_ (
  .A1({ S4909 }),
  .A2({ S4803 }),
  .A3({ S5373 }),
  .ZN({ S5374 })
);
NAND2_X1 #() 
NAND2_X1_5735_ (
  .A1({ S4811 }),
  .A2({ S25957[650] }),
  .ZN({ S5375 })
);
NAND3_X1 #() 
NAND3_X1_6215_ (
  .A1({ S4826 }),
  .A2({ S25957[651] }),
  .A3({ S5375 }),
  .ZN({ S5376 })
);
INV_X1 #() 
INV_X1_1856_ (
  .A({ S5376 }),
  .ZN({ S5377 })
);
NAND2_X1 #() 
NAND2_X1_5736_ (
  .A1({ S4851 }),
  .A2({ S113 }),
  .ZN({ S5378 })
);
OAI21_X1 #() 
OAI21_X1_2989_ (
  .A({ S25957[652] }),
  .B1({ S5378 }),
  .B2({ S25957[649] }),
  .ZN({ S5379 })
);
OAI211_X1 #() 
OAI211_X1_2028_ (
  .A({ S5374 }),
  .B({ S4798 }),
  .C1({ S5377 }),
  .C2({ S5379 }),
  .ZN({ S5380 })
);
NAND3_X1 #() 
NAND3_X1_6216_ (
  .A1({ S5372 }),
  .A2({ S5380 }),
  .A3({ S25957[654] }),
  .ZN({ S5381 })
);
NOR3_X1 #() 
NOR3_X1_180_ (
  .A1({ S4903 }),
  .A2({ S4794 }),
  .A3({ S113 }),
  .ZN({ S5382 })
);
NOR3_X1 #() 
NOR3_X1_181_ (
  .A1({ S5382 }),
  .A2({ S5166 }),
  .A3({ S4803 }),
  .ZN({ S5383 })
);
AOI21_X1 #() 
AOI21_X1_3296_ (
  .A({ S25957[651] }),
  .B1({ S5 }),
  .B2({ S25957[650] }),
  .ZN({ S5384 })
);
INV_X1 #() 
INV_X1_1857_ (
  .A({ S5384 }),
  .ZN({ S5385 })
);
NAND2_X1 #() 
NAND2_X1_5737_ (
  .A1({ S4928 }),
  .A2({ S25957[651] }),
  .ZN({ S5386 })
);
OAI21_X1 #() 
OAI21_X1_2990_ (
  .A({ S5385 }),
  .B1({ S4833 }),
  .B2({ S5386 }),
  .ZN({ S5387 })
);
OAI21_X1 #() 
OAI21_X1_2991_ (
  .A({ S25957[653] }),
  .B1({ S5387 }),
  .B2({ S25957[652] }),
  .ZN({ S5388 })
);
AND3_X1 #() 
AND3_X1_249_ (
  .A1({ S25957[649] }),
  .A2({ S25957[651] }),
  .A3({ S4851 }),
  .ZN({ S5389 })
);
OAI21_X1 #() 
OAI21_X1_2992_ (
  .A({ S25957[652] }),
  .B1({ S5389 }),
  .B2({ S5088 }),
  .ZN({ S5390 })
);
OAI21_X1 #() 
OAI21_X1_2993_ (
  .A({ S5390 }),
  .B1({ S4943 }),
  .B2({ S25957[652] }),
  .ZN({ S5391 })
);
NAND2_X1 #() 
NAND2_X1_5738_ (
  .A1({ S5391 }),
  .A2({ S4798 }),
  .ZN({ S5392 })
);
OAI211_X1 #() 
OAI211_X1_2029_ (
  .A({ S5392 }),
  .B({ S4862 }),
  .C1({ S5383 }),
  .C2({ S5388 }),
  .ZN({ S5393 })
);
NAND3_X1 #() 
NAND3_X1_6217_ (
  .A1({ S5393 }),
  .A2({ S5381 }),
  .A3({ S25957[655] }),
  .ZN({ S5394 })
);
INV_X1 #() 
INV_X1_1858_ (
  .A({ S4965 }),
  .ZN({ S5395 })
);
NAND2_X1 #() 
NAND2_X1_5739_ (
  .A1({ S5021 }),
  .A2({ S25957[652] }),
  .ZN({ S5396 })
);
AOI21_X1 #() 
AOI21_X1_3297_ (
  .A({ S113 }),
  .B1({ S5396 }),
  .B2({ S5395 }),
  .ZN({ S5397 })
);
NAND4_X1 #() 
NAND4_X1_686_ (
  .A1({ S4853 }),
  .A2({ S4928 }),
  .A3({ S25957[652] }),
  .A4({ S113 }),
  .ZN({ S5398 })
);
OAI211_X1 #() 
OAI211_X1_2030_ (
  .A({ S5398 }),
  .B({ S4798 }),
  .C1({ S5252 }),
  .C2({ S25957[652] }),
  .ZN({ S5399 })
);
NAND3_X1 #() 
NAND3_X1_6218_ (
  .A1({ S4908 }),
  .A2({ S113 }),
  .A3({ S25957[648] }),
  .ZN({ S5400 })
);
NAND2_X1 #() 
NAND2_X1_5740_ (
  .A1({ S5400 }),
  .A2({ S4803 }),
  .ZN({ S5401 })
);
AOI21_X1 #() 
AOI21_X1_3298_ (
  .A({ S5401 }),
  .B1({ S4829 }),
  .B2({ S4826 }),
  .ZN({ S5402 })
);
OAI211_X1 #() 
OAI211_X1_2031_ (
  .A({ S3407 }),
  .B({ S3410 }),
  .C1({ S4816 }),
  .C2({ S25957[648] }),
  .ZN({ S5403 })
);
AOI22_X1 #() 
AOI22_X1_647_ (
  .A1({ S5403 }),
  .A2({ S25957[651] }),
  .B1({ S4825 }),
  .B2({ S5163 }),
  .ZN({ S5404 })
);
OAI21_X1 #() 
OAI21_X1_2994_ (
  .A({ S25957[653] }),
  .B1({ S5404 }),
  .B2({ S4803 }),
  .ZN({ S5405 })
);
OAI22_X1 #() 
OAI22_X1_149_ (
  .A1({ S5402 }),
  .A2({ S5405 }),
  .B1({ S5399 }),
  .B2({ S5397 }),
  .ZN({ S5406 })
);
NAND2_X1 #() 
NAND2_X1_5741_ (
  .A1({ S5406 }),
  .A2({ S25957[654] }),
  .ZN({ S5407 })
);
OAI22_X1 #() 
OAI22_X1_150_ (
  .A1({ S4932 }),
  .A2({ S4867 }),
  .B1({ S5010 }),
  .B2({ S25957[651] }),
  .ZN({ S5408 })
);
NAND2_X1 #() 
NAND2_X1_5742_ (
  .A1({ S4808 }),
  .A2({ S4864 }),
  .ZN({ S5409 })
);
NAND3_X1 #() 
NAND3_X1_6219_ (
  .A1({ S5148 }),
  .A2({ S5409 }),
  .A3({ S25957[652] }),
  .ZN({ S5410 })
);
OAI211_X1 #() 
OAI211_X1_2032_ (
  .A({ S5410 }),
  .B({ S25957[653] }),
  .C1({ S5408 }),
  .C2({ S25957[652] }),
  .ZN({ S5411 })
);
AOI21_X1 #() 
AOI21_X1_3299_ (
  .A({ S5389 }),
  .B1({ S4997 }),
  .B2({ S113 }),
  .ZN({ S5412 })
);
NAND4_X1 #() 
NAND4_X1_687_ (
  .A1({ S4826 }),
  .A2({ S4823 }),
  .A3({ S113 }),
  .A4({ S4803 }),
  .ZN({ S5413 })
);
OAI211_X1 #() 
OAI211_X1_2033_ (
  .A({ S5413 }),
  .B({ S4979 }),
  .C1({ S5412 }),
  .C2({ S4803 }),
  .ZN({ S5414 })
);
NAND2_X1 #() 
NAND2_X1_5743_ (
  .A1({ S5414 }),
  .A2({ S4798 }),
  .ZN({ S5415 })
);
NAND3_X1 #() 
NAND3_X1_6220_ (
  .A1({ S5415 }),
  .A2({ S4862 }),
  .A3({ S5411 }),
  .ZN({ S5416 })
);
NAND3_X1 #() 
NAND3_X1_6221_ (
  .A1({ S5416 }),
  .A2({ S5407 }),
  .A3({ S3020 }),
  .ZN({ S5417 })
);
NAND3_X1 #() 
NAND3_X1_6222_ (
  .A1({ S5417 }),
  .A2({ S5394 }),
  .A3({ S25957[754] }),
  .ZN({ S5418 })
);
INV_X1 #() 
INV_X1_1859_ (
  .A({ S25957[754] }),
  .ZN({ S5419 })
);
OAI21_X1 #() 
OAI21_X1_2995_ (
  .A({ S25957[652] }),
  .B1({ S5258 }),
  .B2({ S4866 }),
  .ZN({ S5420 })
);
OAI21_X1 #() 
OAI21_X1_2996_ (
  .A({ S4906 }),
  .B1({ S5033 }),
  .B2({ S5367 }),
  .ZN({ S5421 })
);
AOI21_X1 #() 
AOI21_X1_3300_ (
  .A({ S4798 }),
  .B1({ S5421 }),
  .B2({ S4803 }),
  .ZN({ S5422 })
);
NAND2_X1 #() 
NAND2_X1_5744_ (
  .A1({ S5422 }),
  .A2({ S5420 }),
  .ZN({ S5423 })
);
INV_X1 #() 
INV_X1_1860_ (
  .A({ S5374 }),
  .ZN({ S5424 })
);
AOI21_X1 #() 
AOI21_X1_3301_ (
  .A({ S5379 }),
  .B1({ S4815 }),
  .B2({ S25957[651] }),
  .ZN({ S5425 })
);
OAI21_X1 #() 
OAI21_X1_2997_ (
  .A({ S4798 }),
  .B1({ S5425 }),
  .B2({ S5424 }),
  .ZN({ S5426 })
);
NAND3_X1 #() 
NAND3_X1_6223_ (
  .A1({ S5423 }),
  .A2({ S5426 }),
  .A3({ S25957[654] }),
  .ZN({ S5427 })
);
OAI211_X1 #() 
OAI211_X1_2034_ (
  .A({ S5390 }),
  .B({ S4798 }),
  .C1({ S4943 }),
  .C2({ S25957[652] }),
  .ZN({ S5428 })
);
OAI21_X1 #() 
OAI21_X1_2998_ (
  .A({ S25957[652] }),
  .B1({ S5382 }),
  .B2({ S5166 }),
  .ZN({ S5429 })
);
NOR2_X1 #() 
NOR2_X1_1437_ (
  .A1({ S5386 }),
  .A2({ S4833 }),
  .ZN({ S5430 })
);
OAI21_X1 #() 
OAI21_X1_2999_ (
  .A({ S4803 }),
  .B1({ S5430 }),
  .B2({ S5384 }),
  .ZN({ S5431 })
);
NAND3_X1 #() 
NAND3_X1_6224_ (
  .A1({ S5429 }),
  .A2({ S5431 }),
  .A3({ S25957[653] }),
  .ZN({ S5432 })
);
NAND3_X1 #() 
NAND3_X1_6225_ (
  .A1({ S5432 }),
  .A2({ S5428 }),
  .A3({ S4862 }),
  .ZN({ S5433 })
);
NAND3_X1 #() 
NAND3_X1_6226_ (
  .A1({ S5427 }),
  .A2({ S25957[655] }),
  .A3({ S5433 }),
  .ZN({ S5434 })
);
AOI21_X1 #() 
AOI21_X1_3302_ (
  .A({ S4965 }),
  .B1({ S5021 }),
  .B2({ S25957[652] }),
  .ZN({ S5435 })
);
NAND3_X1 #() 
NAND3_X1_6227_ (
  .A1({ S5375 }),
  .A2({ S4812 }),
  .A3({ S4851 }),
  .ZN({ S5436 })
);
NAND3_X1 #() 
NAND3_X1_6228_ (
  .A1({ S5436 }),
  .A2({ S4803 }),
  .A3({ S113 }),
  .ZN({ S5437 })
);
AND2_X1 #() 
AND2_X1_360_ (
  .A1({ S4928 }),
  .A2({ S25957[652] }),
  .ZN({ S5438 })
);
AOI21_X1 #() 
AOI21_X1_3303_ (
  .A({ S25957[653] }),
  .B1({ S5438 }),
  .B2({ S4893 }),
  .ZN({ S5439 })
);
OAI211_X1 #() 
OAI211_X1_2035_ (
  .A({ S5437 }),
  .B({ S5439 }),
  .C1({ S5435 }),
  .C2({ S113 }),
  .ZN({ S5440 })
);
OAI211_X1 #() 
OAI211_X1_2036_ (
  .A({ S5440 }),
  .B({ S25957[654] }),
  .C1({ S5402 }),
  .C2({ S5405 }),
  .ZN({ S5441 })
);
AOI21_X1 #() 
AOI21_X1_3304_ (
  .A({ S25957[653] }),
  .B1({ S4978 }),
  .B2({ S4857 }),
  .ZN({ S5442 })
);
OAI211_X1 #() 
OAI211_X1_2037_ (
  .A({ S5442 }),
  .B({ S5413 }),
  .C1({ S5412 }),
  .C2({ S4803 }),
  .ZN({ S5443 })
);
NAND2_X1 #() 
NAND2_X1_5745_ (
  .A1({ S5148 }),
  .A2({ S5409 }),
  .ZN({ S5444 })
);
NAND2_X1 #() 
NAND2_X1_5746_ (
  .A1({ S5444 }),
  .A2({ S25957[652] }),
  .ZN({ S5445 })
);
NAND2_X1 #() 
NAND2_X1_5747_ (
  .A1({ S5408 }),
  .A2({ S4803 }),
  .ZN({ S5446 })
);
NAND3_X1 #() 
NAND3_X1_6229_ (
  .A1({ S5445 }),
  .A2({ S5446 }),
  .A3({ S25957[653] }),
  .ZN({ S5447 })
);
NAND3_X1 #() 
NAND3_X1_6230_ (
  .A1({ S5447 }),
  .A2({ S4862 }),
  .A3({ S5443 }),
  .ZN({ S5448 })
);
NAND3_X1 #() 
NAND3_X1_6231_ (
  .A1({ S5448 }),
  .A2({ S5441 }),
  .A3({ S3020 }),
  .ZN({ S5449 })
);
NAND3_X1 #() 
NAND3_X1_6232_ (
  .A1({ S5434 }),
  .A2({ S5419 }),
  .A3({ S5449 }),
  .ZN({ S5450 })
);
NAND3_X1 #() 
NAND3_X1_6233_ (
  .A1({ S5418 }),
  .A2({ S5450 }),
  .A3({ S5363 }),
  .ZN({ S5451 })
);
NAND3_X1 #() 
NAND3_X1_6234_ (
  .A1({ S5417 }),
  .A2({ S5394 }),
  .A3({ S5419 }),
  .ZN({ S5452 })
);
NAND3_X1 #() 
NAND3_X1_6235_ (
  .A1({ S5434 }),
  .A2({ S25957[754] }),
  .A3({ S5449 }),
  .ZN({ S5453 })
);
NAND3_X1 #() 
NAND3_X1_6236_ (
  .A1({ S5452 }),
  .A2({ S5453 }),
  .A3({ S25957[818] }),
  .ZN({ S5454 })
);
NAND3_X1 #() 
NAND3_X1_6237_ (
  .A1({ S5451 }),
  .A2({ S5454 }),
  .A3({ S25957[658] }),
  .ZN({ S5455 })
);
AOI21_X1 #() 
AOI21_X1_3305_ (
  .A({ S25957[914] }),
  .B1({ S2888 }),
  .B2({ S2889 }),
  .ZN({ S5456 })
);
AND3_X1 #() 
AND3_X1_250_ (
  .A1({ S2888 }),
  .A2({ S25957[914] }),
  .A3({ S2889 }),
  .ZN({ S5457 })
);
NOR2_X1 #() 
NOR2_X1_1438_ (
  .A1({ S5457 }),
  .A2({ S5456 }),
  .ZN({ S5458 })
);
AOI21_X1 #() 
AOI21_X1_3306_ (
  .A({ S25957[818] }),
  .B1({ S5452 }),
  .B2({ S5453 }),
  .ZN({ S5459 })
);
AOI21_X1 #() 
AOI21_X1_3307_ (
  .A({ S5363 }),
  .B1({ S5418 }),
  .B2({ S5450 }),
  .ZN({ S5460 })
);
OAI21_X1 #() 
OAI21_X1_3000_ (
  .A({ S5458 }),
  .B1({ S5459 }),
  .B2({ S5460 }),
  .ZN({ S5461 })
);
NAND2_X1 #() 
NAND2_X1_5748_ (
  .A1({ S5461 }),
  .A2({ S5455 }),
  .ZN({ S25957[530] })
);
OAI21_X1 #() 
OAI21_X1_3001_ (
  .A({ S490 }),
  .B1({ S4060 }),
  .B2({ S4061 }),
  .ZN({ S5462 })
);
NAND3_X1 #() 
NAND3_X1_6238_ (
  .A1({ S4077 }),
  .A2({ S25957[897] }),
  .A3({ S4063 }),
  .ZN({ S5463 })
);
NAND2_X1 #() 
NAND2_X1_5749_ (
  .A1({ S5462 }),
  .A2({ S5463 }),
  .ZN({ S5464 })
);
AOI21_X1 #() 
AOI21_X1_3308_ (
  .A({ S5464 }),
  .B1({ S4021 }),
  .B2({ S4018 }),
  .ZN({ S7 })
);
NAND3_X1 #() 
NAND3_X1_6239_ (
  .A1({ S4018 }),
  .A2({ S4021 }),
  .A3({ S5464 }),
  .ZN({ S8 })
);
XOR2_X1 #() 
XOR2_X1_98_ (
  .A({ S25957[847] }),
  .B({ S25957[943] }),
  .Z({ S25957[815] })
);
INV_X1 #() 
INV_X1_1861_ (
  .A({ S25957[646] }),
  .ZN({ S5465 })
);
NAND2_X1 #() 
NAND2_X1_5750_ (
  .A1({ S25957[643] }),
  .A2({ S5464 }),
  .ZN({ S5466 })
);
NAND4_X1 #() 
NAND4_X1_688_ (
  .A1({ S25957[640] }),
  .A2({ S3926 }),
  .A3({ S3929 }),
  .A4({ S25957[642] }),
  .ZN({ S5467 })
);
NAND2_X1 #() 
NAND2_X1_5751_ (
  .A1({ S5466 }),
  .A2({ S5467 }),
  .ZN({ S5468 })
);
AOI21_X1 #() 
AOI21_X1_3309_ (
  .A({ S25957[898] }),
  .B1({ S4162 }),
  .B2({ S4161 }),
  .ZN({ S5469 })
);
AND3_X1 #() 
AND3_X1_251_ (
  .A1({ S4162 }),
  .A2({ S4161 }),
  .A3({ S25957[898] }),
  .ZN({ S5470 })
);
NOR2_X1 #() 
NOR2_X1_1439_ (
  .A1({ S5470 }),
  .A2({ S5469 }),
  .ZN({ S5471 })
);
AOI21_X1 #() 
AOI21_X1_3310_ (
  .A({ S5471 }),
  .B1({ S4021 }),
  .B2({ S4018 }),
  .ZN({ S5472 })
);
NAND3_X1 #() 
NAND3_X1_6240_ (
  .A1({ S3930 }),
  .A2({ S3931 }),
  .A3({ S25957[641] }),
  .ZN({ S5473 })
);
OAI21_X1 #() 
OAI21_X1_3002_ (
  .A({ S25957[644] }),
  .B1({ S5472 }),
  .B2({ S5473 }),
  .ZN({ S5474 })
);
NAND3_X1 #() 
NAND3_X1_6241_ (
  .A1({ S5471 }),
  .A2({ S4018 }),
  .A3({ S4021 }),
  .ZN({ S5475 })
);
AOI22_X1 #() 
AOI22_X1_648_ (
  .A1({ S0 }),
  .A2({ S5475 }),
  .B1({ S3849 }),
  .B2({ S3846 }),
  .ZN({ S5476 })
);
AOI21_X1 #() 
AOI21_X1_3311_ (
  .A({ S25957[896] }),
  .B1({ S4019 }),
  .B2({ S4020 }),
  .ZN({ S5477 })
);
AOI21_X1 #() 
AOI21_X1_3312_ (
  .A({ S499 }),
  .B1({ S4013 }),
  .B2({ S4017 }),
  .ZN({ S5478 })
);
NOR2_X1 #() 
NOR2_X1_1440_ (
  .A1({ S5477 }),
  .A2({ S5478 }),
  .ZN({ S5479 })
);
NAND2_X1 #() 
NAND2_X1_5752_ (
  .A1({ S25957[643] }),
  .A2({ S5479 }),
  .ZN({ S5480 })
);
INV_X1 #() 
INV_X1_1862_ (
  .A({ S5480 }),
  .ZN({ S5481 })
);
OAI21_X1 #() 
OAI21_X1_3003_ (
  .A({ S5476 }),
  .B1({ S5481 }),
  .B2({ S5464 }),
  .ZN({ S5482 })
);
OAI211_X1 #() 
OAI211_X1_2038_ (
  .A({ S5482 }),
  .B({ S25957[645] }),
  .C1({ S5468 }),
  .C2({ S5474 }),
  .ZN({ S5483 })
);
NAND3_X1 #() 
NAND3_X1_6242_ (
  .A1({ S25957[642] }),
  .A2({ S4018 }),
  .A3({ S4021 }),
  .ZN({ S5484 })
);
NAND2_X1 #() 
NAND2_X1_5753_ (
  .A1({ S25957[642] }),
  .A2({ S25957[641] }),
  .ZN({ S5485 })
);
NAND2_X1 #() 
NAND2_X1_5754_ (
  .A1({ S5484 }),
  .A2({ S5485 }),
  .ZN({ S5486 })
);
INV_X1 #() 
INV_X1_1863_ (
  .A({ S5486 }),
  .ZN({ S5487 })
);
OAI21_X1 #() 
OAI21_X1_3004_ (
  .A({ S25957[641] }),
  .B1({ S5477 }),
  .B2({ S5478 }),
  .ZN({ S5488 })
);
NAND3_X1 #() 
NAND3_X1_6243_ (
  .A1({ S5488 }),
  .A2({ S5471 }),
  .A3({ S8 }),
  .ZN({ S5489 })
);
NAND3_X1 #() 
NAND3_X1_6244_ (
  .A1({ S5487 }),
  .A2({ S5489 }),
  .A3({ S0 }),
  .ZN({ S5490 })
);
NOR2_X1 #() 
NOR2_X1_1441_ (
  .A1({ S25957[642] }),
  .A2({ S25957[641] }),
  .ZN({ S5491 })
);
NAND2_X1 #() 
NAND2_X1_5755_ (
  .A1({ S25957[643] }),
  .A2({ S5491 }),
  .ZN({ S5492 })
);
AOI21_X1 #() 
AOI21_X1_3313_ (
  .A({ S25957[644] }),
  .B1({ S5490 }),
  .B2({ S5492 }),
  .ZN({ S5493 })
);
NAND2_X1 #() 
NAND2_X1_5756_ (
  .A1({ S3751 }),
  .A2({ S3754 }),
  .ZN({ S5494 })
);
NAND2_X1 #() 
NAND2_X1_5757_ (
  .A1({ S3846 }),
  .A2({ S3849 }),
  .ZN({ S5495 })
);
AOI22_X1 #() 
AOI22_X1_649_ (
  .A1({ S4160 }),
  .A2({ S4163 }),
  .B1({ S4062 }),
  .B2({ S4078 }),
  .ZN({ S5496 })
);
NAND3_X1 #() 
NAND3_X1_6245_ (
  .A1({ S4018 }),
  .A2({ S4021 }),
  .A3({ S25957[641] }),
  .ZN({ S5497 })
);
OAI21_X1 #() 
OAI21_X1_3005_ (
  .A({ S5464 }),
  .B1({ S5477 }),
  .B2({ S5478 }),
  .ZN({ S5498 })
);
AOI21_X1 #() 
AOI21_X1_3314_ (
  .A({ S25957[642] }),
  .B1({ S5498 }),
  .B2({ S5497 }),
  .ZN({ S5499 })
);
NAND4_X1 #() 
NAND4_X1_689_ (
  .A1({ S25957[642] }),
  .A2({ S5464 }),
  .A3({ S4021 }),
  .A4({ S4018 }),
  .ZN({ S5500 })
);
NAND2_X1 #() 
NAND2_X1_5758_ (
  .A1({ S25957[640] }),
  .A2({ S5496 }),
  .ZN({ S5501 })
);
NAND3_X1 #() 
NAND3_X1_6246_ (
  .A1({ S5501 }),
  .A2({ S25957[643] }),
  .A3({ S5500 }),
  .ZN({ S5502 })
);
NAND2_X1 #() 
NAND2_X1_5759_ (
  .A1({ S25957[640] }),
  .A2({ S5471 }),
  .ZN({ S5503 })
);
NAND2_X1 #() 
NAND2_X1_5760_ (
  .A1({ S5503 }),
  .A2({ S0 }),
  .ZN({ S5504 })
);
OAI22_X1 #() 
OAI22_X1_151_ (
  .A1({ S5499 }),
  .A2({ S5502 }),
  .B1({ S5504 }),
  .B2({ S5496 }),
  .ZN({ S5505 })
);
OAI21_X1 #() 
OAI21_X1_3006_ (
  .A({ S5494 }),
  .B1({ S5505 }),
  .B2({ S5495 }),
  .ZN({ S5506 })
);
OAI211_X1 #() 
OAI211_X1_2039_ (
  .A({ S5465 }),
  .B({ S5483 }),
  .C1({ S5506 }),
  .C2({ S5493 }),
  .ZN({ S5507 })
);
NAND3_X1 #() 
NAND3_X1_6247_ (
  .A1({ S5464 }),
  .A2({ S4160 }),
  .A3({ S4163 }),
  .ZN({ S5508 })
);
OAI211_X1 #() 
OAI211_X1_2040_ (
  .A({ S25957[643] }),
  .B({ S5484 }),
  .C1({ S5479 }),
  .C2({ S5508 }),
  .ZN({ S5509 })
);
OAI21_X1 #() 
OAI21_X1_3007_ (
  .A({ S25957[641] }),
  .B1({ S25957[640] }),
  .B2({ S25957[642] }),
  .ZN({ S5510 })
);
OAI21_X1 #() 
OAI21_X1_3008_ (
  .A({ S5509 }),
  .B1({ S25957[643] }),
  .B2({ S5510 }),
  .ZN({ S5511 })
);
NAND4_X1 #() 
NAND4_X1_690_ (
  .A1({ S25957[642] }),
  .A2({ S25957[641] }),
  .A3({ S4021 }),
  .A4({ S4018 }),
  .ZN({ S5512 })
);
NAND3_X1 #() 
NAND3_X1_6248_ (
  .A1({ S5498 }),
  .A2({ S25957[643] }),
  .A3({ S5512 }),
  .ZN({ S5513 })
);
NAND2_X1 #() 
NAND2_X1_5761_ (
  .A1({ S8 }),
  .A2({ S25957[642] }),
  .ZN({ S5514 })
);
NAND2_X1 #() 
NAND2_X1_5762_ (
  .A1({ S5488 }),
  .A2({ S5471 }),
  .ZN({ S5515 })
);
NAND2_X1 #() 
NAND2_X1_5763_ (
  .A1({ S5515 }),
  .A2({ S5514 }),
  .ZN({ S5516 })
);
AOI21_X1 #() 
AOI21_X1_3315_ (
  .A({ S25957[644] }),
  .B1({ S5516 }),
  .B2({ S0 }),
  .ZN({ S5517 })
);
AOI22_X1 #() 
AOI22_X1_650_ (
  .A1({ S5517 }),
  .A2({ S5513 }),
  .B1({ S5511 }),
  .B2({ S25957[644] }),
  .ZN({ S5518 })
);
AOI21_X1 #() 
AOI21_X1_3316_ (
  .A({ S25957[641] }),
  .B1({ S4160 }),
  .B2({ S4163 }),
  .ZN({ S5519 })
);
NOR2_X1 #() 
NOR2_X1_1442_ (
  .A1({ S0 }),
  .A2({ S5519 }),
  .ZN({ S5520 })
);
INV_X1 #() 
INV_X1_1864_ (
  .A({ S5497 }),
  .ZN({ S5521 })
);
NOR2_X1 #() 
NOR2_X1_1443_ (
  .A1({ S5521 }),
  .A2({ S25957[643] }),
  .ZN({ S5522 })
);
AOI211_X1 #() 
AOI211_X1_101_ (
  .A({ S5495 }),
  .B({ S5522 }),
  .C1({ S5488 }),
  .C2({ S5520 }),
  .ZN({ S5523 })
);
AOI21_X1 #() 
AOI21_X1_3317_ (
  .A({ S25957[641] }),
  .B1({ S4021 }),
  .B2({ S4018 }),
  .ZN({ S5524 })
);
NAND2_X1 #() 
NAND2_X1_5764_ (
  .A1({ S8 }),
  .A2({ S5471 }),
  .ZN({ S5525 })
);
AOI22_X1 #() 
AOI22_X1_651_ (
  .A1({ S5525 }),
  .A2({ S5500 }),
  .B1({ S25957[643] }),
  .B2({ S5524 }),
  .ZN({ S5526 })
);
OAI21_X1 #() 
OAI21_X1_3009_ (
  .A({ S5494 }),
  .B1({ S5526 }),
  .B2({ S25957[644] }),
  .ZN({ S5527 })
);
OAI22_X1 #() 
OAI22_X1_152_ (
  .A1({ S5518 }),
  .A2({ S5494 }),
  .B1({ S5523 }),
  .B2({ S5527 }),
  .ZN({ S5528 })
);
OAI211_X1 #() 
OAI211_X1_2041_ (
  .A({ S25957[647] }),
  .B({ S5507 }),
  .C1({ S5528 }),
  .C2({ S5465 }),
  .ZN({ S5529 })
);
AND2_X1 #() 
AND2_X1_361_ (
  .A1({ S3604 }),
  .A2({ S3601 }),
  .ZN({ S5530 })
);
INV_X1 #() 
INV_X1_1865_ (
  .A({ S5475 }),
  .ZN({ S5531 })
);
NAND2_X1 #() 
NAND2_X1_5765_ (
  .A1({ S0 }),
  .A2({ S5512 }),
  .ZN({ S5532 })
);
OAI21_X1 #() 
OAI21_X1_3010_ (
  .A({ S25957[644] }),
  .B1({ S5532 }),
  .B2({ S5531 }),
  .ZN({ S5533 })
);
AOI21_X1 #() 
AOI21_X1_3318_ (
  .A({ S5533 }),
  .B1({ S5516 }),
  .B2({ S25957[643] }),
  .ZN({ S5534 })
);
NAND2_X1 #() 
NAND2_X1_5766_ (
  .A1({ S5491 }),
  .A2({ S25957[640] }),
  .ZN({ S5535 })
);
NAND3_X1 #() 
NAND3_X1_6249_ (
  .A1({ S5535 }),
  .A2({ S25957[643] }),
  .A3({ S5485 }),
  .ZN({ S5536 })
);
NAND2_X1 #() 
NAND2_X1_5767_ (
  .A1({ S25957[642] }),
  .A2({ S5464 }),
  .ZN({ S5537 })
);
NAND2_X1 #() 
NAND2_X1_5768_ (
  .A1({ S5484 }),
  .A2({ S5537 }),
  .ZN({ S5538 })
);
NAND2_X1 #() 
NAND2_X1_5769_ (
  .A1({ S5538 }),
  .A2({ S0 }),
  .ZN({ S5539 })
);
AOI21_X1 #() 
AOI21_X1_3319_ (
  .A({ S25957[644] }),
  .B1({ S5536 }),
  .B2({ S5539 }),
  .ZN({ S5540 })
);
OAI21_X1 #() 
OAI21_X1_3011_ (
  .A({ S25957[645] }),
  .B1({ S5534 }),
  .B2({ S5540 }),
  .ZN({ S5541 })
);
NAND2_X1 #() 
NAND2_X1_5770_ (
  .A1({ S5488 }),
  .A2({ S25957[642] }),
  .ZN({ S5542 })
);
NAND2_X1 #() 
NAND2_X1_5771_ (
  .A1({ S5479 }),
  .A2({ S5508 }),
  .ZN({ S5543 })
);
NAND4_X1 #() 
NAND4_X1_691_ (
  .A1({ S4160 }),
  .A2({ S4163 }),
  .A3({ S5462 }),
  .A4({ S5463 }),
  .ZN({ S5544 })
);
NAND2_X1 #() 
NAND2_X1_5772_ (
  .A1({ S25957[640] }),
  .A2({ S5544 }),
  .ZN({ S5545 })
);
NAND2_X1 #() 
NAND2_X1_5773_ (
  .A1({ S5543 }),
  .A2({ S5545 }),
  .ZN({ S5546 })
);
AOI21_X1 #() 
AOI21_X1_3320_ (
  .A({ S0 }),
  .B1({ S5546 }),
  .B2({ S5542 }),
  .ZN({ S5547 })
);
NAND3_X1 #() 
NAND3_X1_6250_ (
  .A1({ S5498 }),
  .A2({ S25957[642] }),
  .A3({ S5497 }),
  .ZN({ S5548 })
);
AOI21_X1 #() 
AOI21_X1_3321_ (
  .A({ S25957[643] }),
  .B1({ S5548 }),
  .B2({ S5475 }),
  .ZN({ S5549 })
);
OR3_X1 #() 
OR3_X1_38_ (
  .A1({ S5547 }),
  .A2({ S5549 }),
  .A3({ S5495 }),
  .ZN({ S5550 })
);
INV_X1 #() 
INV_X1_1866_ (
  .A({ S5544 }),
  .ZN({ S5551 })
);
NOR2_X1 #() 
NOR2_X1_1444_ (
  .A1({ S5472 }),
  .A2({ S0 }),
  .ZN({ S5552 })
);
INV_X1 #() 
INV_X1_1867_ (
  .A({ S5552 }),
  .ZN({ S5553 })
);
NAND3_X1 #() 
NAND3_X1_6251_ (
  .A1({ S5537 }),
  .A2({ S25957[640] }),
  .A3({ S5544 }),
  .ZN({ S5554 })
);
AOI21_X1 #() 
AOI21_X1_3322_ (
  .A({ S25957[644] }),
  .B1({ S0 }),
  .B2({ S5554 }),
  .ZN({ S5555 })
);
OAI21_X1 #() 
OAI21_X1_3012_ (
  .A({ S5555 }),
  .B1({ S5551 }),
  .B2({ S5553 }),
  .ZN({ S5556 })
);
NAND3_X1 #() 
NAND3_X1_6252_ (
  .A1({ S5550 }),
  .A2({ S5494 }),
  .A3({ S5556 }),
  .ZN({ S5557 })
);
AOI21_X1 #() 
AOI21_X1_3323_ (
  .A({ S5465 }),
  .B1({ S5557 }),
  .B2({ S5541 }),
  .ZN({ S5558 })
);
NOR2_X1 #() 
NOR2_X1_1445_ (
  .A1({ S25957[643] }),
  .A2({ S5496 }),
  .ZN({ S5559 })
);
NAND2_X1 #() 
NAND2_X1_5774_ (
  .A1({ S8 }),
  .A2({ S5485 }),
  .ZN({ S5560 })
);
NAND2_X1 #() 
NAND2_X1_5775_ (
  .A1({ S5560 }),
  .A2({ S25957[643] }),
  .ZN({ S5561 })
);
INV_X1 #() 
INV_X1_1868_ (
  .A({ S5561 }),
  .ZN({ S5562 })
);
AOI21_X1 #() 
AOI21_X1_3324_ (
  .A({ S5562 }),
  .B1({ S5559 }),
  .B2({ S5515 }),
  .ZN({ S5563 })
);
NAND2_X1 #() 
NAND2_X1_5776_ (
  .A1({ S0 }),
  .A2({ S25957[640] }),
  .ZN({ S5564 })
);
NAND2_X1 #() 
NAND2_X1_5777_ (
  .A1({ S25957[640] }),
  .A2({ S25957[642] }),
  .ZN({ S5565 })
);
NAND3_X1 #() 
NAND3_X1_6253_ (
  .A1({ S5565 }),
  .A2({ S25957[643] }),
  .A3({ S5508 }),
  .ZN({ S5566 })
);
NAND3_X1 #() 
NAND3_X1_6254_ (
  .A1({ S5566 }),
  .A2({ S25957[644] }),
  .A3({ S5564 }),
  .ZN({ S5567 })
);
OAI211_X1 #() 
OAI211_X1_2042_ (
  .A({ S25957[645] }),
  .B({ S5567 }),
  .C1({ S5563 }),
  .C2({ S25957[644] }),
  .ZN({ S5568 })
);
NOR2_X1 #() 
NOR2_X1_1446_ (
  .A1({ S5542 }),
  .A2({ S0 }),
  .ZN({ S5569 })
);
NAND4_X1 #() 
NAND4_X1_692_ (
  .A1({ S5498 }),
  .A2({ S0 }),
  .A3({ S5497 }),
  .A4({ S25957[642] }),
  .ZN({ S5570 })
);
NAND2_X1 #() 
NAND2_X1_5778_ (
  .A1({ S5570 }),
  .A2({ S5495 }),
  .ZN({ S5571 })
);
INV_X1 #() 
INV_X1_1869_ (
  .A({ S5512 }),
  .ZN({ S5572 })
);
NAND3_X1 #() 
NAND3_X1_6255_ (
  .A1({ S25957[640] }),
  .A2({ S25957[641] }),
  .A3({ S5471 }),
  .ZN({ S5573 })
);
OAI211_X1 #() 
OAI211_X1_2043_ (
  .A({ S0 }),
  .B({ S5573 }),
  .C1({ S5514 }),
  .C2({ S7 }),
  .ZN({ S5574 })
);
OAI211_X1 #() 
OAI211_X1_2044_ (
  .A({ S5574 }),
  .B({ S25957[644] }),
  .C1({ S0 }),
  .C2({ S5572 }),
  .ZN({ S5575 })
);
OAI211_X1 #() 
OAI211_X1_2045_ (
  .A({ S5575 }),
  .B({ S5494 }),
  .C1({ S5569 }),
  .C2({ S5571 }),
  .ZN({ S5576 })
);
AND3_X1 #() 
AND3_X1_252_ (
  .A1({ S5568 }),
  .A2({ S5465 }),
  .A3({ S5576 }),
  .ZN({ S5577 })
);
OAI21_X1 #() 
OAI21_X1_3013_ (
  .A({ S5530 }),
  .B1({ S5558 }),
  .B2({ S5577 }),
  .ZN({ S5578 })
);
NAND2_X1 #() 
NAND2_X1_5779_ (
  .A1({ S5578 }),
  .A2({ S5529 }),
  .ZN({ S5579 })
);
XNOR2_X1 #() 
XNOR2_X1_215_ (
  .A({ S5579 }),
  .B({ S25957[751] }),
  .ZN({ S25957[623] })
);
AND2_X1 #() 
AND2_X1_362_ (
  .A1({ S25957[623] }),
  .A2({ S25957[815] }),
  .ZN({ S5580 })
);
NOR2_X1 #() 
NOR2_X1_1447_ (
  .A1({ S25957[623] }),
  .A2({ S25957[815] }),
  .ZN({ S5581 })
);
NOR2_X1 #() 
NOR2_X1_1448_ (
  .A1({ S5580 }),
  .A2({ S5581 }),
  .ZN({ S25957[559] })
);
INV_X1 #() 
INV_X1_1870_ (
  .A({ S25957[559] }),
  .ZN({ S5582 })
);
NAND2_X1 #() 
NAND2_X1_5780_ (
  .A1({ S5582 }),
  .A2({ S25957[655] }),
  .ZN({ S5583 })
);
NAND2_X1 #() 
NAND2_X1_5781_ (
  .A1({ S25957[559] }),
  .A2({ S3020 }),
  .ZN({ S5584 })
);
NAND2_X1 #() 
NAND2_X1_5782_ (
  .A1({ S5583 }),
  .A2({ S5584 }),
  .ZN({ S25957[527] })
);
NOR2_X1 #() 
NOR2_X1_1449_ (
  .A1({ S556 }),
  .A2({ S552 }),
  .ZN({ S25957[814] })
);
XNOR2_X1 #() 
XNOR2_X1_216_ (
  .A({ S3084 }),
  .B({ S23548 }),
  .ZN({ S25957[718] })
);
XOR2_X1 #() 
XOR2_X1_99_ (
  .A({ S25957[718] }),
  .B({ S25957[814] }),
  .Z({ S25957[686] })
);
NAND2_X1 #() 
NAND2_X1_5783_ (
  .A1({ S549 }),
  .A2({ S550 }),
  .ZN({ S25957[878] })
);
XOR2_X1 #() 
XOR2_X1_100_ (
  .A({ S3084 }),
  .B({ S25957[878] }),
  .Z({ S25957[750] })
);
NAND3_X1 #() 
NAND3_X1_6256_ (
  .A1({ S5537 }),
  .A2({ S3926 }),
  .A3({ S3929 }),
  .ZN({ S5585 })
);
AND2_X1 #() 
AND2_X1_363_ (
  .A1({ S5495 }),
  .A2({ S5473 }),
  .ZN({ S5586 })
);
OAI21_X1 #() 
OAI21_X1_3014_ (
  .A({ S5586 }),
  .B1({ S7 }),
  .B2({ S5585 }),
  .ZN({ S5587 })
);
INV_X1 #() 
INV_X1_1871_ (
  .A({ S5503 }),
  .ZN({ S5588 })
);
OAI21_X1 #() 
OAI21_X1_3015_ (
  .A({ S25957[643] }),
  .B1({ S5588 }),
  .B2({ S5486 }),
  .ZN({ S5589 })
);
NAND2_X1 #() 
NAND2_X1_5784_ (
  .A1({ S5514 }),
  .A2({ S0 }),
  .ZN({ S5590 })
);
AOI21_X1 #() 
AOI21_X1_3325_ (
  .A({ S5495 }),
  .B1({ S25957[643] }),
  .B2({ S5551 }),
  .ZN({ S5591 })
);
NAND3_X1 #() 
NAND3_X1_6257_ (
  .A1({ S5589 }),
  .A2({ S5591 }),
  .A3({ S5590 }),
  .ZN({ S5592 })
);
NAND3_X1 #() 
NAND3_X1_6258_ (
  .A1({ S5592 }),
  .A2({ S5587 }),
  .A3({ S25957[645] }),
  .ZN({ S5593 })
);
NAND2_X1 #() 
NAND2_X1_5785_ (
  .A1({ S0 }),
  .A2({ S5484 }),
  .ZN({ S5594 })
);
INV_X1 #() 
INV_X1_1872_ (
  .A({ S5594 }),
  .ZN({ S5595 })
);
NAND2_X1 #() 
NAND2_X1_5786_ (
  .A1({ S5546 }),
  .A2({ S5595 }),
  .ZN({ S5596 })
);
NAND3_X1 #() 
NAND3_X1_6259_ (
  .A1({ S5596 }),
  .A2({ S25957[644] }),
  .A3({ S5589 }),
  .ZN({ S5597 })
);
NOR2_X1 #() 
NOR2_X1_1450_ (
  .A1({ S5510 }),
  .A2({ S0 }),
  .ZN({ S5598 })
);
NAND2_X1 #() 
NAND2_X1_5787_ (
  .A1({ S5555 }),
  .A2({ S5467 }),
  .ZN({ S5599 })
);
OAI211_X1 #() 
OAI211_X1_2046_ (
  .A({ S5597 }),
  .B({ S5494 }),
  .C1({ S5599 }),
  .C2({ S5598 }),
  .ZN({ S5600 })
);
NAND3_X1 #() 
NAND3_X1_6260_ (
  .A1({ S5600 }),
  .A2({ S25957[646] }),
  .A3({ S5593 }),
  .ZN({ S5601 })
);
NAND2_X1 #() 
NAND2_X1_5788_ (
  .A1({ S5498 }),
  .A2({ S5497 }),
  .ZN({ S5602 })
);
NOR2_X1 #() 
NOR2_X1_1451_ (
  .A1({ S5504 }),
  .A2({ S5602 }),
  .ZN({ S5603 })
);
NAND2_X1 #() 
NAND2_X1_5789_ (
  .A1({ S5497 }),
  .A2({ S5471 }),
  .ZN({ S5604 })
);
NAND2_X1 #() 
NAND2_X1_5790_ (
  .A1({ S5604 }),
  .A2({ S5485 }),
  .ZN({ S5605 })
);
AOI21_X1 #() 
AOI21_X1_3326_ (
  .A({ S5603 }),
  .B1({ S25957[643] }),
  .B2({ S5605 }),
  .ZN({ S5606 })
);
NAND2_X1 #() 
NAND2_X1_5791_ (
  .A1({ S25957[643] }),
  .A2({ S5496 }),
  .ZN({ S5607 })
);
NOR2_X1 #() 
NOR2_X1_1452_ (
  .A1({ S25957[640] }),
  .A2({ S5544 }),
  .ZN({ S5608 })
);
NAND2_X1 #() 
NAND2_X1_5792_ (
  .A1({ S5608 }),
  .A2({ S0 }),
  .ZN({ S5609 })
);
NAND4_X1 #() 
NAND4_X1_693_ (
  .A1({ S5570 }),
  .A2({ S5609 }),
  .A3({ S25957[644] }),
  .A4({ S5607 }),
  .ZN({ S5610 })
);
OAI21_X1 #() 
OAI21_X1_3016_ (
  .A({ S5610 }),
  .B1({ S5606 }),
  .B2({ S25957[644] }),
  .ZN({ S5611 })
);
OAI21_X1 #() 
OAI21_X1_3017_ (
  .A({ S25957[643] }),
  .B1({ S5588 }),
  .B2({ S5572 }),
  .ZN({ S5612 })
);
NAND3_X1 #() 
NAND3_X1_6261_ (
  .A1({ S5596 }),
  .A2({ S5495 }),
  .A3({ S5612 }),
  .ZN({ S5613 })
);
AOI21_X1 #() 
AOI21_X1_3327_ (
  .A({ S25957[643] }),
  .B1({ S5544 }),
  .B2({ S5475 }),
  .ZN({ S5614 })
);
OAI21_X1 #() 
OAI21_X1_3018_ (
  .A({ S25957[644] }),
  .B1({ S5468 }),
  .B2({ S5614 }),
  .ZN({ S5615 })
);
NAND3_X1 #() 
NAND3_X1_6262_ (
  .A1({ S5613 }),
  .A2({ S5494 }),
  .A3({ S5615 }),
  .ZN({ S5616 })
);
OAI211_X1 #() 
OAI211_X1_2047_ (
  .A({ S5465 }),
  .B({ S5616 }),
  .C1({ S5611 }),
  .C2({ S5494 }),
  .ZN({ S5617 })
);
NAND3_X1 #() 
NAND3_X1_6263_ (
  .A1({ S5617 }),
  .A2({ S5601 }),
  .A3({ S25957[647] }),
  .ZN({ S5618 })
);
NAND4_X1 #() 
NAND4_X1_694_ (
  .A1({ S5503 }),
  .A2({ S0 }),
  .A3({ S5484 }),
  .A4({ S5537 }),
  .ZN({ S5619 })
);
NAND3_X1 #() 
NAND3_X1_6264_ (
  .A1({ S5503 }),
  .A2({ S25957[643] }),
  .A3({ S8 }),
  .ZN({ S5620 })
);
AND3_X1 #() 
AND3_X1_253_ (
  .A1({ S5619 }),
  .A2({ S25957[644] }),
  .A3({ S5620 }),
  .ZN({ S5621 })
);
INV_X1 #() 
INV_X1_1873_ (
  .A({ S5467 }),
  .ZN({ S5622 })
);
NAND2_X1 #() 
NAND2_X1_5793_ (
  .A1({ S5497 }),
  .A2({ S5485 }),
  .ZN({ S5623 })
);
OAI21_X1 #() 
OAI21_X1_3019_ (
  .A({ S5495 }),
  .B1({ S5622 }),
  .B2({ S5623 }),
  .ZN({ S5624 })
);
INV_X1 #() 
INV_X1_1874_ (
  .A({ S5624 }),
  .ZN({ S5625 })
);
OAI21_X1 #() 
OAI21_X1_3020_ (
  .A({ S25957[645] }),
  .B1({ S5625 }),
  .B2({ S5621 }),
  .ZN({ S5626 })
);
NOR2_X1 #() 
NOR2_X1_1453_ (
  .A1({ S5514 }),
  .A2({ S7 }),
  .ZN({ S5627 })
);
OAI211_X1 #() 
OAI211_X1_2048_ (
  .A({ S5589 }),
  .B({ S5495 }),
  .C1({ S25957[643] }),
  .C2({ S5627 }),
  .ZN({ S5629 })
);
OAI21_X1 #() 
OAI21_X1_3021_ (
  .A({ S5591 }),
  .B1({ S25957[643] }),
  .B2({ S5543 }),
  .ZN({ S5630 })
);
NAND3_X1 #() 
NAND3_X1_6265_ (
  .A1({ S5629 }),
  .A2({ S5494 }),
  .A3({ S5630 }),
  .ZN({ S5631 })
);
NAND3_X1 #() 
NAND3_X1_6266_ (
  .A1({ S5631 }),
  .A2({ S5626 }),
  .A3({ S25957[646] }),
  .ZN({ S5632 })
);
OAI21_X1 #() 
OAI21_X1_3022_ (
  .A({ S25957[643] }),
  .B1({ S5602 }),
  .B2({ S5531 }),
  .ZN({ S5633 })
);
NAND3_X1 #() 
NAND3_X1_6267_ (
  .A1({ S5633 }),
  .A2({ S25957[644] }),
  .A3({ S5504 }),
  .ZN({ S5634 })
);
NAND2_X1 #() 
NAND2_X1_5794_ (
  .A1({ S5537 }),
  .A2({ S5544 }),
  .ZN({ S5635 })
);
NAND2_X1 #() 
NAND2_X1_5795_ (
  .A1({ S5559 }),
  .A2({ S5535 }),
  .ZN({ S5636 })
);
OAI211_X1 #() 
OAI211_X1_2049_ (
  .A({ S5636 }),
  .B({ S5495 }),
  .C1({ S0 }),
  .C2({ S5635 }),
  .ZN({ S5637 })
);
NAND3_X1 #() 
NAND3_X1_6268_ (
  .A1({ S5637 }),
  .A2({ S5634 }),
  .A3({ S25957[645] }),
  .ZN({ S5638 })
);
OAI211_X1 #() 
OAI211_X1_2050_ (
  .A({ S5536 }),
  .B({ S25957[644] }),
  .C1({ S25957[643] }),
  .C2({ S5535 }),
  .ZN({ S5640 })
);
NAND3_X1 #() 
NAND3_X1_6269_ (
  .A1({ S5503 }),
  .A2({ S5508 }),
  .A3({ S5512 }),
  .ZN({ S5641 })
);
NAND2_X1 #() 
NAND2_X1_5796_ (
  .A1({ S5641 }),
  .A2({ S25957[643] }),
  .ZN({ S5642 })
);
NAND2_X1 #() 
NAND2_X1_5797_ (
  .A1({ S5642 }),
  .A2({ S5495 }),
  .ZN({ S5643 })
);
NAND3_X1 #() 
NAND3_X1_6270_ (
  .A1({ S5640 }),
  .A2({ S5643 }),
  .A3({ S5494 }),
  .ZN({ S5644 })
);
NAND3_X1 #() 
NAND3_X1_6271_ (
  .A1({ S5638 }),
  .A2({ S5465 }),
  .A3({ S5644 }),
  .ZN({ S5645 })
);
NAND3_X1 #() 
NAND3_X1_6272_ (
  .A1({ S5632 }),
  .A2({ S5645 }),
  .A3({ S5530 }),
  .ZN({ S5646 })
);
NAND2_X1 #() 
NAND2_X1_5798_ (
  .A1({ S5618 }),
  .A2({ S5646 }),
  .ZN({ S5647 })
);
NAND2_X1 #() 
NAND2_X1_5799_ (
  .A1({ S5647 }),
  .A2({ S25957[750] }),
  .ZN({ S5648 })
);
INV_X1 #() 
INV_X1_1875_ (
  .A({ S25957[750] }),
  .ZN({ S5649 })
);
NAND3_X1 #() 
NAND3_X1_6273_ (
  .A1({ S5618 }),
  .A2({ S5649 }),
  .A3({ S5646 }),
  .ZN({ S5650 })
);
NAND2_X1 #() 
NAND2_X1_5800_ (
  .A1({ S5648 }),
  .A2({ S5650 }),
  .ZN({ S25957[622] })
);
NOR2_X1 #() 
NOR2_X1_1454_ (
  .A1({ S25957[622] }),
  .A2({ S25957[718] }),
  .ZN({ S5651 })
);
INV_X1 #() 
INV_X1_1876_ (
  .A({ S25957[718] }),
  .ZN({ S5652 })
);
AOI21_X1 #() 
AOI21_X1_3328_ (
  .A({ S5652 }),
  .B1({ S5648 }),
  .B2({ S5650 }),
  .ZN({ S5653 })
);
OAI21_X1 #() 
OAI21_X1_3023_ (
  .A({ S25957[686] }),
  .B1({ S5651 }),
  .B2({ S5653 }),
  .ZN({ S5654 })
);
INV_X1 #() 
INV_X1_1877_ (
  .A({ S25957[686] }),
  .ZN({ S5655 })
);
NOR2_X1 #() 
NOR2_X1_1455_ (
  .A1({ S5651 }),
  .A2({ S5653 }),
  .ZN({ S25957[590] })
);
NAND2_X1 #() 
NAND2_X1_5801_ (
  .A1({ S25957[590] }),
  .A2({ S5655 }),
  .ZN({ S5656 })
);
NAND2_X1 #() 
NAND2_X1_5802_ (
  .A1({ S5656 }),
  .A2({ S5654 }),
  .ZN({ S25957[558] })
);
NAND2_X1 #() 
NAND2_X1_5803_ (
  .A1({ S25957[558] }),
  .A2({ S4862 }),
  .ZN({ S5658 })
);
NAND3_X1 #() 
NAND3_X1_6274_ (
  .A1({ S5656 }),
  .A2({ S25957[654] }),
  .A3({ S5654 }),
  .ZN({ S5659 })
);
NAND2_X1 #() 
NAND2_X1_5804_ (
  .A1({ S5658 }),
  .A2({ S5659 }),
  .ZN({ S25957[526] })
);
NAND2_X1 #() 
NAND2_X1_5805_ (
  .A1({ S23627 }),
  .A2({ S23628 }),
  .ZN({ S25957[941] })
);
XNOR2_X1 #() 
XNOR2_X1_217_ (
  .A({ S633 }),
  .B({ S25957[941] }),
  .ZN({ S25957[813] })
);
NAND4_X1 #() 
NAND4_X1_695_ (
  .A1({ S5471 }),
  .A2({ S25957[641] }),
  .A3({ S4021 }),
  .A4({ S4018 }),
  .ZN({ S5660 })
);
NAND4_X1 #() 
NAND4_X1_696_ (
  .A1({ S5501 }),
  .A2({ S5660 }),
  .A3({ S5500 }),
  .A4({ S25957[643] }),
  .ZN({ S5661 })
);
NAND2_X1 #() 
NAND2_X1_5806_ (
  .A1({ S5485 }),
  .A2({ S5508 }),
  .ZN({ S5662 })
);
NAND3_X1 #() 
NAND3_X1_6275_ (
  .A1({ S5662 }),
  .A2({ S0 }),
  .A3({ S5475 }),
  .ZN({ S5663 })
);
NAND3_X1 #() 
NAND3_X1_6276_ (
  .A1({ S5661 }),
  .A2({ S5663 }),
  .A3({ S25957[644] }),
  .ZN({ S5664 })
);
NAND3_X1 #() 
NAND3_X1_6277_ (
  .A1({ S5503 }),
  .A2({ S0 }),
  .A3({ S5497 }),
  .ZN({ S5665 })
);
NAND2_X1 #() 
NAND2_X1_5807_ (
  .A1({ S5665 }),
  .A2({ S5480 }),
  .ZN({ S5666 })
);
NAND2_X1 #() 
NAND2_X1_5808_ (
  .A1({ S5666 }),
  .A2({ S5495 }),
  .ZN({ S5667 })
);
AOI21_X1 #() 
AOI21_X1_3329_ (
  .A({ S5494 }),
  .B1({ S5667 }),
  .B2({ S5664 }),
  .ZN({ S5668 })
);
NAND4_X1 #() 
NAND4_X1_697_ (
  .A1({ S5501 }),
  .A2({ S0 }),
  .A3({ S5475 }),
  .A4({ S5508 }),
  .ZN({ S5669 })
);
NAND2_X1 #() 
NAND2_X1_5809_ (
  .A1({ S5475 }),
  .A2({ S5544 }),
  .ZN({ S5670 })
);
NAND2_X1 #() 
NAND2_X1_5810_ (
  .A1({ S5670 }),
  .A2({ S25957[643] }),
  .ZN({ S5671 })
);
NAND3_X1 #() 
NAND3_X1_6278_ (
  .A1({ S5671 }),
  .A2({ S25957[644] }),
  .A3({ S5669 }),
  .ZN({ S5672 })
);
AOI21_X1 #() 
AOI21_X1_3330_ (
  .A({ S0 }),
  .B1({ S5501 }),
  .B2({ S5475 }),
  .ZN({ S5673 })
);
AOI21_X1 #() 
AOI21_X1_3331_ (
  .A({ S25957[643] }),
  .B1({ S5604 }),
  .B2({ S5484 }),
  .ZN({ S5674 })
);
OAI21_X1 #() 
OAI21_X1_3024_ (
  .A({ S5495 }),
  .B1({ S5674 }),
  .B2({ S5673 }),
  .ZN({ S5676 })
);
AOI21_X1 #() 
AOI21_X1_3332_ (
  .A({ S25957[645] }),
  .B1({ S5676 }),
  .B2({ S5672 }),
  .ZN({ S5677 })
);
OAI21_X1 #() 
OAI21_X1_3025_ (
  .A({ S25957[646] }),
  .B1({ S5677 }),
  .B2({ S5668 }),
  .ZN({ S5678 })
);
AND3_X1 #() 
AND3_X1_254_ (
  .A1({ S5548 }),
  .A2({ S5535 }),
  .A3({ S25957[643] }),
  .ZN({ S5679 })
);
NAND4_X1 #() 
NAND4_X1_698_ (
  .A1({ S5498 }),
  .A2({ S0 }),
  .A3({ S5475 }),
  .A4({ S5497 }),
  .ZN({ S5680 })
);
NAND2_X1 #() 
NAND2_X1_5811_ (
  .A1({ S5680 }),
  .A2({ S25957[644] }),
  .ZN({ S5681 })
);
NAND2_X1 #() 
NAND2_X1_5812_ (
  .A1({ S0 }),
  .A2({ S7 }),
  .ZN({ S5682 })
);
OAI22_X1 #() 
OAI22_X1_153_ (
  .A1({ S5682 }),
  .A2({ S5471 }),
  .B1({ S0 }),
  .B2({ S5498 }),
  .ZN({ S5683 })
);
AOI21_X1 #() 
AOI21_X1_3333_ (
  .A({ S25957[645] }),
  .B1({ S5683 }),
  .B2({ S5495 }),
  .ZN({ S5684 })
);
OAI21_X1 #() 
OAI21_X1_3026_ (
  .A({ S5684 }),
  .B1({ S5679 }),
  .B2({ S5681 }),
  .ZN({ S5685 })
);
AOI21_X1 #() 
AOI21_X1_3334_ (
  .A({ S25957[642] }),
  .B1({ S3926 }),
  .B2({ S3929 }),
  .ZN({ S5687 })
);
NOR2_X1 #() 
NOR2_X1_1456_ (
  .A1({ S5687 }),
  .A2({ S5472 }),
  .ZN({ S5688 })
);
NAND2_X1 #() 
NAND2_X1_5813_ (
  .A1({ S5475 }),
  .A2({ S5508 }),
  .ZN({ S5689 })
);
OAI211_X1 #() 
OAI211_X1_2051_ (
  .A({ S5609 }),
  .B({ S25957[644] }),
  .C1({ S5689 }),
  .C2({ S0 }),
  .ZN({ S5690 })
);
OAI211_X1 #() 
OAI211_X1_2052_ (
  .A({ S5690 }),
  .B({ S25957[645] }),
  .C1({ S5624 }),
  .C2({ S5688 }),
  .ZN({ S5691 })
);
NAND3_X1 #() 
NAND3_X1_6279_ (
  .A1({ S5685 }),
  .A2({ S5465 }),
  .A3({ S5691 }),
  .ZN({ S5692 })
);
NAND2_X1 #() 
NAND2_X1_5814_ (
  .A1({ S5692 }),
  .A2({ S5678 }),
  .ZN({ S5693 })
);
NAND2_X1 #() 
NAND2_X1_5815_ (
  .A1({ S5693 }),
  .A2({ S5530 }),
  .ZN({ S5694 })
);
NAND2_X1 #() 
NAND2_X1_5816_ (
  .A1({ S5543 }),
  .A2({ S25957[643] }),
  .ZN({ S5695 })
);
NAND3_X1 #() 
NAND3_X1_6280_ (
  .A1({ S5545 }),
  .A2({ S0 }),
  .A3({ S5537 }),
  .ZN({ S5696 })
);
NAND3_X1 #() 
NAND3_X1_6281_ (
  .A1({ S5695 }),
  .A2({ S25957[644] }),
  .A3({ S5696 }),
  .ZN({ S5698 })
);
NAND3_X1 #() 
NAND3_X1_6282_ (
  .A1({ S5488 }),
  .A2({ S25957[643] }),
  .A3({ S5485 }),
  .ZN({ S5699 })
);
NAND3_X1 #() 
NAND3_X1_6283_ (
  .A1({ S5586 }),
  .A2({ S5565 }),
  .A3({ S5699 }),
  .ZN({ S5700 })
);
NAND3_X1 #() 
NAND3_X1_6284_ (
  .A1({ S5700 }),
  .A2({ S25957[645] }),
  .A3({ S5698 }),
  .ZN({ S5701 })
);
NAND3_X1 #() 
NAND3_X1_6285_ (
  .A1({ S5589 }),
  .A2({ S5495 }),
  .A3({ S5570 }),
  .ZN({ S5702 })
);
NAND2_X1 #() 
NAND2_X1_5817_ (
  .A1({ S5604 }),
  .A2({ S25957[643] }),
  .ZN({ S5703 })
);
NAND2_X1 #() 
NAND2_X1_5818_ (
  .A1({ S5497 }),
  .A2({ S25957[642] }),
  .ZN({ S5704 })
);
INV_X1 #() 
INV_X1_1878_ (
  .A({ S5704 }),
  .ZN({ S5705 })
);
NAND2_X1 #() 
NAND2_X1_5819_ (
  .A1({ S5705 }),
  .A2({ S0 }),
  .ZN({ S5706 })
);
NAND3_X1 #() 
NAND3_X1_6286_ (
  .A1({ S5706 }),
  .A2({ S25957[644] }),
  .A3({ S5703 }),
  .ZN({ S5707 })
);
NAND3_X1 #() 
NAND3_X1_6287_ (
  .A1({ S5702 }),
  .A2({ S5707 }),
  .A3({ S5494 }),
  .ZN({ S5709 })
);
NAND3_X1 #() 
NAND3_X1_6288_ (
  .A1({ S5709 }),
  .A2({ S25957[646] }),
  .A3({ S5701 }),
  .ZN({ S5710 })
);
NAND4_X1 #() 
NAND4_X1_699_ (
  .A1({ S5488 }),
  .A2({ S25957[643] }),
  .A3({ S5471 }),
  .A4({ S8 }),
  .ZN({ S5711 })
);
AOI21_X1 #() 
AOI21_X1_3335_ (
  .A({ S25957[641] }),
  .B1({ S25957[640] }),
  .B2({ S5471 }),
  .ZN({ S5712 })
);
AOI21_X1 #() 
AOI21_X1_3336_ (
  .A({ S5495 }),
  .B1({ S5712 }),
  .B2({ S0 }),
  .ZN({ S5713 })
);
NAND4_X1 #() 
NAND4_X1_700_ (
  .A1({ S5471 }),
  .A2({ S5464 }),
  .A3({ S4021 }),
  .A4({ S4018 }),
  .ZN({ S5714 })
);
OAI211_X1 #() 
OAI211_X1_2053_ (
  .A({ S25957[643] }),
  .B({ S5714 }),
  .C1({ S5514 }),
  .C2({ S7 }),
  .ZN({ S5715 })
);
AOI22_X1 #() 
AOI22_X1_652_ (
  .A1({ S5687 }),
  .A2({ S7 }),
  .B1({ S3849 }),
  .B2({ S3846 }),
  .ZN({ S5716 })
);
AOI22_X1 #() 
AOI22_X1_653_ (
  .A1({ S5713 }),
  .A2({ S5711 }),
  .B1({ S5715 }),
  .B2({ S5716 }),
  .ZN({ S5717 })
);
INV_X1 #() 
INV_X1_1879_ (
  .A({ S5484 }),
  .ZN({ S5718 })
);
OAI21_X1 #() 
OAI21_X1_3027_ (
  .A({ S0 }),
  .B1({ S5718 }),
  .B2({ S5524 }),
  .ZN({ S5720 })
);
OAI211_X1 #() 
OAI211_X1_2054_ (
  .A({ S5720 }),
  .B({ S25957[644] }),
  .C1({ S0 }),
  .C2({ S5554 }),
  .ZN({ S5721 })
);
AOI22_X1 #() 
AOI22_X1_654_ (
  .A1({ S3926 }),
  .A2({ S3929 }),
  .B1({ S5471 }),
  .B2({ S5464 }),
  .ZN({ S5722 })
);
NAND2_X1 #() 
NAND2_X1_5820_ (
  .A1({ S5722 }),
  .A2({ S5497 }),
  .ZN({ S5723 })
);
AOI22_X1 #() 
AOI22_X1_655_ (
  .A1({ S25957[643] }),
  .A2({ S5464 }),
  .B1({ S3849 }),
  .B2({ S3846 }),
  .ZN({ S5724 })
);
AOI21_X1 #() 
AOI21_X1_3337_ (
  .A({ S5494 }),
  .B1({ S5723 }),
  .B2({ S5724 }),
  .ZN({ S5725 })
);
NAND2_X1 #() 
NAND2_X1_5821_ (
  .A1({ S5721 }),
  .A2({ S5725 }),
  .ZN({ S5726 })
);
OAI211_X1 #() 
OAI211_X1_2055_ (
  .A({ S5465 }),
  .B({ S5726 }),
  .C1({ S25957[645] }),
  .C2({ S5717 }),
  .ZN({ S5727 })
);
NAND3_X1 #() 
NAND3_X1_6289_ (
  .A1({ S5727 }),
  .A2({ S5710 }),
  .A3({ S25957[647] }),
  .ZN({ S5728 })
);
NAND3_X1 #() 
NAND3_X1_6290_ (
  .A1({ S5694 }),
  .A2({ S25957[749] }),
  .A3({ S5728 }),
  .ZN({ S5729 })
);
INV_X1 #() 
INV_X1_1880_ (
  .A({ S25957[749] }),
  .ZN({ S5731 })
);
AOI21_X1 #() 
AOI21_X1_3338_ (
  .A({ S25957[647] }),
  .B1({ S5692 }),
  .B2({ S5678 }),
  .ZN({ S5732 })
);
INV_X1 #() 
INV_X1_1881_ (
  .A({ S5728 }),
  .ZN({ S5733 })
);
OAI21_X1 #() 
OAI21_X1_3028_ (
  .A({ S5731 }),
  .B1({ S5733 }),
  .B2({ S5732 }),
  .ZN({ S5734 })
);
NAND3_X1 #() 
NAND3_X1_6291_ (
  .A1({ S5734 }),
  .A2({ S5729 }),
  .A3({ S25957[813] }),
  .ZN({ S5735 })
);
INV_X1 #() 
INV_X1_1882_ (
  .A({ S25957[813] }),
  .ZN({ S5736 })
);
NAND3_X1 #() 
NAND3_X1_6292_ (
  .A1({ S5694 }),
  .A2({ S5731 }),
  .A3({ S5728 }),
  .ZN({ S5737 })
);
OAI21_X1 #() 
OAI21_X1_3029_ (
  .A({ S25957[749] }),
  .B1({ S5733 }),
  .B2({ S5732 }),
  .ZN({ S5738 })
);
NAND3_X1 #() 
NAND3_X1_6293_ (
  .A1({ S5738 }),
  .A2({ S5737 }),
  .A3({ S5736 }),
  .ZN({ S5739 })
);
NAND3_X1 #() 
NAND3_X1_6294_ (
  .A1({ S5735 }),
  .A2({ S5739 }),
  .A3({ S25957[653] }),
  .ZN({ S5740 })
);
NAND3_X1 #() 
NAND3_X1_6295_ (
  .A1({ S5738 }),
  .A2({ S5737 }),
  .A3({ S25957[813] }),
  .ZN({ S5742 })
);
NAND3_X1 #() 
NAND3_X1_6296_ (
  .A1({ S5734 }),
  .A2({ S5729 }),
  .A3({ S5736 }),
  .ZN({ S5743 })
);
NAND3_X1 #() 
NAND3_X1_6297_ (
  .A1({ S5742 }),
  .A2({ S5743 }),
  .A3({ S4798 }),
  .ZN({ S5744 })
);
AND2_X1 #() 
AND2_X1_364_ (
  .A1({ S5744 }),
  .A2({ S5740 }),
  .ZN({ S25957[525] })
);
NOR2_X1 #() 
NOR2_X1_1457_ (
  .A1({ S3206 }),
  .A2({ S3204 }),
  .ZN({ S5745 })
);
XNOR2_X1 #() 
XNOR2_X1_218_ (
  .A({ S5745 }),
  .B({ S25957[812] }),
  .ZN({ S25957[684] })
);
INV_X1 #() 
INV_X1_1883_ (
  .A({ S25957[812] }),
  .ZN({ S5746 })
);
NAND2_X1 #() 
NAND2_X1_5822_ (
  .A1({ S3203 }),
  .A2({ S3175 }),
  .ZN({ S5747 })
);
XOR2_X1 #() 
XOR2_X1_101_ (
  .A({ S5747 }),
  .B({ S25957[876] }),
  .Z({ S25957[748] })
);
OAI22_X1 #() 
OAI22_X1_154_ (
  .A1({ S5604 }),
  .A2({ S5524 }),
  .B1({ S7 }),
  .B2({ S5471 }),
  .ZN({ S5748 })
);
NAND2_X1 #() 
NAND2_X1_5823_ (
  .A1({ S5748 }),
  .A2({ S0 }),
  .ZN({ S5750 })
);
NAND2_X1 #() 
NAND2_X1_5824_ (
  .A1({ S5520 }),
  .A2({ S5545 }),
  .ZN({ S5751 })
);
NAND3_X1 #() 
NAND3_X1_6298_ (
  .A1({ S5750 }),
  .A2({ S5495 }),
  .A3({ S5751 }),
  .ZN({ S5752 })
);
OAI21_X1 #() 
OAI21_X1_3030_ (
  .A({ S5660 }),
  .B1({ S5687 }),
  .B2({ S5498 }),
  .ZN({ S5753 })
);
AOI21_X1 #() 
AOI21_X1_3339_ (
  .A({ S5494 }),
  .B1({ S5753 }),
  .B2({ S25957[644] }),
  .ZN({ S5754 })
);
NAND2_X1 #() 
NAND2_X1_5825_ (
  .A1({ S5752 }),
  .A2({ S5754 }),
  .ZN({ S5755 })
);
OAI21_X1 #() 
OAI21_X1_3031_ (
  .A({ S0 }),
  .B1({ S5510 }),
  .B2({ S5472 }),
  .ZN({ S5756 })
);
OAI211_X1 #() 
OAI211_X1_2056_ (
  .A({ S5756 }),
  .B({ S25957[644] }),
  .C1({ S5635 }),
  .C2({ S5553 }),
  .ZN({ S5757 })
);
NAND2_X1 #() 
NAND2_X1_5826_ (
  .A1({ S5641 }),
  .A2({ S0 }),
  .ZN({ S5758 })
);
AOI21_X1 #() 
AOI21_X1_3340_ (
  .A({ S25957[641] }),
  .B1({ S3930 }),
  .B2({ S3931 }),
  .ZN({ S5759 })
);
AOI21_X1 #() 
AOI21_X1_3341_ (
  .A({ S25957[644] }),
  .B1({ S5565 }),
  .B2({ S5759 }),
  .ZN({ S5761 })
);
AOI21_X1 #() 
AOI21_X1_3342_ (
  .A({ S25957[645] }),
  .B1({ S5761 }),
  .B2({ S5758 }),
  .ZN({ S5762 })
);
NAND2_X1 #() 
NAND2_X1_5827_ (
  .A1({ S5757 }),
  .A2({ S5762 }),
  .ZN({ S5763 })
);
NAND3_X1 #() 
NAND3_X1_6299_ (
  .A1({ S5763 }),
  .A2({ S5755 }),
  .A3({ S5465 }),
  .ZN({ S5764 })
);
AOI21_X1 #() 
AOI21_X1_3343_ (
  .A({ S0 }),
  .B1({ S5544 }),
  .B2({ S5475 }),
  .ZN({ S5765 })
);
AND2_X1 #() 
AND2_X1_365_ (
  .A1({ S0 }),
  .A2({ S5500 }),
  .ZN({ S5766 })
);
OAI21_X1 #() 
OAI21_X1_3032_ (
  .A({ S25957[644] }),
  .B1({ S5765 }),
  .B2({ S5766 }),
  .ZN({ S5767 })
);
NAND3_X1 #() 
NAND3_X1_6300_ (
  .A1({ S0 }),
  .A2({ S5479 }),
  .A3({ S5544 }),
  .ZN({ S5768 })
);
NAND2_X1 #() 
NAND2_X1_5828_ (
  .A1({ S5566 }),
  .A2({ S5768 }),
  .ZN({ S5769 })
);
NAND2_X1 #() 
NAND2_X1_5829_ (
  .A1({ S5769 }),
  .A2({ S5495 }),
  .ZN({ S5770 })
);
AND3_X1 #() 
AND3_X1_255_ (
  .A1({ S5770 }),
  .A2({ S5767 }),
  .A3({ S25957[645] }),
  .ZN({ S5772 })
);
INV_X1 #() 
INV_X1_1884_ (
  .A({ S5722 }),
  .ZN({ S5773 })
);
OAI211_X1 #() 
OAI211_X1_2057_ (
  .A({ S5561 }),
  .B({ S5495 }),
  .C1({ S5773 }),
  .C2({ S5718 }),
  .ZN({ S5774 })
);
OAI211_X1 #() 
OAI211_X1_2058_ (
  .A({ S5723 }),
  .B({ S25957[644] }),
  .C1({ S5588 }),
  .C2({ S5466 }),
  .ZN({ S5775 })
);
AOI21_X1 #() 
AOI21_X1_3344_ (
  .A({ S25957[645] }),
  .B1({ S5775 }),
  .B2({ S5774 }),
  .ZN({ S5776 })
);
OAI21_X1 #() 
OAI21_X1_3033_ (
  .A({ S25957[646] }),
  .B1({ S5772 }),
  .B2({ S5776 }),
  .ZN({ S5777 })
);
NAND3_X1 #() 
NAND3_X1_6301_ (
  .A1({ S5764 }),
  .A2({ S5777 }),
  .A3({ S25957[647] }),
  .ZN({ S5778 })
);
OAI21_X1 #() 
OAI21_X1_3034_ (
  .A({ S25957[643] }),
  .B1({ S5472 }),
  .B2({ S5464 }),
  .ZN({ S5779 })
);
NAND2_X1 #() 
NAND2_X1_5830_ (
  .A1({ S5722 }),
  .A2({ S5514 }),
  .ZN({ S5780 })
);
AOI21_X1 #() 
AOI21_X1_3345_ (
  .A({ S5495 }),
  .B1({ S5779 }),
  .B2({ S5780 }),
  .ZN({ S5781 })
);
NAND3_X1 #() 
NAND3_X1_6302_ (
  .A1({ S3926 }),
  .A2({ S3929 }),
  .A3({ S25957[642] }),
  .ZN({ S5783 })
);
NAND2_X1 #() 
NAND2_X1_5831_ (
  .A1({ S5594 }),
  .A2({ S5783 }),
  .ZN({ S5784 })
);
AND2_X1 #() 
AND2_X1_366_ (
  .A1({ S5716 }),
  .A2({ S5784 }),
  .ZN({ S5785 })
);
OAI21_X1 #() 
OAI21_X1_3035_ (
  .A({ S5494 }),
  .B1({ S5785 }),
  .B2({ S5781 }),
  .ZN({ S5786 })
);
AOI21_X1 #() 
AOI21_X1_3346_ (
  .A({ S25957[643] }),
  .B1({ S5489 }),
  .B2({ S5704 }),
  .ZN({ S5787 })
);
NAND4_X1 #() 
NAND4_X1_701_ (
  .A1({ S5503 }),
  .A2({ S25957[643] }),
  .A3({ S5484 }),
  .A4({ S5537 }),
  .ZN({ S5788 })
);
NAND2_X1 #() 
NAND2_X1_5832_ (
  .A1({ S5788 }),
  .A2({ S5495 }),
  .ZN({ S5789 })
);
NAND2_X1 #() 
NAND2_X1_5833_ (
  .A1({ S5471 }),
  .A2({ S137 }),
  .ZN({ S5790 })
);
NAND2_X1 #() 
NAND2_X1_5834_ (
  .A1({ S25957[644] }),
  .A2({ S5790 }),
  .ZN({ S5791 })
);
OAI211_X1 #() 
OAI211_X1_2059_ (
  .A({ S25957[645] }),
  .B({ S5791 }),
  .C1({ S5787 }),
  .C2({ S5789 }),
  .ZN({ S5792 })
);
NAND3_X1 #() 
NAND3_X1_6303_ (
  .A1({ S5786 }),
  .A2({ S25957[646] }),
  .A3({ S5792 }),
  .ZN({ S5794 })
);
AOI21_X1 #() 
AOI21_X1_3347_ (
  .A({ S25957[644] }),
  .B1({ S5711 }),
  .B2({ S5682 }),
  .ZN({ S5795 })
);
NAND2_X1 #() 
NAND2_X1_5835_ (
  .A1({ S5704 }),
  .A2({ S0 }),
  .ZN({ S5796 })
);
AOI21_X1 #() 
AOI21_X1_3348_ (
  .A({ S5495 }),
  .B1({ S5536 }),
  .B2({ S5796 }),
  .ZN({ S5797 })
);
OAI21_X1 #() 
OAI21_X1_3036_ (
  .A({ S25957[645] }),
  .B1({ S5797 }),
  .B2({ S5795 }),
  .ZN({ S5798 })
);
NAND3_X1 #() 
NAND3_X1_6304_ (
  .A1({ S5565 }),
  .A2({ S25957[643] }),
  .A3({ S8 }),
  .ZN({ S5799 })
);
NAND3_X1 #() 
NAND3_X1_6305_ (
  .A1({ S5525 }),
  .A2({ S0 }),
  .A3({ S5500 }),
  .ZN({ S5800 })
);
AOI21_X1 #() 
AOI21_X1_3349_ (
  .A({ S25957[644] }),
  .B1({ S5800 }),
  .B2({ S5799 }),
  .ZN({ S5801 })
);
NAND2_X1 #() 
NAND2_X1_5836_ (
  .A1({ S5497 }),
  .A2({ S5508 }),
  .ZN({ S5802 })
);
NAND2_X1 #() 
NAND2_X1_5837_ (
  .A1({ S5802 }),
  .A2({ S0 }),
  .ZN({ S5803 })
);
AOI21_X1 #() 
AOI21_X1_3350_ (
  .A({ S5495 }),
  .B1({ S5509 }),
  .B2({ S5803 }),
  .ZN({ S5805 })
);
OAI21_X1 #() 
OAI21_X1_3037_ (
  .A({ S5494 }),
  .B1({ S5801 }),
  .B2({ S5805 }),
  .ZN({ S5806 })
);
NAND3_X1 #() 
NAND3_X1_6306_ (
  .A1({ S5798 }),
  .A2({ S5806 }),
  .A3({ S5465 }),
  .ZN({ S5807 })
);
NAND3_X1 #() 
NAND3_X1_6307_ (
  .A1({ S5794 }),
  .A2({ S5807 }),
  .A3({ S5530 }),
  .ZN({ S5808 })
);
NAND3_X1 #() 
NAND3_X1_6308_ (
  .A1({ S5778 }),
  .A2({ S5808 }),
  .A3({ S25957[748] }),
  .ZN({ S5809 })
);
INV_X1 #() 
INV_X1_1885_ (
  .A({ S25957[748] }),
  .ZN({ S5810 })
);
NAND2_X1 #() 
NAND2_X1_5838_ (
  .A1({ S5779 }),
  .A2({ S5780 }),
  .ZN({ S5811 })
);
NAND2_X1 #() 
NAND2_X1_5839_ (
  .A1({ S5811 }),
  .A2({ S25957[644] }),
  .ZN({ S5812 })
);
AOI21_X1 #() 
AOI21_X1_3351_ (
  .A({ S25957[645] }),
  .B1({ S5716 }),
  .B2({ S5784 }),
  .ZN({ S5813 })
);
NAND2_X1 #() 
NAND2_X1_5840_ (
  .A1({ S5812 }),
  .A2({ S5813 }),
  .ZN({ S5814 })
);
OAI21_X1 #() 
OAI21_X1_3038_ (
  .A({ S0 }),
  .B1({ S5499 }),
  .B2({ S5705 }),
  .ZN({ S5816 })
);
NOR2_X1 #() 
NOR2_X1_1458_ (
  .A1({ S5673 }),
  .A2({ S25957[644] }),
  .ZN({ S5817 })
);
AOI22_X1 #() 
AOI22_X1_656_ (
  .A1({ S5816 }),
  .A2({ S5817 }),
  .B1({ S25957[644] }),
  .B2({ S5790 }),
  .ZN({ S5818 })
);
OAI211_X1 #() 
OAI211_X1_2060_ (
  .A({ S5814 }),
  .B({ S25957[646] }),
  .C1({ S5818 }),
  .C2({ S5494 }),
  .ZN({ S5819 })
);
OR2_X1 #() 
OR2_X1_76_ (
  .A1({ S5801 }),
  .A2({ S5805 }),
  .ZN({ S5820 })
);
NAND2_X1 #() 
NAND2_X1_5841_ (
  .A1({ S5711 }),
  .A2({ S5682 }),
  .ZN({ S5821 })
);
NAND2_X1 #() 
NAND2_X1_5842_ (
  .A1({ S5821 }),
  .A2({ S5495 }),
  .ZN({ S5822 })
);
OAI211_X1 #() 
OAI211_X1_2061_ (
  .A({ S5706 }),
  .B({ S25957[644] }),
  .C1({ S5670 }),
  .C2({ S5585 }),
  .ZN({ S5823 })
);
NAND3_X1 #() 
NAND3_X1_6309_ (
  .A1({ S5823 }),
  .A2({ S5822 }),
  .A3({ S25957[645] }),
  .ZN({ S5824 })
);
OAI211_X1 #() 
OAI211_X1_2062_ (
  .A({ S5824 }),
  .B({ S5465 }),
  .C1({ S5820 }),
  .C2({ S25957[645] }),
  .ZN({ S5825 })
);
NAND3_X1 #() 
NAND3_X1_6310_ (
  .A1({ S5825 }),
  .A2({ S5819 }),
  .A3({ S5530 }),
  .ZN({ S5827 })
);
AOI22_X1 #() 
AOI22_X1_657_ (
  .A1({ S5762 }),
  .A2({ S5757 }),
  .B1({ S5752 }),
  .B2({ S5754 }),
  .ZN({ S5828 })
);
NAND3_X1 #() 
NAND3_X1_6311_ (
  .A1({ S5770 }),
  .A2({ S5767 }),
  .A3({ S25957[645] }),
  .ZN({ S5829 })
);
NAND2_X1 #() 
NAND2_X1_5843_ (
  .A1({ S5775 }),
  .A2({ S5774 }),
  .ZN({ S5830 })
);
NAND2_X1 #() 
NAND2_X1_5844_ (
  .A1({ S5830 }),
  .A2({ S5494 }),
  .ZN({ S5831 })
);
NAND3_X1 #() 
NAND3_X1_6312_ (
  .A1({ S5831 }),
  .A2({ S5829 }),
  .A3({ S25957[646] }),
  .ZN({ S5832 })
);
OAI211_X1 #() 
OAI211_X1_2063_ (
  .A({ S5832 }),
  .B({ S25957[647] }),
  .C1({ S5828 }),
  .C2({ S25957[646] }),
  .ZN({ S5833 })
);
NAND3_X1 #() 
NAND3_X1_6313_ (
  .A1({ S5833 }),
  .A2({ S5827 }),
  .A3({ S5810 }),
  .ZN({ S5834 })
);
NAND3_X1 #() 
NAND3_X1_6314_ (
  .A1({ S5834 }),
  .A2({ S5809 }),
  .A3({ S5746 }),
  .ZN({ S5835 })
);
NAND3_X1 #() 
NAND3_X1_6315_ (
  .A1({ S5778 }),
  .A2({ S5808 }),
  .A3({ S5810 }),
  .ZN({ S5836 })
);
NAND3_X1 #() 
NAND3_X1_6316_ (
  .A1({ S5833 }),
  .A2({ S5827 }),
  .A3({ S25957[748] }),
  .ZN({ S5838 })
);
NAND3_X1 #() 
NAND3_X1_6317_ (
  .A1({ S5838 }),
  .A2({ S5836 }),
  .A3({ S25957[812] }),
  .ZN({ S5839 })
);
AOI21_X1 #() 
AOI21_X1_3352_ (
  .A({ S4803 }),
  .B1({ S5835 }),
  .B2({ S5839 }),
  .ZN({ S5840 })
);
AND3_X1 #() 
AND3_X1_256_ (
  .A1({ S5839 }),
  .A2({ S5835 }),
  .A3({ S4803 }),
  .ZN({ S5841 })
);
NOR2_X1 #() 
NOR2_X1_1459_ (
  .A1({ S5841 }),
  .A2({ S5840 }),
  .ZN({ S25957[524] })
);
NAND2_X1 #() 
NAND2_X1_5845_ (
  .A1({ S786 }),
  .A2({ S785 }),
  .ZN({ S25957[875] })
);
XNOR2_X1 #() 
XNOR2_X1_219_ (
  .A({ S25957[875] }),
  .B({ S3210 }),
  .ZN({ S25957[843] })
);
INV_X1 #() 
INV_X1_1886_ (
  .A({ S25957[843] }),
  .ZN({ S5842 })
);
OAI221_X1 #() 
OAI221_X1_170_ (
  .A({ S25957[645] }),
  .B1({ S5602 }),
  .B2({ S5594 }),
  .C1({ S5486 }),
  .C2({ S5703 }),
  .ZN({ S5843 })
);
NAND3_X1 #() 
NAND3_X1_6318_ (
  .A1({ S5783 }),
  .A2({ S5503 }),
  .A3({ S8 }),
  .ZN({ S5844 })
);
AOI21_X1 #() 
AOI21_X1_3353_ (
  .A({ S25957[644] }),
  .B1({ S5844 }),
  .B2({ S5494 }),
  .ZN({ S5846 })
);
NAND3_X1 #() 
NAND3_X1_6319_ (
  .A1({ S5548 }),
  .A2({ S0 }),
  .A3({ S5535 }),
  .ZN({ S5847 })
);
NAND3_X1 #() 
NAND3_X1_6320_ (
  .A1({ S5847 }),
  .A2({ S5494 }),
  .A3({ S5699 }),
  .ZN({ S5848 })
);
OAI21_X1 #() 
OAI21_X1_3039_ (
  .A({ S5799 }),
  .B1({ S5532 }),
  .B2({ S5524 }),
  .ZN({ S5849 })
);
AOI21_X1 #() 
AOI21_X1_3354_ (
  .A({ S5495 }),
  .B1({ S5849 }),
  .B2({ S25957[645] }),
  .ZN({ S5850 })
);
AOI22_X1 #() 
AOI22_X1_658_ (
  .A1({ S5850 }),
  .A2({ S5848 }),
  .B1({ S5843 }),
  .B2({ S5846 }),
  .ZN({ S5851 })
);
NAND3_X1 #() 
NAND3_X1_6321_ (
  .A1({ S5503 }),
  .A2({ S0 }),
  .A3({ S8 }),
  .ZN({ S5852 })
);
NAND4_X1 #() 
NAND4_X1_702_ (
  .A1({ S5498 }),
  .A2({ S25957[643] }),
  .A3({ S5497 }),
  .A4({ S25957[642] }),
  .ZN({ S5853 })
);
NAND3_X1 #() 
NAND3_X1_6322_ (
  .A1({ S5853 }),
  .A2({ S5852 }),
  .A3({ S5492 }),
  .ZN({ S5854 })
);
NAND2_X1 #() 
NAND2_X1_5846_ (
  .A1({ S5854 }),
  .A2({ S5495 }),
  .ZN({ S5855 })
);
NAND3_X1 #() 
NAND3_X1_6323_ (
  .A1({ S5573 }),
  .A2({ S25957[643] }),
  .A3({ S5714 }),
  .ZN({ S5857 })
);
AOI21_X1 #() 
AOI21_X1_3355_ (
  .A({ S5495 }),
  .B1({ S5722 }),
  .B2({ S5484 }),
  .ZN({ S5858 })
);
AOI21_X1 #() 
AOI21_X1_3356_ (
  .A({ S25957[645] }),
  .B1({ S5858 }),
  .B2({ S5857 }),
  .ZN({ S5859 })
);
NAND2_X1 #() 
NAND2_X1_5847_ (
  .A1({ S5855 }),
  .A2({ S5859 }),
  .ZN({ S5860 })
);
OAI21_X1 #() 
OAI21_X1_3040_ (
  .A({ S0 }),
  .B1({ S5588 }),
  .B2({ S5486 }),
  .ZN({ S5861 })
);
AND2_X1 #() 
AND2_X1_367_ (
  .A1({ S25957[643] }),
  .A2({ S5500 }),
  .ZN({ S5862 })
);
NAND2_X1 #() 
NAND2_X1_5848_ (
  .A1({ S5862 }),
  .A2({ S5489 }),
  .ZN({ S5863 })
);
NAND3_X1 #() 
NAND3_X1_6324_ (
  .A1({ S5863 }),
  .A2({ S5861 }),
  .A3({ S25957[644] }),
  .ZN({ S5864 })
);
NAND3_X1 #() 
NAND3_X1_6325_ (
  .A1({ S5623 }),
  .A2({ S25957[643] }),
  .A3({ S5484 }),
  .ZN({ S5865 })
);
OAI211_X1 #() 
OAI211_X1_2064_ (
  .A({ S5865 }),
  .B({ S5495 }),
  .C1({ S5627 }),
  .C2({ S5773 }),
  .ZN({ S5866 })
);
NAND3_X1 #() 
NAND3_X1_6326_ (
  .A1({ S5864 }),
  .A2({ S25957[645] }),
  .A3({ S5866 }),
  .ZN({ S5868 })
);
NAND3_X1 #() 
NAND3_X1_6327_ (
  .A1({ S5868 }),
  .A2({ S5860 }),
  .A3({ S5465 }),
  .ZN({ S5869 })
);
OAI211_X1 #() 
OAI211_X1_2065_ (
  .A({ S5869 }),
  .B({ S25957[647] }),
  .C1({ S5851 }),
  .C2({ S5465 }),
  .ZN({ S5870 })
);
NOR2_X1 #() 
NOR2_X1_1460_ (
  .A1({ S5554 }),
  .A2({ S25957[643] }),
  .ZN({ S5871 })
);
NAND2_X1 #() 
NAND2_X1_5849_ (
  .A1({ S5509 }),
  .A2({ S5495 }),
  .ZN({ S5872 })
);
AOI22_X1 #() 
AOI22_X1_659_ (
  .A1({ S5508 }),
  .A2({ S25957[640] }),
  .B1({ S3926 }),
  .B2({ S3929 }),
  .ZN({ S5873 })
);
OR2_X1 #() 
OR2_X1_77_ (
  .A1({ S5873 }),
  .A2({ S5495 }),
  .ZN({ S5874 })
);
OAI211_X1 #() 
OAI211_X1_2066_ (
  .A({ S5874 }),
  .B({ S5494 }),
  .C1({ S5872 }),
  .C2({ S5871 }),
  .ZN({ S5875 })
);
AND3_X1 #() 
AND3_X1_257_ (
  .A1({ S5589 }),
  .A2({ S5574 }),
  .A3({ S25957[644] }),
  .ZN({ S5876 })
);
NAND3_X1 #() 
NAND3_X1_6328_ (
  .A1({ S25957[643] }),
  .A2({ S5479 }),
  .A3({ S5485 }),
  .ZN({ S5877 })
);
NAND2_X1 #() 
NAND2_X1_5850_ (
  .A1({ S5560 }),
  .A2({ S0 }),
  .ZN({ S5879 })
);
NAND3_X1 #() 
NAND3_X1_6329_ (
  .A1({ S5879 }),
  .A2({ S5495 }),
  .A3({ S5877 }),
  .ZN({ S5880 })
);
NAND2_X1 #() 
NAND2_X1_5851_ (
  .A1({ S5880 }),
  .A2({ S25957[645] }),
  .ZN({ S5881 })
);
OAI21_X1 #() 
OAI21_X1_3041_ (
  .A({ S5875 }),
  .B1({ S5876 }),
  .B2({ S5881 }),
  .ZN({ S5882 })
);
NAND2_X1 #() 
NAND2_X1_5852_ (
  .A1({ S5882 }),
  .A2({ S25957[646] }),
  .ZN({ S5883 })
);
AOI21_X1 #() 
AOI21_X1_3357_ (
  .A({ S0 }),
  .B1({ S5515 }),
  .B2({ S5565 }),
  .ZN({ S5884 })
);
OAI21_X1 #() 
OAI21_X1_3042_ (
  .A({ S5495 }),
  .B1({ S5549 }),
  .B2({ S5884 }),
  .ZN({ S5885 })
);
NAND4_X1 #() 
NAND4_X1_703_ (
  .A1({ S5565 }),
  .A2({ S5498 }),
  .A3({ S25957[643] }),
  .A4({ S5497 }),
  .ZN({ S5886 })
);
NAND3_X1 #() 
NAND3_X1_6330_ (
  .A1({ S5636 }),
  .A2({ S25957[644] }),
  .A3({ S5886 }),
  .ZN({ S5887 })
);
NAND3_X1 #() 
NAND3_X1_6331_ (
  .A1({ S5885 }),
  .A2({ S5494 }),
  .A3({ S5887 }),
  .ZN({ S5888 })
);
OAI211_X1 #() 
OAI211_X1_2067_ (
  .A({ S5570 }),
  .B({ S25957[644] }),
  .C1({ S8 }),
  .C2({ S5783 }),
  .ZN({ S5890 })
);
OAI21_X1 #() 
OAI21_X1_3043_ (
  .A({ S5495 }),
  .B1({ S5520 }),
  .B2({ S5545 }),
  .ZN({ S5891 })
);
NAND3_X1 #() 
NAND3_X1_6332_ (
  .A1({ S5890 }),
  .A2({ S25957[645] }),
  .A3({ S5891 }),
  .ZN({ S5892 })
);
NAND3_X1 #() 
NAND3_X1_6333_ (
  .A1({ S5888 }),
  .A2({ S5465 }),
  .A3({ S5892 }),
  .ZN({ S5893 })
);
NAND3_X1 #() 
NAND3_X1_6334_ (
  .A1({ S5893 }),
  .A2({ S5883 }),
  .A3({ S5530 }),
  .ZN({ S5894 })
);
NAND3_X1 #() 
NAND3_X1_6335_ (
  .A1({ S5894 }),
  .A2({ S5870 }),
  .A3({ S5842 }),
  .ZN({ S5895 })
);
INV_X1 #() 
INV_X1_1887_ (
  .A({ S5895 }),
  .ZN({ S5896 })
);
AOI21_X1 #() 
AOI21_X1_3358_ (
  .A({ S5842 }),
  .B1({ S5894 }),
  .B2({ S5870 }),
  .ZN({ S5897 })
);
OAI21_X1 #() 
OAI21_X1_3044_ (
  .A({ S101 }),
  .B1({ S5896 }),
  .B2({ S5897 }),
  .ZN({ S5898 })
);
NAND2_X1 #() 
NAND2_X1_5853_ (
  .A1({ S5894 }),
  .A2({ S5870 }),
  .ZN({ S5899 })
);
NAND2_X1 #() 
NAND2_X1_5854_ (
  .A1({ S5899 }),
  .A2({ S25957[843] }),
  .ZN({ S5901 })
);
NAND3_X1 #() 
NAND3_X1_6336_ (
  .A1({ S5901 }),
  .A2({ S25957[779] }),
  .A3({ S5895 }),
  .ZN({ S5902 })
);
NAND2_X1 #() 
NAND2_X1_5855_ (
  .A1({ S5898 }),
  .A2({ S5902 }),
  .ZN({ S9 })
);
AND2_X1 #() 
AND2_X1_368_ (
  .A1({ S5898 }),
  .A2({ S5902 }),
  .ZN({ S25957[523] })
);
NAND2_X1 #() 
NAND2_X1_5856_ (
  .A1({ S3278 }),
  .A2({ S25957[1064] }),
  .ZN({ S5903 })
);
NAND2_X1 #() 
NAND2_X1_5857_ (
  .A1({ S25957[872] }),
  .A2({ S3276 }),
  .ZN({ S5904 })
);
NAND2_X1 #() 
NAND2_X1_5858_ (
  .A1({ S5904 }),
  .A2({ S5903 }),
  .ZN({ S25957[808] })
);
NAND2_X1 #() 
NAND2_X1_5859_ (
  .A1({ S3348 }),
  .A2({ S3349 }),
  .ZN({ S25957[744] })
);
INV_X1 #() 
INV_X1_1888_ (
  .A({ S25957[744] }),
  .ZN({ S5905 })
);
NAND3_X1 #() 
NAND3_X1_6337_ (
  .A1({ S5548 }),
  .A2({ S25957[643] }),
  .A3({ S5515 }),
  .ZN({ S5906 })
);
AOI21_X1 #() 
AOI21_X1_3359_ (
  .A({ S5495 }),
  .B1({ S5543 }),
  .B2({ S0 }),
  .ZN({ S5908 })
);
AOI22_X1 #() 
AOI22_X1_660_ (
  .A1({ S5906 }),
  .A2({ S5908 }),
  .B1({ S5642 }),
  .B2({ S5476 }),
  .ZN({ S5909 })
);
AOI21_X1 #() 
AOI21_X1_3360_ (
  .A({ S25957[643] }),
  .B1({ S5565 }),
  .B2({ S5464 }),
  .ZN({ S5910 })
);
NAND3_X1 #() 
NAND3_X1_6338_ (
  .A1({ S5605 }),
  .A2({ S25957[644] }),
  .A3({ S5480 }),
  .ZN({ S5911 })
);
OAI211_X1 #() 
OAI211_X1_2068_ (
  .A({ S5911 }),
  .B({ S5494 }),
  .C1({ S5789 }),
  .C2({ S5910 }),
  .ZN({ S5912 })
);
OAI211_X1 #() 
OAI211_X1_2069_ (
  .A({ S5912 }),
  .B({ S25957[646] }),
  .C1({ S5909 }),
  .C2({ S5494 }),
  .ZN({ S5913 })
);
NAND3_X1 #() 
NAND3_X1_6339_ (
  .A1({ S5759 }),
  .A2({ S5484 }),
  .A3({ S5503 }),
  .ZN({ S5914 })
);
NAND2_X1 #() 
NAND2_X1_5860_ (
  .A1({ S5680 }),
  .A2({ S5914 }),
  .ZN({ S5915 })
);
NAND2_X1 #() 
NAND2_X1_5861_ (
  .A1({ S5915 }),
  .A2({ S5495 }),
  .ZN({ S5916 })
);
NAND2_X1 #() 
NAND2_X1_5862_ (
  .A1({ S5665 }),
  .A2({ S5799 }),
  .ZN({ S5917 })
);
AOI21_X1 #() 
AOI21_X1_3361_ (
  .A({ S5494 }),
  .B1({ S5917 }),
  .B2({ S25957[644] }),
  .ZN({ S5919 })
);
NAND2_X1 #() 
NAND2_X1_5863_ (
  .A1({ S0 }),
  .A2({ S5491 }),
  .ZN({ S5920 })
);
NAND3_X1 #() 
NAND3_X1_6340_ (
  .A1({ S5857 }),
  .A2({ S5570 }),
  .A3({ S5920 }),
  .ZN({ S5921 })
);
NAND2_X1 #() 
NAND2_X1_5864_ (
  .A1({ S5921 }),
  .A2({ S25957[644] }),
  .ZN({ S5922 })
);
NAND3_X1 #() 
NAND3_X1_6341_ (
  .A1({ S5501 }),
  .A2({ S25957[643] }),
  .A3({ S8 }),
  .ZN({ S5923 })
);
AOI21_X1 #() 
AOI21_X1_3362_ (
  .A({ S25957[644] }),
  .B1({ S5766 }),
  .B2({ S5535 }),
  .ZN({ S5924 })
);
AOI21_X1 #() 
AOI21_X1_3363_ (
  .A({ S25957[645] }),
  .B1({ S5924 }),
  .B2({ S5923 }),
  .ZN({ S5925 })
);
AOI22_X1 #() 
AOI22_X1_661_ (
  .A1({ S5925 }),
  .A2({ S5922 }),
  .B1({ S5919 }),
  .B2({ S5916 }),
  .ZN({ S5926 })
);
OAI211_X1 #() 
OAI211_X1_2070_ (
  .A({ S5913 }),
  .B({ S5530 }),
  .C1({ S5926 }),
  .C2({ S25957[646] }),
  .ZN({ S5927 })
);
NAND3_X1 #() 
NAND3_X1_6342_ (
  .A1({ S25957[643] }),
  .A2({ S25957[642] }),
  .A3({ S5497 }),
  .ZN({ S5928 })
);
AOI21_X1 #() 
AOI21_X1_3364_ (
  .A({ S5495 }),
  .B1({ S5800 }),
  .B2({ S5928 }),
  .ZN({ S5930 })
);
NAND3_X1 #() 
NAND3_X1_6343_ (
  .A1({ S5554 }),
  .A2({ S0 }),
  .A3({ S5497 }),
  .ZN({ S5931 })
);
AND3_X1 #() 
AND3_X1_258_ (
  .A1({ S5931 }),
  .A2({ S5509 }),
  .A3({ S5495 }),
  .ZN({ S5932 })
);
OAI21_X1 #() 
OAI21_X1_3045_ (
  .A({ S25957[645] }),
  .B1({ S5932 }),
  .B2({ S5930 }),
  .ZN({ S5933 })
);
AOI21_X1 #() 
AOI21_X1_3365_ (
  .A({ S25957[643] }),
  .B1({ S5487 }),
  .B2({ S5604 }),
  .ZN({ S5934 })
);
NAND3_X1 #() 
NAND3_X1_6344_ (
  .A1({ S5542 }),
  .A2({ S5503 }),
  .A3({ S5473 }),
  .ZN({ S5935 })
);
NAND2_X1 #() 
NAND2_X1_5865_ (
  .A1({ S5935 }),
  .A2({ S5476 }),
  .ZN({ S5936 })
);
NAND2_X1 #() 
NAND2_X1_5866_ (
  .A1({ S5853 }),
  .A2({ S25957[644] }),
  .ZN({ S5937 })
);
OAI211_X1 #() 
OAI211_X1_2071_ (
  .A({ S5936 }),
  .B({ S5494 }),
  .C1({ S5934 }),
  .C2({ S5937 }),
  .ZN({ S5938 })
);
NAND3_X1 #() 
NAND3_X1_6345_ (
  .A1({ S5933 }),
  .A2({ S25957[646] }),
  .A3({ S5938 }),
  .ZN({ S5939 })
);
INV_X1 #() 
INV_X1_1889_ (
  .A({ S5862 }),
  .ZN({ S5941 })
);
NOR2_X1 #() 
NOR2_X1_1461_ (
  .A1({ S5479 }),
  .A2({ S5508 }),
  .ZN({ S5942 })
);
OAI21_X1 #() 
OAI21_X1_3046_ (
  .A({ S0 }),
  .B1({ S5942 }),
  .B2({ S5572 }),
  .ZN({ S5943 })
);
NAND3_X1 #() 
NAND3_X1_6346_ (
  .A1({ S5943 }),
  .A2({ S5941 }),
  .A3({ S25957[644] }),
  .ZN({ S5944 })
);
AOI22_X1 #() 
AOI22_X1_662_ (
  .A1({ S0 }),
  .A2({ S5500 }),
  .B1({ S3849 }),
  .B2({ S3846 }),
  .ZN({ S5945 })
);
AOI21_X1 #() 
AOI21_X1_3366_ (
  .A({ S5494 }),
  .B1({ S5751 }),
  .B2({ S5945 }),
  .ZN({ S5946 })
);
NAND2_X1 #() 
NAND2_X1_5867_ (
  .A1({ S5944 }),
  .A2({ S5946 }),
  .ZN({ S5947 })
);
NAND4_X1 #() 
NAND4_X1_704_ (
  .A1({ S5565 }),
  .A2({ S0 }),
  .A3({ S5475 }),
  .A4({ S8 }),
  .ZN({ S5948 })
);
AOI21_X1 #() 
AOI21_X1_3367_ (
  .A({ S25957[644] }),
  .B1({ S5948 }),
  .B2({ S5877 }),
  .ZN({ S5949 })
);
AND3_X1 #() 
AND3_X1_259_ (
  .A1({ S5687 }),
  .A2({ S8 }),
  .A3({ S5488 }),
  .ZN({ S5950 })
);
NAND2_X1 #() 
NAND2_X1_5868_ (
  .A1({ S25957[644] }),
  .A2({ S5607 }),
  .ZN({ S5952 })
);
NOR2_X1 #() 
NOR2_X1_1462_ (
  .A1({ S5950 }),
  .A2({ S5952 }),
  .ZN({ S5953 })
);
OAI21_X1 #() 
OAI21_X1_3047_ (
  .A({ S5494 }),
  .B1({ S5953 }),
  .B2({ S5949 }),
  .ZN({ S5954 })
);
NAND3_X1 #() 
NAND3_X1_6347_ (
  .A1({ S5954 }),
  .A2({ S5947 }),
  .A3({ S5465 }),
  .ZN({ S5955 })
);
NAND3_X1 #() 
NAND3_X1_6348_ (
  .A1({ S5939 }),
  .A2({ S5955 }),
  .A3({ S25957[647] }),
  .ZN({ S5956 })
);
NAND3_X1 #() 
NAND3_X1_6349_ (
  .A1({ S5927 }),
  .A2({ S5956 }),
  .A3({ S5905 }),
  .ZN({ S5957 })
);
NAND2_X1 #() 
NAND2_X1_5869_ (
  .A1({ S5906 }),
  .A2({ S5908 }),
  .ZN({ S5958 })
);
NAND2_X1 #() 
NAND2_X1_5870_ (
  .A1({ S5642 }),
  .A2({ S5476 }),
  .ZN({ S5959 })
);
NAND3_X1 #() 
NAND3_X1_6350_ (
  .A1({ S5958 }),
  .A2({ S5959 }),
  .A3({ S25957[645] }),
  .ZN({ S5960 })
);
NAND3_X1 #() 
NAND3_X1_6351_ (
  .A1({ S5480 }),
  .A2({ S5537 }),
  .A3({ S5660 }),
  .ZN({ S5961 })
);
NAND2_X1 #() 
NAND2_X1_5871_ (
  .A1({ S5961 }),
  .A2({ S25957[644] }),
  .ZN({ S5963 })
);
OAI21_X1 #() 
OAI21_X1_3048_ (
  .A({ S5495 }),
  .B1({ S5673 }),
  .B2({ S5910 }),
  .ZN({ S5964 })
);
NAND3_X1 #() 
NAND3_X1_6352_ (
  .A1({ S5964 }),
  .A2({ S5494 }),
  .A3({ S5963 }),
  .ZN({ S5965 })
);
NAND3_X1 #() 
NAND3_X1_6353_ (
  .A1({ S5960 }),
  .A2({ S5965 }),
  .A3({ S25957[646] }),
  .ZN({ S5966 })
);
NAND2_X1 #() 
NAND2_X1_5872_ (
  .A1({ S5919 }),
  .A2({ S5916 }),
  .ZN({ S5967 })
);
NOR2_X1 #() 
NOR2_X1_1463_ (
  .A1({ S25957[644] }),
  .A2({ S5535 }),
  .ZN({ S5968 })
);
OAI21_X1 #() 
OAI21_X1_3049_ (
  .A({ S5923 }),
  .B1({ S5968 }),
  .B2({ S5945 }),
  .ZN({ S5969 })
);
NAND3_X1 #() 
NAND3_X1_6354_ (
  .A1({ S5922 }),
  .A2({ S5969 }),
  .A3({ S5494 }),
  .ZN({ S5970 })
);
NAND3_X1 #() 
NAND3_X1_6355_ (
  .A1({ S5970 }),
  .A2({ S5465 }),
  .A3({ S5967 }),
  .ZN({ S5971 })
);
NAND3_X1 #() 
NAND3_X1_6356_ (
  .A1({ S5971 }),
  .A2({ S5530 }),
  .A3({ S5966 }),
  .ZN({ S5972 })
);
NAND2_X1 #() 
NAND2_X1_5873_ (
  .A1({ S5488 }),
  .A2({ S8 }),
  .ZN({ S5974 })
);
INV_X1 #() 
INV_X1_1890_ (
  .A({ S5783 }),
  .ZN({ S5975 })
);
NAND4_X1 #() 
NAND4_X1_705_ (
  .A1({ S5503 }),
  .A2({ S5484 }),
  .A3({ S5485 }),
  .A4({ S5508 }),
  .ZN({ S5976 })
);
AOI22_X1 #() 
AOI22_X1_663_ (
  .A1({ S5976 }),
  .A2({ S0 }),
  .B1({ S5975 }),
  .B2({ S5974 }),
  .ZN({ S5977 })
);
NOR2_X1 #() 
NOR2_X1_1464_ (
  .A1({ S5608 }),
  .A2({ S25957[643] }),
  .ZN({ S5978 })
);
OAI21_X1 #() 
OAI21_X1_3050_ (
  .A({ S5495 }),
  .B1({ S5673 }),
  .B2({ S5978 }),
  .ZN({ S5979 })
);
OAI211_X1 #() 
OAI211_X1_2072_ (
  .A({ S5979 }),
  .B({ S5494 }),
  .C1({ S5977 }),
  .C2({ S5495 }),
  .ZN({ S5980 })
);
AOI21_X1 #() 
AOI21_X1_3368_ (
  .A({ S25957[643] }),
  .B1({ S5514 }),
  .B2({ S5714 }),
  .ZN({ S5981 })
);
NOR2_X1 #() 
NOR2_X1_1465_ (
  .A1({ S5521 }),
  .A2({ S5783 }),
  .ZN({ S5982 })
);
OAI21_X1 #() 
OAI21_X1_3051_ (
  .A({ S25957[644] }),
  .B1({ S5981 }),
  .B2({ S5982 }),
  .ZN({ S5983 })
);
NAND3_X1 #() 
NAND3_X1_6357_ (
  .A1({ S5931 }),
  .A2({ S5495 }),
  .A3({ S5509 }),
  .ZN({ S5985 })
);
NAND3_X1 #() 
NAND3_X1_6358_ (
  .A1({ S5983 }),
  .A2({ S25957[645] }),
  .A3({ S5985 }),
  .ZN({ S5986 })
);
NAND3_X1 #() 
NAND3_X1_6359_ (
  .A1({ S5980 }),
  .A2({ S25957[646] }),
  .A3({ S5986 }),
  .ZN({ S5987 })
);
NAND3_X1 #() 
NAND3_X1_6360_ (
  .A1({ S0 }),
  .A2({ S5479 }),
  .A3({ S5485 }),
  .ZN({ S5988 })
);
OAI211_X1 #() 
OAI211_X1_2073_ (
  .A({ S25957[644] }),
  .B({ S5988 }),
  .C1({ S5862 }),
  .C2({ S5873 }),
  .ZN({ S5989 })
);
AND3_X1 #() 
AND3_X1_260_ (
  .A1({ S5545 }),
  .A2({ S5537 }),
  .A3({ S25957[643] }),
  .ZN({ S5990 })
);
OAI21_X1 #() 
OAI21_X1_3052_ (
  .A({ S5495 }),
  .B1({ S5990 }),
  .B2({ S5766 }),
  .ZN({ S5991 })
);
NAND3_X1 #() 
NAND3_X1_6361_ (
  .A1({ S5991 }),
  .A2({ S5989 }),
  .A3({ S25957[645] }),
  .ZN({ S5992 })
);
NAND2_X1 #() 
NAND2_X1_5874_ (
  .A1({ S5948 }),
  .A2({ S5877 }),
  .ZN({ S5993 })
);
NAND2_X1 #() 
NAND2_X1_5875_ (
  .A1({ S5993 }),
  .A2({ S5495 }),
  .ZN({ S5994 })
);
NAND2_X1 #() 
NAND2_X1_5876_ (
  .A1({ S5602 }),
  .A2({ S5687 }),
  .ZN({ S5996 })
);
AOI21_X1 #() 
AOI21_X1_3369_ (
  .A({ S5495 }),
  .B1({ S25957[643] }),
  .B2({ S5496 }),
  .ZN({ S5997 })
);
AOI21_X1 #() 
AOI21_X1_3370_ (
  .A({ S25957[645] }),
  .B1({ S5997 }),
  .B2({ S5996 }),
  .ZN({ S5998 })
);
NAND2_X1 #() 
NAND2_X1_5877_ (
  .A1({ S5998 }),
  .A2({ S5994 }),
  .ZN({ S5999 })
);
NAND3_X1 #() 
NAND3_X1_6362_ (
  .A1({ S5999 }),
  .A2({ S5992 }),
  .A3({ S5465 }),
  .ZN({ S6000 })
);
NAND3_X1 #() 
NAND3_X1_6363_ (
  .A1({ S5987 }),
  .A2({ S6000 }),
  .A3({ S25957[647] }),
  .ZN({ S6001 })
);
NAND3_X1 #() 
NAND3_X1_6364_ (
  .A1({ S5972 }),
  .A2({ S6001 }),
  .A3({ S25957[744] }),
  .ZN({ S6002 })
);
NAND3_X1 #() 
NAND3_X1_6365_ (
  .A1({ S5957 }),
  .A2({ S6002 }),
  .A3({ S25957[808] }),
  .ZN({ S6003 })
);
INV_X1 #() 
INV_X1_1891_ (
  .A({ S25957[808] }),
  .ZN({ S6004 })
);
NAND3_X1 #() 
NAND3_X1_6366_ (
  .A1({ S5927 }),
  .A2({ S5956 }),
  .A3({ S25957[744] }),
  .ZN({ S6005 })
);
NAND3_X1 #() 
NAND3_X1_6367_ (
  .A1({ S5972 }),
  .A2({ S6001 }),
  .A3({ S5905 }),
  .ZN({ S6007 })
);
NAND3_X1 #() 
NAND3_X1_6368_ (
  .A1({ S6005 }),
  .A2({ S6007 }),
  .A3({ S6004 }),
  .ZN({ S6008 })
);
NAND3_X1 #() 
NAND3_X1_6369_ (
  .A1({ S6003 }),
  .A2({ S6008 }),
  .A3({ S25957[648] }),
  .ZN({ S6009 })
);
AOI21_X1 #() 
AOI21_X1_3371_ (
  .A({ S6004 }),
  .B1({ S6005 }),
  .B2({ S6007 }),
  .ZN({ S6010 })
);
AOI21_X1 #() 
AOI21_X1_3372_ (
  .A({ S25957[808] }),
  .B1({ S5957 }),
  .B2({ S6002 }),
  .ZN({ S6011 })
);
OAI21_X1 #() 
OAI21_X1_3053_ (
  .A({ S4794 }),
  .B1({ S6010 }),
  .B2({ S6011 }),
  .ZN({ S6012 })
);
NAND2_X1 #() 
NAND2_X1_5878_ (
  .A1({ S6012 }),
  .A2({ S6009 }),
  .ZN({ S25957[520] })
);
NAND2_X1 #() 
NAND2_X1_5879_ (
  .A1({ S3398 }),
  .A2({ S3396 }),
  .ZN({ S25957[745] })
);
INV_X1 #() 
INV_X1_1892_ (
  .A({ S25957[745] }),
  .ZN({ S6013 })
);
OAI21_X1 #() 
OAI21_X1_3054_ (
  .A({ S5532 }),
  .B1({ S5502 }),
  .B2({ S5689 }),
  .ZN({ S6014 })
);
NAND3_X1 #() 
NAND3_X1_6370_ (
  .A1({ S0 }),
  .A2({ S5484 }),
  .A3({ S5537 }),
  .ZN({ S6016 })
);
NAND3_X1 #() 
NAND3_X1_6371_ (
  .A1({ S5699 }),
  .A2({ S6016 }),
  .A3({ S25957[644] }),
  .ZN({ S6017 })
);
OAI211_X1 #() 
OAI211_X1_2074_ (
  .A({ S6017 }),
  .B({ S25957[645] }),
  .C1({ S6014 }),
  .C2({ S25957[644] }),
  .ZN({ S6018 })
);
NAND2_X1 #() 
NAND2_X1_5880_ (
  .A1({ S5661 }),
  .A2({ S5988 }),
  .ZN({ S6019 })
);
NAND3_X1 #() 
NAND3_X1_6372_ (
  .A1({ S5488 }),
  .A2({ S25957[643] }),
  .A3({ S5484 }),
  .ZN({ S6020 })
);
NAND4_X1 #() 
NAND4_X1_706_ (
  .A1({ S5565 }),
  .A2({ S5714 }),
  .A3({ S5488 }),
  .A4({ S0 }),
  .ZN({ S6021 })
);
NAND3_X1 #() 
NAND3_X1_6373_ (
  .A1({ S6021 }),
  .A2({ S6020 }),
  .A3({ S5495 }),
  .ZN({ S6022 })
);
OAI211_X1 #() 
OAI211_X1_2075_ (
  .A({ S6022 }),
  .B({ S5494 }),
  .C1({ S6019 }),
  .C2({ S5495 }),
  .ZN({ S6023 })
);
NAND3_X1 #() 
NAND3_X1_6374_ (
  .A1({ S6023 }),
  .A2({ S6018 }),
  .A3({ S25957[646] }),
  .ZN({ S6024 })
);
AOI21_X1 #() 
AOI21_X1_3373_ (
  .A({ S0 }),
  .B1({ S5548 }),
  .B2({ S5475 }),
  .ZN({ S6025 })
);
NAND3_X1 #() 
NAND3_X1_6375_ (
  .A1({ S5879 }),
  .A2({ S5703 }),
  .A3({ S5495 }),
  .ZN({ S6027 })
);
OAI211_X1 #() 
OAI211_X1_2076_ (
  .A({ S6027 }),
  .B({ S25957[645] }),
  .C1({ S6025 }),
  .C2({ S5533 }),
  .ZN({ S6028 })
);
NAND2_X1 #() 
NAND2_X1_5881_ (
  .A1({ S25957[643] }),
  .A2({ S5551 }),
  .ZN({ S6029 })
);
NAND2_X1 #() 
NAND2_X1_5882_ (
  .A1({ S5660 }),
  .A2({ S5537 }),
  .ZN({ S6030 })
);
OAI211_X1 #() 
OAI211_X1_2077_ (
  .A({ S25957[644] }),
  .B({ S6029 }),
  .C1({ S6030 }),
  .C2({ S25957[643] }),
  .ZN({ S6031 })
);
NAND2_X1 #() 
NAND2_X1_5883_ (
  .A1({ S5758 }),
  .A2({ S5495 }),
  .ZN({ S6032 })
);
OAI211_X1 #() 
OAI211_X1_2078_ (
  .A({ S5494 }),
  .B({ S6031 }),
  .C1({ S6032 }),
  .C2({ S5547 }),
  .ZN({ S6033 })
);
NAND3_X1 #() 
NAND3_X1_6376_ (
  .A1({ S6033 }),
  .A2({ S5465 }),
  .A3({ S6028 }),
  .ZN({ S6034 })
);
NAND3_X1 #() 
NAND3_X1_6377_ (
  .A1({ S6034 }),
  .A2({ S25957[647] }),
  .A3({ S6024 }),
  .ZN({ S6035 })
);
NAND2_X1 #() 
NAND2_X1_5884_ (
  .A1({ S5865 }),
  .A2({ S5768 }),
  .ZN({ S6036 })
);
AOI21_X1 #() 
AOI21_X1_3374_ (
  .A({ S5555 }),
  .B1({ S6036 }),
  .B2({ S25957[644] }),
  .ZN({ S6038 })
);
NAND2_X1 #() 
NAND2_X1_5885_ (
  .A1({ S5858 }),
  .A2({ S5779 }),
  .ZN({ S6039 })
);
OAI211_X1 #() 
OAI211_X1_2079_ (
  .A({ S5492 }),
  .B({ S5495 }),
  .C1({ S5554 }),
  .C2({ S25957[643] }),
  .ZN({ S6040 })
);
NAND3_X1 #() 
NAND3_X1_6378_ (
  .A1({ S6039 }),
  .A2({ S5494 }),
  .A3({ S6040 }),
  .ZN({ S6041 })
);
OAI211_X1 #() 
OAI211_X1_2080_ (
  .A({ S5465 }),
  .B({ S6041 }),
  .C1({ S6038 }),
  .C2({ S5494 }),
  .ZN({ S6042 })
);
NAND3_X1 #() 
NAND3_X1_6379_ (
  .A1({ S5501 }),
  .A2({ S5714 }),
  .A3({ S0 }),
  .ZN({ S6043 })
);
OAI211_X1 #() 
OAI211_X1_2081_ (
  .A({ S6043 }),
  .B({ S25957[644] }),
  .C1({ S5502 }),
  .C2({ S5689 }),
  .ZN({ S6044 })
);
NAND3_X1 #() 
NAND3_X1_6380_ (
  .A1({ S5619 }),
  .A2({ S5853 }),
  .A3({ S5495 }),
  .ZN({ S6045 })
);
NAND3_X1 #() 
NAND3_X1_6381_ (
  .A1({ S6044 }),
  .A2({ S6045 }),
  .A3({ S5494 }),
  .ZN({ S6046 })
);
NAND3_X1 #() 
NAND3_X1_6382_ (
  .A1({ S5503 }),
  .A2({ S0 }),
  .A3({ S5500 }),
  .ZN({ S6047 })
);
NAND3_X1 #() 
NAND3_X1_6383_ (
  .A1({ S5886 }),
  .A2({ S25957[644] }),
  .A3({ S6047 }),
  .ZN({ S6049 })
);
NAND3_X1 #() 
NAND3_X1_6384_ (
  .A1({ S5724 }),
  .A2({ S5565 }),
  .A3({ S5714 }),
  .ZN({ S6050 })
);
NAND3_X1 #() 
NAND3_X1_6385_ (
  .A1({ S6049 }),
  .A2({ S6050 }),
  .A3({ S25957[645] }),
  .ZN({ S6051 })
);
NAND3_X1 #() 
NAND3_X1_6386_ (
  .A1({ S6046 }),
  .A2({ S6051 }),
  .A3({ S25957[646] }),
  .ZN({ S6052 })
);
NAND3_X1 #() 
NAND3_X1_6387_ (
  .A1({ S6042 }),
  .A2({ S5530 }),
  .A3({ S6052 }),
  .ZN({ S6053 })
);
NAND3_X1 #() 
NAND3_X1_6388_ (
  .A1({ S6035 }),
  .A2({ S6053 }),
  .A3({ S6013 }),
  .ZN({ S6054 })
);
NAND2_X1 #() 
NAND2_X1_5886_ (
  .A1({ S6046 }),
  .A2({ S6051 }),
  .ZN({ S6055 })
);
NAND2_X1 #() 
NAND2_X1_5887_ (
  .A1({ S6055 }),
  .A2({ S25957[646] }),
  .ZN({ S6056 })
);
NAND2_X1 #() 
NAND2_X1_5888_ (
  .A1({ S6036 }),
  .A2({ S25957[644] }),
  .ZN({ S6057 })
);
NAND2_X1 #() 
NAND2_X1_5889_ (
  .A1({ S5554 }),
  .A2({ S0 }),
  .ZN({ S6058 })
);
AOI21_X1 #() 
AOI21_X1_3375_ (
  .A({ S5494 }),
  .B1({ S6058 }),
  .B2({ S5495 }),
  .ZN({ S6060 })
);
NAND2_X1 #() 
NAND2_X1_5890_ (
  .A1({ S6057 }),
  .A2({ S6060 }),
  .ZN({ S6061 })
);
NAND2_X1 #() 
NAND2_X1_5891_ (
  .A1({ S5484 }),
  .A2({ S5508 }),
  .ZN({ S6062 })
);
NOR2_X1 #() 
NOR2_X1_1466_ (
  .A1({ S6062 }),
  .A2({ S25957[643] }),
  .ZN({ S6063 })
);
OAI21_X1 #() 
OAI21_X1_3055_ (
  .A({ S25957[644] }),
  .B1({ S5468 }),
  .B2({ S6063 }),
  .ZN({ S6064 })
);
INV_X1 #() 
INV_X1_1893_ (
  .A({ S5492 }),
  .ZN({ S6065 })
);
OAI21_X1 #() 
OAI21_X1_3056_ (
  .A({ S5495 }),
  .B1({ S5871 }),
  .B2({ S6065 }),
  .ZN({ S6066 })
);
NAND3_X1 #() 
NAND3_X1_6389_ (
  .A1({ S6064 }),
  .A2({ S6066 }),
  .A3({ S5494 }),
  .ZN({ S6067 })
);
NAND3_X1 #() 
NAND3_X1_6390_ (
  .A1({ S6067 }),
  .A2({ S6061 }),
  .A3({ S5465 }),
  .ZN({ S6068 })
);
NAND3_X1 #() 
NAND3_X1_6391_ (
  .A1({ S6056 }),
  .A2({ S5530 }),
  .A3({ S6068 }),
  .ZN({ S6069 })
);
NAND2_X1 #() 
NAND2_X1_5892_ (
  .A1({ S6021 }),
  .A2({ S6020 }),
  .ZN({ S6071 })
);
NAND2_X1 #() 
NAND2_X1_5893_ (
  .A1({ S6071 }),
  .A2({ S5494 }),
  .ZN({ S6072 })
);
NAND2_X1 #() 
NAND2_X1_5894_ (
  .A1({ S6014 }),
  .A2({ S25957[645] }),
  .ZN({ S6073 })
);
NAND3_X1 #() 
NAND3_X1_6392_ (
  .A1({ S6073 }),
  .A2({ S6072 }),
  .A3({ S5495 }),
  .ZN({ S6074 })
);
NAND2_X1 #() 
NAND2_X1_5895_ (
  .A1({ S6019 }),
  .A2({ S5494 }),
  .ZN({ S6075 })
);
NAND2_X1 #() 
NAND2_X1_5896_ (
  .A1({ S5699 }),
  .A2({ S6016 }),
  .ZN({ S6076 })
);
BUF_X1 #() 
BUF_X1_1_ (
  .A({ key[0] }),
  .Z({ S25956[0] })
);
BUF_X1 #() 
BUF_X1_2_ (
  .A({ key[1] }),
  .Z({ S25956[1] })
);
BUF_X1 #() 
BUF_X1_3_ (
  .A({ key[10] }),
  .Z({ S25956[10] })
);
BUF_X1 #() 
BUF_X1_4_ (
  .A({ key[100] }),
  .Z({ S25956[100] })
);
BUF_X1 #() 
BUF_X1_5_ (
  .A({ key[101] }),
  .Z({ S25956[101] })
);
BUF_X1 #() 
BUF_X1_6_ (
  .A({ key[102] }),
  .Z({ S25956[102] })
);
BUF_X1 #() 
BUF_X1_7_ (
  .A({ key[103] }),
  .Z({ S25956[103] })
);
BUF_X1 #() 
BUF_X1_8_ (
  .A({ key[104] }),
  .Z({ S25956[104] })
);
BUF_X1 #() 
BUF_X1_9_ (
  .A({ key[105] }),
  .Z({ S25956[105] })
);
BUF_X1 #() 
BUF_X1_10_ (
  .A({ key[106] }),
  .Z({ S25956[106] })
);
BUF_X1 #() 
BUF_X1_11_ (
  .A({ key[107] }),
  .Z({ S25956[107] })
);
BUF_X1 #() 
BUF_X1_12_ (
  .A({ key[108] }),
  .Z({ S25956[108] })
);
BUF_X1 #() 
BUF_X1_13_ (
  .A({ key[109] }),
  .Z({ S25956[109] })
);
BUF_X1 #() 
BUF_X1_14_ (
  .A({ key[11] }),
  .Z({ S25956[11] })
);
BUF_X1 #() 
BUF_X1_15_ (
  .A({ key[110] }),
  .Z({ S25956[110] })
);
BUF_X1 #() 
BUF_X1_16_ (
  .A({ key[111] }),
  .Z({ S25956[111] })
);
BUF_X1 #() 
BUF_X1_17_ (
  .A({ key[112] }),
  .Z({ S25956[112] })
);
BUF_X1 #() 
BUF_X1_18_ (
  .A({ key[113] }),
  .Z({ S25956[113] })
);
BUF_X1 #() 
BUF_X1_19_ (
  .A({ key[114] }),
  .Z({ S25956[114] })
);
BUF_X1 #() 
BUF_X1_20_ (
  .A({ key[115] }),
  .Z({ S25956[115] })
);
BUF_X1 #() 
BUF_X1_21_ (
  .A({ key[116] }),
  .Z({ S25956[116] })
);
BUF_X1 #() 
BUF_X1_22_ (
  .A({ key[117] }),
  .Z({ S25956[117] })
);
BUF_X1 #() 
BUF_X1_23_ (
  .A({ key[118] }),
  .Z({ S25956[118] })
);
BUF_X1 #() 
BUF_X1_24_ (
  .A({ key[119] }),
  .Z({ S25956[119] })
);
BUF_X1 #() 
BUF_X1_25_ (
  .A({ key[12] }),
  .Z({ S25956[12] })
);
BUF_X1 #() 
BUF_X1_26_ (
  .A({ key[120] }),
  .Z({ S25956[120] })
);
BUF_X1 #() 
BUF_X1_27_ (
  .A({ key[121] }),
  .Z({ S25956[121] })
);
BUF_X1 #() 
BUF_X1_28_ (
  .A({ key[122] }),
  .Z({ S25956[122] })
);
BUF_X1 #() 
BUF_X1_29_ (
  .A({ key[123] }),
  .Z({ S25956[123] })
);
BUF_X1 #() 
BUF_X1_30_ (
  .A({ key[124] }),
  .Z({ S25956[124] })
);
BUF_X1 #() 
BUF_X1_31_ (
  .A({ key[125] }),
  .Z({ S25956[125] })
);
BUF_X1 #() 
BUF_X1_32_ (
  .A({ key[126] }),
  .Z({ S25956[126] })
);
BUF_X1 #() 
BUF_X1_33_ (
  .A({ key[127] }),
  .Z({ S25956[127] })
);
BUF_X1 #() 
BUF_X1_34_ (
  .A({ key[13] }),
  .Z({ S25956[13] })
);
BUF_X1 #() 
BUF_X1_35_ (
  .A({ key[14] }),
  .Z({ S25956[14] })
);
BUF_X1 #() 
BUF_X1_36_ (
  .A({ key[15] }),
  .Z({ S25956[15] })
);
BUF_X1 #() 
BUF_X1_37_ (
  .A({ key[16] }),
  .Z({ S25956[16] })
);
BUF_X1 #() 
BUF_X1_38_ (
  .A({ key[17] }),
  .Z({ S25956[17] })
);
BUF_X1 #() 
BUF_X1_39_ (
  .A({ key[18] }),
  .Z({ S25956[18] })
);
BUF_X1 #() 
BUF_X1_40_ (
  .A({ key[19] }),
  .Z({ S25956[19] })
);
BUF_X1 #() 
BUF_X1_41_ (
  .A({ key[2] }),
  .Z({ S25956[2] })
);
BUF_X1 #() 
BUF_X1_42_ (
  .A({ key[20] }),
  .Z({ S25956[20] })
);
BUF_X1 #() 
BUF_X1_43_ (
  .A({ key[21] }),
  .Z({ S25956[21] })
);
BUF_X1 #() 
BUF_X1_44_ (
  .A({ key[22] }),
  .Z({ S25956[22] })
);
BUF_X1 #() 
BUF_X1_45_ (
  .A({ key[23] }),
  .Z({ S25956[23] })
);
BUF_X1 #() 
BUF_X1_46_ (
  .A({ key[24] }),
  .Z({ S25956[24] })
);
BUF_X1 #() 
BUF_X1_47_ (
  .A({ key[25] }),
  .Z({ S25956[25] })
);
BUF_X1 #() 
BUF_X1_48_ (
  .A({ key[26] }),
  .Z({ S25956[26] })
);
BUF_X1 #() 
BUF_X1_49_ (
  .A({ key[27] }),
  .Z({ S25956[27] })
);
BUF_X1 #() 
BUF_X1_50_ (
  .A({ key[28] }),
  .Z({ S25956[28] })
);
BUF_X1 #() 
BUF_X1_51_ (
  .A({ key[29] }),
  .Z({ S25956[29] })
);
BUF_X1 #() 
BUF_X1_52_ (
  .A({ key[3] }),
  .Z({ S25956[3] })
);
BUF_X1 #() 
BUF_X1_53_ (
  .A({ key[30] }),
  .Z({ S25956[30] })
);
BUF_X1 #() 
BUF_X1_54_ (
  .A({ key[31] }),
  .Z({ S25956[31] })
);
BUF_X1 #() 
BUF_X1_55_ (
  .A({ key[32] }),
  .Z({ S25956[32] })
);
BUF_X1 #() 
BUF_X1_56_ (
  .A({ key[33] }),
  .Z({ S25956[33] })
);
BUF_X1 #() 
BUF_X1_57_ (
  .A({ key[34] }),
  .Z({ S25956[34] })
);
BUF_X1 #() 
BUF_X1_58_ (
  .A({ key[35] }),
  .Z({ S25956[35] })
);
BUF_X1 #() 
BUF_X1_59_ (
  .A({ key[36] }),
  .Z({ S25956[36] })
);
BUF_X1 #() 
BUF_X1_60_ (
  .A({ key[37] }),
  .Z({ S25956[37] })
);
BUF_X1 #() 
BUF_X1_61_ (
  .A({ key[38] }),
  .Z({ S25956[38] })
);
BUF_X1 #() 
BUF_X1_62_ (
  .A({ key[39] }),
  .Z({ S25956[39] })
);
BUF_X1 #() 
BUF_X1_63_ (
  .A({ key[4] }),
  .Z({ S25956[4] })
);
BUF_X1 #() 
BUF_X1_64_ (
  .A({ key[40] }),
  .Z({ S25956[40] })
);
BUF_X1 #() 
BUF_X1_65_ (
  .A({ key[41] }),
  .Z({ S25956[41] })
);
BUF_X1 #() 
BUF_X1_66_ (
  .A({ key[42] }),
  .Z({ S25956[42] })
);
BUF_X1 #() 
BUF_X1_67_ (
  .A({ key[43] }),
  .Z({ S25956[43] })
);
BUF_X1 #() 
BUF_X1_68_ (
  .A({ key[44] }),
  .Z({ S25956[44] })
);
BUF_X1 #() 
BUF_X1_69_ (
  .A({ key[45] }),
  .Z({ S25956[45] })
);
BUF_X1 #() 
BUF_X1_70_ (
  .A({ key[46] }),
  .Z({ S25956[46] })
);
BUF_X1 #() 
BUF_X1_71_ (
  .A({ key[47] }),
  .Z({ S25956[47] })
);
BUF_X1 #() 
BUF_X1_72_ (
  .A({ key[48] }),
  .Z({ S25956[48] })
);
BUF_X1 #() 
BUF_X1_73_ (
  .A({ key[49] }),
  .Z({ S25956[49] })
);
BUF_X1 #() 
BUF_X1_74_ (
  .A({ key[5] }),
  .Z({ S25956[5] })
);
BUF_X1 #() 
BUF_X1_75_ (
  .A({ key[50] }),
  .Z({ S25956[50] })
);
BUF_X1 #() 
BUF_X1_76_ (
  .A({ key[51] }),
  .Z({ S25956[51] })
);
BUF_X1 #() 
BUF_X1_77_ (
  .A({ key[52] }),
  .Z({ S25956[52] })
);
BUF_X1 #() 
BUF_X1_78_ (
  .A({ key[53] }),
  .Z({ S25956[53] })
);
BUF_X1 #() 
BUF_X1_79_ (
  .A({ key[54] }),
  .Z({ S25956[54] })
);
BUF_X1 #() 
BUF_X1_80_ (
  .A({ key[55] }),
  .Z({ S25956[55] })
);
BUF_X1 #() 
BUF_X1_81_ (
  .A({ key[56] }),
  .Z({ S25956[56] })
);
BUF_X1 #() 
BUF_X1_82_ (
  .A({ key[57] }),
  .Z({ S25956[57] })
);
BUF_X1 #() 
BUF_X1_83_ (
  .A({ key[58] }),
  .Z({ S25956[58] })
);
BUF_X1 #() 
BUF_X1_84_ (
  .A({ key[59] }),
  .Z({ S25956[59] })
);
BUF_X1 #() 
BUF_X1_85_ (
  .A({ key[6] }),
  .Z({ S25956[6] })
);
BUF_X1 #() 
BUF_X1_86_ (
  .A({ key[60] }),
  .Z({ S25956[60] })
);
BUF_X1 #() 
BUF_X1_87_ (
  .A({ key[61] }),
  .Z({ S25956[61] })
);
BUF_X1 #() 
BUF_X1_88_ (
  .A({ key[62] }),
  .Z({ S25956[62] })
);
BUF_X1 #() 
BUF_X1_89_ (
  .A({ key[63] }),
  .Z({ S25956[63] })
);
BUF_X1 #() 
BUF_X1_90_ (
  .A({ key[64] }),
  .Z({ S25956[64] })
);
BUF_X1 #() 
BUF_X1_91_ (
  .A({ key[65] }),
  .Z({ S25956[65] })
);
BUF_X1 #() 
BUF_X1_92_ (
  .A({ key[66] }),
  .Z({ S25956[66] })
);
BUF_X1 #() 
BUF_X1_93_ (
  .A({ key[67] }),
  .Z({ S25956[67] })
);
BUF_X1 #() 
BUF_X1_94_ (
  .A({ key[68] }),
  .Z({ S25956[68] })
);
BUF_X1 #() 
BUF_X1_95_ (
  .A({ key[69] }),
  .Z({ S25956[69] })
);
BUF_X1 #() 
BUF_X1_96_ (
  .A({ key[7] }),
  .Z({ S25956[7] })
);
BUF_X1 #() 
BUF_X1_97_ (
  .A({ key[70] }),
  .Z({ S25956[70] })
);
BUF_X1 #() 
BUF_X1_98_ (
  .A({ key[71] }),
  .Z({ S25956[71] })
);
BUF_X1 #() 
BUF_X1_99_ (
  .A({ key[72] }),
  .Z({ S25956[72] })
);
BUF_X1 #() 
BUF_X1_100_ (
  .A({ key[73] }),
  .Z({ S25956[73] })
);
BUF_X1 #() 
BUF_X1_101_ (
  .A({ key[74] }),
  .Z({ S25956[74] })
);
BUF_X1 #() 
BUF_X1_102_ (
  .A({ key[75] }),
  .Z({ S25956[75] })
);
BUF_X1 #() 
BUF_X1_103_ (
  .A({ key[76] }),
  .Z({ S25956[76] })
);
BUF_X1 #() 
BUF_X1_104_ (
  .A({ key[77] }),
  .Z({ S25956[77] })
);
BUF_X1 #() 
BUF_X1_105_ (
  .A({ key[78] }),
  .Z({ S25956[78] })
);
BUF_X1 #() 
BUF_X1_106_ (
  .A({ key[79] }),
  .Z({ S25956[79] })
);
BUF_X1 #() 
BUF_X1_107_ (
  .A({ key[8] }),
  .Z({ S25956[8] })
);
BUF_X1 #() 
BUF_X1_108_ (
  .A({ key[80] }),
  .Z({ S25956[80] })
);
BUF_X1 #() 
BUF_X1_109_ (
  .A({ key[81] }),
  .Z({ S25956[81] })
);
BUF_X1 #() 
BUF_X1_110_ (
  .A({ key[82] }),
  .Z({ S25956[82] })
);
BUF_X1 #() 
BUF_X1_111_ (
  .A({ key[83] }),
  .Z({ S25956[83] })
);
BUF_X1 #() 
BUF_X1_112_ (
  .A({ key[84] }),
  .Z({ S25956[84] })
);
BUF_X1 #() 
BUF_X1_113_ (
  .A({ key[85] }),
  .Z({ S25956[85] })
);
BUF_X1 #() 
BUF_X1_114_ (
  .A({ key[86] }),
  .Z({ S25956[86] })
);
BUF_X1 #() 
BUF_X1_115_ (
  .A({ key[87] }),
  .Z({ S25956[87] })
);
BUF_X1 #() 
BUF_X1_116_ (
  .A({ key[88] }),
  .Z({ S25956[88] })
);
BUF_X1 #() 
BUF_X1_117_ (
  .A({ key[89] }),
  .Z({ S25956[89] })
);
BUF_X1 #() 
BUF_X1_118_ (
  .A({ key[9] }),
  .Z({ S25956[9] })
);
BUF_X1 #() 
BUF_X1_119_ (
  .A({ key[90] }),
  .Z({ S25956[90] })
);
BUF_X1 #() 
BUF_X1_120_ (
  .A({ key[91] }),
  .Z({ S25956[91] })
);
BUF_X1 #() 
BUF_X1_121_ (
  .A({ key[92] }),
  .Z({ S25956[92] })
);
BUF_X1 #() 
BUF_X1_122_ (
  .A({ key[93] }),
  .Z({ S25956[93] })
);
BUF_X1 #() 
BUF_X1_123_ (
  .A({ key[94] }),
  .Z({ S25956[94] })
);
BUF_X1 #() 
BUF_X1_124_ (
  .A({ key[95] }),
  .Z({ S25956[95] })
);
BUF_X1 #() 
BUF_X1_125_ (
  .A({ key[96] }),
  .Z({ S25956[96] })
);
BUF_X1 #() 
BUF_X1_126_ (
  .A({ key[97] }),
  .Z({ S25956[97] })
);
BUF_X1 #() 
BUF_X1_127_ (
  .A({ key[98] }),
  .Z({ S25956[98] })
);
BUF_X1 #() 
BUF_X1_128_ (
  .A({ key[99] }),
  .Z({ S25956[99] })
);
BUF_X1 #() 
BUF_X1_129_ (
  .A({ S25957[0] }),
  .Z({ w[0] })
);
BUF_X1 #() 
BUF_X1_130_ (
  .A({ S25957[1] }),
  .Z({ w[1] })
);
BUF_X1 #() 
BUF_X1_131_ (
  .A({ S25957[10] }),
  .Z({ w[10] })
);
BUF_X1 #() 
BUF_X1_132_ (
  .A({ S25957[100] }),
  .Z({ w[100] })
);
BUF_X1 #() 
BUF_X1_133_ (
  .A({ S25957[1000] }),
  .Z({ w[1000] })
);
BUF_X1 #() 
BUF_X1_134_ (
  .A({ S25957[1001] }),
  .Z({ w[1001] })
);
BUF_X1 #() 
BUF_X1_135_ (
  .A({ S25957[1002] }),
  .Z({ w[1002] })
);
BUF_X1 #() 
BUF_X1_136_ (
  .A({ S25957[1003] }),
  .Z({ w[1003] })
);
BUF_X1 #() 
BUF_X1_137_ (
  .A({ S25957[1004] }),
  .Z({ w[1004] })
);
BUF_X1 #() 
BUF_X1_138_ (
  .A({ S25957[1005] }),
  .Z({ w[1005] })
);
BUF_X1 #() 
BUF_X1_139_ (
  .A({ S25957[1006] }),
  .Z({ w[1006] })
);
BUF_X1 #() 
BUF_X1_140_ (
  .A({ S25957[1007] }),
  .Z({ w[1007] })
);
BUF_X1 #() 
BUF_X1_141_ (
  .A({ S25957[1008] }),
  .Z({ w[1008] })
);
BUF_X1 #() 
BUF_X1_142_ (
  .A({ S25957[1009] }),
  .Z({ w[1009] })
);
BUF_X1 #() 
BUF_X1_143_ (
  .A({ S25957[101] }),
  .Z({ w[101] })
);
BUF_X1 #() 
BUF_X1_144_ (
  .A({ S25957[1010] }),
  .Z({ w[1010] })
);
BUF_X1 #() 
BUF_X1_145_ (
  .A({ S25957[1011] }),
  .Z({ w[1011] })
);
BUF_X1 #() 
BUF_X1_146_ (
  .A({ S25957[1012] }),
  .Z({ w[1012] })
);
BUF_X1 #() 
BUF_X1_147_ (
  .A({ S25957[1013] }),
  .Z({ w[1013] })
);
BUF_X1 #() 
BUF_X1_148_ (
  .A({ S25957[1014] }),
  .Z({ w[1014] })
);
BUF_X1 #() 
BUF_X1_149_ (
  .A({ S25957[1015] }),
  .Z({ w[1015] })
);
BUF_X1 #() 
BUF_X1_150_ (
  .A({ S25957[1016] }),
  .Z({ w[1016] })
);
BUF_X1 #() 
BUF_X1_151_ (
  .A({ S25957[1017] }),
  .Z({ w[1017] })
);
BUF_X1 #() 
BUF_X1_152_ (
  .A({ S25957[1018] }),
  .Z({ w[1018] })
);
BUF_X1 #() 
BUF_X1_153_ (
  .A({ S25957[1019] }),
  .Z({ w[1019] })
);
BUF_X1 #() 
BUF_X1_154_ (
  .A({ S25957[102] }),
  .Z({ w[102] })
);
BUF_X1 #() 
BUF_X1_155_ (
  .A({ S25957[1020] }),
  .Z({ w[1020] })
);
BUF_X1 #() 
BUF_X1_156_ (
  .A({ S25957[1021] }),
  .Z({ w[1021] })
);
BUF_X1 #() 
BUF_X1_157_ (
  .A({ S25957[1022] }),
  .Z({ w[1022] })
);
BUF_X1 #() 
BUF_X1_158_ (
  .A({ S25957[1023] }),
  .Z({ w[1023] })
);
BUF_X1 #() 
BUF_X1_159_ (
  .A({ S25957[1024] }),
  .Z({ w[1024] })
);
BUF_X1 #() 
BUF_X1_160_ (
  .A({ S25957[1025] }),
  .Z({ w[1025] })
);
BUF_X1 #() 
BUF_X1_161_ (
  .A({ S25957[1026] }),
  .Z({ w[1026] })
);
BUF_X1 #() 
BUF_X1_162_ (
  .A({ S25957[1027] }),
  .Z({ w[1027] })
);
BUF_X1 #() 
BUF_X1_163_ (
  .A({ S25957[1028] }),
  .Z({ w[1028] })
);
BUF_X1 #() 
BUF_X1_164_ (
  .A({ S25957[1029] }),
  .Z({ w[1029] })
);
BUF_X1 #() 
BUF_X1_165_ (
  .A({ S25957[103] }),
  .Z({ w[103] })
);
BUF_X1 #() 
BUF_X1_166_ (
  .A({ S25957[1030] }),
  .Z({ w[1030] })
);
BUF_X1 #() 
BUF_X1_167_ (
  .A({ S25957[1031] }),
  .Z({ w[1031] })
);
BUF_X1 #() 
BUF_X1_168_ (
  .A({ S25957[1032] }),
  .Z({ w[1032] })
);
BUF_X1 #() 
BUF_X1_169_ (
  .A({ S25957[1033] }),
  .Z({ w[1033] })
);
BUF_X1 #() 
BUF_X1_170_ (
  .A({ S25957[1034] }),
  .Z({ w[1034] })
);
BUF_X1 #() 
BUF_X1_171_ (
  .A({ S25957[1035] }),
  .Z({ w[1035] })
);
BUF_X1 #() 
BUF_X1_172_ (
  .A({ S25957[1036] }),
  .Z({ w[1036] })
);
BUF_X1 #() 
BUF_X1_173_ (
  .A({ S25957[1037] }),
  .Z({ w[1037] })
);
BUF_X1 #() 
BUF_X1_174_ (
  .A({ S25957[1038] }),
  .Z({ w[1038] })
);
BUF_X1 #() 
BUF_X1_175_ (
  .A({ S25957[1039] }),
  .Z({ w[1039] })
);
BUF_X1 #() 
BUF_X1_176_ (
  .A({ S25957[104] }),
  .Z({ w[104] })
);
BUF_X1 #() 
BUF_X1_177_ (
  .A({ S25957[1040] }),
  .Z({ w[1040] })
);
BUF_X1 #() 
BUF_X1_178_ (
  .A({ S25957[1041] }),
  .Z({ w[1041] })
);
BUF_X1 #() 
BUF_X1_179_ (
  .A({ S25957[1042] }),
  .Z({ w[1042] })
);
BUF_X1 #() 
BUF_X1_180_ (
  .A({ S25957[1043] }),
  .Z({ w[1043] })
);
BUF_X1 #() 
BUF_X1_181_ (
  .A({ S25957[1044] }),
  .Z({ w[1044] })
);
BUF_X1 #() 
BUF_X1_182_ (
  .A({ S25957[1045] }),
  .Z({ w[1045] })
);
BUF_X1 #() 
BUF_X1_183_ (
  .A({ S25957[1046] }),
  .Z({ w[1046] })
);
BUF_X1 #() 
BUF_X1_184_ (
  .A({ S25957[1047] }),
  .Z({ w[1047] })
);
BUF_X1 #() 
BUF_X1_185_ (
  .A({ S25957[1048] }),
  .Z({ w[1048] })
);
BUF_X1 #() 
BUF_X1_186_ (
  .A({ S25957[1049] }),
  .Z({ w[1049] })
);
BUF_X1 #() 
BUF_X1_187_ (
  .A({ S25957[105] }),
  .Z({ w[105] })
);
BUF_X1 #() 
BUF_X1_188_ (
  .A({ S25957[1050] }),
  .Z({ w[1050] })
);
BUF_X1 #() 
BUF_X1_189_ (
  .A({ S25957[1051] }),
  .Z({ w[1051] })
);
BUF_X1 #() 
BUF_X1_190_ (
  .A({ S25957[1052] }),
  .Z({ w[1052] })
);
BUF_X1 #() 
BUF_X1_191_ (
  .A({ S25957[1053] }),
  .Z({ w[1053] })
);
BUF_X1 #() 
BUF_X1_192_ (
  .A({ S25957[1054] }),
  .Z({ w[1054] })
);
BUF_X1 #() 
BUF_X1_193_ (
  .A({ S25957[1055] }),
  .Z({ w[1055] })
);
BUF_X1 #() 
BUF_X1_194_ (
  .A({ S25957[1056] }),
  .Z({ w[1056] })
);
BUF_X1 #() 
BUF_X1_195_ (
  .A({ S25957[1057] }),
  .Z({ w[1057] })
);
BUF_X1 #() 
BUF_X1_196_ (
  .A({ S25957[1058] }),
  .Z({ w[1058] })
);
BUF_X1 #() 
BUF_X1_197_ (
  .A({ S25957[1059] }),
  .Z({ w[1059] })
);
BUF_X1 #() 
BUF_X1_198_ (
  .A({ S25957[106] }),
  .Z({ w[106] })
);
BUF_X1 #() 
BUF_X1_199_ (
  .A({ S25957[1060] }),
  .Z({ w[1060] })
);
BUF_X1 #() 
BUF_X1_200_ (
  .A({ S25957[1061] }),
  .Z({ w[1061] })
);
BUF_X1 #() 
BUF_X1_201_ (
  .A({ S25957[1062] }),
  .Z({ w[1062] })
);
BUF_X1 #() 
BUF_X1_202_ (
  .A({ S25957[1063] }),
  .Z({ w[1063] })
);
BUF_X1 #() 
BUF_X1_203_ (
  .A({ S25957[1064] }),
  .Z({ w[1064] })
);
BUF_X1 #() 
BUF_X1_204_ (
  .A({ S25957[1065] }),
  .Z({ w[1065] })
);
BUF_X1 #() 
BUF_X1_205_ (
  .A({ S25957[1066] }),
  .Z({ w[1066] })
);
BUF_X1 #() 
BUF_X1_206_ (
  .A({ S25957[1067] }),
  .Z({ w[1067] })
);
BUF_X1 #() 
BUF_X1_207_ (
  .A({ S25957[1068] }),
  .Z({ w[1068] })
);
BUF_X1 #() 
BUF_X1_208_ (
  .A({ S25957[1069] }),
  .Z({ w[1069] })
);
BUF_X1 #() 
BUF_X1_209_ (
  .A({ S25957[107] }),
  .Z({ w[107] })
);
BUF_X1 #() 
BUF_X1_210_ (
  .A({ S25957[1070] }),
  .Z({ w[1070] })
);
BUF_X1 #() 
BUF_X1_211_ (
  .A({ S25957[1071] }),
  .Z({ w[1071] })
);
BUF_X1 #() 
BUF_X1_212_ (
  .A({ S25957[1072] }),
  .Z({ w[1072] })
);
BUF_X1 #() 
BUF_X1_213_ (
  .A({ S25957[1073] }),
  .Z({ w[1073] })
);
BUF_X1 #() 
BUF_X1_214_ (
  .A({ S25957[1074] }),
  .Z({ w[1074] })
);
BUF_X1 #() 
BUF_X1_215_ (
  .A({ S25957[1075] }),
  .Z({ w[1075] })
);
BUF_X1 #() 
BUF_X1_216_ (
  .A({ S25957[1076] }),
  .Z({ w[1076] })
);
BUF_X1 #() 
BUF_X1_217_ (
  .A({ S25957[1077] }),
  .Z({ w[1077] })
);
BUF_X1 #() 
BUF_X1_218_ (
  .A({ S25957[1078] }),
  .Z({ w[1078] })
);
BUF_X1 #() 
BUF_X1_219_ (
  .A({ S25957[1079] }),
  .Z({ w[1079] })
);
BUF_X1 #() 
BUF_X1_220_ (
  .A({ S25957[108] }),
  .Z({ w[108] })
);
BUF_X1 #() 
BUF_X1_221_ (
  .A({ S25957[1080] }),
  .Z({ w[1080] })
);
BUF_X1 #() 
BUF_X1_222_ (
  .A({ S25957[1081] }),
  .Z({ w[1081] })
);
BUF_X1 #() 
BUF_X1_223_ (
  .A({ S25957[1082] }),
  .Z({ w[1082] })
);
BUF_X1 #() 
BUF_X1_224_ (
  .A({ S25957[1083] }),
  .Z({ w[1083] })
);
BUF_X1 #() 
BUF_X1_225_ (
  .A({ S25957[1084] }),
  .Z({ w[1084] })
);
BUF_X1 #() 
BUF_X1_226_ (
  .A({ S25957[1085] }),
  .Z({ w[1085] })
);
BUF_X1 #() 
BUF_X1_227_ (
  .A({ S25957[1086] }),
  .Z({ w[1086] })
);
BUF_X1 #() 
BUF_X1_228_ (
  .A({ S25957[1087] }),
  .Z({ w[1087] })
);
BUF_X1 #() 
BUF_X1_229_ (
  .A({ S25957[1088] }),
  .Z({ w[1088] })
);
BUF_X1 #() 
BUF_X1_230_ (
  .A({ S25957[1089] }),
  .Z({ w[1089] })
);
BUF_X1 #() 
BUF_X1_231_ (
  .A({ S25957[109] }),
  .Z({ w[109] })
);
BUF_X1 #() 
BUF_X1_232_ (
  .A({ S25957[1090] }),
  .Z({ w[1090] })
);
BUF_X1 #() 
BUF_X1_233_ (
  .A({ S25957[1091] }),
  .Z({ w[1091] })
);
BUF_X1 #() 
BUF_X1_234_ (
  .A({ S25957[1092] }),
  .Z({ w[1092] })
);
BUF_X1 #() 
BUF_X1_235_ (
  .A({ S25957[1093] }),
  .Z({ w[1093] })
);
BUF_X1 #() 
BUF_X1_236_ (
  .A({ S25957[1094] }),
  .Z({ w[1094] })
);
BUF_X1 #() 
BUF_X1_237_ (
  .A({ S25957[1095] }),
  .Z({ w[1095] })
);
BUF_X1 #() 
BUF_X1_238_ (
  .A({ S25957[1096] }),
  .Z({ w[1096] })
);
BUF_X1 #() 
BUF_X1_239_ (
  .A({ S25957[1097] }),
  .Z({ w[1097] })
);
BUF_X1 #() 
BUF_X1_240_ (
  .A({ S25957[1098] }),
  .Z({ w[1098] })
);
BUF_X1 #() 
BUF_X1_241_ (
  .A({ S25957[1099] }),
  .Z({ w[1099] })
);
BUF_X1 #() 
BUF_X1_242_ (
  .A({ S25957[11] }),
  .Z({ w[11] })
);
BUF_X1 #() 
BUF_X1_243_ (
  .A({ S25957[110] }),
  .Z({ w[110] })
);
BUF_X1 #() 
BUF_X1_244_ (
  .A({ S25957[1100] }),
  .Z({ w[1100] })
);
BUF_X1 #() 
BUF_X1_245_ (
  .A({ S25957[1101] }),
  .Z({ w[1101] })
);
BUF_X1 #() 
BUF_X1_246_ (
  .A({ S25957[1102] }),
  .Z({ w[1102] })
);
BUF_X1 #() 
BUF_X1_247_ (
  .A({ S25957[1103] }),
  .Z({ w[1103] })
);
BUF_X1 #() 
BUF_X1_248_ (
  .A({ S25957[1104] }),
  .Z({ w[1104] })
);
BUF_X1 #() 
BUF_X1_249_ (
  .A({ S25957[1105] }),
  .Z({ w[1105] })
);
BUF_X1 #() 
BUF_X1_250_ (
  .A({ S25957[1106] }),
  .Z({ w[1106] })
);
BUF_X1 #() 
BUF_X1_251_ (
  .A({ S25957[1107] }),
  .Z({ w[1107] })
);
BUF_X1 #() 
BUF_X1_252_ (
  .A({ S25957[1108] }),
  .Z({ w[1108] })
);
BUF_X1 #() 
BUF_X1_253_ (
  .A({ S25957[1109] }),
  .Z({ w[1109] })
);
BUF_X1 #() 
BUF_X1_254_ (
  .A({ S25957[111] }),
  .Z({ w[111] })
);
BUF_X1 #() 
BUF_X1_255_ (
  .A({ S25957[1110] }),
  .Z({ w[1110] })
);
BUF_X1 #() 
BUF_X1_256_ (
  .A({ S25957[1111] }),
  .Z({ w[1111] })
);
BUF_X1 #() 
BUF_X1_257_ (
  .A({ S25957[1112] }),
  .Z({ w[1112] })
);
BUF_X1 #() 
BUF_X1_258_ (
  .A({ S25957[1113] }),
  .Z({ w[1113] })
);
BUF_X1 #() 
BUF_X1_259_ (
  .A({ S25957[1114] }),
  .Z({ w[1114] })
);
BUF_X1 #() 
BUF_X1_260_ (
  .A({ S25957[1115] }),
  .Z({ w[1115] })
);
BUF_X1 #() 
BUF_X1_261_ (
  .A({ S25957[1116] }),
  .Z({ w[1116] })
);
BUF_X1 #() 
BUF_X1_262_ (
  .A({ S25957[1117] }),
  .Z({ w[1117] })
);
BUF_X1 #() 
BUF_X1_263_ (
  .A({ S25957[1118] }),
  .Z({ w[1118] })
);
BUF_X1 #() 
BUF_X1_264_ (
  .A({ S25957[1119] }),
  .Z({ w[1119] })
);
BUF_X1 #() 
BUF_X1_265_ (
  .A({ S25957[112] }),
  .Z({ w[112] })
);
BUF_X1 #() 
BUF_X1_266_ (
  .A({ S25957[1120] }),
  .Z({ w[1120] })
);
BUF_X1 #() 
BUF_X1_267_ (
  .A({ S25957[1121] }),
  .Z({ w[1121] })
);
BUF_X1 #() 
BUF_X1_268_ (
  .A({ S25957[1122] }),
  .Z({ w[1122] })
);
BUF_X1 #() 
BUF_X1_269_ (
  .A({ S25957[1123] }),
  .Z({ w[1123] })
);
BUF_X1 #() 
BUF_X1_270_ (
  .A({ S25957[1124] }),
  .Z({ w[1124] })
);
BUF_X1 #() 
BUF_X1_271_ (
  .A({ S25957[1125] }),
  .Z({ w[1125] })
);
BUF_X1 #() 
BUF_X1_272_ (
  .A({ S25957[1126] }),
  .Z({ w[1126] })
);
BUF_X1 #() 
BUF_X1_273_ (
  .A({ S25957[1127] }),
  .Z({ w[1127] })
);
BUF_X1 #() 
BUF_X1_274_ (
  .A({ S25957[1128] }),
  .Z({ w[1128] })
);
BUF_X1 #() 
BUF_X1_275_ (
  .A({ S25957[1129] }),
  .Z({ w[1129] })
);
BUF_X1 #() 
BUF_X1_276_ (
  .A({ S25957[113] }),
  .Z({ w[113] })
);
BUF_X1 #() 
BUF_X1_277_ (
  .A({ S25957[1130] }),
  .Z({ w[1130] })
);
BUF_X1 #() 
BUF_X1_278_ (
  .A({ S25957[1131] }),
  .Z({ w[1131] })
);
BUF_X1 #() 
BUF_X1_279_ (
  .A({ S25957[1132] }),
  .Z({ w[1132] })
);
BUF_X1 #() 
BUF_X1_280_ (
  .A({ S25957[1133] }),
  .Z({ w[1133] })
);
BUF_X1 #() 
BUF_X1_281_ (
  .A({ S25957[1134] }),
  .Z({ w[1134] })
);
BUF_X1 #() 
BUF_X1_282_ (
  .A({ S25957[1135] }),
  .Z({ w[1135] })
);
BUF_X1 #() 
BUF_X1_283_ (
  .A({ S25957[1136] }),
  .Z({ w[1136] })
);
BUF_X1 #() 
BUF_X1_284_ (
  .A({ S25957[1137] }),
  .Z({ w[1137] })
);
BUF_X1 #() 
BUF_X1_285_ (
  .A({ S25957[1138] }),
  .Z({ w[1138] })
);
BUF_X1 #() 
BUF_X1_286_ (
  .A({ S25957[1139] }),
  .Z({ w[1139] })
);
BUF_X1 #() 
BUF_X1_287_ (
  .A({ S25957[114] }),
  .Z({ w[114] })
);
BUF_X1 #() 
BUF_X1_288_ (
  .A({ S25957[1140] }),
  .Z({ w[1140] })
);
BUF_X1 #() 
BUF_X1_289_ (
  .A({ S25957[1141] }),
  .Z({ w[1141] })
);
BUF_X1 #() 
BUF_X1_290_ (
  .A({ S25957[1142] }),
  .Z({ w[1142] })
);
BUF_X1 #() 
BUF_X1_291_ (
  .A({ S25957[1143] }),
  .Z({ w[1143] })
);
BUF_X1 #() 
BUF_X1_292_ (
  .A({ S25957[1144] }),
  .Z({ w[1144] })
);
BUF_X1 #() 
BUF_X1_293_ (
  .A({ S25957[1145] }),
  .Z({ w[1145] })
);
BUF_X1 #() 
BUF_X1_294_ (
  .A({ S25957[1146] }),
  .Z({ w[1146] })
);
BUF_X1 #() 
BUF_X1_295_ (
  .A({ S25957[1147] }),
  .Z({ w[1147] })
);
BUF_X1 #() 
BUF_X1_296_ (
  .A({ S25957[1148] }),
  .Z({ w[1148] })
);
BUF_X1 #() 
BUF_X1_297_ (
  .A({ S25957[1149] }),
  .Z({ w[1149] })
);
BUF_X1 #() 
BUF_X1_298_ (
  .A({ S25957[115] }),
  .Z({ w[115] })
);
BUF_X1 #() 
BUF_X1_299_ (
  .A({ S25957[1150] }),
  .Z({ w[1150] })
);
BUF_X1 #() 
BUF_X1_300_ (
  .A({ S25957[1151] }),
  .Z({ w[1151] })
);
BUF_X1 #() 
BUF_X1_301_ (
  .A({ S25957[1152] }),
  .Z({ w[1152] })
);
BUF_X1 #() 
BUF_X1_302_ (
  .A({ S25957[1153] }),
  .Z({ w[1153] })
);
BUF_X1 #() 
BUF_X1_303_ (
  .A({ S25957[1154] }),
  .Z({ w[1154] })
);
BUF_X1 #() 
BUF_X1_304_ (
  .A({ S25957[1155] }),
  .Z({ w[1155] })
);
BUF_X1 #() 
BUF_X1_305_ (
  .A({ S25957[1156] }),
  .Z({ w[1156] })
);
BUF_X1 #() 
BUF_X1_306_ (
  .A({ S25957[1157] }),
  .Z({ w[1157] })
);
BUF_X1 #() 
BUF_X1_307_ (
  .A({ S25957[1158] }),
  .Z({ w[1158] })
);
BUF_X1 #() 
BUF_X1_308_ (
  .A({ S25957[1159] }),
  .Z({ w[1159] })
);
BUF_X1 #() 
BUF_X1_309_ (
  .A({ S25957[116] }),
  .Z({ w[116] })
);
BUF_X1 #() 
BUF_X1_310_ (
  .A({ S25957[1160] }),
  .Z({ w[1160] })
);
BUF_X1 #() 
BUF_X1_311_ (
  .A({ S25957[1161] }),
  .Z({ w[1161] })
);
BUF_X1 #() 
BUF_X1_312_ (
  .A({ S25957[1162] }),
  .Z({ w[1162] })
);
BUF_X1 #() 
BUF_X1_313_ (
  .A({ S25957[1163] }),
  .Z({ w[1163] })
);
BUF_X1 #() 
BUF_X1_314_ (
  .A({ S25957[1164] }),
  .Z({ w[1164] })
);
BUF_X1 #() 
BUF_X1_315_ (
  .A({ S25957[1165] }),
  .Z({ w[1165] })
);
BUF_X1 #() 
BUF_X1_316_ (
  .A({ S25957[1166] }),
  .Z({ w[1166] })
);
BUF_X1 #() 
BUF_X1_317_ (
  .A({ S25957[1167] }),
  .Z({ w[1167] })
);
BUF_X1 #() 
BUF_X1_318_ (
  .A({ S25957[1168] }),
  .Z({ w[1168] })
);
BUF_X1 #() 
BUF_X1_319_ (
  .A({ S25957[1169] }),
  .Z({ w[1169] })
);
BUF_X1 #() 
BUF_X1_320_ (
  .A({ S25957[117] }),
  .Z({ w[117] })
);
BUF_X1 #() 
BUF_X1_321_ (
  .A({ S25957[1170] }),
  .Z({ w[1170] })
);
BUF_X1 #() 
BUF_X1_322_ (
  .A({ S25957[1171] }),
  .Z({ w[1171] })
);
BUF_X1 #() 
BUF_X1_323_ (
  .A({ S25957[1172] }),
  .Z({ w[1172] })
);
BUF_X1 #() 
BUF_X1_324_ (
  .A({ S25957[1173] }),
  .Z({ w[1173] })
);
BUF_X1 #() 
BUF_X1_325_ (
  .A({ S25957[1174] }),
  .Z({ w[1174] })
);
BUF_X1 #() 
BUF_X1_326_ (
  .A({ S25957[1175] }),
  .Z({ w[1175] })
);
BUF_X1 #() 
BUF_X1_327_ (
  .A({ S25957[1176] }),
  .Z({ w[1176] })
);
BUF_X1 #() 
BUF_X1_328_ (
  .A({ S25957[1177] }),
  .Z({ w[1177] })
);
BUF_X1 #() 
BUF_X1_329_ (
  .A({ S25957[1178] }),
  .Z({ w[1178] })
);
BUF_X1 #() 
BUF_X1_330_ (
  .A({ S25957[1179] }),
  .Z({ w[1179] })
);
BUF_X1 #() 
BUF_X1_331_ (
  .A({ S25957[118] }),
  .Z({ w[118] })
);
BUF_X1 #() 
BUF_X1_332_ (
  .A({ S25957[1180] }),
  .Z({ w[1180] })
);
BUF_X1 #() 
BUF_X1_333_ (
  .A({ S25957[1181] }),
  .Z({ w[1181] })
);
BUF_X1 #() 
BUF_X1_334_ (
  .A({ S25957[1182] }),
  .Z({ w[1182] })
);
BUF_X1 #() 
BUF_X1_335_ (
  .A({ S25957[1183] }),
  .Z({ w[1183] })
);
BUF_X1 #() 
BUF_X1_336_ (
  .A({ S25957[1184] }),
  .Z({ w[1184] })
);
BUF_X1 #() 
BUF_X1_337_ (
  .A({ S25957[1185] }),
  .Z({ w[1185] })
);
BUF_X1 #() 
BUF_X1_338_ (
  .A({ S25957[1186] }),
  .Z({ w[1186] })
);
BUF_X1 #() 
BUF_X1_339_ (
  .A({ S25957[1187] }),
  .Z({ w[1187] })
);
BUF_X1 #() 
BUF_X1_340_ (
  .A({ S25957[1188] }),
  .Z({ w[1188] })
);
BUF_X1 #() 
BUF_X1_341_ (
  .A({ S25957[1189] }),
  .Z({ w[1189] })
);
BUF_X1 #() 
BUF_X1_342_ (
  .A({ S25957[119] }),
  .Z({ w[119] })
);
BUF_X1 #() 
BUF_X1_343_ (
  .A({ S25957[1190] }),
  .Z({ w[1190] })
);
BUF_X1 #() 
BUF_X1_344_ (
  .A({ S25957[1191] }),
  .Z({ w[1191] })
);
BUF_X1 #() 
BUF_X1_345_ (
  .A({ S25957[1192] }),
  .Z({ w[1192] })
);
BUF_X1 #() 
BUF_X1_346_ (
  .A({ S25957[1193] }),
  .Z({ w[1193] })
);
BUF_X1 #() 
BUF_X1_347_ (
  .A({ S25957[1194] }),
  .Z({ w[1194] })
);
BUF_X1 #() 
BUF_X1_348_ (
  .A({ S25957[1195] }),
  .Z({ w[1195] })
);
BUF_X1 #() 
BUF_X1_349_ (
  .A({ S25957[1196] }),
  .Z({ w[1196] })
);
BUF_X1 #() 
BUF_X1_350_ (
  .A({ S25957[1197] }),
  .Z({ w[1197] })
);
BUF_X1 #() 
BUF_X1_351_ (
  .A({ S25957[1198] }),
  .Z({ w[1198] })
);
BUF_X1 #() 
BUF_X1_352_ (
  .A({ S25957[1199] }),
  .Z({ w[1199] })
);
BUF_X1 #() 
BUF_X1_353_ (
  .A({ S25957[12] }),
  .Z({ w[12] })
);
BUF_X1 #() 
BUF_X1_354_ (
  .A({ S25957[120] }),
  .Z({ w[120] })
);
BUF_X1 #() 
BUF_X1_355_ (
  .A({ S25957[1200] }),
  .Z({ w[1200] })
);
BUF_X1 #() 
BUF_X1_356_ (
  .A({ S25957[1201] }),
  .Z({ w[1201] })
);
BUF_X1 #() 
BUF_X1_357_ (
  .A({ S25957[1202] }),
  .Z({ w[1202] })
);
BUF_X1 #() 
BUF_X1_358_ (
  .A({ S25957[1203] }),
  .Z({ w[1203] })
);
BUF_X1 #() 
BUF_X1_359_ (
  .A({ S25957[1204] }),
  .Z({ w[1204] })
);
BUF_X1 #() 
BUF_X1_360_ (
  .A({ S25957[1205] }),
  .Z({ w[1205] })
);
BUF_X1 #() 
BUF_X1_361_ (
  .A({ S25957[1206] }),
  .Z({ w[1206] })
);
BUF_X1 #() 
BUF_X1_362_ (
  .A({ S25957[1207] }),
  .Z({ w[1207] })
);
BUF_X1 #() 
BUF_X1_363_ (
  .A({ S25957[1208] }),
  .Z({ w[1208] })
);
BUF_X1 #() 
BUF_X1_364_ (
  .A({ S25957[1209] }),
  .Z({ w[1209] })
);
BUF_X1 #() 
BUF_X1_365_ (
  .A({ S25957[121] }),
  .Z({ w[121] })
);
BUF_X1 #() 
BUF_X1_366_ (
  .A({ S25957[1210] }),
  .Z({ w[1210] })
);
BUF_X1 #() 
BUF_X1_367_ (
  .A({ S25957[1211] }),
  .Z({ w[1211] })
);
BUF_X1 #() 
BUF_X1_368_ (
  .A({ S25957[1212] }),
  .Z({ w[1212] })
);
BUF_X1 #() 
BUF_X1_369_ (
  .A({ S25957[1213] }),
  .Z({ w[1213] })
);
BUF_X1 #() 
BUF_X1_370_ (
  .A({ S25957[1214] }),
  .Z({ w[1214] })
);
BUF_X1 #() 
BUF_X1_371_ (
  .A({ S25957[1215] }),
  .Z({ w[1215] })
);
BUF_X1 #() 
BUF_X1_372_ (
  .A({ S25957[1216] }),
  .Z({ w[1216] })
);
BUF_X1 #() 
BUF_X1_373_ (
  .A({ S25957[1217] }),
  .Z({ w[1217] })
);
BUF_X1 #() 
BUF_X1_374_ (
  .A({ S25957[1218] }),
  .Z({ w[1218] })
);
BUF_X1 #() 
BUF_X1_375_ (
  .A({ S25957[1219] }),
  .Z({ w[1219] })
);
BUF_X1 #() 
BUF_X1_376_ (
  .A({ S25957[122] }),
  .Z({ w[122] })
);
BUF_X1 #() 
BUF_X1_377_ (
  .A({ S25957[1220] }),
  .Z({ w[1220] })
);
BUF_X1 #() 
BUF_X1_378_ (
  .A({ S25957[1221] }),
  .Z({ w[1221] })
);
BUF_X1 #() 
BUF_X1_379_ (
  .A({ S25957[1222] }),
  .Z({ w[1222] })
);
BUF_X1 #() 
BUF_X1_380_ (
  .A({ S25957[1223] }),
  .Z({ w[1223] })
);
BUF_X1 #() 
BUF_X1_381_ (
  .A({ S25957[1224] }),
  .Z({ w[1224] })
);
BUF_X1 #() 
BUF_X1_382_ (
  .A({ S25957[1225] }),
  .Z({ w[1225] })
);
BUF_X1 #() 
BUF_X1_383_ (
  .A({ S25957[1226] }),
  .Z({ w[1226] })
);
BUF_X1 #() 
BUF_X1_384_ (
  .A({ S25957[1227] }),
  .Z({ w[1227] })
);
BUF_X1 #() 
BUF_X1_385_ (
  .A({ S25957[1228] }),
  .Z({ w[1228] })
);
BUF_X1 #() 
BUF_X1_386_ (
  .A({ S25957[1229] }),
  .Z({ w[1229] })
);
BUF_X1 #() 
BUF_X1_387_ (
  .A({ S25957[123] }),
  .Z({ w[123] })
);
BUF_X1 #() 
BUF_X1_388_ (
  .A({ S25957[1230] }),
  .Z({ w[1230] })
);
BUF_X1 #() 
BUF_X1_389_ (
  .A({ S25957[1231] }),
  .Z({ w[1231] })
);
BUF_X1 #() 
BUF_X1_390_ (
  .A({ S25957[1232] }),
  .Z({ w[1232] })
);
BUF_X1 #() 
BUF_X1_391_ (
  .A({ S25957[1233] }),
  .Z({ w[1233] })
);
BUF_X1 #() 
BUF_X1_392_ (
  .A({ S25957[1234] }),
  .Z({ w[1234] })
);
BUF_X1 #() 
BUF_X1_393_ (
  .A({ S25957[1235] }),
  .Z({ w[1235] })
);
BUF_X1 #() 
BUF_X1_394_ (
  .A({ S25957[1236] }),
  .Z({ w[1236] })
);
BUF_X1 #() 
BUF_X1_395_ (
  .A({ S25957[1237] }),
  .Z({ w[1237] })
);
BUF_X1 #() 
BUF_X1_396_ (
  .A({ S25957[1238] }),
  .Z({ w[1238] })
);
BUF_X1 #() 
BUF_X1_397_ (
  .A({ S25957[1239] }),
  .Z({ w[1239] })
);
BUF_X1 #() 
BUF_X1_398_ (
  .A({ S25957[124] }),
  .Z({ w[124] })
);
BUF_X1 #() 
BUF_X1_399_ (
  .A({ S25957[1240] }),
  .Z({ w[1240] })
);
BUF_X1 #() 
BUF_X1_400_ (
  .A({ S25957[1241] }),
  .Z({ w[1241] })
);
BUF_X1 #() 
BUF_X1_401_ (
  .A({ S25957[1242] }),
  .Z({ w[1242] })
);
BUF_X1 #() 
BUF_X1_402_ (
  .A({ S25957[1243] }),
  .Z({ w[1243] })
);
BUF_X1 #() 
BUF_X1_403_ (
  .A({ S25957[1244] }),
  .Z({ w[1244] })
);
BUF_X1 #() 
BUF_X1_404_ (
  .A({ S25957[1245] }),
  .Z({ w[1245] })
);
BUF_X1 #() 
BUF_X1_405_ (
  .A({ S25957[1246] }),
  .Z({ w[1246] })
);
BUF_X1 #() 
BUF_X1_406_ (
  .A({ S25957[1247] }),
  .Z({ w[1247] })
);
BUF_X1 #() 
BUF_X1_407_ (
  .A({ S25957[1248] }),
  .Z({ w[1248] })
);
BUF_X1 #() 
BUF_X1_408_ (
  .A({ S25957[1249] }),
  .Z({ w[1249] })
);
BUF_X1 #() 
BUF_X1_409_ (
  .A({ S25957[125] }),
  .Z({ w[125] })
);
BUF_X1 #() 
BUF_X1_410_ (
  .A({ S25957[1250] }),
  .Z({ w[1250] })
);
BUF_X1 #() 
BUF_X1_411_ (
  .A({ S25957[1251] }),
  .Z({ w[1251] })
);
BUF_X1 #() 
BUF_X1_412_ (
  .A({ S25957[1252] }),
  .Z({ w[1252] })
);
BUF_X1 #() 
BUF_X1_413_ (
  .A({ S25957[1253] }),
  .Z({ w[1253] })
);
BUF_X1 #() 
BUF_X1_414_ (
  .A({ S25957[1254] }),
  .Z({ w[1254] })
);
BUF_X1 #() 
BUF_X1_415_ (
  .A({ S25957[1255] }),
  .Z({ w[1255] })
);
BUF_X1 #() 
BUF_X1_416_ (
  .A({ S25957[1256] }),
  .Z({ w[1256] })
);
BUF_X1 #() 
BUF_X1_417_ (
  .A({ S25957[1257] }),
  .Z({ w[1257] })
);
BUF_X1 #() 
BUF_X1_418_ (
  .A({ S25957[1258] }),
  .Z({ w[1258] })
);
BUF_X1 #() 
BUF_X1_419_ (
  .A({ S25957[1259] }),
  .Z({ w[1259] })
);
BUF_X1 #() 
BUF_X1_420_ (
  .A({ S25957[126] }),
  .Z({ w[126] })
);
BUF_X1 #() 
BUF_X1_421_ (
  .A({ S25957[1260] }),
  .Z({ w[1260] })
);
BUF_X1 #() 
BUF_X1_422_ (
  .A({ S25957[1261] }),
  .Z({ w[1261] })
);
BUF_X1 #() 
BUF_X1_423_ (
  .A({ S25957[1262] }),
  .Z({ w[1262] })
);
BUF_X1 #() 
BUF_X1_424_ (
  .A({ S25957[1263] }),
  .Z({ w[1263] })
);
BUF_X1 #() 
BUF_X1_425_ (
  .A({ S25957[1264] }),
  .Z({ w[1264] })
);
BUF_X1 #() 
BUF_X1_426_ (
  .A({ S25957[1265] }),
  .Z({ w[1265] })
);
BUF_X1 #() 
BUF_X1_427_ (
  .A({ S25957[1266] }),
  .Z({ w[1266] })
);
BUF_X1 #() 
BUF_X1_428_ (
  .A({ S25957[1267] }),
  .Z({ w[1267] })
);
BUF_X1 #() 
BUF_X1_429_ (
  .A({ S25957[1268] }),
  .Z({ w[1268] })
);
BUF_X1 #() 
BUF_X1_430_ (
  .A({ S25957[1269] }),
  .Z({ w[1269] })
);
BUF_X1 #() 
BUF_X1_431_ (
  .A({ S25957[127] }),
  .Z({ w[127] })
);
BUF_X1 #() 
BUF_X1_432_ (
  .A({ S25957[1270] }),
  .Z({ w[1270] })
);
BUF_X1 #() 
BUF_X1_433_ (
  .A({ S25957[1271] }),
  .Z({ w[1271] })
);
BUF_X1 #() 
BUF_X1_434_ (
  .A({ S25957[1272] }),
  .Z({ w[1272] })
);
BUF_X1 #() 
BUF_X1_435_ (
  .A({ S25957[1273] }),
  .Z({ w[1273] })
);
BUF_X1 #() 
BUF_X1_436_ (
  .A({ S25957[1274] }),
  .Z({ w[1274] })
);
BUF_X1 #() 
BUF_X1_437_ (
  .A({ S25957[1275] }),
  .Z({ w[1275] })
);
BUF_X1 #() 
BUF_X1_438_ (
  .A({ S25957[1276] }),
  .Z({ w[1276] })
);
BUF_X1 #() 
BUF_X1_439_ (
  .A({ S25957[1277] }),
  .Z({ w[1277] })
);
BUF_X1 #() 
BUF_X1_440_ (
  .A({ S25957[1278] }),
  .Z({ w[1278] })
);
BUF_X1 #() 
BUF_X1_441_ (
  .A({ S25957[1279] }),
  .Z({ w[1279] })
);
BUF_X1 #() 
BUF_X1_442_ (
  .A({ S25957[128] }),
  .Z({ w[128] })
);
BUF_X1 #() 
BUF_X1_443_ (
  .A({ S25957[129] }),
  .Z({ w[129] })
);
BUF_X1 #() 
BUF_X1_444_ (
  .A({ S25957[13] }),
  .Z({ w[13] })
);
BUF_X1 #() 
BUF_X1_445_ (
  .A({ S25957[130] }),
  .Z({ w[130] })
);
BUF_X1 #() 
BUF_X1_446_ (
  .A({ S25957[131] }),
  .Z({ w[131] })
);
BUF_X1 #() 
BUF_X1_447_ (
  .A({ S25957[132] }),
  .Z({ w[132] })
);
BUF_X1 #() 
BUF_X1_448_ (
  .A({ S25957[133] }),
  .Z({ w[133] })
);
BUF_X1 #() 
BUF_X1_449_ (
  .A({ S25957[134] }),
  .Z({ w[134] })
);
BUF_X1 #() 
BUF_X1_450_ (
  .A({ S25957[135] }),
  .Z({ w[135] })
);
BUF_X1 #() 
BUF_X1_451_ (
  .A({ S25957[136] }),
  .Z({ w[136] })
);
BUF_X1 #() 
BUF_X1_452_ (
  .A({ S25957[137] }),
  .Z({ w[137] })
);
BUF_X1 #() 
BUF_X1_453_ (
  .A({ S25957[138] }),
  .Z({ w[138] })
);
BUF_X1 #() 
BUF_X1_454_ (
  .A({ S25957[139] }),
  .Z({ w[139] })
);
BUF_X1 #() 
BUF_X1_455_ (
  .A({ S25957[14] }),
  .Z({ w[14] })
);
BUF_X1 #() 
BUF_X1_456_ (
  .A({ S25957[140] }),
  .Z({ w[140] })
);
BUF_X1 #() 
BUF_X1_457_ (
  .A({ S25957[141] }),
  .Z({ w[141] })
);
BUF_X1 #() 
BUF_X1_458_ (
  .A({ S25957[142] }),
  .Z({ w[142] })
);
BUF_X1 #() 
BUF_X1_459_ (
  .A({ S25957[143] }),
  .Z({ w[143] })
);
BUF_X1 #() 
BUF_X1_460_ (
  .A({ S25957[144] }),
  .Z({ w[144] })
);
BUF_X1 #() 
BUF_X1_461_ (
  .A({ S25957[145] }),
  .Z({ w[145] })
);
BUF_X1 #() 
BUF_X1_462_ (
  .A({ S25957[146] }),
  .Z({ w[146] })
);
BUF_X1 #() 
BUF_X1_463_ (
  .A({ S25957[147] }),
  .Z({ w[147] })
);
BUF_X1 #() 
BUF_X1_464_ (
  .A({ S25957[148] }),
  .Z({ w[148] })
);
BUF_X1 #() 
BUF_X1_465_ (
  .A({ S25957[149] }),
  .Z({ w[149] })
);
BUF_X1 #() 
BUF_X1_466_ (
  .A({ S25957[15] }),
  .Z({ w[15] })
);
BUF_X1 #() 
BUF_X1_467_ (
  .A({ S25957[150] }),
  .Z({ w[150] })
);
BUF_X1 #() 
BUF_X1_468_ (
  .A({ S25957[151] }),
  .Z({ w[151] })
);
BUF_X1 #() 
BUF_X1_469_ (
  .A({ S25957[152] }),
  .Z({ w[152] })
);
BUF_X1 #() 
BUF_X1_470_ (
  .A({ S25957[153] }),
  .Z({ w[153] })
);
BUF_X1 #() 
BUF_X1_471_ (
  .A({ S25957[154] }),
  .Z({ w[154] })
);
BUF_X1 #() 
BUF_X1_472_ (
  .A({ S25957[155] }),
  .Z({ w[155] })
);
BUF_X1 #() 
BUF_X1_473_ (
  .A({ S25957[156] }),
  .Z({ w[156] })
);
BUF_X1 #() 
BUF_X1_474_ (
  .A({ S25957[157] }),
  .Z({ w[157] })
);
BUF_X1 #() 
BUF_X1_475_ (
  .A({ S25957[158] }),
  .Z({ w[158] })
);
BUF_X1 #() 
BUF_X1_476_ (
  .A({ S25957[159] }),
  .Z({ w[159] })
);
BUF_X1 #() 
BUF_X1_477_ (
  .A({ S25957[16] }),
  .Z({ w[16] })
);
BUF_X1 #() 
BUF_X1_478_ (
  .A({ S25957[160] }),
  .Z({ w[160] })
);
BUF_X1 #() 
BUF_X1_479_ (
  .A({ S25957[161] }),
  .Z({ w[161] })
);
BUF_X1 #() 
BUF_X1_480_ (
  .A({ S25957[162] }),
  .Z({ w[162] })
);
BUF_X1 #() 
BUF_X1_481_ (
  .A({ S25957[163] }),
  .Z({ w[163] })
);
BUF_X1 #() 
BUF_X1_482_ (
  .A({ S25957[164] }),
  .Z({ w[164] })
);
BUF_X1 #() 
BUF_X1_483_ (
  .A({ S25957[165] }),
  .Z({ w[165] })
);
BUF_X1 #() 
BUF_X1_484_ (
  .A({ S25957[166] }),
  .Z({ w[166] })
);
BUF_X1 #() 
BUF_X1_485_ (
  .A({ S25957[167] }),
  .Z({ w[167] })
);
BUF_X1 #() 
BUF_X1_486_ (
  .A({ S25957[168] }),
  .Z({ w[168] })
);
BUF_X1 #() 
BUF_X1_487_ (
  .A({ S25957[169] }),
  .Z({ w[169] })
);
BUF_X1 #() 
BUF_X1_488_ (
  .A({ S25957[17] }),
  .Z({ w[17] })
);
BUF_X1 #() 
BUF_X1_489_ (
  .A({ S25957[170] }),
  .Z({ w[170] })
);
BUF_X1 #() 
BUF_X1_490_ (
  .A({ S25957[171] }),
  .Z({ w[171] })
);
BUF_X1 #() 
BUF_X1_491_ (
  .A({ S25957[172] }),
  .Z({ w[172] })
);
BUF_X1 #() 
BUF_X1_492_ (
  .A({ S25957[173] }),
  .Z({ w[173] })
);
BUF_X1 #() 
BUF_X1_493_ (
  .A({ S25957[174] }),
  .Z({ w[174] })
);
BUF_X1 #() 
BUF_X1_494_ (
  .A({ S25957[175] }),
  .Z({ w[175] })
);
BUF_X1 #() 
BUF_X1_495_ (
  .A({ S25957[176] }),
  .Z({ w[176] })
);
BUF_X1 #() 
BUF_X1_496_ (
  .A({ S25957[177] }),
  .Z({ w[177] })
);
BUF_X1 #() 
BUF_X1_497_ (
  .A({ S25957[178] }),
  .Z({ w[178] })
);
BUF_X1 #() 
BUF_X1_498_ (
  .A({ S25957[179] }),
  .Z({ w[179] })
);
BUF_X1 #() 
BUF_X1_499_ (
  .A({ S25957[18] }),
  .Z({ w[18] })
);
BUF_X1 #() 
BUF_X1_500_ (
  .A({ S25957[180] }),
  .Z({ w[180] })
);
BUF_X1 #() 
BUF_X1_501_ (
  .A({ S25957[181] }),
  .Z({ w[181] })
);
BUF_X1 #() 
BUF_X1_502_ (
  .A({ S25957[182] }),
  .Z({ w[182] })
);
BUF_X1 #() 
BUF_X1_503_ (
  .A({ S25957[183] }),
  .Z({ w[183] })
);
BUF_X1 #() 
BUF_X1_504_ (
  .A({ S25957[184] }),
  .Z({ w[184] })
);
BUF_X1 #() 
BUF_X1_505_ (
  .A({ S25957[185] }),
  .Z({ w[185] })
);
BUF_X1 #() 
BUF_X1_506_ (
  .A({ S25957[186] }),
  .Z({ w[186] })
);
BUF_X1 #() 
BUF_X1_507_ (
  .A({ S25957[187] }),
  .Z({ w[187] })
);
BUF_X1 #() 
BUF_X1_508_ (
  .A({ S25957[188] }),
  .Z({ w[188] })
);
BUF_X1 #() 
BUF_X1_509_ (
  .A({ S25957[189] }),
  .Z({ w[189] })
);
BUF_X1 #() 
BUF_X1_510_ (
  .A({ S25957[19] }),
  .Z({ w[19] })
);
BUF_X1 #() 
BUF_X1_511_ (
  .A({ S25957[190] }),
  .Z({ w[190] })
);
BUF_X1 #() 
BUF_X1_512_ (
  .A({ S25957[191] }),
  .Z({ w[191] })
);
BUF_X1 #() 
BUF_X1_513_ (
  .A({ S25957[192] }),
  .Z({ w[192] })
);
BUF_X1 #() 
BUF_X1_514_ (
  .A({ S25957[193] }),
  .Z({ w[193] })
);
BUF_X1 #() 
BUF_X1_515_ (
  .A({ S25957[194] }),
  .Z({ w[194] })
);
BUF_X1 #() 
BUF_X1_516_ (
  .A({ S25957[195] }),
  .Z({ w[195] })
);
BUF_X1 #() 
BUF_X1_517_ (
  .A({ S25957[196] }),
  .Z({ w[196] })
);
BUF_X1 #() 
BUF_X1_518_ (
  .A({ S25957[197] }),
  .Z({ w[197] })
);
BUF_X1 #() 
BUF_X1_519_ (
  .A({ S25957[198] }),
  .Z({ w[198] })
);
BUF_X1 #() 
BUF_X1_520_ (
  .A({ S25957[199] }),
  .Z({ w[199] })
);
BUF_X1 #() 
BUF_X1_521_ (
  .A({ S25957[2] }),
  .Z({ w[2] })
);
BUF_X1 #() 
BUF_X1_522_ (
  .A({ S25957[20] }),
  .Z({ w[20] })
);
BUF_X1 #() 
BUF_X1_523_ (
  .A({ S25957[200] }),
  .Z({ w[200] })
);
BUF_X1 #() 
BUF_X1_524_ (
  .A({ S25957[201] }),
  .Z({ w[201] })
);
BUF_X1 #() 
BUF_X1_525_ (
  .A({ S25957[202] }),
  .Z({ w[202] })
);
BUF_X1 #() 
BUF_X1_526_ (
  .A({ S25957[203] }),
  .Z({ w[203] })
);
BUF_X1 #() 
BUF_X1_527_ (
  .A({ S25957[204] }),
  .Z({ w[204] })
);
BUF_X1 #() 
BUF_X1_528_ (
  .A({ S25957[205] }),
  .Z({ w[205] })
);
BUF_X1 #() 
BUF_X1_529_ (
  .A({ S25957[206] }),
  .Z({ w[206] })
);
BUF_X1 #() 
BUF_X1_530_ (
  .A({ S25957[207] }),
  .Z({ w[207] })
);
BUF_X1 #() 
BUF_X1_531_ (
  .A({ S25957[208] }),
  .Z({ w[208] })
);
BUF_X1 #() 
BUF_X1_532_ (
  .A({ S25957[209] }),
  .Z({ w[209] })
);
BUF_X1 #() 
BUF_X1_533_ (
  .A({ S25957[21] }),
  .Z({ w[21] })
);
BUF_X1 #() 
BUF_X1_534_ (
  .A({ S25957[210] }),
  .Z({ w[210] })
);
BUF_X1 #() 
BUF_X1_535_ (
  .A({ S25957[211] }),
  .Z({ w[211] })
);
BUF_X1 #() 
BUF_X1_536_ (
  .A({ S25957[212] }),
  .Z({ w[212] })
);
BUF_X1 #() 
BUF_X1_537_ (
  .A({ S25957[213] }),
  .Z({ w[213] })
);
BUF_X1 #() 
BUF_X1_538_ (
  .A({ S25957[214] }),
  .Z({ w[214] })
);
BUF_X1 #() 
BUF_X1_539_ (
  .A({ S25957[215] }),
  .Z({ w[215] })
);
BUF_X1 #() 
BUF_X1_540_ (
  .A({ S25957[216] }),
  .Z({ w[216] })
);
BUF_X1 #() 
BUF_X1_541_ (
  .A({ S25957[217] }),
  .Z({ w[217] })
);
BUF_X1 #() 
BUF_X1_542_ (
  .A({ S25957[218] }),
  .Z({ w[218] })
);
BUF_X1 #() 
BUF_X1_543_ (
  .A({ S25957[219] }),
  .Z({ w[219] })
);
BUF_X1 #() 
BUF_X1_544_ (
  .A({ S25957[22] }),
  .Z({ w[22] })
);
BUF_X1 #() 
BUF_X1_545_ (
  .A({ S25957[220] }),
  .Z({ w[220] })
);
BUF_X1 #() 
BUF_X1_546_ (
  .A({ S25957[221] }),
  .Z({ w[221] })
);
BUF_X1 #() 
BUF_X1_547_ (
  .A({ S25957[222] }),
  .Z({ w[222] })
);
BUF_X1 #() 
BUF_X1_548_ (
  .A({ S25957[223] }),
  .Z({ w[223] })
);
BUF_X1 #() 
BUF_X1_549_ (
  .A({ S25957[224] }),
  .Z({ w[224] })
);
BUF_X1 #() 
BUF_X1_550_ (
  .A({ S25957[225] }),
  .Z({ w[225] })
);
BUF_X1 #() 
BUF_X1_551_ (
  .A({ S25957[226] }),
  .Z({ w[226] })
);
BUF_X1 #() 
BUF_X1_552_ (
  .A({ S25957[227] }),
  .Z({ w[227] })
);
BUF_X1 #() 
BUF_X1_553_ (
  .A({ S25957[228] }),
  .Z({ w[228] })
);
BUF_X1 #() 
BUF_X1_554_ (
  .A({ S25957[229] }),
  .Z({ w[229] })
);
BUF_X1 #() 
BUF_X1_555_ (
  .A({ S25957[23] }),
  .Z({ w[23] })
);
BUF_X1 #() 
BUF_X1_556_ (
  .A({ S25957[230] }),
  .Z({ w[230] })
);
BUF_X1 #() 
BUF_X1_557_ (
  .A({ S25957[231] }),
  .Z({ w[231] })
);
BUF_X1 #() 
BUF_X1_558_ (
  .A({ S25957[232] }),
  .Z({ w[232] })
);
BUF_X1 #() 
BUF_X1_559_ (
  .A({ S25957[233] }),
  .Z({ w[233] })
);
BUF_X1 #() 
BUF_X1_560_ (
  .A({ S25957[234] }),
  .Z({ w[234] })
);
BUF_X1 #() 
BUF_X1_561_ (
  .A({ S25957[235] }),
  .Z({ w[235] })
);
BUF_X1 #() 
BUF_X1_562_ (
  .A({ S25957[236] }),
  .Z({ w[236] })
);
BUF_X1 #() 
BUF_X1_563_ (
  .A({ S25957[237] }),
  .Z({ w[237] })
);
BUF_X1 #() 
BUF_X1_564_ (
  .A({ S25957[238] }),
  .Z({ w[238] })
);
BUF_X1 #() 
BUF_X1_565_ (
  .A({ S25957[239] }),
  .Z({ w[239] })
);
BUF_X1 #() 
BUF_X1_566_ (
  .A({ S25957[24] }),
  .Z({ w[24] })
);
BUF_X1 #() 
BUF_X1_567_ (
  .A({ S25957[240] }),
  .Z({ w[240] })
);
BUF_X1 #() 
BUF_X1_568_ (
  .A({ S25957[241] }),
  .Z({ w[241] })
);
BUF_X1 #() 
BUF_X1_569_ (
  .A({ S25957[242] }),
  .Z({ w[242] })
);
BUF_X1 #() 
BUF_X1_570_ (
  .A({ S25957[243] }),
  .Z({ w[243] })
);
BUF_X1 #() 
BUF_X1_571_ (
  .A({ S25957[244] }),
  .Z({ w[244] })
);
BUF_X1 #() 
BUF_X1_572_ (
  .A({ S25957[245] }),
  .Z({ w[245] })
);
BUF_X1 #() 
BUF_X1_573_ (
  .A({ S25957[246] }),
  .Z({ w[246] })
);
BUF_X1 #() 
BUF_X1_574_ (
  .A({ S25957[247] }),
  .Z({ w[247] })
);
BUF_X1 #() 
BUF_X1_575_ (
  .A({ S25957[248] }),
  .Z({ w[248] })
);
BUF_X1 #() 
BUF_X1_576_ (
  .A({ S25957[249] }),
  .Z({ w[249] })
);
BUF_X1 #() 
BUF_X1_577_ (
  .A({ S25957[25] }),
  .Z({ w[25] })
);
BUF_X1 #() 
BUF_X1_578_ (
  .A({ S25957[250] }),
  .Z({ w[250] })
);
BUF_X1 #() 
BUF_X1_579_ (
  .A({ S25957[251] }),
  .Z({ w[251] })
);
BUF_X1 #() 
BUF_X1_580_ (
  .A({ S25957[252] }),
  .Z({ w[252] })
);
BUF_X1 #() 
BUF_X1_581_ (
  .A({ S25957[253] }),
  .Z({ w[253] })
);
BUF_X1 #() 
BUF_X1_582_ (
  .A({ S25957[254] }),
  .Z({ w[254] })
);
BUF_X1 #() 
BUF_X1_583_ (
  .A({ S25957[255] }),
  .Z({ w[255] })
);
BUF_X1 #() 
BUF_X1_584_ (
  .A({ S25957[256] }),
  .Z({ w[256] })
);
BUF_X1 #() 
BUF_X1_585_ (
  .A({ S25957[257] }),
  .Z({ w[257] })
);
BUF_X1 #() 
BUF_X1_586_ (
  .A({ S25957[258] }),
  .Z({ w[258] })
);
BUF_X1 #() 
BUF_X1_587_ (
  .A({ S25957[259] }),
  .Z({ w[259] })
);
BUF_X1 #() 
BUF_X1_588_ (
  .A({ S25957[26] }),
  .Z({ w[26] })
);
BUF_X1 #() 
BUF_X1_589_ (
  .A({ S25957[260] }),
  .Z({ w[260] })
);
BUF_X1 #() 
BUF_X1_590_ (
  .A({ S25957[261] }),
  .Z({ w[261] })
);
BUF_X1 #() 
BUF_X1_591_ (
  .A({ S25957[262] }),
  .Z({ w[262] })
);
BUF_X1 #() 
BUF_X1_592_ (
  .A({ S25957[263] }),
  .Z({ w[263] })
);
BUF_X1 #() 
BUF_X1_593_ (
  .A({ S25957[264] }),
  .Z({ w[264] })
);
BUF_X1 #() 
BUF_X1_594_ (
  .A({ S25957[265] }),
  .Z({ w[265] })
);
BUF_X1 #() 
BUF_X1_595_ (
  .A({ S25957[266] }),
  .Z({ w[266] })
);
BUF_X1 #() 
BUF_X1_596_ (
  .A({ S25957[267] }),
  .Z({ w[267] })
);
BUF_X1 #() 
BUF_X1_597_ (
  .A({ S25957[268] }),
  .Z({ w[268] })
);
BUF_X1 #() 
BUF_X1_598_ (
  .A({ S25957[269] }),
  .Z({ w[269] })
);
BUF_X1 #() 
BUF_X1_599_ (
  .A({ S25957[27] }),
  .Z({ w[27] })
);
BUF_X1 #() 
BUF_X1_600_ (
  .A({ S25957[270] }),
  .Z({ w[270] })
);
BUF_X1 #() 
BUF_X1_601_ (
  .A({ S25957[271] }),
  .Z({ w[271] })
);
BUF_X1 #() 
BUF_X1_602_ (
  .A({ S25957[272] }),
  .Z({ w[272] })
);
BUF_X1 #() 
BUF_X1_603_ (
  .A({ S25957[273] }),
  .Z({ w[273] })
);
BUF_X1 #() 
BUF_X1_604_ (
  .A({ S25957[274] }),
  .Z({ w[274] })
);
BUF_X1 #() 
BUF_X1_605_ (
  .A({ S25957[275] }),
  .Z({ w[275] })
);
BUF_X1 #() 
BUF_X1_606_ (
  .A({ S25957[276] }),
  .Z({ w[276] })
);
BUF_X1 #() 
BUF_X1_607_ (
  .A({ S25957[277] }),
  .Z({ w[277] })
);
BUF_X1 #() 
BUF_X1_608_ (
  .A({ S25957[278] }),
  .Z({ w[278] })
);
BUF_X1 #() 
BUF_X1_609_ (
  .A({ S25957[279] }),
  .Z({ w[279] })
);
BUF_X1 #() 
BUF_X1_610_ (
  .A({ S25957[28] }),
  .Z({ w[28] })
);
BUF_X1 #() 
BUF_X1_611_ (
  .A({ S25957[280] }),
  .Z({ w[280] })
);
BUF_X1 #() 
BUF_X1_612_ (
  .A({ S25957[281] }),
  .Z({ w[281] })
);
BUF_X1 #() 
BUF_X1_613_ (
  .A({ S25957[282] }),
  .Z({ w[282] })
);
BUF_X1 #() 
BUF_X1_614_ (
  .A({ S25957[283] }),
  .Z({ w[283] })
);
BUF_X1 #() 
BUF_X1_615_ (
  .A({ S25957[284] }),
  .Z({ w[284] })
);
BUF_X1 #() 
BUF_X1_616_ (
  .A({ S25957[285] }),
  .Z({ w[285] })
);
BUF_X1 #() 
BUF_X1_617_ (
  .A({ S25957[286] }),
  .Z({ w[286] })
);
BUF_X1 #() 
BUF_X1_618_ (
  .A({ S25957[287] }),
  .Z({ w[287] })
);
BUF_X1 #() 
BUF_X1_619_ (
  .A({ S25957[288] }),
  .Z({ w[288] })
);
BUF_X1 #() 
BUF_X1_620_ (
  .A({ S25957[289] }),
  .Z({ w[289] })
);
BUF_X1 #() 
BUF_X1_621_ (
  .A({ S25957[29] }),
  .Z({ w[29] })
);
BUF_X1 #() 
BUF_X1_622_ (
  .A({ S25957[290] }),
  .Z({ w[290] })
);
BUF_X1 #() 
BUF_X1_623_ (
  .A({ S25957[291] }),
  .Z({ w[291] })
);
BUF_X1 #() 
BUF_X1_624_ (
  .A({ S25957[292] }),
  .Z({ w[292] })
);
BUF_X1 #() 
BUF_X1_625_ (
  .A({ S25957[293] }),
  .Z({ w[293] })
);
BUF_X1 #() 
BUF_X1_626_ (
  .A({ S25957[294] }),
  .Z({ w[294] })
);
BUF_X1 #() 
BUF_X1_627_ (
  .A({ S25957[295] }),
  .Z({ w[295] })
);
BUF_X1 #() 
BUF_X1_628_ (
  .A({ S25957[296] }),
  .Z({ w[296] })
);
BUF_X1 #() 
BUF_X1_629_ (
  .A({ S25957[297] }),
  .Z({ w[297] })
);
BUF_X1 #() 
BUF_X1_630_ (
  .A({ S25957[298] }),
  .Z({ w[298] })
);
BUF_X1 #() 
BUF_X1_631_ (
  .A({ S25957[299] }),
  .Z({ w[299] })
);
BUF_X1 #() 
BUF_X1_632_ (
  .A({ S25957[3] }),
  .Z({ w[3] })
);
BUF_X1 #() 
BUF_X1_633_ (
  .A({ S25957[30] }),
  .Z({ w[30] })
);
BUF_X1 #() 
BUF_X1_634_ (
  .A({ S25957[300] }),
  .Z({ w[300] })
);
BUF_X1 #() 
BUF_X1_635_ (
  .A({ S25957[301] }),
  .Z({ w[301] })
);
BUF_X1 #() 
BUF_X1_636_ (
  .A({ S25957[302] }),
  .Z({ w[302] })
);
BUF_X1 #() 
BUF_X1_637_ (
  .A({ S25957[303] }),
  .Z({ w[303] })
);
BUF_X1 #() 
BUF_X1_638_ (
  .A({ S25957[304] }),
  .Z({ w[304] })
);
BUF_X1 #() 
BUF_X1_639_ (
  .A({ S25957[305] }),
  .Z({ w[305] })
);
BUF_X1 #() 
BUF_X1_640_ (
  .A({ S25957[306] }),
  .Z({ w[306] })
);
BUF_X1 #() 
BUF_X1_641_ (
  .A({ S25957[307] }),
  .Z({ w[307] })
);
BUF_X1 #() 
BUF_X1_642_ (
  .A({ S25957[308] }),
  .Z({ w[308] })
);
BUF_X1 #() 
BUF_X1_643_ (
  .A({ S25957[309] }),
  .Z({ w[309] })
);
BUF_X1 #() 
BUF_X1_644_ (
  .A({ S25957[31] }),
  .Z({ w[31] })
);
BUF_X1 #() 
BUF_X1_645_ (
  .A({ S25957[310] }),
  .Z({ w[310] })
);
BUF_X1 #() 
BUF_X1_646_ (
  .A({ S25957[311] }),
  .Z({ w[311] })
);
BUF_X1 #() 
BUF_X1_647_ (
  .A({ S25957[312] }),
  .Z({ w[312] })
);
BUF_X1 #() 
BUF_X1_648_ (
  .A({ S25957[313] }),
  .Z({ w[313] })
);
BUF_X1 #() 
BUF_X1_649_ (
  .A({ S25957[314] }),
  .Z({ w[314] })
);
BUF_X1 #() 
BUF_X1_650_ (
  .A({ S25957[315] }),
  .Z({ w[315] })
);
BUF_X1 #() 
BUF_X1_651_ (
  .A({ S25957[316] }),
  .Z({ w[316] })
);
BUF_X1 #() 
BUF_X1_652_ (
  .A({ S25957[317] }),
  .Z({ w[317] })
);
BUF_X1 #() 
BUF_X1_653_ (
  .A({ S25957[318] }),
  .Z({ w[318] })
);
BUF_X1 #() 
BUF_X1_654_ (
  .A({ S25957[319] }),
  .Z({ w[319] })
);
BUF_X1 #() 
BUF_X1_655_ (
  .A({ S25957[32] }),
  .Z({ w[32] })
);
BUF_X1 #() 
BUF_X1_656_ (
  .A({ S25957[320] }),
  .Z({ w[320] })
);
BUF_X1 #() 
BUF_X1_657_ (
  .A({ S25957[321] }),
  .Z({ w[321] })
);
BUF_X1 #() 
BUF_X1_658_ (
  .A({ S25957[322] }),
  .Z({ w[322] })
);
BUF_X1 #() 
BUF_X1_659_ (
  .A({ S25957[323] }),
  .Z({ w[323] })
);
BUF_X1 #() 
BUF_X1_660_ (
  .A({ S25957[324] }),
  .Z({ w[324] })
);
BUF_X1 #() 
BUF_X1_661_ (
  .A({ S25957[325] }),
  .Z({ w[325] })
);
BUF_X1 #() 
BUF_X1_662_ (
  .A({ S25957[326] }),
  .Z({ w[326] })
);
BUF_X1 #() 
BUF_X1_663_ (
  .A({ S25957[327] }),
  .Z({ w[327] })
);
BUF_X1 #() 
BUF_X1_664_ (
  .A({ S25957[328] }),
  .Z({ w[328] })
);
BUF_X1 #() 
BUF_X1_665_ (
  .A({ S25957[329] }),
  .Z({ w[329] })
);
BUF_X1 #() 
BUF_X1_666_ (
  .A({ S25957[33] }),
  .Z({ w[33] })
);
BUF_X1 #() 
BUF_X1_667_ (
  .A({ S25957[330] }),
  .Z({ w[330] })
);
BUF_X1 #() 
BUF_X1_668_ (
  .A({ S25957[331] }),
  .Z({ w[331] })
);
BUF_X1 #() 
BUF_X1_669_ (
  .A({ S25957[332] }),
  .Z({ w[332] })
);
BUF_X1 #() 
BUF_X1_670_ (
  .A({ S25957[333] }),
  .Z({ w[333] })
);
BUF_X1 #() 
BUF_X1_671_ (
  .A({ S25957[334] }),
  .Z({ w[334] })
);
BUF_X1 #() 
BUF_X1_672_ (
  .A({ S25957[335] }),
  .Z({ w[335] })
);
BUF_X1 #() 
BUF_X1_673_ (
  .A({ S25957[336] }),
  .Z({ w[336] })
);
BUF_X1 #() 
BUF_X1_674_ (
  .A({ S25957[337] }),
  .Z({ w[337] })
);
BUF_X1 #() 
BUF_X1_675_ (
  .A({ S25957[338] }),
  .Z({ w[338] })
);
BUF_X1 #() 
BUF_X1_676_ (
  .A({ S25957[339] }),
  .Z({ w[339] })
);
BUF_X1 #() 
BUF_X1_677_ (
  .A({ S25957[34] }),
  .Z({ w[34] })
);
BUF_X1 #() 
BUF_X1_678_ (
  .A({ S25957[340] }),
  .Z({ w[340] })
);
BUF_X1 #() 
BUF_X1_679_ (
  .A({ S25957[341] }),
  .Z({ w[341] })
);
BUF_X1 #() 
BUF_X1_680_ (
  .A({ S25957[342] }),
  .Z({ w[342] })
);
BUF_X1 #() 
BUF_X1_681_ (
  .A({ S25957[343] }),
  .Z({ w[343] })
);
BUF_X1 #() 
BUF_X1_682_ (
  .A({ S25957[344] }),
  .Z({ w[344] })
);
BUF_X1 #() 
BUF_X1_683_ (
  .A({ S25957[345] }),
  .Z({ w[345] })
);
BUF_X1 #() 
BUF_X1_684_ (
  .A({ S25957[346] }),
  .Z({ w[346] })
);
BUF_X1 #() 
BUF_X1_685_ (
  .A({ S25957[347] }),
  .Z({ w[347] })
);
BUF_X1 #() 
BUF_X1_686_ (
  .A({ S25957[348] }),
  .Z({ w[348] })
);
BUF_X1 #() 
BUF_X1_687_ (
  .A({ S25957[349] }),
  .Z({ w[349] })
);
BUF_X1 #() 
BUF_X1_688_ (
  .A({ S25957[35] }),
  .Z({ w[35] })
);
BUF_X1 #() 
BUF_X1_689_ (
  .A({ S25957[350] }),
  .Z({ w[350] })
);
BUF_X1 #() 
BUF_X1_690_ (
  .A({ S25957[351] }),
  .Z({ w[351] })
);
BUF_X1 #() 
BUF_X1_691_ (
  .A({ S25957[352] }),
  .Z({ w[352] })
);
BUF_X1 #() 
BUF_X1_692_ (
  .A({ S25957[353] }),
  .Z({ w[353] })
);
BUF_X1 #() 
BUF_X1_693_ (
  .A({ S25957[354] }),
  .Z({ w[354] })
);
BUF_X1 #() 
BUF_X1_694_ (
  .A({ S25957[355] }),
  .Z({ w[355] })
);
BUF_X1 #() 
BUF_X1_695_ (
  .A({ S25957[356] }),
  .Z({ w[356] })
);
BUF_X1 #() 
BUF_X1_696_ (
  .A({ S25957[357] }),
  .Z({ w[357] })
);
BUF_X1 #() 
BUF_X1_697_ (
  .A({ S25957[358] }),
  .Z({ w[358] })
);
BUF_X1 #() 
BUF_X1_698_ (
  .A({ S25957[359] }),
  .Z({ w[359] })
);
BUF_X1 #() 
BUF_X1_699_ (
  .A({ S25957[36] }),
  .Z({ w[36] })
);
BUF_X1 #() 
BUF_X1_700_ (
  .A({ S25957[360] }),
  .Z({ w[360] })
);
BUF_X1 #() 
BUF_X1_701_ (
  .A({ S25957[361] }),
  .Z({ w[361] })
);
BUF_X1 #() 
BUF_X1_702_ (
  .A({ S25957[362] }),
  .Z({ w[362] })
);
BUF_X1 #() 
BUF_X1_703_ (
  .A({ S25957[363] }),
  .Z({ w[363] })
);
BUF_X1 #() 
BUF_X1_704_ (
  .A({ S25957[364] }),
  .Z({ w[364] })
);
BUF_X1 #() 
BUF_X1_705_ (
  .A({ S25957[365] }),
  .Z({ w[365] })
);
BUF_X1 #() 
BUF_X1_706_ (
  .A({ S25957[366] }),
  .Z({ w[366] })
);
BUF_X1 #() 
BUF_X1_707_ (
  .A({ S25957[367] }),
  .Z({ w[367] })
);
BUF_X1 #() 
BUF_X1_708_ (
  .A({ S25957[368] }),
  .Z({ w[368] })
);
BUF_X1 #() 
BUF_X1_709_ (
  .A({ S25957[369] }),
  .Z({ w[369] })
);
BUF_X1 #() 
BUF_X1_710_ (
  .A({ S25957[37] }),
  .Z({ w[37] })
);
BUF_X1 #() 
BUF_X1_711_ (
  .A({ S25957[370] }),
  .Z({ w[370] })
);
BUF_X1 #() 
BUF_X1_712_ (
  .A({ S25957[371] }),
  .Z({ w[371] })
);
BUF_X1 #() 
BUF_X1_713_ (
  .A({ S25957[372] }),
  .Z({ w[372] })
);
BUF_X1 #() 
BUF_X1_714_ (
  .A({ S25957[373] }),
  .Z({ w[373] })
);
BUF_X1 #() 
BUF_X1_715_ (
  .A({ S25957[374] }),
  .Z({ w[374] })
);
BUF_X1 #() 
BUF_X1_716_ (
  .A({ S25957[375] }),
  .Z({ w[375] })
);
BUF_X1 #() 
BUF_X1_717_ (
  .A({ S25957[376] }),
  .Z({ w[376] })
);
BUF_X1 #() 
BUF_X1_718_ (
  .A({ S25957[377] }),
  .Z({ w[377] })
);
BUF_X1 #() 
BUF_X1_719_ (
  .A({ S25957[378] }),
  .Z({ w[378] })
);
BUF_X1 #() 
BUF_X1_720_ (
  .A({ S25957[379] }),
  .Z({ w[379] })
);
BUF_X1 #() 
BUF_X1_721_ (
  .A({ S25957[38] }),
  .Z({ w[38] })
);
BUF_X1 #() 
BUF_X1_722_ (
  .A({ S25957[380] }),
  .Z({ w[380] })
);
BUF_X1 #() 
BUF_X1_723_ (
  .A({ S25957[381] }),
  .Z({ w[381] })
);
BUF_X1 #() 
BUF_X1_724_ (
  .A({ S25957[382] }),
  .Z({ w[382] })
);
BUF_X1 #() 
BUF_X1_725_ (
  .A({ S25957[383] }),
  .Z({ w[383] })
);
BUF_X1 #() 
BUF_X1_726_ (
  .A({ S25957[384] }),
  .Z({ w[384] })
);
BUF_X1 #() 
BUF_X1_727_ (
  .A({ S25957[385] }),
  .Z({ w[385] })
);
BUF_X1 #() 
BUF_X1_728_ (
  .A({ S25957[386] }),
  .Z({ w[386] })
);
BUF_X1 #() 
BUF_X1_729_ (
  .A({ S25957[387] }),
  .Z({ w[387] })
);
BUF_X1 #() 
BUF_X1_730_ (
  .A({ S25957[388] }),
  .Z({ w[388] })
);
BUF_X1 #() 
BUF_X1_731_ (
  .A({ S25957[389] }),
  .Z({ w[389] })
);
BUF_X1 #() 
BUF_X1_732_ (
  .A({ S25957[39] }),
  .Z({ w[39] })
);
BUF_X1 #() 
BUF_X1_733_ (
  .A({ S25957[390] }),
  .Z({ w[390] })
);
BUF_X1 #() 
BUF_X1_734_ (
  .A({ S25957[391] }),
  .Z({ w[391] })
);
BUF_X1 #() 
BUF_X1_735_ (
  .A({ S25957[392] }),
  .Z({ w[392] })
);
BUF_X1 #() 
BUF_X1_736_ (
  .A({ S25957[393] }),
  .Z({ w[393] })
);
BUF_X1 #() 
BUF_X1_737_ (
  .A({ S25957[394] }),
  .Z({ w[394] })
);
BUF_X1 #() 
BUF_X1_738_ (
  .A({ S25957[395] }),
  .Z({ w[395] })
);
BUF_X1 #() 
BUF_X1_739_ (
  .A({ S25957[396] }),
  .Z({ w[396] })
);
BUF_X1 #() 
BUF_X1_740_ (
  .A({ S25957[397] }),
  .Z({ w[397] })
);
BUF_X1 #() 
BUF_X1_741_ (
  .A({ S25957[398] }),
  .Z({ w[398] })
);
BUF_X1 #() 
BUF_X1_742_ (
  .A({ S25957[399] }),
  .Z({ w[399] })
);
BUF_X1 #() 
BUF_X1_743_ (
  .A({ S25957[4] }),
  .Z({ w[4] })
);
BUF_X1 #() 
BUF_X1_744_ (
  .A({ S25957[40] }),
  .Z({ w[40] })
);
BUF_X1 #() 
BUF_X1_745_ (
  .A({ S25957[400] }),
  .Z({ w[400] })
);
BUF_X1 #() 
BUF_X1_746_ (
  .A({ S25957[401] }),
  .Z({ w[401] })
);
BUF_X1 #() 
BUF_X1_747_ (
  .A({ S25957[402] }),
  .Z({ w[402] })
);
BUF_X1 #() 
BUF_X1_748_ (
  .A({ S25957[403] }),
  .Z({ w[403] })
);
BUF_X1 #() 
BUF_X1_749_ (
  .A({ S25957[404] }),
  .Z({ w[404] })
);
BUF_X1 #() 
BUF_X1_750_ (
  .A({ S25957[405] }),
  .Z({ w[405] })
);
BUF_X1 #() 
BUF_X1_751_ (
  .A({ S25957[406] }),
  .Z({ w[406] })
);
BUF_X1 #() 
BUF_X1_752_ (
  .A({ S25957[407] }),
  .Z({ w[407] })
);
BUF_X1 #() 
BUF_X1_753_ (
  .A({ S25957[408] }),
  .Z({ w[408] })
);
BUF_X1 #() 
BUF_X1_754_ (
  .A({ S25957[409] }),
  .Z({ w[409] })
);
BUF_X1 #() 
BUF_X1_755_ (
  .A({ S25957[41] }),
  .Z({ w[41] })
);
BUF_X1 #() 
BUF_X1_756_ (
  .A({ S25957[410] }),
  .Z({ w[410] })
);
BUF_X1 #() 
BUF_X1_757_ (
  .A({ S25957[411] }),
  .Z({ w[411] })
);
BUF_X1 #() 
BUF_X1_758_ (
  .A({ S25957[412] }),
  .Z({ w[412] })
);
BUF_X1 #() 
BUF_X1_759_ (
  .A({ S25957[413] }),
  .Z({ w[413] })
);
BUF_X1 #() 
BUF_X1_760_ (
  .A({ S25957[414] }),
  .Z({ w[414] })
);
BUF_X1 #() 
BUF_X1_761_ (
  .A({ S25957[415] }),
  .Z({ w[415] })
);
BUF_X1 #() 
BUF_X1_762_ (
  .A({ S25957[416] }),
  .Z({ w[416] })
);
BUF_X1 #() 
BUF_X1_763_ (
  .A({ S25957[417] }),
  .Z({ w[417] })
);
BUF_X1 #() 
BUF_X1_764_ (
  .A({ S25957[418] }),
  .Z({ w[418] })
);
BUF_X1 #() 
BUF_X1_765_ (
  .A({ S25957[419] }),
  .Z({ w[419] })
);
BUF_X1 #() 
BUF_X1_766_ (
  .A({ S25957[42] }),
  .Z({ w[42] })
);
BUF_X1 #() 
BUF_X1_767_ (
  .A({ S25957[420] }),
  .Z({ w[420] })
);
BUF_X1 #() 
BUF_X1_768_ (
  .A({ S25957[421] }),
  .Z({ w[421] })
);
BUF_X1 #() 
BUF_X1_769_ (
  .A({ S25957[422] }),
  .Z({ w[422] })
);
BUF_X1 #() 
BUF_X1_770_ (
  .A({ S25957[423] }),
  .Z({ w[423] })
);
BUF_X1 #() 
BUF_X1_771_ (
  .A({ S25957[424] }),
  .Z({ w[424] })
);
BUF_X1 #() 
BUF_X1_772_ (
  .A({ S25957[425] }),
  .Z({ w[425] })
);
BUF_X1 #() 
BUF_X1_773_ (
  .A({ S25957[426] }),
  .Z({ w[426] })
);
BUF_X1 #() 
BUF_X1_774_ (
  .A({ S25957[427] }),
  .Z({ w[427] })
);
BUF_X1 #() 
BUF_X1_775_ (
  .A({ S25957[428] }),
  .Z({ w[428] })
);
BUF_X1 #() 
BUF_X1_776_ (
  .A({ S25957[429] }),
  .Z({ w[429] })
);
BUF_X1 #() 
BUF_X1_777_ (
  .A({ S25957[43] }),
  .Z({ w[43] })
);
BUF_X1 #() 
BUF_X1_778_ (
  .A({ S25957[430] }),
  .Z({ w[430] })
);
BUF_X1 #() 
BUF_X1_779_ (
  .A({ S25957[431] }),
  .Z({ w[431] })
);
BUF_X1 #() 
BUF_X1_780_ (
  .A({ S25957[432] }),
  .Z({ w[432] })
);
BUF_X1 #() 
BUF_X1_781_ (
  .A({ S25957[433] }),
  .Z({ w[433] })
);
BUF_X1 #() 
BUF_X1_782_ (
  .A({ S25957[434] }),
  .Z({ w[434] })
);
BUF_X1 #() 
BUF_X1_783_ (
  .A({ S25957[435] }),
  .Z({ w[435] })
);
BUF_X1 #() 
BUF_X1_784_ (
  .A({ S25957[436] }),
  .Z({ w[436] })
);
BUF_X1 #() 
BUF_X1_785_ (
  .A({ S25957[437] }),
  .Z({ w[437] })
);
BUF_X1 #() 
BUF_X1_786_ (
  .A({ S25957[438] }),
  .Z({ w[438] })
);
BUF_X1 #() 
BUF_X1_787_ (
  .A({ S25957[439] }),
  .Z({ w[439] })
);
BUF_X1 #() 
BUF_X1_788_ (
  .A({ S25957[44] }),
  .Z({ w[44] })
);
BUF_X1 #() 
BUF_X1_789_ (
  .A({ S25957[440] }),
  .Z({ w[440] })
);
BUF_X1 #() 
BUF_X1_790_ (
  .A({ S25957[441] }),
  .Z({ w[441] })
);
BUF_X1 #() 
BUF_X1_791_ (
  .A({ S25957[442] }),
  .Z({ w[442] })
);
BUF_X1 #() 
BUF_X1_792_ (
  .A({ S25957[443] }),
  .Z({ w[443] })
);
BUF_X1 #() 
BUF_X1_793_ (
  .A({ S25957[444] }),
  .Z({ w[444] })
);
BUF_X1 #() 
BUF_X1_794_ (
  .A({ S25957[445] }),
  .Z({ w[445] })
);
BUF_X1 #() 
BUF_X1_795_ (
  .A({ S25957[446] }),
  .Z({ w[446] })
);
BUF_X1 #() 
BUF_X1_796_ (
  .A({ S25957[447] }),
  .Z({ w[447] })
);
BUF_X1 #() 
BUF_X1_797_ (
  .A({ S25957[448] }),
  .Z({ w[448] })
);
BUF_X1 #() 
BUF_X1_798_ (
  .A({ S25957[449] }),
  .Z({ w[449] })
);
BUF_X1 #() 
BUF_X1_799_ (
  .A({ S25957[45] }),
  .Z({ w[45] })
);
BUF_X1 #() 
BUF_X1_800_ (
  .A({ S25957[450] }),
  .Z({ w[450] })
);
BUF_X1 #() 
BUF_X1_801_ (
  .A({ S25957[451] }),
  .Z({ w[451] })
);
BUF_X1 #() 
BUF_X1_802_ (
  .A({ S25957[452] }),
  .Z({ w[452] })
);
BUF_X1 #() 
BUF_X1_803_ (
  .A({ S25957[453] }),
  .Z({ w[453] })
);
BUF_X1 #() 
BUF_X1_804_ (
  .A({ S25957[454] }),
  .Z({ w[454] })
);
BUF_X1 #() 
BUF_X1_805_ (
  .A({ S25957[455] }),
  .Z({ w[455] })
);
BUF_X1 #() 
BUF_X1_806_ (
  .A({ S25957[456] }),
  .Z({ w[456] })
);
BUF_X1 #() 
BUF_X1_807_ (
  .A({ S25957[457] }),
  .Z({ w[457] })
);
BUF_X1 #() 
BUF_X1_808_ (
  .A({ S25957[458] }),
  .Z({ w[458] })
);
BUF_X1 #() 
BUF_X1_809_ (
  .A({ S25957[459] }),
  .Z({ w[459] })
);
BUF_X1 #() 
BUF_X1_810_ (
  .A({ S25957[46] }),
  .Z({ w[46] })
);
BUF_X1 #() 
BUF_X1_811_ (
  .A({ S25957[460] }),
  .Z({ w[460] })
);
BUF_X1 #() 
BUF_X1_812_ (
  .A({ S25957[461] }),
  .Z({ w[461] })
);
BUF_X1 #() 
BUF_X1_813_ (
  .A({ S25957[462] }),
  .Z({ w[462] })
);
BUF_X1 #() 
BUF_X1_814_ (
  .A({ S25957[463] }),
  .Z({ w[463] })
);
BUF_X1 #() 
BUF_X1_815_ (
  .A({ S25957[464] }),
  .Z({ w[464] })
);
BUF_X1 #() 
BUF_X1_816_ (
  .A({ S25957[465] }),
  .Z({ w[465] })
);
BUF_X1 #() 
BUF_X1_817_ (
  .A({ S25957[466] }),
  .Z({ w[466] })
);
BUF_X1 #() 
BUF_X1_818_ (
  .A({ S25957[467] }),
  .Z({ w[467] })
);
BUF_X1 #() 
BUF_X1_819_ (
  .A({ S25957[468] }),
  .Z({ w[468] })
);
BUF_X1 #() 
BUF_X1_820_ (
  .A({ S25957[469] }),
  .Z({ w[469] })
);
BUF_X1 #() 
BUF_X1_821_ (
  .A({ S25957[47] }),
  .Z({ w[47] })
);
BUF_X1 #() 
BUF_X1_822_ (
  .A({ S25957[470] }),
  .Z({ w[470] })
);
BUF_X1 #() 
BUF_X1_823_ (
  .A({ S25957[471] }),
  .Z({ w[471] })
);
BUF_X1 #() 
BUF_X1_824_ (
  .A({ S25957[472] }),
  .Z({ w[472] })
);
BUF_X1 #() 
BUF_X1_825_ (
  .A({ S25957[473] }),
  .Z({ w[473] })
);
BUF_X1 #() 
BUF_X1_826_ (
  .A({ S25957[474] }),
  .Z({ w[474] })
);
BUF_X1 #() 
BUF_X1_827_ (
  .A({ S25957[475] }),
  .Z({ w[475] })
);
BUF_X1 #() 
BUF_X1_828_ (
  .A({ S25957[476] }),
  .Z({ w[476] })
);
BUF_X1 #() 
BUF_X1_829_ (
  .A({ S25957[477] }),
  .Z({ w[477] })
);
BUF_X1 #() 
BUF_X1_830_ (
  .A({ S25957[478] }),
  .Z({ w[478] })
);
BUF_X1 #() 
BUF_X1_831_ (
  .A({ S25957[479] }),
  .Z({ w[479] })
);
BUF_X1 #() 
BUF_X1_832_ (
  .A({ S25957[48] }),
  .Z({ w[48] })
);
BUF_X1 #() 
BUF_X1_833_ (
  .A({ S25957[480] }),
  .Z({ w[480] })
);
BUF_X1 #() 
BUF_X1_834_ (
  .A({ S25957[481] }),
  .Z({ w[481] })
);
BUF_X1 #() 
BUF_X1_835_ (
  .A({ S25957[482] }),
  .Z({ w[482] })
);
BUF_X1 #() 
BUF_X1_836_ (
  .A({ S25957[483] }),
  .Z({ w[483] })
);
BUF_X1 #() 
BUF_X1_837_ (
  .A({ S25957[484] }),
  .Z({ w[484] })
);
BUF_X1 #() 
BUF_X1_838_ (
  .A({ S25957[485] }),
  .Z({ w[485] })
);
BUF_X1 #() 
BUF_X1_839_ (
  .A({ S25957[486] }),
  .Z({ w[486] })
);
BUF_X1 #() 
BUF_X1_840_ (
  .A({ S25957[487] }),
  .Z({ w[487] })
);
BUF_X1 #() 
BUF_X1_841_ (
  .A({ S25957[488] }),
  .Z({ w[488] })
);
BUF_X1 #() 
BUF_X1_842_ (
  .A({ S25957[489] }),
  .Z({ w[489] })
);
BUF_X1 #() 
BUF_X1_843_ (
  .A({ S25957[49] }),
  .Z({ w[49] })
);
BUF_X1 #() 
BUF_X1_844_ (
  .A({ S25957[490] }),
  .Z({ w[490] })
);
BUF_X1 #() 
BUF_X1_845_ (
  .A({ S25957[491] }),
  .Z({ w[491] })
);
BUF_X1 #() 
BUF_X1_846_ (
  .A({ S25957[492] }),
  .Z({ w[492] })
);
BUF_X1 #() 
BUF_X1_847_ (
  .A({ S25957[493] }),
  .Z({ w[493] })
);
BUF_X1 #() 
BUF_X1_848_ (
  .A({ S25957[494] }),
  .Z({ w[494] })
);
BUF_X1 #() 
BUF_X1_849_ (
  .A({ S25957[495] }),
  .Z({ w[495] })
);
BUF_X1 #() 
BUF_X1_850_ (
  .A({ S25957[496] }),
  .Z({ w[496] })
);
BUF_X1 #() 
BUF_X1_851_ (
  .A({ S25957[497] }),
  .Z({ w[497] })
);
BUF_X1 #() 
BUF_X1_852_ (
  .A({ S25957[498] }),
  .Z({ w[498] })
);
BUF_X1 #() 
BUF_X1_853_ (
  .A({ S25957[499] }),
  .Z({ w[499] })
);
BUF_X1 #() 
BUF_X1_854_ (
  .A({ S25957[5] }),
  .Z({ w[5] })
);
BUF_X1 #() 
BUF_X1_855_ (
  .A({ S25957[50] }),
  .Z({ w[50] })
);
BUF_X1 #() 
BUF_X1_856_ (
  .A({ S25957[500] }),
  .Z({ w[500] })
);
BUF_X1 #() 
BUF_X1_857_ (
  .A({ S25957[501] }),
  .Z({ w[501] })
);
BUF_X1 #() 
BUF_X1_858_ (
  .A({ S25957[502] }),
  .Z({ w[502] })
);
BUF_X1 #() 
BUF_X1_859_ (
  .A({ S25957[503] }),
  .Z({ w[503] })
);
BUF_X1 #() 
BUF_X1_860_ (
  .A({ S25957[504] }),
  .Z({ w[504] })
);
BUF_X1 #() 
BUF_X1_861_ (
  .A({ S25957[505] }),
  .Z({ w[505] })
);
BUF_X1 #() 
BUF_X1_862_ (
  .A({ S25957[506] }),
  .Z({ w[506] })
);
BUF_X1 #() 
BUF_X1_863_ (
  .A({ S25957[507] }),
  .Z({ w[507] })
);
BUF_X1 #() 
BUF_X1_864_ (
  .A({ S25957[508] }),
  .Z({ w[508] })
);
BUF_X1 #() 
BUF_X1_865_ (
  .A({ S25957[509] }),
  .Z({ w[509] })
);
BUF_X1 #() 
BUF_X1_866_ (
  .A({ S25957[51] }),
  .Z({ w[51] })
);
BUF_X1 #() 
BUF_X1_867_ (
  .A({ S25957[510] }),
  .Z({ w[510] })
);
BUF_X1 #() 
BUF_X1_868_ (
  .A({ S25957[511] }),
  .Z({ w[511] })
);
BUF_X1 #() 
BUF_X1_869_ (
  .A({ S25957[512] }),
  .Z({ w[512] })
);
BUF_X1 #() 
BUF_X1_870_ (
  .A({ S25957[513] }),
  .Z({ w[513] })
);
BUF_X1 #() 
BUF_X1_871_ (
  .A({ S25957[514] }),
  .Z({ w[514] })
);
BUF_X1 #() 
BUF_X1_872_ (
  .A({ S25957[515] }),
  .Z({ w[515] })
);
BUF_X1 #() 
BUF_X1_873_ (
  .A({ S25957[516] }),
  .Z({ w[516] })
);
BUF_X1 #() 
BUF_X1_874_ (
  .A({ S25957[517] }),
  .Z({ w[517] })
);
BUF_X1 #() 
BUF_X1_875_ (
  .A({ S25957[518] }),
  .Z({ w[518] })
);
BUF_X1 #() 
BUF_X1_876_ (
  .A({ S25957[519] }),
  .Z({ w[519] })
);
BUF_X1 #() 
BUF_X1_877_ (
  .A({ S25957[52] }),
  .Z({ w[52] })
);
BUF_X1 #() 
BUF_X1_878_ (
  .A({ S25957[520] }),
  .Z({ w[520] })
);
BUF_X1 #() 
BUF_X1_879_ (
  .A({ S25957[521] }),
  .Z({ w[521] })
);
BUF_X1 #() 
BUF_X1_880_ (
  .A({ S25957[522] }),
  .Z({ w[522] })
);
BUF_X1 #() 
BUF_X1_881_ (
  .A({ S25957[523] }),
  .Z({ w[523] })
);
BUF_X1 #() 
BUF_X1_882_ (
  .A({ S25957[524] }),
  .Z({ w[524] })
);
BUF_X1 #() 
BUF_X1_883_ (
  .A({ S25957[525] }),
  .Z({ w[525] })
);
BUF_X1 #() 
BUF_X1_884_ (
  .A({ S25957[526] }),
  .Z({ w[526] })
);
BUF_X1 #() 
BUF_X1_885_ (
  .A({ S25957[527] }),
  .Z({ w[527] })
);
BUF_X1 #() 
BUF_X1_886_ (
  .A({ S25957[528] }),
  .Z({ w[528] })
);
BUF_X1 #() 
BUF_X1_887_ (
  .A({ S25957[529] }),
  .Z({ w[529] })
);
BUF_X1 #() 
BUF_X1_888_ (
  .A({ S25957[53] }),
  .Z({ w[53] })
);
BUF_X1 #() 
BUF_X1_889_ (
  .A({ S25957[530] }),
  .Z({ w[530] })
);
BUF_X1 #() 
BUF_X1_890_ (
  .A({ S25957[531] }),
  .Z({ w[531] })
);
BUF_X1 #() 
BUF_X1_891_ (
  .A({ S25957[532] }),
  .Z({ w[532] })
);
BUF_X1 #() 
BUF_X1_892_ (
  .A({ S25957[533] }),
  .Z({ w[533] })
);
BUF_X1 #() 
BUF_X1_893_ (
  .A({ S25957[534] }),
  .Z({ w[534] })
);
BUF_X1 #() 
BUF_X1_894_ (
  .A({ S25957[535] }),
  .Z({ w[535] })
);
BUF_X1 #() 
BUF_X1_895_ (
  .A({ S25957[536] }),
  .Z({ w[536] })
);
BUF_X1 #() 
BUF_X1_896_ (
  .A({ S25957[537] }),
  .Z({ w[537] })
);
BUF_X1 #() 
BUF_X1_897_ (
  .A({ S25957[538] }),
  .Z({ w[538] })
);
BUF_X1 #() 
BUF_X1_898_ (
  .A({ S25957[539] }),
  .Z({ w[539] })
);
BUF_X1 #() 
BUF_X1_899_ (
  .A({ S25957[54] }),
  .Z({ w[54] })
);
BUF_X1 #() 
BUF_X1_900_ (
  .A({ S25957[540] }),
  .Z({ w[540] })
);
BUF_X1 #() 
BUF_X1_901_ (
  .A({ S25957[541] }),
  .Z({ w[541] })
);
BUF_X1 #() 
BUF_X1_902_ (
  .A({ S25957[542] }),
  .Z({ w[542] })
);
BUF_X1 #() 
BUF_X1_903_ (
  .A({ S25957[543] }),
  .Z({ w[543] })
);
BUF_X1 #() 
BUF_X1_904_ (
  .A({ S25957[544] }),
  .Z({ w[544] })
);
BUF_X1 #() 
BUF_X1_905_ (
  .A({ S25957[545] }),
  .Z({ w[545] })
);
BUF_X1 #() 
BUF_X1_906_ (
  .A({ S25957[546] }),
  .Z({ w[546] })
);
BUF_X1 #() 
BUF_X1_907_ (
  .A({ S25957[547] }),
  .Z({ w[547] })
);
BUF_X1 #() 
BUF_X1_908_ (
  .A({ S25957[548] }),
  .Z({ w[548] })
);
BUF_X1 #() 
BUF_X1_909_ (
  .A({ S25957[549] }),
  .Z({ w[549] })
);
BUF_X1 #() 
BUF_X1_910_ (
  .A({ S25957[55] }),
  .Z({ w[55] })
);
BUF_X1 #() 
BUF_X1_911_ (
  .A({ S25957[550] }),
  .Z({ w[550] })
);
BUF_X1 #() 
BUF_X1_912_ (
  .A({ S25957[551] }),
  .Z({ w[551] })
);
BUF_X1 #() 
BUF_X1_913_ (
  .A({ S25957[552] }),
  .Z({ w[552] })
);
BUF_X1 #() 
BUF_X1_914_ (
  .A({ S25957[553] }),
  .Z({ w[553] })
);
BUF_X1 #() 
BUF_X1_915_ (
  .A({ S25957[554] }),
  .Z({ w[554] })
);
BUF_X1 #() 
BUF_X1_916_ (
  .A({ S25957[555] }),
  .Z({ w[555] })
);
BUF_X1 #() 
BUF_X1_917_ (
  .A({ S25957[556] }),
  .Z({ w[556] })
);
BUF_X1 #() 
BUF_X1_918_ (
  .A({ S25957[557] }),
  .Z({ w[557] })
);
BUF_X1 #() 
BUF_X1_919_ (
  .A({ S25957[558] }),
  .Z({ w[558] })
);
BUF_X1 #() 
BUF_X1_920_ (
  .A({ S25957[559] }),
  .Z({ w[559] })
);
BUF_X1 #() 
BUF_X1_921_ (
  .A({ S25957[56] }),
  .Z({ w[56] })
);
BUF_X1 #() 
BUF_X1_922_ (
  .A({ S25957[560] }),
  .Z({ w[560] })
);
BUF_X1 #() 
BUF_X1_923_ (
  .A({ S25957[561] }),
  .Z({ w[561] })
);
BUF_X1 #() 
BUF_X1_924_ (
  .A({ S25957[562] }),
  .Z({ w[562] })
);
BUF_X1 #() 
BUF_X1_925_ (
  .A({ S25957[563] }),
  .Z({ w[563] })
);
BUF_X1 #() 
BUF_X1_926_ (
  .A({ S25957[564] }),
  .Z({ w[564] })
);
BUF_X1 #() 
BUF_X1_927_ (
  .A({ S25957[565] }),
  .Z({ w[565] })
);
BUF_X1 #() 
BUF_X1_928_ (
  .A({ S25957[566] }),
  .Z({ w[566] })
);
BUF_X1 #() 
BUF_X1_929_ (
  .A({ S25957[567] }),
  .Z({ w[567] })
);
BUF_X1 #() 
BUF_X1_930_ (
  .A({ S25957[568] }),
  .Z({ w[568] })
);
BUF_X1 #() 
BUF_X1_931_ (
  .A({ S25957[569] }),
  .Z({ w[569] })
);
BUF_X1 #() 
BUF_X1_932_ (
  .A({ S25957[57] }),
  .Z({ w[57] })
);
BUF_X1 #() 
BUF_X1_933_ (
  .A({ S25957[570] }),
  .Z({ w[570] })
);
BUF_X1 #() 
BUF_X1_934_ (
  .A({ S25957[571] }),
  .Z({ w[571] })
);
BUF_X1 #() 
BUF_X1_935_ (
  .A({ S25957[572] }),
  .Z({ w[572] })
);
BUF_X1 #() 
BUF_X1_936_ (
  .A({ S25957[573] }),
  .Z({ w[573] })
);
BUF_X1 #() 
BUF_X1_937_ (
  .A({ S25957[574] }),
  .Z({ w[574] })
);
BUF_X1 #() 
BUF_X1_938_ (
  .A({ S25957[575] }),
  .Z({ w[575] })
);
BUF_X1 #() 
BUF_X1_939_ (
  .A({ S25957[576] }),
  .Z({ w[576] })
);
BUF_X1 #() 
BUF_X1_940_ (
  .A({ S25957[577] }),
  .Z({ w[577] })
);
BUF_X1 #() 
BUF_X1_941_ (
  .A({ S25957[578] }),
  .Z({ w[578] })
);
BUF_X1 #() 
BUF_X1_942_ (
  .A({ S25957[579] }),
  .Z({ w[579] })
);
BUF_X1 #() 
BUF_X1_943_ (
  .A({ S25957[58] }),
  .Z({ w[58] })
);
BUF_X1 #() 
BUF_X1_944_ (
  .A({ S25957[580] }),
  .Z({ w[580] })
);
BUF_X1 #() 
BUF_X1_945_ (
  .A({ S25957[581] }),
  .Z({ w[581] })
);
BUF_X1 #() 
BUF_X1_946_ (
  .A({ S25957[582] }),
  .Z({ w[582] })
);
BUF_X1 #() 
BUF_X1_947_ (
  .A({ S25957[583] }),
  .Z({ w[583] })
);
BUF_X1 #() 
BUF_X1_948_ (
  .A({ S25957[584] }),
  .Z({ w[584] })
);
BUF_X1 #() 
BUF_X1_949_ (
  .A({ S25957[585] }),
  .Z({ w[585] })
);
BUF_X1 #() 
BUF_X1_950_ (
  .A({ S25957[586] }),
  .Z({ w[586] })
);
BUF_X1 #() 
BUF_X1_951_ (
  .A({ S25957[587] }),
  .Z({ w[587] })
);
BUF_X1 #() 
BUF_X1_952_ (
  .A({ S25957[588] }),
  .Z({ w[588] })
);
BUF_X1 #() 
BUF_X1_953_ (
  .A({ S25957[589] }),
  .Z({ w[589] })
);
BUF_X1 #() 
BUF_X1_954_ (
  .A({ S25957[59] }),
  .Z({ w[59] })
);
BUF_X1 #() 
BUF_X1_955_ (
  .A({ S25957[590] }),
  .Z({ w[590] })
);
BUF_X1 #() 
BUF_X1_956_ (
  .A({ S25957[591] }),
  .Z({ w[591] })
);
BUF_X1 #() 
BUF_X1_957_ (
  .A({ S25957[592] }),
  .Z({ w[592] })
);
BUF_X1 #() 
BUF_X1_958_ (
  .A({ S25957[593] }),
  .Z({ w[593] })
);
BUF_X1 #() 
BUF_X1_959_ (
  .A({ S25957[594] }),
  .Z({ w[594] })
);
BUF_X1 #() 
BUF_X1_960_ (
  .A({ S25957[595] }),
  .Z({ w[595] })
);
BUF_X1 #() 
BUF_X1_961_ (
  .A({ S25957[596] }),
  .Z({ w[596] })
);
BUF_X1 #() 
BUF_X1_962_ (
  .A({ S25957[597] }),
  .Z({ w[597] })
);
BUF_X1 #() 
BUF_X1_963_ (
  .A({ S25957[598] }),
  .Z({ w[598] })
);
BUF_X1 #() 
BUF_X1_964_ (
  .A({ S25957[599] }),
  .Z({ w[599] })
);
BUF_X1 #() 
BUF_X1_965_ (
  .A({ S25957[6] }),
  .Z({ w[6] })
);
BUF_X1 #() 
BUF_X1_966_ (
  .A({ S25957[60] }),
  .Z({ w[60] })
);
BUF_X1 #() 
BUF_X1_967_ (
  .A({ S25957[600] }),
  .Z({ w[600] })
);
BUF_X1 #() 
BUF_X1_968_ (
  .A({ S25957[601] }),
  .Z({ w[601] })
);
BUF_X1 #() 
BUF_X1_969_ (
  .A({ S25957[602] }),
  .Z({ w[602] })
);
BUF_X1 #() 
BUF_X1_970_ (
  .A({ S25957[603] }),
  .Z({ w[603] })
);
BUF_X1 #() 
BUF_X1_971_ (
  .A({ S25957[604] }),
  .Z({ w[604] })
);
BUF_X1 #() 
BUF_X1_972_ (
  .A({ S25957[605] }),
  .Z({ w[605] })
);
BUF_X1 #() 
BUF_X1_973_ (
  .A({ S25957[606] }),
  .Z({ w[606] })
);
BUF_X1 #() 
BUF_X1_974_ (
  .A({ S25957[607] }),
  .Z({ w[607] })
);
BUF_X1 #() 
BUF_X1_975_ (
  .A({ S25957[608] }),
  .Z({ w[608] })
);
BUF_X1 #() 
BUF_X1_976_ (
  .A({ S25957[609] }),
  .Z({ w[609] })
);
BUF_X1 #() 
BUF_X1_977_ (
  .A({ S25957[61] }),
  .Z({ w[61] })
);
BUF_X1 #() 
BUF_X1_978_ (
  .A({ S25957[610] }),
  .Z({ w[610] })
);
BUF_X1 #() 
BUF_X1_979_ (
  .A({ S25957[611] }),
  .Z({ w[611] })
);
BUF_X1 #() 
BUF_X1_980_ (
  .A({ S25957[612] }),
  .Z({ w[612] })
);
BUF_X1 #() 
BUF_X1_981_ (
  .A({ S25957[613] }),
  .Z({ w[613] })
);
BUF_X1 #() 
BUF_X1_982_ (
  .A({ S25957[614] }),
  .Z({ w[614] })
);
BUF_X1 #() 
BUF_X1_983_ (
  .A({ S25957[615] }),
  .Z({ w[615] })
);
BUF_X1 #() 
BUF_X1_984_ (
  .A({ S25957[616] }),
  .Z({ w[616] })
);
BUF_X1 #() 
BUF_X1_985_ (
  .A({ S25957[617] }),
  .Z({ w[617] })
);
BUF_X1 #() 
BUF_X1_986_ (
  .A({ S25957[618] }),
  .Z({ w[618] })
);
BUF_X1 #() 
BUF_X1_987_ (
  .A({ S25957[619] }),
  .Z({ w[619] })
);
BUF_X1 #() 
BUF_X1_988_ (
  .A({ S25957[62] }),
  .Z({ w[62] })
);
BUF_X1 #() 
BUF_X1_989_ (
  .A({ S25957[620] }),
  .Z({ w[620] })
);
BUF_X1 #() 
BUF_X1_990_ (
  .A({ S25957[621] }),
  .Z({ w[621] })
);
BUF_X1 #() 
BUF_X1_991_ (
  .A({ S25957[622] }),
  .Z({ w[622] })
);
BUF_X1 #() 
BUF_X1_992_ (
  .A({ S25957[623] }),
  .Z({ w[623] })
);
BUF_X1 #() 
BUF_X1_993_ (
  .A({ S25957[624] }),
  .Z({ w[624] })
);
BUF_X1 #() 
BUF_X1_994_ (
  .A({ S25957[625] }),
  .Z({ w[625] })
);
BUF_X1 #() 
BUF_X1_995_ (
  .A({ S25957[626] }),
  .Z({ w[626] })
);
BUF_X1 #() 
BUF_X1_996_ (
  .A({ S25957[627] }),
  .Z({ w[627] })
);
BUF_X1 #() 
BUF_X1_997_ (
  .A({ S25957[628] }),
  .Z({ w[628] })
);
BUF_X1 #() 
BUF_X1_998_ (
  .A({ S25957[629] }),
  .Z({ w[629] })
);
BUF_X1 #() 
BUF_X1_999_ (
  .A({ S25957[63] }),
  .Z({ w[63] })
);
BUF_X1 #() 
BUF_X1_1000_ (
  .A({ S25957[630] }),
  .Z({ w[630] })
);
BUF_X1 #() 
BUF_X1_1001_ (
  .A({ S25957[631] }),
  .Z({ w[631] })
);
BUF_X1 #() 
BUF_X1_1002_ (
  .A({ S25957[632] }),
  .Z({ w[632] })
);
BUF_X1 #() 
BUF_X1_1003_ (
  .A({ S25957[633] }),
  .Z({ w[633] })
);
BUF_X1 #() 
BUF_X1_1004_ (
  .A({ S25957[634] }),
  .Z({ w[634] })
);
BUF_X1 #() 
BUF_X1_1005_ (
  .A({ S25957[635] }),
  .Z({ w[635] })
);
BUF_X1 #() 
BUF_X1_1006_ (
  .A({ S25957[636] }),
  .Z({ w[636] })
);
BUF_X1 #() 
BUF_X1_1007_ (
  .A({ S25957[637] }),
  .Z({ w[637] })
);
BUF_X1 #() 
BUF_X1_1008_ (
  .A({ S25957[638] }),
  .Z({ w[638] })
);
BUF_X1 #() 
BUF_X1_1009_ (
  .A({ S25957[639] }),
  .Z({ w[639] })
);
BUF_X1 #() 
BUF_X1_1010_ (
  .A({ S25957[64] }),
  .Z({ w[64] })
);
BUF_X1 #() 
BUF_X1_1011_ (
  .A({ S25957[640] }),
  .Z({ w[640] })
);
BUF_X1 #() 
BUF_X1_1012_ (
  .A({ S25957[641] }),
  .Z({ w[641] })
);
BUF_X1 #() 
BUF_X1_1013_ (
  .A({ S25957[642] }),
  .Z({ w[642] })
);
BUF_X1 #() 
BUF_X1_1014_ (
  .A({ S25957[643] }),
  .Z({ w[643] })
);
BUF_X1 #() 
BUF_X1_1015_ (
  .A({ S25957[644] }),
  .Z({ w[644] })
);
BUF_X1 #() 
BUF_X1_1016_ (
  .A({ S25957[645] }),
  .Z({ w[645] })
);
BUF_X1 #() 
BUF_X1_1017_ (
  .A({ S25957[646] }),
  .Z({ w[646] })
);
BUF_X1 #() 
BUF_X1_1018_ (
  .A({ S25957[647] }),
  .Z({ w[647] })
);
BUF_X1 #() 
BUF_X1_1019_ (
  .A({ S25957[648] }),
  .Z({ w[648] })
);
BUF_X1 #() 
BUF_X1_1020_ (
  .A({ S25957[649] }),
  .Z({ w[649] })
);
BUF_X1 #() 
BUF_X1_1021_ (
  .A({ S25957[65] }),
  .Z({ w[65] })
);
BUF_X1 #() 
BUF_X1_1022_ (
  .A({ S25957[650] }),
  .Z({ w[650] })
);
BUF_X1 #() 
BUF_X1_1023_ (
  .A({ S25957[651] }),
  .Z({ w[651] })
);
BUF_X1 #() 
BUF_X1_1024_ (
  .A({ S25957[652] }),
  .Z({ w[652] })
);
BUF_X1 #() 
BUF_X1_1025_ (
  .A({ S25957[653] }),
  .Z({ w[653] })
);
BUF_X1 #() 
BUF_X1_1026_ (
  .A({ S25957[654] }),
  .Z({ w[654] })
);
BUF_X1 #() 
BUF_X1_1027_ (
  .A({ S25957[655] }),
  .Z({ w[655] })
);
BUF_X1 #() 
BUF_X1_1028_ (
  .A({ S25957[656] }),
  .Z({ w[656] })
);
BUF_X1 #() 
BUF_X1_1029_ (
  .A({ S25957[657] }),
  .Z({ w[657] })
);
BUF_X1 #() 
BUF_X1_1030_ (
  .A({ S25957[658] }),
  .Z({ w[658] })
);
BUF_X1 #() 
BUF_X1_1031_ (
  .A({ S25957[659] }),
  .Z({ w[659] })
);
BUF_X1 #() 
BUF_X1_1032_ (
  .A({ S25957[66] }),
  .Z({ w[66] })
);
BUF_X1 #() 
BUF_X1_1033_ (
  .A({ S25957[660] }),
  .Z({ w[660] })
);
BUF_X1 #() 
BUF_X1_1034_ (
  .A({ S25957[661] }),
  .Z({ w[661] })
);
BUF_X1 #() 
BUF_X1_1035_ (
  .A({ S25957[662] }),
  .Z({ w[662] })
);
BUF_X1 #() 
BUF_X1_1036_ (
  .A({ S25957[663] }),
  .Z({ w[663] })
);
BUF_X1 #() 
BUF_X1_1037_ (
  .A({ S25957[664] }),
  .Z({ w[664] })
);
BUF_X1 #() 
BUF_X1_1038_ (
  .A({ S25957[665] }),
  .Z({ w[665] })
);
BUF_X1 #() 
BUF_X1_1039_ (
  .A({ S25957[666] }),
  .Z({ w[666] })
);
BUF_X1 #() 
BUF_X1_1040_ (
  .A({ S25957[667] }),
  .Z({ w[667] })
);
BUF_X1 #() 
BUF_X1_1041_ (
  .A({ S25957[668] }),
  .Z({ w[668] })
);
BUF_X1 #() 
BUF_X1_1042_ (
  .A({ S25957[669] }),
  .Z({ w[669] })
);
BUF_X1 #() 
BUF_X1_1043_ (
  .A({ S25957[67] }),
  .Z({ w[67] })
);
BUF_X1 #() 
BUF_X1_1044_ (
  .A({ S25957[670] }),
  .Z({ w[670] })
);
BUF_X1 #() 
BUF_X1_1045_ (
  .A({ S25957[671] }),
  .Z({ w[671] })
);
BUF_X1 #() 
BUF_X1_1046_ (
  .A({ S25957[672] }),
  .Z({ w[672] })
);
BUF_X1 #() 
BUF_X1_1047_ (
  .A({ S25957[673] }),
  .Z({ w[673] })
);
BUF_X1 #() 
BUF_X1_1048_ (
  .A({ S25957[674] }),
  .Z({ w[674] })
);
BUF_X1 #() 
BUF_X1_1049_ (
  .A({ S25957[675] }),
  .Z({ w[675] })
);
BUF_X1 #() 
BUF_X1_1050_ (
  .A({ S25957[676] }),
  .Z({ w[676] })
);
BUF_X1 #() 
BUF_X1_1051_ (
  .A({ S25957[677] }),
  .Z({ w[677] })
);
BUF_X1 #() 
BUF_X1_1052_ (
  .A({ S25957[678] }),
  .Z({ w[678] })
);
BUF_X1 #() 
BUF_X1_1053_ (
  .A({ S25957[679] }),
  .Z({ w[679] })
);
BUF_X1 #() 
BUF_X1_1054_ (
  .A({ S25957[68] }),
  .Z({ w[68] })
);
BUF_X1 #() 
BUF_X1_1055_ (
  .A({ S25957[680] }),
  .Z({ w[680] })
);
BUF_X1 #() 
BUF_X1_1056_ (
  .A({ S25957[681] }),
  .Z({ w[681] })
);
BUF_X1 #() 
BUF_X1_1057_ (
  .A({ S25957[682] }),
  .Z({ w[682] })
);
BUF_X1 #() 
BUF_X1_1058_ (
  .A({ S25957[683] }),
  .Z({ w[683] })
);
BUF_X1 #() 
BUF_X1_1059_ (
  .A({ S25957[684] }),
  .Z({ w[684] })
);
BUF_X1 #() 
BUF_X1_1060_ (
  .A({ S25957[685] }),
  .Z({ w[685] })
);
BUF_X1 #() 
BUF_X1_1061_ (
  .A({ S25957[686] }),
  .Z({ w[686] })
);
BUF_X1 #() 
BUF_X1_1062_ (
  .A({ S25957[687] }),
  .Z({ w[687] })
);
BUF_X1 #() 
BUF_X1_1063_ (
  .A({ S25957[688] }),
  .Z({ w[688] })
);
BUF_X1 #() 
BUF_X1_1064_ (
  .A({ S25957[689] }),
  .Z({ w[689] })
);
BUF_X1 #() 
BUF_X1_1065_ (
  .A({ S25957[69] }),
  .Z({ w[69] })
);
BUF_X1 #() 
BUF_X1_1066_ (
  .A({ S25957[690] }),
  .Z({ w[690] })
);
BUF_X1 #() 
BUF_X1_1067_ (
  .A({ S25957[691] }),
  .Z({ w[691] })
);
BUF_X1 #() 
BUF_X1_1068_ (
  .A({ S25957[692] }),
  .Z({ w[692] })
);
BUF_X1 #() 
BUF_X1_1069_ (
  .A({ S25957[693] }),
  .Z({ w[693] })
);
BUF_X1 #() 
BUF_X1_1070_ (
  .A({ S25957[694] }),
  .Z({ w[694] })
);
BUF_X1 #() 
BUF_X1_1071_ (
  .A({ S25957[695] }),
  .Z({ w[695] })
);
BUF_X1 #() 
BUF_X1_1072_ (
  .A({ S25957[696] }),
  .Z({ w[696] })
);
BUF_X1 #() 
BUF_X1_1073_ (
  .A({ S25957[697] }),
  .Z({ w[697] })
);
BUF_X1 #() 
BUF_X1_1074_ (
  .A({ S25957[698] }),
  .Z({ w[698] })
);
BUF_X1 #() 
BUF_X1_1075_ (
  .A({ S25957[699] }),
  .Z({ w[699] })
);
BUF_X1 #() 
BUF_X1_1076_ (
  .A({ S25957[7] }),
  .Z({ w[7] })
);
BUF_X1 #() 
BUF_X1_1077_ (
  .A({ S25957[70] }),
  .Z({ w[70] })
);
BUF_X1 #() 
BUF_X1_1078_ (
  .A({ S25957[700] }),
  .Z({ w[700] })
);
BUF_X1 #() 
BUF_X1_1079_ (
  .A({ S25957[701] }),
  .Z({ w[701] })
);
BUF_X1 #() 
BUF_X1_1080_ (
  .A({ S25957[702] }),
  .Z({ w[702] })
);
BUF_X1 #() 
BUF_X1_1081_ (
  .A({ S25957[703] }),
  .Z({ w[703] })
);
BUF_X1 #() 
BUF_X1_1082_ (
  .A({ S25957[704] }),
  .Z({ w[704] })
);
BUF_X1 #() 
BUF_X1_1083_ (
  .A({ S25957[705] }),
  .Z({ w[705] })
);
BUF_X1 #() 
BUF_X1_1084_ (
  .A({ S25957[706] }),
  .Z({ w[706] })
);
BUF_X1 #() 
BUF_X1_1085_ (
  .A({ S25957[707] }),
  .Z({ w[707] })
);
BUF_X1 #() 
BUF_X1_1086_ (
  .A({ S25957[708] }),
  .Z({ w[708] })
);
BUF_X1 #() 
BUF_X1_1087_ (
  .A({ S25957[709] }),
  .Z({ w[709] })
);
BUF_X1 #() 
BUF_X1_1088_ (
  .A({ S25957[71] }),
  .Z({ w[71] })
);
BUF_X1 #() 
BUF_X1_1089_ (
  .A({ S25957[710] }),
  .Z({ w[710] })
);
BUF_X1 #() 
BUF_X1_1090_ (
  .A({ S25957[711] }),
  .Z({ w[711] })
);
BUF_X1 #() 
BUF_X1_1091_ (
  .A({ S25957[712] }),
  .Z({ w[712] })
);
BUF_X1 #() 
BUF_X1_1092_ (
  .A({ S25957[713] }),
  .Z({ w[713] })
);
BUF_X1 #() 
BUF_X1_1093_ (
  .A({ S25957[714] }),
  .Z({ w[714] })
);
BUF_X1 #() 
BUF_X1_1094_ (
  .A({ S25957[715] }),
  .Z({ w[715] })
);
BUF_X1 #() 
BUF_X1_1095_ (
  .A({ S25957[716] }),
  .Z({ w[716] })
);
BUF_X1 #() 
BUF_X1_1096_ (
  .A({ S25957[717] }),
  .Z({ w[717] })
);
BUF_X1 #() 
BUF_X1_1097_ (
  .A({ S25957[718] }),
  .Z({ w[718] })
);
BUF_X1 #() 
BUF_X1_1098_ (
  .A({ S25957[719] }),
  .Z({ w[719] })
);
BUF_X1 #() 
BUF_X1_1099_ (
  .A({ S25957[72] }),
  .Z({ w[72] })
);
BUF_X1 #() 
BUF_X1_1100_ (
  .A({ S25957[720] }),
  .Z({ w[720] })
);
BUF_X1 #() 
BUF_X1_1101_ (
  .A({ S25957[721] }),
  .Z({ w[721] })
);
BUF_X1 #() 
BUF_X1_1102_ (
  .A({ S25957[722] }),
  .Z({ w[722] })
);
BUF_X1 #() 
BUF_X1_1103_ (
  .A({ S25957[723] }),
  .Z({ w[723] })
);
BUF_X1 #() 
BUF_X1_1104_ (
  .A({ S25957[724] }),
  .Z({ w[724] })
);
BUF_X1 #() 
BUF_X1_1105_ (
  .A({ S25957[725] }),
  .Z({ w[725] })
);
BUF_X1 #() 
BUF_X1_1106_ (
  .A({ S25957[726] }),
  .Z({ w[726] })
);
BUF_X1 #() 
BUF_X1_1107_ (
  .A({ S25957[727] }),
  .Z({ w[727] })
);
BUF_X1 #() 
BUF_X1_1108_ (
  .A({ S25957[728] }),
  .Z({ w[728] })
);
BUF_X1 #() 
BUF_X1_1109_ (
  .A({ S25957[729] }),
  .Z({ w[729] })
);
BUF_X1 #() 
BUF_X1_1110_ (
  .A({ S25957[73] }),
  .Z({ w[73] })
);
BUF_X1 #() 
BUF_X1_1111_ (
  .A({ S25957[730] }),
  .Z({ w[730] })
);
BUF_X1 #() 
BUF_X1_1112_ (
  .A({ S25957[731] }),
  .Z({ w[731] })
);
BUF_X1 #() 
BUF_X1_1113_ (
  .A({ S25957[732] }),
  .Z({ w[732] })
);
BUF_X1 #() 
BUF_X1_1114_ (
  .A({ S25957[733] }),
  .Z({ w[733] })
);
BUF_X1 #() 
BUF_X1_1115_ (
  .A({ S25957[734] }),
  .Z({ w[734] })
);
BUF_X1 #() 
BUF_X1_1116_ (
  .A({ S25957[735] }),
  .Z({ w[735] })
);
BUF_X1 #() 
BUF_X1_1117_ (
  .A({ S25957[736] }),
  .Z({ w[736] })
);
BUF_X1 #() 
BUF_X1_1118_ (
  .A({ S25957[737] }),
  .Z({ w[737] })
);
BUF_X1 #() 
BUF_X1_1119_ (
  .A({ S25957[738] }),
  .Z({ w[738] })
);
BUF_X1 #() 
BUF_X1_1120_ (
  .A({ S25957[739] }),
  .Z({ w[739] })
);
BUF_X1 #() 
BUF_X1_1121_ (
  .A({ S25957[74] }),
  .Z({ w[74] })
);
BUF_X1 #() 
BUF_X1_1122_ (
  .A({ S25957[740] }),
  .Z({ w[740] })
);
BUF_X1 #() 
BUF_X1_1123_ (
  .A({ S25957[741] }),
  .Z({ w[741] })
);
BUF_X1 #() 
BUF_X1_1124_ (
  .A({ S25957[742] }),
  .Z({ w[742] })
);
BUF_X1 #() 
BUF_X1_1125_ (
  .A({ S25957[743] }),
  .Z({ w[743] })
);
BUF_X1 #() 
BUF_X1_1126_ (
  .A({ S25957[744] }),
  .Z({ w[744] })
);
BUF_X1 #() 
BUF_X1_1127_ (
  .A({ S25957[745] }),
  .Z({ w[745] })
);
BUF_X1 #() 
BUF_X1_1128_ (
  .A({ S25957[746] }),
  .Z({ w[746] })
);
BUF_X1 #() 
BUF_X1_1129_ (
  .A({ S25957[747] }),
  .Z({ w[747] })
);
BUF_X1 #() 
BUF_X1_1130_ (
  .A({ S25957[748] }),
  .Z({ w[748] })
);
BUF_X1 #() 
BUF_X1_1131_ (
  .A({ S25957[749] }),
  .Z({ w[749] })
);
BUF_X1 #() 
BUF_X1_1132_ (
  .A({ S25957[75] }),
  .Z({ w[75] })
);
BUF_X1 #() 
BUF_X1_1133_ (
  .A({ S25957[750] }),
  .Z({ w[750] })
);
BUF_X1 #() 
BUF_X1_1134_ (
  .A({ S25957[751] }),
  .Z({ w[751] })
);
BUF_X1 #() 
BUF_X1_1135_ (
  .A({ S25957[752] }),
  .Z({ w[752] })
);
BUF_X1 #() 
BUF_X1_1136_ (
  .A({ S25957[753] }),
  .Z({ w[753] })
);
BUF_X1 #() 
BUF_X1_1137_ (
  .A({ S25957[754] }),
  .Z({ w[754] })
);
BUF_X1 #() 
BUF_X1_1138_ (
  .A({ S25957[755] }),
  .Z({ w[755] })
);
BUF_X1 #() 
BUF_X1_1139_ (
  .A({ S25957[756] }),
  .Z({ w[756] })
);
BUF_X1 #() 
BUF_X1_1140_ (
  .A({ S25957[757] }),
  .Z({ w[757] })
);
BUF_X1 #() 
BUF_X1_1141_ (
  .A({ S25957[758] }),
  .Z({ w[758] })
);
BUF_X1 #() 
BUF_X1_1142_ (
  .A({ S25957[759] }),
  .Z({ w[759] })
);
BUF_X1 #() 
BUF_X1_1143_ (
  .A({ S25957[76] }),
  .Z({ w[76] })
);
BUF_X1 #() 
BUF_X1_1144_ (
  .A({ S25957[760] }),
  .Z({ w[760] })
);
BUF_X1 #() 
BUF_X1_1145_ (
  .A({ S25957[761] }),
  .Z({ w[761] })
);
BUF_X1 #() 
BUF_X1_1146_ (
  .A({ S25957[762] }),
  .Z({ w[762] })
);
BUF_X1 #() 
BUF_X1_1147_ (
  .A({ S25957[763] }),
  .Z({ w[763] })
);
BUF_X1 #() 
BUF_X1_1148_ (
  .A({ S25957[764] }),
  .Z({ w[764] })
);
BUF_X1 #() 
BUF_X1_1149_ (
  .A({ S25957[765] }),
  .Z({ w[765] })
);
BUF_X1 #() 
BUF_X1_1150_ (
  .A({ S25957[766] }),
  .Z({ w[766] })
);
BUF_X1 #() 
BUF_X1_1151_ (
  .A({ S25957[767] }),
  .Z({ w[767] })
);
BUF_X1 #() 
BUF_X1_1152_ (
  .A({ S25957[768] }),
  .Z({ w[768] })
);
BUF_X1 #() 
BUF_X1_1153_ (
  .A({ S25957[769] }),
  .Z({ w[769] })
);
BUF_X1 #() 
BUF_X1_1154_ (
  .A({ S25957[77] }),
  .Z({ w[77] })
);
BUF_X1 #() 
BUF_X1_1155_ (
  .A({ S25957[770] }),
  .Z({ w[770] })
);
BUF_X1 #() 
BUF_X1_1156_ (
  .A({ S25957[771] }),
  .Z({ w[771] })
);
BUF_X1 #() 
BUF_X1_1157_ (
  .A({ S25957[772] }),
  .Z({ w[772] })
);
BUF_X1 #() 
BUF_X1_1158_ (
  .A({ S25957[773] }),
  .Z({ w[773] })
);
BUF_X1 #() 
BUF_X1_1159_ (
  .A({ S25957[774] }),
  .Z({ w[774] })
);
BUF_X1 #() 
BUF_X1_1160_ (
  .A({ S25957[775] }),
  .Z({ w[775] })
);
BUF_X1 #() 
BUF_X1_1161_ (
  .A({ S25957[776] }),
  .Z({ w[776] })
);
BUF_X1 #() 
BUF_X1_1162_ (
  .A({ S25957[777] }),
  .Z({ w[777] })
);
BUF_X1 #() 
BUF_X1_1163_ (
  .A({ S25957[778] }),
  .Z({ w[778] })
);
BUF_X1 #() 
BUF_X1_1164_ (
  .A({ S25957[779] }),
  .Z({ w[779] })
);
BUF_X1 #() 
BUF_X1_1165_ (
  .A({ S25957[78] }),
  .Z({ w[78] })
);
BUF_X1 #() 
BUF_X1_1166_ (
  .A({ S25957[780] }),
  .Z({ w[780] })
);
BUF_X1 #() 
BUF_X1_1167_ (
  .A({ S25957[781] }),
  .Z({ w[781] })
);
BUF_X1 #() 
BUF_X1_1168_ (
  .A({ S25957[782] }),
  .Z({ w[782] })
);
BUF_X1 #() 
BUF_X1_1169_ (
  .A({ S25957[783] }),
  .Z({ w[783] })
);
BUF_X1 #() 
BUF_X1_1170_ (
  .A({ S25957[784] }),
  .Z({ w[784] })
);
BUF_X1 #() 
BUF_X1_1171_ (
  .A({ S25957[785] }),
  .Z({ w[785] })
);
BUF_X1 #() 
BUF_X1_1172_ (
  .A({ S25957[786] }),
  .Z({ w[786] })
);
BUF_X1 #() 
BUF_X1_1173_ (
  .A({ S25957[787] }),
  .Z({ w[787] })
);
BUF_X1 #() 
BUF_X1_1174_ (
  .A({ S25957[788] }),
  .Z({ w[788] })
);
BUF_X1 #() 
BUF_X1_1175_ (
  .A({ S25957[789] }),
  .Z({ w[789] })
);
BUF_X1 #() 
BUF_X1_1176_ (
  .A({ S25957[79] }),
  .Z({ w[79] })
);
BUF_X1 #() 
BUF_X1_1177_ (
  .A({ S25957[790] }),
  .Z({ w[790] })
);
BUF_X1 #() 
BUF_X1_1178_ (
  .A({ S25957[791] }),
  .Z({ w[791] })
);
BUF_X1 #() 
BUF_X1_1179_ (
  .A({ S25957[792] }),
  .Z({ w[792] })
);
BUF_X1 #() 
BUF_X1_1180_ (
  .A({ S25957[793] }),
  .Z({ w[793] })
);
BUF_X1 #() 
BUF_X1_1181_ (
  .A({ S25957[794] }),
  .Z({ w[794] })
);
BUF_X1 #() 
BUF_X1_1182_ (
  .A({ S25957[795] }),
  .Z({ w[795] })
);
BUF_X1 #() 
BUF_X1_1183_ (
  .A({ S25957[796] }),
  .Z({ w[796] })
);
BUF_X1 #() 
BUF_X1_1184_ (
  .A({ S25957[797] }),
  .Z({ w[797] })
);
BUF_X1 #() 
BUF_X1_1185_ (
  .A({ S25957[798] }),
  .Z({ w[798] })
);
BUF_X1 #() 
BUF_X1_1186_ (
  .A({ S25957[799] }),
  .Z({ w[799] })
);
BUF_X1 #() 
BUF_X1_1187_ (
  .A({ S25957[8] }),
  .Z({ w[8] })
);
BUF_X1 #() 
BUF_X1_1188_ (
  .A({ S25957[80] }),
  .Z({ w[80] })
);
BUF_X1 #() 
BUF_X1_1189_ (
  .A({ S25957[800] }),
  .Z({ w[800] })
);
BUF_X1 #() 
BUF_X1_1190_ (
  .A({ S25957[801] }),
  .Z({ w[801] })
);
BUF_X1 #() 
BUF_X1_1191_ (
  .A({ S25957[802] }),
  .Z({ w[802] })
);
BUF_X1 #() 
BUF_X1_1192_ (
  .A({ S25957[803] }),
  .Z({ w[803] })
);
BUF_X1 #() 
BUF_X1_1193_ (
  .A({ S25957[804] }),
  .Z({ w[804] })
);
BUF_X1 #() 
BUF_X1_1194_ (
  .A({ S25957[805] }),
  .Z({ w[805] })
);
BUF_X1 #() 
BUF_X1_1195_ (
  .A({ S25957[806] }),
  .Z({ w[806] })
);
BUF_X1 #() 
BUF_X1_1196_ (
  .A({ S25957[807] }),
  .Z({ w[807] })
);
BUF_X1 #() 
BUF_X1_1197_ (
  .A({ S25957[808] }),
  .Z({ w[808] })
);
BUF_X1 #() 
BUF_X1_1198_ (
  .A({ S25957[809] }),
  .Z({ w[809] })
);
BUF_X1 #() 
BUF_X1_1199_ (
  .A({ S25957[81] }),
  .Z({ w[81] })
);
BUF_X1 #() 
BUF_X1_1200_ (
  .A({ S25957[810] }),
  .Z({ w[810] })
);
BUF_X1 #() 
BUF_X1_1201_ (
  .A({ S25957[811] }),
  .Z({ w[811] })
);
BUF_X1 #() 
BUF_X1_1202_ (
  .A({ S25957[812] }),
  .Z({ w[812] })
);
BUF_X1 #() 
BUF_X1_1203_ (
  .A({ S25957[813] }),
  .Z({ w[813] })
);
BUF_X1 #() 
BUF_X1_1204_ (
  .A({ S25957[814] }),
  .Z({ w[814] })
);
BUF_X1 #() 
BUF_X1_1205_ (
  .A({ S25957[815] }),
  .Z({ w[815] })
);
BUF_X1 #() 
BUF_X1_1206_ (
  .A({ S25957[816] }),
  .Z({ w[816] })
);
BUF_X1 #() 
BUF_X1_1207_ (
  .A({ S25957[817] }),
  .Z({ w[817] })
);
BUF_X1 #() 
BUF_X1_1208_ (
  .A({ S25957[818] }),
  .Z({ w[818] })
);
BUF_X1 #() 
BUF_X1_1209_ (
  .A({ S25957[819] }),
  .Z({ w[819] })
);
BUF_X1 #() 
BUF_X1_1210_ (
  .A({ S25957[82] }),
  .Z({ w[82] })
);
BUF_X1 #() 
BUF_X1_1211_ (
  .A({ S25957[820] }),
  .Z({ w[820] })
);
BUF_X1 #() 
BUF_X1_1212_ (
  .A({ S25957[821] }),
  .Z({ w[821] })
);
BUF_X1 #() 
BUF_X1_1213_ (
  .A({ S25957[822] }),
  .Z({ w[822] })
);
BUF_X1 #() 
BUF_X1_1214_ (
  .A({ S25957[823] }),
  .Z({ w[823] })
);
BUF_X1 #() 
BUF_X1_1215_ (
  .A({ S25957[824] }),
  .Z({ w[824] })
);
BUF_X1 #() 
BUF_X1_1216_ (
  .A({ S25957[825] }),
  .Z({ w[825] })
);
BUF_X1 #() 
BUF_X1_1217_ (
  .A({ S25957[826] }),
  .Z({ w[826] })
);
BUF_X1 #() 
BUF_X1_1218_ (
  .A({ S25957[827] }),
  .Z({ w[827] })
);
BUF_X1 #() 
BUF_X1_1219_ (
  .A({ S25957[828] }),
  .Z({ w[828] })
);
BUF_X1 #() 
BUF_X1_1220_ (
  .A({ S25957[829] }),
  .Z({ w[829] })
);
BUF_X1 #() 
BUF_X1_1221_ (
  .A({ S25957[83] }),
  .Z({ w[83] })
);
BUF_X1 #() 
BUF_X1_1222_ (
  .A({ S25957[830] }),
  .Z({ w[830] })
);
BUF_X1 #() 
BUF_X1_1223_ (
  .A({ S25957[831] }),
  .Z({ w[831] })
);
BUF_X1 #() 
BUF_X1_1224_ (
  .A({ S25957[832] }),
  .Z({ w[832] })
);
BUF_X1 #() 
BUF_X1_1225_ (
  .A({ S25957[833] }),
  .Z({ w[833] })
);
BUF_X1 #() 
BUF_X1_1226_ (
  .A({ S25957[834] }),
  .Z({ w[834] })
);
BUF_X1 #() 
BUF_X1_1227_ (
  .A({ S25957[835] }),
  .Z({ w[835] })
);
BUF_X1 #() 
BUF_X1_1228_ (
  .A({ S25957[836] }),
  .Z({ w[836] })
);
BUF_X1 #() 
BUF_X1_1229_ (
  .A({ S25957[837] }),
  .Z({ w[837] })
);
BUF_X1 #() 
BUF_X1_1230_ (
  .A({ S25957[838] }),
  .Z({ w[838] })
);
BUF_X1 #() 
BUF_X1_1231_ (
  .A({ S25957[839] }),
  .Z({ w[839] })
);
BUF_X1 #() 
BUF_X1_1232_ (
  .A({ S25957[84] }),
  .Z({ w[84] })
);
BUF_X1 #() 
BUF_X1_1233_ (
  .A({ S25957[840] }),
  .Z({ w[840] })
);
BUF_X1 #() 
BUF_X1_1234_ (
  .A({ S25957[841] }),
  .Z({ w[841] })
);
BUF_X1 #() 
BUF_X1_1235_ (
  .A({ S25957[842] }),
  .Z({ w[842] })
);
BUF_X1 #() 
BUF_X1_1236_ (
  .A({ S25957[843] }),
  .Z({ w[843] })
);
BUF_X1 #() 
BUF_X1_1237_ (
  .A({ S25957[844] }),
  .Z({ w[844] })
);
BUF_X1 #() 
BUF_X1_1238_ (
  .A({ S25957[845] }),
  .Z({ w[845] })
);
BUF_X1 #() 
BUF_X1_1239_ (
  .A({ S25957[846] }),
  .Z({ w[846] })
);
BUF_X1 #() 
BUF_X1_1240_ (
  .A({ S25957[847] }),
  .Z({ w[847] })
);
BUF_X1 #() 
BUF_X1_1241_ (
  .A({ S25957[848] }),
  .Z({ w[848] })
);
BUF_X1 #() 
BUF_X1_1242_ (
  .A({ S25957[849] }),
  .Z({ w[849] })
);
BUF_X1 #() 
BUF_X1_1243_ (
  .A({ S25957[85] }),
  .Z({ w[85] })
);
BUF_X1 #() 
BUF_X1_1244_ (
  .A({ S25957[850] }),
  .Z({ w[850] })
);
BUF_X1 #() 
BUF_X1_1245_ (
  .A({ S25957[851] }),
  .Z({ w[851] })
);
BUF_X1 #() 
BUF_X1_1246_ (
  .A({ S25957[852] }),
  .Z({ w[852] })
);
BUF_X1 #() 
BUF_X1_1247_ (
  .A({ S25957[853] }),
  .Z({ w[853] })
);
BUF_X1 #() 
BUF_X1_1248_ (
  .A({ S25957[854] }),
  .Z({ w[854] })
);
BUF_X1 #() 
BUF_X1_1249_ (
  .A({ S25957[855] }),
  .Z({ w[855] })
);
BUF_X1 #() 
BUF_X1_1250_ (
  .A({ S25957[856] }),
  .Z({ w[856] })
);
BUF_X1 #() 
BUF_X1_1251_ (
  .A({ S25957[857] }),
  .Z({ w[857] })
);
BUF_X1 #() 
BUF_X1_1252_ (
  .A({ S25957[858] }),
  .Z({ w[858] })
);
BUF_X1 #() 
BUF_X1_1253_ (
  .A({ S25957[859] }),
  .Z({ w[859] })
);
BUF_X1 #() 
BUF_X1_1254_ (
  .A({ S25957[86] }),
  .Z({ w[86] })
);
BUF_X1 #() 
BUF_X1_1255_ (
  .A({ S25957[860] }),
  .Z({ w[860] })
);
BUF_X1 #() 
BUF_X1_1256_ (
  .A({ S25957[861] }),
  .Z({ w[861] })
);
BUF_X1 #() 
BUF_X1_1257_ (
  .A({ S25957[862] }),
  .Z({ w[862] })
);
BUF_X1 #() 
BUF_X1_1258_ (
  .A({ S25957[863] }),
  .Z({ w[863] })
);
BUF_X1 #() 
BUF_X1_1259_ (
  .A({ S25957[864] }),
  .Z({ w[864] })
);
BUF_X1 #() 
BUF_X1_1260_ (
  .A({ S25957[865] }),
  .Z({ w[865] })
);
BUF_X1 #() 
BUF_X1_1261_ (
  .A({ S25957[866] }),
  .Z({ w[866] })
);
BUF_X1 #() 
BUF_X1_1262_ (
  .A({ S25957[867] }),
  .Z({ w[867] })
);
BUF_X1 #() 
BUF_X1_1263_ (
  .A({ S25957[868] }),
  .Z({ w[868] })
);
BUF_X1 #() 
BUF_X1_1264_ (
  .A({ S25957[869] }),
  .Z({ w[869] })
);
BUF_X1 #() 
BUF_X1_1265_ (
  .A({ S25957[87] }),
  .Z({ w[87] })
);
BUF_X1 #() 
BUF_X1_1266_ (
  .A({ S25957[870] }),
  .Z({ w[870] })
);
BUF_X1 #() 
BUF_X1_1267_ (
  .A({ S25957[871] }),
  .Z({ w[871] })
);
BUF_X1 #() 
BUF_X1_1268_ (
  .A({ S25957[872] }),
  .Z({ w[872] })
);
BUF_X1 #() 
BUF_X1_1269_ (
  .A({ S25957[873] }),
  .Z({ w[873] })
);
BUF_X1 #() 
BUF_X1_1270_ (
  .A({ S25957[874] }),
  .Z({ w[874] })
);
BUF_X1 #() 
BUF_X1_1271_ (
  .A({ S25957[875] }),
  .Z({ w[875] })
);
BUF_X1 #() 
BUF_X1_1272_ (
  .A({ S25957[876] }),
  .Z({ w[876] })
);
BUF_X1 #() 
BUF_X1_1273_ (
  .A({ S25957[877] }),
  .Z({ w[877] })
);
BUF_X1 #() 
BUF_X1_1274_ (
  .A({ S25957[878] }),
  .Z({ w[878] })
);
BUF_X1 #() 
BUF_X1_1275_ (
  .A({ S25957[879] }),
  .Z({ w[879] })
);
BUF_X1 #() 
BUF_X1_1276_ (
  .A({ S25957[88] }),
  .Z({ w[88] })
);
BUF_X1 #() 
BUF_X1_1277_ (
  .A({ S25957[880] }),
  .Z({ w[880] })
);
BUF_X1 #() 
BUF_X1_1278_ (
  .A({ S25957[881] }),
  .Z({ w[881] })
);
BUF_X1 #() 
BUF_X1_1279_ (
  .A({ S25957[882] }),
  .Z({ w[882] })
);
BUF_X1 #() 
BUF_X1_1280_ (
  .A({ S25957[883] }),
  .Z({ w[883] })
);
BUF_X1 #() 
BUF_X1_1281_ (
  .A({ S25957[884] }),
  .Z({ w[884] })
);
BUF_X1 #() 
BUF_X1_1282_ (
  .A({ S25957[885] }),
  .Z({ w[885] })
);
BUF_X1 #() 
BUF_X1_1283_ (
  .A({ S25957[886] }),
  .Z({ w[886] })
);
BUF_X1 #() 
BUF_X1_1284_ (
  .A({ S25957[887] }),
  .Z({ w[887] })
);
BUF_X1 #() 
BUF_X1_1285_ (
  .A({ S25957[888] }),
  .Z({ w[888] })
);
BUF_X1 #() 
BUF_X1_1286_ (
  .A({ S25957[889] }),
  .Z({ w[889] })
);
BUF_X1 #() 
BUF_X1_1287_ (
  .A({ S25957[89] }),
  .Z({ w[89] })
);
BUF_X1 #() 
BUF_X1_1288_ (
  .A({ S25957[890] }),
  .Z({ w[890] })
);
BUF_X1 #() 
BUF_X1_1289_ (
  .A({ S25957[891] }),
  .Z({ w[891] })
);
BUF_X1 #() 
BUF_X1_1290_ (
  .A({ S25957[892] }),
  .Z({ w[892] })
);
BUF_X1 #() 
BUF_X1_1291_ (
  .A({ S25957[893] }),
  .Z({ w[893] })
);
BUF_X1 #() 
BUF_X1_1292_ (
  .A({ S25957[894] }),
  .Z({ w[894] })
);
BUF_X1 #() 
BUF_X1_1293_ (
  .A({ S25957[895] }),
  .Z({ w[895] })
);
BUF_X1 #() 
BUF_X1_1294_ (
  .A({ S25957[896] }),
  .Z({ w[896] })
);
BUF_X1 #() 
BUF_X1_1295_ (
  .A({ S25957[897] }),
  .Z({ w[897] })
);
BUF_X1 #() 
BUF_X1_1296_ (
  .A({ S25957[898] }),
  .Z({ w[898] })
);
BUF_X1 #() 
BUF_X1_1297_ (
  .A({ S25957[899] }),
  .Z({ w[899] })
);
BUF_X1 #() 
BUF_X1_1298_ (
  .A({ S25957[9] }),
  .Z({ w[9] })
);
BUF_X1 #() 
BUF_X1_1299_ (
  .A({ S25957[90] }),
  .Z({ w[90] })
);
BUF_X1 #() 
BUF_X1_1300_ (
  .A({ S25957[900] }),
  .Z({ w[900] })
);
BUF_X1 #() 
BUF_X1_1301_ (
  .A({ S25957[901] }),
  .Z({ w[901] })
);
BUF_X1 #() 
BUF_X1_1302_ (
  .A({ S25957[902] }),
  .Z({ w[902] })
);
BUF_X1 #() 
BUF_X1_1303_ (
  .A({ S25957[903] }),
  .Z({ w[903] })
);
BUF_X1 #() 
BUF_X1_1304_ (
  .A({ S25957[904] }),
  .Z({ w[904] })
);
BUF_X1 #() 
BUF_X1_1305_ (
  .A({ S25957[905] }),
  .Z({ w[905] })
);
BUF_X1 #() 
BUF_X1_1306_ (
  .A({ S25957[906] }),
  .Z({ w[906] })
);
BUF_X1 #() 
BUF_X1_1307_ (
  .A({ S25957[907] }),
  .Z({ w[907] })
);
BUF_X1 #() 
BUF_X1_1308_ (
  .A({ S25957[908] }),
  .Z({ w[908] })
);
BUF_X1 #() 
BUF_X1_1309_ (
  .A({ S25957[909] }),
  .Z({ w[909] })
);
BUF_X1 #() 
BUF_X1_1310_ (
  .A({ S25957[91] }),
  .Z({ w[91] })
);
BUF_X1 #() 
BUF_X1_1311_ (
  .A({ S25957[910] }),
  .Z({ w[910] })
);
BUF_X1 #() 
BUF_X1_1312_ (
  .A({ S25957[911] }),
  .Z({ w[911] })
);
BUF_X1 #() 
BUF_X1_1313_ (
  .A({ S25957[912] }),
  .Z({ w[912] })
);
BUF_X1 #() 
BUF_X1_1314_ (
  .A({ S25957[913] }),
  .Z({ w[913] })
);
BUF_X1 #() 
BUF_X1_1315_ (
  .A({ S25957[914] }),
  .Z({ w[914] })
);
BUF_X1 #() 
BUF_X1_1316_ (
  .A({ S25957[915] }),
  .Z({ w[915] })
);
BUF_X1 #() 
BUF_X1_1317_ (
  .A({ S25957[916] }),
  .Z({ w[916] })
);
BUF_X1 #() 
BUF_X1_1318_ (
  .A({ S25957[917] }),
  .Z({ w[917] })
);
BUF_X1 #() 
BUF_X1_1319_ (
  .A({ S25957[918] }),
  .Z({ w[918] })
);
BUF_X1 #() 
BUF_X1_1320_ (
  .A({ S25957[919] }),
  .Z({ w[919] })
);
BUF_X1 #() 
BUF_X1_1321_ (
  .A({ S25957[92] }),
  .Z({ w[92] })
);
BUF_X1 #() 
BUF_X1_1322_ (
  .A({ S25957[920] }),
  .Z({ w[920] })
);
BUF_X1 #() 
BUF_X1_1323_ (
  .A({ S25957[921] }),
  .Z({ w[921] })
);
BUF_X1 #() 
BUF_X1_1324_ (
  .A({ S25957[922] }),
  .Z({ w[922] })
);
BUF_X1 #() 
BUF_X1_1325_ (
  .A({ S25957[923] }),
  .Z({ w[923] })
);
BUF_X1 #() 
BUF_X1_1326_ (
  .A({ S25957[924] }),
  .Z({ w[924] })
);
BUF_X1 #() 
BUF_X1_1327_ (
  .A({ S25957[925] }),
  .Z({ w[925] })
);
BUF_X1 #() 
BUF_X1_1328_ (
  .A({ S25957[926] }),
  .Z({ w[926] })
);
BUF_X1 #() 
BUF_X1_1329_ (
  .A({ S25957[927] }),
  .Z({ w[927] })
);
BUF_X1 #() 
BUF_X1_1330_ (
  .A({ S25957[928] }),
  .Z({ w[928] })
);
BUF_X1 #() 
BUF_X1_1331_ (
  .A({ S25957[929] }),
  .Z({ w[929] })
);
BUF_X1 #() 
BUF_X1_1332_ (
  .A({ S25957[93] }),
  .Z({ w[93] })
);
BUF_X1 #() 
BUF_X1_1333_ (
  .A({ S25957[930] }),
  .Z({ w[930] })
);
BUF_X1 #() 
BUF_X1_1334_ (
  .A({ S25957[931] }),
  .Z({ w[931] })
);
BUF_X1 #() 
BUF_X1_1335_ (
  .A({ S25957[932] }),
  .Z({ w[932] })
);
BUF_X1 #() 
BUF_X1_1336_ (
  .A({ S25957[933] }),
  .Z({ w[933] })
);
BUF_X1 #() 
BUF_X1_1337_ (
  .A({ S25957[934] }),
  .Z({ w[934] })
);
BUF_X1 #() 
BUF_X1_1338_ (
  .A({ S25957[935] }),
  .Z({ w[935] })
);
BUF_X1 #() 
BUF_X1_1339_ (
  .A({ S25957[936] }),
  .Z({ w[936] })
);
BUF_X1 #() 
BUF_X1_1340_ (
  .A({ S25957[937] }),
  .Z({ w[937] })
);
BUF_X1 #() 
BUF_X1_1341_ (
  .A({ S25957[938] }),
  .Z({ w[938] })
);
BUF_X1 #() 
BUF_X1_1342_ (
  .A({ S25957[939] }),
  .Z({ w[939] })
);
BUF_X1 #() 
BUF_X1_1343_ (
  .A({ S25957[94] }),
  .Z({ w[94] })
);
BUF_X1 #() 
BUF_X1_1344_ (
  .A({ S25957[940] }),
  .Z({ w[940] })
);
BUF_X1 #() 
BUF_X1_1345_ (
  .A({ S25957[941] }),
  .Z({ w[941] })
);
BUF_X1 #() 
BUF_X1_1346_ (
  .A({ S25957[942] }),
  .Z({ w[942] })
);
BUF_X1 #() 
BUF_X1_1347_ (
  .A({ S25957[943] }),
  .Z({ w[943] })
);
BUF_X1 #() 
BUF_X1_1348_ (
  .A({ S25957[944] }),
  .Z({ w[944] })
);
BUF_X1 #() 
BUF_X1_1349_ (
  .A({ S25957[945] }),
  .Z({ w[945] })
);
BUF_X1 #() 
BUF_X1_1350_ (
  .A({ S25957[946] }),
  .Z({ w[946] })
);
BUF_X1 #() 
BUF_X1_1351_ (
  .A({ S25957[947] }),
  .Z({ w[947] })
);
BUF_X1 #() 
BUF_X1_1352_ (
  .A({ S25957[948] }),
  .Z({ w[948] })
);
BUF_X1 #() 
BUF_X1_1353_ (
  .A({ S25957[949] }),
  .Z({ w[949] })
);
BUF_X1 #() 
BUF_X1_1354_ (
  .A({ S25957[95] }),
  .Z({ w[95] })
);
BUF_X1 #() 
BUF_X1_1355_ (
  .A({ S25957[950] }),
  .Z({ w[950] })
);
BUF_X1 #() 
BUF_X1_1356_ (
  .A({ S25957[951] }),
  .Z({ w[951] })
);
BUF_X1 #() 
BUF_X1_1357_ (
  .A({ S25957[952] }),
  .Z({ w[952] })
);
BUF_X1 #() 
BUF_X1_1358_ (
  .A({ S25957[953] }),
  .Z({ w[953] })
);
BUF_X1 #() 
BUF_X1_1359_ (
  .A({ S25957[954] }),
  .Z({ w[954] })
);
BUF_X1 #() 
BUF_X1_1360_ (
  .A({ S25957[955] }),
  .Z({ w[955] })
);
BUF_X1 #() 
BUF_X1_1361_ (
  .A({ S25957[956] }),
  .Z({ w[956] })
);
BUF_X1 #() 
BUF_X1_1362_ (
  .A({ S25957[957] }),
  .Z({ w[957] })
);
BUF_X1 #() 
BUF_X1_1363_ (
  .A({ S25957[958] }),
  .Z({ w[958] })
);
BUF_X1 #() 
BUF_X1_1364_ (
  .A({ S25957[959] }),
  .Z({ w[959] })
);
BUF_X1 #() 
BUF_X1_1365_ (
  .A({ S25957[96] }),
  .Z({ w[96] })
);
BUF_X1 #() 
BUF_X1_1366_ (
  .A({ S25957[960] }),
  .Z({ w[960] })
);
BUF_X1 #() 
BUF_X1_1367_ (
  .A({ S25957[961] }),
  .Z({ w[961] })
);
BUF_X1 #() 
BUF_X1_1368_ (
  .A({ S25957[962] }),
  .Z({ w[962] })
);
BUF_X1 #() 
BUF_X1_1369_ (
  .A({ S25957[963] }),
  .Z({ w[963] })
);
BUF_X1 #() 
BUF_X1_1370_ (
  .A({ S25957[964] }),
  .Z({ w[964] })
);
BUF_X1 #() 
BUF_X1_1371_ (
  .A({ S25957[965] }),
  .Z({ w[965] })
);
BUF_X1 #() 
BUF_X1_1372_ (
  .A({ S25957[966] }),
  .Z({ w[966] })
);
BUF_X1 #() 
BUF_X1_1373_ (
  .A({ S25957[967] }),
  .Z({ w[967] })
);
BUF_X1 #() 
BUF_X1_1374_ (
  .A({ S25957[968] }),
  .Z({ w[968] })
);
BUF_X1 #() 
BUF_X1_1375_ (
  .A({ S25957[969] }),
  .Z({ w[969] })
);
BUF_X1 #() 
BUF_X1_1376_ (
  .A({ S25957[97] }),
  .Z({ w[97] })
);
BUF_X1 #() 
BUF_X1_1377_ (
  .A({ S25957[970] }),
  .Z({ w[970] })
);
BUF_X1 #() 
BUF_X1_1378_ (
  .A({ S25957[971] }),
  .Z({ w[971] })
);
BUF_X1 #() 
BUF_X1_1379_ (
  .A({ S25957[972] }),
  .Z({ w[972] })
);
BUF_X1 #() 
BUF_X1_1380_ (
  .A({ S25957[973] }),
  .Z({ w[973] })
);
BUF_X1 #() 
BUF_X1_1381_ (
  .A({ S25957[974] }),
  .Z({ w[974] })
);
BUF_X1 #() 
BUF_X1_1382_ (
  .A({ S25957[975] }),
  .Z({ w[975] })
);
BUF_X1 #() 
BUF_X1_1383_ (
  .A({ S25957[976] }),
  .Z({ w[976] })
);
BUF_X1 #() 
BUF_X1_1384_ (
  .A({ S25957[977] }),
  .Z({ w[977] })
);
BUF_X1 #() 
BUF_X1_1385_ (
  .A({ S25957[978] }),
  .Z({ w[978] })
);
BUF_X1 #() 
BUF_X1_1386_ (
  .A({ S25957[979] }),
  .Z({ w[979] })
);
BUF_X1 #() 
BUF_X1_1387_ (
  .A({ S25957[98] }),
  .Z({ w[98] })
);
BUF_X1 #() 
BUF_X1_1388_ (
  .A({ S25957[980] }),
  .Z({ w[980] })
);
BUF_X1 #() 
BUF_X1_1389_ (
  .A({ S25957[981] }),
  .Z({ w[981] })
);
BUF_X1 #() 
BUF_X1_1390_ (
  .A({ S25957[982] }),
  .Z({ w[982] })
);
BUF_X1 #() 
BUF_X1_1391_ (
  .A({ S25957[983] }),
  .Z({ w[983] })
);
BUF_X1 #() 
BUF_X1_1392_ (
  .A({ S25957[984] }),
  .Z({ w[984] })
);
BUF_X1 #() 
BUF_X1_1393_ (
  .A({ S25957[985] }),
  .Z({ w[985] })
);
BUF_X1 #() 
BUF_X1_1394_ (
  .A({ S25957[986] }),
  .Z({ w[986] })
);
BUF_X1 #() 
BUF_X1_1395_ (
  .A({ S25957[987] }),
  .Z({ w[987] })
);
BUF_X1 #() 
BUF_X1_1396_ (
  .A({ S25957[988] }),
  .Z({ w[988] })
);
BUF_X1 #() 
BUF_X1_1397_ (
  .A({ S25957[989] }),
  .Z({ w[989] })
);
BUF_X1 #() 
BUF_X1_1398_ (
  .A({ S25957[99] }),
  .Z({ w[99] })
);
BUF_X1 #() 
BUF_X1_1399_ (
  .A({ S25957[990] }),
  .Z({ w[990] })
);
BUF_X1 #() 
BUF_X1_1400_ (
  .A({ S25957[991] }),
  .Z({ w[991] })
);
BUF_X1 #() 
BUF_X1_1401_ (
  .A({ S25957[992] }),
  .Z({ w[992] })
);
BUF_X1 #() 
BUF_X1_1402_ (
  .A({ S25957[993] }),
  .Z({ w[993] })
);
BUF_X1 #() 
BUF_X1_1403_ (
  .A({ S25957[994] }),
  .Z({ w[994] })
);
BUF_X1 #() 
BUF_X1_1404_ (
  .A({ S25957[995] }),
  .Z({ w[995] })
);
BUF_X1 #() 
BUF_X1_1405_ (
  .A({ S25957[996] }),
  .Z({ w[996] })
);
BUF_X1 #() 
BUF_X1_1406_ (
  .A({ S25957[997] }),
  .Z({ w[997] })
);
BUF_X1 #() 
BUF_X1_1407_ (
  .A({ S25957[998] }),
  .Z({ w[998] })
);
BUF_X1 #() 
BUF_X1_1408_ (
  .A({ S25957[999] }),
  .Z({ w[999] })
);

endmodule