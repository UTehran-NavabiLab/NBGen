LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

ENTITY TopLevel IS
    PORT (
        clk : IN STD_LOGIC;
        rst : IN STD_LOGIC;
        writeMEM : OUT STD_LOGIC;
        readMEM : OUT STD_LOGIC;
                addrBus : OUT STD_LOGIC_VECTOR (15 DOWNTO 0));
END ENTITY TopLevel;

ARCHITECTURE arch OF TopLevel IS
    SIGNAL S0 : STD_LOGIC;
    SIGNAL S1 : STD_LOGIC;
    SIGNAL S2 : STD_LOGIC;
    SIGNAL S3 : STD_LOGIC;
    SIGNAL S4 : STD_LOGIC;
    SIGNAL S5 : STD_LOGIC;
    SIGNAL S6 : STD_LOGIC;
    SIGNAL S7 : STD_LOGIC;
    SIGNAL S8 : STD_LOGIC;
    SIGNAL S9 : STD_LOGIC;
    SIGNAL S10 : STD_LOGIC;
    SIGNAL S11 : STD_LOGIC;
    SIGNAL S12 : STD_LOGIC;
    SIGNAL S13 : STD_LOGIC;
    SIGNAL S14 : STD_LOGIC;
    SIGNAL S15 : STD_LOGIC;
    SIGNAL S16 : STD_LOGIC;
    SIGNAL S17 : STD_LOGIC;
    SIGNAL S18 : STD_LOGIC;
    SIGNAL S19 : STD_LOGIC;
    SIGNAL S20 : STD_LOGIC;
    SIGNAL S21 : STD_LOGIC;
    SIGNAL S22 : STD_LOGIC;
    SIGNAL S23 : STD_LOGIC;
    SIGNAL S24 : STD_LOGIC;
    SIGNAL S25 : STD_LOGIC;
    SIGNAL S26 : STD_LOGIC;
    SIGNAL S27 : STD_LOGIC;
    SIGNAL S28 : STD_LOGIC;
    SIGNAL S29 : STD_LOGIC;
    SIGNAL S30 : STD_LOGIC;
    SIGNAL S31 : STD_LOGIC;
    SIGNAL S32 : STD_LOGIC;
    SIGNAL S33 : STD_LOGIC;
    SIGNAL S34 : STD_LOGIC;
    SIGNAL S35 : STD_LOGIC;
    SIGNAL S36 : STD_LOGIC;
    SIGNAL S37 : STD_LOGIC;
    SIGNAL S38 : STD_LOGIC;
    SIGNAL S39 : STD_LOGIC;
    SIGNAL S40 : STD_LOGIC;
    SIGNAL S41 : STD_LOGIC;
    SIGNAL S42 : STD_LOGIC;
    SIGNAL S43 : STD_LOGIC;
    SIGNAL S44 : STD_LOGIC;
    SIGNAL S45 : STD_LOGIC;
    SIGNAL S46 : STD_LOGIC;
    SIGNAL S47 : STD_LOGIC;
    SIGNAL S48 : STD_LOGIC;
    SIGNAL S49 : STD_LOGIC;
    SIGNAL S50 : STD_LOGIC;
    SIGNAL S51 : STD_LOGIC;
    SIGNAL S52 : STD_LOGIC;
    SIGNAL S53 : STD_LOGIC;
    SIGNAL S54 : STD_LOGIC;
    SIGNAL S55 : STD_LOGIC;
    SIGNAL S56 : STD_LOGIC;
    SIGNAL S57 : STD_LOGIC;
    SIGNAL S58 : STD_LOGIC;
    SIGNAL S59 : STD_LOGIC;
    SIGNAL S60 : STD_LOGIC;
    SIGNAL S61 : STD_LOGIC;
    SIGNAL S62 : STD_LOGIC;
    SIGNAL S63 : STD_LOGIC;
    SIGNAL S64 : STD_LOGIC;
    SIGNAL S65 : STD_LOGIC;
    SIGNAL S66 : STD_LOGIC;
    SIGNAL S67 : STD_LOGIC;
    SIGNAL S68 : STD_LOGIC;
    SIGNAL S69 : STD_LOGIC;
    SIGNAL S70 : STD_LOGIC;
    SIGNAL S71 : STD_LOGIC;
    SIGNAL S72 : STD_LOGIC;
    SIGNAL S73 : STD_LOGIC;
    SIGNAL S74 : STD_LOGIC;
    SIGNAL S75 : STD_LOGIC;
    SIGNAL S76 : STD_LOGIC;
    SIGNAL S77 : STD_LOGIC;
    SIGNAL S78 : STD_LOGIC;
    SIGNAL S79 : STD_LOGIC;
    SIGNAL S80 : STD_LOGIC;
    SIGNAL S81 : STD_LOGIC;
    SIGNAL S82 : STD_LOGIC;
    SIGNAL S83 : STD_LOGIC;
    SIGNAL S84 : STD_LOGIC;
    SIGNAL S85 : STD_LOGIC;
    SIGNAL S86 : STD_LOGIC;
    SIGNAL S87 : STD_LOGIC;
    SIGNAL S88 : STD_LOGIC;
    SIGNAL S89 : STD_LOGIC;
    SIGNAL S90 : STD_LOGIC;
    SIGNAL S91 : STD_LOGIC;
    SIGNAL S92 : STD_LOGIC;
    SIGNAL S93 : STD_LOGIC;
    SIGNAL S94 : STD_LOGIC;
    SIGNAL S95 : STD_LOGIC;
    SIGNAL S96 : STD_LOGIC;
    SIGNAL S97 : STD_LOGIC;
    SIGNAL S98 : STD_LOGIC;
    SIGNAL S99 : STD_LOGIC;
    SIGNAL S100 : STD_LOGIC;
    SIGNAL S101 : STD_LOGIC;
    SIGNAL S102 : STD_LOGIC;
    SIGNAL S103 : STD_LOGIC;
    SIGNAL S104 : STD_LOGIC;
    SIGNAL S105 : STD_LOGIC;
    SIGNAL S106 : STD_LOGIC;
    SIGNAL S107 : STD_LOGIC;
    SIGNAL S108 : STD_LOGIC;
    SIGNAL S109 : STD_LOGIC;
    SIGNAL S110 : STD_LOGIC;
    SIGNAL S111 : STD_LOGIC;
    SIGNAL S112 : STD_LOGIC;
    SIGNAL S113 : STD_LOGIC;
    SIGNAL S114 : STD_LOGIC;
    SIGNAL S115 : STD_LOGIC;
    SIGNAL S116 : STD_LOGIC;
    SIGNAL S117 : STD_LOGIC;
    SIGNAL S118 : STD_LOGIC;
    SIGNAL S119 : STD_LOGIC;
    SIGNAL S120 : STD_LOGIC;
    SIGNAL S121 : STD_LOGIC;
    SIGNAL S122 : STD_LOGIC;
    SIGNAL S123 : STD_LOGIC;
    SIGNAL S124 : STD_LOGIC;
    SIGNAL S125 : STD_LOGIC;
    SIGNAL S126 : STD_LOGIC;
    SIGNAL S127 : STD_LOGIC;
    SIGNAL S128 : STD_LOGIC;
    SIGNAL S129 : STD_LOGIC;
    SIGNAL S130 : STD_LOGIC;
    SIGNAL S131 : STD_LOGIC;
    SIGNAL S132 : STD_LOGIC;
    SIGNAL S133 : STD_LOGIC;
    SIGNAL S134 : STD_LOGIC;
    SIGNAL S135 : STD_LOGIC;
    SIGNAL S136 : STD_LOGIC;
    SIGNAL S137 : STD_LOGIC;
    SIGNAL S138 : STD_LOGIC;
    SIGNAL S139 : STD_LOGIC;
    SIGNAL S140 : STD_LOGIC;
    SIGNAL S141 : STD_LOGIC;
    SIGNAL S142 : STD_LOGIC;
    SIGNAL S143 : STD_LOGIC;
    SIGNAL S144 : STD_LOGIC;
    SIGNAL S145 : STD_LOGIC;
    SIGNAL S146 : STD_LOGIC;
    SIGNAL S147 : STD_LOGIC;
    SIGNAL S148 : STD_LOGIC;
    SIGNAL S149 : STD_LOGIC;
    SIGNAL S150 : STD_LOGIC;
    SIGNAL S151 : STD_LOGIC;
    SIGNAL S152 : STD_LOGIC;
    SIGNAL S153 : STD_LOGIC;
    SIGNAL S154 : STD_LOGIC;
    SIGNAL S155 : STD_LOGIC;
    SIGNAL S156 : STD_LOGIC;
    SIGNAL S157 : STD_LOGIC;
    SIGNAL S158 : STD_LOGIC;
    SIGNAL S159 : STD_LOGIC;
    SIGNAL S160 : STD_LOGIC;
    SIGNAL S161 : STD_LOGIC;
    SIGNAL S162 : STD_LOGIC;
    SIGNAL S163 : STD_LOGIC;
    SIGNAL S164 : STD_LOGIC;
    SIGNAL S165 : STD_LOGIC;
    SIGNAL S166 : STD_LOGIC;
    SIGNAL S167 : STD_LOGIC;
    SIGNAL S168 : STD_LOGIC;
    SIGNAL S169 : STD_LOGIC;
    SIGNAL S170 : STD_LOGIC;
    SIGNAL S171 : STD_LOGIC;
    SIGNAL S172 : STD_LOGIC;
    SIGNAL S173 : STD_LOGIC;
    SIGNAL S174 : STD_LOGIC;
    SIGNAL S175 : STD_LOGIC;
    SIGNAL S176 : STD_LOGIC;
    SIGNAL S177 : STD_LOGIC;
    SIGNAL S178 : STD_LOGIC;
    SIGNAL S179 : STD_LOGIC;
    SIGNAL S180 : STD_LOGIC;
    SIGNAL S181 : STD_LOGIC;
    SIGNAL S182 : STD_LOGIC;
    SIGNAL S183 : STD_LOGIC;
    SIGNAL S184 : STD_LOGIC;
    SIGNAL S185 : STD_LOGIC;
    SIGNAL S186 : STD_LOGIC;
    SIGNAL S187 : STD_LOGIC;
    SIGNAL S188 : STD_LOGIC;
    SIGNAL S189 : STD_LOGIC;
    SIGNAL S190 : STD_LOGIC;
    SIGNAL S191 : STD_LOGIC;
    SIGNAL S192 : STD_LOGIC;
    SIGNAL S193 : STD_LOGIC;
    SIGNAL S194 : STD_LOGIC;
    SIGNAL S195 : STD_LOGIC;
    SIGNAL S196 : STD_LOGIC;
    SIGNAL S197 : STD_LOGIC;
    SIGNAL S198 : STD_LOGIC;
    SIGNAL S199 : STD_LOGIC;
    SIGNAL S200 : STD_LOGIC;
    SIGNAL S201 : STD_LOGIC;
    SIGNAL S202 : STD_LOGIC;
    SIGNAL S203 : STD_LOGIC;
    SIGNAL S204 : STD_LOGIC;
    SIGNAL S205 : STD_LOGIC;
    SIGNAL S206 : STD_LOGIC;
    SIGNAL S207 : STD_LOGIC;
    SIGNAL S208 : STD_LOGIC;
    SIGNAL S209 : STD_LOGIC;
    SIGNAL S210 : STD_LOGIC;
    SIGNAL S211 : STD_LOGIC;
    SIGNAL S212 : STD_LOGIC;
    SIGNAL S213 : STD_LOGIC;
    SIGNAL S214 : STD_LOGIC;
    SIGNAL S215 : STD_LOGIC;
    SIGNAL S216 : STD_LOGIC;
    SIGNAL S217 : STD_LOGIC;
    SIGNAL S218 : STD_LOGIC;
    SIGNAL S219 : STD_LOGIC;
    SIGNAL S220 : STD_LOGIC;
    SIGNAL S221 : STD_LOGIC;
    SIGNAL S222 : STD_LOGIC;
    SIGNAL S223 : STD_LOGIC;
    SIGNAL S224 : STD_LOGIC;
    SIGNAL S225 : STD_LOGIC;
    SIGNAL S226 : STD_LOGIC;
    SIGNAL S227 : STD_LOGIC;
    SIGNAL S228 : STD_LOGIC;
    SIGNAL S229 : STD_LOGIC;
    SIGNAL S230 : STD_LOGIC;
    SIGNAL S231 : STD_LOGIC;
    SIGNAL S232 : STD_LOGIC;
    SIGNAL S233 : STD_LOGIC;
    SIGNAL S234 : STD_LOGIC;
    SIGNAL S235 : STD_LOGIC;
    SIGNAL S236 : STD_LOGIC;
    SIGNAL S237 : STD_LOGIC;
    SIGNAL S238 : STD_LOGIC;
    SIGNAL S239 : STD_LOGIC;
    SIGNAL S240 : STD_LOGIC;
    SIGNAL S241 : STD_LOGIC;
    SIGNAL S242 : STD_LOGIC;
    SIGNAL S243 : STD_LOGIC;
    SIGNAL S244 : STD_LOGIC;
    SIGNAL S245 : STD_LOGIC;
    SIGNAL S246 : STD_LOGIC;
    SIGNAL S247 : STD_LOGIC;
    SIGNAL S248 : STD_LOGIC;
    SIGNAL S249 : STD_LOGIC;
    SIGNAL S250 : STD_LOGIC;
    SIGNAL S251 : STD_LOGIC;
    SIGNAL S252 : STD_LOGIC;
    SIGNAL S253 : STD_LOGIC;
    SIGNAL S254 : STD_LOGIC;
    SIGNAL S255 : STD_LOGIC;
    SIGNAL S256 : STD_LOGIC;
    SIGNAL S257 : STD_LOGIC;
    SIGNAL S258 : STD_LOGIC;
    SIGNAL S259 : STD_LOGIC;
    SIGNAL S260 : STD_LOGIC;
    SIGNAL S261 : STD_LOGIC;
    SIGNAL S262 : STD_LOGIC;
    SIGNAL S263 : STD_LOGIC;
    SIGNAL S264 : STD_LOGIC;
    SIGNAL S265 : STD_LOGIC;
    SIGNAL S266 : STD_LOGIC;
    SIGNAL S267 : STD_LOGIC;
    SIGNAL S268 : STD_LOGIC;
    SIGNAL S269 : STD_LOGIC;
    SIGNAL S270 : STD_LOGIC;
    SIGNAL S271 : STD_LOGIC;
    SIGNAL S272 : STD_LOGIC;
    SIGNAL S273 : STD_LOGIC;
    SIGNAL S274 : STD_LOGIC;
    SIGNAL S275 : STD_LOGIC;
    SIGNAL S276 : STD_LOGIC;
    SIGNAL S277 : STD_LOGIC;
    SIGNAL S278 : STD_LOGIC;
    SIGNAL S279 : STD_LOGIC;
    SIGNAL S280 : STD_LOGIC;
    SIGNAL S281 : STD_LOGIC;
    SIGNAL S282 : STD_LOGIC;
    SIGNAL S283 : STD_LOGIC;
    SIGNAL S284 : STD_LOGIC;
    SIGNAL S285 : STD_LOGIC;
    SIGNAL S286 : STD_LOGIC;
    SIGNAL S287 : STD_LOGIC;
    SIGNAL S288 : STD_LOGIC;
    SIGNAL S289 : STD_LOGIC;
    SIGNAL S290 : STD_LOGIC;
    SIGNAL S291 : STD_LOGIC;
    SIGNAL S292 : STD_LOGIC;
    SIGNAL S293 : STD_LOGIC;
    SIGNAL S294 : STD_LOGIC;
    SIGNAL S295 : STD_LOGIC;
    SIGNAL S296 : STD_LOGIC;
    SIGNAL S297 : STD_LOGIC;
    SIGNAL S298 : STD_LOGIC;
    SIGNAL S299 : STD_LOGIC;
    SIGNAL S300 : STD_LOGIC;
    SIGNAL S301 : STD_LOGIC;
    SIGNAL S302 : STD_LOGIC;
    SIGNAL S303 : STD_LOGIC;
    SIGNAL S304 : STD_LOGIC;
    SIGNAL S305 : STD_LOGIC;
    SIGNAL S306 : STD_LOGIC;
    SIGNAL S307 : STD_LOGIC;
    SIGNAL S308 : STD_LOGIC;
    SIGNAL S309 : STD_LOGIC;
    SIGNAL S310 : STD_LOGIC;
    SIGNAL S311 : STD_LOGIC;
    SIGNAL S312 : STD_LOGIC;
    SIGNAL S313 : STD_LOGIC;
    SIGNAL S314 : STD_LOGIC;
    SIGNAL S315 : STD_LOGIC;
    SIGNAL S316 : STD_LOGIC;
    SIGNAL S317 : STD_LOGIC;
    SIGNAL S318 : STD_LOGIC;
    SIGNAL S319 : STD_LOGIC;
    SIGNAL S320 : STD_LOGIC;
    SIGNAL S321 : STD_LOGIC;
    SIGNAL S322 : STD_LOGIC;
    SIGNAL S323 : STD_LOGIC;
    SIGNAL S324 : STD_LOGIC;
    SIGNAL S325 : STD_LOGIC;
    SIGNAL S326 : STD_LOGIC;
    SIGNAL S327 : STD_LOGIC;
    SIGNAL S328 : STD_LOGIC;
    SIGNAL S329 : STD_LOGIC;
    SIGNAL S330 : STD_LOGIC;
    SIGNAL S331 : STD_LOGIC;
    SIGNAL S332 : STD_LOGIC;
    SIGNAL S333 : STD_LOGIC;
    SIGNAL S334 : STD_LOGIC;
    SIGNAL S335 : STD_LOGIC;
    SIGNAL S336 : STD_LOGIC;
    SIGNAL S337 : STD_LOGIC;
    SIGNAL S338 : STD_LOGIC;
    SIGNAL S339 : STD_LOGIC;
    SIGNAL S340 : STD_LOGIC;
    SIGNAL S341 : STD_LOGIC;
    SIGNAL S342 : STD_LOGIC;
    SIGNAL S343 : STD_LOGIC;
    SIGNAL S344 : STD_LOGIC;
    SIGNAL S345 : STD_LOGIC;
    SIGNAL S346 : STD_LOGIC;
    SIGNAL S347 : STD_LOGIC;
    SIGNAL S348 : STD_LOGIC;
    SIGNAL S349 : STD_LOGIC;
    SIGNAL S350 : STD_LOGIC;
    SIGNAL S351 : STD_LOGIC;
    SIGNAL S352 : STD_LOGIC;
    SIGNAL S353 : STD_LOGIC;
    SIGNAL S354 : STD_LOGIC;
    SIGNAL S355 : STD_LOGIC;
    SIGNAL S356 : STD_LOGIC;
    SIGNAL S357 : STD_LOGIC;
    SIGNAL S358 : STD_LOGIC;
    SIGNAL S359 : STD_LOGIC;
    SIGNAL S360 : STD_LOGIC;
    SIGNAL S361 : STD_LOGIC;
    SIGNAL S362 : STD_LOGIC;
    SIGNAL S363 : STD_LOGIC;
    SIGNAL S364 : STD_LOGIC;
    SIGNAL S365 : STD_LOGIC;
    SIGNAL S366 : STD_LOGIC;
    SIGNAL S367 : STD_LOGIC;
    SIGNAL S368 : STD_LOGIC;
    SIGNAL S369 : STD_LOGIC;
    SIGNAL S370 : STD_LOGIC;
    SIGNAL S371 : STD_LOGIC;
    SIGNAL S372 : STD_LOGIC;
    SIGNAL S373 : STD_LOGIC;
    SIGNAL S374 : STD_LOGIC;
    SIGNAL S375 : STD_LOGIC;
    SIGNAL S376 : STD_LOGIC;
    SIGNAL S377 : STD_LOGIC;
    SIGNAL S378 : STD_LOGIC;
    SIGNAL S379 : STD_LOGIC;
    SIGNAL S380 : STD_LOGIC;
    SIGNAL S381 : STD_LOGIC;
    SIGNAL S382 : STD_LOGIC;
    SIGNAL S383 : STD_LOGIC;
    SIGNAL S384 : STD_LOGIC;
    SIGNAL S385 : STD_LOGIC;
    SIGNAL S386 : STD_LOGIC;
    SIGNAL S387 : STD_LOGIC;
    SIGNAL S388 : STD_LOGIC;
    SIGNAL S389 : STD_LOGIC;
    SIGNAL S390 : STD_LOGIC;
    SIGNAL S391 : STD_LOGIC;
    SIGNAL S392 : STD_LOGIC;
    SIGNAL S393 : STD_LOGIC;
    SIGNAL S394 : STD_LOGIC;
    SIGNAL S395 : STD_LOGIC;
    SIGNAL S396 : STD_LOGIC;
    SIGNAL S397 : STD_LOGIC;
    SIGNAL S398 : STD_LOGIC;
    SIGNAL S399 : STD_LOGIC;
    SIGNAL S400 : STD_LOGIC;
    SIGNAL S401 : STD_LOGIC;
    SIGNAL S402 : STD_LOGIC;
    SIGNAL S403 : STD_LOGIC;
    SIGNAL S404 : STD_LOGIC;
    SIGNAL S405 : STD_LOGIC;
    SIGNAL S406 : STD_LOGIC;
    SIGNAL S407 : STD_LOGIC;
    SIGNAL S408 : STD_LOGIC;
    SIGNAL S409 : STD_LOGIC;
    SIGNAL S410 : STD_LOGIC;
    SIGNAL S411 : STD_LOGIC;
    SIGNAL S412 : STD_LOGIC;
    SIGNAL S413 : STD_LOGIC;
    SIGNAL S414 : STD_LOGIC;
    SIGNAL S415 : STD_LOGIC;
    SIGNAL S416 : STD_LOGIC;
    SIGNAL S417 : STD_LOGIC;
    SIGNAL S418 : STD_LOGIC;
    SIGNAL S419 : STD_LOGIC;
    SIGNAL S420 : STD_LOGIC;
    SIGNAL S421 : STD_LOGIC;
    SIGNAL S422 : STD_LOGIC;
    SIGNAL S423 : STD_LOGIC;
    SIGNAL S424 : STD_LOGIC;
    SIGNAL S425 : STD_LOGIC;
    SIGNAL S426 : STD_LOGIC;
    SIGNAL S427 : STD_LOGIC;
    SIGNAL S428 : STD_LOGIC;
    SIGNAL S429 : STD_LOGIC;
    SIGNAL S430 : STD_LOGIC;
    SIGNAL S431 : STD_LOGIC;
    SIGNAL S432 : STD_LOGIC;
    SIGNAL S433 : STD_LOGIC;
    SIGNAL S434 : STD_LOGIC;
    SIGNAL S435 : STD_LOGIC;
    SIGNAL S436 : STD_LOGIC;
    SIGNAL S437 : STD_LOGIC;
    SIGNAL S438 : STD_LOGIC;
    SIGNAL S439 : STD_LOGIC;
    SIGNAL S440 : STD_LOGIC;
    SIGNAL S441 : STD_LOGIC;
    SIGNAL S442 : STD_LOGIC;
    SIGNAL S443 : STD_LOGIC;
    SIGNAL S444 : STD_LOGIC;
    SIGNAL S445 : STD_LOGIC;
    SIGNAL S446 : STD_LOGIC;
    SIGNAL S447 : STD_LOGIC;
    SIGNAL S448 : STD_LOGIC;
    SIGNAL S449 : STD_LOGIC;
    SIGNAL S450 : STD_LOGIC;
    SIGNAL S451 : STD_LOGIC;
    SIGNAL S452 : STD_LOGIC;
    SIGNAL S453 : STD_LOGIC;
    SIGNAL S454 : STD_LOGIC;
    SIGNAL S455 : STD_LOGIC;
    SIGNAL S456 : STD_LOGIC;
    SIGNAL S457 : STD_LOGIC;
    SIGNAL S458 : STD_LOGIC;
    SIGNAL S459 : STD_LOGIC;
    SIGNAL S460 : STD_LOGIC;
    SIGNAL S461 : STD_LOGIC;
    SIGNAL S462 : STD_LOGIC;
    SIGNAL S463 : STD_LOGIC;
    SIGNAL S464 : STD_LOGIC;
    SIGNAL S465 : STD_LOGIC;
    SIGNAL S466 : STD_LOGIC;
    SIGNAL S467 : STD_LOGIC;
    SIGNAL S468 : STD_LOGIC;
    SIGNAL S469 : STD_LOGIC;
    SIGNAL S470 : STD_LOGIC;
    SIGNAL S471 : STD_LOGIC;
    SIGNAL S472 : STD_LOGIC;
    SIGNAL S473 : STD_LOGIC;
    SIGNAL S474 : STD_LOGIC;
    SIGNAL S475 : STD_LOGIC;
    SIGNAL S476 : STD_LOGIC;
    SIGNAL S477 : STD_LOGIC;
    SIGNAL S478 : STD_LOGIC;
    SIGNAL S479 : STD_LOGIC;
    SIGNAL S480 : STD_LOGIC;
    SIGNAL S481 : STD_LOGIC;
    SIGNAL S482 : STD_LOGIC;
    SIGNAL S483 : STD_LOGIC;
    SIGNAL S484 : STD_LOGIC;
    SIGNAL S485 : STD_LOGIC;
    SIGNAL S486 : STD_LOGIC;
    SIGNAL S487 : STD_LOGIC;
    SIGNAL S488 : STD_LOGIC;
    SIGNAL S489 : STD_LOGIC;
    SIGNAL S490 : STD_LOGIC;
    SIGNAL S491 : STD_LOGIC;
    SIGNAL S492 : STD_LOGIC;
    SIGNAL S493 : STD_LOGIC;
    SIGNAL S494 : STD_LOGIC;
    SIGNAL S495 : STD_LOGIC;
    SIGNAL S496 : STD_LOGIC;
    SIGNAL S497 : STD_LOGIC;
    SIGNAL S498 : STD_LOGIC;
    SIGNAL S499 : STD_LOGIC;
    SIGNAL S500 : STD_LOGIC;
    SIGNAL S501 : STD_LOGIC;
    SIGNAL S502 : STD_LOGIC;
    SIGNAL S503 : STD_LOGIC;
    SIGNAL S504 : STD_LOGIC;
    SIGNAL S505 : STD_LOGIC;
    SIGNAL S506 : STD_LOGIC;
    SIGNAL S507 : STD_LOGIC;
    SIGNAL S508 : STD_LOGIC;
    SIGNAL S509 : STD_LOGIC;
    SIGNAL S510 : STD_LOGIC;
    SIGNAL S511 : STD_LOGIC;
    SIGNAL S512 : STD_LOGIC;
    SIGNAL S513 : STD_LOGIC;
    SIGNAL S514 : STD_LOGIC;
    SIGNAL S515 : STD_LOGIC;
    SIGNAL S516 : STD_LOGIC;
    SIGNAL S517 : STD_LOGIC;
    SIGNAL S518 : STD_LOGIC;
    SIGNAL S519 : STD_LOGIC;
    SIGNAL S520 : STD_LOGIC;
    SIGNAL S521 : STD_LOGIC;
    SIGNAL S522 : STD_LOGIC;
    SIGNAL S523 : STD_LOGIC;
    SIGNAL S524 : STD_LOGIC;
    SIGNAL S525 : STD_LOGIC;
    SIGNAL S526 : STD_LOGIC;
    SIGNAL S527 : STD_LOGIC;
    SIGNAL S528 : STD_LOGIC;
    SIGNAL S529 : STD_LOGIC;
    SIGNAL S530 : STD_LOGIC;
    SIGNAL S531 : STD_LOGIC;
    SIGNAL S532 : STD_LOGIC;
    SIGNAL S533 : STD_LOGIC;
    SIGNAL S534 : STD_LOGIC;
    SIGNAL S535 : STD_LOGIC;
    SIGNAL S536 : STD_LOGIC;
    SIGNAL S537 : STD_LOGIC;
    SIGNAL S538 : STD_LOGIC;
    SIGNAL S539 : STD_LOGIC;
    SIGNAL S540 : STD_LOGIC;
    SIGNAL S541 : STD_LOGIC;
    SIGNAL S542 : STD_LOGIC;
    SIGNAL S543 : STD_LOGIC;
    SIGNAL S544 : STD_LOGIC;
    SIGNAL S545 : STD_LOGIC;
    SIGNAL S546 : STD_LOGIC;
    SIGNAL S547 : STD_LOGIC;
    SIGNAL S548 : STD_LOGIC;
    SIGNAL S549 : STD_LOGIC;
    SIGNAL S550 : STD_LOGIC;
    SIGNAL S551 : STD_LOGIC;
    SIGNAL S552 : STD_LOGIC;
    SIGNAL S553 : STD_LOGIC;
    SIGNAL S554 : STD_LOGIC;
    SIGNAL S555 : STD_LOGIC;
    SIGNAL S556 : STD_LOGIC;
    SIGNAL S557 : STD_LOGIC;
    SIGNAL S558 : STD_LOGIC;
    SIGNAL S559 : STD_LOGIC;
    SIGNAL S560 : STD_LOGIC;
    SIGNAL S561 : STD_LOGIC;
    SIGNAL S562 : STD_LOGIC;
    SIGNAL S563 : STD_LOGIC;
    SIGNAL S564 : STD_LOGIC;
    SIGNAL S565 : STD_LOGIC;
    SIGNAL S566 : STD_LOGIC;
    SIGNAL S567 : STD_LOGIC;
    SIGNAL S568 : STD_LOGIC;
    SIGNAL S569 : STD_LOGIC;
    SIGNAL S570 : STD_LOGIC;
    SIGNAL S571 : STD_LOGIC;
    SIGNAL S572 : STD_LOGIC;
    SIGNAL S573 : STD_LOGIC;
    SIGNAL S574 : STD_LOGIC;
    SIGNAL S575 : STD_LOGIC;
    SIGNAL S576 : STD_LOGIC;
    SIGNAL S577 : STD_LOGIC;
    SIGNAL S578 : STD_LOGIC;
    SIGNAL S579 : STD_LOGIC;
    SIGNAL S580 : STD_LOGIC;
    SIGNAL S581 : STD_LOGIC;
    SIGNAL S582 : STD_LOGIC;
    SIGNAL S583 : STD_LOGIC;
    SIGNAL S584 : STD_LOGIC;
    SIGNAL S585 : STD_LOGIC;
    SIGNAL S586 : STD_LOGIC;
    SIGNAL S587 : STD_LOGIC;
    SIGNAL S588 : STD_LOGIC;
    SIGNAL S589 : STD_LOGIC;
    SIGNAL S590 : STD_LOGIC;
    SIGNAL S591 : STD_LOGIC;
    SIGNAL S592 : STD_LOGIC;
    SIGNAL S593 : STD_LOGIC;
    SIGNAL S594 : STD_LOGIC;
    SIGNAL S595 : STD_LOGIC;
    SIGNAL S596 : STD_LOGIC;
    SIGNAL S597 : STD_LOGIC;
    SIGNAL S598 : STD_LOGIC;
    SIGNAL S599 : STD_LOGIC;
    SIGNAL S600 : STD_LOGIC;
    SIGNAL S601 : STD_LOGIC;
    SIGNAL S602 : STD_LOGIC;
    SIGNAL S603 : STD_LOGIC;
    SIGNAL S604 : STD_LOGIC;
    SIGNAL S605 : STD_LOGIC;
    SIGNAL S606 : STD_LOGIC;
    SIGNAL S607 : STD_LOGIC;
    SIGNAL S608 : STD_LOGIC;
    SIGNAL S609 : STD_LOGIC;
    SIGNAL S610 : STD_LOGIC;
    SIGNAL S611 : STD_LOGIC;
    SIGNAL S612 : STD_LOGIC;
    SIGNAL S613 : STD_LOGIC;
    SIGNAL S614 : STD_LOGIC;
    SIGNAL S615 : STD_LOGIC;
    SIGNAL S616 : STD_LOGIC;
    SIGNAL S617 : STD_LOGIC;
    SIGNAL S618 : STD_LOGIC;
    SIGNAL S619 : STD_LOGIC;
    SIGNAL S620 : STD_LOGIC;
    SIGNAL S621 : STD_LOGIC;
    SIGNAL S622 : STD_LOGIC;
    SIGNAL S623 : STD_LOGIC;
    SIGNAL S624 : STD_LOGIC;
    SIGNAL S625 : STD_LOGIC;
    SIGNAL S626 : STD_LOGIC;
    SIGNAL S627 : STD_LOGIC;
    SIGNAL S628 : STD_LOGIC;
    SIGNAL S629 : STD_LOGIC;
    SIGNAL S630 : STD_LOGIC;
    SIGNAL S631 : STD_LOGIC;
    SIGNAL S632 : STD_LOGIC;
    SIGNAL S633 : STD_LOGIC;
    SIGNAL S634 : STD_LOGIC;
    SIGNAL S635 : STD_LOGIC;
    SIGNAL S636 : STD_LOGIC;
    SIGNAL S637 : STD_LOGIC;
    SIGNAL S638 : STD_LOGIC;
    SIGNAL S639 : STD_LOGIC;
    SIGNAL S640 : STD_LOGIC;
    SIGNAL S641 : STD_LOGIC;
    SIGNAL S642 : STD_LOGIC;
    SIGNAL S643 : STD_LOGIC;
    SIGNAL S644 : STD_LOGIC;
    SIGNAL S645 : STD_LOGIC;
    SIGNAL S646 : STD_LOGIC;
    SIGNAL S647 : STD_LOGIC;
    SIGNAL S648 : STD_LOGIC;
    SIGNAL S649 : STD_LOGIC;
    SIGNAL S650 : STD_LOGIC;
    SIGNAL S651 : STD_LOGIC;
    SIGNAL S652 : STD_LOGIC;
    SIGNAL S653 : STD_LOGIC;
    SIGNAL S654 : STD_LOGIC;
    SIGNAL S655 : STD_LOGIC;
    SIGNAL S656 : STD_LOGIC;
    SIGNAL S657 : STD_LOGIC;
    SIGNAL S658 : STD_LOGIC;
    SIGNAL S659 : STD_LOGIC;
    SIGNAL S660 : STD_LOGIC;
    SIGNAL S661 : STD_LOGIC;
    SIGNAL S662 : STD_LOGIC;
    SIGNAL S663 : STD_LOGIC;
    SIGNAL S664 : STD_LOGIC;
    SIGNAL S665 : STD_LOGIC;
    SIGNAL S666 : STD_LOGIC;
    SIGNAL S667 : STD_LOGIC;
    SIGNAL S668 : STD_LOGIC;
    SIGNAL S669 : STD_LOGIC;
    SIGNAL S670 : STD_LOGIC;
    SIGNAL S671 : STD_LOGIC;
    SIGNAL S672 : STD_LOGIC;
    SIGNAL S673 : STD_LOGIC;
    SIGNAL S674 : STD_LOGIC;
    SIGNAL S675 : STD_LOGIC;
    SIGNAL S676 : STD_LOGIC;
    SIGNAL S677 : STD_LOGIC;
    SIGNAL S678 : STD_LOGIC;
    SIGNAL S679 : STD_LOGIC;
    SIGNAL S680 : STD_LOGIC;
    SIGNAL S681 : STD_LOGIC;
    SIGNAL S682 : STD_LOGIC;
    SIGNAL S683 : STD_LOGIC;
    SIGNAL S684 : STD_LOGIC;
    SIGNAL S685 : STD_LOGIC;
    SIGNAL S686 : STD_LOGIC;
    SIGNAL S687 : STD_LOGIC;
    SIGNAL S688 : STD_LOGIC;
    SIGNAL S689 : STD_LOGIC;
    SIGNAL S690 : STD_LOGIC;
    SIGNAL S691 : STD_LOGIC;
    SIGNAL S692 : STD_LOGIC;
    SIGNAL S693 : STD_LOGIC;
    SIGNAL S694 : STD_LOGIC;
    SIGNAL S695 : STD_LOGIC;
    SIGNAL S696 : STD_LOGIC;
    SIGNAL S697 : STD_LOGIC;
    SIGNAL S698 : STD_LOGIC;
    SIGNAL S699 : STD_LOGIC;
    SIGNAL S700 : STD_LOGIC;
    SIGNAL S701 : STD_LOGIC;
    SIGNAL S702 : STD_LOGIC;
    SIGNAL S703 : STD_LOGIC;
    SIGNAL S704 : STD_LOGIC;
    SIGNAL S705 : STD_LOGIC;
    SIGNAL S706 : STD_LOGIC;
    SIGNAL S707 : STD_LOGIC;
    SIGNAL S708 : STD_LOGIC;
    SIGNAL S709 : STD_LOGIC;
    SIGNAL S710 : STD_LOGIC;
    SIGNAL S711 : STD_LOGIC;
    SIGNAL S712 : STD_LOGIC;
    SIGNAL S713 : STD_LOGIC;
    SIGNAL S714 : STD_LOGIC;
    SIGNAL S715 : STD_LOGIC;
    SIGNAL S716 : STD_LOGIC;
    SIGNAL S717 : STD_LOGIC;
    SIGNAL S718 : STD_LOGIC;
    SIGNAL S719 : STD_LOGIC;
    SIGNAL S720 : STD_LOGIC;
    SIGNAL S721 : STD_LOGIC;
    SIGNAL S722 : STD_LOGIC;
    SIGNAL S723 : STD_LOGIC;
    SIGNAL S724 : STD_LOGIC;
    SIGNAL S725 : STD_LOGIC;
    SIGNAL S726 : STD_LOGIC;
    SIGNAL S727 : STD_LOGIC;
    SIGNAL S728 : STD_LOGIC;
    SIGNAL S729 : STD_LOGIC;
    SIGNAL S730 : STD_LOGIC;
    SIGNAL S731 : STD_LOGIC;
    SIGNAL S732 : STD_LOGIC;
    SIGNAL S733 : STD_LOGIC;
    SIGNAL S734 : STD_LOGIC;
    SIGNAL S735 : STD_LOGIC;
    SIGNAL S736 : STD_LOGIC;
    SIGNAL S737 : STD_LOGIC;
    SIGNAL S738 : STD_LOGIC;
    SIGNAL S739 : STD_LOGIC;
    SIGNAL S740 : STD_LOGIC;
    SIGNAL S741 : STD_LOGIC;
    SIGNAL S742 : STD_LOGIC;
    SIGNAL S743 : STD_LOGIC;
    SIGNAL S744 : STD_LOGIC;
    SIGNAL S745 : STD_LOGIC;
    SIGNAL S746 : STD_LOGIC;
    SIGNAL S747 : STD_LOGIC;
    SIGNAL S748 : STD_LOGIC;
    SIGNAL S749 : STD_LOGIC;
    SIGNAL S750 : STD_LOGIC;
    SIGNAL S751 : STD_LOGIC;
    SIGNAL S752 : STD_LOGIC;
    SIGNAL S753 : STD_LOGIC;
    SIGNAL S754 : STD_LOGIC;
    SIGNAL S755 : STD_LOGIC;
    SIGNAL S756 : STD_LOGIC;
    SIGNAL S757 : STD_LOGIC;
    SIGNAL S758 : STD_LOGIC;
    SIGNAL S759 : STD_LOGIC;
    SIGNAL S760 : STD_LOGIC;
    SIGNAL S761 : STD_LOGIC;
    SIGNAL S762 : STD_LOGIC;
    SIGNAL S763 : STD_LOGIC;
    SIGNAL S764 : STD_LOGIC;
    SIGNAL S765 : STD_LOGIC;
    SIGNAL S766 : STD_LOGIC;
    SIGNAL S767 : STD_LOGIC;
    SIGNAL S768 : STD_LOGIC;
    SIGNAL S769 : STD_LOGIC;
    SIGNAL S770 : STD_LOGIC;
    SIGNAL S771 : STD_LOGIC;
    SIGNAL S772 : STD_LOGIC;
    SIGNAL S773 : STD_LOGIC;
    SIGNAL S774 : STD_LOGIC;
    SIGNAL S775 : STD_LOGIC;
    SIGNAL S776 : STD_LOGIC;
    SIGNAL S777 : STD_LOGIC;
    SIGNAL S778 : STD_LOGIC;
    SIGNAL S779 : STD_LOGIC;
    SIGNAL S780 : STD_LOGIC;
    SIGNAL S781 : STD_LOGIC;
    SIGNAL S782 : STD_LOGIC;
    SIGNAL S783 : STD_LOGIC;
    SIGNAL S784 : STD_LOGIC;
    SIGNAL S785 : STD_LOGIC;
    SIGNAL S786 : STD_LOGIC;
    SIGNAL S787 : STD_LOGIC;
    SIGNAL S788 : STD_LOGIC;
    SIGNAL S789 : STD_LOGIC;
    SIGNAL S790 : STD_LOGIC;
    SIGNAL S791 : STD_LOGIC;
    SIGNAL S792 : STD_LOGIC;
    SIGNAL S793 : STD_LOGIC;
    SIGNAL S794 : STD_LOGIC;
    SIGNAL S795 : STD_LOGIC;
    SIGNAL S796 : STD_LOGIC;
    SIGNAL S797 : STD_LOGIC;
    SIGNAL S798 : STD_LOGIC;
    SIGNAL S799 : STD_LOGIC;
    SIGNAL S800 : STD_LOGIC;
    SIGNAL S801 : STD_LOGIC;
    SIGNAL S802 : STD_LOGIC;
    SIGNAL S803 : STD_LOGIC;
    SIGNAL S804 : STD_LOGIC;
    SIGNAL S805 : STD_LOGIC;
    SIGNAL S806 : STD_LOGIC;
    SIGNAL S807 : STD_LOGIC;
    SIGNAL S808 : STD_LOGIC;
    SIGNAL S809 : STD_LOGIC;
    SIGNAL S810 : STD_LOGIC;
    SIGNAL S811 : STD_LOGIC;
    SIGNAL S812 : STD_LOGIC;
    SIGNAL S813 : STD_LOGIC;
    SIGNAL S814 : STD_LOGIC;
    SIGNAL S815 : STD_LOGIC;
    SIGNAL S816 : STD_LOGIC;
    SIGNAL S817 : STD_LOGIC;
    SIGNAL S818 : STD_LOGIC;
    SIGNAL S819 : STD_LOGIC;
    SIGNAL S820 : STD_LOGIC;
    SIGNAL S821 : STD_LOGIC;
    SIGNAL S822 : STD_LOGIC;
    SIGNAL S823 : STD_LOGIC;
    SIGNAL S824 : STD_LOGIC;
    SIGNAL S825 : STD_LOGIC;
    SIGNAL S826 : STD_LOGIC;
    SIGNAL S827 : STD_LOGIC;
    SIGNAL S828 : STD_LOGIC;
    SIGNAL S829 : STD_LOGIC;
    SIGNAL S830 : STD_LOGIC;
    SIGNAL S831 : STD_LOGIC;
    SIGNAL S832 : STD_LOGIC;
    SIGNAL S833 : STD_LOGIC;
    SIGNAL S834 : STD_LOGIC;
    SIGNAL S835 : STD_LOGIC;
    SIGNAL S836 : STD_LOGIC;
    SIGNAL S837 : STD_LOGIC;
    SIGNAL S838 : STD_LOGIC;
    SIGNAL S839 : STD_LOGIC;
    SIGNAL S840 : STD_LOGIC;
    SIGNAL S841 : STD_LOGIC;
    SIGNAL S842 : STD_LOGIC;
    SIGNAL S843 : STD_LOGIC;
    SIGNAL S844 : STD_LOGIC;
    SIGNAL S845 : STD_LOGIC;
    SIGNAL S846 : STD_LOGIC;
    SIGNAL S847 : STD_LOGIC;
    SIGNAL S848 : STD_LOGIC;
    SIGNAL S849 : STD_LOGIC;
    SIGNAL S850 : STD_LOGIC;
    SIGNAL S851 : STD_LOGIC;
    SIGNAL S852 : STD_LOGIC;
    SIGNAL S853 : STD_LOGIC;
    SIGNAL S854 : STD_LOGIC;
    SIGNAL S855 : STD_LOGIC;
    SIGNAL S856 : STD_LOGIC;
    SIGNAL S857 : STD_LOGIC;
    SIGNAL S858 : STD_LOGIC;
    SIGNAL S859 : STD_LOGIC;
    SIGNAL S860 : STD_LOGIC;
    SIGNAL S861 : STD_LOGIC;
    SIGNAL S862 : STD_LOGIC;
    SIGNAL S863 : STD_LOGIC;
    SIGNAL S864 : STD_LOGIC;
    SIGNAL S865 : STD_LOGIC;
    SIGNAL S866 : STD_LOGIC;
    SIGNAL S867 : STD_LOGIC;
    SIGNAL S868 : STD_LOGIC;
    SIGNAL S869 : STD_LOGIC;
    SIGNAL S870 : STD_LOGIC;
    SIGNAL S871 : STD_LOGIC;
    SIGNAL S872 : STD_LOGIC;
    SIGNAL S873 : STD_LOGIC;
    SIGNAL S874 : STD_LOGIC;
    SIGNAL S875 : STD_LOGIC;
    SIGNAL S876 : STD_LOGIC;
    SIGNAL S877 : STD_LOGIC;
    SIGNAL S878 : STD_LOGIC;
    SIGNAL S879 : STD_LOGIC;
    SIGNAL S880 : STD_LOGIC;
    SIGNAL S881 : STD_LOGIC;
    SIGNAL S882 : STD_LOGIC;
    SIGNAL S883 : STD_LOGIC;
    SIGNAL S884 : STD_LOGIC;
    SIGNAL S885 : STD_LOGIC;
    SIGNAL S886 : STD_LOGIC;
    SIGNAL S887 : STD_LOGIC;
    SIGNAL S888 : STD_LOGIC;
    SIGNAL S889 : STD_LOGIC;
    SIGNAL S890 : STD_LOGIC;
    SIGNAL S891 : STD_LOGIC;
    SIGNAL S892 : STD_LOGIC;
    SIGNAL S893 : STD_LOGIC;
    SIGNAL S894 : STD_LOGIC;
    SIGNAL S895 : STD_LOGIC;
    SIGNAL S896 : STD_LOGIC;
    SIGNAL S897 : STD_LOGIC;
    SIGNAL S898 : STD_LOGIC;
    SIGNAL S899 : STD_LOGIC;
    SIGNAL S900 : STD_LOGIC;
    SIGNAL S901 : STD_LOGIC;
    SIGNAL S902 : STD_LOGIC;
    SIGNAL S903 : STD_LOGIC;
    SIGNAL S904 : STD_LOGIC;
    SIGNAL S905 : STD_LOGIC;
    SIGNAL S906 : STD_LOGIC;
    SIGNAL S907 : STD_LOGIC;
    SIGNAL S908 : STD_LOGIC;
    SIGNAL S909 : STD_LOGIC;
    SIGNAL S910 : STD_LOGIC;
    SIGNAL S911 : STD_LOGIC;
    SIGNAL S912 : STD_LOGIC;
    SIGNAL S913 : STD_LOGIC;
    SIGNAL S914 : STD_LOGIC;
    SIGNAL S915 : STD_LOGIC;
    SIGNAL S916 : STD_LOGIC;
    SIGNAL S917 : STD_LOGIC;
    SIGNAL S918 : STD_LOGIC;
    SIGNAL S919 : STD_LOGIC;
    SIGNAL S920 : STD_LOGIC;
    SIGNAL S921 : STD_LOGIC;
    SIGNAL S922 : STD_LOGIC;
    SIGNAL S923 : STD_LOGIC;
    SIGNAL S924 : STD_LOGIC;
    SIGNAL S925 : STD_LOGIC;
    SIGNAL S926 : STD_LOGIC;
    SIGNAL S927 : STD_LOGIC;
    SIGNAL S928 : STD_LOGIC;
    SIGNAL S929 : STD_LOGIC;
    SIGNAL S930 : STD_LOGIC;
    SIGNAL S931 : STD_LOGIC;
    SIGNAL S932 : STD_LOGIC;
    SIGNAL S933 : STD_LOGIC;
    SIGNAL S934 : STD_LOGIC;
    SIGNAL S935 : STD_LOGIC;
    SIGNAL S936 : STD_LOGIC;
    SIGNAL S937 : STD_LOGIC;
    SIGNAL S938 : STD_LOGIC;
    SIGNAL S939 : STD_LOGIC;
    SIGNAL S940 : STD_LOGIC;
    SIGNAL S941 : STD_LOGIC;
    SIGNAL S942 : STD_LOGIC;
    SIGNAL S943 : STD_LOGIC;
    SIGNAL S944 : STD_LOGIC;
    SIGNAL S945 : STD_LOGIC;
    SIGNAL S946 : STD_LOGIC;
    SIGNAL S947 : STD_LOGIC;
    SIGNAL S948 : STD_LOGIC;
    SIGNAL S949 : STD_LOGIC;
    SIGNAL S950 : STD_LOGIC;
    SIGNAL S951 : STD_LOGIC;
    SIGNAL S952 : STD_LOGIC;
    SIGNAL S953 : STD_LOGIC;
    SIGNAL S954 : STD_LOGIC;
    SIGNAL S955 : STD_LOGIC;
    SIGNAL S956 : STD_LOGIC;
    SIGNAL S957 : STD_LOGIC;
    SIGNAL S958 : STD_LOGIC;
    SIGNAL S959 : STD_LOGIC;
    SIGNAL S960 : STD_LOGIC;
    SIGNAL S961 : STD_LOGIC;
    SIGNAL S962 : STD_LOGIC;
    SIGNAL S963 : STD_LOGIC;
    SIGNAL S964 : STD_LOGIC;
    SIGNAL S965 : STD_LOGIC;
    SIGNAL S966 : STD_LOGIC;
    SIGNAL S967 : STD_LOGIC;
    SIGNAL S968 : STD_LOGIC;
    SIGNAL S969 : STD_LOGIC;
    SIGNAL S970 : STD_LOGIC;
    SIGNAL S971 : STD_LOGIC;
    SIGNAL S972 : STD_LOGIC;
    SIGNAL S973 : STD_LOGIC;
    SIGNAL S974 : STD_LOGIC;
    SIGNAL S975 : STD_LOGIC;
    SIGNAL S976 : STD_LOGIC;
    SIGNAL S977 : STD_LOGIC;
    SIGNAL S978 : STD_LOGIC;
    SIGNAL S979 : STD_LOGIC;
    SIGNAL S980 : STD_LOGIC;
    SIGNAL S981 : STD_LOGIC;
    SIGNAL S982 : STD_LOGIC;
    SIGNAL S983 : STD_LOGIC;
    SIGNAL S984 : STD_LOGIC;
    SIGNAL S985 : STD_LOGIC;
    SIGNAL S986 : STD_LOGIC;
    SIGNAL S987 : STD_LOGIC;
    SIGNAL S988 : STD_LOGIC;
    SIGNAL S989 : STD_LOGIC;
    SIGNAL S990 : STD_LOGIC;
    SIGNAL S991 : STD_LOGIC;
    SIGNAL S992 : STD_LOGIC;
    SIGNAL S993 : STD_LOGIC;
    SIGNAL S994 : STD_LOGIC;
    SIGNAL S995 : STD_LOGIC;
    SIGNAL S996 : STD_LOGIC;
    SIGNAL S997 : STD_LOGIC;
    SIGNAL S998 : STD_LOGIC;
    SIGNAL S999 : STD_LOGIC;
    SIGNAL S1000 : STD_LOGIC;
    SIGNAL S1001 : STD_LOGIC;
    SIGNAL S1002 : STD_LOGIC;
    SIGNAL S1003 : STD_LOGIC;
    SIGNAL S1004 : STD_LOGIC;
    SIGNAL S1005 : STD_LOGIC;
    SIGNAL S1006 : STD_LOGIC;
    SIGNAL S1007 : STD_LOGIC;
    SIGNAL S1008 : STD_LOGIC;
    SIGNAL S1009 : STD_LOGIC;
    SIGNAL S1010 : STD_LOGIC;
    SIGNAL S1011 : STD_LOGIC;
    SIGNAL S1012 : STD_LOGIC;
    SIGNAL S1013 : STD_LOGIC;
    SIGNAL S1014 : STD_LOGIC;
    SIGNAL S1015 : STD_LOGIC;
    SIGNAL S1016 : STD_LOGIC;
    SIGNAL S1017 : STD_LOGIC;
    SIGNAL S1018 : STD_LOGIC;
    SIGNAL S1019 : STD_LOGIC;
    SIGNAL S1020 : STD_LOGIC;
    SIGNAL S1021 : STD_LOGIC;
    SIGNAL S1022 : STD_LOGIC;
    SIGNAL S1023 : STD_LOGIC;
    SIGNAL S1024 : STD_LOGIC;
    SIGNAL S1025 : STD_LOGIC;
    SIGNAL S1026 : STD_LOGIC;
    SIGNAL S1027 : STD_LOGIC;
    SIGNAL S1028 : STD_LOGIC;
    SIGNAL S1029 : STD_LOGIC;
    SIGNAL S1030 : STD_LOGIC;
    SIGNAL S1031 : STD_LOGIC;
    SIGNAL S1032 : STD_LOGIC;
    SIGNAL S1033 : STD_LOGIC;
    SIGNAL S1034 : STD_LOGIC;
    SIGNAL S1035 : STD_LOGIC;
    SIGNAL S1036 : STD_LOGIC;
    SIGNAL S1037 : STD_LOGIC;
    SIGNAL S1038 : STD_LOGIC;
    SIGNAL S1039 : STD_LOGIC;
    SIGNAL S1040 : STD_LOGIC;
    SIGNAL S1041 : STD_LOGIC;
    SIGNAL S1042 : STD_LOGIC;
    SIGNAL S1043 : STD_LOGIC;
    SIGNAL S1044 : STD_LOGIC;
    SIGNAL S1045 : STD_LOGIC;
    SIGNAL S1046 : STD_LOGIC;
    SIGNAL S1047 : STD_LOGIC;
    SIGNAL S1048 : STD_LOGIC;
    SIGNAL S1049 : STD_LOGIC;
    SIGNAL S1050 : STD_LOGIC;
    SIGNAL S1051 : STD_LOGIC;
    SIGNAL S1052 : STD_LOGIC;
    SIGNAL S1053 : STD_LOGIC;
    SIGNAL S1054 : STD_LOGIC;
    SIGNAL S1055 : STD_LOGIC;
    SIGNAL S1056 : STD_LOGIC;
    SIGNAL S1057 : STD_LOGIC;
    SIGNAL S1058 : STD_LOGIC;
    SIGNAL S1059 : STD_LOGIC;
    SIGNAL S1060 : STD_LOGIC;
    SIGNAL S1061 : STD_LOGIC;
    SIGNAL S1062 : STD_LOGIC;
    SIGNAL S1063 : STD_LOGIC;
    SIGNAL S1064 : STD_LOGIC;
    SIGNAL S1065 : STD_LOGIC;
    SIGNAL S1066 : STD_LOGIC;
    SIGNAL S1067 : STD_LOGIC;
    SIGNAL S1068 : STD_LOGIC;
    SIGNAL S1069 : STD_LOGIC;
    SIGNAL S1070 : STD_LOGIC;
    SIGNAL S1071 : STD_LOGIC;
    SIGNAL S1072 : STD_LOGIC;
    SIGNAL S1073 : STD_LOGIC;
    SIGNAL S1074 : STD_LOGIC;
    SIGNAL S1075 : STD_LOGIC;
    SIGNAL S1076 : STD_LOGIC;
    SIGNAL S1077 : STD_LOGIC;
    SIGNAL S1078 : STD_LOGIC;
    SIGNAL S1079 : STD_LOGIC;
    SIGNAL S1080 : STD_LOGIC;
    SIGNAL S1081 : STD_LOGIC;
    SIGNAL S1082 : STD_LOGIC;
    SIGNAL S1083 : STD_LOGIC;
    SIGNAL S1084 : STD_LOGIC;
    SIGNAL S1085 : STD_LOGIC;
    SIGNAL S1086 : STD_LOGIC;
    SIGNAL S1087 : STD_LOGIC;
    SIGNAL S1088 : STD_LOGIC;
    SIGNAL S1089 : STD_LOGIC;
    SIGNAL S1090 : STD_LOGIC;
    SIGNAL S1091 : STD_LOGIC;
    SIGNAL S1092 : STD_LOGIC;
    SIGNAL S1093 : STD_LOGIC;
    SIGNAL S1094 : STD_LOGIC;
    SIGNAL S1095 : STD_LOGIC;
    SIGNAL S1096 : STD_LOGIC;
    SIGNAL S1097 : STD_LOGIC;
    SIGNAL S1098 : STD_LOGIC;
    SIGNAL S1099 : STD_LOGIC;
    SIGNAL S1100 : STD_LOGIC;
    SIGNAL S1101 : STD_LOGIC;
    SIGNAL S1102 : STD_LOGIC;
    SIGNAL S1103 : STD_LOGIC;
    SIGNAL S1104 : STD_LOGIC;
    SIGNAL S1105 : STD_LOGIC;
    SIGNAL S1106 : STD_LOGIC;
    SIGNAL S1107 : STD_LOGIC;
    SIGNAL S1108 : STD_LOGIC;
    SIGNAL S1109 : STD_LOGIC;
    SIGNAL S1110 : STD_LOGIC;
    SIGNAL S1111 : STD_LOGIC;
    SIGNAL S1112 : STD_LOGIC;
    SIGNAL S1113 : STD_LOGIC;
    SIGNAL S1114 : STD_LOGIC;
    SIGNAL S1115 : STD_LOGIC;
    SIGNAL S1116 : STD_LOGIC;
    SIGNAL S1117 : STD_LOGIC;
    SIGNAL S1118 : STD_LOGIC;
    SIGNAL S1119 : STD_LOGIC;
    SIGNAL S1120 : STD_LOGIC;
    SIGNAL S1121 : STD_LOGIC;
    SIGNAL S1122 : STD_LOGIC;
    SIGNAL S1123 : STD_LOGIC;
    SIGNAL S1124 : STD_LOGIC;
    SIGNAL S1125 : STD_LOGIC;
    SIGNAL S1126 : STD_LOGIC;
    SIGNAL S1127 : STD_LOGIC;
    SIGNAL S1128 : STD_LOGIC;
    SIGNAL S1129 : STD_LOGIC;
    SIGNAL S1130 : STD_LOGIC;
    SIGNAL S1131 : STD_LOGIC;
    SIGNAL S1132 : STD_LOGIC;
    SIGNAL S1133 : STD_LOGIC;
    SIGNAL S1134 : STD_LOGIC;
    SIGNAL S1135 : STD_LOGIC;
    SIGNAL S1136 : STD_LOGIC;
    SIGNAL S1137 : STD_LOGIC;
    SIGNAL S1138 : STD_LOGIC;
    SIGNAL S1139 : STD_LOGIC;
    SIGNAL S1140 : STD_LOGIC;
    SIGNAL S1141 : STD_LOGIC;
    SIGNAL S1142 : STD_LOGIC;
    SIGNAL S1143 : STD_LOGIC;
    SIGNAL S1144 : STD_LOGIC;
    SIGNAL S1145 : STD_LOGIC;
    SIGNAL S1146 : STD_LOGIC;
    SIGNAL S1147 : STD_LOGIC;
    SIGNAL S1148 : STD_LOGIC;
    SIGNAL S1149 : STD_LOGIC;
    SIGNAL S1150 : STD_LOGIC;
    SIGNAL S1151 : STD_LOGIC;
    SIGNAL S1152 : STD_LOGIC;
    SIGNAL S1153 : STD_LOGIC;
    SIGNAL S1154 : STD_LOGIC;
    SIGNAL S1155 : STD_LOGIC;
    SIGNAL S1156 : STD_LOGIC;
    SIGNAL S1157 : STD_LOGIC;
    SIGNAL S1158 : STD_LOGIC;
    SIGNAL S1159 : STD_LOGIC;
    SIGNAL S1160 : STD_LOGIC;
    SIGNAL S1161 : STD_LOGIC;
    SIGNAL S1162 : STD_LOGIC;
    SIGNAL S1163 : STD_LOGIC;
    SIGNAL S1164 : STD_LOGIC;
    SIGNAL S1165 : STD_LOGIC;
    SIGNAL S1166 : STD_LOGIC;
    SIGNAL S1167 : STD_LOGIC;
    SIGNAL S1168 : STD_LOGIC;
    SIGNAL S1169 : STD_LOGIC;
    SIGNAL S1170 : STD_LOGIC;
    SIGNAL S1171 : STD_LOGIC;
    SIGNAL S1172 : STD_LOGIC;
    SIGNAL S1173 : STD_LOGIC;
    SIGNAL S1174 : STD_LOGIC;
    SIGNAL S1175 : STD_LOGIC;
    SIGNAL S1176 : STD_LOGIC;
    SIGNAL S1177 : STD_LOGIC;
    SIGNAL S1178 : STD_LOGIC;
    SIGNAL S1179 : STD_LOGIC;
    SIGNAL S1180 : STD_LOGIC;
    SIGNAL S1181 : STD_LOGIC;
    SIGNAL S1182 : STD_LOGIC;
    SIGNAL S1183 : STD_LOGIC;
    SIGNAL S1184 : STD_LOGIC;
    SIGNAL S1185 : STD_LOGIC;
    SIGNAL S1186 : STD_LOGIC;
    SIGNAL S1187 : STD_LOGIC;
    SIGNAL S1188 : STD_LOGIC;
    SIGNAL S1189 : STD_LOGIC;
    SIGNAL S1190 : STD_LOGIC;
    SIGNAL S1191 : STD_LOGIC;
    SIGNAL S1192 : STD_LOGIC;
    SIGNAL S1193 : STD_LOGIC;
    SIGNAL S1194 : STD_LOGIC;
    SIGNAL S1195 : STD_LOGIC;
    SIGNAL S1196 : STD_LOGIC;
    SIGNAL S1197 : STD_LOGIC;
    SIGNAL S1198 : STD_LOGIC;
    SIGNAL S1199 : STD_LOGIC;
    SIGNAL S1200 : STD_LOGIC;
    SIGNAL S1201 : STD_LOGIC;
    SIGNAL S1202 : STD_LOGIC;
    SIGNAL S1203 : STD_LOGIC;
    SIGNAL S1204 : STD_LOGIC;
    SIGNAL S1205 : STD_LOGIC;
    SIGNAL S1206 : STD_LOGIC;
    SIGNAL S1207 : STD_LOGIC;
    SIGNAL S1208 : STD_LOGIC;
    SIGNAL S1209 : STD_LOGIC;
    SIGNAL S1210 : STD_LOGIC;
    SIGNAL S1211 : STD_LOGIC;
    SIGNAL S1212 : STD_LOGIC;
    SIGNAL S1213 : STD_LOGIC;
    SIGNAL S1214 : STD_LOGIC;
    SIGNAL S1215 : STD_LOGIC;
    SIGNAL S1216 : STD_LOGIC;
    SIGNAL S1217 : STD_LOGIC;
    SIGNAL S1218 : STD_LOGIC;
    SIGNAL S1219 : STD_LOGIC;
    SIGNAL S1220 : STD_LOGIC;
    SIGNAL S1221 : STD_LOGIC;
    SIGNAL S1222 : STD_LOGIC;
    SIGNAL S1223 : STD_LOGIC;
    SIGNAL S1224 : STD_LOGIC;
    SIGNAL S1225 : STD_LOGIC;
    SIGNAL S1226 : STD_LOGIC;
    SIGNAL S1227 : STD_LOGIC;
    SIGNAL S1228 : STD_LOGIC;
    SIGNAL S1229 : STD_LOGIC;
    SIGNAL S1230 : STD_LOGIC;
    SIGNAL S1231 : STD_LOGIC;
    SIGNAL S1232 : STD_LOGIC;
    SIGNAL S1233 : STD_LOGIC;
    SIGNAL S1234 : STD_LOGIC;
    SIGNAL S1235 : STD_LOGIC;
    SIGNAL S1236 : STD_LOGIC;
    SIGNAL S1237 : STD_LOGIC;
    SIGNAL S1238 : STD_LOGIC;
    SIGNAL S1239 : STD_LOGIC;
    SIGNAL S1240 : STD_LOGIC;
    SIGNAL S1241 : STD_LOGIC;
    SIGNAL S1242 : STD_LOGIC;
    SIGNAL S1243 : STD_LOGIC;
    SIGNAL S1244 : STD_LOGIC;
    SIGNAL S1245 : STD_LOGIC;
    SIGNAL S1246 : STD_LOGIC;
    SIGNAL S1247 : STD_LOGIC;
    SIGNAL S1248 : STD_LOGIC;
    SIGNAL S1249 : STD_LOGIC;
    SIGNAL S1250 : STD_LOGIC;
    SIGNAL S1251 : STD_LOGIC;
    SIGNAL S1252 : STD_LOGIC;
    SIGNAL S1253 : STD_LOGIC;
    SIGNAL S1254 : STD_LOGIC;
    SIGNAL S1255 : STD_LOGIC;
    SIGNAL S1256 : STD_LOGIC;
    SIGNAL S1257 : STD_LOGIC;
    SIGNAL S1258 : STD_LOGIC;
    SIGNAL S1259 : STD_LOGIC;
    SIGNAL S1260 : STD_LOGIC;
    SIGNAL S1261 : STD_LOGIC;
    SIGNAL S1262 : STD_LOGIC;
    SIGNAL S1263 : STD_LOGIC;
    SIGNAL S1264 : STD_LOGIC;
    SIGNAL S1265 : STD_LOGIC;
    SIGNAL S1266 : STD_LOGIC;
    SIGNAL S1267 : STD_LOGIC;
    SIGNAL S1268 : STD_LOGIC;
    SIGNAL S1269 : STD_LOGIC;
    SIGNAL S1270 : STD_LOGIC;
    SIGNAL S1271 : STD_LOGIC;
    SIGNAL S1272 : STD_LOGIC;
    SIGNAL S1273 : STD_LOGIC;
    SIGNAL S1274 : STD_LOGIC;
    SIGNAL S1275 : STD_LOGIC;
    SIGNAL S1276 : STD_LOGIC;
    SIGNAL S1277 : STD_LOGIC;
    SIGNAL S1278 : STD_LOGIC;
    SIGNAL S1279 : STD_LOGIC;
    SIGNAL S1280 : STD_LOGIC;
    SIGNAL S1281 : STD_LOGIC;
    SIGNAL S1282 : STD_LOGIC;
    SIGNAL S1283 : STD_LOGIC;
    SIGNAL S1284 : STD_LOGIC;
    SIGNAL S1285 : STD_LOGIC;
    SIGNAL S1286 : STD_LOGIC;
    SIGNAL S1287 : STD_LOGIC;
    SIGNAL S1288 : STD_LOGIC;
    SIGNAL S1289 : STD_LOGIC;
    SIGNAL S1290 : STD_LOGIC;
    SIGNAL S1291 : STD_LOGIC;
    SIGNAL S1292 : STD_LOGIC;
    SIGNAL S1293 : STD_LOGIC;
    SIGNAL S1294 : STD_LOGIC;
    SIGNAL S1295 : STD_LOGIC;
    SIGNAL S1296 : STD_LOGIC;
    SIGNAL S1297 : STD_LOGIC;
    SIGNAL S1298 : STD_LOGIC;
    SIGNAL S1299 : STD_LOGIC;
    SIGNAL S1300 : STD_LOGIC;
    SIGNAL S1301 : STD_LOGIC;
    SIGNAL S1302 : STD_LOGIC;
    SIGNAL S1303 : STD_LOGIC;
    SIGNAL S1304 : STD_LOGIC;
    SIGNAL S1305 : STD_LOGIC;
    SIGNAL S1306 : STD_LOGIC;
    SIGNAL S1307 : STD_LOGIC;
    SIGNAL S1308 : STD_LOGIC;
    SIGNAL S1309 : STD_LOGIC;
    SIGNAL S1310 : STD_LOGIC;
    SIGNAL S1311 : STD_LOGIC;
    SIGNAL S1312 : STD_LOGIC;
    SIGNAL S1313 : STD_LOGIC;
    SIGNAL S1314 : STD_LOGIC;
    SIGNAL S1315 : STD_LOGIC;
    SIGNAL S1316 : STD_LOGIC;
    SIGNAL S1317 : STD_LOGIC;
    SIGNAL S1318 : STD_LOGIC;
    SIGNAL S1319 : STD_LOGIC;
    SIGNAL S1320 : STD_LOGIC;
    SIGNAL S1321 : STD_LOGIC;
    SIGNAL S1322 : STD_LOGIC;
    SIGNAL S1323 : STD_LOGIC;
    SIGNAL S1324 : STD_LOGIC;
    SIGNAL S1325 : STD_LOGIC;
    SIGNAL S1326 : STD_LOGIC;
    SIGNAL S1327 : STD_LOGIC;
    SIGNAL S1328 : STD_LOGIC;
    SIGNAL S1329 : STD_LOGIC;
    SIGNAL S1330 : STD_LOGIC;
    SIGNAL S1331 : STD_LOGIC;
    SIGNAL S1332 : STD_LOGIC;
    SIGNAL S1333 : STD_LOGIC;
    SIGNAL S1334 : STD_LOGIC;
    SIGNAL S1335 : STD_LOGIC;
    SIGNAL S1336 : STD_LOGIC;
    SIGNAL S1337 : STD_LOGIC;
    SIGNAL S1338 : STD_LOGIC;
    SIGNAL S1339 : STD_LOGIC;
    SIGNAL S1340 : STD_LOGIC;
    SIGNAL S1341 : STD_LOGIC;
    SIGNAL S1342 : STD_LOGIC;
    SIGNAL S1343 : STD_LOGIC;
    SIGNAL S1344 : STD_LOGIC;
    SIGNAL S1345 : STD_LOGIC;
    SIGNAL S1346 : STD_LOGIC;
    SIGNAL S1347 : STD_LOGIC;
    SIGNAL S1348 : STD_LOGIC;
    SIGNAL S1349 : STD_LOGIC;
    SIGNAL S1350 : STD_LOGIC;
    SIGNAL S1351 : STD_LOGIC;
    SIGNAL S1352 : STD_LOGIC;
    SIGNAL S1353 : STD_LOGIC;
    SIGNAL S1354 : STD_LOGIC;
    SIGNAL S1355 : STD_LOGIC;
    SIGNAL S1356 : STD_LOGIC;
    SIGNAL S1357 : STD_LOGIC;
    SIGNAL S1358 : STD_LOGIC;
    SIGNAL S1359 : STD_LOGIC;
    SIGNAL S1360 : STD_LOGIC;
    SIGNAL S1361 : STD_LOGIC;
    SIGNAL S1362 : STD_LOGIC;
    SIGNAL S1363 : STD_LOGIC;
    SIGNAL S1364 : STD_LOGIC;
    SIGNAL S1365 : STD_LOGIC;
    SIGNAL S1366 : STD_LOGIC;
    SIGNAL S1367 : STD_LOGIC;
    SIGNAL S1368 : STD_LOGIC;
    SIGNAL S1369 : STD_LOGIC;
    SIGNAL S1370 : STD_LOGIC;
    SIGNAL S1371 : STD_LOGIC;
    SIGNAL S1372 : STD_LOGIC;
    SIGNAL S1373 : STD_LOGIC;
    SIGNAL S1374 : STD_LOGIC;
    SIGNAL S1375 : STD_LOGIC;
    SIGNAL S1376 : STD_LOGIC;
    SIGNAL S1377 : STD_LOGIC;
    SIGNAL S1378 : STD_LOGIC;
    SIGNAL S1379 : STD_LOGIC;
    SIGNAL S1380 : STD_LOGIC;
    SIGNAL S1381 : STD_LOGIC;
    SIGNAL S1382 : STD_LOGIC;
    SIGNAL S1383 : STD_LOGIC;
    SIGNAL S1384 : STD_LOGIC;
    SIGNAL S1385 : STD_LOGIC;
    SIGNAL S1386 : STD_LOGIC;
    SIGNAL S1387 : STD_LOGIC;
    SIGNAL S1388 : STD_LOGIC;
    SIGNAL S1389 : STD_LOGIC;
    SIGNAL S1390 : STD_LOGIC;
    SIGNAL S1391 : STD_LOGIC;
    SIGNAL S1392 : STD_LOGIC;
    SIGNAL S1393 : STD_LOGIC;
    SIGNAL S1394 : STD_LOGIC;
    SIGNAL S1395 : STD_LOGIC;
    SIGNAL S1396 : STD_LOGIC;
    SIGNAL S1397 : STD_LOGIC;
    SIGNAL S1398 : STD_LOGIC;
    SIGNAL S1399 : STD_LOGIC;
    SIGNAL S1400 : STD_LOGIC;
    SIGNAL S1401 : STD_LOGIC;
    SIGNAL S1402 : STD_LOGIC;
    SIGNAL S1403 : STD_LOGIC;
    SIGNAL S1404 : STD_LOGIC;
    SIGNAL S1405 : STD_LOGIC;
    SIGNAL S1406 : STD_LOGIC;
    SIGNAL S1407 : STD_LOGIC;
    SIGNAL S1408 : STD_LOGIC;
    SIGNAL S1409 : STD_LOGIC;
    SIGNAL S1410 : STD_LOGIC;
    SIGNAL S1411 : STD_LOGIC;
    SIGNAL S1412 : STD_LOGIC;
    SIGNAL S1413 : STD_LOGIC;
    SIGNAL S1414 : STD_LOGIC;
    SIGNAL S1415 : STD_LOGIC;
    SIGNAL S1416 : STD_LOGIC;
    SIGNAL S1417 : STD_LOGIC;
    SIGNAL S1418 : STD_LOGIC;
    SIGNAL S1419 : STD_LOGIC;
    SIGNAL S1420 : STD_LOGIC;
    SIGNAL S1421 : STD_LOGIC;
    SIGNAL S1422 : STD_LOGIC;
    SIGNAL S1423 : STD_LOGIC;
    SIGNAL S1424 : STD_LOGIC;
    SIGNAL S1425 : STD_LOGIC;
    SIGNAL S1426 : STD_LOGIC;
    SIGNAL S1427 : STD_LOGIC;
    SIGNAL S1428 : STD_LOGIC;
    SIGNAL S1429 : STD_LOGIC;
    SIGNAL S1430 : STD_LOGIC;
    SIGNAL S1431 : STD_LOGIC;
    SIGNAL S1432 : STD_LOGIC;
    SIGNAL S1433 : STD_LOGIC;
    SIGNAL S1434 : STD_LOGIC;
    SIGNAL S1435 : STD_LOGIC;
    SIGNAL S1436 : STD_LOGIC;
    SIGNAL S1437 : STD_LOGIC;
    SIGNAL S1438 : STD_LOGIC;
    SIGNAL S1439 : STD_LOGIC;
    SIGNAL S1440 : STD_LOGIC;
    SIGNAL S1441 : STD_LOGIC;
    SIGNAL S1442 : STD_LOGIC;
    SIGNAL S1443 : STD_LOGIC;
    SIGNAL S1444 : STD_LOGIC;
    SIGNAL S1445 : STD_LOGIC;
    SIGNAL S1446 : STD_LOGIC;
    SIGNAL S1447 : STD_LOGIC;
    SIGNAL S1448 : STD_LOGIC;
    SIGNAL S1449 : STD_LOGIC;
    SIGNAL S1450 : STD_LOGIC;
    SIGNAL S1451 : STD_LOGIC;
    SIGNAL S1452 : STD_LOGIC;
    SIGNAL S1453 : STD_LOGIC;
    SIGNAL S1454 : STD_LOGIC;
    SIGNAL S1455 : STD_LOGIC;
    SIGNAL S1456 : STD_LOGIC;
    SIGNAL S1457 : STD_LOGIC;
    SIGNAL S1458 : STD_LOGIC;
    SIGNAL S1459 : STD_LOGIC;
    SIGNAL S1460 : STD_LOGIC;
    SIGNAL S1461 : STD_LOGIC;
    SIGNAL S1462 : STD_LOGIC;
    SIGNAL S1463 : STD_LOGIC;
    SIGNAL S1464 : STD_LOGIC;
    SIGNAL S1465 : STD_LOGIC;
    SIGNAL S1466 : STD_LOGIC;
    SIGNAL S1467 : STD_LOGIC;
    SIGNAL S1468 : STD_LOGIC;
    SIGNAL S1469 : STD_LOGIC;
    SIGNAL S1470 : STD_LOGIC;
    SIGNAL S1471 : STD_LOGIC;
    SIGNAL S1472 : STD_LOGIC;
    SIGNAL S1473 : STD_LOGIC;
    SIGNAL S1474 : STD_LOGIC;
    SIGNAL S1475 : STD_LOGIC;
    SIGNAL S1476 : STD_LOGIC;
    SIGNAL S1477 : STD_LOGIC;
    SIGNAL S1478 : STD_LOGIC;
    SIGNAL S1479 : STD_LOGIC;
    SIGNAL S1480 : STD_LOGIC;
    SIGNAL S1481 : STD_LOGIC;
    SIGNAL S1482 : STD_LOGIC;
    SIGNAL S1483 : STD_LOGIC;
    SIGNAL S1484 : STD_LOGIC;
    SIGNAL S1485 : STD_LOGIC;
    SIGNAL S1486 : STD_LOGIC;
    SIGNAL S1487 : STD_LOGIC;
    SIGNAL S1488 : STD_LOGIC;
    SIGNAL S1489 : STD_LOGIC;
    SIGNAL S1490 : STD_LOGIC;
    SIGNAL S1491 : STD_LOGIC;
    SIGNAL S1492 : STD_LOGIC;
    SIGNAL S1493 : STD_LOGIC;
    SIGNAL S1494 : STD_LOGIC;
    SIGNAL S1495 : STD_LOGIC;
    SIGNAL S1496 : STD_LOGIC;
    SIGNAL S1497 : STD_LOGIC;
    SIGNAL S1498 : STD_LOGIC;
    SIGNAL S1499 : STD_LOGIC;
    SIGNAL S1500 : STD_LOGIC;
    SIGNAL S1501 : STD_LOGIC;
    SIGNAL S1502 : STD_LOGIC;
    SIGNAL S1503 : STD_LOGIC;
    SIGNAL S1504 : STD_LOGIC;
    SIGNAL S1505 : STD_LOGIC;
    SIGNAL S1506 : STD_LOGIC;
    SIGNAL S1507 : STD_LOGIC;
    SIGNAL S1508 : STD_LOGIC;
    SIGNAL S1509 : STD_LOGIC;
    SIGNAL S1510 : STD_LOGIC;
    SIGNAL S1511 : STD_LOGIC;
    SIGNAL S1512 : STD_LOGIC;
    SIGNAL S1513 : STD_LOGIC;
    SIGNAL S1514 : STD_LOGIC;
    SIGNAL S1515 : STD_LOGIC;
    SIGNAL S1516 : STD_LOGIC;
    SIGNAL S1517 : STD_LOGIC;
    SIGNAL S1518 : STD_LOGIC;
    SIGNAL S1519 : STD_LOGIC;
    SIGNAL S1520 : STD_LOGIC;
    SIGNAL S1521 : STD_LOGIC;
    SIGNAL S1522 : STD_LOGIC;
    SIGNAL S1523 : STD_LOGIC;
    SIGNAL S1524 : STD_LOGIC;
    SIGNAL S1525 : STD_LOGIC;
    SIGNAL S1526 : STD_LOGIC;
    SIGNAL S1527 : STD_LOGIC;
    SIGNAL S1528 : STD_LOGIC;
    SIGNAL S1529 : STD_LOGIC;
    SIGNAL S1530 : STD_LOGIC;
    SIGNAL S1531 : STD_LOGIC;
    SIGNAL S1532 : STD_LOGIC;
    SIGNAL S1533 : STD_LOGIC;
    SIGNAL S1534 : STD_LOGIC;
    SIGNAL S1535 : STD_LOGIC;
    SIGNAL S1536 : STD_LOGIC;
    SIGNAL S1537 : STD_LOGIC;
    SIGNAL S1538 : STD_LOGIC;
    SIGNAL S1539 : STD_LOGIC;
    SIGNAL S1540 : STD_LOGIC;
    SIGNAL S1541 : STD_LOGIC;
    SIGNAL S1542 : STD_LOGIC;
    SIGNAL S1543 : STD_LOGIC;
    SIGNAL S1544 : STD_LOGIC;
    SIGNAL S1545 : STD_LOGIC;
    SIGNAL S1546 : STD_LOGIC;
    SIGNAL S1547 : STD_LOGIC;
    SIGNAL S1548 : STD_LOGIC;
    SIGNAL S1549 : STD_LOGIC;
    SIGNAL S1550 : STD_LOGIC;
    SIGNAL S1551 : STD_LOGIC;
    SIGNAL S1552 : STD_LOGIC;
    SIGNAL S1553 : STD_LOGIC;
    SIGNAL S1554 : STD_LOGIC;
    SIGNAL S1555 : STD_LOGIC;
    SIGNAL S1556 : STD_LOGIC;
    SIGNAL S1557 : STD_LOGIC;
    SIGNAL S1558 : STD_LOGIC;
    SIGNAL S1559 : STD_LOGIC;
    SIGNAL S1560 : STD_LOGIC;
    SIGNAL S1561 : STD_LOGIC;
    SIGNAL S1562 : STD_LOGIC;
    SIGNAL S1563 : STD_LOGIC;
    SIGNAL S1564 : STD_LOGIC;
    SIGNAL S1565 : STD_LOGIC;
    SIGNAL S1566 : STD_LOGIC;
    SIGNAL S1567 : STD_LOGIC;
    SIGNAL S1568 : STD_LOGIC;
    SIGNAL S1569 : STD_LOGIC;
    SIGNAL S1570 : STD_LOGIC;
    SIGNAL S1571 : STD_LOGIC;
    SIGNAL S1572 : STD_LOGIC;
    SIGNAL S1573 : STD_LOGIC;
    SIGNAL S1574 : STD_LOGIC;
    SIGNAL S1575 : STD_LOGIC;
    SIGNAL S1576 : STD_LOGIC;
    SIGNAL S1577 : STD_LOGIC;
    SIGNAL S1578 : STD_LOGIC;
    SIGNAL S1579 : STD_LOGIC;
    SIGNAL S1580 : STD_LOGIC;
    SIGNAL S1581 : STD_LOGIC;
    SIGNAL S1582 : STD_LOGIC;
    SIGNAL S1583 : STD_LOGIC;
    SIGNAL S1584 : STD_LOGIC;
    SIGNAL S1585 : STD_LOGIC;
    SIGNAL S1586 : STD_LOGIC;
    SIGNAL S1587 : STD_LOGIC;
    SIGNAL S1588 : STD_LOGIC;
    SIGNAL S1589 : STD_LOGIC;
    SIGNAL S1590 : STD_LOGIC;
    SIGNAL S1591 : STD_LOGIC;
    SIGNAL S1592 : STD_LOGIC;
    SIGNAL S1593 : STD_LOGIC;
    SIGNAL S1594 : STD_LOGIC;
    SIGNAL S1595 : STD_LOGIC;
    SIGNAL S1596 : STD_LOGIC;
    SIGNAL S1597 : STD_LOGIC;
    SIGNAL S1598 : STD_LOGIC;
    SIGNAL S1599 : STD_LOGIC;
    SIGNAL S1600 : STD_LOGIC;
    SIGNAL S1601 : STD_LOGIC;
    SIGNAL S1602 : STD_LOGIC;
    SIGNAL S1603 : STD_LOGIC;
    SIGNAL S1604 : STD_LOGIC;
    SIGNAL S1605 : STD_LOGIC;
    SIGNAL S1606 : STD_LOGIC;
    SIGNAL S1607 : STD_LOGIC;
    SIGNAL S1608 : STD_LOGIC;
    SIGNAL S1609 : STD_LOGIC;
    SIGNAL S1610 : STD_LOGIC;
    SIGNAL S1611 : STD_LOGIC;
    SIGNAL S1612 : STD_LOGIC;
    SIGNAL S1613 : STD_LOGIC;
    SIGNAL S1614 : STD_LOGIC;
    SIGNAL S1615 : STD_LOGIC;
    SIGNAL S1616 : STD_LOGIC;
    SIGNAL S1617 : STD_LOGIC;
    SIGNAL S1618 : STD_LOGIC;
    SIGNAL S1619 : STD_LOGIC;
    SIGNAL S1620 : STD_LOGIC;
    SIGNAL S1621 : STD_LOGIC;
    SIGNAL S1622 : STD_LOGIC;
    SIGNAL S1623 : STD_LOGIC;
    SIGNAL S1624 : STD_LOGIC;
    SIGNAL S1625 : STD_LOGIC;
    SIGNAL S1626 : STD_LOGIC;
    SIGNAL S1627 : STD_LOGIC;
    SIGNAL S1628 : STD_LOGIC;
    SIGNAL S1629 : STD_LOGIC;
    SIGNAL S1630 : STD_LOGIC;
    SIGNAL S1631 : STD_LOGIC;
    SIGNAL S1632 : STD_LOGIC;
    SIGNAL S1633 : STD_LOGIC;
    SIGNAL S1634 : STD_LOGIC;
    SIGNAL S1635 : STD_LOGIC;
    SIGNAL S1636 : STD_LOGIC;
    SIGNAL S1637 : STD_LOGIC;
    SIGNAL S1638 : STD_LOGIC;
    SIGNAL S1639 : STD_LOGIC;
    SIGNAL S1640 : STD_LOGIC;
    SIGNAL S1641 : STD_LOGIC;
    SIGNAL S1642 : STD_LOGIC;
    SIGNAL S1643 : STD_LOGIC;
    SIGNAL S1644 : STD_LOGIC;
    SIGNAL S1645 : STD_LOGIC;
    SIGNAL S1646 : STD_LOGIC;
    SIGNAL S1647 : STD_LOGIC;
    SIGNAL S1648 : STD_LOGIC;
    SIGNAL S1649 : STD_LOGIC;
    SIGNAL S1650 : STD_LOGIC;
    SIGNAL S1651 : STD_LOGIC;
    SIGNAL S1652 : STD_LOGIC;
    SIGNAL S1653 : STD_LOGIC;
    SIGNAL S1654 : STD_LOGIC;
    SIGNAL S1655 : STD_LOGIC;
    SIGNAL S1656 : STD_LOGIC;
    SIGNAL S1657 : STD_LOGIC;
    SIGNAL S1658 : STD_LOGIC;
    SIGNAL S1659 : STD_LOGIC;
    SIGNAL S1660 : STD_LOGIC;
    SIGNAL S1661 : STD_LOGIC;
    SIGNAL S1662 : STD_LOGIC;
    SIGNAL S1663 : STD_LOGIC;
    SIGNAL S1664 : STD_LOGIC;
    SIGNAL S1665 : STD_LOGIC;
    SIGNAL S1666 : STD_LOGIC;
    SIGNAL S1667 : STD_LOGIC;
    SIGNAL S1668 : STD_LOGIC;
    SIGNAL S1669 : STD_LOGIC;
    SIGNAL S1670 : STD_LOGIC;
    SIGNAL S1671 : STD_LOGIC;
    SIGNAL S1672 : STD_LOGIC;
    SIGNAL S1673 : STD_LOGIC;
    SIGNAL S1674 : STD_LOGIC;
    SIGNAL S1675 : STD_LOGIC;
    SIGNAL S1676 : STD_LOGIC;
    SIGNAL S1677 : STD_LOGIC;
    SIGNAL S1678 : STD_LOGIC;
    SIGNAL S1679 : STD_LOGIC;
    SIGNAL S1680 : STD_LOGIC;
    SIGNAL S1681 : STD_LOGIC;
    SIGNAL S1682 : STD_LOGIC;
    SIGNAL S1683 : STD_LOGIC;
    SIGNAL S1684 : STD_LOGIC;
    SIGNAL S1685 : STD_LOGIC;
    SIGNAL S1686 : STD_LOGIC;
    SIGNAL S1687 : STD_LOGIC;
    SIGNAL S1688 : STD_LOGIC;
    SIGNAL S1689 : STD_LOGIC;
    SIGNAL S1690 : STD_LOGIC;
    SIGNAL S1691 : STD_LOGIC;
    SIGNAL S1692 : STD_LOGIC;
    SIGNAL S1693 : STD_LOGIC;
    SIGNAL S1694 : STD_LOGIC;
    SIGNAL S1695 : STD_LOGIC;
    SIGNAL S1696 : STD_LOGIC;
    SIGNAL S1697 : STD_LOGIC;
    SIGNAL S1698 : STD_LOGIC;
    SIGNAL S1699 : STD_LOGIC;
    SIGNAL S1700 : STD_LOGIC;
    SIGNAL S1701 : STD_LOGIC;
    SIGNAL S1702 : STD_LOGIC;
    SIGNAL S1703 : STD_LOGIC;
    SIGNAL S1704 : STD_LOGIC;
    SIGNAL S1705 : STD_LOGIC;
    SIGNAL S1706 : STD_LOGIC;
    SIGNAL S1707 : STD_LOGIC;
    SIGNAL S1708 : STD_LOGIC;
    SIGNAL S1709 : STD_LOGIC;
    SIGNAL S1710 : STD_LOGIC;
    SIGNAL S1711 : STD_LOGIC;
    SIGNAL S1712 : STD_LOGIC;
    SIGNAL S1713 : STD_LOGIC;
    SIGNAL S1714 : STD_LOGIC;
    SIGNAL S1715 : STD_LOGIC;
    SIGNAL S1716 : STD_LOGIC;
    SIGNAL S1717 : STD_LOGIC;
    SIGNAL S1718 : STD_LOGIC;
    SIGNAL S1719 : STD_LOGIC;
    SIGNAL S1720 : STD_LOGIC;
    SIGNAL S1721 : STD_LOGIC;
    SIGNAL S1722 : STD_LOGIC;
    SIGNAL S1723 : STD_LOGIC;
    SIGNAL S1724 : STD_LOGIC;
    SIGNAL S1725 : STD_LOGIC;
    SIGNAL S1726 : STD_LOGIC;
    SIGNAL S1727 : STD_LOGIC;
    SIGNAL S1728 : STD_LOGIC;
    SIGNAL S1729 : STD_LOGIC;
    SIGNAL S1730 : STD_LOGIC;
    SIGNAL S1731 : STD_LOGIC;
    SIGNAL S1732 : STD_LOGIC;
    SIGNAL S1733 : STD_LOGIC;
    SIGNAL S1734 : STD_LOGIC;
    SIGNAL S1735 : STD_LOGIC;
    SIGNAL S1736 : STD_LOGIC;
    SIGNAL S1737 : STD_LOGIC;
    SIGNAL S1738 : STD_LOGIC;
    SIGNAL S1739 : STD_LOGIC;
    SIGNAL S1740 : STD_LOGIC;
    SIGNAL S1741 : STD_LOGIC;
    SIGNAL S1742 : STD_LOGIC;
    SIGNAL S1743 : STD_LOGIC;
    SIGNAL S1744 : STD_LOGIC;
    SIGNAL S1745 : STD_LOGIC;
    SIGNAL S1746 : STD_LOGIC;
    SIGNAL S1747 : STD_LOGIC;
    SIGNAL S1748 : STD_LOGIC;
    SIGNAL S1749 : STD_LOGIC;
    SIGNAL S1750 : STD_LOGIC;
    SIGNAL S1751 : STD_LOGIC;
    SIGNAL S1752 : STD_LOGIC;
    SIGNAL S1753 : STD_LOGIC;
    SIGNAL S1754 : STD_LOGIC;
    SIGNAL S1755 : STD_LOGIC;
    SIGNAL S1756 : STD_LOGIC;
    SIGNAL S1757 : STD_LOGIC;
    SIGNAL S1758 : STD_LOGIC;
    SIGNAL S1759 : STD_LOGIC;
    SIGNAL S1760 : STD_LOGIC;
    SIGNAL S1761 : STD_LOGIC;
    SIGNAL S1762 : STD_LOGIC;
    SIGNAL S1763 : STD_LOGIC;
    SIGNAL S1764 : STD_LOGIC;
    SIGNAL S1765 : STD_LOGIC;
    SIGNAL S1766 : STD_LOGIC;
    SIGNAL S1767 : STD_LOGIC;
    SIGNAL S1768 : STD_LOGIC;
    SIGNAL S1769 : STD_LOGIC;
    SIGNAL S1770 : STD_LOGIC;
    SIGNAL S1771 : STD_LOGIC;
    SIGNAL S1772 : STD_LOGIC;
    SIGNAL S1773 : STD_LOGIC;
    SIGNAL S1774 : STD_LOGIC;
    SIGNAL S1775 : STD_LOGIC;
    SIGNAL S1776 : STD_LOGIC;
    SIGNAL S1777 : STD_LOGIC;
    SIGNAL S1778 : STD_LOGIC;
    SIGNAL S1779 : STD_LOGIC;
    SIGNAL S1780 : STD_LOGIC;
    SIGNAL S1781 : STD_LOGIC;
    SIGNAL S1782 : STD_LOGIC;
    SIGNAL S1783 : STD_LOGIC;
    SIGNAL S1784 : STD_LOGIC;
    SIGNAL S1785 : STD_LOGIC;
    SIGNAL S1786 : STD_LOGIC;
    SIGNAL S1787 : STD_LOGIC;
    SIGNAL S1788 : STD_LOGIC;
    SIGNAL S1789 : STD_LOGIC;
    SIGNAL S1790 : STD_LOGIC;
    SIGNAL S1791 : STD_LOGIC;
    SIGNAL S1792 : STD_LOGIC;
    SIGNAL S1793 : STD_LOGIC;
    SIGNAL S1794 : STD_LOGIC;
    SIGNAL S1795 : STD_LOGIC;
    SIGNAL S1796 : STD_LOGIC;
    SIGNAL S1797 : STD_LOGIC;
    SIGNAL S1798 : STD_LOGIC;
    SIGNAL S1799 : STD_LOGIC;
    SIGNAL S1800 : STD_LOGIC;
    SIGNAL S1801 : STD_LOGIC;
    SIGNAL S1802 : STD_LOGIC;
    SIGNAL S1803 : STD_LOGIC;
    SIGNAL S1804 : STD_LOGIC;
    SIGNAL S1805 : STD_LOGIC;
    SIGNAL S1806 : STD_LOGIC;
    SIGNAL S1807 : STD_LOGIC;
    SIGNAL S1808 : STD_LOGIC;
    SIGNAL S1809 : STD_LOGIC;
    SIGNAL S1810 : STD_LOGIC;
    SIGNAL S1811 : STD_LOGIC;
    SIGNAL S1812 : STD_LOGIC;
    SIGNAL S1813 : STD_LOGIC;
    SIGNAL S1814 : STD_LOGIC;
    SIGNAL S1815 : STD_LOGIC;
    SIGNAL S1816 : STD_LOGIC;
    SIGNAL S1817 : STD_LOGIC;
    SIGNAL S1818 : STD_LOGIC;
    SIGNAL S1819 : STD_LOGIC;
    SIGNAL S1820 : STD_LOGIC;
    SIGNAL S1821 : STD_LOGIC;
    SIGNAL S1822 : STD_LOGIC;
    SIGNAL S1823 : STD_LOGIC;
    SIGNAL S1824 : STD_LOGIC;
    SIGNAL S1825 : STD_LOGIC;
    SIGNAL S1826 : STD_LOGIC;
    SIGNAL S1827 : STD_LOGIC;
    SIGNAL S1828 : STD_LOGIC;
    SIGNAL S1829 : STD_LOGIC;
    SIGNAL S1830 : STD_LOGIC;
    SIGNAL S1831 : STD_LOGIC;
    SIGNAL S1832 : STD_LOGIC;
    SIGNAL S1833 : STD_LOGIC;
    SIGNAL S1834 : STD_LOGIC;
    SIGNAL S1835 : STD_LOGIC;
    SIGNAL S1836 : STD_LOGIC;
    SIGNAL S1837 : STD_LOGIC;
    SIGNAL S1838 : STD_LOGIC;
    SIGNAL S1839 : STD_LOGIC;
    SIGNAL S1840 : STD_LOGIC;
    SIGNAL S1841 : STD_LOGIC;
    SIGNAL S1842 : STD_LOGIC;
    SIGNAL S1843 : STD_LOGIC;
    SIGNAL S1844 : STD_LOGIC;
    SIGNAL S1845 : STD_LOGIC;
    SIGNAL S1846 : STD_LOGIC;
    SIGNAL S1847 : STD_LOGIC;
    SIGNAL S1848 : STD_LOGIC;
    SIGNAL S1849 : STD_LOGIC;
    SIGNAL S1850 : STD_LOGIC;
    SIGNAL S1851 : STD_LOGIC;
    SIGNAL S1852 : STD_LOGIC;
    SIGNAL S1853 : STD_LOGIC;
    SIGNAL S1854 : STD_LOGIC;
    SIGNAL S1855 : STD_LOGIC;
    SIGNAL S1856 : STD_LOGIC;
    SIGNAL S1857 : STD_LOGIC;
    SIGNAL S1858 : STD_LOGIC;
    SIGNAL S1859 : STD_LOGIC;
    SIGNAL S1860 : STD_LOGIC;
    SIGNAL S1861 : STD_LOGIC;
    SIGNAL S1862 : STD_LOGIC;
    SIGNAL S1863 : STD_LOGIC;
    SIGNAL S1864 : STD_LOGIC;
    SIGNAL S1865 : STD_LOGIC;
    SIGNAL S1866 : STD_LOGIC;
    SIGNAL S1867 : STD_LOGIC;
    SIGNAL S1868 : STD_LOGIC;
    SIGNAL S1869 : STD_LOGIC;
    SIGNAL S1870 : STD_LOGIC;
    SIGNAL S1871 : STD_LOGIC;
    SIGNAL S1872 : STD_LOGIC;
    SIGNAL S1873 : STD_LOGIC;
    SIGNAL S1874 : STD_LOGIC;
    SIGNAL S1875 : STD_LOGIC;
    SIGNAL S1876 : STD_LOGIC;
    SIGNAL S1877 : STD_LOGIC;
    SIGNAL S1878 : STD_LOGIC;
    SIGNAL S1879 : STD_LOGIC;
    SIGNAL S1880 : STD_LOGIC;
    SIGNAL S1881 : STD_LOGIC;
    SIGNAL S1882 : STD_LOGIC;
    SIGNAL S1883 : STD_LOGIC;
    SIGNAL S1884 : STD_LOGIC;
    SIGNAL S1885 : STD_LOGIC;
    SIGNAL S1886 : STD_LOGIC;
    SIGNAL S1887 : STD_LOGIC;
    SIGNAL S1888 : STD_LOGIC;
    SIGNAL S1889 : STD_LOGIC;
    SIGNAL S1890 : STD_LOGIC;
    SIGNAL S1891 : STD_LOGIC;
    SIGNAL S1892 : STD_LOGIC;
    SIGNAL S1893 : STD_LOGIC;
    SIGNAL S1894 : STD_LOGIC;
    SIGNAL S1895 : STD_LOGIC;
    SIGNAL S1896 : STD_LOGIC;
    SIGNAL S1897 : STD_LOGIC;
    SIGNAL S1898 : STD_LOGIC;
    SIGNAL S1899 : STD_LOGIC;
    SIGNAL S1900 : STD_LOGIC;
    SIGNAL S1901 : STD_LOGIC;
    SIGNAL S1902 : STD_LOGIC;
    SIGNAL S1903 : STD_LOGIC;
    SIGNAL S1904 : STD_LOGIC;
    SIGNAL S1905 : STD_LOGIC;
    SIGNAL S1906 : STD_LOGIC;
    SIGNAL S1907 : STD_LOGIC;
    SIGNAL S1908 : STD_LOGIC;
    SIGNAL S1909 : STD_LOGIC;
    SIGNAL S1910 : STD_LOGIC;
    SIGNAL S1911 : STD_LOGIC;
    SIGNAL S1912 : STD_LOGIC;
    SIGNAL S1913 : STD_LOGIC;
    SIGNAL S1914 : STD_LOGIC;
    SIGNAL S1915 : STD_LOGIC;
    SIGNAL S1916 : STD_LOGIC;
    SIGNAL S1917 : STD_LOGIC;
    SIGNAL S1918 : STD_LOGIC;
    SIGNAL S1919 : STD_LOGIC;
    SIGNAL S1920 : STD_LOGIC;
    SIGNAL S1921 : STD_LOGIC;
    SIGNAL S1922 : STD_LOGIC;
    SIGNAL S1923 : STD_LOGIC;
    SIGNAL S1924 : STD_LOGIC;
    SIGNAL S1925 : STD_LOGIC;
    SIGNAL S1926 : STD_LOGIC;
    SIGNAL S1927 : STD_LOGIC;
    SIGNAL S1928 : STD_LOGIC;
    SIGNAL S1929 : STD_LOGIC;
    SIGNAL S1930 : STD_LOGIC;
    SIGNAL S1931 : STD_LOGIC;
    SIGNAL S1932 : STD_LOGIC;
    SIGNAL S1933 : STD_LOGIC;
    SIGNAL S1934 : STD_LOGIC;
    SIGNAL S1935 : STD_LOGIC;
    SIGNAL S1936 : STD_LOGIC;
    SIGNAL S1937 : STD_LOGIC;
    SIGNAL S1938 : STD_LOGIC;
    SIGNAL S1939 : STD_LOGIC;
    SIGNAL S1940 : STD_LOGIC;
    SIGNAL S1941 : STD_LOGIC;
    SIGNAL S1942 : STD_LOGIC;
    SIGNAL S1943 : STD_LOGIC;
    SIGNAL S1944 : STD_LOGIC;
    SIGNAL S1945 : STD_LOGIC;
    SIGNAL S1946 : STD_LOGIC;
    SIGNAL S1947 : STD_LOGIC;
    SIGNAL S1948 : STD_LOGIC;
    SIGNAL S1949 : STD_LOGIC;
    SIGNAL S1950 : STD_LOGIC;
    SIGNAL S1951 : STD_LOGIC;
    SIGNAL S1952 : STD_LOGIC;
    SIGNAL S1953 : STD_LOGIC;
    SIGNAL S1954 : STD_LOGIC;
    SIGNAL S1955 : STD_LOGIC;
    SIGNAL S1956 : STD_LOGIC;
    SIGNAL S1957 : STD_LOGIC;
    SIGNAL S1958 : STD_LOGIC;
    SIGNAL S1959 : STD_LOGIC;
    SIGNAL S1960 : STD_LOGIC;
    SIGNAL S1961 : STD_LOGIC;
    SIGNAL S1962 : STD_LOGIC;
    SIGNAL S1963 : STD_LOGIC;
    SIGNAL S1964 : STD_LOGIC;
    SIGNAL S1965 : STD_LOGIC;
    SIGNAL S1966 : STD_LOGIC;
    SIGNAL S1967 : STD_LOGIC;
    SIGNAL S1968 : STD_LOGIC;
    SIGNAL S1969 : STD_LOGIC;
    SIGNAL S1970 : STD_LOGIC;
    SIGNAL S1971 : STD_LOGIC;
    SIGNAL S1972 : STD_LOGIC;
    SIGNAL S1973 : STD_LOGIC;
    SIGNAL S1974 : STD_LOGIC;
    SIGNAL S1975 : STD_LOGIC;
    SIGNAL S1976 : STD_LOGIC;
    SIGNAL S1977 : STD_LOGIC;
    SIGNAL S1978 : STD_LOGIC;
    SIGNAL S1979 : STD_LOGIC;
    SIGNAL S1980 : STD_LOGIC;
    SIGNAL S1981 : STD_LOGIC;
    SIGNAL S1982 : STD_LOGIC;
    SIGNAL S1983 : STD_LOGIC;
    SIGNAL S1984 : STD_LOGIC;
    SIGNAL S1985 : STD_LOGIC;
    SIGNAL S1986 : STD_LOGIC;
    SIGNAL S1987 : STD_LOGIC;
    SIGNAL S1988 : STD_LOGIC;
    SIGNAL S1989 : STD_LOGIC;
    SIGNAL S1990 : STD_LOGIC;
    SIGNAL S1991 : STD_LOGIC;
    SIGNAL S1992 : STD_LOGIC;
    SIGNAL S1993 : STD_LOGIC;
    SIGNAL S1994 : STD_LOGIC;
    SIGNAL S1995 : STD_LOGIC;
    SIGNAL S1996 : STD_LOGIC;
    SIGNAL S1997 : STD_LOGIC;
    SIGNAL S1998 : STD_LOGIC;
    SIGNAL S1999 : STD_LOGIC;
    SIGNAL S2000 : STD_LOGIC;
    SIGNAL S2001 : STD_LOGIC;
    SIGNAL S2002 : STD_LOGIC;
    SIGNAL S2003 : STD_LOGIC;
    SIGNAL S2004 : STD_LOGIC;
    SIGNAL S2005 : STD_LOGIC;
    SIGNAL S2006 : STD_LOGIC;
    SIGNAL S2007 : STD_LOGIC;
    SIGNAL S2008 : STD_LOGIC;
    SIGNAL S2009 : STD_LOGIC;
    SIGNAL S2010 : STD_LOGIC;
    SIGNAL S2011 : STD_LOGIC;
    SIGNAL S2012 : STD_LOGIC;
    SIGNAL S2013 : STD_LOGIC;
    SIGNAL S2014 : STD_LOGIC;
    SIGNAL S2015 : STD_LOGIC;
    SIGNAL S2016 : STD_LOGIC;
    SIGNAL S2017 : STD_LOGIC;
    SIGNAL S2018 : STD_LOGIC;
    SIGNAL S2019 : STD_LOGIC;
    SIGNAL S2020 : STD_LOGIC;
    SIGNAL S2021 : STD_LOGIC;
    SIGNAL S2022 : STD_LOGIC;
    SIGNAL S2023 : STD_LOGIC;
    SIGNAL S2024 : STD_LOGIC;
    SIGNAL S2025 : STD_LOGIC;
    SIGNAL S2026 : STD_LOGIC;
    SIGNAL S2027 : STD_LOGIC;
    SIGNAL S2028 : STD_LOGIC;
    SIGNAL S2029 : STD_LOGIC;
    SIGNAL S2030 : STD_LOGIC;
    SIGNAL S2031 : STD_LOGIC;
    SIGNAL S2032 : STD_LOGIC;
    SIGNAL S2033 : STD_LOGIC;
    SIGNAL S2034 : STD_LOGIC;
    SIGNAL S2035 : STD_LOGIC;
    SIGNAL S2036 : STD_LOGIC;
    SIGNAL S2037 : STD_LOGIC;
    SIGNAL S2038 : STD_LOGIC;
    SIGNAL S2039 : STD_LOGIC;
    SIGNAL S2040 : STD_LOGIC;
    SIGNAL S2041 : STD_LOGIC;
    SIGNAL S2042 : STD_LOGIC;
    SIGNAL S2043 : STD_LOGIC;
    SIGNAL S2044 : STD_LOGIC;
    SIGNAL S2045 : STD_LOGIC;
    SIGNAL S2046 : STD_LOGIC;
    SIGNAL S2047 : STD_LOGIC;
    SIGNAL S2048 : STD_LOGIC;
    SIGNAL S2049 : STD_LOGIC;
    SIGNAL S2050 : STD_LOGIC;
    SIGNAL S2051 : STD_LOGIC;
    SIGNAL S2052 : STD_LOGIC;
    SIGNAL S2053 : STD_LOGIC;
    SIGNAL S2054 : STD_LOGIC;
    SIGNAL S2055 : STD_LOGIC;
    SIGNAL S2056 : STD_LOGIC;
    SIGNAL S2057 : STD_LOGIC;
    SIGNAL S2058 : STD_LOGIC;
    SIGNAL S2059 : STD_LOGIC;
    SIGNAL S2060 : STD_LOGIC;
    SIGNAL S2061 : STD_LOGIC;
    SIGNAL S2062 : STD_LOGIC;
    SIGNAL S2063 : STD_LOGIC;
    SIGNAL S2064 : STD_LOGIC;
    SIGNAL S2065 : STD_LOGIC;
    SIGNAL S2066 : STD_LOGIC;
    SIGNAL S2067 : STD_LOGIC;
    SIGNAL S2068 : STD_LOGIC;
    SIGNAL S2069 : STD_LOGIC;
    SIGNAL S2070 : STD_LOGIC;
    SIGNAL S2071 : STD_LOGIC;
    SIGNAL S2072 : STD_LOGIC;
    SIGNAL S2073 : STD_LOGIC;
    SIGNAL S2074 : STD_LOGIC;
    SIGNAL S2075 : STD_LOGIC;
    SIGNAL S2076 : STD_LOGIC;
    SIGNAL S2077 : STD_LOGIC;
    SIGNAL S2078 : STD_LOGIC;
    SIGNAL S2079 : STD_LOGIC;
    SIGNAL S2080 : STD_LOGIC;
    SIGNAL S2081 : STD_LOGIC;
    SIGNAL S2082 : STD_LOGIC;
    SIGNAL S2083 : STD_LOGIC;
    SIGNAL S2084 : STD_LOGIC;
    SIGNAL S2085 : STD_LOGIC;
    SIGNAL S2086 : STD_LOGIC;
    SIGNAL S2087 : STD_LOGIC;
    SIGNAL S2088 : STD_LOGIC;
    SIGNAL S2089 : STD_LOGIC;
    SIGNAL S2090 : STD_LOGIC;
    SIGNAL S2091 : STD_LOGIC;
    SIGNAL S2092 : STD_LOGIC;
    SIGNAL S2093 : STD_LOGIC;
    SIGNAL S2094 : STD_LOGIC;
    SIGNAL S2095 : STD_LOGIC;
    SIGNAL S2096 : STD_LOGIC;
    SIGNAL S2097 : STD_LOGIC;
    SIGNAL S2098 : STD_LOGIC;
    SIGNAL S2099 : STD_LOGIC;
    SIGNAL S2100 : STD_LOGIC;
    SIGNAL S2101 : STD_LOGIC;
    SIGNAL S2102 : STD_LOGIC;
    SIGNAL S2103 : STD_LOGIC;
    SIGNAL S2104 : STD_LOGIC;
    SIGNAL S2105 : STD_LOGIC;
    SIGNAL S2106 : STD_LOGIC;
    SIGNAL S2107 : STD_LOGIC;
    SIGNAL S2108 : STD_LOGIC;
    SIGNAL S2109 : STD_LOGIC;
    SIGNAL S2110 : STD_LOGIC;
    SIGNAL S2111 : STD_LOGIC;
    SIGNAL S2112 : STD_LOGIC;
    SIGNAL S2113 : STD_LOGIC;
    SIGNAL S2114 : STD_LOGIC;
    SIGNAL S2115 : STD_LOGIC;
    SIGNAL S2116 : STD_LOGIC;
    SIGNAL S2117 : STD_LOGIC;
    SIGNAL S2118 : STD_LOGIC;
    SIGNAL S2119 : STD_LOGIC;
    SIGNAL S2120 : STD_LOGIC;
    SIGNAL S2121 : STD_LOGIC;
    SIGNAL S2122 : STD_LOGIC;
    SIGNAL S2123 : STD_LOGIC;
    SIGNAL S2124 : STD_LOGIC;
    SIGNAL S2125 : STD_LOGIC;
    SIGNAL S2126 : STD_LOGIC;
    SIGNAL S2127 : STD_LOGIC;
    SIGNAL S2128 : STD_LOGIC;
    SIGNAL S2129 : STD_LOGIC;
    SIGNAL S2130 : STD_LOGIC;
    SIGNAL S2131 : STD_LOGIC;
    SIGNAL S2132 : STD_LOGIC;
    SIGNAL S2133 : STD_LOGIC;
    SIGNAL S2134 : STD_LOGIC;
    SIGNAL S2135 : STD_LOGIC;
    SIGNAL S2136 : STD_LOGIC;
    SIGNAL S2137 : STD_LOGIC;
    SIGNAL S2138 : STD_LOGIC;
    SIGNAL S2139 : STD_LOGIC;
    SIGNAL S2140 : STD_LOGIC;
    SIGNAL S2141 : STD_LOGIC;
    SIGNAL S2142 : STD_LOGIC;
    SIGNAL S2143 : STD_LOGIC;
    SIGNAL S2144 : STD_LOGIC;
    SIGNAL S2145 : STD_LOGIC;
    SIGNAL S2146 : STD_LOGIC;
    SIGNAL S2147 : STD_LOGIC;
    SIGNAL S2148 : STD_LOGIC;
    SIGNAL S2149 : STD_LOGIC;
    SIGNAL S2150 : STD_LOGIC;
    SIGNAL S2151 : STD_LOGIC;
    SIGNAL S2152 : STD_LOGIC;
    SIGNAL S2153 : STD_LOGIC;
    SIGNAL S2154 : STD_LOGIC;
    SIGNAL S2155 : STD_LOGIC;
    SIGNAL S2156 : STD_LOGIC;
    SIGNAL S2157 : STD_LOGIC;
    SIGNAL S2158 : STD_LOGIC;
    SIGNAL S2159 : STD_LOGIC;
    SIGNAL S2160 : STD_LOGIC;
    SIGNAL S2161 : STD_LOGIC;
    SIGNAL S2162 : STD_LOGIC;
    SIGNAL S2163 : STD_LOGIC;
    SIGNAL S2164 : STD_LOGIC;
    SIGNAL S2165 : STD_LOGIC;
    SIGNAL S2166 : STD_LOGIC;
    SIGNAL S2167 : STD_LOGIC;
    SIGNAL S2168 : STD_LOGIC;
    SIGNAL S2169 : STD_LOGIC;
    SIGNAL S2170 : STD_LOGIC;
    SIGNAL S2171 : STD_LOGIC;
    SIGNAL S2172 : STD_LOGIC;
    SIGNAL S2173 : STD_LOGIC;
    SIGNAL S2174 : STD_LOGIC;
    SIGNAL S2175 : STD_LOGIC;
    SIGNAL S2176 : STD_LOGIC;
    SIGNAL S2177 : STD_LOGIC;
    SIGNAL S2178 : STD_LOGIC;
    SIGNAL S2179 : STD_LOGIC;
    SIGNAL S2180 : STD_LOGIC;
    SIGNAL S2181 : STD_LOGIC;
    SIGNAL S2182 : STD_LOGIC;
    SIGNAL S2183 : STD_LOGIC;
    SIGNAL S2184 : STD_LOGIC;
    SIGNAL S2185 : STD_LOGIC;
    SIGNAL S2186 : STD_LOGIC;
    SIGNAL S2187 : STD_LOGIC;
    SIGNAL S2188 : STD_LOGIC;
    SIGNAL S2189 : STD_LOGIC;
    SIGNAL S2190 : STD_LOGIC;
    SIGNAL S2191 : STD_LOGIC;
    SIGNAL S2192 : STD_LOGIC;
    SIGNAL S2193 : STD_LOGIC;
    SIGNAL S2194 : STD_LOGIC;
    SIGNAL S2195 : STD_LOGIC;
    SIGNAL S2196 : STD_LOGIC;
    SIGNAL S2197 : STD_LOGIC;
    SIGNAL S2198 : STD_LOGIC;
    SIGNAL S2199 : STD_LOGIC;
    SIGNAL S2200 : STD_LOGIC;
    SIGNAL S2201 : STD_LOGIC;
    SIGNAL S2202 : STD_LOGIC;
    SIGNAL S2203 : STD_LOGIC;
    SIGNAL S2204 : STD_LOGIC;
    SIGNAL S2205 : STD_LOGIC;
    SIGNAL S2206 : STD_LOGIC;
    SIGNAL S2207 : STD_LOGIC;
    SIGNAL S2208 : STD_LOGIC;
    SIGNAL S2209 : STD_LOGIC;
    SIGNAL S2210 : STD_LOGIC;
    SIGNAL S2211 : STD_LOGIC;
    SIGNAL S2212 : STD_LOGIC;
    SIGNAL S2213 : STD_LOGIC;
    SIGNAL S2214 : STD_LOGIC;
    SIGNAL S2215 : STD_LOGIC;
    SIGNAL S2216 : STD_LOGIC;
    SIGNAL S2217 : STD_LOGIC;
    SIGNAL S2218 : STD_LOGIC;
    SIGNAL S2219 : STD_LOGIC;
    SIGNAL S2220 : STD_LOGIC;
    SIGNAL S2221 : STD_LOGIC;
    SIGNAL S2222 : STD_LOGIC;
    SIGNAL S2223 : STD_LOGIC;
    SIGNAL S2224 : STD_LOGIC;
    SIGNAL S2225 : STD_LOGIC;
    SIGNAL S2226 : STD_LOGIC;
    SIGNAL S2227 : STD_LOGIC;
    SIGNAL S2228 : STD_LOGIC;
    SIGNAL S2229 : STD_LOGIC;
    SIGNAL S2230 : STD_LOGIC;
    SIGNAL S2231 : STD_LOGIC;
    SIGNAL S2232 : STD_LOGIC;
    SIGNAL S2233 : STD_LOGIC;
    SIGNAL S2234 : STD_LOGIC;
    SIGNAL S2235 : STD_LOGIC;
    SIGNAL S2236 : STD_LOGIC;
    SIGNAL S2237 : STD_LOGIC;
    SIGNAL S2238 : STD_LOGIC;
    SIGNAL S2239 : STD_LOGIC;
    SIGNAL S2240 : STD_LOGIC;
    SIGNAL S2241 : STD_LOGIC;
    SIGNAL S2242 : STD_LOGIC;
    SIGNAL S2243 : STD_LOGIC;
    SIGNAL S2244 : STD_LOGIC;
    SIGNAL S2245 : STD_LOGIC;
    SIGNAL S2246 : STD_LOGIC;
    SIGNAL S2247 : STD_LOGIC;
    SIGNAL S2248 : STD_LOGIC;
    SIGNAL S2249 : STD_LOGIC;
    SIGNAL S2250 : STD_LOGIC;
    SIGNAL S2251 : STD_LOGIC;
    SIGNAL S2252 : STD_LOGIC;
    SIGNAL S2253 : STD_LOGIC;
    SIGNAL S2254 : STD_LOGIC;
    SIGNAL S2255 : STD_LOGIC;
    SIGNAL S2256 : STD_LOGIC;
    SIGNAL S2257 : STD_LOGIC;
    SIGNAL S2258 : STD_LOGIC;
    SIGNAL S2259 : STD_LOGIC;
    SIGNAL S2260 : STD_LOGIC;
    SIGNAL S2261 : STD_LOGIC;
    SIGNAL S2262 : STD_LOGIC;
    SIGNAL S2263 : STD_LOGIC;
    SIGNAL S2264 : STD_LOGIC;
    SIGNAL S2265 : STD_LOGIC;
    SIGNAL S2266 : STD_LOGIC;
    SIGNAL S2267 : STD_LOGIC;
    SIGNAL S2268 : STD_LOGIC;
    SIGNAL S2269 : STD_LOGIC;
    SIGNAL S2270 : STD_LOGIC;
    SIGNAL S2271 : STD_LOGIC;
    SIGNAL S2272 : STD_LOGIC;
    SIGNAL S2273 : STD_LOGIC;
    SIGNAL S2274 : STD_LOGIC;
    SIGNAL S2275 : STD_LOGIC;
    SIGNAL S2276 : STD_LOGIC;
    SIGNAL S2277 : STD_LOGIC;
    SIGNAL S2278 : STD_LOGIC;
    SIGNAL S2279 : STD_LOGIC;
    SIGNAL S2280 : STD_LOGIC;
    SIGNAL S2281 : STD_LOGIC;
    SIGNAL S2282 : STD_LOGIC;
    SIGNAL S2283 : STD_LOGIC;
    SIGNAL S2284 : STD_LOGIC;
    SIGNAL S2285 : STD_LOGIC;
    SIGNAL S2286 : STD_LOGIC;
    SIGNAL S2287 : STD_LOGIC;
    SIGNAL S2288 : STD_LOGIC;
    SIGNAL S2289 : STD_LOGIC;
    SIGNAL S2290 : STD_LOGIC;
    SIGNAL S2291 : STD_LOGIC;
    SIGNAL S2292 : STD_LOGIC;
    SIGNAL S2293 : STD_LOGIC;
    SIGNAL S2294 : STD_LOGIC;
    SIGNAL S2295 : STD_LOGIC;
    SIGNAL S2296 : STD_LOGIC;
    SIGNAL S2297 : STD_LOGIC;
    SIGNAL S2298 : STD_LOGIC;
    SIGNAL S2299 : STD_LOGIC;
    SIGNAL S2300 : STD_LOGIC;
    SIGNAL S2301 : STD_LOGIC;
    SIGNAL S2302 : STD_LOGIC;
    SIGNAL S2303 : STD_LOGIC;
    SIGNAL S2304 : STD_LOGIC;
    SIGNAL S2305 : STD_LOGIC;
    SIGNAL S2306 : STD_LOGIC;
    SIGNAL S2307 : STD_LOGIC;
    SIGNAL S2308 : STD_LOGIC;
    SIGNAL S2309 : STD_LOGIC;
    SIGNAL S2310 : STD_LOGIC;
    SIGNAL S2311 : STD_LOGIC;
    SIGNAL S2312 : STD_LOGIC;
    SIGNAL S2313 : STD_LOGIC;
    SIGNAL S2314 : STD_LOGIC;
    SIGNAL S2315 : STD_LOGIC;
    SIGNAL S2316 : STD_LOGIC;
    SIGNAL S2317 : STD_LOGIC;
    SIGNAL S2318 : STD_LOGIC;
    SIGNAL S2319 : STD_LOGIC;
    SIGNAL S2320 : STD_LOGIC;
    SIGNAL S2321 : STD_LOGIC;
    SIGNAL S2322 : STD_LOGIC;
    SIGNAL S2323 : STD_LOGIC;
    SIGNAL S2324 : STD_LOGIC;
    SIGNAL S2325 : STD_LOGIC;
    SIGNAL S2326 : STD_LOGIC;
    SIGNAL S2327 : STD_LOGIC;
    SIGNAL S2328 : STD_LOGIC;
    SIGNAL S2329 : STD_LOGIC;
    SIGNAL S2330 : STD_LOGIC;
    SIGNAL S2331 : STD_LOGIC;
    SIGNAL S2332 : STD_LOGIC;
    SIGNAL S2333 : STD_LOGIC;
    SIGNAL S2334 : STD_LOGIC;
    SIGNAL S2335 : STD_LOGIC;
    SIGNAL S2336 : STD_LOGIC;
    SIGNAL S2337 : STD_LOGIC;
    SIGNAL S2338 : STD_LOGIC;
    SIGNAL S2339 : STD_LOGIC;
    SIGNAL S2340 : STD_LOGIC;
    SIGNAL S2341 : STD_LOGIC;
    SIGNAL S2342 : STD_LOGIC;
    SIGNAL S2343 : STD_LOGIC;
    SIGNAL S2344 : STD_LOGIC;
    SIGNAL S2345 : STD_LOGIC;
    SIGNAL S2346 : STD_LOGIC;
    SIGNAL S2347 : STD_LOGIC;
    SIGNAL S2348 : STD_LOGIC;
    SIGNAL S2349 : STD_LOGIC;
    SIGNAL S2350 : STD_LOGIC;
    SIGNAL S2351 : STD_LOGIC;
    SIGNAL S2352 : STD_LOGIC;
    SIGNAL S2353 : STD_LOGIC;
    SIGNAL S2354 : STD_LOGIC;
    SIGNAL S2355 : STD_LOGIC;
    SIGNAL S2356 : STD_LOGIC;
    SIGNAL S2357 : STD_LOGIC;
    SIGNAL S2358 : STD_LOGIC;
    SIGNAL S2359 : STD_LOGIC;
    SIGNAL S2360 : STD_LOGIC;
    SIGNAL S2361 : STD_LOGIC;
    SIGNAL S2362 : STD_LOGIC;
    SIGNAL S2363 : STD_LOGIC;
    SIGNAL S2364 : STD_LOGIC;
    SIGNAL S2365 : STD_LOGIC;
    SIGNAL S2366 : STD_LOGIC;
    SIGNAL S2367 : STD_LOGIC;
    SIGNAL S2368 : STD_LOGIC;
    SIGNAL S2369 : STD_LOGIC;
    SIGNAL S2370 : STD_LOGIC;
    SIGNAL S2371 : STD_LOGIC;
    SIGNAL S2372 : STD_LOGIC;
    SIGNAL S2373 : STD_LOGIC;
    SIGNAL S2374 : STD_LOGIC;
    SIGNAL S2375 : STD_LOGIC;
    SIGNAL S2376 : STD_LOGIC;
    SIGNAL S2377 : STD_LOGIC;
    SIGNAL S2378 : STD_LOGIC;
    SIGNAL S2379 : STD_LOGIC;
    SIGNAL S2380 : STD_LOGIC;
    SIGNAL S2381 : STD_LOGIC;
    SIGNAL S2382 : STD_LOGIC;
    SIGNAL S2383 : STD_LOGIC;
    SIGNAL S2384 : STD_LOGIC;
    SIGNAL S2385 : STD_LOGIC;
    SIGNAL S2386 : STD_LOGIC;
    SIGNAL S2387 : STD_LOGIC;
    SIGNAL S2388 : STD_LOGIC;
    SIGNAL S2389 : STD_LOGIC;
    SIGNAL S2390 : STD_LOGIC;
    SIGNAL S2391 : STD_LOGIC;
    SIGNAL S2392 : STD_LOGIC;
    SIGNAL S2393 : STD_LOGIC;
    SIGNAL S2394 : STD_LOGIC;
    SIGNAL S2395 : STD_LOGIC;
    SIGNAL S2396 : STD_LOGIC;
    SIGNAL S2397 : STD_LOGIC;
    SIGNAL S2398 : STD_LOGIC;
    SIGNAL S2399 : STD_LOGIC;
    SIGNAL S2400 : STD_LOGIC;
    SIGNAL S2401 : STD_LOGIC;
    SIGNAL S2402 : STD_LOGIC;
    SIGNAL S2403 : STD_LOGIC;
    SIGNAL S2404 : STD_LOGIC;
    SIGNAL S2405 : STD_LOGIC;
    SIGNAL S2406 : STD_LOGIC;
    SIGNAL S2407 : STD_LOGIC;
    SIGNAL S2408 : STD_LOGIC;
    SIGNAL S2409 : STD_LOGIC;
    SIGNAL S2410 : STD_LOGIC;
    SIGNAL S2411 : STD_LOGIC;
    SIGNAL S2412 : STD_LOGIC;
    SIGNAL S2413 : STD_LOGIC;
    SIGNAL S2414 : STD_LOGIC;
    SIGNAL S2415 : STD_LOGIC;
    SIGNAL S2416 : STD_LOGIC;
    SIGNAL S2417 : STD_LOGIC;
    SIGNAL S2418 : STD_LOGIC;
    SIGNAL S2419 : STD_LOGIC;
    SIGNAL S2420 : STD_LOGIC;
    SIGNAL S2421 : STD_LOGIC;
    SIGNAL S2422 : STD_LOGIC;
    SIGNAL S2423 : STD_LOGIC;
    SIGNAL S2424 : STD_LOGIC;
    SIGNAL S2425 : STD_LOGIC;
    SIGNAL S2426 : STD_LOGIC;
    SIGNAL S2427 : STD_LOGIC;
    SIGNAL S2428 : STD_LOGIC;
    SIGNAL S2429 : STD_LOGIC;
    SIGNAL S2430 : STD_LOGIC;
    SIGNAL S2431 : STD_LOGIC;
    SIGNAL S2432 : STD_LOGIC;
    SIGNAL S2433 : STD_LOGIC;
    SIGNAL S2434 : STD_LOGIC;
    SIGNAL S2435 : STD_LOGIC;
    SIGNAL S2436 : STD_LOGIC;
    SIGNAL S2437 : STD_LOGIC;
    SIGNAL S2438 : STD_LOGIC;
    SIGNAL S2439 : STD_LOGIC;
    SIGNAL S2440 : STD_LOGIC;
    SIGNAL S2441 : STD_LOGIC;
    SIGNAL S2442 : STD_LOGIC;
    SIGNAL S2443 : STD_LOGIC;
    SIGNAL S2444 : STD_LOGIC;
    SIGNAL S2445 : STD_LOGIC;
    SIGNAL S2446 : STD_LOGIC;
    SIGNAL S2447 : STD_LOGIC;
    SIGNAL S2448 : STD_LOGIC;
    SIGNAL S2449 : STD_LOGIC;
    SIGNAL S2450 : STD_LOGIC;
    SIGNAL S2451 : STD_LOGIC;
    SIGNAL S2452 : STD_LOGIC;
    SIGNAL S2453 : STD_LOGIC;
    SIGNAL S2454 : STD_LOGIC;
    SIGNAL S2455 : STD_LOGIC;
    SIGNAL S2456 : STD_LOGIC;
    SIGNAL S2457 : STD_LOGIC;
    SIGNAL S2458 : STD_LOGIC;
    SIGNAL S2459 : STD_LOGIC;
    SIGNAL S2460 : STD_LOGIC;
    SIGNAL S2461 : STD_LOGIC;
    SIGNAL S2462 : STD_LOGIC;
    SIGNAL S2463 : STD_LOGIC;
    SIGNAL S2464 : STD_LOGIC;
    SIGNAL S2465 : STD_LOGIC;
    SIGNAL S2466 : STD_LOGIC;
    SIGNAL S2467 : STD_LOGIC;
    SIGNAL S2468 : STD_LOGIC;
    SIGNAL S2469 : STD_LOGIC;
    SIGNAL S2470 : STD_LOGIC;
    SIGNAL S2471 : STD_LOGIC;
    SIGNAL S2472 : STD_LOGIC;
    SIGNAL S2473 : STD_LOGIC;
    SIGNAL S2474 : STD_LOGIC;
    SIGNAL S2475 : STD_LOGIC;
    SIGNAL S2476 : STD_LOGIC;
    SIGNAL S2477 : STD_LOGIC;
    SIGNAL S2478 : STD_LOGIC;
    SIGNAL S2479 : STD_LOGIC;
    SIGNAL S2480 : STD_LOGIC;
    SIGNAL S2481 : STD_LOGIC;
    SIGNAL S2482 : STD_LOGIC;
    SIGNAL S2483 : STD_LOGIC;
    SIGNAL S2484 : STD_LOGIC;
    SIGNAL S2485 : STD_LOGIC;
    SIGNAL S2486 : STD_LOGIC;
    SIGNAL S2487 : STD_LOGIC;
    SIGNAL S2488 : STD_LOGIC;
    SIGNAL S2489 : STD_LOGIC;
    SIGNAL S2490 : STD_LOGIC;
    SIGNAL S2491 : STD_LOGIC;
    SIGNAL S2492 : STD_LOGIC;
    SIGNAL S2493 : STD_LOGIC;
    SIGNAL S2494 : STD_LOGIC;
    SIGNAL S2495 : STD_LOGIC;
    SIGNAL S2496 : STD_LOGIC;
    SIGNAL S2497 : STD_LOGIC;
    SIGNAL S2498 : STD_LOGIC;
    SIGNAL S2499 : STD_LOGIC;
    SIGNAL S2500 : STD_LOGIC;
    SIGNAL S2501 : STD_LOGIC;
    SIGNAL S2502 : STD_LOGIC;
    SIGNAL S2503 : STD_LOGIC;
    SIGNAL S2504 : STD_LOGIC;
    SIGNAL S2505 : STD_LOGIC;
    SIGNAL S2506 : STD_LOGIC;
    SIGNAL S2507 : STD_LOGIC;
    SIGNAL S2508 : STD_LOGIC;
    SIGNAL S2509 : STD_LOGIC;
    SIGNAL S2510 : STD_LOGIC;
    SIGNAL S2511 : STD_LOGIC;
    SIGNAL S2512 : STD_LOGIC;
    SIGNAL S2513 : STD_LOGIC;
    SIGNAL S2514 : STD_LOGIC;
    SIGNAL S2515 : STD_LOGIC;
    SIGNAL S2516 : STD_LOGIC;
    SIGNAL S2517 : STD_LOGIC;
    SIGNAL S2518 : STD_LOGIC;
    SIGNAL S2519 : STD_LOGIC;
    SIGNAL S2520 : STD_LOGIC;
    SIGNAL S2521 : STD_LOGIC;
    SIGNAL S2522 : STD_LOGIC;
    SIGNAL S2523 : STD_LOGIC;
    SIGNAL S2524 : STD_LOGIC;
    SIGNAL S2525 : STD_LOGIC;
    SIGNAL S2526 : STD_LOGIC;
    SIGNAL S2527 : STD_LOGIC;
    SIGNAL S2528 : STD_LOGIC;
    SIGNAL S2529 : STD_LOGIC;
    SIGNAL S2530 : STD_LOGIC;
    SIGNAL S2531 : STD_LOGIC;
    SIGNAL S2532 : STD_LOGIC;
    SIGNAL S2533 : STD_LOGIC;
    SIGNAL S2534 : STD_LOGIC;
    SIGNAL S2535 : STD_LOGIC;
    SIGNAL S2536 : STD_LOGIC;
    SIGNAL S2537 : STD_LOGIC;
    SIGNAL S2538 : STD_LOGIC;
    SIGNAL S2539 : STD_LOGIC;
    SIGNAL S2540 : STD_LOGIC;
    SIGNAL S2541 : STD_LOGIC;
    SIGNAL S2542 : STD_LOGIC;
    SIGNAL S2543 : STD_LOGIC;
    SIGNAL S2544 : STD_LOGIC;
    SIGNAL S2545 : STD_LOGIC;
    SIGNAL S2546 : STD_LOGIC;
    SIGNAL S2547 : STD_LOGIC;
    SIGNAL S2548 : STD_LOGIC;
    SIGNAL S2549 : STD_LOGIC;
    SIGNAL S2550 : STD_LOGIC;
    SIGNAL S2551 : STD_LOGIC;
    SIGNAL S2552 : STD_LOGIC;
    SIGNAL S2553 : STD_LOGIC;
    SIGNAL S2554 : STD_LOGIC;
    SIGNAL S2555 : STD_LOGIC;
    SIGNAL S2556 : STD_LOGIC;
    SIGNAL S2557 : STD_LOGIC;
    SIGNAL S2558 : STD_LOGIC;
    SIGNAL S2559 : STD_LOGIC;
    SIGNAL S2560 : STD_LOGIC;
    SIGNAL S2561 : STD_LOGIC;
    SIGNAL S2562 : STD_LOGIC;
    SIGNAL S2563 : STD_LOGIC;
    SIGNAL S2564 : STD_LOGIC;
    SIGNAL S2565 : STD_LOGIC;
    SIGNAL S2566 : STD_LOGIC;
    SIGNAL S2567 : STD_LOGIC;
    SIGNAL S2568 : STD_LOGIC;
    SIGNAL S2569 : STD_LOGIC;
    SIGNAL S2570 : STD_LOGIC;
    SIGNAL S2571 : STD_LOGIC;
    SIGNAL S2572 : STD_LOGIC;
    SIGNAL S2573 : STD_LOGIC;
    SIGNAL S2574 : STD_LOGIC;
    SIGNAL S2575 : STD_LOGIC;
    SIGNAL S2576 : STD_LOGIC;
    SIGNAL S2577 : STD_LOGIC;
    SIGNAL S2578 : STD_LOGIC;
    SIGNAL S2579 : STD_LOGIC;
    SIGNAL S2580 : STD_LOGIC;
    SIGNAL S2581 : STD_LOGIC;
    SIGNAL S2582 : STD_LOGIC;
    SIGNAL S2583 : STD_LOGIC;
    SIGNAL S2584 : STD_LOGIC;
    SIGNAL S2585 : STD_LOGIC;
    SIGNAL S2586 : STD_LOGIC;
    SIGNAL S2587 : STD_LOGIC;
    SIGNAL S2588 : STD_LOGIC;
    SIGNAL S2589 : STD_LOGIC;
    SIGNAL S2590 : STD_LOGIC;
    SIGNAL S2591 : STD_LOGIC;
    SIGNAL S2592 : STD_LOGIC;
    SIGNAL S2593 : STD_LOGIC;
    SIGNAL S2594 : STD_LOGIC;
    SIGNAL S2595 : STD_LOGIC;
    SIGNAL S2596 : STD_LOGIC;
    SIGNAL S2597 : STD_LOGIC;
    SIGNAL S2598 : STD_LOGIC;
    SIGNAL S2599 : STD_LOGIC;
    SIGNAL S2600 : STD_LOGIC;
    SIGNAL S2601 : STD_LOGIC;
    SIGNAL S2602 : STD_LOGIC;
    SIGNAL S2603 : STD_LOGIC;
    SIGNAL S2604 : STD_LOGIC;
    SIGNAL S2605 : STD_LOGIC;
    SIGNAL S2606 : STD_LOGIC;
    SIGNAL S2607 : STD_LOGIC;
    SIGNAL S2608 : STD_LOGIC;
    SIGNAL S2609 : STD_LOGIC;
    SIGNAL S2610 : STD_LOGIC;
    SIGNAL S2611 : STD_LOGIC;
    SIGNAL S2612 : STD_LOGIC;
    SIGNAL S2613 : STD_LOGIC;
    SIGNAL S2614 : STD_LOGIC;
    SIGNAL S2615 : STD_LOGIC;
    SIGNAL S2616 : STD_LOGIC;
    SIGNAL S2617 : STD_LOGIC;
    SIGNAL S2618 : STD_LOGIC;
    SIGNAL S2619 : STD_LOGIC;
    SIGNAL S2620 : STD_LOGIC;
    SIGNAL S2621 : STD_LOGIC;
    SIGNAL S2622 : STD_LOGIC;
    SIGNAL S2623 : STD_LOGIC;
    SIGNAL S2624 : STD_LOGIC;
    SIGNAL S2625 : STD_LOGIC;
    SIGNAL S2626 : STD_LOGIC;
    SIGNAL S2627 : STD_LOGIC;
    SIGNAL S2628 : STD_LOGIC;
    SIGNAL S2629 : STD_LOGIC;
    SIGNAL S2630 : STD_LOGIC;
    SIGNAL S2631 : STD_LOGIC;
    SIGNAL S2632 : STD_LOGIC;
    SIGNAL S2633 : STD_LOGIC;
    SIGNAL S2634 : STD_LOGIC;
    SIGNAL S2635 : STD_LOGIC;
    SIGNAL S2636 : STD_LOGIC;
    SIGNAL S2637 : STD_LOGIC;
    SIGNAL S2638 : STD_LOGIC;
    SIGNAL S2639 : STD_LOGIC;
    SIGNAL S2640 : STD_LOGIC;
    SIGNAL S2641 : STD_LOGIC;
    SIGNAL S2642 : STD_LOGIC;
    SIGNAL S2643 : STD_LOGIC;
    SIGNAL S2644 : STD_LOGIC;
    SIGNAL S2645 : STD_LOGIC;
    SIGNAL S2646 : STD_LOGIC;
    SIGNAL S2647 : STD_LOGIC;
    SIGNAL S2648 : STD_LOGIC;
    SIGNAL S2649 : STD_LOGIC;
    SIGNAL S2650 : STD_LOGIC;
    SIGNAL S2651 : STD_LOGIC;
    SIGNAL S2652 : STD_LOGIC;
    SIGNAL S2653 : STD_LOGIC;
    SIGNAL S2654 : STD_LOGIC;
    SIGNAL S2655 : STD_LOGIC;
    SIGNAL S2656 : STD_LOGIC;
    SIGNAL S2657 : STD_LOGIC;
    SIGNAL S2658 : STD_LOGIC;
    SIGNAL S2659 : STD_LOGIC;
    SIGNAL S2660 : STD_LOGIC;
    SIGNAL S2661 : STD_LOGIC;
    SIGNAL S2662 : STD_LOGIC;
    SIGNAL S2663 : STD_LOGIC;
    SIGNAL S2664 : STD_LOGIC;
    SIGNAL S2665 : STD_LOGIC;
    SIGNAL S2666 : STD_LOGIC;
    SIGNAL S2667 : STD_LOGIC;
    SIGNAL S2668 : STD_LOGIC;
    SIGNAL S2669 : STD_LOGIC;
    SIGNAL S2670 : STD_LOGIC;
    SIGNAL S2671 : STD_LOGIC;
    SIGNAL S2672 : STD_LOGIC;
    SIGNAL S2673 : STD_LOGIC;
    SIGNAL S2674 : STD_LOGIC;
    SIGNAL S2675 : STD_LOGIC;
    SIGNAL S2676 : STD_LOGIC;
    SIGNAL S2677 : STD_LOGIC;
    SIGNAL S2678 : STD_LOGIC;
    SIGNAL S2679 : STD_LOGIC;
    SIGNAL S2680 : STD_LOGIC;
    SIGNAL S2681 : STD_LOGIC;
    SIGNAL S2682 : STD_LOGIC;
    SIGNAL S2683 : STD_LOGIC;
    SIGNAL S2684 : STD_LOGIC;
    SIGNAL S2685 : STD_LOGIC;
    SIGNAL S2686 : STD_LOGIC;
    SIGNAL S2687 : STD_LOGIC;
    SIGNAL S2688 : STD_LOGIC;
    SIGNAL S2689 : STD_LOGIC;
    SIGNAL S2690 : STD_LOGIC;
    SIGNAL S2691 : STD_LOGIC;
    SIGNAL S2692 : STD_LOGIC;
    SIGNAL S2693 : STD_LOGIC;
    SIGNAL S2694 : STD_LOGIC;
    SIGNAL S2695 : STD_LOGIC;
    SIGNAL S2696 : STD_LOGIC;
    SIGNAL S2697 : STD_LOGIC;
    SIGNAL S2698 : STD_LOGIC;
    SIGNAL S2699 : STD_LOGIC;
    SIGNAL S2700 : STD_LOGIC;
    SIGNAL S2701 : STD_LOGIC;
    SIGNAL S2702 : STD_LOGIC;
    SIGNAL S2703 : STD_LOGIC;
    SIGNAL S2704 : STD_LOGIC;
    SIGNAL S2705 : STD_LOGIC;
    SIGNAL S2706 : STD_LOGIC;
    SIGNAL S2707 : STD_LOGIC;
    SIGNAL S2708 : STD_LOGIC;
    SIGNAL S2709 : STD_LOGIC;
    SIGNAL S2710 : STD_LOGIC;
    SIGNAL S2711 : STD_LOGIC;
    SIGNAL S2712 : STD_LOGIC;
    SIGNAL S2713 : STD_LOGIC;
    SIGNAL S2714 : STD_LOGIC;
    SIGNAL S2715 : STD_LOGIC;
    SIGNAL S2716 : STD_LOGIC;
    SIGNAL S2717 : STD_LOGIC;
    SIGNAL S2718 : STD_LOGIC;
    SIGNAL S2719 : STD_LOGIC;
    SIGNAL S2720 : STD_LOGIC;
    SIGNAL S2721 : STD_LOGIC;
    SIGNAL S2722 : STD_LOGIC;
    SIGNAL S2723 : STD_LOGIC;
    SIGNAL S2724 : STD_LOGIC;
    SIGNAL S2725 : STD_LOGIC;
    SIGNAL S2726 : STD_LOGIC;
    SIGNAL S2727 : STD_LOGIC;
    SIGNAL S2728 : STD_LOGIC;
    SIGNAL S2729 : STD_LOGIC;
    SIGNAL S2730 : STD_LOGIC;
    SIGNAL S2731 : STD_LOGIC;
    SIGNAL S2732 : STD_LOGIC;
    SIGNAL S2733 : STD_LOGIC;
    SIGNAL S2734 : STD_LOGIC;
    SIGNAL S2735 : STD_LOGIC;
    SIGNAL S2736 : STD_LOGIC;
    SIGNAL S2737 : STD_LOGIC;
    SIGNAL S2738 : STD_LOGIC;
    SIGNAL S2739 : STD_LOGIC;
    SIGNAL S2740 : STD_LOGIC;
    SIGNAL S2741 : STD_LOGIC;
    SIGNAL S2742 : STD_LOGIC;
    SIGNAL S2743 : STD_LOGIC;
    SIGNAL S2744 : STD_LOGIC;
    SIGNAL S2745 : STD_LOGIC;
    SIGNAL S2746 : STD_LOGIC;
    SIGNAL S2747 : STD_LOGIC;
    SIGNAL S2748 : STD_LOGIC;
    SIGNAL S2749 : STD_LOGIC;
    SIGNAL S2750 : STD_LOGIC;
    SIGNAL S2751 : STD_LOGIC;
    SIGNAL S2752 : STD_LOGIC;
    SIGNAL S2753 : STD_LOGIC;
    SIGNAL S2754 : STD_LOGIC;
    SIGNAL S2755 : STD_LOGIC;
    SIGNAL S2756 : STD_LOGIC;
    SIGNAL S2757 : STD_LOGIC;
    SIGNAL S2758 : STD_LOGIC;
    SIGNAL S2759 : STD_LOGIC;
    SIGNAL S2760 : STD_LOGIC;
    SIGNAL S2761 : STD_LOGIC;
    SIGNAL S2762 : STD_LOGIC;
    SIGNAL S2763 : STD_LOGIC;
    SIGNAL S2764 : STD_LOGIC;
    SIGNAL S2765 : STD_LOGIC;
    SIGNAL S2766 : STD_LOGIC;
    SIGNAL S2767 : STD_LOGIC;
    SIGNAL S2768 : STD_LOGIC;
    SIGNAL S2769 : STD_LOGIC;
    SIGNAL S2770 : STD_LOGIC;
    SIGNAL S2771 : STD_LOGIC;
    SIGNAL S2772 : STD_LOGIC;
    SIGNAL S2773 : STD_LOGIC;
    SIGNAL S2774 : STD_LOGIC;
    SIGNAL S2775 : STD_LOGIC;
    SIGNAL S2776 : STD_LOGIC;
    SIGNAL S2777 : STD_LOGIC;
    SIGNAL S2778 : STD_LOGIC;
    SIGNAL S2779 : STD_LOGIC;
    SIGNAL S2780 : STD_LOGIC;
    SIGNAL S2781 : STD_LOGIC;
    SIGNAL S2782 : STD_LOGIC;
    SIGNAL S2783 : STD_LOGIC;
    SIGNAL S2784 : STD_LOGIC;
    SIGNAL S2785 : STD_LOGIC;
    SIGNAL S2786 : STD_LOGIC;
    SIGNAL S2787 : STD_LOGIC;
    SIGNAL S2788 : STD_LOGIC;
    SIGNAL S2789 : STD_LOGIC;
    SIGNAL S2790 : STD_LOGIC;
    SIGNAL S2791 : STD_LOGIC;
    SIGNAL S2792 : STD_LOGIC;
    SIGNAL S2793 : STD_LOGIC;
    SIGNAL S2794 : STD_LOGIC;
    SIGNAL S2795 : STD_LOGIC;
    SIGNAL S2796 : STD_LOGIC;
    SIGNAL S2797 : STD_LOGIC;
    SIGNAL S2798 : STD_LOGIC;
    SIGNAL S2799 : STD_LOGIC;
    SIGNAL S2800 : STD_LOGIC;
    SIGNAL S2801 : STD_LOGIC;
    SIGNAL S2802 : STD_LOGIC;
    SIGNAL S2803 : STD_LOGIC;
    SIGNAL S2804 : STD_LOGIC;
    SIGNAL S2805 : STD_LOGIC;
    SIGNAL S2806 : STD_LOGIC;
    SIGNAL S2807 : STD_LOGIC;
    SIGNAL S2808 : STD_LOGIC;
    SIGNAL S2809 : STD_LOGIC;
    SIGNAL S2810 : STD_LOGIC;
    SIGNAL S2811 : STD_LOGIC;
    SIGNAL S2812 : STD_LOGIC;
    SIGNAL S2813 : STD_LOGIC;
    SIGNAL S2814 : STD_LOGIC;
    SIGNAL S2815 : STD_LOGIC;
    SIGNAL S2816 : STD_LOGIC;
    SIGNAL S2817 : STD_LOGIC;
    SIGNAL S2818 : STD_LOGIC;
    SIGNAL S2819 : STD_LOGIC;
    SIGNAL S2820 : STD_LOGIC;
    SIGNAL S2821 : STD_LOGIC;
    SIGNAL S2822 : STD_LOGIC;
    SIGNAL S2823 : STD_LOGIC;
    SIGNAL S2824 : STD_LOGIC;
    SIGNAL S2825 : STD_LOGIC;
    SIGNAL S2826 : STD_LOGIC;
    SIGNAL S2827 : STD_LOGIC;
    SIGNAL S2828 : STD_LOGIC;
    SIGNAL S2829 : STD_LOGIC;
    SIGNAL S2830 : STD_LOGIC;
    SIGNAL S2831 : STD_LOGIC;
    SIGNAL S2832 : STD_LOGIC;
    SIGNAL S2833 : STD_LOGIC;
    SIGNAL S2834 : STD_LOGIC;
    SIGNAL S2835 : STD_LOGIC;
    SIGNAL S2836 : STD_LOGIC;
    SIGNAL S2837 : STD_LOGIC;
    SIGNAL S2838 : STD_LOGIC;
    SIGNAL S2839 : STD_LOGIC;
    SIGNAL S2840 : STD_LOGIC;
    SIGNAL S2841 : STD_LOGIC;
    SIGNAL S2842 : STD_LOGIC;
    SIGNAL S2843 : STD_LOGIC;
    SIGNAL S2844 : STD_LOGIC;
    SIGNAL S2845 : STD_LOGIC;
    SIGNAL S2846 : STD_LOGIC;
    SIGNAL S2847 : STD_LOGIC;
    SIGNAL S2848 : STD_LOGIC;
    SIGNAL S2849 : STD_LOGIC;
    SIGNAL S2850 : STD_LOGIC;
    SIGNAL S2851 : STD_LOGIC;
    SIGNAL S2852 : STD_LOGIC;
    SIGNAL S2853 : STD_LOGIC;
    SIGNAL S2854 : STD_LOGIC;
    SIGNAL S2855 : STD_LOGIC;
    SIGNAL S2856 : STD_LOGIC;
    SIGNAL S2857 : STD_LOGIC;
    SIGNAL S2858 : STD_LOGIC;
    SIGNAL S2859 : STD_LOGIC;
    SIGNAL S2860 : STD_LOGIC;
    SIGNAL S2861 : STD_LOGIC;
    SIGNAL S2862 : STD_LOGIC;
    SIGNAL S2863 : STD_LOGIC;
    SIGNAL S2864 : STD_LOGIC;
    SIGNAL S2865 : STD_LOGIC;
    SIGNAL S2866 : STD_LOGIC;
    SIGNAL S2867 : STD_LOGIC;
    SIGNAL S2868 : STD_LOGIC;
    SIGNAL S2869 : STD_LOGIC;
    SIGNAL S2870 : STD_LOGIC;
    SIGNAL S2871 : STD_LOGIC;
    SIGNAL S2872 : STD_LOGIC;
    SIGNAL S2873 : STD_LOGIC;
    SIGNAL S2874 : STD_LOGIC;
    SIGNAL S2875 : STD_LOGIC;
    SIGNAL S2876 : STD_LOGIC;
    SIGNAL S2877 : STD_LOGIC;
    SIGNAL S2878 : STD_LOGIC;
    SIGNAL S2879 : STD_LOGIC;
    SIGNAL S2880 : STD_LOGIC;
    SIGNAL S2881 : STD_LOGIC;
    SIGNAL S2882 : STD_LOGIC;
    SIGNAL S2883 : STD_LOGIC;
    SIGNAL S2884 : STD_LOGIC;
    SIGNAL S2885 : STD_LOGIC;
    SIGNAL S2886 : STD_LOGIC;
    SIGNAL S2887 : STD_LOGIC;
    SIGNAL S2888 : STD_LOGIC;
    SIGNAL S2889 : STD_LOGIC;
    SIGNAL S2890 : STD_LOGIC;
    SIGNAL S2891 : STD_LOGIC;
    SIGNAL S2892 : STD_LOGIC;
    SIGNAL S2893 : STD_LOGIC;
    SIGNAL S2894 : STD_LOGIC;
    SIGNAL S2895 : STD_LOGIC;
    SIGNAL S2896 : STD_LOGIC;
    SIGNAL S2897 : STD_LOGIC;
    SIGNAL S2898 : STD_LOGIC;
    SIGNAL S2899 : STD_LOGIC;
    SIGNAL S2900 : STD_LOGIC;
    SIGNAL S2901 : STD_LOGIC;
    SIGNAL S2902 : STD_LOGIC;
    SIGNAL S2903 : STD_LOGIC;
    SIGNAL S2904 : STD_LOGIC;
    SIGNAL S2905 : STD_LOGIC;
    SIGNAL S2906 : STD_LOGIC;
    SIGNAL S2907 : STD_LOGIC;
    SIGNAL S2908 : STD_LOGIC;
    SIGNAL S2909 : STD_LOGIC;
    SIGNAL S2910 : STD_LOGIC;
    SIGNAL S2911 : STD_LOGIC;
    SIGNAL S2912 : STD_LOGIC;
    SIGNAL S2913 : STD_LOGIC;
    SIGNAL S2914 : STD_LOGIC;
    SIGNAL S2915 : STD_LOGIC;
    SIGNAL S2916 : STD_LOGIC;
    SIGNAL S2917 : STD_LOGIC;
    SIGNAL S2918 : STD_LOGIC;
    SIGNAL S2919 : STD_LOGIC;
    SIGNAL S2920 : STD_LOGIC;
    SIGNAL S2921 : STD_LOGIC;
    SIGNAL S2922 : STD_LOGIC;
    SIGNAL S2923 : STD_LOGIC;
    SIGNAL S2924 : STD_LOGIC;
    SIGNAL S2925 : STD_LOGIC;
    SIGNAL S2926 : STD_LOGIC;
    SIGNAL S2927 : STD_LOGIC;
    SIGNAL S2928 : STD_LOGIC;
    SIGNAL S2929 : STD_LOGIC;
    SIGNAL S2930 : STD_LOGIC;
    SIGNAL S2931 : STD_LOGIC;
    SIGNAL S2932 : STD_LOGIC;
    SIGNAL S2933 : STD_LOGIC;
    SIGNAL S2934 : STD_LOGIC;
    SIGNAL S2935 : STD_LOGIC;
    SIGNAL S2936 : STD_LOGIC;
    SIGNAL S2937 : STD_LOGIC;
    SIGNAL S2938 : STD_LOGIC;
    SIGNAL S2939 : STD_LOGIC;
    SIGNAL S2940 : STD_LOGIC;
    SIGNAL S2941 : STD_LOGIC;
    SIGNAL S2942 : STD_LOGIC;
    SIGNAL S2943 : STD_LOGIC;
    SIGNAL S2944 : STD_LOGIC;
    SIGNAL S2945 : STD_LOGIC;
    SIGNAL S2946 : STD_LOGIC;
    SIGNAL S2947 : STD_LOGIC;
    SIGNAL S2948 : STD_LOGIC;
    SIGNAL S2949 : STD_LOGIC;
    SIGNAL S2950 : STD_LOGIC;
    SIGNAL S2951 : STD_LOGIC;
    SIGNAL S2952 : STD_LOGIC;
    SIGNAL S2953 : STD_LOGIC;
    SIGNAL S2954 : STD_LOGIC;
    SIGNAL S2955 : STD_LOGIC;
    SIGNAL S2956 : STD_LOGIC;
    SIGNAL S2957 : STD_LOGIC;
    SIGNAL S2958 : STD_LOGIC;
    SIGNAL S2959 : STD_LOGIC;
    SIGNAL S2960 : STD_LOGIC;
    SIGNAL S2961 : STD_LOGIC;
    SIGNAL S2962 : STD_LOGIC;
    SIGNAL S2963 : STD_LOGIC;
    SIGNAL S2964 : STD_LOGIC;
    SIGNAL S2965 : STD_LOGIC;
    SIGNAL S2966 : STD_LOGIC;
    SIGNAL S2967 : STD_LOGIC;
    SIGNAL S2968 : STD_LOGIC;
    SIGNAL S2969 : STD_LOGIC;
    SIGNAL S2970 : STD_LOGIC;
    SIGNAL S2971 : STD_LOGIC;
    SIGNAL S2972 : STD_LOGIC;
    SIGNAL S2973 : STD_LOGIC;
    SIGNAL S2974 : STD_LOGIC;
    SIGNAL S2975 : STD_LOGIC;
    SIGNAL S2976 : STD_LOGIC;
    SIGNAL S2977 : STD_LOGIC;
    SIGNAL S2978 : STD_LOGIC;
    SIGNAL S2979 : STD_LOGIC;
    SIGNAL S2980 : STD_LOGIC;
    SIGNAL S2981 : STD_LOGIC;
    SIGNAL S2982 : STD_LOGIC;
    SIGNAL S2983 : STD_LOGIC;
    SIGNAL S2984 : STD_LOGIC;
    SIGNAL S2985 : STD_LOGIC;
    SIGNAL S2986 : STD_LOGIC;
    SIGNAL S2987 : STD_LOGIC;
    SIGNAL S2988 : STD_LOGIC;
    SIGNAL S2989 : STD_LOGIC;
    SIGNAL S2990 : STD_LOGIC;
    SIGNAL S2991 : STD_LOGIC;
    SIGNAL S2992 : STD_LOGIC;
    SIGNAL S2993 : STD_LOGIC;
    SIGNAL S2994 : STD_LOGIC;
    SIGNAL S2995 : STD_LOGIC;
    SIGNAL S2996 : STD_LOGIC;
    SIGNAL S2997 : STD_LOGIC;
    SIGNAL S2998 : STD_LOGIC;
    SIGNAL S2999 : STD_LOGIC;
    SIGNAL S3000 : STD_LOGIC;
    SIGNAL S3001 : STD_LOGIC;
    SIGNAL S3002 : STD_LOGIC;
    SIGNAL S3003 : STD_LOGIC;
    SIGNAL S3004 : STD_LOGIC;
    SIGNAL S3005 : STD_LOGIC;
    SIGNAL S3006 : STD_LOGIC;
    SIGNAL S3007 : STD_LOGIC;
    SIGNAL S3008 : STD_LOGIC;
    SIGNAL S3009 : STD_LOGIC;
    SIGNAL S3010 : STD_LOGIC;
    SIGNAL S3011 : STD_LOGIC;
    SIGNAL S3012 : STD_LOGIC;
    SIGNAL S3013 : STD_LOGIC;
    SIGNAL S3014 : STD_LOGIC;
    SIGNAL S3015 : STD_LOGIC;
    SIGNAL S3016 : STD_LOGIC;
    SIGNAL S3017 : STD_LOGIC;
    SIGNAL S3018 : STD_LOGIC;
    SIGNAL S3019 : STD_LOGIC;
    SIGNAL S3020 : STD_LOGIC;
    SIGNAL S3021 : STD_LOGIC;
    SIGNAL S3022 : STD_LOGIC;
    SIGNAL S3023 : STD_LOGIC;
    SIGNAL S3024 : STD_LOGIC;
    SIGNAL S3025 : STD_LOGIC;
    SIGNAL S3026 : STD_LOGIC;
    SIGNAL S3027 : STD_LOGIC;
    SIGNAL S3028 : STD_LOGIC;
    SIGNAL S3029 : STD_LOGIC;
    SIGNAL S3030 : STD_LOGIC;
    SIGNAL S3031 : STD_LOGIC;
    SIGNAL S3032 : STD_LOGIC;
    SIGNAL S3033 : STD_LOGIC;
    SIGNAL S3034 : STD_LOGIC;
    SIGNAL S3035 : STD_LOGIC;
    SIGNAL S3036 : STD_LOGIC;
    SIGNAL S3037 : STD_LOGIC;
    SIGNAL S3038 : STD_LOGIC;
    SIGNAL S3039 : STD_LOGIC;
    SIGNAL S3040 : STD_LOGIC;
    SIGNAL S3041 : STD_LOGIC;
    SIGNAL S3042 : STD_LOGIC;
    SIGNAL S3043 : STD_LOGIC;
    SIGNAL S3044 : STD_LOGIC;
    SIGNAL S3045 : STD_LOGIC;
    SIGNAL S3046 : STD_LOGIC;
    SIGNAL S3047 : STD_LOGIC;
    SIGNAL S3048 : STD_LOGIC;
    SIGNAL S3049 : STD_LOGIC;
    SIGNAL S3050 : STD_LOGIC;
    SIGNAL S3051 : STD_LOGIC;
    SIGNAL S3052 : STD_LOGIC;
    SIGNAL S3053 : STD_LOGIC;
    SIGNAL S3054 : STD_LOGIC;
    SIGNAL S3055 : STD_LOGIC;
    SIGNAL S3056 : STD_LOGIC;
    SIGNAL S3057 : STD_LOGIC;
    SIGNAL S3058 : STD_LOGIC;
    SIGNAL S3059 : STD_LOGIC;
    SIGNAL S3060 : STD_LOGIC;
    SIGNAL S3061 : STD_LOGIC;
    SIGNAL S3062 : STD_LOGIC;
    SIGNAL S3063 : STD_LOGIC;
    SIGNAL S3064 : STD_LOGIC;
    SIGNAL S3065 : STD_LOGIC;
    SIGNAL S3066 : STD_LOGIC;
    SIGNAL S3067 : STD_LOGIC;
    SIGNAL S3068 : STD_LOGIC;
    SIGNAL S3069 : STD_LOGIC;
    SIGNAL S3070 : STD_LOGIC;
    SIGNAL S3071 : STD_LOGIC;
    SIGNAL S3072 : STD_LOGIC;
    SIGNAL S3073 : STD_LOGIC;
    SIGNAL S3074 : STD_LOGIC;
    SIGNAL S3075 : STD_LOGIC;
    SIGNAL S3076 : STD_LOGIC;
    SIGNAL S3077 : STD_LOGIC;
    SIGNAL S3078 : STD_LOGIC;
    SIGNAL S3079 : STD_LOGIC;
    SIGNAL S3080 : STD_LOGIC;
    SIGNAL S3081 : STD_LOGIC;
    SIGNAL S3082 : STD_LOGIC;
    SIGNAL S3083 : STD_LOGIC;
    SIGNAL S3084 : STD_LOGIC;
    SIGNAL S3085 : STD_LOGIC;
    SIGNAL S3086 : STD_LOGIC;
    SIGNAL S3087 : STD_LOGIC;
    SIGNAL S3088 : STD_LOGIC;
    SIGNAL S3089 : STD_LOGIC;
    SIGNAL S3090 : STD_LOGIC;
    SIGNAL S3091 : STD_LOGIC;
    SIGNAL S3092 : STD_LOGIC;
    SIGNAL S3093 : STD_LOGIC;
    SIGNAL S3094 : STD_LOGIC;
    SIGNAL S3095 : STD_LOGIC;
    SIGNAL S3096 : STD_LOGIC;
    SIGNAL S3097 : STD_LOGIC;
    SIGNAL S3098 : STD_LOGIC;
    SIGNAL S3099 : STD_LOGIC;
    SIGNAL S3100 : STD_LOGIC;
    SIGNAL S3101 : STD_LOGIC;
    SIGNAL S3102 : STD_LOGIC;
    SIGNAL S3103 : STD_LOGIC;
    SIGNAL S3104 : STD_LOGIC;
    SIGNAL S3105 : STD_LOGIC;
    SIGNAL S3106 : STD_LOGIC;
    SIGNAL S3107 : STD_LOGIC;
    SIGNAL S3108 : STD_LOGIC;
    SIGNAL S3109 : STD_LOGIC;
    SIGNAL S3110 : STD_LOGIC;
    SIGNAL S3111 : STD_LOGIC;
    SIGNAL S3112 : STD_LOGIC;
    SIGNAL S3113 : STD_LOGIC;
    SIGNAL S3114 : STD_LOGIC;
    SIGNAL S3115 : STD_LOGIC;
    SIGNAL S3116 : STD_LOGIC;
    SIGNAL S3117 : STD_LOGIC;
    SIGNAL S3118 : STD_LOGIC;
    SIGNAL S3119 : STD_LOGIC;
    SIGNAL S3120 : STD_LOGIC;
    SIGNAL S3121 : STD_LOGIC;
    SIGNAL S3122 : STD_LOGIC;
    SIGNAL S3123 : STD_LOGIC;
    SIGNAL S3124 : STD_LOGIC;
    SIGNAL S3125 : STD_LOGIC;
    SIGNAL S3126 : STD_LOGIC;
    SIGNAL S3127 : STD_LOGIC;
    SIGNAL S3128 : STD_LOGIC;
    SIGNAL S3129 : STD_LOGIC;
    SIGNAL S3130 : STD_LOGIC;
    SIGNAL S3131 : STD_LOGIC;
    SIGNAL S3132 : STD_LOGIC;
    SIGNAL S3133 : STD_LOGIC;
    SIGNAL S3134 : STD_LOGIC;
    SIGNAL S3135 : STD_LOGIC;
    SIGNAL S3136 : STD_LOGIC;
    SIGNAL S3137 : STD_LOGIC;
    SIGNAL S3138 : STD_LOGIC;
    SIGNAL S3139 : STD_LOGIC;
    SIGNAL S3140 : STD_LOGIC;
    SIGNAL S3141 : STD_LOGIC;
    SIGNAL S3142 : STD_LOGIC;
    SIGNAL S3143 : STD_LOGIC;
    SIGNAL S3144 : STD_LOGIC;
    SIGNAL S3145 : STD_LOGIC;
    SIGNAL S3146 : STD_LOGIC;
    SIGNAL S3147 : STD_LOGIC;
    SIGNAL S3148 : STD_LOGIC;
    SIGNAL S3149 : STD_LOGIC;
    SIGNAL S3150 : STD_LOGIC;
    SIGNAL S3151 : STD_LOGIC;
    SIGNAL S3152 : STD_LOGIC;
    SIGNAL S3153 : STD_LOGIC;
    SIGNAL S3154 : STD_LOGIC;
    SIGNAL S3155 : STD_LOGIC;
    SIGNAL S3156 : STD_LOGIC;
    SIGNAL S3157 : STD_LOGIC;
    SIGNAL S3158 : STD_LOGIC;
    SIGNAL S3159 : STD_LOGIC;
    SIGNAL S3160 : STD_LOGIC;
    SIGNAL S3161 : STD_LOGIC;
    SIGNAL S3162 : STD_LOGIC;
    SIGNAL S3163 : STD_LOGIC;
    SIGNAL S3164 : STD_LOGIC;
    SIGNAL S3165 : STD_LOGIC;
    SIGNAL S3166 : STD_LOGIC;
    SIGNAL S3167 : STD_LOGIC;
    SIGNAL S3168 : STD_LOGIC;
    SIGNAL S3169 : STD_LOGIC;
    SIGNAL S3170 : STD_LOGIC;
    SIGNAL S3171 : STD_LOGIC;
    SIGNAL S3172 : STD_LOGIC;
    SIGNAL S3173 : STD_LOGIC;
    SIGNAL S3174 : STD_LOGIC;
    SIGNAL S3175 : STD_LOGIC;
    SIGNAL S3176 : STD_LOGIC;
    SIGNAL S3177 : STD_LOGIC;
    SIGNAL S3178 : STD_LOGIC;
    SIGNAL S3179 : STD_LOGIC;
    SIGNAL S3180 : STD_LOGIC;
    SIGNAL S3181 : STD_LOGIC;
    SIGNAL S3182 : STD_LOGIC;
    SIGNAL S3183 : STD_LOGIC;
    SIGNAL S3184 : STD_LOGIC;
    SIGNAL S3185 : STD_LOGIC;
    SIGNAL S3186 : STD_LOGIC;
    SIGNAL S3187 : STD_LOGIC;
    SIGNAL S3188 : STD_LOGIC;
    SIGNAL S3189 : STD_LOGIC;
    SIGNAL S3190 : STD_LOGIC;
    SIGNAL S3191 : STD_LOGIC;
    SIGNAL S3192 : STD_LOGIC;
    SIGNAL S3193 : STD_LOGIC;
    SIGNAL S3194 : STD_LOGIC;
    SIGNAL S3195 : STD_LOGIC;
    SIGNAL S3196 : STD_LOGIC;
    SIGNAL S3197 : STD_LOGIC;
    SIGNAL S3198 : STD_LOGIC;
    SIGNAL S3199 : STD_LOGIC;
    SIGNAL S3200 : STD_LOGIC;
    SIGNAL S3201 : STD_LOGIC;
    SIGNAL S3202 : STD_LOGIC;
    SIGNAL S3203 : STD_LOGIC;
    SIGNAL S3204 : STD_LOGIC;
    SIGNAL S3205 : STD_LOGIC;
    SIGNAL S3206 : STD_LOGIC;
    SIGNAL S3207 : STD_LOGIC;
    SIGNAL S3208 : STD_LOGIC;
    SIGNAL S3209 : STD_LOGIC;
    SIGNAL S3210 : STD_LOGIC;
    SIGNAL S3211 : STD_LOGIC;
    SIGNAL S3212 : STD_LOGIC;
    SIGNAL S3213 : STD_LOGIC;
    SIGNAL S3214 : STD_LOGIC;
    SIGNAL S3215 : STD_LOGIC;
    SIGNAL S3216 : STD_LOGIC;
    SIGNAL S3217 : STD_LOGIC;
    SIGNAL S3218 : STD_LOGIC;
    SIGNAL S3219 : STD_LOGIC;
    SIGNAL S3220 : STD_LOGIC;
    SIGNAL S3221 : STD_LOGIC;
    SIGNAL S3222 : STD_LOGIC;
    SIGNAL S3223 : STD_LOGIC;
    SIGNAL S3224 : STD_LOGIC;
    SIGNAL S3225 : STD_LOGIC;
    SIGNAL S3226 : STD_LOGIC;
    SIGNAL S3227 : STD_LOGIC;
    SIGNAL S3228 : STD_LOGIC;
    SIGNAL S3229 : STD_LOGIC;
    SIGNAL S3230 : STD_LOGIC;
    SIGNAL S3231 : STD_LOGIC;
    SIGNAL S3232 : STD_LOGIC;
    SIGNAL S3233 : STD_LOGIC;
    SIGNAL S3234 : STD_LOGIC;
    SIGNAL S3235 : STD_LOGIC;
    SIGNAL S3236 : STD_LOGIC;
    SIGNAL S3237 : STD_LOGIC;
    SIGNAL S3238 : STD_LOGIC;
    SIGNAL S3239 : STD_LOGIC;
    SIGNAL S3240 : STD_LOGIC;
    SIGNAL S3241 : STD_LOGIC;
    SIGNAL S3242 : STD_LOGIC;
    SIGNAL S3243 : STD_LOGIC;
    SIGNAL S3244 : STD_LOGIC;
    SIGNAL S3245 : STD_LOGIC;
    SIGNAL S3246 : STD_LOGIC;
    SIGNAL S3247 : STD_LOGIC;
    SIGNAL S3248 : STD_LOGIC;
    SIGNAL S3249 : STD_LOGIC;
    SIGNAL S3250 : STD_LOGIC;
    SIGNAL S3251 : STD_LOGIC;
    SIGNAL S3252 : STD_LOGIC;
    SIGNAL S3253 : STD_LOGIC;
    SIGNAL S3254 : STD_LOGIC;
    SIGNAL S3255 : STD_LOGIC;
    SIGNAL S3256 : STD_LOGIC;
    SIGNAL S3257 : STD_LOGIC;
    SIGNAL S3258 : STD_LOGIC;
    SIGNAL S3259 : STD_LOGIC;
    SIGNAL S3260 : STD_LOGIC;
    SIGNAL S3261 : STD_LOGIC;
    SIGNAL S3262 : STD_LOGIC;
    SIGNAL S3263 : STD_LOGIC;
    SIGNAL S3264 : STD_LOGIC;
    SIGNAL S3265 : STD_LOGIC;
    SIGNAL S3266 : STD_LOGIC;
    SIGNAL S3267 : STD_LOGIC;
    SIGNAL S3268 : STD_LOGIC;
    SIGNAL S3269 : STD_LOGIC;
    SIGNAL S3270 : STD_LOGIC;
    SIGNAL S3271 : STD_LOGIC;
    SIGNAL S3272 : STD_LOGIC;
    SIGNAL S3273 : STD_LOGIC;
    SIGNAL S3274 : STD_LOGIC;
    SIGNAL S3275 : STD_LOGIC;
    SIGNAL S3276 : STD_LOGIC;
    SIGNAL S3277 : STD_LOGIC;
    SIGNAL S3278 : STD_LOGIC;
    SIGNAL S3279 : STD_LOGIC;
    SIGNAL S3280 : STD_LOGIC;
    SIGNAL S3281 : STD_LOGIC;
    SIGNAL S3282 : STD_LOGIC;
    SIGNAL S3283 : STD_LOGIC;
    SIGNAL S3284 : STD_LOGIC;
    SIGNAL S3285 : STD_LOGIC;
    SIGNAL S3286 : STD_LOGIC;
    SIGNAL S3287 : STD_LOGIC;
    SIGNAL S3288 : STD_LOGIC;
    SIGNAL S3289 : STD_LOGIC;
    SIGNAL S3290 : STD_LOGIC;
    SIGNAL S3291 : STD_LOGIC;
    SIGNAL S3292 : STD_LOGIC;
    SIGNAL S3293 : STD_LOGIC;
    SIGNAL S3294 : STD_LOGIC;
    SIGNAL S3295 : STD_LOGIC;
    SIGNAL S3296 : STD_LOGIC;
    SIGNAL S3297 : STD_LOGIC;
    SIGNAL S3298 : STD_LOGIC;
    SIGNAL S3299 : STD_LOGIC;
    SIGNAL S3300 : STD_LOGIC;
    SIGNAL S3301 : STD_LOGIC;
    SIGNAL S3302 : STD_LOGIC;
    SIGNAL S3303 : STD_LOGIC;
    SIGNAL S3304 : STD_LOGIC;
    SIGNAL S3305 : STD_LOGIC;
    SIGNAL S3306 : STD_LOGIC;
    SIGNAL S3307 : STD_LOGIC;
    SIGNAL S3308 : STD_LOGIC;
    SIGNAL S3309 : STD_LOGIC;
    SIGNAL S3310 : STD_LOGIC;
    SIGNAL S3311 : STD_LOGIC;
    SIGNAL S3312 : STD_LOGIC;
    SIGNAL S3313 : STD_LOGIC;
    SIGNAL S3314 : STD_LOGIC;
    SIGNAL S3315 : STD_LOGIC;
    SIGNAL S3316 : STD_LOGIC;
    SIGNAL S3317 : STD_LOGIC;
    SIGNAL S3318 : STD_LOGIC;
    SIGNAL S3319 : STD_LOGIC;
    SIGNAL S3320 : STD_LOGIC;
    SIGNAL S3321 : STD_LOGIC;
    SIGNAL S3322 : STD_LOGIC;
    SIGNAL S3323 : STD_LOGIC;
    SIGNAL S3324 : STD_LOGIC;
    SIGNAL S3325 : STD_LOGIC;
    SIGNAL S3326 : STD_LOGIC;
    SIGNAL S3327 : STD_LOGIC;
    SIGNAL S3328 : STD_LOGIC;
    SIGNAL S3329 : STD_LOGIC;
    SIGNAL S3330 : STD_LOGIC;
    SIGNAL S3331 : STD_LOGIC;
    SIGNAL S3332 : STD_LOGIC;
    SIGNAL S3333 : STD_LOGIC;
    SIGNAL S3334 : STD_LOGIC;
    SIGNAL S3335 : STD_LOGIC;
    SIGNAL S3336 : STD_LOGIC;
    SIGNAL S3337 : STD_LOGIC;
    SIGNAL S3338 : STD_LOGIC;
    SIGNAL S3339 : STD_LOGIC;
    SIGNAL S3340 : STD_LOGIC;
    SIGNAL S3341 : STD_LOGIC;
    SIGNAL S3342 : STD_LOGIC;
    SIGNAL S3343 : STD_LOGIC;
    SIGNAL S3344 : STD_LOGIC;
    SIGNAL S3345 : STD_LOGIC;
    SIGNAL S3346 : STD_LOGIC;
    SIGNAL S3347 : STD_LOGIC;
    SIGNAL S3348 : STD_LOGIC;
    SIGNAL S3349 : STD_LOGIC;
    SIGNAL S3350 : STD_LOGIC;
    SIGNAL S3351 : STD_LOGIC;
    SIGNAL S3352 : STD_LOGIC;
    SIGNAL S3353 : STD_LOGIC;
    SIGNAL S3354 : STD_LOGIC;
    SIGNAL S3355 : STD_LOGIC;
    SIGNAL S3356 : STD_LOGIC;
    SIGNAL S3357 : STD_LOGIC;
    SIGNAL S3358 : STD_LOGIC;
    SIGNAL S3359 : STD_LOGIC;
    SIGNAL S3360 : STD_LOGIC;
    SIGNAL S3361 : STD_LOGIC;
    SIGNAL S3362 : STD_LOGIC;
    SIGNAL S3363 : STD_LOGIC;
    SIGNAL S3364 : STD_LOGIC;
    SIGNAL S3365 : STD_LOGIC;
    SIGNAL S3366 : STD_LOGIC;
    SIGNAL CU_ADD : STD_LOGIC;
    SIGNAL CU_AND : STD_LOGIC;
    SIGNAL CU_INC1 : STD_LOGIC;
    SIGNAL CU_INC2 : STD_LOGIC;
    SIGNAL CU_LSB0E : STD_LOGIC;
    SIGNAL CU_MUL : STD_LOGIC;
    SIGNAL CU_NOT : STD_LOGIC;
    SIGNAL CU_SE12bits : STD_LOGIC;
    SIGNAL CU_SE4bits : STD_LOGIC;
    SIGNAL CU_SHF_0 : STD_LOGIC;
    SIGNAL CU_SHF_1 : STD_LOGIC;
    SIGNAL CU_clk : STD_LOGIC;
    SIGNAL CU_conOF : STD_LOGIC;
    SIGNAL CU_enSKP : STD_LOGIC;
    SIGNAL CU_inst_0 : STD_LOGIC;
    SIGNAL CU_inst_10 : STD_LOGIC;
    SIGNAL CU_inst_11 : STD_LOGIC;
    SIGNAL CU_inst_12 : STD_LOGIC;
    SIGNAL CU_inst_13 : STD_LOGIC;
    SIGNAL CU_inst_14 : STD_LOGIC;
    SIGNAL CU_inst_15 : STD_LOGIC;
    SIGNAL CU_inst_1 : STD_LOGIC;
    SIGNAL CU_inst_2 : STD_LOGIC;
    SIGNAL CU_inst_3 : STD_LOGIC;
    SIGNAL CU_inst_4 : STD_LOGIC;
    SIGNAL CU_inst_5 : STD_LOGIC;
    SIGNAL CU_inst_6 : STD_LOGIC;
    SIGNAL CU_inst_7 : STD_LOGIC;
    SIGNAL CU_inst_8 : STD_LOGIC;
    SIGNAL CU_inst_9 : STD_LOGIC;
    SIGNAL CU_ldAC : STD_LOGIC;
    SIGNAL CU_ldIN : STD_LOGIC;
    SIGNAL CU_ldIR : STD_LOGIC;
    SIGNAL CU_ldOF : STD_LOGIC;
    SIGNAL CU_ldPC : STD_LOGIC;
    SIGNAL CU_ldSR_0 : STD_LOGIC;
    SIGNAL CU_ldSR_1 : STD_LOGIC;
    SIGNAL CU_ldSR_2 : STD_LOGIC;
    SIGNAL CU_ldSR_3 : STD_LOGIC;
    SIGNAL CU_nstate_0 : STD_LOGIC;
    SIGNAL CU_nstate_1 : STD_LOGIC;
    SIGNAL CU_pstate_0 : STD_LOGIC;
    SIGNAL CU_pstate_1 : STD_LOGIC;
    SIGNAL CU_readMEM : STD_LOGIC;
    SIGNAL CU_rst : STD_LOGIC;
    SIGNAL CU_sel1_ARU : STD_LOGIC;
    SIGNAL CU_selAC_MEM : STD_LOGIC;
    SIGNAL CU_selARU_AC : STD_LOGIC;
    SIGNAL CU_selARU_SR : STD_LOGIC;
    SIGNAL CU_selIMM_AC : STD_LOGIC;
    SIGNAL CU_selIMM_LGU : STD_LOGIC;
    SIGNAL CU_selIMM_OF : STD_LOGIC;
    SIGNAL CU_selIMM_PC : STD_LOGIC;
    SIGNAL CU_selINC_IN : STD_LOGIC;
    SIGNAL CU_selINC_PC : STD_LOGIC;
    SIGNAL CU_selIN_ADR : STD_LOGIC;
    SIGNAL CU_selIN_MEM : STD_LOGIC;
    SIGNAL CU_selIR_ADR : STD_LOGIC;
    SIGNAL CU_selLGU_AC : STD_LOGIC;
    SIGNAL CU_selLGU_SR : STD_LOGIC;
    SIGNAL CU_selMEM_AC : STD_LOGIC;
    SIGNAL CU_selMEM_IN : STD_LOGIC;
    SIGNAL CU_selMEM_LGU : STD_LOGIC;
    SIGNAL CU_selMEM_PC : STD_LOGIC;
    SIGNAL CU_selPC_MEM : STD_LOGIC;
    SIGNAL CU_selPC_OF : STD_LOGIC;
    SIGNAL CU_selSET_SR : STD_LOGIC;
    SIGNAL CU_seldataBus : STD_LOGIC;
    SIGNAL CU_zeroAC : STD_LOGIC;
    SIGNAL DP_AC_in_0 : STD_LOGIC;
    SIGNAL DP_AC_in_10 : STD_LOGIC;
    SIGNAL DP_AC_in_11 : STD_LOGIC;
    SIGNAL DP_AC_in_12 : STD_LOGIC;
    SIGNAL DP_AC_in_13 : STD_LOGIC;
    SIGNAL DP_AC_in_14 : STD_LOGIC;
    SIGNAL DP_AC_in_15 : STD_LOGIC;
    SIGNAL DP_AC_in_1 : STD_LOGIC;
    SIGNAL DP_AC_in_2 : STD_LOGIC;
    SIGNAL DP_AC_in_3 : STD_LOGIC;
    SIGNAL DP_AC_in_4 : STD_LOGIC;
    SIGNAL DP_AC_in_5 : STD_LOGIC;
    SIGNAL DP_AC_in_6 : STD_LOGIC;
    SIGNAL DP_AC_in_7 : STD_LOGIC;
    SIGNAL DP_AC_in_8 : STD_LOGIC;
    SIGNAL DP_AC_in_9 : STD_LOGIC;
    SIGNAL DP_AC_out_0 : STD_LOGIC;
    SIGNAL DP_AC_out_10 : STD_LOGIC;
    SIGNAL DP_AC_out_11 : STD_LOGIC;
    SIGNAL DP_AC_out_12 : STD_LOGIC;
    SIGNAL DP_AC_out_13 : STD_LOGIC;
    SIGNAL DP_AC_out_14 : STD_LOGIC;
    SIGNAL DP_AC_out_15 : STD_LOGIC;
    SIGNAL DP_AC_out_1 : STD_LOGIC;
    SIGNAL DP_AC_out_2 : STD_LOGIC;
    SIGNAL DP_AC_out_3 : STD_LOGIC;
    SIGNAL DP_AC_out_4 : STD_LOGIC;
    SIGNAL DP_AC_out_5 : STD_LOGIC;
    SIGNAL DP_AC_out_6 : STD_LOGIC;
    SIGNAL DP_AC_out_7 : STD_LOGIC;
    SIGNAL DP_AC_out_8 : STD_LOGIC;
    SIGNAL DP_AC_out_9 : STD_LOGIC;
    SIGNAL DP_ARU1_C : STD_LOGIC;
    SIGNAL DP_ARU1_N : STD_LOGIC;
    SIGNAL DP_ARU1_V : STD_LOGIC;
    SIGNAL DP_ARU1_Z : STD_LOGIC;
    SIGNAL DP_ARU1_in1_0 : STD_LOGIC;
    SIGNAL DP_ARU1_in1_10 : STD_LOGIC;
    SIGNAL DP_ARU1_in1_11 : STD_LOGIC;
    SIGNAL DP_ARU1_in1_12 : STD_LOGIC;
    SIGNAL DP_ARU1_in1_13 : STD_LOGIC;
    SIGNAL DP_ARU1_in1_14 : STD_LOGIC;
    SIGNAL DP_ARU1_in1_15 : STD_LOGIC;
    SIGNAL DP_ARU1_in1_1 : STD_LOGIC;
    SIGNAL DP_ARU1_in1_2 : STD_LOGIC;
    SIGNAL DP_ARU1_in1_3 : STD_LOGIC;
    SIGNAL DP_ARU1_in1_4 : STD_LOGIC;
    SIGNAL DP_ARU1_in1_5 : STD_LOGIC;
    SIGNAL DP_ARU1_in1_6 : STD_LOGIC;
    SIGNAL DP_ARU1_in1_7 : STD_LOGIC;
    SIGNAL DP_ARU1_in1_8 : STD_LOGIC;
    SIGNAL DP_ARU1_in1_9 : STD_LOGIC;
    SIGNAL DP_ARU1_out_0 : STD_LOGIC;
    SIGNAL DP_ARU1_out_10 : STD_LOGIC;
    SIGNAL DP_ARU1_out_11 : STD_LOGIC;
    SIGNAL DP_ARU1_out_12 : STD_LOGIC;
    SIGNAL DP_ARU1_out_13 : STD_LOGIC;
    SIGNAL DP_ARU1_out_14 : STD_LOGIC;
    SIGNAL DP_ARU1_out_1 : STD_LOGIC;
    SIGNAL DP_ARU1_out_2 : STD_LOGIC;
    SIGNAL DP_ARU1_out_3 : STD_LOGIC;
    SIGNAL DP_ARU1_out_4 : STD_LOGIC;
    SIGNAL DP_ARU1_out_5 : STD_LOGIC;
    SIGNAL DP_ARU1_out_6 : STD_LOGIC;
    SIGNAL DP_ARU1_out_7 : STD_LOGIC;
    SIGNAL DP_ARU1_out_8 : STD_LOGIC;
    SIGNAL DP_ARU1_out_9 : STD_LOGIC;
    SIGNAL DP_IMM1_in1_0 : STD_LOGIC;
    SIGNAL DP_IMM1_in1_1 : STD_LOGIC;
    SIGNAL DP_IMM1_in1_2 : STD_LOGIC;
    SIGNAL DP_IMM1_in1_3 : STD_LOGIC;
    SIGNAL DP_IMM1_out_0 : STD_LOGIC;
    SIGNAL DP_IMM1_out_10 : STD_LOGIC;
    SIGNAL DP_IMM1_out_11 : STD_LOGIC;
    SIGNAL DP_IMM1_out_12 : STD_LOGIC;
    SIGNAL DP_IMM1_out_13 : STD_LOGIC;
    SIGNAL DP_IMM1_out_14 : STD_LOGIC;
    SIGNAL DP_IMM1_out_15 : STD_LOGIC;
    SIGNAL DP_IMM1_out_1 : STD_LOGIC;
    SIGNAL DP_IMM1_out_2 : STD_LOGIC;
    SIGNAL DP_IMM1_out_3 : STD_LOGIC;
    SIGNAL DP_IMM1_out_4 : STD_LOGIC;
    SIGNAL DP_IMM1_out_5 : STD_LOGIC;
    SIGNAL DP_IMM1_out_6 : STD_LOGIC;
    SIGNAL DP_IMM1_out_7 : STD_LOGIC;
    SIGNAL DP_IMM1_out_8 : STD_LOGIC;
    SIGNAL DP_IMM1_out_9 : STD_LOGIC;
    SIGNAL DP_IN_in_0 : STD_LOGIC;
    SIGNAL DP_IN_in_10 : STD_LOGIC;
    SIGNAL DP_IN_in_11 : STD_LOGIC;
    SIGNAL DP_IN_in_12 : STD_LOGIC;
    SIGNAL DP_IN_in_13 : STD_LOGIC;
    SIGNAL DP_IN_in_14 : STD_LOGIC;
    SIGNAL DP_IN_in_15 : STD_LOGIC;
    SIGNAL DP_IN_in_1 : STD_LOGIC;
    SIGNAL DP_IN_in_2 : STD_LOGIC;
    SIGNAL DP_IN_in_3 : STD_LOGIC;
    SIGNAL DP_IN_in_4 : STD_LOGIC;
    SIGNAL DP_IN_in_5 : STD_LOGIC;
    SIGNAL DP_IN_in_6 : STD_LOGIC;
    SIGNAL DP_IN_in_7 : STD_LOGIC;
    SIGNAL DP_IN_in_8 : STD_LOGIC;
    SIGNAL DP_IN_in_9 : STD_LOGIC;
    SIGNAL DP_IN_out_0 : STD_LOGIC;
    SIGNAL DP_IN_out_10 : STD_LOGIC;
    SIGNAL DP_IN_out_11 : STD_LOGIC;
    SIGNAL DP_IN_out_12 : STD_LOGIC;
    SIGNAL DP_IN_out_13 : STD_LOGIC;
    SIGNAL DP_IN_out_14 : STD_LOGIC;
    SIGNAL DP_IN_out_15 : STD_LOGIC;
    SIGNAL DP_IN_out_1 : STD_LOGIC;
    SIGNAL DP_IN_out_2 : STD_LOGIC;
    SIGNAL DP_IN_out_3 : STD_LOGIC;
    SIGNAL DP_IN_out_4 : STD_LOGIC;
    SIGNAL DP_IN_out_5 : STD_LOGIC;
    SIGNAL DP_IN_out_6 : STD_LOGIC;
    SIGNAL DP_IN_out_7 : STD_LOGIC;
    SIGNAL DP_IN_out_8 : STD_LOGIC;
    SIGNAL DP_IN_out_9 : STD_LOGIC;
    SIGNAL DP_INC2_out_0 : STD_LOGIC;
    SIGNAL DP_INC2_out_10 : STD_LOGIC;
    SIGNAL DP_INC2_out_11 : STD_LOGIC;
    SIGNAL DP_INC2_out_12 : STD_LOGIC;
    SIGNAL DP_INC2_out_13 : STD_LOGIC;
    SIGNAL DP_INC2_out_14 : STD_LOGIC;
    SIGNAL DP_INC2_out_15 : STD_LOGIC;
    SIGNAL DP_INC2_out_1 : STD_LOGIC;
    SIGNAL DP_INC2_out_2 : STD_LOGIC;
    SIGNAL DP_INC2_out_3 : STD_LOGIC;
    SIGNAL DP_INC2_out_4 : STD_LOGIC;
    SIGNAL DP_INC2_out_5 : STD_LOGIC;
    SIGNAL DP_INC2_out_6 : STD_LOGIC;
    SIGNAL DP_INC2_out_7 : STD_LOGIC;
    SIGNAL DP_INC2_out_8 : STD_LOGIC;
    SIGNAL DP_INC2_out_9 : STD_LOGIC;
    SIGNAL DP_INC_1_in_0 : STD_LOGIC;
    SIGNAL DP_INC_1_in_10 : STD_LOGIC;
    SIGNAL DP_INC_1_in_11 : STD_LOGIC;
    SIGNAL DP_INC_1_in_12 : STD_LOGIC;
    SIGNAL DP_INC_1_in_13 : STD_LOGIC;
    SIGNAL DP_INC_1_in_14 : STD_LOGIC;
    SIGNAL DP_INC_1_in_15 : STD_LOGIC;
    SIGNAL DP_INC_1_in_1 : STD_LOGIC;
    SIGNAL DP_INC_1_in_2 : STD_LOGIC;
    SIGNAL DP_INC_1_in_3 : STD_LOGIC;
    SIGNAL DP_INC_1_in_4 : STD_LOGIC;
    SIGNAL DP_INC_1_in_5 : STD_LOGIC;
    SIGNAL DP_INC_1_in_6 : STD_LOGIC;
    SIGNAL DP_INC_1_in_7 : STD_LOGIC;
    SIGNAL DP_INC_1_in_8 : STD_LOGIC;
    SIGNAL DP_INC_1_in_9 : STD_LOGIC;
    SIGNAL DP_INC_1_inc_val_0 : STD_LOGIC;
    SIGNAL DP_INC_1_inc_val_1 : STD_LOGIC;
    SIGNAL DP_INC_1_out_0 : STD_LOGIC;
    SIGNAL DP_INC_1_out_10 : STD_LOGIC;
    SIGNAL DP_INC_1_out_11 : STD_LOGIC;
    SIGNAL DP_INC_1_out_12 : STD_LOGIC;
    SIGNAL DP_INC_1_out_13 : STD_LOGIC;
    SIGNAL DP_INC_1_out_14 : STD_LOGIC;
    SIGNAL DP_INC_1_out_15 : STD_LOGIC;
    SIGNAL DP_INC_1_out_1 : STD_LOGIC;
    SIGNAL DP_INC_1_out_2 : STD_LOGIC;
    SIGNAL DP_INC_1_out_3 : STD_LOGIC;
    SIGNAL DP_INC_1_out_4 : STD_LOGIC;
    SIGNAL DP_INC_1_out_5 : STD_LOGIC;
    SIGNAL DP_INC_1_out_6 : STD_LOGIC;
    SIGNAL DP_INC_1_out_7 : STD_LOGIC;
    SIGNAL DP_INC_1_out_8 : STD_LOGIC;
    SIGNAL DP_INC_1_out_9 : STD_LOGIC;
    SIGNAL DP_LGU1_N : STD_LOGIC;
    SIGNAL DP_LGU1_Z : STD_LOGIC;
    SIGNAL DP_LGU1_in1_0 : STD_LOGIC;
    SIGNAL DP_LGU1_in1_10 : STD_LOGIC;
    SIGNAL DP_LGU1_in1_11 : STD_LOGIC;
    SIGNAL DP_LGU1_in1_12 : STD_LOGIC;
    SIGNAL DP_LGU1_in1_13 : STD_LOGIC;
    SIGNAL DP_LGU1_in1_14 : STD_LOGIC;
    SIGNAL DP_LGU1_in1_15 : STD_LOGIC;
    SIGNAL DP_LGU1_in1_1 : STD_LOGIC;
    SIGNAL DP_LGU1_in1_2 : STD_LOGIC;
    SIGNAL DP_LGU1_in1_3 : STD_LOGIC;
    SIGNAL DP_LGU1_in1_4 : STD_LOGIC;
    SIGNAL DP_LGU1_in1_5 : STD_LOGIC;
    SIGNAL DP_LGU1_in1_6 : STD_LOGIC;
    SIGNAL DP_LGU1_in1_7 : STD_LOGIC;
    SIGNAL DP_LGU1_in1_8 : STD_LOGIC;
    SIGNAL DP_LGU1_in1_9 : STD_LOGIC;
    SIGNAL DP_LGU1_out_0 : STD_LOGIC;
    SIGNAL DP_LGU1_out_10 : STD_LOGIC;
    SIGNAL DP_LGU1_out_11 : STD_LOGIC;
    SIGNAL DP_LGU1_out_12 : STD_LOGIC;
    SIGNAL DP_LGU1_out_13 : STD_LOGIC;
    SIGNAL DP_LGU1_out_14 : STD_LOGIC;
    SIGNAL DP_LGU1_out_1 : STD_LOGIC;
    SIGNAL DP_LGU1_out_2 : STD_LOGIC;
    SIGNAL DP_LGU1_out_3 : STD_LOGIC;
    SIGNAL DP_LGU1_out_4 : STD_LOGIC;
    SIGNAL DP_LGU1_out_5 : STD_LOGIC;
    SIGNAL DP_LGU1_out_6 : STD_LOGIC;
    SIGNAL DP_LGU1_out_7 : STD_LOGIC;
    SIGNAL DP_LGU1_out_8 : STD_LOGIC;
    SIGNAL DP_LGU1_out_9 : STD_LOGIC;
    SIGNAL DP_OF_in_0 : STD_LOGIC;
    SIGNAL DP_OF_in_1 : STD_LOGIC;
    SIGNAL DP_OF_in_2 : STD_LOGIC;
    SIGNAL DP_OF_in_3 : STD_LOGIC;
    SIGNAL DP_PC_in_0 : STD_LOGIC;
    SIGNAL DP_PC_in_10 : STD_LOGIC;
    SIGNAL DP_PC_in_11 : STD_LOGIC;
    SIGNAL DP_PC_in_12 : STD_LOGIC;
    SIGNAL DP_PC_in_13 : STD_LOGIC;
    SIGNAL DP_PC_in_14 : STD_LOGIC;
    SIGNAL DP_PC_in_15 : STD_LOGIC;
    SIGNAL DP_PC_in_1 : STD_LOGIC;
    SIGNAL DP_PC_in_2 : STD_LOGIC;
    SIGNAL DP_PC_in_3 : STD_LOGIC;
    SIGNAL DP_PC_in_4 : STD_LOGIC;
    SIGNAL DP_PC_in_5 : STD_LOGIC;
    SIGNAL DP_PC_in_6 : STD_LOGIC;
    SIGNAL DP_PC_in_7 : STD_LOGIC;
    SIGNAL DP_PC_in_8 : STD_LOGIC;
    SIGNAL DP_PC_in_9 : STD_LOGIC;
    SIGNAL DP_SR_C_in : STD_LOGIC;
    SIGNAL DP_SR_C_out : STD_LOGIC;
    SIGNAL DP_SR_N_in : STD_LOGIC;
    SIGNAL DP_SR_N_out : STD_LOGIC;
    SIGNAL DP_SR_V_in : STD_LOGIC;
    SIGNAL DP_SR_V_out : STD_LOGIC;
    SIGNAL DP_SR_Z_in : STD_LOGIC;
    SIGNAL DP_SR_Z_out : STD_LOGIC;
    SIGNAL DP_addrBus_0 : STD_LOGIC;
    SIGNAL DP_addrBus_10 : STD_LOGIC;
    SIGNAL DP_addrBus_11 : STD_LOGIC;
    SIGNAL DP_addrBus_12 : STD_LOGIC;
    SIGNAL DP_addrBus_13 : STD_LOGIC;
    SIGNAL DP_addrBus_14 : STD_LOGIC;
    SIGNAL DP_addrBus_15 : STD_LOGIC;
    SIGNAL DP_addrBus_1 : STD_LOGIC;
    SIGNAL DP_addrBus_2 : STD_LOGIC;
    SIGNAL DP_addrBus_3 : STD_LOGIC;
    SIGNAL DP_addrBus_4 : STD_LOGIC;
    SIGNAL DP_addrBus_5 : STD_LOGIC;
    SIGNAL DP_addrBus_6 : STD_LOGIC;
    SIGNAL DP_addrBus_7 : STD_LOGIC;
    SIGNAL DP_addrBus_8 : STD_LOGIC;
    SIGNAL DP_addrBus_9 : STD_LOGIC;

BEGIN
bufg_1: ENTITY WORK.bufg
    PORT MAP (
        in1 => '1',
        out1 => S0
    );
bufg_2: ENTITY WORK.bufg
    PORT MAP (
        in1 => '1',
        out1 => S1
    );
bufg_3: ENTITY WORK.bufg
    PORT MAP (
        in1 => '1',
        out1 => S2
    );
bufg_4: ENTITY WORK.bufg
    PORT MAP (
        in1 => '1',
        out1 => S3
    );
bufg_5: ENTITY WORK.bufg
    PORT MAP (
        in1 => '1',
        out1 => S4
    );
bufg_6: ENTITY WORK.bufg
    PORT MAP (
        in1 => '1',
        out1 => S5
    );
bufg_7: ENTITY WORK.bufg
    PORT MAP (
        in1 => '0',
        out1 => S6
    );
bufg_8: ENTITY WORK.bufg
    PORT MAP (
        in1 => '0',
        out1 => S7
    );
bufg_9: ENTITY WORK.bufg
    PORT MAP (
        in1 => '0',
        out1 => S8
    );
bufg_10: ENTITY WORK.bufg
    PORT MAP (
        in1 => '0',
        out1 => S9
    );
bufg_11: ENTITY WORK.bufg
    PORT MAP (
        in1 => '0',
        out1 => S10
    );
bufg_12: ENTITY WORK.bufg
    PORT MAP (
        in1 => '0',
        out1 => S11
    );
bufg_13: ENTITY WORK.bufg
    PORT MAP (
        in1 => '0',
        out1 => S12
    );
bufg_14: ENTITY WORK.bufg
    PORT MAP (
        in1 => '0',
        out1 => S13
    );
bufg_15: ENTITY WORK.bufg
    PORT MAP (
        in1 => '0',
        out1 => S14
    );
bufg_16: ENTITY WORK.bufg
    PORT MAP (
        in1 => '0',
        out1 => S15
    );
bufg_17: ENTITY WORK.bufg
    PORT MAP (
        in1 => '0',
        out1 => S16
    );
bufg_18: ENTITY WORK.bufg
    PORT MAP (
        in1 => '0',
        out1 => S17
    );
bufg_19: ENTITY WORK.bufg
    PORT MAP (
        in1 => '0',
        out1 => S18
    );
bufg_20: ENTITY WORK.bufg
    PORT MAP (
        in1 => '0',
        out1 => S19
    );
bufg_21: ENTITY WORK.bufg
    PORT MAP (
        in1 => '0',
        out1 => S20
    );
bufg_22: ENTITY WORK.bufg
    PORT MAP (
        in1 => '0',
        out1 => S21
    );
bufg_23: ENTITY WORK.bufg
    PORT MAP (
        in1 => '0',
        out1 => S22
    );
bufg_24: ENTITY WORK.bufg
    PORT MAP (
        in1 => '0',
        out1 => S23
    );
bufg_25: ENTITY WORK.bufg
    PORT MAP (
        in1 => '0',
        out1 => S24
    );
bufg_26: ENTITY WORK.bufg
    PORT MAP (
        in1 => '0',
        out1 => S25
    );
bufg_27: ENTITY WORK.bufg
    PORT MAP (
        in1 => '0',
        out1 => S26
    );
bufg_28: ENTITY WORK.bufg
    PORT MAP (
        in1 => '0',
        out1 => S27
    );
bufg_29: ENTITY WORK.bufg
    PORT MAP (
        in1 => '0',
        out1 => S28
    );
bufg_30: ENTITY WORK.bufg
    PORT MAP (
        in1 => '0',
        out1 => S29
    );
bufg_31: ENTITY WORK.bufg
    PORT MAP (
        in1 => '0',
        out1 => S30
    );
bufg_32: ENTITY WORK.bufg
    PORT MAP (
        in1 => '0',
        out1 => S31
    );
bufg_33: ENTITY WORK.bufg
    PORT MAP (
        in1 => '0',
        out1 => S32
    );
bufg_34: ENTITY WORK.bufg
    PORT MAP (
        in1 => '0',
        out1 => S33
    );
bufg_35: ENTITY WORK.bufg
    PORT MAP (
        in1 => '0',
        out1 => S34
    );
bufg_36: ENTITY WORK.bufg
    PORT MAP (
        in1 => '0',
        out1 => S35
    );
bufg_37: ENTITY WORK.bufg
    PORT MAP (
        in1 => '0',
        out1 => S36
    );
bufg_38: ENTITY WORK.bufg
    PORT MAP (
        in1 => '0',
        out1 => S37
    );
nand_n_1: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S130,
        in1(1) => S129,
        out1 => S131
    );
nor_n_1: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S70,
        in1(1) => CU_ldIR,
        out1 => S132
    );
nand_n_2: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S132,
        in1(1) => S131,
        out1 => CU_readMEM
    );
nor_n_2: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S129,
        in1(1) => CU_selIN_MEM,
        out1 => S133
    );
notg_1: ENTITY WORK.notg
    PORT MAP (
        in1 => S133,
        out1 => CU_conOF
    );
nor_n_3: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S240,
        in1(1) => CU_inst_13,
        out1 => S134
    );
notg_2: ENTITY WORK.notg
    PORT MAP (
        in1 => S134,
        out1 => S135
    );
nor_n_4: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S135,
        in1(1) => CU_inst_12,
        out1 => S136
    );
nor_n_5: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S136,
        in1(1) => S133,
        out1 => CU_selIR_ADR
    );
nor_n_6: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => CU_inst_14,
        in1(1) => S220,
        out1 => S137
    );
nand_n_3: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S50,
        in1(1) => CU_inst_12,
        out1 => S138
    );
nor_n_7: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S138,
        in1(1) => CU_inst_13,
        out1 => S139
    );
nor_n_8: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S134,
        in1(1) => S120,
        out1 => S140
    );
nor_n_9: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S134,
        in1(1) => S121,
        out1 => S141
    );
nor_n_10: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S139,
        in1(1) => S124,
        out1 => S142
    );
nand_n_4: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S142,
        in1(1) => S141,
        out1 => S143
    );
nand_n_5: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S106,
        in1(1) => S74,
        out1 => S144
    );
nand_n_6: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S144,
        in1(1) => S60,
        out1 => S145
    );
nand_n_7: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S65,
        in1(1) => S238,
        out1 => S146
    );
nor_n_11: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S146,
        in1(1) => S143,
        out1 => S147
    );
nand_n_8: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S147,
        in1(1) => S145,
        out1 => S148
    );
nand_n_9: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S148,
        in1(1) => S235,
        out1 => CU_seldataBus
    );
nand_n_10: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S68,
        in1(1) => S230,
        out1 => S149
    );
nor_n_12: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S92,
        in1(1) => CU_inst_1,
        out1 => S150
    );
notg_3: ENTITY WORK.notg
    PORT MAP (
        in1 => S150,
        out1 => S151
    );
nand_n_11: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S150,
        in1(1) => S100,
        out1 => S152
    );
nor_n_13: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S88,
        in1(1) => S245,
        out1 => S153
    );
nand_n_12: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S89,
        in1(1) => S244,
        out1 => S154
    );
nand_n_13: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S153,
        in1(1) => S152,
        out1 => S155
    );
nor_n_14: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => CU_inst_9,
        in1(1) => S224,
        out1 => S156
    );
nor_n_15: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S44,
        in1(1) => S229,
        out1 => S157
    );
nand_n_14: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S156,
        in1(1) => CU_enSKP,
        out1 => S158
    );
nor_n_16: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S158,
        in1(1) => S44,
        out1 => S159
    );
nand_n_15: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S157,
        in1(1) => S156,
        out1 => S160
    );
nand_n_16: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S88,
        in1(1) => S244,
        out1 => S161
    );
nor_n_17: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S161,
        in1(1) => S159,
        out1 => S162
    );
nand_n_17: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S60,
        in1(1) => CU_inst_14,
        out1 => S163
    );
nand_n_18: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S163,
        in1(1) => S64,
        out1 => S164
    );
nand_n_19: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S164,
        in1(1) => S49,
        out1 => S165
    );
nor_n_18: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S165,
        in1(1) => S162,
        out1 => S166
    );
nand_n_20: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S166,
        in1(1) => S155,
        out1 => S167
    );
nand_n_21: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S167,
        in1(1) => S238,
        out1 => S168
    );
nand_n_22: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S168,
        in1(1) => S149,
        out1 => CU_INC1
    );
nand_n_23: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S113,
        in1(1) => S71,
        out1 => CU_selARU_SR
    );
nor_n_19: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S154,
        in1(1) => S152,
        out1 => S169
    );
notg_4: ENTITY WORK.notg
    PORT MAP (
        in1 => S169,
        out1 => S170
    );
nand_n_24: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S135,
        in1(1) => S238,
        out1 => S171
    );
nor_n_20: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S171,
        in1(1) => S169,
        out1 => S172
    );
nand_n_25: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S172,
        in1(1) => S67,
        out1 => S173
    );
nand_n_26: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S173,
        in1(1) => S149,
        out1 => CU_selINC_PC
    );
nand_n_27: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S149,
        in1(1) => S146,
        out1 => CU_ldPC
    );
nand_n_28: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S84,
        in1(1) => CU_inst_2,
        out1 => S174
    );
nor_n_21: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S174,
        in1(1) => S88,
        out1 => S175
    );
nand_n_29: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S175,
        in1(1) => S150,
        out1 => S176
    );
nand_n_30: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S176,
        in1(1) => S244,
        out1 => S177
    );
notg_5: ENTITY WORK.notg
    PORT MAP (
        in1 => S177,
        out1 => S178
    );
nand_n_31: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S140,
        in1(1) => S67,
        out1 => S179
    );
nor_n_22: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S179,
        in1(1) => S239,
        out1 => S180
    );
nand_n_32: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S138,
        in1(1) => S106,
        out1 => S181
    );
nand_n_33: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S177,
        in1(1) => S138,
        out1 => S182
    );
nor_n_23: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S182,
        in1(1) => S107,
        out1 => S183
    );
nand_n_34: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S183,
        in1(1) => S180,
        out1 => S184
    );
nand_n_35: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S184,
        in1(1) => S71,
        out1 => CU_selARU_AC
    );
nor_n_24: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S69,
        in1(1) => CU_inst_15,
        out1 => S185
    );
notg_6: ENTITY WORK.notg
    PORT MAP (
        in1 => S185,
        out1 => S186
    );
nand_n_36: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S139,
        in1(1) => S238,
        out1 => S187
    );
nand_n_37: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S187,
        in1(1) => S186,
        out1 => CU_selMEM_AC
    );
nand_n_38: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S47,
        in1(1) => S42,
        out1 => S188
    );
nor_n_25: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S188,
        in1(1) => S102,
        out1 => S189
    );
nand_n_39: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S189,
        in1(1) => S178,
        out1 => S190
    );
nand_n_40: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S134,
        in1(1) => CU_inst_12,
        out1 => S191
    );
nand_n_41: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S191,
        in1(1) => S130,
        out1 => S192
    );
nor_n_26: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S192,
        in1(1) => S146,
        out1 => S193
    );
nand_n_42: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S193,
        in1(1) => S190,
        out1 => S194
    );
nand_n_43: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S194,
        in1(1) => S69,
        out1 => CU_ldAC
    );
nand_n_44: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S144,
        in1(1) => S122,
        out1 => S195
    );
nand_n_45: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S195,
        in1(1) => S71,
        out1 => CU_selMEM_LGU
    );
nand_n_46: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S73,
        in1(1) => S242,
        out1 => S196
    );
nor_n_27: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S181,
        in1(1) => S239,
        out1 => S197
    );
nand_n_47: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S196,
        in1(1) => S177,
        out1 => S198
    );
nor_n_28: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S198,
        in1(1) => S179,
        out1 => S199
    );
nand_n_48: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S199,
        in1(1) => S197,
        out1 => S200
    );
nand_n_49: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S200,
        in1(1) => S71,
        out1 => CU_ADD
    );
nor_n_29: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S137,
        in1(1) => S75,
        out1 => S201
    );
nand_n_50: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S201,
        in1(1) => S180,
        out1 => S202
    );
nand_n_51: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S98,
        in1(1) => S244,
        out1 => S203
    );
nor_n_30: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S203,
        in1(1) => S102,
        out1 => S204
    );
nor_n_31: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S204,
        in1(1) => S202,
        out1 => CU_selLGU_SR
    );
nor_n_32: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S160,
        in1(1) => S40,
        out1 => CU_INC2
    );
nor_n_33: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S63,
        in1(1) => S55,
        out1 => S205
    );
nand_n_52: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S69,
        in1(1) => S56,
        out1 => CU_selIN_ADR
    );
nand_n_53: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S156,
        in1(1) => S41,
        out1 => S206
    );
notg_7: ENTITY WORK.notg
    PORT MAP (
        in1 => S206,
        out1 => CU_selIMM_OF
    );
nand_n_54: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S87,
        in1(1) => S238,
        out1 => S207
    );
nor_n_34: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S207,
        in1(1) => S151,
        out1 => S208
    );
nand_n_55: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S208,
        in1(1) => S153,
        out1 => S209
    );
notg_8: ENTITY WORK.notg
    PORT MAP (
        in1 => S209,
        out1 => CU_selPC_OF
    );
nand_n_56: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S209,
        in1(1) => S206,
        out1 => CU_ldOF
    );
nor_n_35: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S205,
        in1(1) => S239,
        out1 => CU_selMEM_IN
    );
nor_n_36: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S123,
        in1(1) => S234,
        out1 => CU_selINC_IN
    );
nor_n_37: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S170,
        in1(1) => S239,
        out1 => CU_LSB0E
    );
nor_n_38: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S169,
        in1(1) => S58,
        out1 => S210
    );
nor_n_39: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S210,
        in1(1) => S239,
        out1 => CU_selIMM_PC
    );
nor_n_40: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S135,
        in1(1) => S123,
        out1 => CU_selMEM_PC
    );
nand_n_57: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S189,
        in1(1) => S244,
        out1 => S211
    );
notg_9: ENTITY WORK.notg
    PORT MAP (
        in1 => S211,
        out1 => S212
    );
nor_n_41: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S212,
        in1(1) => S202,
        out1 => CU_selLGU_AC
    );
nor_n_42: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S119,
        in1(1) => S239,
        out1 => CU_selIMM_AC
    );
nor_n_43: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S188,
        in1(1) => S245,
        out1 => S213
    );
nor_n_44: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S137,
        in1(1) => S48,
        out1 => S214
    );
nand_n_58: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S214,
        in1(1) => S180,
        out1 => S215
    );
nor_n_45: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S215,
        in1(1) => S213,
        out1 => CU_selIMM_LGU
    );
nor_n_46: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S176,
        in1(1) => S40,
        out1 => CU_sel1_ARU
    );
nand_n_59: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S214,
        in1(1) => S240,
        out1 => S216
    );
nor_n_47: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S216,
        in1(1) => S146,
        out1 => CU_SE4bits
    );
nand_n_60: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S188,
        in1(1) => S39,
        out1 => S217
    );
nand_n_61: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S217,
        in1(1) => S206,
        out1 => CU_SE12bits
    );
nor_n_48: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S196,
        in1(1) => S239,
        out1 => CU_MUL
    );
notg_10: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_pstate_0,
        out1 => S218
    );
notg_11: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_pstate_1,
        out1 => S219
    );
notg_12: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_inst_12,
        out1 => S220
    );
notg_13: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_inst_13,
        out1 => S221
    );
notg_14: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_inst_14,
        out1 => S222
    );
notg_15: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_inst_15,
        out1 => S223
    );
notg_16: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_inst_8,
        out1 => S224
    );
notg_17: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_inst_11,
        out1 => S225
    );
notg_18: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_rst,
        out1 => S226
    );
notg_19: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_inst_1,
        out1 => S227
    );
notg_20: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_inst_3,
        out1 => S228
    );
notg_21: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_enSKP,
        out1 => S229
    );
nor_n_49: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => CU_pstate_1,
        in1(1) => CU_pstate_0,
        out1 => CU_ldIR
    );
nor_n_50: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S219,
        in1(1) => CU_pstate_0,
        out1 => S230
    );
nor_n_51: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => CU_inst_15,
        in1(1) => S222,
        out1 => S231
    );
nand_n_62: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S223,
        in1(1) => CU_inst_14,
        out1 => S232
    );
nor_n_52: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S232,
        in1(1) => CU_inst_13,
        out1 => S233
    );
nand_n_63: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S231,
        in1(1) => S221,
        out1 => S234
    );
nand_n_64: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S233,
        in1(1) => S230,
        out1 => S235
    );
nor_n_53: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S235,
        in1(1) => S220,
        out1 => CU_selIN_MEM
    );
nor_n_54: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => CU_inst_10,
        in1(1) => CU_inst_11,
        out1 => S236
    );
notg_22: ENTITY WORK.notg
    PORT MAP (
        in1 => S236,
        out1 => S237
    );
nor_n_55: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => CU_pstate_1,
        in1(1) => S218,
        out1 => S238
    );
nand_n_65: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S219,
        in1(1) => CU_pstate_0,
        out1 => S239
    );
nand_n_66: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_inst_15,
        in1(1) => CU_inst_14,
        out1 => S240
    );
notg_23: ENTITY WORK.notg
    PORT MAP (
        in1 => S240,
        out1 => S241
    );
nor_n_56: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S221,
        in1(1) => S220,
        out1 => S242
    );
nand_n_67: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_inst_13,
        in1(1) => CU_inst_12,
        out1 => S243
    );
nor_n_57: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S243,
        in1(1) => S240,
        out1 => S244
    );
nand_n_68: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S242,
        in1(1) => S241,
        out1 => S245
    );
nor_n_58: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S245,
        in1(1) => S239,
        out1 => S39
    );
nand_n_69: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S244,
        in1(1) => S238,
        out1 => S40
    );
nor_n_59: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S40,
        in1(1) => S237,
        out1 => S41
    );
nand_n_70: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S236,
        in1(1) => CU_inst_9,
        out1 => S42
    );
nand_n_71: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S39,
        in1(1) => CU_inst_8,
        out1 => S43
    );
nor_n_60: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S43,
        in1(1) => S42,
        out1 => CU_SHF_0
    );
nand_n_72: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_inst_10,
        in1(1) => S225,
        out1 => S44
    );
notg_24: ENTITY WORK.notg
    PORT MAP (
        in1 => S44,
        out1 => S45
    );
nor_n_61: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => CU_inst_9,
        in1(1) => CU_inst_8,
        out1 => S46
    );
nand_n_73: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S46,
        in1(1) => S45,
        out1 => S47
    );
nor_n_62: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S47,
        in1(1) => S40,
        out1 => CU_SHF_1
    );
nor_n_63: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S243,
        in1(1) => CU_inst_15,
        out1 => S48
    );
nand_n_74: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S242,
        in1(1) => S223,
        out1 => S49
    );
nor_n_64: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => CU_inst_15,
        in1(1) => CU_inst_14,
        out1 => S50
    );
nor_n_65: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S49,
        in1(1) => CU_inst_14,
        out1 => S51
    );
nand_n_75: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S51,
        in1(1) => S238,
        out1 => S52
    );
nor_n_66: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => CU_inst_13,
        in1(1) => CU_inst_12,
        out1 => S53
    );
nand_n_76: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S221,
        in1(1) => S220,
        out1 => S54
    );
nor_n_67: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S54,
        in1(1) => S232,
        out1 => S55
    );
nand_n_77: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S55,
        in1(1) => S230,
        out1 => S56
    );
nand_n_78: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S56,
        in1(1) => S52,
        out1 => CU_selAC_MEM
    );
nand_n_79: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S239,
        in1(1) => S226,
        out1 => S57
    );
nor_n_68: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S57,
        in1(1) => S230,
        out1 => S246
    );
nor_n_69: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S240,
        in1(1) => CU_inst_12,
        out1 => S58
    );
nor_n_70: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S221,
        in1(1) => CU_inst_12,
        out1 => S59
    );
nand_n_80: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_inst_13,
        in1(1) => S220,
        out1 => S60
    );
nand_n_81: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S58,
        in1(1) => CU_inst_13,
        out1 => S61
    );
notg_25: ENTITY WORK.notg
    PORT MAP (
        in1 => S61,
        out1 => S62
    );
nor_n_71: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S61,
        in1(1) => S239,
        out1 => CU_selPC_MEM
    );
nor_n_72: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S60,
        in1(1) => CU_inst_14,
        out1 => S63
    );
nand_n_82: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S59,
        in1(1) => S222,
        out1 => S64
    );
nor_n_73: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S63,
        in1(1) => S233,
        out1 => S65
    );
nand_n_83: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S64,
        in1(1) => S234,
        out1 => S66
    );
nor_n_74: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S65,
        in1(1) => S239,
        out1 => CU_ldIN
    );
nor_n_75: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S66,
        in1(1) => S62,
        out1 => S67
    );
nand_n_84: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S65,
        in1(1) => S61,
        out1 => S68
    );
nor_n_76: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S67,
        in1(1) => S239,
        out1 => S247
    );
nand_n_85: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S63,
        in1(1) => S230,
        out1 => S69
    );
notg_26: ENTITY WORK.notg
    PORT MAP (
        in1 => S69,
        out1 => S70
    );
nand_n_86: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S70,
        in1(1) => CU_inst_15,
        out1 => S71
    );
notg_27: ENTITY WORK.notg
    PORT MAP (
        in1 => S71,
        out1 => S72
    );
nor_n_77: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S223,
        in1(1) => CU_inst_14,
        out1 => S73
    );
nand_n_87: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_inst_15,
        in1(1) => S222,
        out1 => S74
    );
nor_n_78: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S74,
        in1(1) => CU_inst_13,
        out1 => S75
    );
notg_28: ENTITY WORK.notg
    PORT MAP (
        in1 => S75,
        out1 => S76
    );
nor_n_79: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S76,
        in1(1) => S239,
        out1 => S77
    );
nand_n_88: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S75,
        in1(1) => S238,
        out1 => S78
    );
nor_n_80: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S77,
        in1(1) => S72,
        out1 => S79
    );
nor_n_81: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S44,
        in1(1) => CU_inst_8,
        out1 => S80
    );
nand_n_89: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S80,
        in1(1) => CU_inst_9,
        out1 => S81
    );
nor_n_82: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S81,
        in1(1) => S40,
        out1 => CU_selSET_SR
    );
nand_n_90: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_selSET_SR,
        in1(1) => CU_inst_4,
        out1 => S82
    );
nand_n_91: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S82,
        in1(1) => S79,
        out1 => CU_ldSR_0
    );
nand_n_92: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_selSET_SR,
        in1(1) => CU_inst_5,
        out1 => S83
    );
nand_n_93: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S83,
        in1(1) => S79,
        out1 => CU_ldSR_1
    );
nor_n_83: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => CU_inst_3,
        in1(1) => CU_inst_0,
        out1 => S84
    );
notg_29: ENTITY WORK.notg
    PORT MAP (
        in1 => S84,
        out1 => S85
    );
nor_n_84: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => CU_inst_2,
        in1(1) => CU_inst_3,
        out1 => S86
    );
nor_n_85: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S85,
        in1(1) => CU_inst_2,
        out1 => S87
    );
nand_n_94: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S46,
        in1(1) => S236,
        out1 => S88
    );
notg_30: ENTITY WORK.notg
    PORT MAP (
        in1 => S88,
        out1 => S89
    );
nor_n_86: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => CU_inst_5,
        in1(1) => CU_inst_4,
        out1 => S90
    );
nor_n_87: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => CU_inst_7,
        in1(1) => CU_inst_6,
        out1 => S91
    );
nand_n_95: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S91,
        in1(1) => S90,
        out1 => S92
    );
notg_31: ENTITY WORK.notg
    PORT MAP (
        in1 => S92,
        out1 => S93
    );
nor_n_88: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S92,
        in1(1) => S227,
        out1 => S94
    );
nand_n_96: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S93,
        in1(1) => CU_inst_1,
        out1 => S95
    );
nor_n_89: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S95,
        in1(1) => S88,
        out1 => S96
    );
nand_n_97: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S94,
        in1(1) => S89,
        out1 => S97
    );
nand_n_98: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S96,
        in1(1) => S87,
        out1 => S98
    );
nor_n_90: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S98,
        in1(1) => S40,
        out1 => CU_zeroAC
    );
nand_n_99: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S228,
        in1(1) => CU_inst_0,
        out1 => S99
    );
nor_n_91: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S99,
        in1(1) => CU_inst_2,
        out1 => S100
    );
nand_n_100: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S86,
        in1(1) => CU_inst_0,
        out1 => S101
    );
nor_n_92: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S101,
        in1(1) => S97,
        out1 => S102
    );
nand_n_101: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S102,
        in1(1) => S39,
        out1 => S103
    );
notg_32: ENTITY WORK.notg
    PORT MAP (
        in1 => S103,
        out1 => CU_NOT
    );
nand_n_102: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S103,
        in1(1) => S71,
        out1 => S104
    );
nor_n_93: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S104,
        in1(1) => CU_zeroAC,
        out1 => S105
    );
nand_n_103: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S231,
        in1(1) => CU_inst_13,
        out1 => S106
    );
notg_33: ENTITY WORK.notg
    PORT MAP (
        in1 => S106,
        out1 => S107
    );
nor_n_94: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S106,
        in1(1) => S239,
        out1 => CU_AND
    );
notg_34: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_AND,
        out1 => S108
    );
nand_n_104: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_selSET_SR,
        in1(1) => CU_inst_6,
        out1 => S109
    );
nand_n_105: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S109,
        in1(1) => S78,
        out1 => S110
    );
nor_n_95: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S110,
        in1(1) => CU_AND,
        out1 => S111
    );
nand_n_106: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S111,
        in1(1) => S105,
        out1 => CU_ldSR_2
    );
nor_n_96: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S74,
        in1(1) => S59,
        out1 => S112
    );
nand_n_107: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S112,
        in1(1) => S238,
        out1 => S113
    );
nand_n_108: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S113,
        in1(1) => S108,
        out1 => S114
    );
nand_n_109: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_selSET_SR,
        in1(1) => CU_inst_7,
        out1 => S115
    );
notg_35: ENTITY WORK.notg
    PORT MAP (
        in1 => S115,
        out1 => S116
    );
nor_n_97: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S116,
        in1(1) => S114,
        out1 => S117
    );
nand_n_110: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S117,
        in1(1) => S105,
        out1 => CU_ldSR_3
    );
nand_n_111: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_pstate_1,
        in1(1) => CU_pstate_0,
        out1 => S118
    );
notg_36: ENTITY WORK.notg
    PORT MAP (
        in1 => S118,
        out1 => S38
    );
nand_n_112: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S53,
        in1(1) => S50,
        out1 => S119
    );
notg_37: ENTITY WORK.notg
    PORT MAP (
        in1 => S119,
        out1 => S120
    );
nand_n_113: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S119,
        in1(1) => S245,
        out1 => S121
    );
nor_n_98: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S239,
        in1(1) => S220,
        out1 => S122
    );
nand_n_114: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S238,
        in1(1) => CU_inst_12,
        out1 => S123
    );
nor_n_99: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S60,
        in1(1) => S232,
        out1 => S124
    );
nor_n_100: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S74,
        in1(1) => S54,
        out1 => S125
    );
nor_n_101: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S125,
        in1(1) => S124,
        out1 => S126
    );
nor_n_102: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S121,
        in1(1) => S239,
        out1 => S127
    );
nand_n_115: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S127,
        in1(1) => S126,
        out1 => S128
    );
notg_38: ENTITY WORK.notg
    PORT MAP (
        in1 => S128,
        out1 => S129
    );
nor_n_103: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S58,
        in1(1) => S51,
        out1 => S130
    );
$_DLATCH_N__1: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S246,
        E => S38,
        Q => CU_nstate_0
    );
$_DLATCH_N__2: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S247,
        E => S38,
        Q => CU_nstate_1
    );
dff_1: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => CU_nstate_0,
        NbarT => '0',
        PRE => '0',
        Q => CU_pstate_0,
        Si => S3365,
        global_reset => '0'
    );
dff_2: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => CU_nstate_1,
        NbarT => '0',
        PRE => '0',
        Q => CU_pstate_1,
        Si => S3366,
        global_reset => '0'
    );
notg_39: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_SR_V_out,
        out1 => S248
    );
notg_40: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_SR_C_out,
        out1 => S249
    );
notg_41: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_SR_N_out,
        out1 => S250
    );
notg_42: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_SR_Z_out,
        out1 => S251
    );
nor_n_104: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S250,
        in1(1) => CU_inst_2,
        out1 => S252
    );
nand_n_116: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S250,
        in1(1) => CU_inst_2,
        out1 => S253
    );
nand_n_117: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S253,
        in1(1) => CU_inst_6,
        out1 => S254
    );
nor_n_105: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S254,
        in1(1) => S252,
        out1 => S255
    );
nor_n_106: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S251,
        in1(1) => CU_inst_3,
        out1 => S256
    );
nand_n_118: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S251,
        in1(1) => CU_inst_3,
        out1 => S257
    );
nand_n_119: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S257,
        in1(1) => CU_inst_7,
        out1 => S258
    );
nor_n_107: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S258,
        in1(1) => S256,
        out1 => S259
    );
nor_n_108: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S259,
        in1(1) => S255,
        out1 => S260
    );
nor_n_109: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S248,
        in1(1) => CU_inst_0,
        out1 => S261
    );
nand_n_120: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S248,
        in1(1) => CU_inst_0,
        out1 => S262
    );
nand_n_121: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S262,
        in1(1) => CU_inst_4,
        out1 => S263
    );
nor_n_110: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S263,
        in1(1) => S261,
        out1 => S264
    );
nor_n_111: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S249,
        in1(1) => CU_inst_1,
        out1 => S265
    );
nand_n_122: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S249,
        in1(1) => CU_inst_1,
        out1 => S266
    );
nand_n_123: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S266,
        in1(1) => CU_inst_5,
        out1 => S267
    );
nor_n_112: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S267,
        in1(1) => S265,
        out1 => S268
    );
nor_n_113: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S268,
        in1(1) => S264,
        out1 => S269
    );
nand_n_124: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S269,
        in1(1) => S260,
        out1 => CU_enSKP
    );
notg_43: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_ldAC,
        out1 => S287
    );
nor_n_114: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => CU_ldAC,
        in1(1) => CU_zeroAC,
        out1 => S288
    );
nand_n_125: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S288,
        in1(1) => DP_AC_out_0,
        out1 => S289
    );
nor_n_115: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S287,
        in1(1) => CU_zeroAC,
        out1 => S290
    );
nand_n_126: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S290,
        in1(1) => DP_AC_in_0,
        out1 => S291
    );
nand_n_127: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S291,
        in1(1) => S289,
        out1 => S270
    );
nand_n_128: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S288,
        in1(1) => DP_AC_out_1,
        out1 => S292
    );
nand_n_129: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S290,
        in1(1) => DP_AC_in_1,
        out1 => S293
    );
nand_n_130: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S293,
        in1(1) => S292,
        out1 => S271
    );
nand_n_131: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S288,
        in1(1) => DP_AC_out_2,
        out1 => S294
    );
nand_n_132: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S290,
        in1(1) => DP_AC_in_2,
        out1 => S295
    );
nand_n_133: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S295,
        in1(1) => S294,
        out1 => S272
    );
nand_n_134: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S288,
        in1(1) => DP_AC_out_3,
        out1 => S296
    );
nand_n_135: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S290,
        in1(1) => DP_AC_in_3,
        out1 => S297
    );
nand_n_136: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S297,
        in1(1) => S296,
        out1 => S273
    );
nand_n_137: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S288,
        in1(1) => DP_AC_out_4,
        out1 => S298
    );
nand_n_138: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S290,
        in1(1) => DP_AC_in_4,
        out1 => S299
    );
nand_n_139: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S299,
        in1(1) => S298,
        out1 => S274
    );
nand_n_140: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S288,
        in1(1) => DP_AC_out_5,
        out1 => S300
    );
nand_n_141: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S290,
        in1(1) => DP_AC_in_5,
        out1 => S301
    );
nand_n_142: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S301,
        in1(1) => S300,
        out1 => S275
    );
nand_n_143: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S288,
        in1(1) => DP_AC_out_6,
        out1 => S302
    );
nand_n_144: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S290,
        in1(1) => DP_AC_in_6,
        out1 => S303
    );
nand_n_145: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S303,
        in1(1) => S302,
        out1 => S276
    );
nand_n_146: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S288,
        in1(1) => DP_AC_out_7,
        out1 => S304
    );
nand_n_147: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S290,
        in1(1) => DP_AC_in_7,
        out1 => S305
    );
nand_n_148: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S305,
        in1(1) => S304,
        out1 => S277
    );
nand_n_149: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S288,
        in1(1) => DP_AC_out_8,
        out1 => S306
    );
nand_n_150: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S290,
        in1(1) => DP_AC_in_8,
        out1 => S307
    );
nand_n_151: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S307,
        in1(1) => S306,
        out1 => S278
    );
nand_n_152: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S288,
        in1(1) => DP_AC_out_9,
        out1 => S308
    );
nand_n_153: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S290,
        in1(1) => DP_AC_in_9,
        out1 => S309
    );
nand_n_154: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S309,
        in1(1) => S308,
        out1 => S279
    );
nand_n_155: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S288,
        in1(1) => DP_AC_out_10,
        out1 => S310
    );
nand_n_156: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S290,
        in1(1) => DP_AC_in_10,
        out1 => S311
    );
nand_n_157: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S311,
        in1(1) => S310,
        out1 => S280
    );
nand_n_158: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S288,
        in1(1) => DP_AC_out_11,
        out1 => S312
    );
nand_n_159: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S290,
        in1(1) => DP_AC_in_11,
        out1 => S313
    );
nand_n_160: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S313,
        in1(1) => S312,
        out1 => S281
    );
nand_n_161: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S288,
        in1(1) => DP_AC_out_12,
        out1 => S314
    );
nand_n_162: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S290,
        in1(1) => DP_AC_in_12,
        out1 => S315
    );
nand_n_163: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S315,
        in1(1) => S314,
        out1 => S282
    );
nand_n_164: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S288,
        in1(1) => DP_AC_out_13,
        out1 => S316
    );
nand_n_165: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S290,
        in1(1) => DP_AC_in_13,
        out1 => S317
    );
nand_n_166: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S317,
        in1(1) => S316,
        out1 => S283
    );
nand_n_167: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S288,
        in1(1) => DP_AC_out_14,
        out1 => S318
    );
nand_n_168: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S290,
        in1(1) => DP_AC_in_14,
        out1 => S319
    );
nand_n_169: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S319,
        in1(1) => S318,
        out1 => S284
    );
nand_n_170: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S288,
        in1(1) => DP_AC_out_15,
        out1 => S320
    );
nand_n_171: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S290,
        in1(1) => DP_AC_in_15,
        out1 => S286
    );
nand_n_172: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S286,
        in1(1) => S320,
        out1 => S285
    );
dff_3: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S270,
        NbarT => '0',
        PRE => '0',
        Q => DP_AC_out_0,
        Si => S3307,
        global_reset => '0'
    );
dff_4: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S271,
        NbarT => '0',
        PRE => '0',
        Q => DP_AC_out_1,
        Si => S3306,
        global_reset => '0'
    );
dff_5: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S272,
        NbarT => '0',
        PRE => '0',
        Q => DP_AC_out_2,
        Si => S3305,
        global_reset => '0'
    );
dff_6: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S273,
        NbarT => '0',
        PRE => '0',
        Q => DP_AC_out_3,
        Si => S3304,
        global_reset => '0'
    );
dff_7: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S274,
        NbarT => '0',
        PRE => '0',
        Q => DP_AC_out_4,
        Si => S3303,
        global_reset => '0'
    );
dff_8: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S275,
        NbarT => '0',
        PRE => '0',
        Q => DP_AC_out_5,
        Si => S3302,
        global_reset => '0'
    );
dff_9: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S276,
        NbarT => '0',
        PRE => '0',
        Q => DP_AC_out_6,
        Si => S3301,
        global_reset => '0'
    );
dff_10: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S277,
        NbarT => '0',
        PRE => '0',
        Q => DP_AC_out_7,
        Si => S3300,
        global_reset => '0'
    );
dff_11: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S278,
        NbarT => '0',
        PRE => '0',
        Q => DP_AC_out_8,
        Si => S3299,
        global_reset => '0'
    );
dff_12: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S279,
        NbarT => '0',
        PRE => '0',
        Q => DP_AC_out_9,
        Si => S3298,
        global_reset => '0'
    );
dff_13: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S280,
        NbarT => '0',
        PRE => '0',
        Q => DP_AC_out_10,
        Si => S3297,
        global_reset => '0'
    );
dff_14: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S281,
        NbarT => '0',
        PRE => '0',
        Q => DP_AC_out_11,
        Si => S3296,
        global_reset => '0'
    );
dff_15: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S282,
        NbarT => '0',
        PRE => '0',
        Q => DP_AC_out_12,
        Si => S3295,
        global_reset => '0'
    );
dff_16: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S283,
        NbarT => '0',
        PRE => '0',
        Q => DP_AC_out_13,
        Si => S3294,
        global_reset => '0'
    );
dff_17: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S284,
        NbarT => '0',
        PRE => '0',
        Q => DP_AC_out_14,
        Si => S3293,
        global_reset => '0'
    );
dff_18: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S285,
        NbarT => '0',
        PRE => '0',
        Q => DP_AC_out_15,
        Si => S3356,
        global_reset => '0'
    );
notg_44: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_AC_out_0,
        out1 => S966
    );
notg_45: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_ARU1_in1_0,
        out1 => S977
    );
notg_46: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_ADD,
        out1 => S988
    );
notg_47: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_AC_out_1,
        out1 => S998
    );
notg_48: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_ARU1_in1_1,
        out1 => S1009
    );
notg_49: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_AC_out_2,
        out1 => S1020
    );
notg_50: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_ARU1_in1_2,
        out1 => S1031
    );
notg_51: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_AC_out_3,
        out1 => S1042
    );
notg_52: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_ARU1_in1_3,
        out1 => S1053
    );
notg_53: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_AC_out_4,
        out1 => S1064
    );
notg_54: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_ARU1_in1_4,
        out1 => S1075
    );
notg_55: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_AC_out_5,
        out1 => S1085
    );
notg_56: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_ARU1_in1_5,
        out1 => S1096
    );
notg_57: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_AC_out_6,
        out1 => S1107
    );
notg_58: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_ARU1_in1_6,
        out1 => S1118
    );
notg_59: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_AC_out_7,
        out1 => S1129
    );
notg_60: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_ARU1_in1_7,
        out1 => S1140
    );
notg_61: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_AC_out_9,
        out1 => S1150
    );
notg_62: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_ARU1_in1_9,
        out1 => S1161
    );
notg_63: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_AC_out_11,
        out1 => S1172
    );
notg_64: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_ARU1_in1_11,
        out1 => S1183
    );
notg_65: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_AC_out_13,
        out1 => S1194
    );
notg_66: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_ARU1_in1_13,
        out1 => S1205
    );
notg_67: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_AC_out_14,
        out1 => S1215
    );
notg_68: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_ARU1_in1_14,
        out1 => S1226
    );
nor_n_116: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => DP_ARU1_out_7,
        in1(1) => DP_ARU1_out_4,
        out1 => S1237
    );
nor_n_117: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => DP_ARU1_out_2,
        in1(1) => DP_ARU1_out_1,
        out1 => S1248
    );
nand_n_173: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1248,
        in1(1) => S1237,
        out1 => S1258
    );
nor_n_118: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => DP_ARU1_out_14,
        in1(1) => DP_ARU1_out_13,
        out1 => S1269
    );
nor_n_119: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => DP_ARU1_out_11,
        in1(1) => DP_ARU1_out_8,
        out1 => S348
    );
nand_n_174: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S348,
        in1(1) => S1269,
        out1 => S358
    );
nor_n_120: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S358,
        in1(1) => S1258,
        out1 => S359
    );
nor_n_121: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => DP_ARU1_out_6,
        in1(1) => DP_ARU1_out_5,
        out1 => S360
    );
nor_n_122: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => DP_ARU1_out_3,
        in1(1) => DP_ARU1_out_0,
        out1 => S361
    );
nand_n_175: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S361,
        in1(1) => S360,
        out1 => S362
    );
nor_n_123: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => DP_ARU1_N,
        in1(1) => DP_ARU1_out_12,
        out1 => S363
    );
nor_n_124: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => DP_ARU1_out_10,
        in1(1) => DP_ARU1_out_9,
        out1 => S364
    );
nand_n_176: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S364,
        in1(1) => S363,
        out1 => S365
    );
nor_n_125: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S365,
        in1(1) => S362,
        out1 => S366
    );
nand_n_177: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S366,
        in1(1) => S359,
        out1 => S367
    );
notg_69: ENTITY WORK.notg
    PORT MAP (
        in1 => S367,
        out1 => DP_ARU1_Z
    );
nor_n_126: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_15,
        in1(1) => DP_AC_out_15,
        out1 => S368
    );
nand_n_178: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S368,
        in1(1) => DP_ARU1_N,
        out1 => S369
    );
nand_n_179: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_15,
        in1(1) => DP_AC_out_15,
        out1 => S370
    );
notg_70: ENTITY WORK.notg
    PORT MAP (
        in1 => S370,
        out1 => S371
    );
nor_n_127: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S370,
        in1(1) => DP_ARU1_N,
        out1 => S372
    );
notg_71: ENTITY WORK.notg
    PORT MAP (
        in1 => S372,
        out1 => S373
    );
nand_n_180: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S373,
        in1(1) => S369,
        out1 => DP_ARU1_V
    );
nor_n_128: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_0,
        in1(1) => DP_AC_out_0,
        out1 => S374
    );
nor_n_129: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S977,
        in1(1) => S966,
        out1 => S375
    );
nand_n_181: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_0,
        in1(1) => DP_AC_out_0,
        out1 => S376
    );
nor_n_130: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S376,
        in1(1) => S988,
        out1 => S377
    );
nor_n_131: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S374,
        in1(1) => S988,
        out1 => S378
    );
nor_n_132: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S378,
        in1(1) => S375,
        out1 => S379
    );
nor_n_133: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S379,
        in1(1) => S377,
        out1 => S321
    );
nor_n_134: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1009,
        in1(1) => S998,
        out1 => S380
    );
nand_n_182: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_1,
        in1(1) => DP_AC_out_1,
        out1 => S381
    );
nor_n_135: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_1,
        in1(1) => DP_AC_out_1,
        out1 => S382
    );
nor_n_136: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S382,
        in1(1) => S380,
        out1 => S383
    );
nand_n_183: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S383,
        in1(1) => S375,
        out1 => S384
    );
nor_n_137: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S383,
        in1(1) => S375,
        out1 => S385
    );
nand_n_184: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_1,
        in1(1) => DP_AC_out_0,
        out1 => S386
    );
nand_n_185: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_1,
        in1(1) => DP_ARU1_in1_0,
        out1 => S387
    );
nor_n_138: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S381,
        in1(1) => S376,
        out1 => S388
    );
nand_n_186: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S387,
        in1(1) => S386,
        out1 => S389
    );
notg_72: ENTITY WORK.notg
    PORT MAP (
        in1 => S389,
        out1 => S390
    );
nor_n_139: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S390,
        in1(1) => S388,
        out1 => S391
    );
nand_n_187: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S391,
        in1(1) => S988,
        out1 => S392
    );
nor_n_140: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S385,
        in1(1) => S988,
        out1 => S393
    );
nand_n_188: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S393,
        in1(1) => S384,
        out1 => S394
    );
nand_n_189: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S394,
        in1(1) => S392,
        out1 => S328
    );
nand_n_190: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S384,
        in1(1) => S381,
        out1 => S395
    );
nor_n_141: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_2,
        in1(1) => DP_AC_out_2,
        out1 => S396
    );
nor_n_142: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1031,
        in1(1) => S1020,
        out1 => S397
    );
nand_n_191: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_2,
        in1(1) => DP_AC_out_2,
        out1 => S398
    );
nor_n_143: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S397,
        in1(1) => S396,
        out1 => S399
    );
nor_n_144: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S399,
        in1(1) => S395,
        out1 => S400
    );
nand_n_192: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S399,
        in1(1) => S395,
        out1 => S401
    );
notg_73: ENTITY WORK.notg
    PORT MAP (
        in1 => S401,
        out1 => S402
    );
nor_n_145: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S402,
        in1(1) => S400,
        out1 => S403
    );
nand_n_193: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_2,
        in1(1) => DP_AC_out_0,
        out1 => S404
    );
nand_n_194: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_2,
        in1(1) => DP_ARU1_in1_0,
        out1 => S405
    );
nand_n_195: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_2,
        in1(1) => DP_ARU1_in1_1,
        out1 => S406
    );
notg_74: ENTITY WORK.notg
    PORT MAP (
        in1 => S406,
        out1 => S407
    );
nor_n_146: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S405,
        in1(1) => S381,
        out1 => S408
    );
notg_75: ENTITY WORK.notg
    PORT MAP (
        in1 => S408,
        out1 => S409
    );
nand_n_196: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S405,
        in1(1) => S381,
        out1 => S410
    );
nand_n_197: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S410,
        in1(1) => S409,
        out1 => S411
    );
nand_n_198: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S411,
        in1(1) => S404,
        out1 => S412
    );
notg_76: ENTITY WORK.notg
    PORT MAP (
        in1 => S412,
        out1 => S413
    );
nor_n_147: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S411,
        in1(1) => S404,
        out1 => S414
    );
nor_n_148: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S414,
        in1(1) => S413,
        out1 => S415
    );
nand_n_199: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S415,
        in1(1) => S388,
        out1 => S416
    );
nor_n_149: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S415,
        in1(1) => S388,
        out1 => S417
    );
nor_n_150: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S417,
        in1(1) => CU_ADD,
        out1 => S418
    );
nand_n_200: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S418,
        in1(1) => S416,
        out1 => S419
    );
nand_n_201: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S403,
        in1(1) => CU_ADD,
        out1 => S420
    );
nand_n_202: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S420,
        in1(1) => S419,
        out1 => S329
    );
nand_n_203: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S401,
        in1(1) => S398,
        out1 => S421
    );
nor_n_151: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_3,
        in1(1) => DP_AC_out_3,
        out1 => S422
    );
nor_n_152: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1053,
        in1(1) => S1042,
        out1 => S423
    );
nand_n_204: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_3,
        in1(1) => DP_AC_out_3,
        out1 => S424
    );
nor_n_153: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S423,
        in1(1) => S422,
        out1 => S425
    );
nand_n_205: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S425,
        in1(1) => S421,
        out1 => S426
    );
notg_77: ENTITY WORK.notg
    PORT MAP (
        in1 => S426,
        out1 => S427
    );
nor_n_154: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S425,
        in1(1) => S421,
        out1 => S428
    );
nor_n_155: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S428,
        in1(1) => S427,
        out1 => S429
    );
nand_n_206: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S429,
        in1(1) => CU_ADD,
        out1 => S430
    );
nand_n_207: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_3,
        in1(1) => DP_AC_out_0,
        out1 => S431
    );
notg_78: ENTITY WORK.notg
    PORT MAP (
        in1 => S431,
        out1 => S432
    );
nor_n_156: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S414,
        in1(1) => S408,
        out1 => S433
    );
notg_79: ENTITY WORK.notg
    PORT MAP (
        in1 => S433,
        out1 => S434
    );
nand_n_208: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_2,
        in1(1) => DP_AC_out_1,
        out1 => S435
    );
notg_80: ENTITY WORK.notg
    PORT MAP (
        in1 => S435,
        out1 => S436
    );
nand_n_209: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_3,
        in1(1) => DP_ARU1_in1_0,
        out1 => S437
    );
notg_81: ENTITY WORK.notg
    PORT MAP (
        in1 => S437,
        out1 => S438
    );
nand_n_210: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_3,
        in1(1) => DP_ARU1_in1_1,
        out1 => S439
    );
nor_n_157: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S437,
        in1(1) => S406,
        out1 => S440
    );
nand_n_211: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S438,
        in1(1) => S407,
        out1 => S441
    );
nand_n_212: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S437,
        in1(1) => S406,
        out1 => S442
    );
notg_82: ENTITY WORK.notg
    PORT MAP (
        in1 => S442,
        out1 => S443
    );
nor_n_158: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S443,
        in1(1) => S440,
        out1 => S444
    );
nand_n_213: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S442,
        in1(1) => S441,
        out1 => S445
    );
nand_n_214: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S445,
        in1(1) => S435,
        out1 => S446
    );
nor_n_159: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S445,
        in1(1) => S435,
        out1 => S447
    );
nand_n_215: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S444,
        in1(1) => S436,
        out1 => S448
    );
nand_n_216: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S448,
        in1(1) => S446,
        out1 => S449
    );
notg_83: ENTITY WORK.notg
    PORT MAP (
        in1 => S449,
        out1 => S450
    );
nand_n_217: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S450,
        in1(1) => S434,
        out1 => S451
    );
notg_84: ENTITY WORK.notg
    PORT MAP (
        in1 => S451,
        out1 => S452
    );
nand_n_218: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S449,
        in1(1) => S433,
        out1 => S453
    );
nand_n_219: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S453,
        in1(1) => S451,
        out1 => S454
    );
notg_85: ENTITY WORK.notg
    PORT MAP (
        in1 => S454,
        out1 => S455
    );
nand_n_220: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S454,
        in1(1) => S431,
        out1 => S456
    );
nor_n_160: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S454,
        in1(1) => S431,
        out1 => S457
    );
nand_n_221: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S455,
        in1(1) => S432,
        out1 => S458
    );
nand_n_222: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S458,
        in1(1) => S456,
        out1 => S459
    );
nand_n_223: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S459,
        in1(1) => S416,
        out1 => S460
    );
nor_n_161: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S459,
        in1(1) => S416,
        out1 => S461
    );
notg_86: ENTITY WORK.notg
    PORT MAP (
        in1 => S461,
        out1 => S462
    );
nor_n_162: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S461,
        in1(1) => CU_ADD,
        out1 => S463
    );
nand_n_224: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S463,
        in1(1) => S460,
        out1 => S464
    );
nand_n_225: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S464,
        in1(1) => S430,
        out1 => S330
    );
nor_n_163: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_4,
        in1(1) => DP_AC_out_4,
        out1 => S465
    );
nor_n_164: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1075,
        in1(1) => S1064,
        out1 => S466
    );
nand_n_226: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_4,
        in1(1) => DP_AC_out_4,
        out1 => S467
    );
nor_n_165: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S466,
        in1(1) => S465,
        out1 => S468
    );
nor_n_166: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S423,
        in1(1) => S421,
        out1 => S469
    );
nor_n_167: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S469,
        in1(1) => S422,
        out1 => S470
    );
nand_n_227: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S470,
        in1(1) => S468,
        out1 => S471
    );
notg_87: ENTITY WORK.notg
    PORT MAP (
        in1 => S471,
        out1 => S472
    );
nor_n_168: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S470,
        in1(1) => S468,
        out1 => S473
    );
nor_n_169: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S473,
        in1(1) => S472,
        out1 => S474
    );
nor_n_170: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S474,
        in1(1) => S988,
        out1 => S475
    );
nor_n_171: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S457,
        in1(1) => S452,
        out1 => S476
    );
nand_n_228: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S458,
        in1(1) => S451,
        out1 => S477
    );
nand_n_229: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_4,
        in1(1) => DP_AC_out_0,
        out1 => S478
    );
nand_n_230: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_3,
        in1(1) => DP_AC_out_1,
        out1 => S479
    );
nand_n_231: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S479,
        in1(1) => S478,
        out1 => S480
    );
notg_88: ENTITY WORK.notg
    PORT MAP (
        in1 => S480,
        out1 => S481
    );
nand_n_232: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_4,
        in1(1) => DP_AC_out_1,
        out1 => S482
    );
notg_89: ENTITY WORK.notg
    PORT MAP (
        in1 => S482,
        out1 => S483
    );
nor_n_172: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S482,
        in1(1) => S431,
        out1 => S484
    );
nand_n_233: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S483,
        in1(1) => S432,
        out1 => S485
    );
nor_n_173: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S484,
        in1(1) => S481,
        out1 => S486
    );
notg_90: ENTITY WORK.notg
    PORT MAP (
        in1 => S486,
        out1 => S487
    );
nor_n_174: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S447,
        in1(1) => S440,
        out1 => S488
    );
nand_n_234: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S448,
        in1(1) => S441,
        out1 => S489
    );
nand_n_235: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_4,
        in1(1) => DP_ARU1_in1_0,
        out1 => S490
    );
nand_n_236: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_4,
        in1(1) => DP_ARU1_in1_1,
        out1 => S491
    );
notg_91: ENTITY WORK.notg
    PORT MAP (
        in1 => S491,
        out1 => S492
    );
nor_n_175: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S490,
        in1(1) => S439,
        out1 => S493
    );
nand_n_237: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S492,
        in1(1) => S438,
        out1 => S494
    );
nand_n_238: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S490,
        in1(1) => S439,
        out1 => S495
    );
notg_92: ENTITY WORK.notg
    PORT MAP (
        in1 => S495,
        out1 => S496
    );
nor_n_176: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S496,
        in1(1) => S493,
        out1 => S497
    );
nand_n_239: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S495,
        in1(1) => S494,
        out1 => S498
    );
nor_n_177: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S497,
        in1(1) => S397,
        out1 => S499
    );
nand_n_240: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S498,
        in1(1) => S398,
        out1 => S500
    );
nor_n_178: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S498,
        in1(1) => S398,
        out1 => S501
    );
nand_n_241: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S497,
        in1(1) => S397,
        out1 => S502
    );
nor_n_179: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S501,
        in1(1) => S499,
        out1 => S503
    );
nand_n_242: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S502,
        in1(1) => S500,
        out1 => S504
    );
nor_n_180: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S504,
        in1(1) => S488,
        out1 => S505
    );
nand_n_243: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S503,
        in1(1) => S489,
        out1 => S506
    );
nor_n_181: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S503,
        in1(1) => S489,
        out1 => S507
    );
nand_n_244: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S504,
        in1(1) => S488,
        out1 => S508
    );
nor_n_182: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S507,
        in1(1) => S505,
        out1 => S509
    );
nand_n_245: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S508,
        in1(1) => S506,
        out1 => S510
    );
nor_n_183: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S509,
        in1(1) => S486,
        out1 => S511
    );
nor_n_184: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S510,
        in1(1) => S487,
        out1 => S512
    );
nand_n_246: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S509,
        in1(1) => S486,
        out1 => S513
    );
nor_n_185: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S512,
        in1(1) => S511,
        out1 => S514
    );
notg_93: ENTITY WORK.notg
    PORT MAP (
        in1 => S514,
        out1 => S515
    );
nor_n_186: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S515,
        in1(1) => S476,
        out1 => S516
    );
notg_94: ENTITY WORK.notg
    PORT MAP (
        in1 => S516,
        out1 => S517
    );
nor_n_187: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S514,
        in1(1) => S477,
        out1 => S518
    );
nor_n_188: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S518,
        in1(1) => S516,
        out1 => S519
    );
notg_95: ENTITY WORK.notg
    PORT MAP (
        in1 => S519,
        out1 => S520
    );
nor_n_189: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S519,
        in1(1) => S461,
        out1 => S521
    );
nor_n_190: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S520,
        in1(1) => S462,
        out1 => S522
    );
notg_96: ENTITY WORK.notg
    PORT MAP (
        in1 => S522,
        out1 => S523
    );
nor_n_191: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S522,
        in1(1) => S521,
        out1 => S524
    );
nor_n_192: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S524,
        in1(1) => CU_ADD,
        out1 => S525
    );
nor_n_193: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S525,
        in1(1) => S475,
        out1 => S331
    );
nand_n_247: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S471,
        in1(1) => S467,
        out1 => S526
    );
nor_n_194: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_5,
        in1(1) => DP_AC_out_5,
        out1 => S527
    );
nor_n_195: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1096,
        in1(1) => S1085,
        out1 => S528
    );
nand_n_248: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_5,
        in1(1) => DP_AC_out_5,
        out1 => S529
    );
nor_n_196: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S528,
        in1(1) => S527,
        out1 => S530
    );
nor_n_197: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S530,
        in1(1) => S526,
        out1 => S531
    );
nand_n_249: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S530,
        in1(1) => S526,
        out1 => S532
    );
notg_97: ENTITY WORK.notg
    PORT MAP (
        in1 => S532,
        out1 => S533
    );
nor_n_198: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S533,
        in1(1) => S531,
        out1 => S534
    );
nor_n_199: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S534,
        in1(1) => S988,
        out1 => S535
    );
nor_n_200: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S512,
        in1(1) => S505,
        out1 => S536
    );
nand_n_250: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S513,
        in1(1) => S506,
        out1 => S537
    );
nand_n_251: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_5,
        in1(1) => DP_AC_out_0,
        out1 => S538
    );
nand_n_252: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_3,
        in1(1) => DP_AC_out_2,
        out1 => S539
    );
nand_n_253: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_4,
        in1(1) => DP_AC_out_2,
        out1 => S540
    );
nor_n_201: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S539,
        in1(1) => S482,
        out1 => S541
    );
notg_98: ENTITY WORK.notg
    PORT MAP (
        in1 => S541,
        out1 => S542
    );
nand_n_254: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S539,
        in1(1) => S482,
        out1 => S543
    );
nand_n_255: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S543,
        in1(1) => S542,
        out1 => S544
    );
nand_n_256: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S544,
        in1(1) => S538,
        out1 => S545
    );
notg_99: ENTITY WORK.notg
    PORT MAP (
        in1 => S545,
        out1 => S546
    );
nor_n_202: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S544,
        in1(1) => S538,
        out1 => S547
    );
notg_100: ENTITY WORK.notg
    PORT MAP (
        in1 => S547,
        out1 => S548
    );
nor_n_203: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S547,
        in1(1) => S546,
        out1 => S549
    );
nand_n_257: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S548,
        in1(1) => S545,
        out1 => S550
    );
nor_n_204: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S501,
        in1(1) => S493,
        out1 => S551
    );
nand_n_258: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S502,
        in1(1) => S494,
        out1 => S552
    );
nand_n_259: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_3,
        in1(1) => DP_ARU1_in1_2,
        out1 => S553
    );
notg_101: ENTITY WORK.notg
    PORT MAP (
        in1 => S553,
        out1 => S554
    );
nand_n_260: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_5,
        in1(1) => DP_ARU1_in1_0,
        out1 => S555
    );
notg_102: ENTITY WORK.notg
    PORT MAP (
        in1 => S555,
        out1 => S556
    );
nand_n_261: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_5,
        in1(1) => DP_ARU1_in1_1,
        out1 => S557
    );
nor_n_205: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S555,
        in1(1) => S491,
        out1 => S558
    );
nand_n_262: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S556,
        in1(1) => S492,
        out1 => S559
    );
nand_n_263: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S555,
        in1(1) => S491,
        out1 => S560
    );
notg_103: ENTITY WORK.notg
    PORT MAP (
        in1 => S560,
        out1 => S561
    );
nor_n_206: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S561,
        in1(1) => S558,
        out1 => S562
    );
nand_n_264: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S560,
        in1(1) => S559,
        out1 => S563
    );
nor_n_207: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S562,
        in1(1) => S554,
        out1 => S564
    );
nand_n_265: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S563,
        in1(1) => S553,
        out1 => S565
    );
nor_n_208: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S563,
        in1(1) => S553,
        out1 => S566
    );
nand_n_266: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S562,
        in1(1) => S554,
        out1 => S567
    );
nor_n_209: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S566,
        in1(1) => S564,
        out1 => S568
    );
nand_n_267: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S567,
        in1(1) => S565,
        out1 => S569
    );
nor_n_210: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S569,
        in1(1) => S551,
        out1 => S570
    );
nand_n_268: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S568,
        in1(1) => S552,
        out1 => S571
    );
nor_n_211: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S568,
        in1(1) => S552,
        out1 => S572
    );
nand_n_269: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S569,
        in1(1) => S551,
        out1 => S573
    );
nor_n_212: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S572,
        in1(1) => S570,
        out1 => S574
    );
nand_n_270: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S573,
        in1(1) => S571,
        out1 => S575
    );
nor_n_213: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S574,
        in1(1) => S549,
        out1 => S576
    );
nand_n_271: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S575,
        in1(1) => S550,
        out1 => S577
    );
nor_n_214: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S575,
        in1(1) => S550,
        out1 => S578
    );
nand_n_272: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S574,
        in1(1) => S549,
        out1 => S579
    );
nor_n_215: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S578,
        in1(1) => S576,
        out1 => S580
    );
nand_n_273: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S579,
        in1(1) => S577,
        out1 => S581
    );
nor_n_216: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S581,
        in1(1) => S536,
        out1 => S582
    );
nand_n_274: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S580,
        in1(1) => S537,
        out1 => S583
    );
nor_n_217: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S580,
        in1(1) => S537,
        out1 => S584
    );
nand_n_275: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S581,
        in1(1) => S536,
        out1 => S585
    );
nor_n_218: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S584,
        in1(1) => S582,
        out1 => S586
    );
nand_n_276: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S585,
        in1(1) => S583,
        out1 => S587
    );
nor_n_219: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S587,
        in1(1) => S485,
        out1 => S588
    );
nand_n_277: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S586,
        in1(1) => S484,
        out1 => S589
    );
nor_n_220: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S586,
        in1(1) => S484,
        out1 => S590
    );
nand_n_278: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S587,
        in1(1) => S485,
        out1 => S591
    );
nor_n_221: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S590,
        in1(1) => S588,
        out1 => S592
    );
nand_n_279: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S591,
        in1(1) => S589,
        out1 => S593
    );
nor_n_222: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S593,
        in1(1) => S517,
        out1 => S594
    );
nand_n_280: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S592,
        in1(1) => S516,
        out1 => S595
    );
nor_n_223: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S592,
        in1(1) => S516,
        out1 => S596
    );
nor_n_224: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S596,
        in1(1) => S594,
        out1 => S597
    );
notg_104: ENTITY WORK.notg
    PORT MAP (
        in1 => S597,
        out1 => S598
    );
nor_n_225: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S597,
        in1(1) => S522,
        out1 => S599
    );
nor_n_226: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S598,
        in1(1) => S523,
        out1 => S600
    );
nand_n_281: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S597,
        in1(1) => S522,
        out1 => S601
    );
nor_n_227: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S600,
        in1(1) => S599,
        out1 => S602
    );
nor_n_228: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S602,
        in1(1) => CU_ADD,
        out1 => S603
    );
nor_n_229: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S603,
        in1(1) => S535,
        out1 => S332
    );
nand_n_282: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S532,
        in1(1) => S529,
        out1 => S604
    );
nor_n_230: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_6,
        in1(1) => DP_AC_out_6,
        out1 => S605
    );
nor_n_231: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1118,
        in1(1) => S1107,
        out1 => S606
    );
nand_n_283: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_6,
        in1(1) => DP_AC_out_6,
        out1 => S607
    );
nor_n_232: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S606,
        in1(1) => S605,
        out1 => S608
    );
nor_n_233: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S608,
        in1(1) => S604,
        out1 => S609
    );
nand_n_284: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S608,
        in1(1) => S604,
        out1 => S610
    );
nor_n_234: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S588,
        in1(1) => S582,
        out1 => S611
    );
nand_n_285: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S589,
        in1(1) => S583,
        out1 => S612
    );
nand_n_286: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_6,
        in1(1) => DP_AC_out_0,
        out1 => S613
    );
notg_105: ENTITY WORK.notg
    PORT MAP (
        in1 => S613,
        out1 => S614
    );
nor_n_235: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S547,
        in1(1) => S541,
        out1 => S615
    );
notg_106: ENTITY WORK.notg
    PORT MAP (
        in1 => S615,
        out1 => S616
    );
nor_n_236: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S615,
        in1(1) => S613,
        out1 => S617
    );
nand_n_287: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S616,
        in1(1) => S614,
        out1 => S618
    );
nand_n_288: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S615,
        in1(1) => S613,
        out1 => S619
    );
notg_107: ENTITY WORK.notg
    PORT MAP (
        in1 => S619,
        out1 => S620
    );
nor_n_237: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S620,
        in1(1) => S617,
        out1 => S621
    );
nand_n_289: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S619,
        in1(1) => S618,
        out1 => S622
    );
nor_n_238: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S578,
        in1(1) => S570,
        out1 => S623
    );
nand_n_290: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S579,
        in1(1) => S571,
        out1 => S624
    );
nand_n_291: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_5,
        in1(1) => DP_AC_out_1,
        out1 => S625
    );
nand_n_292: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_4,
        in1(1) => DP_AC_out_3,
        out1 => S626
    );
nor_n_239: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S540,
        in1(1) => S424,
        out1 => S627
    );
notg_108: ENTITY WORK.notg
    PORT MAP (
        in1 => S627,
        out1 => S628
    );
nand_n_293: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S540,
        in1(1) => S424,
        out1 => S629
    );
nand_n_294: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S629,
        in1(1) => S628,
        out1 => S630
    );
nand_n_295: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S630,
        in1(1) => S625,
        out1 => S631
    );
notg_109: ENTITY WORK.notg
    PORT MAP (
        in1 => S631,
        out1 => S632
    );
nor_n_240: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S630,
        in1(1) => S625,
        out1 => S633
    );
notg_110: ENTITY WORK.notg
    PORT MAP (
        in1 => S633,
        out1 => S634
    );
nor_n_241: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S633,
        in1(1) => S632,
        out1 => S635
    );
nand_n_296: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S634,
        in1(1) => S631,
        out1 => S636
    );
nor_n_242: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S566,
        in1(1) => S558,
        out1 => S637
    );
nand_n_297: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S567,
        in1(1) => S559,
        out1 => S638
    );
nand_n_298: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_4,
        in1(1) => DP_ARU1_in1_2,
        out1 => S639
    );
notg_111: ENTITY WORK.notg
    PORT MAP (
        in1 => S639,
        out1 => S640
    );
nand_n_299: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_6,
        in1(1) => DP_ARU1_in1_0,
        out1 => S641
    );
nor_n_243: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1107,
        in1(1) => S1009,
        out1 => S642
    );
nand_n_300: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_6,
        in1(1) => DP_ARU1_in1_1,
        out1 => S643
    );
nor_n_244: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S643,
        in1(1) => S555,
        out1 => S644
    );
nand_n_301: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S642,
        in1(1) => S556,
        out1 => S645
    );
nand_n_302: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S641,
        in1(1) => S557,
        out1 => S646
    );
notg_112: ENTITY WORK.notg
    PORT MAP (
        in1 => S646,
        out1 => S647
    );
nor_n_245: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S647,
        in1(1) => S644,
        out1 => S648
    );
nand_n_303: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S646,
        in1(1) => S645,
        out1 => S649
    );
nor_n_246: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S648,
        in1(1) => S640,
        out1 => S650
    );
nand_n_304: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S649,
        in1(1) => S639,
        out1 => S651
    );
nor_n_247: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S649,
        in1(1) => S639,
        out1 => S652
    );
nand_n_305: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S648,
        in1(1) => S640,
        out1 => S653
    );
nor_n_248: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S652,
        in1(1) => S650,
        out1 => S654
    );
nand_n_306: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S653,
        in1(1) => S651,
        out1 => S655
    );
nor_n_249: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S655,
        in1(1) => S637,
        out1 => S656
    );
nand_n_307: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S654,
        in1(1) => S638,
        out1 => S657
    );
nor_n_250: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S654,
        in1(1) => S638,
        out1 => S658
    );
nand_n_308: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S655,
        in1(1) => S637,
        out1 => S659
    );
nor_n_251: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S658,
        in1(1) => S656,
        out1 => S660
    );
nand_n_309: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S659,
        in1(1) => S657,
        out1 => S661
    );
nor_n_252: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S660,
        in1(1) => S635,
        out1 => S662
    );
nand_n_310: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S661,
        in1(1) => S636,
        out1 => S663
    );
nor_n_253: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S661,
        in1(1) => S636,
        out1 => S664
    );
nand_n_311: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S660,
        in1(1) => S635,
        out1 => S665
    );
nor_n_254: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S664,
        in1(1) => S662,
        out1 => S666
    );
nand_n_312: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S665,
        in1(1) => S663,
        out1 => S667
    );
nor_n_255: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S667,
        in1(1) => S623,
        out1 => S668
    );
nand_n_313: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S666,
        in1(1) => S624,
        out1 => S669
    );
nor_n_256: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S666,
        in1(1) => S624,
        out1 => S670
    );
nand_n_314: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S667,
        in1(1) => S623,
        out1 => S671
    );
nor_n_257: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S670,
        in1(1) => S668,
        out1 => S672
    );
nand_n_315: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S671,
        in1(1) => S669,
        out1 => S673
    );
nor_n_258: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S673,
        in1(1) => S622,
        out1 => S674
    );
nand_n_316: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S672,
        in1(1) => S621,
        out1 => S675
    );
nor_n_259: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S672,
        in1(1) => S621,
        out1 => S676
    );
nand_n_317: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S673,
        in1(1) => S622,
        out1 => S677
    );
nor_n_260: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S676,
        in1(1) => S674,
        out1 => S678
    );
nand_n_318: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S677,
        in1(1) => S675,
        out1 => S679
    );
nor_n_261: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S678,
        in1(1) => S612,
        out1 => S680
    );
nand_n_319: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S679,
        in1(1) => S611,
        out1 => S681
    );
nor_n_262: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S679,
        in1(1) => S611,
        out1 => S682
    );
nand_n_320: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S678,
        in1(1) => S612,
        out1 => S683
    );
nor_n_263: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S682,
        in1(1) => S680,
        out1 => S684
    );
nand_n_321: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S683,
        in1(1) => S681,
        out1 => S685
    );
nor_n_264: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S685,
        in1(1) => S595,
        out1 => S686
    );
nand_n_322: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S684,
        in1(1) => S594,
        out1 => S687
    );
nor_n_265: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S684,
        in1(1) => S594,
        out1 => S688
    );
nand_n_323: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S685,
        in1(1) => S595,
        out1 => S689
    );
nor_n_266: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S688,
        in1(1) => S686,
        out1 => S690
    );
nand_n_324: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S689,
        in1(1) => S687,
        out1 => S691
    );
nor_n_267: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S690,
        in1(1) => S600,
        out1 => S692
    );
nor_n_268: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S691,
        in1(1) => S601,
        out1 => S693
    );
nand_n_325: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S690,
        in1(1) => S600,
        out1 => S694
    );
nor_n_269: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S693,
        in1(1) => S692,
        out1 => S695
    );
nor_n_270: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S609,
        in1(1) => S988,
        out1 => S696
    );
nand_n_326: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S696,
        in1(1) => S610,
        out1 => S697
    );
nand_n_327: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S695,
        in1(1) => S988,
        out1 => S698
    );
nand_n_328: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S698,
        in1(1) => S697,
        out1 => S333
    );
nand_n_329: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S610,
        in1(1) => S607,
        out1 => S699
    );
nor_n_271: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_7,
        in1(1) => DP_AC_out_7,
        out1 => S700
    );
nor_n_272: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1140,
        in1(1) => S1129,
        out1 => S701
    );
nand_n_330: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_7,
        in1(1) => DP_AC_out_7,
        out1 => S702
    );
nor_n_273: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S701,
        in1(1) => S700,
        out1 => S703
    );
nand_n_331: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S703,
        in1(1) => S699,
        out1 => S704
    );
notg_113: ENTITY WORK.notg
    PORT MAP (
        in1 => S704,
        out1 => S705
    );
nor_n_274: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S703,
        in1(1) => S699,
        out1 => S706
    );
nor_n_275: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S706,
        in1(1) => S705,
        out1 => S707
    );
nor_n_276: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S693,
        in1(1) => S686,
        out1 => S708
    );
nand_n_332: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S694,
        in1(1) => S687,
        out1 => S709
    );
nor_n_277: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S674,
        in1(1) => S668,
        out1 => S710
    );
nand_n_333: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S675,
        in1(1) => S669,
        out1 => S711
    );
nand_n_334: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_7,
        in1(1) => DP_AC_out_0,
        out1 => S712
    );
nand_n_335: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_6,
        in1(1) => DP_AC_out_1,
        out1 => S713
    );
nor_n_278: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S633,
        in1(1) => S627,
        out1 => S714
    );
nor_n_279: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S714,
        in1(1) => S713,
        out1 => S715
    );
notg_114: ENTITY WORK.notg
    PORT MAP (
        in1 => S715,
        out1 => S716
    );
nand_n_336: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S714,
        in1(1) => S713,
        out1 => S717
    );
nand_n_337: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S717,
        in1(1) => S716,
        out1 => S718
    );
nand_n_338: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S718,
        in1(1) => S712,
        out1 => S719
    );
notg_115: ENTITY WORK.notg
    PORT MAP (
        in1 => S719,
        out1 => S720
    );
nor_n_280: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S718,
        in1(1) => S712,
        out1 => S721
    );
notg_116: ENTITY WORK.notg
    PORT MAP (
        in1 => S721,
        out1 => S722
    );
nor_n_281: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S721,
        in1(1) => S720,
        out1 => S723
    );
nand_n_339: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S722,
        in1(1) => S719,
        out1 => S724
    );
nor_n_282: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S664,
        in1(1) => S656,
        out1 => S725
    );
nand_n_340: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S665,
        in1(1) => S657,
        out1 => S726
    );
nand_n_341: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_5,
        in1(1) => DP_AC_out_2,
        out1 => S727
    );
nand_n_342: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_4,
        in1(1) => DP_ARU1_in1_3,
        out1 => S728
    );
nor_n_283: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S467,
        in1(1) => S424,
        out1 => S729
    );
notg_117: ENTITY WORK.notg
    PORT MAP (
        in1 => S729,
        out1 => S730
    );
nand_n_343: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S728,
        in1(1) => S626,
        out1 => S731
    );
nand_n_344: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S731,
        in1(1) => S730,
        out1 => S732
    );
nand_n_345: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S732,
        in1(1) => S727,
        out1 => S733
    );
notg_118: ENTITY WORK.notg
    PORT MAP (
        in1 => S733,
        out1 => S734
    );
nor_n_284: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S732,
        in1(1) => S727,
        out1 => S735
    );
notg_119: ENTITY WORK.notg
    PORT MAP (
        in1 => S735,
        out1 => S736
    );
nor_n_285: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S735,
        in1(1) => S734,
        out1 => S737
    );
nand_n_346: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S736,
        in1(1) => S733,
        out1 => S738
    );
nor_n_286: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S652,
        in1(1) => S644,
        out1 => S739
    );
nand_n_347: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S653,
        in1(1) => S645,
        out1 => S740
    );
nand_n_348: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_5,
        in1(1) => DP_ARU1_in1_2,
        out1 => S741
    );
notg_120: ENTITY WORK.notg
    PORT MAP (
        in1 => S741,
        out1 => S742
    );
nand_n_349: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_7,
        in1(1) => DP_ARU1_in1_0,
        out1 => S743
    );
nand_n_350: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_7,
        in1(1) => DP_ARU1_in1_1,
        out1 => S744
    );
nor_n_287: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S744,
        in1(1) => S641,
        out1 => S745
    );
notg_121: ENTITY WORK.notg
    PORT MAP (
        in1 => S745,
        out1 => S746
    );
nand_n_351: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S743,
        in1(1) => S643,
        out1 => S747
    );
notg_122: ENTITY WORK.notg
    PORT MAP (
        in1 => S747,
        out1 => S748
    );
nor_n_288: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S748,
        in1(1) => S745,
        out1 => S749
    );
nand_n_352: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S747,
        in1(1) => S746,
        out1 => S750
    );
nor_n_289: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S749,
        in1(1) => S742,
        out1 => S751
    );
nand_n_353: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S750,
        in1(1) => S741,
        out1 => S752
    );
nor_n_290: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S750,
        in1(1) => S741,
        out1 => S753
    );
nand_n_354: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S749,
        in1(1) => S742,
        out1 => S754
    );
nor_n_291: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S753,
        in1(1) => S751,
        out1 => S755
    );
nand_n_355: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S754,
        in1(1) => S752,
        out1 => S756
    );
nor_n_292: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S756,
        in1(1) => S739,
        out1 => S757
    );
nand_n_356: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S755,
        in1(1) => S740,
        out1 => S758
    );
nor_n_293: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S755,
        in1(1) => S740,
        out1 => S759
    );
nand_n_357: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S756,
        in1(1) => S739,
        out1 => S760
    );
nor_n_294: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S759,
        in1(1) => S757,
        out1 => S761
    );
nand_n_358: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S760,
        in1(1) => S758,
        out1 => S762
    );
nor_n_295: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S761,
        in1(1) => S737,
        out1 => S763
    );
nand_n_359: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S762,
        in1(1) => S738,
        out1 => S764
    );
nor_n_296: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S762,
        in1(1) => S738,
        out1 => S765
    );
nand_n_360: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S761,
        in1(1) => S737,
        out1 => S766
    );
nor_n_297: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S765,
        in1(1) => S763,
        out1 => S767
    );
nand_n_361: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S766,
        in1(1) => S764,
        out1 => S768
    );
nor_n_298: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S768,
        in1(1) => S725,
        out1 => S769
    );
nand_n_362: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S767,
        in1(1) => S726,
        out1 => S770
    );
nor_n_299: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S767,
        in1(1) => S726,
        out1 => S771
    );
nand_n_363: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S768,
        in1(1) => S725,
        out1 => S772
    );
nor_n_300: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S771,
        in1(1) => S769,
        out1 => S773
    );
nand_n_364: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S772,
        in1(1) => S770,
        out1 => S774
    );
nor_n_301: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S773,
        in1(1) => S723,
        out1 => S775
    );
nand_n_365: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S774,
        in1(1) => S724,
        out1 => S776
    );
nor_n_302: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S774,
        in1(1) => S724,
        out1 => S777
    );
nand_n_366: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S773,
        in1(1) => S723,
        out1 => S778
    );
nor_n_303: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S777,
        in1(1) => S775,
        out1 => S779
    );
nand_n_367: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S778,
        in1(1) => S776,
        out1 => S780
    );
nor_n_304: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S780,
        in1(1) => S710,
        out1 => S781
    );
nand_n_368: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S779,
        in1(1) => S711,
        out1 => S782
    );
nor_n_305: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S779,
        in1(1) => S711,
        out1 => S783
    );
nand_n_369: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S780,
        in1(1) => S710,
        out1 => S784
    );
nor_n_306: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S783,
        in1(1) => S781,
        out1 => S785
    );
nand_n_370: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S784,
        in1(1) => S782,
        out1 => S786
    );
nor_n_307: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S785,
        in1(1) => S617,
        out1 => S787
    );
nand_n_371: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S786,
        in1(1) => S618,
        out1 => S788
    );
nor_n_308: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S786,
        in1(1) => S618,
        out1 => S789
    );
nand_n_372: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S785,
        in1(1) => S617,
        out1 => S790
    );
nor_n_309: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S789,
        in1(1) => S787,
        out1 => S791
    );
nand_n_373: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S790,
        in1(1) => S788,
        out1 => S792
    );
nor_n_310: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S792,
        in1(1) => S683,
        out1 => S793
    );
nand_n_374: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S791,
        in1(1) => S682,
        out1 => S794
    );
nor_n_311: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S791,
        in1(1) => S682,
        out1 => S795
    );
nand_n_375: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S792,
        in1(1) => S683,
        out1 => S796
    );
nor_n_312: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S795,
        in1(1) => S793,
        out1 => S797
    );
nand_n_376: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S796,
        in1(1) => S794,
        out1 => S798
    );
nor_n_313: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S798,
        in1(1) => S708,
        out1 => S799
    );
nand_n_377: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S797,
        in1(1) => S709,
        out1 => S800
    );
nor_n_314: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S797,
        in1(1) => S709,
        out1 => S801
    );
nor_n_315: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S801,
        in1(1) => S799,
        out1 => S802
    );
nor_n_316: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S802,
        in1(1) => CU_ADD,
        out1 => S803
    );
nor_n_317: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S707,
        in1(1) => S988,
        out1 => S804
    );
nor_n_318: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S804,
        in1(1) => S803,
        out1 => S334
    );
nor_n_319: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_8,
        in1(1) => DP_AC_out_8,
        out1 => S805
    );
nand_n_378: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_8,
        in1(1) => DP_AC_out_8,
        out1 => S806
    );
notg_123: ENTITY WORK.notg
    PORT MAP (
        in1 => S806,
        out1 => S807
    );
nor_n_320: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S807,
        in1(1) => S805,
        out1 => S808
    );
nor_n_321: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S701,
        in1(1) => S699,
        out1 => S809
    );
nor_n_322: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S809,
        in1(1) => S700,
        out1 => S810
    );
nand_n_379: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S810,
        in1(1) => S808,
        out1 => S811
    );
nor_n_323: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S810,
        in1(1) => S808,
        out1 => S812
    );
nor_n_324: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S799,
        in1(1) => S793,
        out1 => S813
    );
nand_n_380: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S800,
        in1(1) => S794,
        out1 => S814
    );
nor_n_325: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S789,
        in1(1) => S781,
        out1 => S815
    );
nand_n_381: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S790,
        in1(1) => S782,
        out1 => S816
    );
nor_n_326: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S721,
        in1(1) => S715,
        out1 => S817
    );
nor_n_327: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S777,
        in1(1) => S769,
        out1 => S818
    );
notg_124: ENTITY WORK.notg
    PORT MAP (
        in1 => S818,
        out1 => S819
    );
nand_n_382: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_7,
        in1(1) => DP_AC_out_1,
        out1 => S820
    );
nand_n_383: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_6,
        in1(1) => DP_AC_out_2,
        out1 => S821
    );
nor_n_328: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S735,
        in1(1) => S729,
        out1 => S822
    );
nor_n_329: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S822,
        in1(1) => S821,
        out1 => S823
    );
notg_125: ENTITY WORK.notg
    PORT MAP (
        in1 => S823,
        out1 => S824
    );
nand_n_384: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S822,
        in1(1) => S821,
        out1 => S825
    );
nand_n_385: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S825,
        in1(1) => S824,
        out1 => S826
    );
nor_n_330: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S826,
        in1(1) => S820,
        out1 => S827
    );
notg_126: ENTITY WORK.notg
    PORT MAP (
        in1 => S827,
        out1 => S828
    );
nand_n_386: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S826,
        in1(1) => S820,
        out1 => S829
    );
notg_127: ENTITY WORK.notg
    PORT MAP (
        in1 => S829,
        out1 => S830
    );
nor_n_331: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S830,
        in1(1) => S827,
        out1 => S831
    );
nand_n_387: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S829,
        in1(1) => S828,
        out1 => S832
    );
nor_n_332: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S765,
        in1(1) => S757,
        out1 => S833
    );
nand_n_388: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S766,
        in1(1) => S758,
        out1 => S834
    );
nand_n_389: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_5,
        in1(1) => DP_AC_out_3,
        out1 => S835
    );
nand_n_390: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_5,
        in1(1) => DP_ARU1_in1_3,
        out1 => S836
    );
nand_n_391: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_5,
        in1(1) => DP_ARU1_in1_4,
        out1 => S837
    );
nor_n_333: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S836,
        in1(1) => S467,
        out1 => S838
    );
notg_128: ENTITY WORK.notg
    PORT MAP (
        in1 => S838,
        out1 => S839
    );
nand_n_392: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S836,
        in1(1) => S467,
        out1 => S840
    );
nand_n_393: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S840,
        in1(1) => S839,
        out1 => S841
    );
nand_n_394: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S841,
        in1(1) => S835,
        out1 => S842
    );
notg_129: ENTITY WORK.notg
    PORT MAP (
        in1 => S842,
        out1 => S843
    );
nor_n_334: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S841,
        in1(1) => S835,
        out1 => S844
    );
notg_130: ENTITY WORK.notg
    PORT MAP (
        in1 => S844,
        out1 => S845
    );
nor_n_335: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S844,
        in1(1) => S843,
        out1 => S846
    );
nand_n_395: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S845,
        in1(1) => S842,
        out1 => S847
    );
nor_n_336: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S753,
        in1(1) => S745,
        out1 => S848
    );
notg_131: ENTITY WORK.notg
    PORT MAP (
        in1 => S848,
        out1 => S849
    );
nand_n_396: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_6,
        in1(1) => DP_ARU1_in1_2,
        out1 => S850
    );
nor_n_337: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1129,
        in1(1) => S1031,
        out1 => S851
    );
nand_n_397: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_7,
        in1(1) => DP_ARU1_in1_2,
        out1 => S852
    );
nor_n_338: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S852,
        in1(1) => S643,
        out1 => S853
    );
nand_n_398: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S851,
        in1(1) => S642,
        out1 => S854
    );
nand_n_399: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S850,
        in1(1) => S744,
        out1 => S855
    );
nand_n_400: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S855,
        in1(1) => S854,
        out1 => S856
    );
notg_132: ENTITY WORK.notg
    PORT MAP (
        in1 => S856,
        out1 => S857
    );
nor_n_339: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S856,
        in1(1) => S848,
        out1 => S858
    );
nand_n_401: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S857,
        in1(1) => S849,
        out1 => S859
    );
nand_n_402: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S856,
        in1(1) => S848,
        out1 => S860
    );
notg_133: ENTITY WORK.notg
    PORT MAP (
        in1 => S860,
        out1 => S861
    );
nor_n_340: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S861,
        in1(1) => S858,
        out1 => S862
    );
nand_n_403: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S860,
        in1(1) => S859,
        out1 => S863
    );
nor_n_341: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S862,
        in1(1) => S846,
        out1 => S864
    );
nand_n_404: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S863,
        in1(1) => S847,
        out1 => S865
    );
nor_n_342: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S863,
        in1(1) => S847,
        out1 => S866
    );
nand_n_405: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S862,
        in1(1) => S846,
        out1 => S867
    );
nor_n_343: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S866,
        in1(1) => S864,
        out1 => S868
    );
nand_n_406: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S867,
        in1(1) => S865,
        out1 => S869
    );
nor_n_344: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S869,
        in1(1) => S833,
        out1 => S870
    );
nand_n_407: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S868,
        in1(1) => S834,
        out1 => S871
    );
nor_n_345: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S868,
        in1(1) => S834,
        out1 => S872
    );
nand_n_408: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S869,
        in1(1) => S833,
        out1 => S873
    );
nor_n_346: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S872,
        in1(1) => S870,
        out1 => S874
    );
nand_n_409: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S873,
        in1(1) => S871,
        out1 => S875
    );
nor_n_347: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S874,
        in1(1) => S831,
        out1 => S876
    );
nand_n_410: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S875,
        in1(1) => S832,
        out1 => S877
    );
nor_n_348: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S875,
        in1(1) => S832,
        out1 => S878
    );
nand_n_411: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S874,
        in1(1) => S831,
        out1 => S879
    );
nor_n_349: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S878,
        in1(1) => S876,
        out1 => S880
    );
nand_n_412: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S879,
        in1(1) => S877,
        out1 => S881
    );
nor_n_350: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S881,
        in1(1) => S818,
        out1 => S882
    );
nand_n_413: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S880,
        in1(1) => S819,
        out1 => S883
    );
nand_n_414: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S881,
        in1(1) => S818,
        out1 => S884
    );
nand_n_415: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S884,
        in1(1) => S883,
        out1 => S885
    );
nand_n_416: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S885,
        in1(1) => S817,
        out1 => S886
    );
notg_134: ENTITY WORK.notg
    PORT MAP (
        in1 => S886,
        out1 => S887
    );
nor_n_351: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S885,
        in1(1) => S817,
        out1 => S888
    );
notg_135: ENTITY WORK.notg
    PORT MAP (
        in1 => S888,
        out1 => S889
    );
nor_n_352: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S888,
        in1(1) => S887,
        out1 => S890
    );
nand_n_417: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S889,
        in1(1) => S886,
        out1 => S891
    );
nor_n_353: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S891,
        in1(1) => S815,
        out1 => S892
    );
nand_n_418: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S890,
        in1(1) => S816,
        out1 => S893
    );
nor_n_354: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S890,
        in1(1) => S816,
        out1 => S894
    );
nand_n_419: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S891,
        in1(1) => S815,
        out1 => S895
    );
nor_n_355: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S894,
        in1(1) => S892,
        out1 => S896
    );
nand_n_420: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S895,
        in1(1) => S893,
        out1 => S897
    );
nand_n_421: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S897,
        in1(1) => S813,
        out1 => S898
    );
nor_n_356: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S897,
        in1(1) => S813,
        out1 => S899
    );
nand_n_422: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S896,
        in1(1) => S814,
        out1 => S900
    );
nand_n_423: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S900,
        in1(1) => S898,
        out1 => S901
    );
nor_n_357: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S901,
        in1(1) => CU_ADD,
        out1 => S902
    );
nand_n_424: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S811,
        in1(1) => CU_ADD,
        out1 => S903
    );
nor_n_358: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S903,
        in1(1) => S812,
        out1 => S904
    );
nor_n_359: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S904,
        in1(1) => S902,
        out1 => S905
    );
notg_136: ENTITY WORK.notg
    PORT MAP (
        in1 => S905,
        out1 => S335
    );
nand_n_425: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S811,
        in1(1) => S806,
        out1 => S906
    );
nand_n_426: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1161,
        in1(1) => S1150,
        out1 => S907
    );
nand_n_427: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_9,
        in1(1) => DP_AC_out_9,
        out1 => S908
    );
nand_n_428: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S908,
        in1(1) => S907,
        out1 => S909
    );
nand_n_429: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S909,
        in1(1) => S906,
        out1 => S910
    );
nor_n_360: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S909,
        in1(1) => S906,
        out1 => S911
    );
notg_137: ENTITY WORK.notg
    PORT MAP (
        in1 => S911,
        out1 => S912
    );
nand_n_430: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S912,
        in1(1) => S910,
        out1 => S913
    );
nor_n_361: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S899,
        in1(1) => S892,
        out1 => S914
    );
nand_n_431: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S900,
        in1(1) => S893,
        out1 => S915
    );
nor_n_362: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S888,
        in1(1) => S882,
        out1 => S916
    );
notg_138: ENTITY WORK.notg
    PORT MAP (
        in1 => S916,
        out1 => S917
    );
nor_n_363: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S827,
        in1(1) => S823,
        out1 => S918
    );
notg_139: ENTITY WORK.notg
    PORT MAP (
        in1 => S918,
        out1 => S919
    );
nor_n_364: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S878,
        in1(1) => S870,
        out1 => S920
    );
nand_n_432: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S879,
        in1(1) => S871,
        out1 => S921
    );
nand_n_433: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_7,
        in1(1) => DP_AC_out_2,
        out1 => S922
    );
nand_n_434: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_6,
        in1(1) => DP_AC_out_3,
        out1 => S923
    );
nor_n_365: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S844,
        in1(1) => S838,
        out1 => S924
    );
nor_n_366: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S924,
        in1(1) => S923,
        out1 => S925
    );
notg_140: ENTITY WORK.notg
    PORT MAP (
        in1 => S925,
        out1 => S926
    );
nand_n_435: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S924,
        in1(1) => S923,
        out1 => S927
    );
nand_n_436: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S927,
        in1(1) => S926,
        out1 => S928
    );
nor_n_367: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S928,
        in1(1) => S922,
        out1 => S929
    );
notg_141: ENTITY WORK.notg
    PORT MAP (
        in1 => S929,
        out1 => S930
    );
nand_n_437: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S928,
        in1(1) => S922,
        out1 => S931
    );
notg_142: ENTITY WORK.notg
    PORT MAP (
        in1 => S931,
        out1 => S932
    );
nor_n_368: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S932,
        in1(1) => S929,
        out1 => S933
    );
nand_n_438: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S931,
        in1(1) => S930,
        out1 => S934
    );
nor_n_369: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S866,
        in1(1) => S858,
        out1 => S935
    );
nand_n_439: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S867,
        in1(1) => S859,
        out1 => S936
    );
nand_n_440: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_5,
        in1(1) => DP_AC_out_4,
        out1 => S937
    );
nand_n_441: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_6,
        in1(1) => DP_ARU1_in1_3,
        out1 => S938
    );
nand_n_442: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_6,
        in1(1) => DP_ARU1_in1_4,
        out1 => S939
    );
notg_143: ENTITY WORK.notg
    PORT MAP (
        in1 => S939,
        out1 => S940
    );
nor_n_370: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S939,
        in1(1) => S836,
        out1 => S941
    );
notg_144: ENTITY WORK.notg
    PORT MAP (
        in1 => S941,
        out1 => S942
    );
nand_n_443: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S938,
        in1(1) => S837,
        out1 => S943
    );
nand_n_444: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S943,
        in1(1) => S942,
        out1 => S944
    );
nand_n_445: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S944,
        in1(1) => S937,
        out1 => S945
    );
notg_145: ENTITY WORK.notg
    PORT MAP (
        in1 => S945,
        out1 => S946
    );
nor_n_371: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S944,
        in1(1) => S937,
        out1 => S947
    );
notg_146: ENTITY WORK.notg
    PORT MAP (
        in1 => S947,
        out1 => S948
    );
nor_n_372: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S947,
        in1(1) => S946,
        out1 => S949
    );
nand_n_446: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S948,
        in1(1) => S945,
        out1 => S950
    );
nor_n_373: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S852,
        in1(1) => S642,
        out1 => S951
    );
nand_n_447: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S851,
        in1(1) => S643,
        out1 => S952
    );
nor_n_374: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S951,
        in1(1) => S949,
        out1 => S953
    );
nand_n_448: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S952,
        in1(1) => S950,
        out1 => S954
    );
nor_n_375: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S952,
        in1(1) => S950,
        out1 => S955
    );
nand_n_449: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S951,
        in1(1) => S949,
        out1 => S956
    );
nor_n_376: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S955,
        in1(1) => S953,
        out1 => S957
    );
nand_n_450: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S956,
        in1(1) => S954,
        out1 => S958
    );
nor_n_377: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S958,
        in1(1) => S935,
        out1 => S959
    );
nand_n_451: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S957,
        in1(1) => S936,
        out1 => S960
    );
nor_n_378: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S957,
        in1(1) => S936,
        out1 => S961
    );
nand_n_452: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S958,
        in1(1) => S935,
        out1 => S962
    );
nor_n_379: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S961,
        in1(1) => S959,
        out1 => S963
    );
nand_n_453: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S962,
        in1(1) => S960,
        out1 => S964
    );
nor_n_380: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S963,
        in1(1) => S933,
        out1 => S965
    );
nand_n_454: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S964,
        in1(1) => S934,
        out1 => S967
    );
nor_n_381: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S964,
        in1(1) => S934,
        out1 => S968
    );
nand_n_455: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S963,
        in1(1) => S933,
        out1 => S969
    );
nor_n_382: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S968,
        in1(1) => S965,
        out1 => S970
    );
nand_n_456: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S969,
        in1(1) => S967,
        out1 => S971
    );
nand_n_457: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S970,
        in1(1) => S921,
        out1 => S972
    );
nand_n_458: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S971,
        in1(1) => S920,
        out1 => S973
    );
nand_n_459: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S973,
        in1(1) => S972,
        out1 => S974
    );
notg_147: ENTITY WORK.notg
    PORT MAP (
        in1 => S974,
        out1 => S975
    );
nand_n_460: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S975,
        in1(1) => S919,
        out1 => S976
    );
nand_n_461: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S974,
        in1(1) => S918,
        out1 => S978
    );
nand_n_462: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S978,
        in1(1) => S976,
        out1 => S979
    );
notg_148: ENTITY WORK.notg
    PORT MAP (
        in1 => S979,
        out1 => S980
    );
nand_n_463: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S979,
        in1(1) => S916,
        out1 => S981
    );
nand_n_464: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S980,
        in1(1) => S917,
        out1 => S982
    );
notg_149: ENTITY WORK.notg
    PORT MAP (
        in1 => S982,
        out1 => S983
    );
nand_n_465: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S982,
        in1(1) => S981,
        out1 => S984
    );
notg_150: ENTITY WORK.notg
    PORT MAP (
        in1 => S984,
        out1 => S985
    );
nor_n_383: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S985,
        in1(1) => S915,
        out1 => S986
    );
nor_n_384: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S984,
        in1(1) => S914,
        out1 => S987
    );
nand_n_466: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S985,
        in1(1) => S915,
        out1 => S989
    );
nor_n_385: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S987,
        in1(1) => S986,
        out1 => S990
    );
nor_n_386: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S990,
        in1(1) => CU_ADD,
        out1 => S991
    );
nor_n_387: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S913,
        in1(1) => S988,
        out1 => S992
    );
nor_n_388: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S992,
        in1(1) => S991,
        out1 => S336
    );
nor_n_389: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_10,
        in1(1) => DP_AC_out_10,
        out1 => S993
    );
nand_n_467: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_10,
        in1(1) => DP_AC_out_10,
        out1 => S994
    );
notg_151: ENTITY WORK.notg
    PORT MAP (
        in1 => S994,
        out1 => S995
    );
nor_n_390: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S995,
        in1(1) => S993,
        out1 => S996
    );
notg_152: ENTITY WORK.notg
    PORT MAP (
        in1 => S996,
        out1 => S997
    );
nand_n_468: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S907,
        in1(1) => S906,
        out1 => S999
    );
nand_n_469: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S999,
        in1(1) => S908,
        out1 => S1000
    );
notg_153: ENTITY WORK.notg
    PORT MAP (
        in1 => S1000,
        out1 => S1001
    );
nor_n_391: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1000,
        in1(1) => S996,
        out1 => S1002
    );
nor_n_392: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1001,
        in1(1) => S997,
        out1 => S1003
    );
notg_154: ENTITY WORK.notg
    PORT MAP (
        in1 => S1003,
        out1 => S1004
    );
nor_n_393: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1003,
        in1(1) => S1002,
        out1 => S1005
    );
nor_n_394: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1005,
        in1(1) => S988,
        out1 => S1006
    );
nor_n_395: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S987,
        in1(1) => S983,
        out1 => S1007
    );
nand_n_470: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S989,
        in1(1) => S982,
        out1 => S1008
    );
nand_n_471: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S976,
        in1(1) => S972,
        out1 => S1010
    );
notg_155: ENTITY WORK.notg
    PORT MAP (
        in1 => S1010,
        out1 => S1011
    );
nor_n_396: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S929,
        in1(1) => S925,
        out1 => S1012
    );
nor_n_397: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S968,
        in1(1) => S959,
        out1 => S1013
    );
nand_n_472: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_7,
        in1(1) => DP_AC_out_3,
        out1 => S1014
    );
nand_n_473: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_6,
        in1(1) => DP_AC_out_4,
        out1 => S1015
    );
nor_n_398: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S947,
        in1(1) => S941,
        out1 => S1016
    );
nor_n_399: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1016,
        in1(1) => S1015,
        out1 => S1017
    );
notg_156: ENTITY WORK.notg
    PORT MAP (
        in1 => S1017,
        out1 => S1018
    );
nand_n_474: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1016,
        in1(1) => S1015,
        out1 => S1019
    );
nand_n_475: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1019,
        in1(1) => S1018,
        out1 => S1021
    );
nor_n_400: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1021,
        in1(1) => S1014,
        out1 => S1022
    );
notg_157: ENTITY WORK.notg
    PORT MAP (
        in1 => S1022,
        out1 => S1023
    );
nand_n_476: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1021,
        in1(1) => S1014,
        out1 => S1024
    );
notg_158: ENTITY WORK.notg
    PORT MAP (
        in1 => S1024,
        out1 => S1025
    );
nor_n_401: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1025,
        in1(1) => S1022,
        out1 => S1026
    );
nand_n_477: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1024,
        in1(1) => S1023,
        out1 => S1027
    );
nor_n_402: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S955,
        in1(1) => S853,
        out1 => S1028
    );
nand_n_478: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S956,
        in1(1) => S854,
        out1 => S1029
    );
nand_n_479: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_7,
        in1(1) => DP_ARU1_in1_3,
        out1 => S1030
    );
nand_n_480: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1030,
        in1(1) => S939,
        out1 => S1032
    );
notg_159: ENTITY WORK.notg
    PORT MAP (
        in1 => S1032,
        out1 => S1033
    );
nand_n_481: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_7,
        in1(1) => DP_ARU1_in1_4,
        out1 => S1034
    );
nor_n_403: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1034,
        in1(1) => S938,
        out1 => S1035
    );
notg_160: ENTITY WORK.notg
    PORT MAP (
        in1 => S1035,
        out1 => S1036
    );
nor_n_404: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1035,
        in1(1) => S1033,
        out1 => S1037
    );
nand_n_482: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1036,
        in1(1) => S1032,
        out1 => S1038
    );
nor_n_405: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1037,
        in1(1) => S528,
        out1 => S1039
    );
nand_n_483: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1038,
        in1(1) => S529,
        out1 => S1040
    );
nor_n_406: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1038,
        in1(1) => S529,
        out1 => S1041
    );
notg_161: ENTITY WORK.notg
    PORT MAP (
        in1 => S1041,
        out1 => S1043
    );
nor_n_407: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1041,
        in1(1) => S1039,
        out1 => S1044
    );
nand_n_484: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1043,
        in1(1) => S1040,
        out1 => S1045
    );
nor_n_408: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1045,
        in1(1) => S1028,
        out1 => S1046
    );
nand_n_485: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1044,
        in1(1) => S1029,
        out1 => S1047
    );
nor_n_409: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1044,
        in1(1) => S1029,
        out1 => S1048
    );
nand_n_486: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1045,
        in1(1) => S1028,
        out1 => S1049
    );
nor_n_410: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1048,
        in1(1) => S1046,
        out1 => S1050
    );
nand_n_487: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1049,
        in1(1) => S1047,
        out1 => S1051
    );
nand_n_488: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1051,
        in1(1) => S1027,
        out1 => S1052
    );
nor_n_411: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1051,
        in1(1) => S1027,
        out1 => S1054
    );
nand_n_489: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1050,
        in1(1) => S1026,
        out1 => S1055
    );
nand_n_490: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1055,
        in1(1) => S1052,
        out1 => S1056
    );
nor_n_412: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1056,
        in1(1) => S1013,
        out1 => S1057
    );
notg_162: ENTITY WORK.notg
    PORT MAP (
        in1 => S1057,
        out1 => S1058
    );
nand_n_491: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1056,
        in1(1) => S1013,
        out1 => S1059
    );
nand_n_492: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1059,
        in1(1) => S1058,
        out1 => S1060
    );
nand_n_493: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1060,
        in1(1) => S1012,
        out1 => S1061
    );
notg_163: ENTITY WORK.notg
    PORT MAP (
        in1 => S1061,
        out1 => S1062
    );
nor_n_413: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1060,
        in1(1) => S1012,
        out1 => S1063
    );
nor_n_414: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1063,
        in1(1) => S1062,
        out1 => S1065
    );
notg_164: ENTITY WORK.notg
    PORT MAP (
        in1 => S1065,
        out1 => S1066
    );
nor_n_415: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1066,
        in1(1) => S1011,
        out1 => S1067
    );
notg_165: ENTITY WORK.notg
    PORT MAP (
        in1 => S1067,
        out1 => S1068
    );
nor_n_416: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1065,
        in1(1) => S1010,
        out1 => S1069
    );
nor_n_417: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1069,
        in1(1) => S1067,
        out1 => S1070
    );
notg_166: ENTITY WORK.notg
    PORT MAP (
        in1 => S1070,
        out1 => S1071
    );
nor_n_418: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1070,
        in1(1) => S1008,
        out1 => S1072
    );
nor_n_419: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1071,
        in1(1) => S1007,
        out1 => S1073
    );
nand_n_494: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1070,
        in1(1) => S1008,
        out1 => S1074
    );
nor_n_420: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1073,
        in1(1) => S1072,
        out1 => S1076
    );
nor_n_421: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1076,
        in1(1) => CU_ADD,
        out1 => S1077
    );
nor_n_422: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1077,
        in1(1) => S1006,
        out1 => S322
    );
nand_n_495: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1004,
        in1(1) => S994,
        out1 => S1078
    );
nand_n_496: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1183,
        in1(1) => S1172,
        out1 => S1079
    );
nand_n_497: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_11,
        in1(1) => DP_AC_out_11,
        out1 => S1080
    );
nand_n_498: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1080,
        in1(1) => S1079,
        out1 => S1081
    );
nand_n_499: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1081,
        in1(1) => S1078,
        out1 => S1082
    );
nor_n_423: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1081,
        in1(1) => S1078,
        out1 => S1083
    );
notg_167: ENTITY WORK.notg
    PORT MAP (
        in1 => S1083,
        out1 => S1084
    );
nand_n_500: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1084,
        in1(1) => S1082,
        out1 => S1086
    );
nor_n_424: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1073,
        in1(1) => S1067,
        out1 => S1087
    );
nand_n_501: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1074,
        in1(1) => S1068,
        out1 => S1088
    );
nor_n_425: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1063,
        in1(1) => S1057,
        out1 => S1089
    );
notg_168: ENTITY WORK.notg
    PORT MAP (
        in1 => S1089,
        out1 => S1090
    );
nor_n_426: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1022,
        in1(1) => S1017,
        out1 => S1091
    );
notg_169: ENTITY WORK.notg
    PORT MAP (
        in1 => S1091,
        out1 => S1092
    );
nor_n_427: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1054,
        in1(1) => S1046,
        out1 => S1093
    );
nand_n_502: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1055,
        in1(1) => S1047,
        out1 => S1094
    );
nand_n_503: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_7,
        in1(1) => DP_AC_out_4,
        out1 => S1095
    );
nand_n_504: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_6,
        in1(1) => DP_AC_out_5,
        out1 => S1097
    );
nor_n_428: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1041,
        in1(1) => S1035,
        out1 => S1098
    );
nor_n_429: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1098,
        in1(1) => S1097,
        out1 => S1099
    );
notg_170: ENTITY WORK.notg
    PORT MAP (
        in1 => S1099,
        out1 => S1100
    );
nand_n_505: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1098,
        in1(1) => S1097,
        out1 => S1101
    );
nand_n_506: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1101,
        in1(1) => S1100,
        out1 => S1102
    );
nor_n_430: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1102,
        in1(1) => S1095,
        out1 => S1103
    );
notg_171: ENTITY WORK.notg
    PORT MAP (
        in1 => S1103,
        out1 => S1104
    );
nand_n_507: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1102,
        in1(1) => S1095,
        out1 => S1105
    );
notg_172: ENTITY WORK.notg
    PORT MAP (
        in1 => S1105,
        out1 => S1106
    );
nor_n_431: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1106,
        in1(1) => S1103,
        out1 => S1108
    );
nand_n_508: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1105,
        in1(1) => S1104,
        out1 => S1109
    );
nand_n_509: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_6,
        in1(1) => DP_ARU1_in1_5,
        out1 => S1110
    );
nand_n_510: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1110,
        in1(1) => S1034,
        out1 => S1111
    );
notg_173: ENTITY WORK.notg
    PORT MAP (
        in1 => S1111,
        out1 => S1112
    );
nor_n_432: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1129,
        in1(1) => S1096,
        out1 => S1113
    );
nand_n_511: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_7,
        in1(1) => DP_ARU1_in1_5,
        out1 => S1114
    );
nor_n_433: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1114,
        in1(1) => S939,
        out1 => S1115
    );
nand_n_512: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1113,
        in1(1) => S940,
        out1 => S1116
    );
nor_n_434: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1115,
        in1(1) => S1112,
        out1 => S1117
    );
nand_n_513: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1116,
        in1(1) => S1111,
        out1 => S1119
    );
nand_n_514: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1119,
        in1(1) => S1109,
        out1 => S1120
    );
nor_n_435: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1119,
        in1(1) => S1109,
        out1 => S1121
    );
nand_n_515: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1117,
        in1(1) => S1108,
        out1 => S1122
    );
nand_n_516: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1122,
        in1(1) => S1120,
        out1 => S1123
    );
notg_174: ENTITY WORK.notg
    PORT MAP (
        in1 => S1123,
        out1 => S1124
    );
nand_n_517: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1124,
        in1(1) => S1094,
        out1 => S1125
    );
nand_n_518: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1123,
        in1(1) => S1093,
        out1 => S1126
    );
nand_n_519: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1126,
        in1(1) => S1125,
        out1 => S1127
    );
notg_175: ENTITY WORK.notg
    PORT MAP (
        in1 => S1127,
        out1 => S1128
    );
nand_n_520: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1127,
        in1(1) => S1091,
        out1 => S1130
    );
nand_n_521: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1128,
        in1(1) => S1092,
        out1 => S1131
    );
nand_n_522: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1131,
        in1(1) => S1130,
        out1 => S1132
    );
notg_176: ENTITY WORK.notg
    PORT MAP (
        in1 => S1132,
        out1 => S1133
    );
nand_n_523: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1133,
        in1(1) => S1090,
        out1 => S1134
    );
notg_177: ENTITY WORK.notg
    PORT MAP (
        in1 => S1134,
        out1 => S1135
    );
nand_n_524: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1132,
        in1(1) => S1089,
        out1 => S1136
    );
nand_n_525: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1136,
        in1(1) => S1134,
        out1 => S1137
    );
notg_178: ENTITY WORK.notg
    PORT MAP (
        in1 => S1137,
        out1 => S1138
    );
nor_n_436: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1138,
        in1(1) => S1088,
        out1 => S1139
    );
nor_n_437: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1137,
        in1(1) => S1087,
        out1 => S1141
    );
nand_n_526: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1138,
        in1(1) => S1088,
        out1 => S1142
    );
nor_n_438: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1141,
        in1(1) => S1139,
        out1 => S1143
    );
nor_n_439: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1143,
        in1(1) => CU_ADD,
        out1 => S1144
    );
nor_n_440: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1086,
        in1(1) => S988,
        out1 => S1145
    );
nor_n_441: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1145,
        in1(1) => S1144,
        out1 => S323
    );
nor_n_442: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_12,
        in1(1) => DP_AC_out_12,
        out1 => S1146
    );
nand_n_527: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_12,
        in1(1) => DP_AC_out_12,
        out1 => S1147
    );
notg_179: ENTITY WORK.notg
    PORT MAP (
        in1 => S1147,
        out1 => S1148
    );
nor_n_443: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1148,
        in1(1) => S1146,
        out1 => S1149
    );
nand_n_528: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1079,
        in1(1) => S1078,
        out1 => S1151
    );
nand_n_529: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1151,
        in1(1) => S1080,
        out1 => S1152
    );
nand_n_530: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1152,
        in1(1) => S1149,
        out1 => S1153
    );
nor_n_444: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1152,
        in1(1) => S1149,
        out1 => S1154
    );
nor_n_445: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1141,
        in1(1) => S1135,
        out1 => S1155
    );
nand_n_531: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1142,
        in1(1) => S1134,
        out1 => S1156
    );
nand_n_532: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1131,
        in1(1) => S1125,
        out1 => S1157
    );
notg_180: ENTITY WORK.notg
    PORT MAP (
        in1 => S1157,
        out1 => S1158
    );
nor_n_446: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1103,
        in1(1) => S1099,
        out1 => S1159
    );
nand_n_533: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_7,
        in1(1) => DP_AC_out_5,
        out1 => S1160
    );
notg_181: ENTITY WORK.notg
    PORT MAP (
        in1 => S1160,
        out1 => S1162
    );
nand_n_534: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1115,
        in1(1) => DP_ARU1_in1_6,
        out1 => S1163
    );
notg_182: ENTITY WORK.notg
    PORT MAP (
        in1 => S1163,
        out1 => S1164
    );
nand_n_535: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1116,
        in1(1) => S607,
        out1 => S1165
    );
nand_n_536: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1165,
        in1(1) => S1163,
        out1 => S1166
    );
notg_183: ENTITY WORK.notg
    PORT MAP (
        in1 => S1166,
        out1 => S1167
    );
nor_n_447: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1166,
        in1(1) => S1160,
        out1 => S1168
    );
nand_n_537: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1167,
        in1(1) => S1162,
        out1 => S1169
    );
nand_n_538: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1166,
        in1(1) => S1160,
        out1 => S1170
    );
notg_184: ENTITY WORK.notg
    PORT MAP (
        in1 => S1170,
        out1 => S1171
    );
nor_n_448: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1171,
        in1(1) => S1168,
        out1 => S1173
    );
nand_n_539: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1170,
        in1(1) => S1169,
        out1 => S1174
    );
nand_n_540: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1174,
        in1(1) => S1114,
        out1 => S1175
    );
nor_n_449: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1174,
        in1(1) => S1114,
        out1 => S1176
    );
nand_n_541: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1173,
        in1(1) => S1113,
        out1 => S1177
    );
nand_n_542: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1177,
        in1(1) => S1175,
        out1 => S1178
    );
notg_185: ENTITY WORK.notg
    PORT MAP (
        in1 => S1178,
        out1 => S1179
    );
nand_n_543: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1179,
        in1(1) => S1121,
        out1 => S1180
    );
notg_186: ENTITY WORK.notg
    PORT MAP (
        in1 => S1180,
        out1 => S1181
    );
nand_n_544: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1178,
        in1(1) => S1122,
        out1 => S1182
    );
nand_n_545: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1182,
        in1(1) => S1180,
        out1 => S1184
    );
nor_n_450: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1184,
        in1(1) => S1159,
        out1 => S1185
    );
notg_187: ENTITY WORK.notg
    PORT MAP (
        in1 => S1185,
        out1 => S1186
    );
nand_n_546: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1184,
        in1(1) => S1159,
        out1 => S1187
    );
notg_188: ENTITY WORK.notg
    PORT MAP (
        in1 => S1187,
        out1 => S1188
    );
nor_n_451: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1188,
        in1(1) => S1185,
        out1 => S1189
    );
notg_189: ENTITY WORK.notg
    PORT MAP (
        in1 => S1189,
        out1 => S1190
    );
nor_n_452: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1190,
        in1(1) => S1158,
        out1 => S1191
    );
notg_190: ENTITY WORK.notg
    PORT MAP (
        in1 => S1191,
        out1 => S1192
    );
nor_n_453: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1189,
        in1(1) => S1157,
        out1 => S1193
    );
nor_n_454: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1193,
        in1(1) => S1191,
        out1 => S1195
    );
notg_191: ENTITY WORK.notg
    PORT MAP (
        in1 => S1195,
        out1 => S1196
    );
nand_n_547: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1196,
        in1(1) => S1155,
        out1 => S1197
    );
notg_192: ENTITY WORK.notg
    PORT MAP (
        in1 => S1197,
        out1 => S1198
    );
nor_n_455: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1196,
        in1(1) => S1155,
        out1 => S1199
    );
nand_n_548: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1195,
        in1(1) => S1156,
        out1 => S1200
    );
nor_n_456: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1199,
        in1(1) => S1198,
        out1 => S1201
    );
nor_n_457: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1154,
        in1(1) => S988,
        out1 => S1202
    );
nand_n_549: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1202,
        in1(1) => S1153,
        out1 => S1203
    );
nand_n_550: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1201,
        in1(1) => S988,
        out1 => S1204
    );
nand_n_551: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1204,
        in1(1) => S1203,
        out1 => S324
    );
nand_n_552: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1153,
        in1(1) => S1147,
        out1 => S1206
    );
nand_n_553: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1205,
        in1(1) => S1194,
        out1 => S1207
    );
nand_n_554: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_13,
        in1(1) => DP_AC_out_13,
        out1 => S1208
    );
nand_n_555: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1208,
        in1(1) => S1207,
        out1 => S1209
    );
nand_n_556: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1209,
        in1(1) => S1206,
        out1 => S1210
    );
nor_n_458: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1209,
        in1(1) => S1206,
        out1 => S1211
    );
nor_n_459: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1199,
        in1(1) => S1191,
        out1 => S1212
    );
nand_n_557: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1200,
        in1(1) => S1192,
        out1 => S1213
    );
nor_n_460: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1185,
        in1(1) => S1181,
        out1 => S1214
    );
nand_n_558: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1186,
        in1(1) => S1180,
        out1 => S1216
    );
nor_n_461: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1168,
        in1(1) => S1164,
        out1 => S1217
    );
nand_n_559: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1169,
        in1(1) => S1163,
        out1 => S1218
    );
nand_n_560: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_7,
        in1(1) => DP_AC_out_6,
        out1 => S1219
    );
nand_n_561: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_7,
        in1(1) => DP_ARU1_in1_6,
        out1 => S1220
    );
nand_n_562: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1220,
        in1(1) => S1219,
        out1 => S1221
    );
notg_193: ENTITY WORK.notg
    PORT MAP (
        in1 => S1221,
        out1 => S1222
    );
nor_n_462: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S702,
        in1(1) => S607,
        out1 => S1223
    );
nand_n_563: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S701,
        in1(1) => S606,
        out1 => S1224
    );
nor_n_463: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1223,
        in1(1) => S1222,
        out1 => S1225
    );
nand_n_564: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1224,
        in1(1) => S1221,
        out1 => S1227
    );
nor_n_464: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1227,
        in1(1) => S1177,
        out1 => S1228
    );
nand_n_565: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1225,
        in1(1) => S1176,
        out1 => S1229
    );
nor_n_465: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1225,
        in1(1) => S1176,
        out1 => S1230
    );
nand_n_566: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1227,
        in1(1) => S1177,
        out1 => S1231
    );
nor_n_466: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1230,
        in1(1) => S1228,
        out1 => S1232
    );
nand_n_567: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1231,
        in1(1) => S1229,
        out1 => S1233
    );
nor_n_467: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1233,
        in1(1) => S1217,
        out1 => S1234
    );
nand_n_568: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1232,
        in1(1) => S1218,
        out1 => S1235
    );
nor_n_468: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1232,
        in1(1) => S1218,
        out1 => S1236
    );
nand_n_569: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1233,
        in1(1) => S1217,
        out1 => S1238
    );
nor_n_469: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1236,
        in1(1) => S1234,
        out1 => S1239
    );
nand_n_570: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1238,
        in1(1) => S1235,
        out1 => S1240
    );
nor_n_470: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1240,
        in1(1) => S1214,
        out1 => S1241
    );
nor_n_471: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1239,
        in1(1) => S1216,
        out1 => S1242
    );
nor_n_472: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1242,
        in1(1) => S1241,
        out1 => S1243
    );
nor_n_473: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1243,
        in1(1) => S1212,
        out1 => S1244
    );
nand_n_571: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1243,
        in1(1) => S1212,
        out1 => S1245
    );
nand_n_572: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1210,
        in1(1) => CU_ADD,
        out1 => S1246
    );
nor_n_474: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1246,
        in1(1) => S1211,
        out1 => S1247
    );
nand_n_573: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1245,
        in1(1) => S988,
        out1 => S1249
    );
nor_n_475: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1249,
        in1(1) => S1244,
        out1 => S1250
    );
nor_n_476: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1250,
        in1(1) => S1247,
        out1 => S325
    );
nor_n_477: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1234,
        in1(1) => S1228,
        out1 => S1251
    );
nand_n_574: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1235,
        in1(1) => S1229,
        out1 => S1252
    );
nor_n_478: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S702,
        in1(1) => S606,
        out1 => S1253
    );
nand_n_575: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S701,
        in1(1) => S607,
        out1 => S1254
    );
nand_n_576: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1253,
        in1(1) => S1252,
        out1 => S1255
    );
nand_n_577: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1254,
        in1(1) => S1251,
        out1 => S1256
    );
nand_n_578: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1256,
        in1(1) => S1255,
        out1 => S1257
    );
notg_194: ENTITY WORK.notg
    PORT MAP (
        in1 => S1257,
        out1 => S1259
    );
nor_n_479: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1242,
        in1(1) => S1212,
        out1 => S1260
    );
nor_n_480: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1241,
        in1(1) => S1213,
        out1 => S1261
    );
nor_n_481: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1260,
        in1(1) => S1241,
        out1 => S1262
    );
nor_n_482: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1261,
        in1(1) => S1242,
        out1 => S1263
    );
nand_n_579: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1262,
        in1(1) => S1257,
        out1 => S1264
    );
nor_n_483: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1262,
        in1(1) => S1257,
        out1 => S1265
    );
nand_n_580: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1263,
        in1(1) => S1259,
        out1 => S1266
    );
nor_n_484: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1265,
        in1(1) => CU_ADD,
        out1 => S1267
    );
nand_n_581: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1266,
        in1(1) => S988,
        out1 => S1268
    );
nand_n_582: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1267,
        in1(1) => S1264,
        out1 => S338
    );
nor_n_485: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => DP_ARU1_in1_14,
        in1(1) => DP_AC_out_14,
        out1 => S339
    );
nor_n_486: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1226,
        in1(1) => S1215,
        out1 => S340
    );
nor_n_487: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S340,
        in1(1) => S339,
        out1 => S341
    );
nand_n_583: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1207,
        in1(1) => S1206,
        out1 => S342
    );
nand_n_584: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S342,
        in1(1) => S1208,
        out1 => S343
    );
nor_n_488: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S343,
        in1(1) => S341,
        out1 => S344
    );
nand_n_585: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S343,
        in1(1) => S341,
        out1 => S345
    );
notg_195: ENTITY WORK.notg
    PORT MAP (
        in1 => S345,
        out1 => S346
    );
nor_n_489: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S344,
        in1(1) => S988,
        out1 => S347
    );
nand_n_586: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S347,
        in1(1) => S345,
        out1 => S349
    );
nand_n_587: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S349,
        in1(1) => S338,
        out1 => S326
    );
nand_n_588: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1255,
        in1(1) => S1224,
        out1 => S350
    );
nor_n_490: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S350,
        in1(1) => S1268,
        out1 => S351
    );
nor_n_491: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S346,
        in1(1) => S340,
        out1 => S352
    );
nor_n_492: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S371,
        in1(1) => S368,
        out1 => S353
    );
nor_n_493: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S353,
        in1(1) => S352,
        out1 => S354
    );
nand_n_589: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S353,
        in1(1) => S352,
        out1 => S355
    );
nand_n_590: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S355,
        in1(1) => CU_ADD,
        out1 => S356
    );
nor_n_494: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S356,
        in1(1) => S354,
        out1 => S357
    );
nor_n_495: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S357,
        in1(1) => S351,
        out1 => S327
    );
nor_n_496: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => CU_MUL,
        in1(1) => CU_ADD,
        out1 => S337
    );
nand_n_591: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S355,
        in1(1) => S370,
        out1 => S1270
    );
$_DLATCH_P__1: ENTITY WORK.$_DLATCH_P_
    PORT MAP (
        D => S1270,
        E => CU_ADD,
        Q => DP_ARU1_C
    );
$_DLATCH_N__3: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S321,
        E => S337,
        Q => DP_ARU1_out_0
    );
$_DLATCH_N__4: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S328,
        E => S337,
        Q => DP_ARU1_out_1
    );
$_DLATCH_N__5: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S329,
        E => S337,
        Q => DP_ARU1_out_2
    );
$_DLATCH_N__6: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S330,
        E => S337,
        Q => DP_ARU1_out_3
    );
$_DLATCH_N__7: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S331,
        E => S337,
        Q => DP_ARU1_out_4
    );
$_DLATCH_N__8: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S332,
        E => S337,
        Q => DP_ARU1_out_5
    );
$_DLATCH_N__9: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S333,
        E => S337,
        Q => DP_ARU1_out_6
    );
$_DLATCH_N__10: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S334,
        E => S337,
        Q => DP_ARU1_out_7
    );
$_DLATCH_N__11: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S335,
        E => S337,
        Q => DP_ARU1_out_8
    );
$_DLATCH_N__12: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S336,
        E => S337,
        Q => DP_ARU1_out_9
    );
$_DLATCH_N__13: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S322,
        E => S337,
        Q => DP_ARU1_out_10
    );
$_DLATCH_N__14: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S323,
        E => S337,
        Q => DP_ARU1_out_11
    );
$_DLATCH_N__15: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S324,
        E => S337,
        Q => DP_ARU1_out_12
    );
$_DLATCH_N__16: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S325,
        E => S337,
        Q => DP_ARU1_out_13
    );
$_DLATCH_N__17: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S326,
        E => S337,
        Q => DP_ARU1_out_14
    );
$_DLATCH_N__18: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S327,
        E => S337,
        Q => DP_ARU1_N
    );
notg_196: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_inst_0,
        out1 => S1290
    );
notg_197: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_LSB0E,
        out1 => S1291
    );
notg_198: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_conOF,
        out1 => S1292
    );
notg_199: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_inst_1,
        out1 => S1293
    );
notg_200: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_inst_2,
        out1 => S1294
    );
notg_201: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_inst_3,
        out1 => S1295
    );
notg_202: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_inst_4,
        out1 => S1296
    );
notg_203: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_SE12bits,
        out1 => S1297
    );
nor_n_497: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => CU_conOF,
        in1(1) => S1291,
        out1 => S1298
    );
nor_n_498: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1298,
        in1(1) => S1290,
        out1 => S1271
    );
nor_n_499: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1298,
        in1(1) => S1293,
        out1 => S1278
    );
nor_n_500: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1298,
        in1(1) => S1294,
        out1 => S1279
    );
nor_n_501: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1298,
        in1(1) => S1295,
        out1 => S1280
    );
nand_n_592: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1292,
        in1(1) => S1291,
        out1 => S1299
    );
nand_n_593: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_SE12bits,
        in1(1) => CU_inst_3,
        out1 => S1300
    );
nand_n_594: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_SE12bits,
        in1(1) => S1292,
        out1 => S1301
    );
nor_n_502: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1300,
        in1(1) => S1299,
        out1 => S1302
    );
notg_204: ENTITY WORK.notg
    PORT MAP (
        in1 => S1302,
        out1 => S1303
    );
nor_n_503: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1298,
        in1(1) => S1296,
        out1 => S1304
    );
nand_n_595: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1304,
        in1(1) => S1301,
        out1 => S1305
    );
nand_n_596: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1305,
        in1(1) => S1303,
        out1 => S1281
    );
nor_n_504: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1299,
        in1(1) => CU_SE12bits,
        out1 => S1306
    );
notg_205: ENTITY WORK.notg
    PORT MAP (
        in1 => S1306,
        out1 => S1307
    );
nand_n_597: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1306,
        in1(1) => CU_inst_5,
        out1 => S1308
    );
nand_n_598: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_inst_5,
        in1(1) => CU_conOF,
        out1 => S1309
    );
notg_206: ENTITY WORK.notg
    PORT MAP (
        in1 => S1309,
        out1 => S1310
    );
nor_n_505: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1310,
        in1(1) => S1302,
        out1 => S1311
    );
nand_n_599: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1311,
        in1(1) => S1308,
        out1 => S1282
    );
nand_n_600: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1306,
        in1(1) => CU_inst_6,
        out1 => S1312
    );
nand_n_601: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_inst_6,
        in1(1) => CU_conOF,
        out1 => S1313
    );
notg_207: ENTITY WORK.notg
    PORT MAP (
        in1 => S1313,
        out1 => S1314
    );
nor_n_506: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1314,
        in1(1) => S1302,
        out1 => S1315
    );
nand_n_602: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1315,
        in1(1) => S1312,
        out1 => S1283
    );
nand_n_603: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1306,
        in1(1) => CU_inst_7,
        out1 => S1316
    );
nand_n_604: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_inst_7,
        in1(1) => CU_conOF,
        out1 => S1317
    );
notg_208: ENTITY WORK.notg
    PORT MAP (
        in1 => S1317,
        out1 => S1318
    );
nor_n_507: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1318,
        in1(1) => S1302,
        out1 => S1319
    );
nand_n_605: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1319,
        in1(1) => S1316,
        out1 => S1284
    );
nand_n_606: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1306,
        in1(1) => CU_inst_8,
        out1 => S1320
    );
nand_n_607: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_inst_8,
        in1(1) => CU_conOF,
        out1 => S1321
    );
notg_209: ENTITY WORK.notg
    PORT MAP (
        in1 => S1321,
        out1 => S1322
    );
nor_n_508: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1322,
        in1(1) => S1302,
        out1 => S1323
    );
nand_n_608: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1323,
        in1(1) => S1320,
        out1 => S1285
    );
nand_n_609: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1306,
        in1(1) => CU_inst_9,
        out1 => S1324
    );
nand_n_610: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_inst_9,
        in1(1) => CU_conOF,
        out1 => S1325
    );
notg_210: ENTITY WORK.notg
    PORT MAP (
        in1 => S1325,
        out1 => S1326
    );
nor_n_509: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1326,
        in1(1) => S1302,
        out1 => S1327
    );
nand_n_611: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1327,
        in1(1) => S1324,
        out1 => S1286
    );
nand_n_612: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1306,
        in1(1) => CU_inst_10,
        out1 => S1328
    );
nand_n_613: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_inst_10,
        in1(1) => CU_conOF,
        out1 => S1329
    );
notg_211: ENTITY WORK.notg
    PORT MAP (
        in1 => S1329,
        out1 => S1330
    );
nor_n_510: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1330,
        in1(1) => S1302,
        out1 => S1331
    );
nand_n_614: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1331,
        in1(1) => S1328,
        out1 => S1272
    );
nand_n_615: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_inst_11,
        in1(1) => CU_conOF,
        out1 => S1332
    );
nand_n_616: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_inst_11,
        in1(1) => S1297,
        out1 => S1333
    );
nor_n_511: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1333,
        in1(1) => S1299,
        out1 => S1334
    );
nor_n_512: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1334,
        in1(1) => S1302,
        out1 => S1335
    );
nand_n_617: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1335,
        in1(1) => S1332,
        out1 => S1273
    );
nand_n_618: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1299,
        in1(1) => DP_IMM1_in1_0,
        out1 => S1336
    );
nand_n_619: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1336,
        in1(1) => S1335,
        out1 => S1274
    );
nand_n_620: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1299,
        in1(1) => DP_IMM1_in1_1,
        out1 => S1337
    );
nand_n_621: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1337,
        in1(1) => S1335,
        out1 => S1275
    );
nand_n_622: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1299,
        in1(1) => DP_IMM1_in1_2,
        out1 => S1288
    );
nand_n_623: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1288,
        in1(1) => S1335,
        out1 => S1276
    );
nand_n_624: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1299,
        in1(1) => DP_IMM1_in1_3,
        out1 => S1289
    );
nand_n_625: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1289,
        in1(1) => S1335,
        out1 => S1277
    );
nor_n_513: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1307,
        in1(1) => CU_SE4bits,
        out1 => S1287
    );
$_DLATCH_N__19: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S1271,
        E => S1287,
        Q => DP_IMM1_out_0
    );
$_DLATCH_N__20: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S1278,
        E => S1287,
        Q => DP_IMM1_out_1
    );
$_DLATCH_N__21: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S1279,
        E => S1287,
        Q => DP_IMM1_out_2
    );
$_DLATCH_N__22: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S1280,
        E => S1287,
        Q => DP_IMM1_out_3
    );
$_DLATCH_N__23: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S1281,
        E => S1287,
        Q => DP_IMM1_out_4
    );
$_DLATCH_N__24: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S1282,
        E => S1287,
        Q => DP_IMM1_out_5
    );
$_DLATCH_N__25: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S1283,
        E => S1287,
        Q => DP_IMM1_out_6
    );
$_DLATCH_N__26: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S1284,
        E => S1287,
        Q => DP_IMM1_out_7
    );
$_DLATCH_N__27: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S1285,
        E => S1287,
        Q => DP_IMM1_out_8
    );
$_DLATCH_N__28: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S1286,
        E => S1287,
        Q => DP_IMM1_out_9
    );
$_DLATCH_N__29: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S1272,
        E => S1287,
        Q => DP_IMM1_out_10
    );
$_DLATCH_N__30: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S1273,
        E => S1287,
        Q => DP_IMM1_out_11
    );
$_DLATCH_N__31: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S1274,
        E => S1287,
        Q => DP_IMM1_out_12
    );
$_DLATCH_N__32: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S1275,
        E => S1287,
        Q => DP_IMM1_out_13
    );
$_DLATCH_N__33: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S1276,
        E => S1287,
        Q => DP_IMM1_out_14
    );
$_DLATCH_N__34: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S1277,
        E => S1287,
        Q => DP_IMM1_out_15
    );
notg_212: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_ldIN,
        out1 => S1355
    );
nor_n_514: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => CU_ldIN,
        in1(1) => S6,
        out1 => S1356
    );
nand_n_626: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1356,
        in1(1) => DP_IN_out_0,
        out1 => S1357
    );
nor_n_515: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1355,
        in1(1) => S7,
        out1 => S1358
    );
nand_n_627: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1358,
        in1(1) => DP_IN_in_0,
        out1 => S1359
    );
nand_n_628: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1359,
        in1(1) => S1357,
        out1 => S1338
    );
nand_n_629: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1356,
        in1(1) => DP_IN_out_1,
        out1 => S1360
    );
nand_n_630: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1358,
        in1(1) => DP_IN_in_1,
        out1 => S1361
    );
nand_n_631: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1361,
        in1(1) => S1360,
        out1 => S1339
    );
nand_n_632: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1356,
        in1(1) => DP_IN_out_2,
        out1 => S1362
    );
nand_n_633: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1358,
        in1(1) => DP_IN_in_2,
        out1 => S1363
    );
nand_n_634: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1363,
        in1(1) => S1362,
        out1 => S1340
    );
nand_n_635: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1356,
        in1(1) => DP_IN_out_3,
        out1 => S1364
    );
nand_n_636: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1358,
        in1(1) => DP_IN_in_3,
        out1 => S1365
    );
nand_n_637: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1365,
        in1(1) => S1364,
        out1 => S1341
    );
nand_n_638: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1356,
        in1(1) => DP_IN_out_4,
        out1 => S1366
    );
nand_n_639: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1358,
        in1(1) => DP_IN_in_4,
        out1 => S1367
    );
nand_n_640: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1367,
        in1(1) => S1366,
        out1 => S1342
    );
nand_n_641: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1356,
        in1(1) => DP_IN_out_5,
        out1 => S1368
    );
nand_n_642: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1358,
        in1(1) => DP_IN_in_5,
        out1 => S1369
    );
nand_n_643: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1369,
        in1(1) => S1368,
        out1 => S1343
    );
nand_n_644: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1356,
        in1(1) => DP_IN_out_6,
        out1 => S1370
    );
nand_n_645: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1358,
        in1(1) => DP_IN_in_6,
        out1 => S1371
    );
nand_n_646: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1371,
        in1(1) => S1370,
        out1 => S1344
    );
nand_n_647: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1356,
        in1(1) => DP_IN_out_7,
        out1 => S1372
    );
nand_n_648: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1358,
        in1(1) => DP_IN_in_7,
        out1 => S1373
    );
nand_n_649: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1373,
        in1(1) => S1372,
        out1 => S1345
    );
nand_n_650: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1356,
        in1(1) => DP_IN_out_8,
        out1 => S1374
    );
nand_n_651: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1358,
        in1(1) => DP_IN_in_8,
        out1 => S1375
    );
nand_n_652: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1375,
        in1(1) => S1374,
        out1 => S1346
    );
nand_n_653: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1356,
        in1(1) => DP_IN_out_9,
        out1 => S1376
    );
nand_n_654: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1358,
        in1(1) => DP_IN_in_9,
        out1 => S1377
    );
nand_n_655: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1377,
        in1(1) => S1376,
        out1 => S1347
    );
nand_n_656: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1356,
        in1(1) => DP_IN_out_10,
        out1 => S1378
    );
nand_n_657: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1358,
        in1(1) => DP_IN_in_10,
        out1 => S1379
    );
nand_n_658: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1379,
        in1(1) => S1378,
        out1 => S1348
    );
nand_n_659: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1356,
        in1(1) => DP_IN_out_11,
        out1 => S1380
    );
nand_n_660: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1358,
        in1(1) => DP_IN_in_11,
        out1 => S1381
    );
nand_n_661: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1381,
        in1(1) => S1380,
        out1 => S1349
    );
nand_n_662: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1356,
        in1(1) => DP_IN_out_12,
        out1 => S1382
    );
nand_n_663: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1358,
        in1(1) => DP_IN_in_12,
        out1 => S1383
    );
nand_n_664: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1383,
        in1(1) => S1382,
        out1 => S1350
    );
nand_n_665: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1356,
        in1(1) => DP_IN_out_13,
        out1 => S1384
    );
nand_n_666: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1358,
        in1(1) => DP_IN_in_13,
        out1 => S1385
    );
nand_n_667: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1385,
        in1(1) => S1384,
        out1 => S1351
    );
nand_n_668: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1356,
        in1(1) => DP_IN_out_14,
        out1 => S1386
    );
nand_n_669: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1358,
        in1(1) => DP_IN_in_14,
        out1 => S1387
    );
nand_n_670: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1387,
        in1(1) => S1386,
        out1 => S1352
    );
nand_n_671: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1356,
        in1(1) => DP_IN_out_15,
        out1 => S1388
    );
nand_n_672: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1358,
        in1(1) => DP_IN_in_15,
        out1 => S1354
    );
nand_n_673: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1354,
        in1(1) => S1388,
        out1 => S1353
    );
dff_19: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S1338,
        NbarT => '0',
        PRE => '0',
        Q => DP_IN_out_0,
        Si => S3322,
        global_reset => '0'
    );
dff_20: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S1339,
        NbarT => '0',
        PRE => '0',
        Q => DP_IN_out_1,
        Si => S3321,
        global_reset => '0'
    );
dff_21: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S1340,
        NbarT => '0',
        PRE => '0',
        Q => DP_IN_out_2,
        Si => S3320,
        global_reset => '0'
    );
dff_22: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S1341,
        NbarT => '0',
        PRE => '0',
        Q => DP_IN_out_3,
        Si => S3319,
        global_reset => '0'
    );
dff_23: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S1342,
        NbarT => '0',
        PRE => '0',
        Q => DP_IN_out_4,
        Si => S3318,
        global_reset => '0'
    );
dff_24: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S1343,
        NbarT => '0',
        PRE => '0',
        Q => DP_IN_out_5,
        Si => S3317,
        global_reset => '0'
    );
dff_25: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S1344,
        NbarT => '0',
        PRE => '0',
        Q => DP_IN_out_6,
        Si => S3316,
        global_reset => '0'
    );
dff_26: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S1345,
        NbarT => '0',
        PRE => '0',
        Q => DP_IN_out_7,
        Si => S3315,
        global_reset => '0'
    );
dff_27: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S1346,
        NbarT => '0',
        PRE => '0',
        Q => DP_IN_out_8,
        Si => S3314,
        global_reset => '0'
    );
dff_28: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S1347,
        NbarT => '0',
        PRE => '0',
        Q => DP_IN_out_9,
        Si => S3313,
        global_reset => '0'
    );
dff_29: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S1348,
        NbarT => '0',
        PRE => '0',
        Q => DP_IN_out_10,
        Si => S3312,
        global_reset => '0'
    );
dff_30: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S1349,
        NbarT => '0',
        PRE => '0',
        Q => DP_IN_out_11,
        Si => S3311,
        global_reset => '0'
    );
dff_31: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S1350,
        NbarT => '0',
        PRE => '0',
        Q => DP_IN_out_12,
        Si => S3310,
        global_reset => '0'
    );
dff_32: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S1351,
        NbarT => '0',
        PRE => '0',
        Q => DP_IN_out_13,
        Si => S3309,
        global_reset => '0'
    );
dff_33: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S1352,
        NbarT => '0',
        PRE => '0',
        Q => DP_IN_out_14,
        Si => S3308,
        global_reset => '0'
    );
dff_34: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S1353,
        NbarT => '0',
        PRE => '0',
        Q => DP_IN_out_15,
        Si => S3357,
        global_reset => '0'
    );
notg_213: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_in_0,
        out1 => S1406
    );
notg_214: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_inc_val_0,
        out1 => S1407
    );
notg_215: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_in_1,
        out1 => S1408
    );
notg_216: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_inc_val_1,
        out1 => S1409
    );
notg_217: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_in_2,
        out1 => S1410
    );
notg_218: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_in_3,
        out1 => S1411
    );
notg_219: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_in_4,
        out1 => S1412
    );
notg_220: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_in_5,
        out1 => S1413
    );
notg_221: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_in_6,
        out1 => S1414
    );
notg_222: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_in_7,
        out1 => S1415
    );
notg_223: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_in_8,
        out1 => S1416
    );
notg_224: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_in_9,
        out1 => S1417
    );
notg_225: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_in_10,
        out1 => S1418
    );
notg_226: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_in_11,
        out1 => S1419
    );
notg_227: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_in_12,
        out1 => S1420
    );
notg_228: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_in_13,
        out1 => S1421
    );
notg_229: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_in_14,
        out1 => S1422
    );
notg_230: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_in_15,
        out1 => S1423
    );
nor_n_516: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1407,
        in1(1) => S1406,
        out1 => S1424
    );
nand_n_674: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_INC_1_inc_val_0,
        in1(1) => DP_INC_1_in_0,
        out1 => S1425
    );
nor_n_517: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => DP_INC_1_inc_val_0,
        in1(1) => DP_INC_1_in_0,
        out1 => S1426
    );
nor_n_518: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1426,
        in1(1) => S1424,
        out1 => DP_INC_1_out_0
    );
nor_n_519: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1409,
        in1(1) => S1408,
        out1 => S1427
    );
nand_n_675: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_INC_1_inc_val_1,
        in1(1) => DP_INC_1_in_1,
        out1 => S1428
    );
nor_n_520: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => DP_INC_1_inc_val_1,
        in1(1) => DP_INC_1_in_1,
        out1 => S1429
    );
notg_231: ENTITY WORK.notg
    PORT MAP (
        in1 => S1429,
        out1 => S1430
    );
nor_n_521: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1429,
        in1(1) => S1427,
        out1 => S1431
    );
nand_n_676: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1430,
        in1(1) => S1428,
        out1 => S1432
    );
nor_n_522: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1432,
        in1(1) => S1425,
        out1 => S1433
    );
nand_n_677: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1431,
        in1(1) => S1424,
        out1 => S1434
    );
nor_n_523: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1431,
        in1(1) => S1424,
        out1 => S1435
    );
nor_n_524: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1435,
        in1(1) => S1433,
        out1 => DP_INC_1_out_1
    );
nor_n_525: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1433,
        in1(1) => S1427,
        out1 => S1436
    );
nand_n_678: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1434,
        in1(1) => S1428,
        out1 => S1437
    );
nor_n_526: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1436,
        in1(1) => S1410,
        out1 => S1438
    );
nand_n_679: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1437,
        in1(1) => DP_INC_1_in_2,
        out1 => S1439
    );
nor_n_527: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1437,
        in1(1) => DP_INC_1_in_2,
        out1 => S1440
    );
nor_n_528: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1440,
        in1(1) => S1438,
        out1 => DP_INC_1_out_2
    );
nor_n_529: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1439,
        in1(1) => S1411,
        out1 => S1441
    );
nand_n_680: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1438,
        in1(1) => DP_INC_1_in_3,
        out1 => S1442
    );
nor_n_530: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1438,
        in1(1) => DP_INC_1_in_3,
        out1 => S1443
    );
nor_n_531: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1443,
        in1(1) => S1441,
        out1 => DP_INC_1_out_3
    );
nor_n_532: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1442,
        in1(1) => S1412,
        out1 => S1444
    );
nand_n_681: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1441,
        in1(1) => DP_INC_1_in_4,
        out1 => S1445
    );
nor_n_533: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1441,
        in1(1) => DP_INC_1_in_4,
        out1 => S1446
    );
nor_n_534: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1446,
        in1(1) => S1444,
        out1 => DP_INC_1_out_4
    );
nor_n_535: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1445,
        in1(1) => S1413,
        out1 => S1447
    );
nand_n_682: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1444,
        in1(1) => DP_INC_1_in_5,
        out1 => S1448
    );
nor_n_536: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1444,
        in1(1) => DP_INC_1_in_5,
        out1 => S1449
    );
nor_n_537: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1449,
        in1(1) => S1447,
        out1 => DP_INC_1_out_5
    );
nor_n_538: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1448,
        in1(1) => S1414,
        out1 => S1450
    );
nand_n_683: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1447,
        in1(1) => DP_INC_1_in_6,
        out1 => S1451
    );
nor_n_539: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1447,
        in1(1) => DP_INC_1_in_6,
        out1 => S1452
    );
nor_n_540: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1452,
        in1(1) => S1450,
        out1 => DP_INC_1_out_6
    );
nor_n_541: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1451,
        in1(1) => S1415,
        out1 => S1453
    );
nand_n_684: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1450,
        in1(1) => DP_INC_1_in_7,
        out1 => S1454
    );
nor_n_542: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1450,
        in1(1) => DP_INC_1_in_7,
        out1 => S1455
    );
nor_n_543: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1455,
        in1(1) => S1453,
        out1 => DP_INC_1_out_7
    );
nor_n_544: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1454,
        in1(1) => S1416,
        out1 => S1456
    );
nand_n_685: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1453,
        in1(1) => DP_INC_1_in_8,
        out1 => S1457
    );
nor_n_545: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1453,
        in1(1) => DP_INC_1_in_8,
        out1 => S1458
    );
nor_n_546: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1458,
        in1(1) => S1456,
        out1 => DP_INC_1_out_8
    );
nor_n_547: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1457,
        in1(1) => S1417,
        out1 => S1459
    );
nand_n_686: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1456,
        in1(1) => DP_INC_1_in_9,
        out1 => S1460
    );
nor_n_548: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1456,
        in1(1) => DP_INC_1_in_9,
        out1 => S1461
    );
nor_n_549: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1461,
        in1(1) => S1459,
        out1 => DP_INC_1_out_9
    );
nor_n_550: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1460,
        in1(1) => S1418,
        out1 => S1389
    );
nand_n_687: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1459,
        in1(1) => DP_INC_1_in_10,
        out1 => S1390
    );
nor_n_551: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1459,
        in1(1) => DP_INC_1_in_10,
        out1 => S1391
    );
nor_n_552: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1391,
        in1(1) => S1389,
        out1 => DP_INC_1_out_10
    );
nor_n_553: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1390,
        in1(1) => S1419,
        out1 => S1392
    );
nand_n_688: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1389,
        in1(1) => DP_INC_1_in_11,
        out1 => S1393
    );
nor_n_554: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1389,
        in1(1) => DP_INC_1_in_11,
        out1 => S1394
    );
nor_n_555: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1394,
        in1(1) => S1392,
        out1 => DP_INC_1_out_11
    );
nor_n_556: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1393,
        in1(1) => S1420,
        out1 => S1395
    );
nand_n_689: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1392,
        in1(1) => DP_INC_1_in_12,
        out1 => S1396
    );
nor_n_557: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1392,
        in1(1) => DP_INC_1_in_12,
        out1 => S1397
    );
nor_n_558: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1397,
        in1(1) => S1395,
        out1 => DP_INC_1_out_12
    );
nor_n_559: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1396,
        in1(1) => S1421,
        out1 => S1398
    );
nand_n_690: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1395,
        in1(1) => DP_INC_1_in_13,
        out1 => S1399
    );
nor_n_560: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1395,
        in1(1) => DP_INC_1_in_13,
        out1 => S1400
    );
nor_n_561: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1400,
        in1(1) => S1398,
        out1 => DP_INC_1_out_13
    );
nor_n_562: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1399,
        in1(1) => S1422,
        out1 => S1401
    );
nand_n_691: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1398,
        in1(1) => DP_INC_1_in_14,
        out1 => S1402
    );
nor_n_563: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1398,
        in1(1) => DP_INC_1_in_14,
        out1 => S1403
    );
nor_n_564: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1403,
        in1(1) => S1401,
        out1 => DP_INC_1_out_14
    );
nor_n_565: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1401,
        in1(1) => DP_INC_1_in_15,
        out1 => S1404
    );
nor_n_566: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1402,
        in1(1) => S1423,
        out1 => S1405
    );
nor_n_567: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1405,
        in1(1) => S1404,
        out1 => DP_INC_1_out_15
    );
notg_232: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(0),
        out1 => S1479
    );
notg_233: ENTITY WORK.notg
    PORT MAP (
        in1 => S0,
        out1 => S1480
    );
notg_234: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(1),
        out1 => S1481
    );
notg_235: ENTITY WORK.notg
    PORT MAP (
        in1 => S8,
        out1 => S1482
    );
notg_236: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(2),
        out1 => S1483
    );
notg_237: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(3),
        out1 => S1484
    );
notg_238: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(4),
        out1 => S1485
    );
notg_239: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(5),
        out1 => S1486
    );
notg_240: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(6),
        out1 => S1487
    );
notg_241: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(7),
        out1 => S1488
    );
notg_242: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(8),
        out1 => S1489
    );
notg_243: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(9),
        out1 => S1490
    );
notg_244: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(10),
        out1 => S1491
    );
notg_245: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(11),
        out1 => S1492
    );
notg_246: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(12),
        out1 => S1493
    );
notg_247: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(13),
        out1 => S1494
    );
notg_248: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(14),
        out1 => S1495
    );
notg_249: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(15),
        out1 => S1496
    );
nor_n_568: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1480,
        in1(1) => S1479,
        out1 => S1497
    );
nand_n_692: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1,
        in1(1) => dataBus(0),
        out1 => S1498
    );
nor_n_569: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2,
        in1(1) => dataBus(0),
        out1 => S1499
    );
nor_n_570: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1499,
        in1(1) => S1497,
        out1 => DP_INC2_out_0
    );
nor_n_571: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1482,
        in1(1) => S1481,
        out1 => S1500
    );
nand_n_693: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S9,
        in1(1) => dataBus(1),
        out1 => S1501
    );
nor_n_572: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S10,
        in1(1) => dataBus(1),
        out1 => S1502
    );
notg_250: ENTITY WORK.notg
    PORT MAP (
        in1 => S1502,
        out1 => S1503
    );
nor_n_573: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1502,
        in1(1) => S1500,
        out1 => S1504
    );
nand_n_694: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1503,
        in1(1) => S1501,
        out1 => S1505
    );
nor_n_574: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1505,
        in1(1) => S1498,
        out1 => S1506
    );
nand_n_695: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1504,
        in1(1) => S1497,
        out1 => S1507
    );
nor_n_575: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1504,
        in1(1) => S1497,
        out1 => S1508
    );
nor_n_576: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1508,
        in1(1) => S1506,
        out1 => DP_INC2_out_1
    );
nor_n_577: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1506,
        in1(1) => S1500,
        out1 => S1509
    );
nand_n_696: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1507,
        in1(1) => S1501,
        out1 => S1510
    );
nor_n_578: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1509,
        in1(1) => S1483,
        out1 => S1511
    );
nand_n_697: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1510,
        in1(1) => dataBus(2),
        out1 => S1512
    );
nor_n_579: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1510,
        in1(1) => dataBus(2),
        out1 => S1513
    );
nor_n_580: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1513,
        in1(1) => S1511,
        out1 => DP_INC2_out_2
    );
nor_n_581: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1512,
        in1(1) => S1484,
        out1 => S1514
    );
nand_n_698: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1511,
        in1(1) => dataBus(3),
        out1 => S1515
    );
nor_n_582: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1511,
        in1(1) => dataBus(3),
        out1 => S1516
    );
nor_n_583: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1516,
        in1(1) => S1514,
        out1 => DP_INC2_out_3
    );
nor_n_584: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1515,
        in1(1) => S1485,
        out1 => S1517
    );
nand_n_699: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1514,
        in1(1) => dataBus(4),
        out1 => S1518
    );
nor_n_585: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1514,
        in1(1) => dataBus(4),
        out1 => S1519
    );
nor_n_586: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1519,
        in1(1) => S1517,
        out1 => DP_INC2_out_4
    );
nor_n_587: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1518,
        in1(1) => S1486,
        out1 => S1520
    );
nand_n_700: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1517,
        in1(1) => dataBus(5),
        out1 => S1521
    );
nor_n_588: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1517,
        in1(1) => dataBus(5),
        out1 => S1522
    );
nor_n_589: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1522,
        in1(1) => S1520,
        out1 => DP_INC2_out_5
    );
nor_n_590: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1521,
        in1(1) => S1487,
        out1 => S1523
    );
nand_n_701: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1520,
        in1(1) => dataBus(6),
        out1 => S1524
    );
nor_n_591: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1520,
        in1(1) => dataBus(6),
        out1 => S1525
    );
nor_n_592: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1525,
        in1(1) => S1523,
        out1 => DP_INC2_out_6
    );
nor_n_593: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1524,
        in1(1) => S1488,
        out1 => S1526
    );
nand_n_702: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1523,
        in1(1) => dataBus(7),
        out1 => S1527
    );
nor_n_594: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1523,
        in1(1) => dataBus(7),
        out1 => S1528
    );
nor_n_595: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1528,
        in1(1) => S1526,
        out1 => DP_INC2_out_7
    );
nor_n_596: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1527,
        in1(1) => S1489,
        out1 => S1529
    );
nand_n_703: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1526,
        in1(1) => dataBus(8),
        out1 => S1530
    );
nor_n_597: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1526,
        in1(1) => dataBus(8),
        out1 => S1531
    );
nor_n_598: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1531,
        in1(1) => S1529,
        out1 => DP_INC2_out_8
    );
nor_n_599: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1530,
        in1(1) => S1490,
        out1 => S1532
    );
nand_n_704: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1529,
        in1(1) => dataBus(9),
        out1 => S1533
    );
nor_n_600: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1529,
        in1(1) => dataBus(9),
        out1 => S1534
    );
nor_n_601: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1534,
        in1(1) => S1532,
        out1 => DP_INC2_out_9
    );
nor_n_602: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1533,
        in1(1) => S1491,
        out1 => S1462
    );
nand_n_705: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1532,
        in1(1) => dataBus(10),
        out1 => S1463
    );
nor_n_603: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1532,
        in1(1) => dataBus(10),
        out1 => S1464
    );
nor_n_604: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1464,
        in1(1) => S1462,
        out1 => DP_INC2_out_10
    );
nor_n_605: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1463,
        in1(1) => S1492,
        out1 => S1465
    );
nand_n_706: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1462,
        in1(1) => dataBus(11),
        out1 => S1466
    );
nor_n_606: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1462,
        in1(1) => dataBus(11),
        out1 => S1467
    );
nor_n_607: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1467,
        in1(1) => S1465,
        out1 => DP_INC2_out_11
    );
nor_n_608: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1466,
        in1(1) => S1493,
        out1 => S1468
    );
nand_n_707: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1465,
        in1(1) => dataBus(12),
        out1 => S1469
    );
nor_n_609: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1465,
        in1(1) => dataBus(12),
        out1 => S1470
    );
nor_n_610: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1470,
        in1(1) => S1468,
        out1 => DP_INC2_out_12
    );
nor_n_611: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1469,
        in1(1) => S1494,
        out1 => S1471
    );
nand_n_708: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1468,
        in1(1) => dataBus(13),
        out1 => S1472
    );
nor_n_612: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1468,
        in1(1) => dataBus(13),
        out1 => S1473
    );
nor_n_613: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1473,
        in1(1) => S1471,
        out1 => DP_INC2_out_13
    );
nor_n_614: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1472,
        in1(1) => S1495,
        out1 => S1474
    );
nand_n_709: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1471,
        in1(1) => dataBus(14),
        out1 => S1475
    );
nor_n_615: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1471,
        in1(1) => dataBus(14),
        out1 => S1476
    );
nor_n_616: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1476,
        in1(1) => S1474,
        out1 => DP_INC2_out_14
    );
nor_n_617: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1474,
        in1(1) => dataBus(15),
        out1 => S1477
    );
nor_n_618: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1475,
        in1(1) => S1496,
        out1 => S1478
    );
nor_n_619: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1478,
        in1(1) => S1477,
        out1 => DP_INC2_out_15
    );
notg_251: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_ldIR,
        out1 => S1552
    );
nor_n_620: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => CU_ldIR,
        in1(1) => S11,
        out1 => S1553
    );
nand_n_710: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1553,
        in1(1) => CU_inst_0,
        out1 => S1554
    );
nor_n_621: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1552,
        in1(1) => S12,
        out1 => S1555
    );
nand_n_711: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1555,
        in1(1) => dataBus(0),
        out1 => S1556
    );
nand_n_712: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1556,
        in1(1) => S1554,
        out1 => S1535
    );
nand_n_713: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1553,
        in1(1) => CU_inst_1,
        out1 => S1557
    );
nand_n_714: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1555,
        in1(1) => dataBus(1),
        out1 => S1558
    );
nand_n_715: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1558,
        in1(1) => S1557,
        out1 => S1536
    );
nand_n_716: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1553,
        in1(1) => CU_inst_2,
        out1 => S1559
    );
nand_n_717: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1555,
        in1(1) => dataBus(2),
        out1 => S1560
    );
nand_n_718: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1560,
        in1(1) => S1559,
        out1 => S1537
    );
nand_n_719: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1553,
        in1(1) => CU_inst_3,
        out1 => S1561
    );
nand_n_720: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1555,
        in1(1) => dataBus(3),
        out1 => S1562
    );
nand_n_721: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1562,
        in1(1) => S1561,
        out1 => S1538
    );
nand_n_722: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1553,
        in1(1) => CU_inst_4,
        out1 => S1563
    );
nand_n_723: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1555,
        in1(1) => dataBus(4),
        out1 => S1564
    );
nand_n_724: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1564,
        in1(1) => S1563,
        out1 => S1539
    );
nand_n_725: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1553,
        in1(1) => CU_inst_5,
        out1 => S1565
    );
nand_n_726: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1555,
        in1(1) => dataBus(5),
        out1 => S1566
    );
nand_n_727: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1566,
        in1(1) => S1565,
        out1 => S1540
    );
nand_n_728: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1553,
        in1(1) => CU_inst_6,
        out1 => S1567
    );
nand_n_729: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1555,
        in1(1) => dataBus(6),
        out1 => S1568
    );
nand_n_730: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1568,
        in1(1) => S1567,
        out1 => S1541
    );
nand_n_731: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1553,
        in1(1) => CU_inst_7,
        out1 => S1569
    );
nand_n_732: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1555,
        in1(1) => dataBus(7),
        out1 => S1570
    );
nand_n_733: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1570,
        in1(1) => S1569,
        out1 => S1542
    );
nand_n_734: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1553,
        in1(1) => CU_inst_8,
        out1 => S1571
    );
nand_n_735: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1555,
        in1(1) => dataBus(8),
        out1 => S1572
    );
nand_n_736: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1572,
        in1(1) => S1571,
        out1 => S1543
    );
nand_n_737: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1553,
        in1(1) => CU_inst_9,
        out1 => S1573
    );
nand_n_738: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1555,
        in1(1) => dataBus(9),
        out1 => S1574
    );
nand_n_739: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1574,
        in1(1) => S1573,
        out1 => S1544
    );
nand_n_740: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1553,
        in1(1) => CU_inst_10,
        out1 => S1575
    );
nand_n_741: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1555,
        in1(1) => dataBus(10),
        out1 => S1576
    );
nand_n_742: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1576,
        in1(1) => S1575,
        out1 => S1545
    );
nand_n_743: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1553,
        in1(1) => CU_inst_11,
        out1 => S1577
    );
nand_n_744: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1555,
        in1(1) => dataBus(11),
        out1 => S1578
    );
nand_n_745: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1578,
        in1(1) => S1577,
        out1 => S1546
    );
nand_n_746: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1553,
        in1(1) => CU_inst_12,
        out1 => S1579
    );
nand_n_747: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1555,
        in1(1) => dataBus(12),
        out1 => S1580
    );
nand_n_748: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1580,
        in1(1) => S1579,
        out1 => S1547
    );
nand_n_749: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1553,
        in1(1) => CU_inst_13,
        out1 => S1581
    );
nand_n_750: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1555,
        in1(1) => dataBus(13),
        out1 => S1582
    );
nand_n_751: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1582,
        in1(1) => S1581,
        out1 => S1548
    );
nand_n_752: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1553,
        in1(1) => CU_inst_14,
        out1 => S1583
    );
nand_n_753: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1555,
        in1(1) => dataBus(14),
        out1 => S1584
    );
nand_n_754: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1584,
        in1(1) => S1583,
        out1 => S1549
    );
nand_n_755: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1553,
        in1(1) => CU_inst_15,
        out1 => S1585
    );
nand_n_756: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1555,
        in1(1) => dataBus(15),
        out1 => S1551
    );
nand_n_757: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1551,
        in1(1) => S1585,
        out1 => S1550
    );
dff_35: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S1535,
        NbarT => '0',
        PRE => '0',
        Q => CU_inst_0,
        Si => S3337,
        global_reset => '0'
    );
dff_36: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S1536,
        NbarT => '0',
        PRE => '0',
        Q => CU_inst_1,
        Si => S3336,
        global_reset => '0'
    );
dff_37: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S1537,
        NbarT => '0',
        PRE => '0',
        Q => CU_inst_2,
        Si => S3335,
        global_reset => '0'
    );
dff_38: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S1538,
        NbarT => '0',
        PRE => '0',
        Q => CU_inst_3,
        Si => S3334,
        global_reset => '0'
    );
dff_39: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S1539,
        NbarT => '0',
        PRE => '0',
        Q => CU_inst_4,
        Si => S3333,
        global_reset => '0'
    );
dff_40: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S1540,
        NbarT => '0',
        PRE => '0',
        Q => CU_inst_5,
        Si => S3332,
        global_reset => '0'
    );
dff_41: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S1541,
        NbarT => '0',
        PRE => '0',
        Q => CU_inst_6,
        Si => S3331,
        global_reset => '0'
    );
dff_42: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S1542,
        NbarT => '0',
        PRE => '0',
        Q => CU_inst_7,
        Si => S3330,
        global_reset => '0'
    );
dff_43: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S1543,
        NbarT => '0',
        PRE => '0',
        Q => CU_inst_8,
        Si => S3329,
        global_reset => '0'
    );
dff_44: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S1544,
        NbarT => '0',
        PRE => '0',
        Q => CU_inst_9,
        Si => S3328,
        global_reset => '0'
    );
dff_45: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S1545,
        NbarT => '0',
        PRE => '0',
        Q => CU_inst_10,
        Si => S3327,
        global_reset => '0'
    );
dff_46: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S1546,
        NbarT => '0',
        PRE => '0',
        Q => CU_inst_11,
        Si => S3326,
        global_reset => '0'
    );
dff_47: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S1547,
        NbarT => '0',
        PRE => '0',
        Q => CU_inst_12,
        Si => S3325,
        global_reset => '0'
    );
dff_48: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S1548,
        NbarT => '0',
        PRE => '0',
        Q => CU_inst_13,
        Si => S3324,
        global_reset => '0'
    );
dff_49: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S1549,
        NbarT => '0',
        PRE => '0',
        Q => CU_inst_14,
        Si => S3323,
        global_reset => '0'
    );
dff_50: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S1550,
        NbarT => '0',
        PRE => '0',
        Q => CU_inst_15,
        Si => S3358,
        global_reset => '0'
    );
notg_252: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_AC_out_15,
        out1 => S1652
    );
notg_253: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_LGU1_in1_0,
        out1 => S1653
    );
notg_254: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_LGU1_in1_1,
        out1 => S1654
    );
notg_255: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_AC_out_4,
        out1 => S1655
    );
notg_256: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_AC_out_5,
        out1 => S1656
    );
notg_257: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_LGU1_in1_2,
        out1 => S1657
    );
notg_258: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_LGU1_in1_3,
        out1 => S1658
    );
notg_259: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_LGU1_in1_4,
        out1 => S1659
    );
notg_260: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_SHF_0,
        out1 => S1660
    );
notg_261: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_SHF_1,
        out1 => S1661
    );
notg_262: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_NOT,
        out1 => S1662
    );
nor_n_622: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => DP_LGU1_out_7,
        in1(1) => DP_LGU1_out_4,
        out1 => S1663
    );
nor_n_623: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => DP_LGU1_out_2,
        in1(1) => DP_LGU1_out_1,
        out1 => S1664
    );
nand_n_758: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1664,
        in1(1) => S1663,
        out1 => S1665
    );
nor_n_624: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => DP_LGU1_out_14,
        in1(1) => DP_LGU1_out_13,
        out1 => S1666
    );
nor_n_625: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => DP_LGU1_out_11,
        in1(1) => DP_LGU1_out_8,
        out1 => S1667
    );
nand_n_759: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1667,
        in1(1) => S1666,
        out1 => S1668
    );
nor_n_626: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1668,
        in1(1) => S1665,
        out1 => S1669
    );
nor_n_627: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => DP_LGU1_out_6,
        in1(1) => DP_LGU1_out_5,
        out1 => S1670
    );
nor_n_628: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => DP_LGU1_out_3,
        in1(1) => DP_LGU1_out_0,
        out1 => S1671
    );
nand_n_760: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1671,
        in1(1) => S1670,
        out1 => S1672
    );
nor_n_629: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => DP_LGU1_N,
        in1(1) => DP_LGU1_out_12,
        out1 => S1673
    );
nor_n_630: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => DP_LGU1_out_10,
        in1(1) => DP_LGU1_out_9,
        out1 => S1674
    );
nand_n_761: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1674,
        in1(1) => S1673,
        out1 => S1675
    );
nor_n_631: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1675,
        in1(1) => S1672,
        out1 => S1676
    );
nand_n_762: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1676,
        in1(1) => S1669,
        out1 => S1677
    );
notg_263: ENTITY WORK.notg
    PORT MAP (
        in1 => S1677,
        out1 => DP_LGU1_Z
    );
nor_n_632: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => DP_LGU1_in1_15,
        in1(1) => DP_LGU1_in1_14,
        out1 => S1678
    );
notg_264: ENTITY WORK.notg
    PORT MAP (
        in1 => S1678,
        out1 => S1679
    );
nor_n_633: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1679,
        in1(1) => DP_LGU1_in1_13,
        out1 => S1680
    );
nor_n_634: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => DP_LGU1_in1_9,
        in1(1) => DP_LGU1_in1_10,
        out1 => S1681
    );
nor_n_635: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => DP_LGU1_in1_11,
        in1(1) => DP_LGU1_in1_12,
        out1 => S1682
    );
nand_n_763: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1682,
        in1(1) => S1681,
        out1 => S1683
    );
nor_n_636: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => DP_LGU1_in1_5,
        in1(1) => DP_LGU1_in1_6,
        out1 => S1684
    );
nor_n_637: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => DP_LGU1_in1_7,
        in1(1) => DP_LGU1_in1_8,
        out1 => S1685
    );
nand_n_764: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1685,
        in1(1) => S1684,
        out1 => S1686
    );
notg_265: ENTITY WORK.notg
    PORT MAP (
        in1 => S1686,
        out1 => S1687
    );
nor_n_638: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1686,
        in1(1) => S1683,
        out1 => S1688
    );
nand_n_765: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1687,
        in1(1) => S1680,
        out1 => S1689
    );
nor_n_639: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1689,
        in1(1) => S1683,
        out1 => S1690
    );
nand_n_766: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1688,
        in1(1) => S1680,
        out1 => S1691
    );
nor_n_640: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1691,
        in1(1) => S1655,
        out1 => S1692
    );
nand_n_767: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1690,
        in1(1) => DP_AC_out_4,
        out1 => S1693
    );
nor_n_641: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1693,
        in1(1) => DP_LGU1_in1_0,
        out1 => S1694
    );
nand_n_768: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1692,
        in1(1) => S1653,
        out1 => S1695
    );
nor_n_642: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1691,
        in1(1) => S1656,
        out1 => S1696
    );
nand_n_769: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1690,
        in1(1) => DP_AC_out_5,
        out1 => S1697
    );
nor_n_643: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1697,
        in1(1) => S1653,
        out1 => S1698
    );
nand_n_770: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1696,
        in1(1) => DP_LGU1_in1_0,
        out1 => S1699
    );
nand_n_771: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1699,
        in1(1) => S1695,
        out1 => S1700
    );
nor_n_644: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1700,
        in1(1) => DP_LGU1_in1_1,
        out1 => S1701
    );
notg_266: ENTITY WORK.notg
    PORT MAP (
        in1 => S1701,
        out1 => S1702
    );
nand_n_772: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1690,
        in1(1) => DP_AC_out_6,
        out1 => S1703
    );
nor_n_645: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1703,
        in1(1) => DP_LGU1_in1_0,
        out1 => S1704
    );
nand_n_773: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1690,
        in1(1) => DP_AC_out_7,
        out1 => S1705
    );
nand_n_774: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1703,
        in1(1) => S1653,
        out1 => S1706
    );
nand_n_775: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1705,
        in1(1) => DP_LGU1_in1_0,
        out1 => S1707
    );
nand_n_776: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1707,
        in1(1) => S1706,
        out1 => S1708
    );
notg_267: ENTITY WORK.notg
    PORT MAP (
        in1 => S1708,
        out1 => S1709
    );
nand_n_777: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1708,
        in1(1) => DP_LGU1_in1_1,
        out1 => S1710
    );
notg_268: ENTITY WORK.notg
    PORT MAP (
        in1 => S1710,
        out1 => S1711
    );
nor_n_646: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1711,
        in1(1) => S1701,
        out1 => S1712
    );
nand_n_778: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1710,
        in1(1) => S1702,
        out1 => S1713
    );
nand_n_779: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1712,
        in1(1) => DP_LGU1_in1_2,
        out1 => S1714
    );
nand_n_780: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1690,
        in1(1) => DP_AC_out_2,
        out1 => S1715
    );
nor_n_647: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1715,
        in1(1) => DP_LGU1_in1_0,
        out1 => S1716
    );
nand_n_781: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1690,
        in1(1) => DP_AC_out_3,
        out1 => S1717
    );
nor_n_648: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1717,
        in1(1) => S1653,
        out1 => S1718
    );
nor_n_649: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1718,
        in1(1) => S1716,
        out1 => S1719
    );
notg_269: ENTITY WORK.notg
    PORT MAP (
        in1 => S1719,
        out1 => S1720
    );
nor_n_650: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1719,
        in1(1) => S1654,
        out1 => S1721
    );
nand_n_782: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1690,
        in1(1) => DP_AC_out_1,
        out1 => S1722
    );
notg_270: ENTITY WORK.notg
    PORT MAP (
        in1 => S1722,
        out1 => S1723
    );
nor_n_651: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1722,
        in1(1) => S1653,
        out1 => S1724
    );
nand_n_783: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1723,
        in1(1) => DP_LGU1_in1_0,
        out1 => S1725
    );
nor_n_652: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1725,
        in1(1) => DP_LGU1_in1_1,
        out1 => S1726
    );
nor_n_653: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1726,
        in1(1) => S1721,
        out1 => S1727
    );
nor_n_654: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1727,
        in1(1) => DP_LGU1_in1_2,
        out1 => S1728
    );
nand_n_784: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1690,
        in1(1) => DP_AC_out_0,
        out1 => S1729
    );
nor_n_655: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1729,
        in1(1) => DP_LGU1_in1_0,
        out1 => S1730
    );
nand_n_785: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1730,
        in1(1) => S1654,
        out1 => S1731
    );
nor_n_656: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1731,
        in1(1) => DP_LGU1_in1_2,
        out1 => S1732
    );
nor_n_657: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1732,
        in1(1) => DP_LGU1_in1_3,
        out1 => S1733
    );
notg_271: ENTITY WORK.notg
    PORT MAP (
        in1 => S1733,
        out1 => S1734
    );
nor_n_658: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1734,
        in1(1) => S1728,
        out1 => S1735
    );
nand_n_786: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1733,
        in1(1) => S1714,
        out1 => S1736
    );
nor_n_659: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1736,
        in1(1) => S1728,
        out1 => S1737
    );
nand_n_787: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1735,
        in1(1) => S1714,
        out1 => S1738
    );
nand_n_788: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1690,
        in1(1) => DP_AC_out_8,
        out1 => S1739
    );
nand_n_789: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1739,
        in1(1) => S1653,
        out1 => S1740
    );
nand_n_790: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1690,
        in1(1) => DP_AC_out_9,
        out1 => S1741
    );
nand_n_791: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1741,
        in1(1) => DP_LGU1_in1_0,
        out1 => S1742
    );
nand_n_792: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1742,
        in1(1) => S1740,
        out1 => S1743
    );
nand_n_793: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1743,
        in1(1) => S1654,
        out1 => S1744
    );
nand_n_794: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1690,
        in1(1) => DP_AC_out_10,
        out1 => S1745
    );
nand_n_795: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1745,
        in1(1) => S1653,
        out1 => S1746
    );
nand_n_796: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1690,
        in1(1) => DP_AC_out_11,
        out1 => S1747
    );
nand_n_797: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1747,
        in1(1) => DP_LGU1_in1_0,
        out1 => S1748
    );
nand_n_798: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1748,
        in1(1) => S1746,
        out1 => S1749
    );
notg_272: ENTITY WORK.notg
    PORT MAP (
        in1 => S1749,
        out1 => S1750
    );
nand_n_799: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1749,
        in1(1) => DP_LGU1_in1_1,
        out1 => S1751
    );
nand_n_800: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1751,
        in1(1) => S1744,
        out1 => S1752
    );
nand_n_801: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1752,
        in1(1) => S1657,
        out1 => S1753
    );
nand_n_802: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1690,
        in1(1) => DP_AC_out_12,
        out1 => S1754
    );
nand_n_803: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1754,
        in1(1) => S1653,
        out1 => S1755
    );
nand_n_804: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1690,
        in1(1) => DP_AC_out_13,
        out1 => S1756
    );
nand_n_805: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1756,
        in1(1) => DP_LGU1_in1_0,
        out1 => S1757
    );
nand_n_806: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1757,
        in1(1) => S1755,
        out1 => S1758
    );
nand_n_807: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1758,
        in1(1) => S1654,
        out1 => S1759
    );
nand_n_808: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1690,
        in1(1) => DP_AC_out_14,
        out1 => S1760
    );
nand_n_809: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1760,
        in1(1) => S1653,
        out1 => S1761
    );
nand_n_810: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1690,
        in1(1) => DP_AC_out_15,
        out1 => S1762
    );
nand_n_811: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1762,
        in1(1) => DP_LGU1_in1_0,
        out1 => S1763
    );
nand_n_812: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1763,
        in1(1) => S1761,
        out1 => S1764
    );
nand_n_813: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1764,
        in1(1) => DP_LGU1_in1_1,
        out1 => S1765
    );
nand_n_814: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1765,
        in1(1) => S1759,
        out1 => S1766
    );
nand_n_815: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1766,
        in1(1) => DP_LGU1_in1_2,
        out1 => S1767
    );
nand_n_816: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1767,
        in1(1) => S1753,
        out1 => S1768
    );
nand_n_817: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1768,
        in1(1) => DP_LGU1_in1_3,
        out1 => S1769
    );
nand_n_818: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1769,
        in1(1) => S1738,
        out1 => S1603
    );
nor_n_660: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => CU_SHF_1,
        in1(1) => S1660,
        out1 => S1604
    );
nand_n_819: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1732,
        in1(1) => S1658,
        out1 => S1605
    );
nand_n_820: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_0,
        in1(1) => CU_AND,
        out1 => S1770
    );
notg_273: ENTITY WORK.notg
    PORT MAP (
        in1 => S1770,
        out1 => S1771
    );
nand_n_821: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1771,
        in1(1) => DP_LGU1_in1_0,
        out1 => S1772
    );
nor_n_661: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => CU_NOT,
        in1(1) => CU_AND,
        out1 => S1773
    );
nand_n_822: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_NOT,
        in1(1) => DP_AC_out_0,
        out1 => S1774
    );
notg_274: ENTITY WORK.notg
    PORT MAP (
        in1 => S1774,
        out1 => S1775
    );
nor_n_662: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1775,
        in1(1) => CU_AND,
        out1 => S1776
    );
nor_n_663: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => CU_SHF_1,
        in1(1) => CU_SHF_0,
        out1 => S1777
    );
nand_n_823: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1661,
        in1(1) => S1660,
        out1 => S1778
    );
nand_n_824: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_in1_0,
        in1(1) => S1652,
        out1 => S1779
    );
nand_n_825: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1779,
        in1(1) => S1761,
        out1 => S1780
    );
nand_n_826: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1780,
        in1(1) => DP_LGU1_in1_1,
        out1 => S1781
    );
nand_n_827: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1781,
        in1(1) => S1759,
        out1 => S1782
    );
nand_n_828: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1782,
        in1(1) => DP_LGU1_in1_2,
        out1 => S1783
    );
nand_n_829: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1783,
        in1(1) => S1753,
        out1 => S1784
    );
nand_n_830: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1784,
        in1(1) => DP_LGU1_in1_3,
        out1 => S1785
    );
nor_n_664: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1737,
        in1(1) => DP_LGU1_in1_4,
        out1 => S1786
    );
nand_n_831: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1786,
        in1(1) => S1785,
        out1 => S1787
    );
nor_n_665: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1659,
        in1(1) => S1652,
        out1 => S1788
    );
nand_n_832: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_in1_4,
        in1(1) => DP_AC_out_15,
        out1 => S1789
    );
nor_n_666: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1690,
        in1(1) => S1652,
        out1 => S1790
    );
nand_n_833: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1691,
        in1(1) => DP_AC_out_15,
        out1 => S1791
    );
nor_n_667: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1790,
        in1(1) => S1788,
        out1 => S1792
    );
nand_n_834: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1792,
        in1(1) => S1787,
        out1 => S1793
    );
nand_n_835: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1793,
        in1(1) => S1777,
        out1 => S1794
    );
nand_n_836: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1778,
        in1(1) => S1659,
        out1 => S1795
    );
nor_n_668: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1795,
        in1(1) => S1636,
        out1 => S1796
    );
nor_n_669: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1796,
        in1(1) => CU_NOT,
        out1 => S1797
    );
nand_n_837: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1797,
        in1(1) => S1794,
        out1 => S1798
    );
nand_n_838: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1798,
        in1(1) => S1776,
        out1 => S1799
    );
nand_n_839: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1799,
        in1(1) => S1772,
        out1 => S1586
    );
nand_n_840: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1722,
        in1(1) => S1653,
        out1 => S1800
    );
nand_n_841: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1715,
        in1(1) => DP_LGU1_in1_0,
        out1 => S1801
    );
nand_n_842: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1801,
        in1(1) => S1800,
        out1 => S1802
    );
nand_n_843: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1802,
        in1(1) => S1654,
        out1 => S1803
    );
nand_n_844: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1717,
        in1(1) => S1653,
        out1 => S1804
    );
nand_n_845: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1693,
        in1(1) => DP_LGU1_in1_0,
        out1 => S1805
    );
nand_n_846: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1805,
        in1(1) => S1804,
        out1 => S1806
    );
nand_n_847: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1806,
        in1(1) => DP_LGU1_in1_1,
        out1 => S1807
    );
nand_n_848: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1807,
        in1(1) => S1803,
        out1 => S1808
    );
nand_n_849: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1808,
        in1(1) => S1657,
        out1 => S1809
    );
nand_n_850: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1697,
        in1(1) => S1653,
        out1 => S1810
    );
nand_n_851: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1703,
        in1(1) => DP_LGU1_in1_0,
        out1 => S1811
    );
nand_n_852: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1811,
        in1(1) => S1810,
        out1 => S1812
    );
nand_n_853: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1812,
        in1(1) => S1654,
        out1 => S1813
    );
nand_n_854: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1705,
        in1(1) => S1653,
        out1 => S1814
    );
nand_n_855: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1739,
        in1(1) => DP_LGU1_in1_0,
        out1 => S1815
    );
nand_n_856: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1815,
        in1(1) => S1814,
        out1 => S1816
    );
nand_n_857: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1816,
        in1(1) => DP_LGU1_in1_1,
        out1 => S1817
    );
nand_n_858: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1817,
        in1(1) => S1813,
        out1 => S1818
    );
nand_n_859: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1818,
        in1(1) => DP_LGU1_in1_2,
        out1 => S1819
    );
nand_n_860: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1819,
        in1(1) => S1809,
        out1 => S1820
    );
nand_n_861: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1820,
        in1(1) => S1658,
        out1 => S1821
    );
nor_n_670: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1745,
        in1(1) => S1653,
        out1 => S1822
    );
nand_n_862: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1741,
        in1(1) => S1653,
        out1 => S1823
    );
nand_n_863: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1745,
        in1(1) => DP_LGU1_in1_0,
        out1 => S1824
    );
nand_n_864: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1824,
        in1(1) => S1823,
        out1 => S1825
    );
notg_275: ENTITY WORK.notg
    PORT MAP (
        in1 => S1825,
        out1 => S1826
    );
nor_n_671: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1826,
        in1(1) => DP_LGU1_in1_1,
        out1 => S1827
    );
nand_n_865: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1825,
        in1(1) => S1654,
        out1 => S1828
    );
nor_n_672: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1754,
        in1(1) => S1653,
        out1 => S1829
    );
nor_n_673: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1747,
        in1(1) => DP_LGU1_in1_0,
        out1 => S1830
    );
nor_n_674: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1830,
        in1(1) => S1829,
        out1 => S1831
    );
nand_n_866: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1831,
        in1(1) => DP_LGU1_in1_1,
        out1 => S1832
    );
notg_276: ENTITY WORK.notg
    PORT MAP (
        in1 => S1832,
        out1 => S1833
    );
nor_n_675: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1833,
        in1(1) => S1827,
        out1 => S1834
    );
nand_n_867: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1832,
        in1(1) => S1828,
        out1 => S1835
    );
nor_n_676: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1834,
        in1(1) => DP_LGU1_in1_2,
        out1 => S1836
    );
nand_n_868: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1835,
        in1(1) => S1657,
        out1 => S1837
    );
nor_n_677: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1760,
        in1(1) => S1653,
        out1 => S1838
    );
nor_n_678: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1756,
        in1(1) => DP_LGU1_in1_0,
        out1 => S1839
    );
nor_n_679: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1839,
        in1(1) => S1838,
        out1 => S1840
    );
nor_n_680: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1840,
        in1(1) => DP_LGU1_in1_1,
        out1 => S1841
    );
nor_n_681: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1762,
        in1(1) => DP_LGU1_in1_0,
        out1 => S1842
    );
nand_n_869: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1842,
        in1(1) => DP_LGU1_in1_1,
        out1 => S1843
    );
notg_277: ENTITY WORK.notg
    PORT MAP (
        in1 => S1843,
        out1 => S1844
    );
nor_n_682: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1844,
        in1(1) => S1841,
        out1 => S1845
    );
nand_n_870: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1845,
        in1(1) => DP_LGU1_in1_2,
        out1 => S1846
    );
nand_n_871: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1846,
        in1(1) => S1837,
        out1 => S1847
    );
nand_n_872: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1847,
        in1(1) => DP_LGU1_in1_3,
        out1 => S1848
    );
nand_n_873: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1848,
        in1(1) => S1821,
        out1 => S1606
    );
nand_n_874: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1729,
        in1(1) => DP_LGU1_in1_0,
        out1 => S1849
    );
nand_n_875: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1849,
        in1(1) => S1800,
        out1 => S1850
    );
notg_278: ENTITY WORK.notg
    PORT MAP (
        in1 => S1850,
        out1 => S1851
    );
nand_n_876: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1851,
        in1(1) => S1654,
        out1 => S1852
    );
nor_n_683: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1852,
        in1(1) => DP_LGU1_in1_2,
        out1 => S1853
    );
notg_279: ENTITY WORK.notg
    PORT MAP (
        in1 => S1853,
        out1 => S1854
    );
nand_n_877: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1853,
        in1(1) => S1658,
        out1 => S1607
    );
nand_n_878: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_1,
        in1(1) => CU_AND,
        out1 => S1855
    );
notg_280: ENTITY WORK.notg
    PORT MAP (
        in1 => S1855,
        out1 => S1856
    );
nand_n_879: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1856,
        in1(1) => DP_LGU1_in1_1,
        out1 => S1857
    );
nor_n_684: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1637,
        in1(1) => DP_LGU1_in1_4,
        out1 => S1858
    );
nor_n_685: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1858,
        in1(1) => S1777,
        out1 => S1859
    );
notg_281: ENTITY WORK.notg
    PORT MAP (
        in1 => S1859,
        out1 => S1860
    );
nor_n_686: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1788,
        in1(1) => S1778,
        out1 => S1861
    );
nand_n_880: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1789,
        in1(1) => S1777,
        out1 => S1862
    );
nor_n_687: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1821,
        in1(1) => S1790,
        out1 => S1863
    );
nor_n_688: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1837,
        in1(1) => S1790,
        out1 => S1864
    );
nand_n_881: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1836,
        in1(1) => S1791,
        out1 => S1865
    );
nor_n_689: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1691,
        in1(1) => DP_LGU1_in1_1,
        out1 => S1866
    );
nor_n_690: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1866,
        in1(1) => S1652,
        out1 => S1867
    );
nor_n_691: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1867,
        in1(1) => S1841,
        out1 => S1868
    );
nand_n_882: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1868,
        in1(1) => DP_LGU1_in1_2,
        out1 => S1869
    );
notg_282: ENTITY WORK.notg
    PORT MAP (
        in1 => S1869,
        out1 => S1870
    );
nor_n_692: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1870,
        in1(1) => S1864,
        out1 => S1871
    );
nand_n_883: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1869,
        in1(1) => S1865,
        out1 => S1872
    );
nor_n_693: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1871,
        in1(1) => S1658,
        out1 => S1873
    );
nor_n_694: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1873,
        in1(1) => S1863,
        out1 => S1874
    );
nand_n_884: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1874,
        in1(1) => S1659,
        out1 => S1875
    );
nand_n_885: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1875,
        in1(1) => S1861,
        out1 => S1876
    );
nand_n_886: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1876,
        in1(1) => S1860,
        out1 => S1877
    );
nand_n_887: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1877,
        in1(1) => S1662,
        out1 => S1878
    );
nand_n_888: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_NOT,
        in1(1) => DP_AC_out_1,
        out1 => S1879
    );
notg_283: ENTITY WORK.notg
    PORT MAP (
        in1 => S1879,
        out1 => S1880
    );
nor_n_695: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1880,
        in1(1) => CU_AND,
        out1 => S1881
    );
nand_n_889: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1881,
        in1(1) => S1878,
        out1 => S1882
    );
nand_n_890: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1882,
        in1(1) => S1857,
        out1 => S1593
    );
nor_n_696: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1700,
        in1(1) => S1654,
        out1 => S1883
    );
nor_n_697: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1720,
        in1(1) => DP_LGU1_in1_1,
        out1 => S1884
    );
nor_n_698: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1884,
        in1(1) => S1883,
        out1 => S1885
    );
nor_n_699: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1885,
        in1(1) => DP_LGU1_in1_2,
        out1 => S1886
    );
nor_n_700: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1709,
        in1(1) => DP_LGU1_in1_1,
        out1 => S1887
    );
nand_n_891: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1708,
        in1(1) => S1654,
        out1 => S1888
    );
nand_n_892: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1743,
        in1(1) => DP_LGU1_in1_1,
        out1 => S1889
    );
notg_284: ENTITY WORK.notg
    PORT MAP (
        in1 => S1889,
        out1 => S1890
    );
nor_n_701: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1890,
        in1(1) => S1887,
        out1 => S1891
    );
nand_n_893: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1889,
        in1(1) => S1888,
        out1 => S1892
    );
nor_n_702: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1891,
        in1(1) => S1657,
        out1 => S1893
    );
nor_n_703: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1893,
        in1(1) => S1886,
        out1 => S1894
    );
nand_n_894: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1891,
        in1(1) => DP_LGU1_in1_2,
        out1 => S1895
    );
nor_n_704: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1884,
        in1(1) => DP_LGU1_in1_2,
        out1 => S1896
    );
notg_285: ENTITY WORK.notg
    PORT MAP (
        in1 => S1896,
        out1 => S1897
    );
nor_n_705: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1897,
        in1(1) => S1883,
        out1 => S1898
    );
nor_n_706: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1898,
        in1(1) => DP_LGU1_in1_3,
        out1 => S1899
    );
nor_n_707: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1894,
        in1(1) => DP_LGU1_in1_3,
        out1 => S1900
    );
nand_n_895: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1899,
        in1(1) => S1895,
        out1 => S1901
    );
nor_n_708: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1750,
        in1(1) => DP_LGU1_in1_1,
        out1 => S1902
    );
nand_n_896: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1749,
        in1(1) => S1654,
        out1 => S1903
    );
nand_n_897: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1758,
        in1(1) => DP_LGU1_in1_1,
        out1 => S1904
    );
notg_286: ENTITY WORK.notg
    PORT MAP (
        in1 => S1904,
        out1 => S1905
    );
nor_n_709: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1905,
        in1(1) => S1902,
        out1 => S1906
    );
nand_n_898: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1904,
        in1(1) => S1903,
        out1 => S1907
    );
nor_n_710: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1906,
        in1(1) => DP_LGU1_in1_2,
        out1 => S1908
    );
nand_n_899: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1907,
        in1(1) => S1657,
        out1 => S1909
    );
nor_n_711: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1764,
        in1(1) => DP_LGU1_in1_1,
        out1 => S1910
    );
notg_287: ENTITY WORK.notg
    PORT MAP (
        in1 => S1910,
        out1 => S1911
    );
nor_n_712: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1910,
        in1(1) => S1657,
        out1 => S1912
    );
nor_n_713: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1912,
        in1(1) => S1908,
        out1 => S1913
    );
notg_288: ENTITY WORK.notg
    PORT MAP (
        in1 => S1913,
        out1 => S1914
    );
nand_n_900: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1914,
        in1(1) => DP_LGU1_in1_3,
        out1 => S1915
    );
nand_n_901: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1915,
        in1(1) => S1901,
        out1 => S1608
    );
nor_n_714: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1724,
        in1(1) => S1716,
        out1 => S1916
    );
nor_n_715: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1916,
        in1(1) => DP_LGU1_in1_1,
        out1 => S1917
    );
nand_n_902: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1730,
        in1(1) => DP_LGU1_in1_1,
        out1 => S1918
    );
notg_289: ENTITY WORK.notg
    PORT MAP (
        in1 => S1918,
        out1 => S1919
    );
nor_n_716: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1919,
        in1(1) => S1917,
        out1 => S1920
    );
nor_n_717: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1920,
        in1(1) => DP_LGU1_in1_2,
        out1 => S1921
    );
notg_290: ENTITY WORK.notg
    PORT MAP (
        in1 => S1921,
        out1 => S1922
    );
nand_n_903: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1921,
        in1(1) => S1658,
        out1 => S1609
    );
nand_n_904: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_2,
        in1(1) => CU_AND,
        out1 => S1923
    );
notg_291: ENTITY WORK.notg
    PORT MAP (
        in1 => S1923,
        out1 => S1924
    );
nand_n_905: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1924,
        in1(1) => DP_LGU1_in1_2,
        out1 => S1925
    );
nor_n_718: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1638,
        in1(1) => DP_LGU1_in1_4,
        out1 => S1926
    );
nor_n_719: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1926,
        in1(1) => S1777,
        out1 => S1927
    );
notg_292: ENTITY WORK.notg
    PORT MAP (
        in1 => S1927,
        out1 => S1928
    );
nand_n_906: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1900,
        in1(1) => S1791,
        out1 => S1929
    );
nor_n_720: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1909,
        in1(1) => S1790,
        out1 => S1930
    );
nand_n_907: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1908,
        in1(1) => S1791,
        out1 => S1931
    );
nor_n_721: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1780,
        in1(1) => DP_LGU1_in1_1,
        out1 => S1932
    );
nor_n_722: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1932,
        in1(1) => S1867,
        out1 => S1933
    );
nand_n_908: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1933,
        in1(1) => DP_LGU1_in1_2,
        out1 => S1934
    );
notg_293: ENTITY WORK.notg
    PORT MAP (
        in1 => S1934,
        out1 => S1935
    );
nor_n_723: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1935,
        in1(1) => S1930,
        out1 => S1936
    );
nand_n_909: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1934,
        in1(1) => S1931,
        out1 => S1937
    );
nor_n_724: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1936,
        in1(1) => S1658,
        out1 => S1938
    );
nor_n_725: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1938,
        in1(1) => DP_LGU1_in1_4,
        out1 => S1939
    );
nand_n_910: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1939,
        in1(1) => S1929,
        out1 => S1940
    );
nand_n_911: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1940,
        in1(1) => S1861,
        out1 => S1941
    );
nand_n_912: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1941,
        in1(1) => S1928,
        out1 => S1942
    );
nand_n_913: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1942,
        in1(1) => S1662,
        out1 => S1943
    );
nand_n_914: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_NOT,
        in1(1) => DP_AC_out_2,
        out1 => S1944
    );
notg_294: ENTITY WORK.notg
    PORT MAP (
        in1 => S1944,
        out1 => S1945
    );
nor_n_726: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1945,
        in1(1) => CU_AND,
        out1 => S1946
    );
nand_n_915: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1946,
        in1(1) => S1943,
        out1 => S1947
    );
nand_n_916: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1947,
        in1(1) => S1925,
        out1 => S1594
    );
nand_n_917: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1806,
        in1(1) => S1654,
        out1 => S1948
    );
nand_n_918: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1812,
        in1(1) => DP_LGU1_in1_1,
        out1 => S1949
    );
nand_n_919: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1949,
        in1(1) => S1948,
        out1 => S1950
    );
nand_n_920: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1950,
        in1(1) => S1657,
        out1 => S1951
    );
nand_n_921: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1816,
        in1(1) => S1654,
        out1 => S1952
    );
nand_n_922: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1825,
        in1(1) => DP_LGU1_in1_1,
        out1 => S1953
    );
nand_n_923: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1953,
        in1(1) => S1952,
        out1 => S1954
    );
nand_n_924: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1954,
        in1(1) => DP_LGU1_in1_2,
        out1 => S1955
    );
nand_n_925: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1955,
        in1(1) => S1951,
        out1 => S1956
    );
nand_n_926: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1956,
        in1(1) => S1658,
        out1 => S1957
    );
nand_n_927: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1842,
        in1(1) => S1654,
        out1 => S1958
    );
nor_n_727: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1958,
        in1(1) => S1657,
        out1 => S1959
    );
nand_n_928: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1831,
        in1(1) => S1654,
        out1 => S1960
    );
nand_n_929: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1840,
        in1(1) => DP_LGU1_in1_1,
        out1 => S1961
    );
nand_n_930: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1961,
        in1(1) => S1960,
        out1 => S1962
    );
nor_n_728: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1962,
        in1(1) => DP_LGU1_in1_2,
        out1 => S1963
    );
nor_n_729: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1963,
        in1(1) => S1959,
        out1 => S1964
    );
nand_n_931: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1964,
        in1(1) => DP_LGU1_in1_3,
        out1 => S1965
    );
nand_n_932: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1965,
        in1(1) => S1957,
        out1 => S1610
    );
nand_n_933: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1804,
        in1(1) => S1801,
        out1 => S1966
    );
nand_n_934: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1966,
        in1(1) => S1654,
        out1 => S1967
    );
nand_n_935: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1850,
        in1(1) => DP_LGU1_in1_1,
        out1 => S1968
    );
nand_n_936: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1968,
        in1(1) => S1967,
        out1 => S1969
    );
nor_n_730: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1969,
        in1(1) => DP_LGU1_in1_2,
        out1 => S1970
    );
notg_295: ENTITY WORK.notg
    PORT MAP (
        in1 => S1970,
        out1 => S1971
    );
nand_n_937: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1970,
        in1(1) => S1658,
        out1 => S1611
    );
nand_n_938: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_3,
        in1(1) => CU_AND,
        out1 => S1972
    );
notg_296: ENTITY WORK.notg
    PORT MAP (
        in1 => S1972,
        out1 => S1973
    );
nand_n_939: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1973,
        in1(1) => DP_LGU1_in1_3,
        out1 => S1974
    );
nor_n_731: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1639,
        in1(1) => DP_LGU1_in1_4,
        out1 => S1975
    );
nor_n_732: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1975,
        in1(1) => S1777,
        out1 => S1976
    );
nor_n_733: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1957,
        in1(1) => S1790,
        out1 => S1977
    );
nand_n_940: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_in1_2,
        in1(1) => DP_AC_out_15,
        out1 => S1978
    );
notg_297: ENTITY WORK.notg
    PORT MAP (
        in1 => S1978,
        out1 => S1979
    );
nand_n_941: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1978,
        in1(1) => S1791,
        out1 => S1980
    );
nor_n_734: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1980,
        in1(1) => S1963,
        out1 => S1981
    );
nand_n_942: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1981,
        in1(1) => DP_LGU1_in1_3,
        out1 => S1982
    );
nand_n_943: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1982,
        in1(1) => S1659,
        out1 => S1983
    );
nor_n_735: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1983,
        in1(1) => S1977,
        out1 => S1984
    );
nor_n_736: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1984,
        in1(1) => S1862,
        out1 => S1985
    );
nor_n_737: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1985,
        in1(1) => S1976,
        out1 => S1986
    );
nor_n_738: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1986,
        in1(1) => CU_NOT,
        out1 => S1987
    );
notg_298: ENTITY WORK.notg
    PORT MAP (
        in1 => S1987,
        out1 => S1988
    );
nand_n_944: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_NOT,
        in1(1) => DP_AC_out_3,
        out1 => S1989
    );
notg_299: ENTITY WORK.notg
    PORT MAP (
        in1 => S1989,
        out1 => S1990
    );
nor_n_739: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1990,
        in1(1) => CU_AND,
        out1 => S1991
    );
nand_n_945: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1991,
        in1(1) => S1988,
        out1 => S1992
    );
nand_n_946: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1992,
        in1(1) => S1974,
        out1 => S1595
    );
nand_n_947: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1713,
        in1(1) => S1657,
        out1 => S1993
    );
nand_n_948: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1752,
        in1(1) => DP_LGU1_in1_2,
        out1 => S1994
    );
nand_n_949: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1994,
        in1(1) => S1993,
        out1 => S1995
    );
nand_n_950: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1995,
        in1(1) => S1658,
        out1 => S1996
    );
nor_n_740: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1766,
        in1(1) => DP_LGU1_in1_2,
        out1 => S1997
    );
notg_300: ENTITY WORK.notg
    PORT MAP (
        in1 => S1997,
        out1 => S1998
    );
nand_n_951: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1998,
        in1(1) => DP_LGU1_in1_3,
        out1 => S1999
    );
nand_n_952: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1999,
        in1(1) => S1996,
        out1 => S1612
    );
nor_n_741: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1718,
        in1(1) => S1694,
        out1 => S2000
    );
nand_n_953: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2000,
        in1(1) => S1654,
        out1 => S2001
    );
nand_n_954: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1916,
        in1(1) => DP_LGU1_in1_1,
        out1 => S2002
    );
nand_n_955: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2002,
        in1(1) => S2001,
        out1 => S2003
    );
nand_n_956: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2003,
        in1(1) => S1657,
        out1 => S2004
    );
nand_n_957: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1731,
        in1(1) => DP_LGU1_in1_2,
        out1 => S2005
    );
nand_n_958: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2005,
        in1(1) => S2004,
        out1 => S2006
    );
nor_n_742: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2006,
        in1(1) => DP_LGU1_in1_3,
        out1 => S2007
    );
notg_301: ENTITY WORK.notg
    PORT MAP (
        in1 => S2007,
        out1 => S1613
    );
nor_n_743: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1659,
        in1(1) => S1655,
        out1 => S2008
    );
nand_n_959: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2008,
        in1(1) => CU_AND,
        out1 => S2009
    );
nor_n_744: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1640,
        in1(1) => DP_LGU1_in1_4,
        out1 => S2010
    );
nor_n_745: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2010,
        in1(1) => S1777,
        out1 => S2011
    );
nor_n_746: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1996,
        in1(1) => S1790,
        out1 => S2012
    );
nor_n_747: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1782,
        in1(1) => DP_LGU1_in1_2,
        out1 => S2013
    );
nor_n_748: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2013,
        in1(1) => S1980,
        out1 => S2014
    );
nand_n_960: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2014,
        in1(1) => DP_LGU1_in1_3,
        out1 => S2015
    );
nand_n_961: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2015,
        in1(1) => S1659,
        out1 => S2016
    );
nor_n_749: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2016,
        in1(1) => S2012,
        out1 => S2017
    );
nor_n_750: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2017,
        in1(1) => S1862,
        out1 => S2018
    );
nor_n_751: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2018,
        in1(1) => S2011,
        out1 => S2019
    );
nor_n_752: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2019,
        in1(1) => CU_NOT,
        out1 => S2020
    );
notg_302: ENTITY WORK.notg
    PORT MAP (
        in1 => S2020,
        out1 => S2021
    );
nand_n_962: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_NOT,
        in1(1) => DP_AC_out_4,
        out1 => S2022
    );
notg_303: ENTITY WORK.notg
    PORT MAP (
        in1 => S2022,
        out1 => S2023
    );
nor_n_753: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2023,
        in1(1) => CU_AND,
        out1 => S2024
    );
nand_n_963: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2024,
        in1(1) => S2021,
        out1 => S2025
    );
nand_n_964: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2025,
        in1(1) => S2009,
        out1 => S1596
    );
nor_n_754: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1818,
        in1(1) => DP_LGU1_in1_2,
        out1 => S2026
    );
nor_n_755: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2026,
        in1(1) => DP_LGU1_in1_3,
        out1 => S2027
    );
nand_n_965: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1834,
        in1(1) => DP_LGU1_in1_2,
        out1 => S2028
    );
nand_n_966: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2028,
        in1(1) => S2027,
        out1 => S2029
    );
nor_n_756: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1845,
        in1(1) => DP_LGU1_in1_2,
        out1 => S2030
    );
notg_304: ENTITY WORK.notg
    PORT MAP (
        in1 => S2030,
        out1 => S2031
    );
nand_n_967: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2031,
        in1(1) => DP_LGU1_in1_3,
        out1 => S2032
    );
nand_n_968: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2032,
        in1(1) => S2029,
        out1 => S1614
    );
nand_n_969: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1810,
        in1(1) => S1805,
        out1 => S2033
    );
nand_n_970: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2033,
        in1(1) => S1654,
        out1 => S2034
    );
nand_n_971: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1966,
        in1(1) => DP_LGU1_in1_1,
        out1 => S2035
    );
nand_n_972: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2035,
        in1(1) => S2034,
        out1 => S2036
    );
nand_n_973: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2036,
        in1(1) => S1657,
        out1 => S2037
    );
nand_n_974: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1852,
        in1(1) => DP_LGU1_in1_2,
        out1 => S2038
    );
nand_n_975: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2038,
        in1(1) => S2037,
        out1 => S2039
    );
nor_n_757: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2039,
        in1(1) => DP_LGU1_in1_3,
        out1 => S2040
    );
notg_305: ENTITY WORK.notg
    PORT MAP (
        in1 => S2040,
        out1 => S1615
    );
nand_n_976: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_in1_5,
        in1(1) => CU_AND,
        out1 => S2041
    );
notg_306: ENTITY WORK.notg
    PORT MAP (
        in1 => S2041,
        out1 => S2042
    );
nand_n_977: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2042,
        in1(1) => DP_AC_out_5,
        out1 => S2043
    );
nor_n_758: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1641,
        in1(1) => DP_LGU1_in1_4,
        out1 => S2044
    );
nor_n_759: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2044,
        in1(1) => S1777,
        out1 => S2045
    );
notg_307: ENTITY WORK.notg
    PORT MAP (
        in1 => S2045,
        out1 => S2046
    );
nor_n_760: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2029,
        in1(1) => S1790,
        out1 => S2047
    );
nor_n_761: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1868,
        in1(1) => DP_LGU1_in1_2,
        out1 => S2048
    );
notg_308: ENTITY WORK.notg
    PORT MAP (
        in1 => S2048,
        out1 => S2049
    );
nor_n_762: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2048,
        in1(1) => S1979,
        out1 => S2050
    );
nand_n_978: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2049,
        in1(1) => S1978,
        out1 => S2051
    );
nor_n_763: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2051,
        in1(1) => S1658,
        out1 => S2052
    );
nor_n_764: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2052,
        in1(1) => S2047,
        out1 => S2053
    );
nand_n_979: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2053,
        in1(1) => S1659,
        out1 => S2054
    );
nand_n_980: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2054,
        in1(1) => S1861,
        out1 => S2055
    );
nand_n_981: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2055,
        in1(1) => S2046,
        out1 => S2056
    );
nand_n_982: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2056,
        in1(1) => S1662,
        out1 => S2057
    );
nand_n_983: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_NOT,
        in1(1) => DP_AC_out_5,
        out1 => S2058
    );
notg_309: ENTITY WORK.notg
    PORT MAP (
        in1 => S2058,
        out1 => S2059
    );
nor_n_765: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2059,
        in1(1) => CU_AND,
        out1 => S2060
    );
nand_n_984: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2060,
        in1(1) => S2057,
        out1 => S2061
    );
nand_n_985: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2061,
        in1(1) => S2043,
        out1 => S1597
    );
nor_n_766: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1892,
        in1(1) => DP_LGU1_in1_2,
        out1 => S2062
    );
nor_n_767: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2062,
        in1(1) => DP_LGU1_in1_3,
        out1 => S2063
    );
nand_n_986: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1906,
        in1(1) => DP_LGU1_in1_2,
        out1 => S2064
    );
nand_n_987: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2064,
        in1(1) => S2063,
        out1 => S2065
    );
nor_n_768: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1911,
        in1(1) => DP_LGU1_in1_2,
        out1 => S2066
    );
nand_n_988: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1910,
        in1(1) => S1657,
        out1 => S2067
    );
nand_n_989: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2067,
        in1(1) => DP_LGU1_in1_3,
        out1 => S2068
    );
nand_n_990: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2068,
        in1(1) => S2065,
        out1 => S1616
    );
nor_n_769: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1704,
        in1(1) => S1698,
        out1 => S2069
    );
nand_n_991: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2069,
        in1(1) => S1654,
        out1 => S2070
    );
nand_n_992: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2000,
        in1(1) => DP_LGU1_in1_1,
        out1 => S2071
    );
nand_n_993: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2071,
        in1(1) => S2070,
        out1 => S2072
    );
nand_n_994: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2072,
        in1(1) => S1657,
        out1 => S2073
    );
nand_n_995: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1920,
        in1(1) => DP_LGU1_in1_2,
        out1 => S2074
    );
nand_n_996: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2074,
        in1(1) => S2073,
        out1 => S2075
    );
nor_n_770: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2075,
        in1(1) => DP_LGU1_in1_3,
        out1 => S2076
    );
notg_310: ENTITY WORK.notg
    PORT MAP (
        in1 => S2076,
        out1 => S1617
    );
nand_n_997: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_in1_6,
        in1(1) => CU_AND,
        out1 => S2077
    );
notg_311: ENTITY WORK.notg
    PORT MAP (
        in1 => S2077,
        out1 => S2078
    );
nand_n_998: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2078,
        in1(1) => DP_AC_out_6,
        out1 => S2079
    );
nor_n_771: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1642,
        in1(1) => DP_LGU1_in1_4,
        out1 => S2080
    );
nor_n_772: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2080,
        in1(1) => S1777,
        out1 => S2081
    );
notg_312: ENTITY WORK.notg
    PORT MAP (
        in1 => S2081,
        out1 => S2082
    );
nor_n_773: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2065,
        in1(1) => S1790,
        out1 => S2083
    );
nor_n_774: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1933,
        in1(1) => DP_LGU1_in1_2,
        out1 => S2084
    );
notg_313: ENTITY WORK.notg
    PORT MAP (
        in1 => S2084,
        out1 => S2085
    );
nor_n_775: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2084,
        in1(1) => S1979,
        out1 => S2086
    );
nand_n_999: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2085,
        in1(1) => S1978,
        out1 => S2087
    );
nor_n_776: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2087,
        in1(1) => S1658,
        out1 => S2088
    );
nor_n_777: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2088,
        in1(1) => S2083,
        out1 => S2089
    );
nand_n_1000: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2089,
        in1(1) => S1659,
        out1 => S2090
    );
nand_n_1001: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2090,
        in1(1) => S1861,
        out1 => S2091
    );
nand_n_1002: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2091,
        in1(1) => S2082,
        out1 => S2092
    );
nand_n_1003: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2092,
        in1(1) => S1662,
        out1 => S2093
    );
nand_n_1004: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_NOT,
        in1(1) => DP_AC_out_6,
        out1 => S2094
    );
notg_314: ENTITY WORK.notg
    PORT MAP (
        in1 => S2094,
        out1 => S2095
    );
nor_n_778: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2095,
        in1(1) => CU_AND,
        out1 => S2096
    );
nand_n_1005: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2096,
        in1(1) => S2093,
        out1 => S2097
    );
nand_n_1006: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2097,
        in1(1) => S2079,
        out1 => S1598
    );
nor_n_779: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1962,
        in1(1) => S1657,
        out1 => S2098
    );
nor_n_780: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1954,
        in1(1) => DP_LGU1_in1_2,
        out1 => S2099
    );
nor_n_781: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2099,
        in1(1) => S2098,
        out1 => S2100
    );
nor_n_782: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2100,
        in1(1) => DP_LGU1_in1_3,
        out1 => S2101
    );
notg_315: ENTITY WORK.notg
    PORT MAP (
        in1 => S2101,
        out1 => S2102
    );
nor_n_783: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1958,
        in1(1) => DP_LGU1_in1_2,
        out1 => S2103
    );
nand_n_1007: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2103,
        in1(1) => DP_LGU1_in1_3,
        out1 => S2104
    );
notg_316: ENTITY WORK.notg
    PORT MAP (
        in1 => S2104,
        out1 => S2105
    );
nor_n_784: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2105,
        in1(1) => S2101,
        out1 => S1618
    );
nand_n_1008: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1814,
        in1(1) => S1811,
        out1 => S2106
    );
nand_n_1009: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2106,
        in1(1) => S1654,
        out1 => S2107
    );
nand_n_1010: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2033,
        in1(1) => DP_LGU1_in1_1,
        out1 => S2108
    );
nand_n_1011: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2108,
        in1(1) => S2107,
        out1 => S2109
    );
nand_n_1012: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2109,
        in1(1) => S1657,
        out1 => S2110
    );
nand_n_1013: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1969,
        in1(1) => DP_LGU1_in1_2,
        out1 => S2111
    );
nand_n_1014: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2111,
        in1(1) => S2110,
        out1 => S2112
    );
nor_n_785: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2112,
        in1(1) => DP_LGU1_in1_3,
        out1 => S2113
    );
notg_317: ENTITY WORK.notg
    PORT MAP (
        in1 => S2113,
        out1 => S1619
    );
nor_n_786: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1643,
        in1(1) => DP_LGU1_in1_4,
        out1 => S2114
    );
nor_n_787: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2114,
        in1(1) => S1777,
        out1 => S2115
    );
nor_n_788: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => DP_LGU1_in1_4,
        in1(1) => DP_LGU1_in1_3,
        out1 => S2116
    );
notg_318: ENTITY WORK.notg
    PORT MAP (
        in1 => S2116,
        out1 => S2117
    );
nor_n_789: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2116,
        in1(1) => S1652,
        out1 => S2118
    );
nor_n_790: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2118,
        in1(1) => S1778,
        out1 => S2119
    );
nand_n_1015: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2119,
        in1(1) => S1791,
        out1 => S2120
    );
nor_n_791: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2102,
        in1(1) => DP_LGU1_in1_4,
        out1 => S2121
    );
nor_n_792: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2121,
        in1(1) => S2120,
        out1 => S2122
    );
nor_n_793: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2122,
        in1(1) => S2115,
        out1 => S2123
    );
nor_n_794: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2123,
        in1(1) => CU_NOT,
        out1 => S2124
    );
notg_319: ENTITY WORK.notg
    PORT MAP (
        in1 => S2124,
        out1 => S2125
    );
nand_n_1016: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_NOT,
        in1(1) => DP_AC_out_7,
        out1 => S2126
    );
notg_320: ENTITY WORK.notg
    PORT MAP (
        in1 => S2126,
        out1 => S2127
    );
nor_n_795: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2127,
        in1(1) => CU_AND,
        out1 => S2128
    );
nand_n_1017: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2128,
        in1(1) => S2125,
        out1 => S2129
    );
nand_n_1018: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_in1_7,
        in1(1) => CU_AND,
        out1 => S2130
    );
notg_321: ENTITY WORK.notg
    PORT MAP (
        in1 => S2130,
        out1 => S2131
    );
nand_n_1019: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2131,
        in1(1) => DP_AC_out_7,
        out1 => S2132
    );
nand_n_1020: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2132,
        in1(1) => S2129,
        out1 => S1599
    );
nor_n_796: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1768,
        in1(1) => DP_LGU1_in1_3,
        out1 => S2133
    );
notg_322: ENTITY WORK.notg
    PORT MAP (
        in1 => S2133,
        out1 => S1620
    );
nor_n_797: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2003,
        in1(1) => S1657,
        out1 => S2134
    );
nand_n_1021: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1740,
        in1(1) => S1707,
        out1 => S2135
    );
nand_n_1022: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2135,
        in1(1) => S1654,
        out1 => S2136
    );
nand_n_1023: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2069,
        in1(1) => DP_LGU1_in1_1,
        out1 => S2137
    );
nand_n_1024: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2137,
        in1(1) => S2136,
        out1 => S2138
    );
nor_n_798: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2138,
        in1(1) => DP_LGU1_in1_2,
        out1 => S2139
    );
nor_n_799: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2139,
        in1(1) => S2134,
        out1 => S2140
    );
nor_n_800: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2140,
        in1(1) => DP_LGU1_in1_3,
        out1 => S2141
    );
nand_n_1025: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1732,
        in1(1) => DP_LGU1_in1_3,
        out1 => S2142
    );
notg_323: ENTITY WORK.notg
    PORT MAP (
        in1 => S2142,
        out1 => S2143
    );
nor_n_801: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2143,
        in1(1) => S2141,
        out1 => S1621
    );
nor_n_802: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1644,
        in1(1) => DP_LGU1_in1_4,
        out1 => S2144
    );
nor_n_803: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2144,
        in1(1) => S1777,
        out1 => S2145
    );
nor_n_804: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2117,
        in1(1) => S1784,
        out1 => S2146
    );
nor_n_805: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2146,
        in1(1) => S2120,
        out1 => S2147
    );
nor_n_806: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2147,
        in1(1) => S2145,
        out1 => S2148
    );
nor_n_807: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2148,
        in1(1) => CU_NOT,
        out1 => S2149
    );
notg_324: ENTITY WORK.notg
    PORT MAP (
        in1 => S2149,
        out1 => S2150
    );
nand_n_1026: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_NOT,
        in1(1) => DP_AC_out_8,
        out1 => S2151
    );
notg_325: ENTITY WORK.notg
    PORT MAP (
        in1 => S2151,
        out1 => S2152
    );
nor_n_808: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2152,
        in1(1) => CU_AND,
        out1 => S2153
    );
nand_n_1027: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2153,
        in1(1) => S2150,
        out1 => S2154
    );
nand_n_1028: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_in1_8,
        in1(1) => CU_AND,
        out1 => S2155
    );
notg_326: ENTITY WORK.notg
    PORT MAP (
        in1 => S2155,
        out1 => S2156
    );
nand_n_1029: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2156,
        in1(1) => DP_AC_out_8,
        out1 => S2157
    );
nand_n_1030: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2157,
        in1(1) => S2154,
        out1 => S1600
    );
nor_n_809: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1847,
        in1(1) => DP_LGU1_in1_3,
        out1 => S2158
    );
notg_327: ENTITY WORK.notg
    PORT MAP (
        in1 => S2158,
        out1 => S1622
    );
nand_n_1031: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1823,
        in1(1) => S1815,
        out1 => S2159
    );
nand_n_1032: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2159,
        in1(1) => S1654,
        out1 => S2160
    );
nand_n_1033: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2106,
        in1(1) => DP_LGU1_in1_1,
        out1 => S2161
    );
nand_n_1034: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2161,
        in1(1) => S2160,
        out1 => S2162
    );
nand_n_1035: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2162,
        in1(1) => S1657,
        out1 => S2163
    );
nand_n_1036: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2036,
        in1(1) => DP_LGU1_in1_2,
        out1 => S2164
    );
nand_n_1037: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2164,
        in1(1) => S2163,
        out1 => S2165
    );
nand_n_1038: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2165,
        in1(1) => S1658,
        out1 => S2166
    );
nand_n_1039: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1854,
        in1(1) => DP_LGU1_in1_3,
        out1 => S2167
    );
nand_n_1040: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2167,
        in1(1) => S2166,
        out1 => S1623
    );
nand_n_1041: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_NOT,
        in1(1) => DP_AC_out_9,
        out1 => S2168
    );
notg_328: ENTITY WORK.notg
    PORT MAP (
        in1 => S2168,
        out1 => S2169
    );
nor_n_810: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2169,
        in1(1) => CU_AND,
        out1 => S2170
    );
nand_n_1042: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2116,
        in1(1) => S1872,
        out1 => S2171
    );
nand_n_1043: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1777,
        in1(1) => DP_AC_out_15,
        out1 => S2172
    );
nor_n_811: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2116,
        in1(1) => DP_AC_out_15,
        out1 => S2173
    );
nor_n_812: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2173,
        in1(1) => S1778,
        out1 => S2174
    );
nand_n_1044: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2174,
        in1(1) => S2171,
        out1 => S2175
    );
nor_n_813: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1795,
        in1(1) => S1645,
        out1 => S2176
    );
nor_n_814: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2176,
        in1(1) => CU_NOT,
        out1 => S2177
    );
nand_n_1045: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2177,
        in1(1) => S2175,
        out1 => S2178
    );
nand_n_1046: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2178,
        in1(1) => S2170,
        out1 => S2179
    );
nand_n_1047: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_in1_9,
        in1(1) => CU_AND,
        out1 => S2180
    );
notg_329: ENTITY WORK.notg
    PORT MAP (
        in1 => S2180,
        out1 => S2181
    );
nand_n_1048: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2181,
        in1(1) => DP_AC_out_9,
        out1 => S2182
    );
nand_n_1049: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2182,
        in1(1) => S2179,
        out1 => S1601
    );
nand_n_1050: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1913,
        in1(1) => S1658,
        out1 => S1624
    );
nand_n_1051: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1746,
        in1(1) => S1742,
        out1 => S2183
    );
nand_n_1052: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2183,
        in1(1) => S1654,
        out1 => S2184
    );
nand_n_1053: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2135,
        in1(1) => DP_LGU1_in1_1,
        out1 => S2185
    );
nand_n_1054: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2185,
        in1(1) => S2184,
        out1 => S2186
    );
nand_n_1055: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2186,
        in1(1) => S1657,
        out1 => S2187
    );
nand_n_1056: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2072,
        in1(1) => DP_LGU1_in1_2,
        out1 => S2188
    );
nand_n_1057: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2188,
        in1(1) => S2187,
        out1 => S2189
    );
nand_n_1058: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2189,
        in1(1) => S1658,
        out1 => S2190
    );
nand_n_1059: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1922,
        in1(1) => DP_LGU1_in1_3,
        out1 => S2191
    );
nand_n_1060: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2191,
        in1(1) => S2190,
        out1 => S1625
    );
nand_n_1061: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_NOT,
        in1(1) => DP_AC_out_10,
        out1 => S2192
    );
notg_330: ENTITY WORK.notg
    PORT MAP (
        in1 => S2192,
        out1 => S2193
    );
nor_n_815: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2193,
        in1(1) => CU_AND,
        out1 => S2194
    );
nand_n_1062: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2116,
        in1(1) => S1937,
        out1 => S2195
    );
nand_n_1063: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2195,
        in1(1) => S2174,
        out1 => S2196
    );
nor_n_816: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1795,
        in1(1) => S1646,
        out1 => S2197
    );
nor_n_817: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2197,
        in1(1) => CU_NOT,
        out1 => S2198
    );
nand_n_1064: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2198,
        in1(1) => S2196,
        out1 => S2199
    );
nand_n_1065: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2199,
        in1(1) => S2194,
        out1 => S2200
    );
nand_n_1066: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_in1_10,
        in1(1) => CU_AND,
        out1 => S2201
    );
notg_331: ENTITY WORK.notg
    PORT MAP (
        in1 => S2201,
        out1 => S2202
    );
nand_n_1067: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2202,
        in1(1) => DP_AC_out_10,
        out1 => S2203
    );
nand_n_1068: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2203,
        in1(1) => S2200,
        out1 => S1587
    );
nor_n_818: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1964,
        in1(1) => DP_LGU1_in1_3,
        out1 => S2204
    );
notg_332: ENTITY WORK.notg
    PORT MAP (
        in1 => S2204,
        out1 => S1626
    );
nor_n_819: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1830,
        in1(1) => S1822,
        out1 => S2205
    );
nand_n_1069: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2205,
        in1(1) => S1654,
        out1 => S2206
    );
nand_n_1070: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2159,
        in1(1) => DP_LGU1_in1_1,
        out1 => S2207
    );
nand_n_1071: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2207,
        in1(1) => S2206,
        out1 => S2208
    );
nand_n_1072: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2208,
        in1(1) => S1657,
        out1 => S2209
    );
nand_n_1073: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2109,
        in1(1) => DP_LGU1_in1_2,
        out1 => S2210
    );
nand_n_1074: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2210,
        in1(1) => S2209,
        out1 => S2211
    );
nand_n_1075: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2211,
        in1(1) => S1658,
        out1 => S2212
    );
nand_n_1076: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1971,
        in1(1) => DP_LGU1_in1_3,
        out1 => S2213
    );
nand_n_1077: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2213,
        in1(1) => S2212,
        out1 => S1627
    );
nand_n_1078: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_NOT,
        in1(1) => DP_AC_out_11,
        out1 => S2214
    );
notg_333: ENTITY WORK.notg
    PORT MAP (
        in1 => S2214,
        out1 => S2215
    );
nor_n_820: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2215,
        in1(1) => CU_AND,
        out1 => S2216
    );
nand_n_1079: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2116,
        in1(1) => S1981,
        out1 => S2217
    );
nand_n_1080: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2217,
        in1(1) => S2174,
        out1 => S2218
    );
nor_n_821: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1795,
        in1(1) => S1647,
        out1 => S2219
    );
nor_n_822: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2219,
        in1(1) => CU_NOT,
        out1 => S2220
    );
nand_n_1081: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2220,
        in1(1) => S2218,
        out1 => S2221
    );
nand_n_1082: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2221,
        in1(1) => S2216,
        out1 => S2222
    );
nand_n_1083: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_in1_11,
        in1(1) => CU_AND,
        out1 => S2223
    );
notg_334: ENTITY WORK.notg
    PORT MAP (
        in1 => S2223,
        out1 => S2224
    );
nand_n_1084: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2224,
        in1(1) => DP_AC_out_11,
        out1 => S2225
    );
nand_n_1085: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2225,
        in1(1) => S2222,
        out1 => S1588
    );
nand_n_1086: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1997,
        in1(1) => S1658,
        out1 => S1628
    );
nand_n_1087: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1755,
        in1(1) => S1748,
        out1 => S2226
    );
nand_n_1088: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2226,
        in1(1) => S1654,
        out1 => S2227
    );
nand_n_1089: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2183,
        in1(1) => DP_LGU1_in1_1,
        out1 => S2228
    );
nand_n_1090: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2228,
        in1(1) => S2227,
        out1 => S2229
    );
nand_n_1091: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2229,
        in1(1) => S1657,
        out1 => S2230
    );
nand_n_1092: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2138,
        in1(1) => DP_LGU1_in1_2,
        out1 => S2231
    );
nand_n_1093: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2231,
        in1(1) => S2230,
        out1 => S2232
    );
nand_n_1094: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2232,
        in1(1) => S1658,
        out1 => S2233
    );
nand_n_1095: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2006,
        in1(1) => DP_LGU1_in1_3,
        out1 => S2234
    );
nand_n_1096: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2234,
        in1(1) => S2233,
        out1 => S1629
    );
nand_n_1097: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_NOT,
        in1(1) => DP_AC_out_12,
        out1 => S2235
    );
notg_335: ENTITY WORK.notg
    PORT MAP (
        in1 => S2235,
        out1 => S2236
    );
nor_n_823: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2236,
        in1(1) => CU_AND,
        out1 => S2237
    );
nand_n_1098: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2116,
        in1(1) => S2014,
        out1 => S2238
    );
nand_n_1099: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2238,
        in1(1) => S2174,
        out1 => S2239
    );
nor_n_824: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1795,
        in1(1) => S1648,
        out1 => S2240
    );
nor_n_825: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2240,
        in1(1) => CU_NOT,
        out1 => S2241
    );
nand_n_1100: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2241,
        in1(1) => S2239,
        out1 => S2242
    );
nand_n_1101: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2242,
        in1(1) => S2237,
        out1 => S2243
    );
nand_n_1102: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_in1_12,
        in1(1) => CU_AND,
        out1 => S2244
    );
notg_336: ENTITY WORK.notg
    PORT MAP (
        in1 => S2244,
        out1 => S2245
    );
nand_n_1103: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2245,
        in1(1) => DP_AC_out_12,
        out1 => S2246
    );
nand_n_1104: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2246,
        in1(1) => S2243,
        out1 => S1589
    );
nand_n_1105: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2030,
        in1(1) => S1658,
        out1 => S1630
    );
nor_n_826: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1839,
        in1(1) => S1829,
        out1 => S2247
    );
nand_n_1106: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2247,
        in1(1) => S1654,
        out1 => S2248
    );
nand_n_1107: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2205,
        in1(1) => DP_LGU1_in1_1,
        out1 => S2249
    );
nand_n_1108: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2249,
        in1(1) => S2248,
        out1 => S2250
    );
nand_n_1109: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2250,
        in1(1) => S1657,
        out1 => S2251
    );
nand_n_1110: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2162,
        in1(1) => DP_LGU1_in1_2,
        out1 => S2252
    );
nand_n_1111: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2252,
        in1(1) => S2251,
        out1 => S2253
    );
nand_n_1112: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2253,
        in1(1) => S1658,
        out1 => S2254
    );
nand_n_1113: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2039,
        in1(1) => DP_LGU1_in1_3,
        out1 => S2255
    );
nand_n_1114: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2255,
        in1(1) => S2254,
        out1 => S1631
    );
nand_n_1115: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_NOT,
        in1(1) => DP_AC_out_13,
        out1 => S2256
    );
notg_337: ENTITY WORK.notg
    PORT MAP (
        in1 => S2256,
        out1 => S2257
    );
nor_n_827: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2257,
        in1(1) => CU_AND,
        out1 => S2258
    );
nand_n_1116: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2116,
        in1(1) => S2050,
        out1 => S2259
    );
nand_n_1117: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2259,
        in1(1) => S2174,
        out1 => S2260
    );
nor_n_828: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1795,
        in1(1) => S1649,
        out1 => S2261
    );
nor_n_829: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2261,
        in1(1) => CU_NOT,
        out1 => S2262
    );
nand_n_1118: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2262,
        in1(1) => S2260,
        out1 => S2263
    );
nand_n_1119: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2263,
        in1(1) => S2258,
        out1 => S2264
    );
nand_n_1120: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_in1_13,
        in1(1) => CU_AND,
        out1 => S2265
    );
notg_338: ENTITY WORK.notg
    PORT MAP (
        in1 => S2265,
        out1 => S2266
    );
nand_n_1121: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2266,
        in1(1) => DP_AC_out_13,
        out1 => S2267
    );
nand_n_1122: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2267,
        in1(1) => S2264,
        out1 => S1590
    );
nand_n_1123: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2066,
        in1(1) => S1658,
        out1 => S1632
    );
nand_n_1124: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1761,
        in1(1) => S1757,
        out1 => S2268
    );
nand_n_1125: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2268,
        in1(1) => S1654,
        out1 => S2269
    );
nand_n_1126: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2226,
        in1(1) => DP_LGU1_in1_1,
        out1 => S2270
    );
nand_n_1127: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2270,
        in1(1) => S2269,
        out1 => S2271
    );
nand_n_1128: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2271,
        in1(1) => S1657,
        out1 => S2272
    );
nand_n_1129: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2186,
        in1(1) => DP_LGU1_in1_2,
        out1 => S2273
    );
nand_n_1130: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2273,
        in1(1) => S2272,
        out1 => S2274
    );
nand_n_1131: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2274,
        in1(1) => S1658,
        out1 => S2275
    );
nand_n_1132: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2075,
        in1(1) => DP_LGU1_in1_3,
        out1 => S2276
    );
nand_n_1133: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2276,
        in1(1) => S2275,
        out1 => S1633
    );
nand_n_1134: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_NOT,
        in1(1) => DP_AC_out_14,
        out1 => S2277
    );
notg_339: ENTITY WORK.notg
    PORT MAP (
        in1 => S2277,
        out1 => S2278
    );
nor_n_830: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2278,
        in1(1) => CU_AND,
        out1 => S2279
    );
nand_n_1135: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2116,
        in1(1) => S2086,
        out1 => S2280
    );
nand_n_1136: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2280,
        in1(1) => S2174,
        out1 => S2281
    );
nor_n_831: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1795,
        in1(1) => S1650,
        out1 => S2282
    );
nor_n_832: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2282,
        in1(1) => CU_NOT,
        out1 => S2283
    );
nand_n_1137: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2283,
        in1(1) => S2281,
        out1 => S2284
    );
nand_n_1138: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2284,
        in1(1) => S2279,
        out1 => S2285
    );
nand_n_1139: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_in1_14,
        in1(1) => CU_AND,
        out1 => S2286
    );
notg_340: ENTITY WORK.notg
    PORT MAP (
        in1 => S2286,
        out1 => S2287
    );
nand_n_1140: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2287,
        in1(1) => DP_AC_out_14,
        out1 => S2288
    );
nand_n_1141: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2288,
        in1(1) => S2285,
        out1 => S1591
    );
nand_n_1142: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2103,
        in1(1) => S1658,
        out1 => S1634
    );
nor_n_833: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2112,
        in1(1) => S1658,
        out1 => S2289
    );
nor_n_834: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2247,
        in1(1) => S1654,
        out1 => S2290
    );
nand_n_1143: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1838,
        in1(1) => S1654,
        out1 => S2291
    );
nand_n_1144: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2291,
        in1(1) => S1958,
        out1 => S2292
    );
nor_n_835: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2292,
        in1(1) => S2290,
        out1 => S2293
    );
nor_n_836: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2293,
        in1(1) => DP_LGU1_in1_2,
        out1 => S2294
    );
nor_n_837: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2208,
        in1(1) => S1657,
        out1 => S2295
    );
nor_n_838: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2295,
        in1(1) => S2294,
        out1 => S2296
    );
nor_n_839: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2296,
        in1(1) => DP_LGU1_in1_3,
        out1 => S2297
    );
nor_n_840: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2297,
        in1(1) => S2289,
        out1 => S1635
    );
nand_n_1145: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_15,
        in1(1) => DP_LGU1_in1_15,
        out1 => S2298
    );
nand_n_1146: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2298,
        in1(1) => CU_AND,
        out1 => S2299
    );
notg_341: ENTITY WORK.notg
    PORT MAP (
        in1 => S2299,
        out1 => S2300
    );
nor_n_841: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1795,
        in1(1) => S1651,
        out1 => S2301
    );
nand_n_1147: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2172,
        in1(1) => S1662,
        out1 => S2302
    );
nor_n_842: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2302,
        in1(1) => S2301,
        out1 => S2303
    );
nand_n_1148: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_NOT,
        in1(1) => DP_AC_out_15,
        out1 => S2304
    );
notg_342: ENTITY WORK.notg
    PORT MAP (
        in1 => S2304,
        out1 => S2305
    );
nor_n_843: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2305,
        in1(1) => S2303,
        out1 => S2306
    );
nor_n_844: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2306,
        in1(1) => CU_AND,
        out1 => S2307
    );
nor_n_845: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2307,
        in1(1) => S2300,
        out1 => S1592
    );
nand_n_1149: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1773,
        in1(1) => CU_SHF_0,
        out1 => S2308
    );
nor_n_846: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2308,
        in1(1) => S1661,
        out1 => S1602
    );
$mux_1: ENTITY WORK.$mux
    PORT MAP (
        A => S1605,
        B => S1603,
        S => S1604,
        Y => S1636
    );
$mux_2: ENTITY WORK.$mux
    PORT MAP (
        A => S1607,
        B => S1606,
        S => S1604,
        Y => S1637
    );
$mux_3: ENTITY WORK.$mux
    PORT MAP (
        A => S1609,
        B => S1608,
        S => S1604,
        Y => S1638
    );
$mux_4: ENTITY WORK.$mux
    PORT MAP (
        A => S1611,
        B => S1610,
        S => S1604,
        Y => S1639
    );
$mux_5: ENTITY WORK.$mux
    PORT MAP (
        A => S1613,
        B => S1612,
        S => S1604,
        Y => S1640
    );
$mux_6: ENTITY WORK.$mux
    PORT MAP (
        A => S1615,
        B => S1614,
        S => S1604,
        Y => S1641
    );
$mux_7: ENTITY WORK.$mux
    PORT MAP (
        A => S1617,
        B => S1616,
        S => S1604,
        Y => S1642
    );
$mux_8: ENTITY WORK.$mux
    PORT MAP (
        A => S1619,
        B => S1618,
        S => S1604,
        Y => S1643
    );
$mux_9: ENTITY WORK.$mux
    PORT MAP (
        A => S1621,
        B => S1620,
        S => S1604,
        Y => S1644
    );
$mux_10: ENTITY WORK.$mux
    PORT MAP (
        A => S1623,
        B => S1622,
        S => S1604,
        Y => S1645
    );
$mux_11: ENTITY WORK.$mux
    PORT MAP (
        A => S1625,
        B => S1624,
        S => S1604,
        Y => S1646
    );
$mux_12: ENTITY WORK.$mux
    PORT MAP (
        A => S1627,
        B => S1626,
        S => S1604,
        Y => S1647
    );
$mux_13: ENTITY WORK.$mux
    PORT MAP (
        A => S1629,
        B => S1628,
        S => S1604,
        Y => S1648
    );
$mux_14: ENTITY WORK.$mux
    PORT MAP (
        A => S1631,
        B => S1630,
        S => S1604,
        Y => S1649
    );
$mux_15: ENTITY WORK.$mux
    PORT MAP (
        A => S1633,
        B => S1632,
        S => S1604,
        Y => S1650
    );
$mux_16: ENTITY WORK.$mux
    PORT MAP (
        A => S1635,
        B => S1634,
        S => S1604,
        Y => S1651
    );
$_DLATCH_N__35: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S1586,
        E => S1602,
        Q => DP_LGU1_out_0
    );
$_DLATCH_N__36: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S1593,
        E => S1602,
        Q => DP_LGU1_out_1
    );
$_DLATCH_N__37: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S1594,
        E => S1602,
        Q => DP_LGU1_out_2
    );
$_DLATCH_N__38: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S1595,
        E => S1602,
        Q => DP_LGU1_out_3
    );
$_DLATCH_N__39: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S1596,
        E => S1602,
        Q => DP_LGU1_out_4
    );
$_DLATCH_N__40: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S1597,
        E => S1602,
        Q => DP_LGU1_out_5
    );
$_DLATCH_N__41: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S1598,
        E => S1602,
        Q => DP_LGU1_out_6
    );
$_DLATCH_N__42: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S1599,
        E => S1602,
        Q => DP_LGU1_out_7
    );
$_DLATCH_N__43: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S1600,
        E => S1602,
        Q => DP_LGU1_out_8
    );
$_DLATCH_N__44: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S1601,
        E => S1602,
        Q => DP_LGU1_out_9
    );
$_DLATCH_N__45: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S1587,
        E => S1602,
        Q => DP_LGU1_out_10
    );
$_DLATCH_N__46: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S1588,
        E => S1602,
        Q => DP_LGU1_out_11
    );
$_DLATCH_N__47: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S1589,
        E => S1602,
        Q => DP_LGU1_out_12
    );
$_DLATCH_N__48: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S1590,
        E => S1602,
        Q => DP_LGU1_out_13
    );
$_DLATCH_N__49: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S1591,
        E => S1602,
        Q => DP_LGU1_out_14
    );
$_DLATCH_N__50: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S1592,
        E => S1602,
        Q => DP_LGU1_N
    );
notg_343: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_ldOF,
        out1 => S2313
    );
nor_n_847: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => CU_ldOF,
        in1(1) => S13,
        out1 => S2314
    );
nand_n_1150: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2314,
        in1(1) => DP_IMM1_in1_0,
        out1 => S2315
    );
nor_n_848: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2313,
        in1(1) => S14,
        out1 => S2316
    );
nand_n_1151: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2316,
        in1(1) => DP_OF_in_0,
        out1 => S2317
    );
nand_n_1152: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2317,
        in1(1) => S2315,
        out1 => S2309
    );
nand_n_1153: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2314,
        in1(1) => DP_IMM1_in1_1,
        out1 => S2318
    );
nand_n_1154: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2316,
        in1(1) => DP_OF_in_1,
        out1 => S2319
    );
nand_n_1155: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2319,
        in1(1) => S2318,
        out1 => S2310
    );
nand_n_1156: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2314,
        in1(1) => DP_IMM1_in1_2,
        out1 => S2320
    );
nand_n_1157: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2316,
        in1(1) => DP_OF_in_2,
        out1 => S2321
    );
nand_n_1158: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2321,
        in1(1) => S2320,
        out1 => S2311
    );
nand_n_1159: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2314,
        in1(1) => DP_IMM1_in1_3,
        out1 => S2322
    );
nand_n_1160: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2316,
        in1(1) => DP_OF_in_3,
        out1 => S2323
    );
nand_n_1161: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2323,
        in1(1) => S2322,
        out1 => S2312
    );
dff_51: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S2309,
        NbarT => '0',
        PRE => '0',
        Q => DP_IMM1_in1_0,
        Si => S3340,
        global_reset => '0'
    );
dff_52: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S2310,
        NbarT => '0',
        PRE => '0',
        Q => DP_IMM1_in1_1,
        Si => S3339,
        global_reset => '0'
    );
dff_53: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S2311,
        NbarT => '0',
        PRE => '0',
        Q => DP_IMM1_in1_2,
        Si => S3338,
        global_reset => '0'
    );
dff_54: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S2312,
        NbarT => '0',
        PRE => '0',
        Q => DP_IMM1_in1_3,
        Si => S3359,
        global_reset => '0'
    );
notg_344: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_ldPC,
        out1 => S2341
    );
nor_n_849: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => CU_ldPC,
        in1(1) => S15,
        out1 => S2342
    );
nand_n_1162: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2342,
        in1(1) => DP_INC_1_in_0,
        out1 => S2343
    );
nor_n_850: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2341,
        in1(1) => S16,
        out1 => S2344
    );
nand_n_1163: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2344,
        in1(1) => DP_PC_in_0,
        out1 => S2345
    );
nand_n_1164: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2345,
        in1(1) => S2343,
        out1 => S2324
    );
nand_n_1165: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2342,
        in1(1) => DP_INC_1_in_1,
        out1 => S2346
    );
nand_n_1166: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2344,
        in1(1) => DP_PC_in_1,
        out1 => S2347
    );
nand_n_1167: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2347,
        in1(1) => S2346,
        out1 => S2325
    );
nand_n_1168: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2342,
        in1(1) => DP_INC_1_in_2,
        out1 => S2348
    );
nand_n_1169: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2344,
        in1(1) => DP_PC_in_2,
        out1 => S2349
    );
nand_n_1170: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2349,
        in1(1) => S2348,
        out1 => S2326
    );
nand_n_1171: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2342,
        in1(1) => DP_INC_1_in_3,
        out1 => S2350
    );
nand_n_1172: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2344,
        in1(1) => DP_PC_in_3,
        out1 => S2351
    );
nand_n_1173: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2351,
        in1(1) => S2350,
        out1 => S2327
    );
nand_n_1174: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2342,
        in1(1) => DP_INC_1_in_4,
        out1 => S2352
    );
nand_n_1175: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2344,
        in1(1) => DP_PC_in_4,
        out1 => S2353
    );
nand_n_1176: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2353,
        in1(1) => S2352,
        out1 => S2328
    );
nand_n_1177: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2342,
        in1(1) => DP_INC_1_in_5,
        out1 => S2354
    );
nand_n_1178: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2344,
        in1(1) => DP_PC_in_5,
        out1 => S2355
    );
nand_n_1179: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2355,
        in1(1) => S2354,
        out1 => S2329
    );
nand_n_1180: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2342,
        in1(1) => DP_INC_1_in_6,
        out1 => S2356
    );
nand_n_1181: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2344,
        in1(1) => DP_PC_in_6,
        out1 => S2357
    );
nand_n_1182: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2357,
        in1(1) => S2356,
        out1 => S2330
    );
nand_n_1183: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2342,
        in1(1) => DP_INC_1_in_7,
        out1 => S2358
    );
nand_n_1184: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2344,
        in1(1) => DP_PC_in_7,
        out1 => S2359
    );
nand_n_1185: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2359,
        in1(1) => S2358,
        out1 => S2331
    );
nand_n_1186: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2342,
        in1(1) => DP_INC_1_in_8,
        out1 => S2360
    );
nand_n_1187: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2344,
        in1(1) => DP_PC_in_8,
        out1 => S2361
    );
nand_n_1188: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2361,
        in1(1) => S2360,
        out1 => S2332
    );
nand_n_1189: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2342,
        in1(1) => DP_INC_1_in_9,
        out1 => S2362
    );
nand_n_1190: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2344,
        in1(1) => DP_PC_in_9,
        out1 => S2363
    );
nand_n_1191: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2363,
        in1(1) => S2362,
        out1 => S2333
    );
nand_n_1192: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2342,
        in1(1) => DP_INC_1_in_10,
        out1 => S2364
    );
nand_n_1193: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2344,
        in1(1) => DP_PC_in_10,
        out1 => S2365
    );
nand_n_1194: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2365,
        in1(1) => S2364,
        out1 => S2334
    );
nand_n_1195: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2342,
        in1(1) => DP_INC_1_in_11,
        out1 => S2366
    );
nand_n_1196: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2344,
        in1(1) => DP_PC_in_11,
        out1 => S2367
    );
nand_n_1197: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2367,
        in1(1) => S2366,
        out1 => S2335
    );
nand_n_1198: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2342,
        in1(1) => DP_INC_1_in_12,
        out1 => S2368
    );
nand_n_1199: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2344,
        in1(1) => DP_PC_in_12,
        out1 => S2369
    );
nand_n_1200: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2369,
        in1(1) => S2368,
        out1 => S2336
    );
nand_n_1201: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2342,
        in1(1) => DP_INC_1_in_13,
        out1 => S2370
    );
nand_n_1202: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2344,
        in1(1) => DP_PC_in_13,
        out1 => S2371
    );
nand_n_1203: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2371,
        in1(1) => S2370,
        out1 => S2337
    );
nand_n_1204: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2342,
        in1(1) => DP_INC_1_in_14,
        out1 => S2372
    );
nand_n_1205: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2344,
        in1(1) => DP_PC_in_14,
        out1 => S2373
    );
nand_n_1206: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2373,
        in1(1) => S2372,
        out1 => S2338
    );
nand_n_1207: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2342,
        in1(1) => DP_INC_1_in_15,
        out1 => S2374
    );
nand_n_1208: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2344,
        in1(1) => DP_PC_in_15,
        out1 => S2340
    );
nand_n_1209: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2340,
        in1(1) => S2374,
        out1 => S2339
    );
dff_55: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S2324,
        NbarT => '0',
        PRE => '0',
        Q => DP_INC_1_in_0,
        Si => S3355,
        global_reset => '0'
    );
dff_56: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S2325,
        NbarT => '0',
        PRE => '0',
        Q => DP_INC_1_in_1,
        Si => S3354,
        global_reset => '0'
    );
dff_57: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S2326,
        NbarT => '0',
        PRE => '0',
        Q => DP_INC_1_in_2,
        Si => S3353,
        global_reset => '0'
    );
dff_58: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S2327,
        NbarT => '0',
        PRE => '0',
        Q => DP_INC_1_in_3,
        Si => S3352,
        global_reset => '0'
    );
dff_59: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S2328,
        NbarT => '0',
        PRE => '0',
        Q => DP_INC_1_in_4,
        Si => S3351,
        global_reset => '0'
    );
dff_60: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S2329,
        NbarT => '0',
        PRE => '0',
        Q => DP_INC_1_in_5,
        Si => S3350,
        global_reset => '0'
    );
dff_61: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S2330,
        NbarT => '0',
        PRE => '0',
        Q => DP_INC_1_in_6,
        Si => S3349,
        global_reset => '0'
    );
dff_62: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S2331,
        NbarT => '0',
        PRE => '0',
        Q => DP_INC_1_in_7,
        Si => S3348,
        global_reset => '0'
    );
dff_63: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S2332,
        NbarT => '0',
        PRE => '0',
        Q => DP_INC_1_in_8,
        Si => S3347,
        global_reset => '0'
    );
dff_64: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S2333,
        NbarT => '0',
        PRE => '0',
        Q => DP_INC_1_in_9,
        Si => S3346,
        global_reset => '0'
    );
dff_65: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S2334,
        NbarT => '0',
        PRE => '0',
        Q => DP_INC_1_in_10,
        Si => S3345,
        global_reset => '0'
    );
dff_66: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S2335,
        NbarT => '0',
        PRE => '0',
        Q => DP_INC_1_in_11,
        Si => S3344,
        global_reset => '0'
    );
dff_67: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S2336,
        NbarT => '0',
        PRE => '0',
        Q => DP_INC_1_in_12,
        Si => S3343,
        global_reset => '0'
    );
dff_68: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S2337,
        NbarT => '0',
        PRE => '0',
        Q => DP_INC_1_in_13,
        Si => S3342,
        global_reset => '0'
    );
dff_69: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S2338,
        NbarT => '0',
        PRE => '0',
        Q => DP_INC_1_in_14,
        Si => S3341,
        global_reset => '0'
    );
dff_70: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S2339,
        NbarT => '0',
        PRE => '0',
        Q => DP_INC_1_in_15,
        Si => S3360,
        global_reset => '0'
    );
notg_345: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_SR_C_out,
        out1 => S2377
    );
nand_n_1210: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_SR_C_in,
        in1(1) => CU_ldSR_1,
        out1 => S2378
    );
notg_346: ENTITY WORK.notg
    PORT MAP (
        in1 => S2378,
        out1 => S2379
    );
nor_n_851: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2377,
        in1(1) => CU_ldSR_1,
        out1 => S2380
    );
nor_n_852: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2380,
        in1(1) => S2379,
        out1 => S2376
    );
nor_n_853: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2376,
        in1(1) => S17,
        out1 => S2375
    );
dff_71: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S2375,
        NbarT => '0',
        PRE => '0',
        Q => DP_SR_C_out,
        Si => S3361,
        global_reset => '0'
    );
notg_347: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_SR_N_out,
        out1 => S2383
    );
nand_n_1211: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_SR_N_in,
        in1(1) => CU_ldSR_2,
        out1 => S2384
    );
notg_348: ENTITY WORK.notg
    PORT MAP (
        in1 => S2384,
        out1 => S2385
    );
nor_n_854: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2383,
        in1(1) => CU_ldSR_2,
        out1 => S2386
    );
nor_n_855: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2386,
        in1(1) => S2385,
        out1 => S2382
    );
nor_n_856: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2382,
        in1(1) => S18,
        out1 => S2381
    );
dff_72: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S2381,
        NbarT => '0',
        PRE => '0',
        Q => DP_SR_N_out,
        Si => S3362,
        global_reset => '0'
    );
notg_349: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_SR_V_out,
        out1 => S2389
    );
nand_n_1212: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_SR_V_in,
        in1(1) => CU_ldSR_0,
        out1 => S2390
    );
notg_350: ENTITY WORK.notg
    PORT MAP (
        in1 => S2390,
        out1 => S2391
    );
nor_n_857: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2389,
        in1(1) => CU_ldSR_0,
        out1 => S2392
    );
nor_n_858: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2392,
        in1(1) => S2391,
        out1 => S2388
    );
nor_n_859: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2388,
        in1(1) => S19,
        out1 => S2387
    );
dff_73: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S2387,
        NbarT => '0',
        PRE => '0',
        Q => DP_SR_V_out,
        Si => S3363,
        global_reset => '0'
    );
notg_351: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_SR_Z_out,
        out1 => S2395
    );
nand_n_1213: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_SR_Z_in,
        in1(1) => CU_ldSR_3,
        out1 => S2396
    );
notg_352: ENTITY WORK.notg
    PORT MAP (
        in1 => S2396,
        out1 => S2397
    );
nor_n_860: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2395,
        in1(1) => CU_ldSR_3,
        out1 => S2398
    );
nor_n_861: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2398,
        in1(1) => S2397,
        out1 => S2394
    );
nor_n_862: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2394,
        in1(1) => S20,
        out1 => S2393
    );
dff_74: ENTITY WORK.dff
    PORT MAP (
        C => CU_clk,
        CE => '1',
        CLR => CU_rst,
        D => S2393,
        NbarT => '0',
        PRE => '0',
        Q => DP_SR_Z_out,
        Si => S3364,
        global_reset => '0'
    );
notg_353: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_sel1_ARU,
        out1 => S2416
    );
nand_n_1214: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_sel1_ARU,
        in1(1) => S3,
        out1 => S2417
    );
nand_n_1215: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2416,
        in1(1) => DP_LGU1_in1_0,
        out1 => S2418
    );
nand_n_1216: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2418,
        in1(1) => S2417,
        out1 => S2399
    );
nand_n_1217: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S21,
        in1(1) => CU_sel1_ARU,
        out1 => S2419
    );
nand_n_1218: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_in1_1,
        in1(1) => S2416,
        out1 => S2420
    );
nand_n_1219: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2420,
        in1(1) => S2419,
        out1 => S2406
    );
nand_n_1220: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S22,
        in1(1) => CU_sel1_ARU,
        out1 => S2421
    );
nand_n_1221: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_in1_2,
        in1(1) => S2416,
        out1 => S2422
    );
nand_n_1222: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2422,
        in1(1) => S2421,
        out1 => S2407
    );
nand_n_1223: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S23,
        in1(1) => CU_sel1_ARU,
        out1 => S2423
    );
nand_n_1224: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_in1_3,
        in1(1) => S2416,
        out1 => S2424
    );
nand_n_1225: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2424,
        in1(1) => S2423,
        out1 => S2408
    );
nand_n_1226: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S24,
        in1(1) => CU_sel1_ARU,
        out1 => S2425
    );
nand_n_1227: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_in1_4,
        in1(1) => S2416,
        out1 => S2426
    );
nand_n_1228: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2426,
        in1(1) => S2425,
        out1 => S2409
    );
nand_n_1229: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S25,
        in1(1) => CU_sel1_ARU,
        out1 => S2427
    );
nand_n_1230: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_in1_5,
        in1(1) => S2416,
        out1 => S2428
    );
nand_n_1231: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2428,
        in1(1) => S2427,
        out1 => S2410
    );
nand_n_1232: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S26,
        in1(1) => CU_sel1_ARU,
        out1 => S2429
    );
nand_n_1233: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_in1_6,
        in1(1) => S2416,
        out1 => S2430
    );
nand_n_1234: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2430,
        in1(1) => S2429,
        out1 => S2411
    );
nand_n_1235: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S27,
        in1(1) => CU_sel1_ARU,
        out1 => S2431
    );
nand_n_1236: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_in1_7,
        in1(1) => S2416,
        out1 => S2432
    );
nand_n_1237: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2432,
        in1(1) => S2431,
        out1 => S2412
    );
nand_n_1238: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S28,
        in1(1) => CU_sel1_ARU,
        out1 => S2433
    );
nand_n_1239: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_in1_8,
        in1(1) => S2416,
        out1 => S2434
    );
nand_n_1240: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2434,
        in1(1) => S2433,
        out1 => S2413
    );
nand_n_1241: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S29,
        in1(1) => CU_sel1_ARU,
        out1 => S2435
    );
nand_n_1242: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_in1_9,
        in1(1) => S2416,
        out1 => S2436
    );
nand_n_1243: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2436,
        in1(1) => S2435,
        out1 => S2414
    );
nand_n_1244: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S30,
        in1(1) => CU_sel1_ARU,
        out1 => S2437
    );
nand_n_1245: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_in1_10,
        in1(1) => S2416,
        out1 => S2438
    );
nand_n_1246: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2438,
        in1(1) => S2437,
        out1 => S2400
    );
nand_n_1247: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S31,
        in1(1) => CU_sel1_ARU,
        out1 => S2439
    );
nand_n_1248: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_in1_11,
        in1(1) => S2416,
        out1 => S2440
    );
nand_n_1249: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2440,
        in1(1) => S2439,
        out1 => S2401
    );
nand_n_1250: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S32,
        in1(1) => CU_sel1_ARU,
        out1 => S2441
    );
nand_n_1251: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_in1_12,
        in1(1) => S2416,
        out1 => S2442
    );
nand_n_1252: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2442,
        in1(1) => S2441,
        out1 => S2402
    );
nand_n_1253: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S33,
        in1(1) => CU_sel1_ARU,
        out1 => S2443
    );
nand_n_1254: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_in1_13,
        in1(1) => S2416,
        out1 => S2444
    );
nand_n_1255: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2444,
        in1(1) => S2443,
        out1 => S2403
    );
nand_n_1256: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S34,
        in1(1) => CU_sel1_ARU,
        out1 => S2445
    );
nand_n_1257: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_in1_14,
        in1(1) => S2416,
        out1 => S2446
    );
nand_n_1258: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2446,
        in1(1) => S2445,
        out1 => S2404
    );
nand_n_1259: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S35,
        in1(1) => CU_sel1_ARU,
        out1 => S2447
    );
nand_n_1260: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_in1_15,
        in1(1) => S2416,
        out1 => S2448
    );
nand_n_1261: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2448,
        in1(1) => S2447,
        out1 => S2405
    );
nor_n_863: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => CU_selARU_SR,
        in1(1) => CU_sel1_ARU,
        out1 => S2415
    );
$_DLATCH_N__51: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2399,
        E => S2415,
        Q => DP_ARU1_in1_0
    );
$_DLATCH_N__52: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2406,
        E => S2415,
        Q => DP_ARU1_in1_1
    );
$_DLATCH_N__53: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2407,
        E => S2415,
        Q => DP_ARU1_in1_2
    );
$_DLATCH_N__54: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2408,
        E => S2415,
        Q => DP_ARU1_in1_3
    );
$_DLATCH_N__55: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2409,
        E => S2415,
        Q => DP_ARU1_in1_4
    );
$_DLATCH_N__56: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2410,
        E => S2415,
        Q => DP_ARU1_in1_5
    );
$_DLATCH_N__57: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2411,
        E => S2415,
        Q => DP_ARU1_in1_6
    );
$_DLATCH_N__58: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2412,
        E => S2415,
        Q => DP_ARU1_in1_7
    );
$_DLATCH_N__59: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2413,
        E => S2415,
        Q => DP_ARU1_in1_8
    );
$_DLATCH_N__60: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2414,
        E => S2415,
        Q => DP_ARU1_in1_9
    );
$_DLATCH_N__61: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2400,
        E => S2415,
        Q => DP_ARU1_in1_10
    );
$_DLATCH_N__62: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2401,
        E => S2415,
        Q => DP_ARU1_in1_11
    );
$_DLATCH_N__63: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2402,
        E => S2415,
        Q => DP_ARU1_in1_12
    );
$_DLATCH_N__64: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2403,
        E => S2415,
        Q => DP_ARU1_in1_13
    );
$_DLATCH_N__65: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2404,
        E => S2415,
        Q => DP_ARU1_in1_14
    );
$_DLATCH_N__66: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2405,
        E => S2415,
        Q => DP_ARU1_in1_15
    );
notg_354: ENTITY WORK.notg
    PORT MAP (
        in1 => 'z',
        out1 => S2454
    );
notg_355: ENTITY WORK.notg
    PORT MAP (
        in1 => 'z',
        out1 => S2455
    );
notg_356: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_selLGU_SR,
        out1 => S2456
    );
notg_357: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_inst_0,
        out1 => S2457
    );
notg_358: ENTITY WORK.notg
    PORT MAP (
        in1 => 'z',
        out1 => S2458
    );
notg_359: ENTITY WORK.notg
    PORT MAP (
        in1 => 'z',
        out1 => S2459
    );
notg_360: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_inst_1,
        out1 => S2460
    );
notg_361: ENTITY WORK.notg
    PORT MAP (
        in1 => 'z',
        out1 => S2461
    );
notg_362: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_LGU1_N,
        out1 => S2462
    );
notg_363: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_inst_2,
        out1 => S2463
    );
notg_364: ENTITY WORK.notg
    PORT MAP (
        in1 => 'z',
        out1 => S2464
    );
notg_365: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_LGU1_Z,
        out1 => S2465
    );
notg_366: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_inst_3,
        out1 => S2466
    );
notg_367: ENTITY WORK.notg
    PORT MAP (
        in1 => 'z',
        out1 => S2467
    );
nor_n_864: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => CU_selSET_SR,
        in1(1) => CU_selLGU_SR,
        out1 => S2468
    );
nor_n_865: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => CU_selARU_SR,
        in1(1) => S2454,
        out1 => S2469
    );
nand_n_1262: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_selARU_SR,
        in1(1) => DP_ARU1_V,
        out1 => S2470
    );
nand_n_1263: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2470,
        in1(1) => S2468,
        out1 => S2471
    );
nor_n_866: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2471,
        in1(1) => S2469,
        out1 => S2472
    );
nand_n_1264: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_selSET_SR,
        in1(1) => S2457,
        out1 => S2473
    );
nor_n_867: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => CU_selSET_SR,
        in1(1) => S2456,
        out1 => S2474
    );
nand_n_1265: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2474,
        in1(1) => S2455,
        out1 => S2475
    );
nand_n_1266: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2475,
        in1(1) => S2473,
        out1 => S2476
    );
nor_n_868: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2476,
        in1(1) => S2472,
        out1 => S2449
    );
nor_n_869: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2458,
        in1(1) => CU_selARU_SR,
        out1 => S2477
    );
nand_n_1267: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_C,
        in1(1) => CU_selARU_SR,
        out1 => S2478
    );
nand_n_1268: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2478,
        in1(1) => S2468,
        out1 => S2479
    );
nor_n_870: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2479,
        in1(1) => S2477,
        out1 => S2480
    );
nand_n_1269: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2460,
        in1(1) => CU_selSET_SR,
        out1 => S2481
    );
nand_n_1270: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2474,
        in1(1) => S2459,
        out1 => S2482
    );
nand_n_1271: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2482,
        in1(1) => S2481,
        out1 => S2483
    );
nor_n_871: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2483,
        in1(1) => S2480,
        out1 => S2450
    );
nor_n_872: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2461,
        in1(1) => CU_selARU_SR,
        out1 => S2484
    );
nand_n_1272: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_N,
        in1(1) => CU_selARU_SR,
        out1 => S2485
    );
nand_n_1273: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2485,
        in1(1) => S2468,
        out1 => S2486
    );
nor_n_873: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2486,
        in1(1) => S2484,
        out1 => S2487
    );
nand_n_1274: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2463,
        in1(1) => CU_selSET_SR,
        out1 => S2488
    );
nand_n_1275: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2474,
        in1(1) => S2462,
        out1 => S2489
    );
nand_n_1276: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2489,
        in1(1) => S2488,
        out1 => S2490
    );
nor_n_874: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2490,
        in1(1) => S2487,
        out1 => S2451
    );
nor_n_875: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2464,
        in1(1) => CU_selARU_SR,
        out1 => S2491
    );
nand_n_1277: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_Z,
        in1(1) => CU_selARU_SR,
        out1 => S2492
    );
nand_n_1278: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2492,
        in1(1) => S2468,
        out1 => S2493
    );
nor_n_876: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2493,
        in1(1) => S2491,
        out1 => S2494
    );
nand_n_1279: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2466,
        in1(1) => CU_selSET_SR,
        out1 => S2495
    );
nand_n_1280: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2474,
        in1(1) => S2465,
        out1 => S2496
    );
nand_n_1281: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2496,
        in1(1) => S2495,
        out1 => S2497
    );
nor_n_877: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2497,
        in1(1) => S2494,
        out1 => S2452
    );
nand_n_1282: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2468,
        in1(1) => S2467,
        out1 => S2498
    );
nor_n_878: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2498,
        in1(1) => CU_selARU_SR,
        out1 => S2453
    );
$_DLATCH_N__67: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2449,
        E => S2453,
        Q => DP_SR_V_in
    );
$_DLATCH_N__68: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2450,
        E => S2453,
        Q => DP_SR_C_in
    );
$_DLATCH_N__69: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2451,
        E => S2453,
        Q => DP_SR_N_in
    );
$_DLATCH_N__70: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2452,
        E => S2453,
        Q => DP_SR_Z_in
    );
notg_368: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_selIMM_LGU,
        out1 => S2516
    );
nand_n_1283: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_selIMM_LGU,
        in1(1) => DP_IMM1_out_0,
        out1 => S2517
    );
nand_n_1284: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2516,
        in1(1) => dataBus(0),
        out1 => S2518
    );
nand_n_1285: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2518,
        in1(1) => S2517,
        out1 => S2499
    );
nand_n_1286: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_IMM1_out_1,
        in1(1) => CU_selIMM_LGU,
        out1 => S2519
    );
nand_n_1287: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => dataBus(1),
        in1(1) => S2516,
        out1 => S2520
    );
nand_n_1288: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2520,
        in1(1) => S2519,
        out1 => S2506
    );
nand_n_1289: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_IMM1_out_2,
        in1(1) => CU_selIMM_LGU,
        out1 => S2521
    );
nand_n_1290: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => dataBus(2),
        in1(1) => S2516,
        out1 => S2522
    );
nand_n_1291: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2522,
        in1(1) => S2521,
        out1 => S2507
    );
nand_n_1292: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_IMM1_out_3,
        in1(1) => CU_selIMM_LGU,
        out1 => S2523
    );
nand_n_1293: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => dataBus(3),
        in1(1) => S2516,
        out1 => S2524
    );
nand_n_1294: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2524,
        in1(1) => S2523,
        out1 => S2508
    );
nand_n_1295: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_IMM1_out_4,
        in1(1) => CU_selIMM_LGU,
        out1 => S2525
    );
nand_n_1296: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => dataBus(4),
        in1(1) => S2516,
        out1 => S2526
    );
nand_n_1297: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2526,
        in1(1) => S2525,
        out1 => S2509
    );
nand_n_1298: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_IMM1_out_5,
        in1(1) => CU_selIMM_LGU,
        out1 => S2527
    );
nand_n_1299: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => dataBus(5),
        in1(1) => S2516,
        out1 => S2528
    );
nand_n_1300: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2528,
        in1(1) => S2527,
        out1 => S2510
    );
nand_n_1301: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_IMM1_out_6,
        in1(1) => CU_selIMM_LGU,
        out1 => S2529
    );
nand_n_1302: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => dataBus(6),
        in1(1) => S2516,
        out1 => S2530
    );
nand_n_1303: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2530,
        in1(1) => S2529,
        out1 => S2511
    );
nand_n_1304: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_IMM1_out_7,
        in1(1) => CU_selIMM_LGU,
        out1 => S2531
    );
nand_n_1305: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => dataBus(7),
        in1(1) => S2516,
        out1 => S2532
    );
nand_n_1306: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2532,
        in1(1) => S2531,
        out1 => S2512
    );
nand_n_1307: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_IMM1_out_8,
        in1(1) => CU_selIMM_LGU,
        out1 => S2533
    );
nand_n_1308: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => dataBus(8),
        in1(1) => S2516,
        out1 => S2534
    );
nand_n_1309: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2534,
        in1(1) => S2533,
        out1 => S2513
    );
nand_n_1310: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_IMM1_out_9,
        in1(1) => CU_selIMM_LGU,
        out1 => S2535
    );
nand_n_1311: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => dataBus(9),
        in1(1) => S2516,
        out1 => S2536
    );
nand_n_1312: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2536,
        in1(1) => S2535,
        out1 => S2514
    );
nand_n_1313: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_IMM1_out_10,
        in1(1) => CU_selIMM_LGU,
        out1 => S2537
    );
nand_n_1314: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => dataBus(10),
        in1(1) => S2516,
        out1 => S2538
    );
nand_n_1315: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2538,
        in1(1) => S2537,
        out1 => S2500
    );
nand_n_1316: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_IMM1_out_11,
        in1(1) => CU_selIMM_LGU,
        out1 => S2539
    );
nand_n_1317: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => dataBus(11),
        in1(1) => S2516,
        out1 => S2540
    );
nand_n_1318: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2540,
        in1(1) => S2539,
        out1 => S2501
    );
nand_n_1319: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_IMM1_out_12,
        in1(1) => CU_selIMM_LGU,
        out1 => S2541
    );
nand_n_1320: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => dataBus(12),
        in1(1) => S2516,
        out1 => S2542
    );
nand_n_1321: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2542,
        in1(1) => S2541,
        out1 => S2502
    );
nand_n_1322: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_IMM1_out_13,
        in1(1) => CU_selIMM_LGU,
        out1 => S2543
    );
nand_n_1323: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => dataBus(13),
        in1(1) => S2516,
        out1 => S2544
    );
nand_n_1324: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2544,
        in1(1) => S2543,
        out1 => S2503
    );
nand_n_1325: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_IMM1_out_14,
        in1(1) => CU_selIMM_LGU,
        out1 => S2545
    );
nand_n_1326: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => dataBus(14),
        in1(1) => S2516,
        out1 => S2546
    );
nand_n_1327: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2546,
        in1(1) => S2545,
        out1 => S2504
    );
nand_n_1328: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_IMM1_out_15,
        in1(1) => CU_selIMM_LGU,
        out1 => S2547
    );
nand_n_1329: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => dataBus(15),
        in1(1) => S2516,
        out1 => S2548
    );
nand_n_1330: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2548,
        in1(1) => S2547,
        out1 => S2505
    );
nor_n_879: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => CU_selMEM_LGU,
        in1(1) => CU_selIMM_LGU,
        out1 => S2515
    );
$_DLATCH_N__71: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2499,
        E => S2515,
        Q => DP_LGU1_in1_0
    );
$_DLATCH_N__72: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2506,
        E => S2515,
        Q => DP_LGU1_in1_1
    );
$_DLATCH_N__73: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2507,
        E => S2515,
        Q => DP_LGU1_in1_2
    );
$_DLATCH_N__74: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2508,
        E => S2515,
        Q => DP_LGU1_in1_3
    );
$_DLATCH_N__75: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2509,
        E => S2515,
        Q => DP_LGU1_in1_4
    );
$_DLATCH_N__76: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2510,
        E => S2515,
        Q => DP_LGU1_in1_5
    );
$_DLATCH_N__77: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2511,
        E => S2515,
        Q => DP_LGU1_in1_6
    );
$_DLATCH_N__78: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2512,
        E => S2515,
        Q => DP_LGU1_in1_7
    );
$_DLATCH_N__79: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2513,
        E => S2515,
        Q => DP_LGU1_in1_8
    );
$_DLATCH_N__80: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2514,
        E => S2515,
        Q => DP_LGU1_in1_9
    );
$_DLATCH_N__81: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2500,
        E => S2515,
        Q => DP_LGU1_in1_10
    );
$_DLATCH_N__82: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2501,
        E => S2515,
        Q => DP_LGU1_in1_11
    );
$_DLATCH_N__83: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2502,
        E => S2515,
        Q => DP_LGU1_in1_12
    );
$_DLATCH_N__84: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2503,
        E => S2515,
        Q => DP_LGU1_in1_13
    );
$_DLATCH_N__85: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2504,
        E => S2515,
        Q => DP_LGU1_in1_14
    );
$_DLATCH_N__86: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2505,
        E => S2515,
        Q => DP_LGU1_in1_15
    );
notg_369: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_selARU_AC,
        out1 => S2703
    );
notg_370: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(0),
        out1 => S2704
    );
notg_371: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_selMEM_AC,
        out1 => S2705
    );
notg_372: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IMM1_out_0,
        out1 => S2706
    );
notg_373: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_selIMM_AC,
        out1 => S2707
    );
notg_374: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(1),
        out1 => S2708
    );
notg_375: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IMM1_out_1,
        out1 => S2709
    );
notg_376: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(2),
        out1 => S2710
    );
notg_377: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IMM1_out_2,
        out1 => S2711
    );
notg_378: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(3),
        out1 => S2712
    );
notg_379: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IMM1_out_3,
        out1 => S2713
    );
notg_380: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(4),
        out1 => S2714
    );
notg_381: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IMM1_out_4,
        out1 => S2715
    );
notg_382: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(5),
        out1 => S2716
    );
notg_383: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IMM1_out_5,
        out1 => S2566
    );
notg_384: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(6),
        out1 => S2567
    );
notg_385: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IMM1_out_6,
        out1 => S2568
    );
notg_386: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(7),
        out1 => S2569
    );
notg_387: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IMM1_out_7,
        out1 => S2570
    );
notg_388: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(8),
        out1 => S2571
    );
notg_389: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IMM1_out_8,
        out1 => S2572
    );
notg_390: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(9),
        out1 => S2573
    );
notg_391: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IMM1_out_9,
        out1 => S2574
    );
notg_392: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(10),
        out1 => S2575
    );
notg_393: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IMM1_out_10,
        out1 => S2576
    );
notg_394: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(11),
        out1 => S2577
    );
notg_395: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IMM1_out_11,
        out1 => S2578
    );
notg_396: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(12),
        out1 => S2579
    );
notg_397: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IMM1_out_12,
        out1 => S2580
    );
notg_398: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(13),
        out1 => S2581
    );
notg_399: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IMM1_out_13,
        out1 => S2582
    );
notg_400: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(14),
        out1 => S2583
    );
notg_401: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IMM1_out_14,
        out1 => S2584
    );
notg_402: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(15),
        out1 => S2585
    );
notg_403: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IMM1_out_15,
        out1 => S2586
    );
notg_404: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_selLGU_AC,
        out1 => S2587
    );
nand_n_1331: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2707,
        in1(1) => S2705,
        out1 => S2588
    );
nand_n_1332: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_selARU_AC,
        in1(1) => DP_ARU1_out_0,
        out1 => S2589
    );
nand_n_1333: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2703,
        in1(1) => DP_LGU1_out_0,
        out1 => S2590
    );
nand_n_1334: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2590,
        in1(1) => S2589,
        out1 => S2591
    );
nor_n_880: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2591,
        in1(1) => S2588,
        out1 => S2592
    );
nand_n_1335: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_selIMM_AC,
        in1(1) => S2706,
        out1 => S2593
    );
nor_n_881: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => CU_selIMM_AC,
        in1(1) => S2705,
        out1 => S2594
    );
nand_n_1336: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2594,
        in1(1) => S2704,
        out1 => S2595
    );
nand_n_1337: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2595,
        in1(1) => S2593,
        out1 => S2596
    );
nor_n_882: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2596,
        in1(1) => S2592,
        out1 => S2549
    );
nand_n_1338: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_out_1,
        in1(1) => S2703,
        out1 => S2597
    );
nand_n_1339: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_out_1,
        in1(1) => CU_selARU_AC,
        out1 => S2598
    );
nand_n_1340: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2598,
        in1(1) => S2597,
        out1 => S2599
    );
nor_n_883: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2599,
        in1(1) => S2588,
        out1 => S2600
    );
nand_n_1341: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2709,
        in1(1) => CU_selIMM_AC,
        out1 => S2601
    );
nand_n_1342: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2594,
        in1(1) => S2708,
        out1 => S2602
    );
nand_n_1343: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2602,
        in1(1) => S2601,
        out1 => S2603
    );
nor_n_884: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2603,
        in1(1) => S2600,
        out1 => S2556
    );
nand_n_1344: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_out_2,
        in1(1) => S2703,
        out1 => S2604
    );
nand_n_1345: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_out_2,
        in1(1) => CU_selARU_AC,
        out1 => S2605
    );
nand_n_1346: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2605,
        in1(1) => S2604,
        out1 => S2606
    );
nor_n_885: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2606,
        in1(1) => S2588,
        out1 => S2607
    );
nand_n_1347: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2711,
        in1(1) => CU_selIMM_AC,
        out1 => S2608
    );
nand_n_1348: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2594,
        in1(1) => S2710,
        out1 => S2609
    );
nand_n_1349: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2609,
        in1(1) => S2608,
        out1 => S2610
    );
nor_n_886: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2610,
        in1(1) => S2607,
        out1 => S2557
    );
nand_n_1350: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_out_3,
        in1(1) => S2703,
        out1 => S2611
    );
nand_n_1351: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_out_3,
        in1(1) => CU_selARU_AC,
        out1 => S2612
    );
nand_n_1352: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2612,
        in1(1) => S2611,
        out1 => S2613
    );
nor_n_887: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2613,
        in1(1) => S2588,
        out1 => S2614
    );
nand_n_1353: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2713,
        in1(1) => CU_selIMM_AC,
        out1 => S2615
    );
nand_n_1354: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2594,
        in1(1) => S2712,
        out1 => S2616
    );
nand_n_1355: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2616,
        in1(1) => S2615,
        out1 => S2617
    );
nor_n_888: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2617,
        in1(1) => S2614,
        out1 => S2558
    );
nand_n_1356: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_out_4,
        in1(1) => S2703,
        out1 => S2618
    );
nand_n_1357: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_out_4,
        in1(1) => CU_selARU_AC,
        out1 => S2619
    );
nand_n_1358: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2619,
        in1(1) => S2618,
        out1 => S2620
    );
nor_n_889: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2620,
        in1(1) => S2588,
        out1 => S2621
    );
nand_n_1359: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2715,
        in1(1) => CU_selIMM_AC,
        out1 => S2622
    );
nand_n_1360: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2594,
        in1(1) => S2714,
        out1 => S2623
    );
nand_n_1361: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2623,
        in1(1) => S2622,
        out1 => S2624
    );
nor_n_890: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2624,
        in1(1) => S2621,
        out1 => S2559
    );
nand_n_1362: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_out_5,
        in1(1) => S2703,
        out1 => S2625
    );
nand_n_1363: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_out_5,
        in1(1) => CU_selARU_AC,
        out1 => S2626
    );
nand_n_1364: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2626,
        in1(1) => S2625,
        out1 => S2627
    );
nor_n_891: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2627,
        in1(1) => S2588,
        out1 => S2628
    );
nand_n_1365: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2566,
        in1(1) => CU_selIMM_AC,
        out1 => S2629
    );
nand_n_1366: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2594,
        in1(1) => S2716,
        out1 => S2630
    );
nand_n_1367: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2630,
        in1(1) => S2629,
        out1 => S2631
    );
nor_n_892: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2631,
        in1(1) => S2628,
        out1 => S2560
    );
nand_n_1368: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_out_6,
        in1(1) => S2703,
        out1 => S2632
    );
nand_n_1369: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_out_6,
        in1(1) => CU_selARU_AC,
        out1 => S2633
    );
nand_n_1370: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2633,
        in1(1) => S2632,
        out1 => S2634
    );
nor_n_893: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2634,
        in1(1) => S2588,
        out1 => S2635
    );
nand_n_1371: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2568,
        in1(1) => CU_selIMM_AC,
        out1 => S2636
    );
nand_n_1372: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2594,
        in1(1) => S2567,
        out1 => S2637
    );
nand_n_1373: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2637,
        in1(1) => S2636,
        out1 => S2638
    );
nor_n_894: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2638,
        in1(1) => S2635,
        out1 => S2561
    );
nand_n_1374: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_out_7,
        in1(1) => S2703,
        out1 => S2639
    );
nand_n_1375: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_out_7,
        in1(1) => CU_selARU_AC,
        out1 => S2640
    );
nand_n_1376: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2640,
        in1(1) => S2639,
        out1 => S2641
    );
nor_n_895: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2641,
        in1(1) => S2588,
        out1 => S2642
    );
nand_n_1377: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2570,
        in1(1) => CU_selIMM_AC,
        out1 => S2643
    );
nand_n_1378: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2594,
        in1(1) => S2569,
        out1 => S2644
    );
nand_n_1379: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2644,
        in1(1) => S2643,
        out1 => S2645
    );
nor_n_896: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2645,
        in1(1) => S2642,
        out1 => S2562
    );
nand_n_1380: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_out_8,
        in1(1) => CU_selARU_AC,
        out1 => S2646
    );
nand_n_1381: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_out_8,
        in1(1) => S2703,
        out1 => S2647
    );
nand_n_1382: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2647,
        in1(1) => S2646,
        out1 => S2648
    );
nor_n_897: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2648,
        in1(1) => S2588,
        out1 => S2649
    );
nand_n_1383: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2572,
        in1(1) => CU_selIMM_AC,
        out1 => S2650
    );
nand_n_1384: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2594,
        in1(1) => S2571,
        out1 => S2651
    );
nand_n_1385: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2651,
        in1(1) => S2650,
        out1 => S2652
    );
nor_n_898: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2652,
        in1(1) => S2649,
        out1 => S2563
    );
nand_n_1386: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_out_9,
        in1(1) => S2703,
        out1 => S2653
    );
nand_n_1387: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_out_9,
        in1(1) => CU_selARU_AC,
        out1 => S2654
    );
nand_n_1388: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2654,
        in1(1) => S2653,
        out1 => S2655
    );
nor_n_899: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2655,
        in1(1) => S2588,
        out1 => S2656
    );
nand_n_1389: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2574,
        in1(1) => CU_selIMM_AC,
        out1 => S2657
    );
nand_n_1390: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2594,
        in1(1) => S2573,
        out1 => S2658
    );
nand_n_1391: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2658,
        in1(1) => S2657,
        out1 => S2659
    );
nor_n_900: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2659,
        in1(1) => S2656,
        out1 => S2564
    );
nand_n_1392: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_out_10,
        in1(1) => CU_selARU_AC,
        out1 => S2660
    );
nand_n_1393: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_out_10,
        in1(1) => S2703,
        out1 => S2661
    );
nand_n_1394: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2661,
        in1(1) => S2660,
        out1 => S2662
    );
nor_n_901: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2662,
        in1(1) => S2588,
        out1 => S2663
    );
nand_n_1395: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2576,
        in1(1) => CU_selIMM_AC,
        out1 => S2664
    );
nand_n_1396: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2594,
        in1(1) => S2575,
        out1 => S2665
    );
nand_n_1397: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2665,
        in1(1) => S2664,
        out1 => S2666
    );
nor_n_902: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2666,
        in1(1) => S2663,
        out1 => S2550
    );
nand_n_1398: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_out_11,
        in1(1) => S2703,
        out1 => S2667
    );
nand_n_1399: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_out_11,
        in1(1) => CU_selARU_AC,
        out1 => S2668
    );
nand_n_1400: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2668,
        in1(1) => S2667,
        out1 => S2669
    );
nor_n_903: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2669,
        in1(1) => S2588,
        out1 => S2670
    );
nand_n_1401: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2578,
        in1(1) => CU_selIMM_AC,
        out1 => S2671
    );
nand_n_1402: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2594,
        in1(1) => S2577,
        out1 => S2672
    );
nand_n_1403: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2672,
        in1(1) => S2671,
        out1 => S2673
    );
nor_n_904: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2673,
        in1(1) => S2670,
        out1 => S2551
    );
nand_n_1404: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_out_12,
        in1(1) => CU_selARU_AC,
        out1 => S2674
    );
nand_n_1405: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_out_12,
        in1(1) => S2703,
        out1 => S2675
    );
nand_n_1406: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2675,
        in1(1) => S2674,
        out1 => S2676
    );
nor_n_905: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2676,
        in1(1) => S2588,
        out1 => S2677
    );
nand_n_1407: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2580,
        in1(1) => CU_selIMM_AC,
        out1 => S2678
    );
nand_n_1408: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2594,
        in1(1) => S2579,
        out1 => S2679
    );
nand_n_1409: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2679,
        in1(1) => S2678,
        out1 => S2680
    );
nor_n_906: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2680,
        in1(1) => S2677,
        out1 => S2552
    );
nand_n_1410: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_out_13,
        in1(1) => S2703,
        out1 => S2681
    );
nand_n_1411: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_out_13,
        in1(1) => CU_selARU_AC,
        out1 => S2682
    );
nand_n_1412: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2682,
        in1(1) => S2681,
        out1 => S2683
    );
nor_n_907: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2683,
        in1(1) => S2588,
        out1 => S2684
    );
nand_n_1413: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2582,
        in1(1) => CU_selIMM_AC,
        out1 => S2685
    );
nand_n_1414: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2594,
        in1(1) => S2581,
        out1 => S2686
    );
nand_n_1415: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2686,
        in1(1) => S2685,
        out1 => S2687
    );
nor_n_908: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2687,
        in1(1) => S2684,
        out1 => S2553
    );
nand_n_1416: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_out_14,
        in1(1) => CU_selARU_AC,
        out1 => S2688
    );
nand_n_1417: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_out_14,
        in1(1) => S2703,
        out1 => S2689
    );
nand_n_1418: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2689,
        in1(1) => S2688,
        out1 => S2690
    );
nor_n_909: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2690,
        in1(1) => S2588,
        out1 => S2691
    );
nand_n_1419: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2584,
        in1(1) => CU_selIMM_AC,
        out1 => S2692
    );
nand_n_1420: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2594,
        in1(1) => S2583,
        out1 => S2693
    );
nand_n_1421: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2693,
        in1(1) => S2692,
        out1 => S2694
    );
nor_n_910: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2694,
        in1(1) => S2691,
        out1 => S2554
    );
nand_n_1422: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_LGU1_N,
        in1(1) => S2703,
        out1 => S2695
    );
nand_n_1423: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_ARU1_N,
        in1(1) => CU_selARU_AC,
        out1 => S2696
    );
nand_n_1424: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2696,
        in1(1) => S2695,
        out1 => S2697
    );
nor_n_911: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2697,
        in1(1) => S2588,
        out1 => S2698
    );
nand_n_1425: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2586,
        in1(1) => CU_selIMM_AC,
        out1 => S2699
    );
nand_n_1426: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2594,
        in1(1) => S2585,
        out1 => S2700
    );
nand_n_1427: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2700,
        in1(1) => S2699,
        out1 => S2701
    );
nor_n_912: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2701,
        in1(1) => S2698,
        out1 => S2555
    );
nand_n_1428: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2587,
        in1(1) => S2703,
        out1 => S2702
    );
nor_n_913: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2702,
        in1(1) => S2588,
        out1 => S2565
    );
$_DLATCH_N__87: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2549,
        E => S2565,
        Q => DP_AC_in_0
    );
$_DLATCH_N__88: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2556,
        E => S2565,
        Q => DP_AC_in_1
    );
$_DLATCH_N__89: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2557,
        E => S2565,
        Q => DP_AC_in_2
    );
$_DLATCH_N__90: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2558,
        E => S2565,
        Q => DP_AC_in_3
    );
$_DLATCH_N__91: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2559,
        E => S2565,
        Q => DP_AC_in_4
    );
$_DLATCH_N__92: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2560,
        E => S2565,
        Q => DP_AC_in_5
    );
$_DLATCH_N__93: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2561,
        E => S2565,
        Q => DP_AC_in_6
    );
$_DLATCH_N__94: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2562,
        E => S2565,
        Q => DP_AC_in_7
    );
$_DLATCH_N__95: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2563,
        E => S2565,
        Q => DP_AC_in_8
    );
$_DLATCH_N__96: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2564,
        E => S2565,
        Q => DP_AC_in_9
    );
$_DLATCH_N__97: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2550,
        E => S2565,
        Q => DP_AC_in_10
    );
$_DLATCH_N__98: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2551,
        E => S2565,
        Q => DP_AC_in_11
    );
$_DLATCH_N__99: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2552,
        E => S2565,
        Q => DP_AC_in_12
    );
$_DLATCH_N__100: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2553,
        E => S2565,
        Q => DP_AC_in_13
    );
$_DLATCH_N__101: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2554,
        E => S2565,
        Q => DP_AC_in_14
    );
$_DLATCH_N__102: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2555,
        E => S2565,
        Q => DP_AC_in_15
    );
notg_405: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_selPC_OF,
        out1 => S2722
    );
nand_n_1429: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_selPC_OF,
        in1(1) => DP_INC_1_in_12,
        out1 => S2723
    );
nand_n_1430: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2722,
        in1(1) => DP_IMM1_out_0,
        out1 => S2724
    );
nand_n_1431: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2724,
        in1(1) => S2723,
        out1 => S2717
    );
nand_n_1432: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_INC_1_in_13,
        in1(1) => CU_selPC_OF,
        out1 => S2725
    );
nand_n_1433: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_IMM1_out_1,
        in1(1) => S2722,
        out1 => S2726
    );
nand_n_1434: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2726,
        in1(1) => S2725,
        out1 => S2718
    );
nand_n_1435: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_INC_1_in_14,
        in1(1) => CU_selPC_OF,
        out1 => S2727
    );
nand_n_1436: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_IMM1_out_2,
        in1(1) => S2722,
        out1 => S2728
    );
nand_n_1437: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2728,
        in1(1) => S2727,
        out1 => S2719
    );
nand_n_1438: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_INC_1_in_15,
        in1(1) => CU_selPC_OF,
        out1 => S2729
    );
nand_n_1439: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_IMM1_out_3,
        in1(1) => S2722,
        out1 => S2730
    );
nand_n_1440: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2730,
        in1(1) => S2729,
        out1 => S2720
    );
nor_n_914: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => CU_selIMM_OF,
        in1(1) => CU_selPC_OF,
        out1 => S2721
    );
$_DLATCH_N__103: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2717,
        E => S2721,
        Q => DP_OF_in_0
    );
$_DLATCH_N__104: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2718,
        E => S2721,
        Q => DP_OF_in_1
    );
$_DLATCH_N__105: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2719,
        E => S2721,
        Q => DP_OF_in_2
    );
$_DLATCH_N__106: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2720,
        E => S2721,
        Q => DP_OF_in_3
    );
notg_406: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_selIMM_PC,
        out1 => S2885
    );
notg_407: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(0),
        out1 => S2886
    );
notg_408: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_selMEM_PC,
        out1 => S2887
    );
notg_409: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_out_0,
        out1 => S2888
    );
notg_410: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_selINC_PC,
        out1 => S2889
    );
notg_411: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(1),
        out1 => S2890
    );
notg_412: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_out_1,
        out1 => S2891
    );
notg_413: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(2),
        out1 => S2892
    );
notg_414: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_out_2,
        out1 => S2893
    );
notg_415: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(3),
        out1 => S2894
    );
notg_416: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_out_3,
        out1 => S2895
    );
notg_417: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(4),
        out1 => S2896
    );
notg_418: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_out_4,
        out1 => S2897
    );
notg_419: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(5),
        out1 => S2898
    );
notg_420: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_out_5,
        out1 => S2748
    );
notg_421: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(6),
        out1 => S2749
    );
notg_422: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_out_6,
        out1 => S2750
    );
notg_423: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(7),
        out1 => S2751
    );
notg_424: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_out_7,
        out1 => S2752
    );
notg_425: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(8),
        out1 => S2753
    );
notg_426: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_out_8,
        out1 => S2754
    );
notg_427: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(9),
        out1 => S2755
    );
notg_428: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_out_9,
        out1 => S2756
    );
notg_429: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(10),
        out1 => S2757
    );
notg_430: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_out_10,
        out1 => S2758
    );
notg_431: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(11),
        out1 => S2759
    );
notg_432: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_out_11,
        out1 => S2760
    );
notg_433: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(12),
        out1 => S2761
    );
notg_434: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_out_12,
        out1 => S2762
    );
notg_435: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(13),
        out1 => S2763
    );
notg_436: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_out_13,
        out1 => S2764
    );
notg_437: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(14),
        out1 => S2765
    );
notg_438: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_out_14,
        out1 => S2766
    );
notg_439: ENTITY WORK.notg
    PORT MAP (
        in1 => dataBus(15),
        out1 => S2767
    );
notg_440: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_out_15,
        out1 => S2768
    );
notg_441: ENTITY WORK.notg
    PORT MAP (
        in1 => 'z',
        out1 => S2769
    );
nand_n_1441: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2889,
        in1(1) => S2887,
        out1 => S2770
    );
nand_n_1442: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_selIMM_PC,
        in1(1) => DP_IMM1_out_0,
        out1 => S2771
    );
nand_n_1443: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2885,
        in1(1) => 'z',
        out1 => S2772
    );
nand_n_1444: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2772,
        in1(1) => S2771,
        out1 => S2773
    );
nor_n_915: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2773,
        in1(1) => S2770,
        out1 => S2774
    );
nand_n_1445: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_selINC_PC,
        in1(1) => S2888,
        out1 => S2775
    );
nor_n_916: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => CU_selINC_PC,
        in1(1) => S2887,
        out1 => S2776
    );
nand_n_1446: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2776,
        in1(1) => S2886,
        out1 => S2777
    );
nand_n_1447: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2777,
        in1(1) => S2775,
        out1 => S2778
    );
nor_n_917: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2778,
        in1(1) => S2774,
        out1 => S2731
    );
nand_n_1448: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S2885,
        out1 => S2779
    );
nand_n_1449: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_IMM1_out_1,
        in1(1) => CU_selIMM_PC,
        out1 => S2780
    );
nand_n_1450: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2780,
        in1(1) => S2779,
        out1 => S2781
    );
nor_n_918: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2781,
        in1(1) => S2770,
        out1 => S2782
    );
nand_n_1451: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2891,
        in1(1) => CU_selINC_PC,
        out1 => S2783
    );
nand_n_1452: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2776,
        in1(1) => S2890,
        out1 => S2784
    );
nand_n_1453: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2784,
        in1(1) => S2783,
        out1 => S2785
    );
nor_n_919: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2785,
        in1(1) => S2782,
        out1 => S2738
    );
nand_n_1454: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S2885,
        out1 => S2786
    );
nand_n_1455: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_IMM1_out_2,
        in1(1) => CU_selIMM_PC,
        out1 => S2787
    );
nand_n_1456: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2787,
        in1(1) => S2786,
        out1 => S2788
    );
nor_n_920: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2788,
        in1(1) => S2770,
        out1 => S2789
    );
nand_n_1457: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2893,
        in1(1) => CU_selINC_PC,
        out1 => S2790
    );
nand_n_1458: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2776,
        in1(1) => S2892,
        out1 => S2791
    );
nand_n_1459: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2791,
        in1(1) => S2790,
        out1 => S2792
    );
nor_n_921: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2792,
        in1(1) => S2789,
        out1 => S2739
    );
nand_n_1460: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S2885,
        out1 => S2793
    );
nand_n_1461: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_IMM1_out_3,
        in1(1) => CU_selIMM_PC,
        out1 => S2794
    );
nand_n_1462: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2794,
        in1(1) => S2793,
        out1 => S2795
    );
nor_n_922: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2795,
        in1(1) => S2770,
        out1 => S2796
    );
nand_n_1463: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2895,
        in1(1) => CU_selINC_PC,
        out1 => S2797
    );
nand_n_1464: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2776,
        in1(1) => S2894,
        out1 => S2798
    );
nand_n_1465: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2798,
        in1(1) => S2797,
        out1 => S2799
    );
nor_n_923: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2799,
        in1(1) => S2796,
        out1 => S2740
    );
nand_n_1466: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S2885,
        out1 => S2800
    );
nand_n_1467: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_IMM1_out_4,
        in1(1) => CU_selIMM_PC,
        out1 => S2801
    );
nand_n_1468: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2801,
        in1(1) => S2800,
        out1 => S2802
    );
nor_n_924: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2802,
        in1(1) => S2770,
        out1 => S2803
    );
nand_n_1469: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2897,
        in1(1) => CU_selINC_PC,
        out1 => S2804
    );
nand_n_1470: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2776,
        in1(1) => S2896,
        out1 => S2805
    );
nand_n_1471: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2805,
        in1(1) => S2804,
        out1 => S2806
    );
nor_n_925: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2806,
        in1(1) => S2803,
        out1 => S2741
    );
nand_n_1472: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S2885,
        out1 => S2807
    );
nand_n_1473: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_IMM1_out_5,
        in1(1) => CU_selIMM_PC,
        out1 => S2808
    );
nand_n_1474: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2808,
        in1(1) => S2807,
        out1 => S2809
    );
nor_n_926: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2809,
        in1(1) => S2770,
        out1 => S2810
    );
nand_n_1475: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2748,
        in1(1) => CU_selINC_PC,
        out1 => S2811
    );
nand_n_1476: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2776,
        in1(1) => S2898,
        out1 => S2812
    );
nand_n_1477: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2812,
        in1(1) => S2811,
        out1 => S2813
    );
nor_n_927: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2813,
        in1(1) => S2810,
        out1 => S2742
    );
nand_n_1478: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S2885,
        out1 => S2814
    );
nand_n_1479: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_IMM1_out_6,
        in1(1) => CU_selIMM_PC,
        out1 => S2815
    );
nand_n_1480: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2815,
        in1(1) => S2814,
        out1 => S2816
    );
nor_n_928: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2816,
        in1(1) => S2770,
        out1 => S2817
    );
nand_n_1481: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2750,
        in1(1) => CU_selINC_PC,
        out1 => S2818
    );
nand_n_1482: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2776,
        in1(1) => S2749,
        out1 => S2819
    );
nand_n_1483: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2819,
        in1(1) => S2818,
        out1 => S2820
    );
nor_n_929: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2820,
        in1(1) => S2817,
        out1 => S2743
    );
nand_n_1484: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S2885,
        out1 => S2821
    );
nand_n_1485: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_IMM1_out_7,
        in1(1) => CU_selIMM_PC,
        out1 => S2822
    );
nand_n_1486: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2822,
        in1(1) => S2821,
        out1 => S2823
    );
nor_n_930: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2823,
        in1(1) => S2770,
        out1 => S2824
    );
nand_n_1487: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2752,
        in1(1) => CU_selINC_PC,
        out1 => S2825
    );
nand_n_1488: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2776,
        in1(1) => S2751,
        out1 => S2826
    );
nand_n_1489: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2826,
        in1(1) => S2825,
        out1 => S2827
    );
nor_n_931: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2827,
        in1(1) => S2824,
        out1 => S2744
    );
nand_n_1490: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_IMM1_out_8,
        in1(1) => CU_selIMM_PC,
        out1 => S2828
    );
nand_n_1491: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S2885,
        out1 => S2829
    );
nand_n_1492: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2829,
        in1(1) => S2828,
        out1 => S2830
    );
nor_n_932: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2830,
        in1(1) => S2770,
        out1 => S2831
    );
nand_n_1493: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2754,
        in1(1) => CU_selINC_PC,
        out1 => S2832
    );
nand_n_1494: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2776,
        in1(1) => S2753,
        out1 => S2833
    );
nand_n_1495: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2833,
        in1(1) => S2832,
        out1 => S2834
    );
nor_n_933: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2834,
        in1(1) => S2831,
        out1 => S2745
    );
nand_n_1496: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S2885,
        out1 => S2835
    );
nand_n_1497: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_IMM1_out_9,
        in1(1) => CU_selIMM_PC,
        out1 => S2836
    );
nand_n_1498: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2836,
        in1(1) => S2835,
        out1 => S2837
    );
nor_n_934: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2837,
        in1(1) => S2770,
        out1 => S2838
    );
nand_n_1499: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2756,
        in1(1) => CU_selINC_PC,
        out1 => S2839
    );
nand_n_1500: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2776,
        in1(1) => S2755,
        out1 => S2840
    );
nand_n_1501: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2840,
        in1(1) => S2839,
        out1 => S2841
    );
nor_n_935: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2841,
        in1(1) => S2838,
        out1 => S2746
    );
nand_n_1502: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_IMM1_out_10,
        in1(1) => CU_selIMM_PC,
        out1 => S2842
    );
nand_n_1503: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S2885,
        out1 => S2843
    );
nand_n_1504: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2843,
        in1(1) => S2842,
        out1 => S2844
    );
nor_n_936: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2844,
        in1(1) => S2770,
        out1 => S2845
    );
nand_n_1505: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2758,
        in1(1) => CU_selINC_PC,
        out1 => S2846
    );
nand_n_1506: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2776,
        in1(1) => S2757,
        out1 => S2847
    );
nand_n_1507: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2847,
        in1(1) => S2846,
        out1 => S2848
    );
nor_n_937: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2848,
        in1(1) => S2845,
        out1 => S2732
    );
nand_n_1508: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S2885,
        out1 => S2849
    );
nand_n_1509: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_IMM1_out_11,
        in1(1) => CU_selIMM_PC,
        out1 => S2850
    );
nand_n_1510: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2850,
        in1(1) => S2849,
        out1 => S2851
    );
nor_n_938: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2851,
        in1(1) => S2770,
        out1 => S2852
    );
nand_n_1511: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2760,
        in1(1) => CU_selINC_PC,
        out1 => S2853
    );
nand_n_1512: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2776,
        in1(1) => S2759,
        out1 => S2854
    );
nand_n_1513: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2854,
        in1(1) => S2853,
        out1 => S2855
    );
nor_n_939: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2855,
        in1(1) => S2852,
        out1 => S2733
    );
nand_n_1514: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_IMM1_out_12,
        in1(1) => CU_selIMM_PC,
        out1 => S2856
    );
nand_n_1515: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S2885,
        out1 => S2857
    );
nand_n_1516: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2857,
        in1(1) => S2856,
        out1 => S2858
    );
nor_n_940: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2858,
        in1(1) => S2770,
        out1 => S2859
    );
nand_n_1517: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2762,
        in1(1) => CU_selINC_PC,
        out1 => S2860
    );
nand_n_1518: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2776,
        in1(1) => S2761,
        out1 => S2861
    );
nand_n_1519: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2861,
        in1(1) => S2860,
        out1 => S2862
    );
nor_n_941: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2862,
        in1(1) => S2859,
        out1 => S2734
    );
nand_n_1520: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S2885,
        out1 => S2863
    );
nand_n_1521: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_IMM1_out_13,
        in1(1) => CU_selIMM_PC,
        out1 => S2864
    );
nand_n_1522: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2864,
        in1(1) => S2863,
        out1 => S2865
    );
nor_n_942: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2865,
        in1(1) => S2770,
        out1 => S2866
    );
nand_n_1523: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2764,
        in1(1) => CU_selINC_PC,
        out1 => S2867
    );
nand_n_1524: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2776,
        in1(1) => S2763,
        out1 => S2868
    );
nand_n_1525: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2868,
        in1(1) => S2867,
        out1 => S2869
    );
nor_n_943: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2869,
        in1(1) => S2866,
        out1 => S2735
    );
nand_n_1526: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_IMM1_out_14,
        in1(1) => CU_selIMM_PC,
        out1 => S2870
    );
nand_n_1527: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S2885,
        out1 => S2871
    );
nand_n_1528: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2871,
        in1(1) => S2870,
        out1 => S2872
    );
nor_n_944: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2872,
        in1(1) => S2770,
        out1 => S2873
    );
nand_n_1529: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2766,
        in1(1) => CU_selINC_PC,
        out1 => S2874
    );
nand_n_1530: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2776,
        in1(1) => S2765,
        out1 => S2875
    );
nand_n_1531: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2875,
        in1(1) => S2874,
        out1 => S2876
    );
nor_n_945: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2876,
        in1(1) => S2873,
        out1 => S2736
    );
nand_n_1532: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S2885,
        out1 => S2877
    );
nand_n_1533: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_IMM1_out_15,
        in1(1) => CU_selIMM_PC,
        out1 => S2878
    );
nand_n_1534: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2878,
        in1(1) => S2877,
        out1 => S2879
    );
nor_n_946: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2879,
        in1(1) => S2770,
        out1 => S2880
    );
nand_n_1535: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2768,
        in1(1) => CU_selINC_PC,
        out1 => S2881
    );
nand_n_1536: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2776,
        in1(1) => S2767,
        out1 => S2882
    );
nand_n_1537: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2882,
        in1(1) => S2881,
        out1 => S2883
    );
nor_n_947: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2883,
        in1(1) => S2880,
        out1 => S2737
    );
nand_n_1538: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2769,
        in1(1) => S2885,
        out1 => S2884
    );
nor_n_948: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2884,
        in1(1) => S2770,
        out1 => S2747
    );
$_DLATCH_N__107: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2731,
        E => S2747,
        Q => DP_PC_in_0
    );
$_DLATCH_N__108: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2738,
        E => S2747,
        Q => DP_PC_in_1
    );
$_DLATCH_N__109: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2739,
        E => S2747,
        Q => DP_PC_in_2
    );
$_DLATCH_N__110: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2740,
        E => S2747,
        Q => DP_PC_in_3
    );
$_DLATCH_N__111: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2741,
        E => S2747,
        Q => DP_PC_in_4
    );
$_DLATCH_N__112: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2742,
        E => S2747,
        Q => DP_PC_in_5
    );
$_DLATCH_N__113: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2743,
        E => S2747,
        Q => DP_PC_in_6
    );
$_DLATCH_N__114: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2744,
        E => S2747,
        Q => DP_PC_in_7
    );
$_DLATCH_N__115: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2745,
        E => S2747,
        Q => DP_PC_in_8
    );
$_DLATCH_N__116: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2746,
        E => S2747,
        Q => DP_PC_in_9
    );
$_DLATCH_N__117: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2732,
        E => S2747,
        Q => DP_PC_in_10
    );
$_DLATCH_N__118: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2733,
        E => S2747,
        Q => DP_PC_in_11
    );
$_DLATCH_N__119: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2734,
        E => S2747,
        Q => DP_PC_in_12
    );
$_DLATCH_N__120: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2735,
        E => S2747,
        Q => DP_PC_in_13
    );
$_DLATCH_N__121: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2736,
        E => S2747,
        Q => DP_PC_in_14
    );
$_DLATCH_N__122: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2737,
        E => S2747,
        Q => DP_PC_in_15
    );
notg_442: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_selINC_IN,
        out1 => S2916
    );
nand_n_1539: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_selINC_IN,
        in1(1) => DP_INC2_out_0,
        out1 => S2917
    );
nand_n_1540: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2916,
        in1(1) => dataBus(0),
        out1 => S2918
    );
nand_n_1541: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2918,
        in1(1) => S2917,
        out1 => S2899
    );
nand_n_1542: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_INC2_out_1,
        in1(1) => CU_selINC_IN,
        out1 => S2919
    );
nand_n_1543: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => dataBus(1),
        in1(1) => S2916,
        out1 => S2920
    );
nand_n_1544: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2920,
        in1(1) => S2919,
        out1 => S2906
    );
nand_n_1545: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_INC2_out_2,
        in1(1) => CU_selINC_IN,
        out1 => S2921
    );
nand_n_1546: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => dataBus(2),
        in1(1) => S2916,
        out1 => S2922
    );
nand_n_1547: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2922,
        in1(1) => S2921,
        out1 => S2907
    );
nand_n_1548: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_INC2_out_3,
        in1(1) => CU_selINC_IN,
        out1 => S2923
    );
nand_n_1549: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => dataBus(3),
        in1(1) => S2916,
        out1 => S2924
    );
nand_n_1550: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2924,
        in1(1) => S2923,
        out1 => S2908
    );
nand_n_1551: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_INC2_out_4,
        in1(1) => CU_selINC_IN,
        out1 => S2925
    );
nand_n_1552: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => dataBus(4),
        in1(1) => S2916,
        out1 => S2926
    );
nand_n_1553: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2926,
        in1(1) => S2925,
        out1 => S2909
    );
nand_n_1554: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_INC2_out_5,
        in1(1) => CU_selINC_IN,
        out1 => S2927
    );
nand_n_1555: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => dataBus(5),
        in1(1) => S2916,
        out1 => S2928
    );
nand_n_1556: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2928,
        in1(1) => S2927,
        out1 => S2910
    );
nand_n_1557: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_INC2_out_6,
        in1(1) => CU_selINC_IN,
        out1 => S2929
    );
nand_n_1558: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => dataBus(6),
        in1(1) => S2916,
        out1 => S2930
    );
nand_n_1559: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2930,
        in1(1) => S2929,
        out1 => S2911
    );
nand_n_1560: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_INC2_out_7,
        in1(1) => CU_selINC_IN,
        out1 => S2931
    );
nand_n_1561: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => dataBus(7),
        in1(1) => S2916,
        out1 => S2932
    );
nand_n_1562: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2932,
        in1(1) => S2931,
        out1 => S2912
    );
nand_n_1563: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_INC2_out_8,
        in1(1) => CU_selINC_IN,
        out1 => S2933
    );
nand_n_1564: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => dataBus(8),
        in1(1) => S2916,
        out1 => S2934
    );
nand_n_1565: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2934,
        in1(1) => S2933,
        out1 => S2913
    );
nand_n_1566: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_INC2_out_9,
        in1(1) => CU_selINC_IN,
        out1 => S2935
    );
nand_n_1567: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => dataBus(9),
        in1(1) => S2916,
        out1 => S2936
    );
nand_n_1568: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2936,
        in1(1) => S2935,
        out1 => S2914
    );
nand_n_1569: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_INC2_out_10,
        in1(1) => CU_selINC_IN,
        out1 => S2937
    );
nand_n_1570: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => dataBus(10),
        in1(1) => S2916,
        out1 => S2938
    );
nand_n_1571: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2938,
        in1(1) => S2937,
        out1 => S2900
    );
nand_n_1572: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_INC2_out_11,
        in1(1) => CU_selINC_IN,
        out1 => S2939
    );
nand_n_1573: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => dataBus(11),
        in1(1) => S2916,
        out1 => S2940
    );
nand_n_1574: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2940,
        in1(1) => S2939,
        out1 => S2901
    );
nand_n_1575: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_INC2_out_12,
        in1(1) => CU_selINC_IN,
        out1 => S2941
    );
nand_n_1576: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => dataBus(12),
        in1(1) => S2916,
        out1 => S2942
    );
nand_n_1577: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2942,
        in1(1) => S2941,
        out1 => S2902
    );
nand_n_1578: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_INC2_out_13,
        in1(1) => CU_selINC_IN,
        out1 => S2943
    );
nand_n_1579: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => dataBus(13),
        in1(1) => S2916,
        out1 => S2944
    );
nand_n_1580: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2944,
        in1(1) => S2943,
        out1 => S2903
    );
nand_n_1581: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_INC2_out_14,
        in1(1) => CU_selINC_IN,
        out1 => S2945
    );
nand_n_1582: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => dataBus(14),
        in1(1) => S2916,
        out1 => S2946
    );
nand_n_1583: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2946,
        in1(1) => S2945,
        out1 => S2904
    );
nand_n_1584: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_INC2_out_15,
        in1(1) => CU_selINC_IN,
        out1 => S2947
    );
nand_n_1585: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => dataBus(15),
        in1(1) => S2916,
        out1 => S2948
    );
nand_n_1586: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2948,
        in1(1) => S2947,
        out1 => S2905
    );
nor_n_949: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => CU_selMEM_IN,
        in1(1) => CU_selINC_IN,
        out1 => S2915
    );
$_DLATCH_N__123: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2899,
        E => S2915,
        Q => DP_IN_in_0
    );
$_DLATCH_N__124: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2906,
        E => S2915,
        Q => DP_IN_in_1
    );
$_DLATCH_N__125: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2907,
        E => S2915,
        Q => DP_IN_in_2
    );
$_DLATCH_N__126: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2908,
        E => S2915,
        Q => DP_IN_in_3
    );
$_DLATCH_N__127: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2909,
        E => S2915,
        Q => DP_IN_in_4
    );
$_DLATCH_N__128: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2910,
        E => S2915,
        Q => DP_IN_in_5
    );
$_DLATCH_N__129: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2911,
        E => S2915,
        Q => DP_IN_in_6
    );
$_DLATCH_N__130: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2912,
        E => S2915,
        Q => DP_IN_in_7
    );
$_DLATCH_N__131: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2913,
        E => S2915,
        Q => DP_IN_in_8
    );
$_DLATCH_N__132: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2914,
        E => S2915,
        Q => DP_IN_in_9
    );
$_DLATCH_N__133: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2900,
        E => S2915,
        Q => DP_IN_in_10
    );
$_DLATCH_N__134: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2901,
        E => S2915,
        Q => DP_IN_in_11
    );
$_DLATCH_N__135: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2902,
        E => S2915,
        Q => DP_IN_in_12
    );
$_DLATCH_N__136: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2903,
        E => S2915,
        Q => DP_IN_in_13
    );
$_DLATCH_N__137: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2904,
        E => S2915,
        Q => DP_IN_in_14
    );
$_DLATCH_N__138: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2905,
        E => S2915,
        Q => DP_IN_in_15
    );
notg_443: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_selAC_MEM,
        out1 => S3103
    );
notg_444: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_out_0,
        out1 => S3104
    );
notg_445: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_selPC_MEM,
        out1 => S3105
    );
notg_446: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IN_out_0,
        out1 => S3106
    );
notg_447: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_selIN_MEM,
        out1 => S3107
    );
notg_448: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_out_1,
        out1 => S3108
    );
notg_449: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IN_out_1,
        out1 => S3109
    );
notg_450: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_out_2,
        out1 => S3110
    );
notg_451: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IN_out_2,
        out1 => S3111
    );
notg_452: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_out_3,
        out1 => S3112
    );
notg_453: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IN_out_3,
        out1 => S3113
    );
notg_454: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_out_4,
        out1 => S3114
    );
notg_455: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IN_out_4,
        out1 => S3115
    );
notg_456: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_out_5,
        out1 => S3116
    );
notg_457: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IN_out_5,
        out1 => S2966
    );
notg_458: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_out_6,
        out1 => S2967
    );
notg_459: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IN_out_6,
        out1 => S2968
    );
notg_460: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_out_7,
        out1 => S2969
    );
notg_461: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IN_out_7,
        out1 => S2970
    );
notg_462: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_out_8,
        out1 => S2971
    );
notg_463: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IN_out_8,
        out1 => S2972
    );
notg_464: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_out_9,
        out1 => S2973
    );
notg_465: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IN_out_9,
        out1 => S2974
    );
notg_466: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_out_10,
        out1 => S2975
    );
notg_467: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IN_out_10,
        out1 => S2976
    );
notg_468: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_out_11,
        out1 => S2977
    );
notg_469: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IN_out_11,
        out1 => S2978
    );
notg_470: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_out_12,
        out1 => S2979
    );
notg_471: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IN_out_12,
        out1 => S2980
    );
notg_472: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_out_13,
        out1 => S2981
    );
notg_473: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IN_out_13,
        out1 => S2982
    );
notg_474: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_out_14,
        out1 => S2983
    );
notg_475: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IN_out_14,
        out1 => S2984
    );
notg_476: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_INC_1_out_15,
        out1 => S2985
    );
notg_477: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IN_out_15,
        out1 => S2986
    );
notg_478: ENTITY WORK.notg
    PORT MAP (
        in1 => 'z',
        out1 => S2987
    );
nand_n_1587: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3107,
        in1(1) => S3105,
        out1 => S2988
    );
nand_n_1588: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_selAC_MEM,
        in1(1) => DP_AC_out_0,
        out1 => S2989
    );
nand_n_1589: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3103,
        in1(1) => 'z',
        out1 => S2990
    );
nand_n_1590: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2990,
        in1(1) => S2989,
        out1 => S2991
    );
nor_n_950: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2991,
        in1(1) => S2988,
        out1 => S2992
    );
nand_n_1591: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_selIN_MEM,
        in1(1) => S3106,
        out1 => S2993
    );
nor_n_951: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => CU_selIN_MEM,
        in1(1) => S3105,
        out1 => S2994
    );
nand_n_1592: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2994,
        in1(1) => S3104,
        out1 => S2995
    );
nand_n_1593: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2995,
        in1(1) => S2993,
        out1 => S2996
    );
nor_n_952: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2996,
        in1(1) => S2992,
        out1 => S2949
    );
nand_n_1594: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S3103,
        out1 => S2997
    );
nand_n_1595: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_1,
        in1(1) => CU_selAC_MEM,
        out1 => S2998
    );
nand_n_1596: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2998,
        in1(1) => S2997,
        out1 => S2999
    );
nor_n_953: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2999,
        in1(1) => S2988,
        out1 => S3000
    );
nand_n_1597: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3109,
        in1(1) => CU_selIN_MEM,
        out1 => S3001
    );
nand_n_1598: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2994,
        in1(1) => S3108,
        out1 => S3002
    );
nand_n_1599: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3002,
        in1(1) => S3001,
        out1 => S3003
    );
nor_n_954: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3003,
        in1(1) => S3000,
        out1 => S2956
    );
nand_n_1600: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S3103,
        out1 => S3004
    );
nand_n_1601: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_2,
        in1(1) => CU_selAC_MEM,
        out1 => S3005
    );
nand_n_1602: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3005,
        in1(1) => S3004,
        out1 => S3006
    );
nor_n_955: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3006,
        in1(1) => S2988,
        out1 => S3007
    );
nand_n_1603: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3111,
        in1(1) => CU_selIN_MEM,
        out1 => S3008
    );
nand_n_1604: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2994,
        in1(1) => S3110,
        out1 => S3009
    );
nand_n_1605: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3009,
        in1(1) => S3008,
        out1 => S3010
    );
nor_n_956: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3010,
        in1(1) => S3007,
        out1 => S2957
    );
nand_n_1606: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S3103,
        out1 => S3011
    );
nand_n_1607: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_3,
        in1(1) => CU_selAC_MEM,
        out1 => S3012
    );
nand_n_1608: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3012,
        in1(1) => S3011,
        out1 => S3013
    );
nor_n_957: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3013,
        in1(1) => S2988,
        out1 => S3014
    );
nand_n_1609: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3113,
        in1(1) => CU_selIN_MEM,
        out1 => S3015
    );
nand_n_1610: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2994,
        in1(1) => S3112,
        out1 => S3016
    );
nand_n_1611: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3016,
        in1(1) => S3015,
        out1 => S3017
    );
nor_n_958: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3017,
        in1(1) => S3014,
        out1 => S2958
    );
nand_n_1612: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S3103,
        out1 => S3018
    );
nand_n_1613: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_4,
        in1(1) => CU_selAC_MEM,
        out1 => S3019
    );
nand_n_1614: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3019,
        in1(1) => S3018,
        out1 => S3020
    );
nor_n_959: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3020,
        in1(1) => S2988,
        out1 => S3021
    );
nand_n_1615: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3115,
        in1(1) => CU_selIN_MEM,
        out1 => S3022
    );
nand_n_1616: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2994,
        in1(1) => S3114,
        out1 => S3023
    );
nand_n_1617: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3023,
        in1(1) => S3022,
        out1 => S3024
    );
nor_n_960: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3024,
        in1(1) => S3021,
        out1 => S2959
    );
nand_n_1618: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S3103,
        out1 => S3025
    );
nand_n_1619: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_5,
        in1(1) => CU_selAC_MEM,
        out1 => S3026
    );
nand_n_1620: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3026,
        in1(1) => S3025,
        out1 => S3027
    );
nor_n_961: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3027,
        in1(1) => S2988,
        out1 => S3028
    );
nand_n_1621: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2966,
        in1(1) => CU_selIN_MEM,
        out1 => S3029
    );
nand_n_1622: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2994,
        in1(1) => S3116,
        out1 => S3030
    );
nand_n_1623: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3030,
        in1(1) => S3029,
        out1 => S3031
    );
nor_n_962: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3031,
        in1(1) => S3028,
        out1 => S2960
    );
nand_n_1624: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S3103,
        out1 => S3032
    );
nand_n_1625: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_6,
        in1(1) => CU_selAC_MEM,
        out1 => S3033
    );
nand_n_1626: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3033,
        in1(1) => S3032,
        out1 => S3034
    );
nor_n_963: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3034,
        in1(1) => S2988,
        out1 => S3035
    );
nand_n_1627: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2968,
        in1(1) => CU_selIN_MEM,
        out1 => S3036
    );
nand_n_1628: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2994,
        in1(1) => S2967,
        out1 => S3037
    );
nand_n_1629: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3037,
        in1(1) => S3036,
        out1 => S3038
    );
nor_n_964: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3038,
        in1(1) => S3035,
        out1 => S2961
    );
nand_n_1630: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S3103,
        out1 => S3039
    );
nand_n_1631: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_7,
        in1(1) => CU_selAC_MEM,
        out1 => S3040
    );
nand_n_1632: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3040,
        in1(1) => S3039,
        out1 => S3041
    );
nor_n_965: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3041,
        in1(1) => S2988,
        out1 => S3042
    );
nand_n_1633: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2970,
        in1(1) => CU_selIN_MEM,
        out1 => S3043
    );
nand_n_1634: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2994,
        in1(1) => S2969,
        out1 => S3044
    );
nand_n_1635: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3044,
        in1(1) => S3043,
        out1 => S3045
    );
nor_n_966: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3045,
        in1(1) => S3042,
        out1 => S2962
    );
nand_n_1636: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_8,
        in1(1) => CU_selAC_MEM,
        out1 => S3046
    );
nand_n_1637: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S3103,
        out1 => S3047
    );
nand_n_1638: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3047,
        in1(1) => S3046,
        out1 => S3048
    );
nor_n_967: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3048,
        in1(1) => S2988,
        out1 => S3049
    );
nand_n_1639: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2972,
        in1(1) => CU_selIN_MEM,
        out1 => S3050
    );
nand_n_1640: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2994,
        in1(1) => S2971,
        out1 => S3051
    );
nand_n_1641: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3051,
        in1(1) => S3050,
        out1 => S3052
    );
nor_n_968: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3052,
        in1(1) => S3049,
        out1 => S2963
    );
nand_n_1642: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S3103,
        out1 => S3053
    );
nand_n_1643: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_9,
        in1(1) => CU_selAC_MEM,
        out1 => S3054
    );
nand_n_1644: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3054,
        in1(1) => S3053,
        out1 => S3055
    );
nor_n_969: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3055,
        in1(1) => S2988,
        out1 => S3056
    );
nand_n_1645: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2974,
        in1(1) => CU_selIN_MEM,
        out1 => S3057
    );
nand_n_1646: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2994,
        in1(1) => S2973,
        out1 => S3058
    );
nand_n_1647: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3058,
        in1(1) => S3057,
        out1 => S3059
    );
nor_n_970: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3059,
        in1(1) => S3056,
        out1 => S2964
    );
nand_n_1648: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_10,
        in1(1) => CU_selAC_MEM,
        out1 => S3060
    );
nand_n_1649: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S3103,
        out1 => S3061
    );
nand_n_1650: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3061,
        in1(1) => S3060,
        out1 => S3062
    );
nor_n_971: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3062,
        in1(1) => S2988,
        out1 => S3063
    );
nand_n_1651: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2976,
        in1(1) => CU_selIN_MEM,
        out1 => S3064
    );
nand_n_1652: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2994,
        in1(1) => S2975,
        out1 => S3065
    );
nand_n_1653: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3065,
        in1(1) => S3064,
        out1 => S3066
    );
nor_n_972: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3066,
        in1(1) => S3063,
        out1 => S2950
    );
nand_n_1654: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S3103,
        out1 => S3067
    );
nand_n_1655: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_11,
        in1(1) => CU_selAC_MEM,
        out1 => S3068
    );
nand_n_1656: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3068,
        in1(1) => S3067,
        out1 => S3069
    );
nor_n_973: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3069,
        in1(1) => S2988,
        out1 => S3070
    );
nand_n_1657: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2978,
        in1(1) => CU_selIN_MEM,
        out1 => S3071
    );
nand_n_1658: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2994,
        in1(1) => S2977,
        out1 => S3072
    );
nand_n_1659: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3072,
        in1(1) => S3071,
        out1 => S3073
    );
nor_n_974: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3073,
        in1(1) => S3070,
        out1 => S2951
    );
nand_n_1660: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_12,
        in1(1) => CU_selAC_MEM,
        out1 => S3074
    );
nand_n_1661: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S3103,
        out1 => S3075
    );
nand_n_1662: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3075,
        in1(1) => S3074,
        out1 => S3076
    );
nor_n_975: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3076,
        in1(1) => S2988,
        out1 => S3077
    );
nand_n_1663: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2980,
        in1(1) => CU_selIN_MEM,
        out1 => S3078
    );
nand_n_1664: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2994,
        in1(1) => S2979,
        out1 => S3079
    );
nand_n_1665: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3079,
        in1(1) => S3078,
        out1 => S3080
    );
nor_n_976: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3080,
        in1(1) => S3077,
        out1 => S2952
    );
nand_n_1666: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S3103,
        out1 => S3081
    );
nand_n_1667: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_13,
        in1(1) => CU_selAC_MEM,
        out1 => S3082
    );
nand_n_1668: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3082,
        in1(1) => S3081,
        out1 => S3083
    );
nor_n_977: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3083,
        in1(1) => S2988,
        out1 => S3084
    );
nand_n_1669: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2982,
        in1(1) => CU_selIN_MEM,
        out1 => S3085
    );
nand_n_1670: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2994,
        in1(1) => S2981,
        out1 => S3086
    );
nand_n_1671: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3086,
        in1(1) => S3085,
        out1 => S3087
    );
nor_n_978: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3087,
        in1(1) => S3084,
        out1 => S2953
    );
nand_n_1672: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_14,
        in1(1) => CU_selAC_MEM,
        out1 => S3088
    );
nand_n_1673: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S3103,
        out1 => S3089
    );
nand_n_1674: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3089,
        in1(1) => S3088,
        out1 => S3090
    );
nor_n_979: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3090,
        in1(1) => S2988,
        out1 => S3091
    );
nand_n_1675: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2984,
        in1(1) => CU_selIN_MEM,
        out1 => S3092
    );
nand_n_1676: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2994,
        in1(1) => S2983,
        out1 => S3093
    );
nand_n_1677: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3093,
        in1(1) => S3092,
        out1 => S3094
    );
nor_n_980: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3094,
        in1(1) => S3091,
        out1 => S2954
    );
nand_n_1678: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S3103,
        out1 => S3095
    );
nand_n_1679: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_AC_out_15,
        in1(1) => CU_selAC_MEM,
        out1 => S3096
    );
nand_n_1680: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3096,
        in1(1) => S3095,
        out1 => S3097
    );
nor_n_981: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3097,
        in1(1) => S2988,
        out1 => S3098
    );
nand_n_1681: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2986,
        in1(1) => CU_selIN_MEM,
        out1 => S3099
    );
nand_n_1682: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2994,
        in1(1) => S2985,
        out1 => S3100
    );
nand_n_1683: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3100,
        in1(1) => S3099,
        out1 => S3101
    );
nor_n_982: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3101,
        in1(1) => S3098,
        out1 => S2955
    );
nand_n_1684: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2987,
        in1(1) => S3103,
        out1 => S3102
    );
nor_n_983: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3102,
        in1(1) => S2988,
        out1 => S2965
    );
$_DLATCH_N__139: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2949,
        E => S2965,
        Q => dataBus(0)
    );
$_DLATCH_N__140: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2956,
        E => S2965,
        Q => dataBus(1)
    );
$_DLATCH_N__141: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2957,
        E => S2965,
        Q => dataBus(2)
    );
$_DLATCH_N__142: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2958,
        E => S2965,
        Q => dataBus(3)
    );
$_DLATCH_N__143: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2959,
        E => S2965,
        Q => dataBus(4)
    );
$_DLATCH_N__144: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2960,
        E => S2965,
        Q => dataBus(5)
    );
$_DLATCH_N__145: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2961,
        E => S2965,
        Q => dataBus(6)
    );
$_DLATCH_N__146: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2962,
        E => S2965,
        Q => dataBus(7)
    );
$_DLATCH_N__147: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2963,
        E => S2965,
        Q => dataBus(8)
    );
$_DLATCH_N__148: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2964,
        E => S2965,
        Q => dataBus(9)
    );
$_DLATCH_N__149: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2950,
        E => S2965,
        Q => dataBus(10)
    );
$_DLATCH_N__150: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2951,
        E => S2965,
        Q => dataBus(11)
    );
$_DLATCH_N__151: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2952,
        E => S2965,
        Q => dataBus(12)
    );
$_DLATCH_N__152: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2953,
        E => S2965,
        Q => dataBus(13)
    );
$_DLATCH_N__153: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2954,
        E => S2965,
        Q => dataBus(14)
    );
$_DLATCH_N__154: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S2955,
        E => S2965,
        Q => dataBus(15)
    );
notg_479: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_ldIR,
        out1 => S3271
    );
notg_480: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IMM1_out_0,
        out1 => S3272
    );
notg_481: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_selIR_ADR,
        out1 => S3273
    );
notg_482: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IN_out_0,
        out1 => S3274
    );
notg_483: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_selIN_ADR,
        out1 => S3275
    );
notg_484: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IMM1_out_1,
        out1 => S3276
    );
notg_485: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IN_out_1,
        out1 => S3277
    );
notg_486: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IMM1_out_2,
        out1 => S3278
    );
notg_487: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IN_out_2,
        out1 => S3279
    );
notg_488: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IMM1_out_3,
        out1 => S3280
    );
notg_489: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IN_out_3,
        out1 => S3281
    );
notg_490: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IMM1_out_4,
        out1 => S3282
    );
notg_491: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IN_out_4,
        out1 => S3283
    );
notg_492: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IMM1_out_5,
        out1 => S3284
    );
notg_493: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IN_out_5,
        out1 => S3134
    );
notg_494: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IMM1_out_6,
        out1 => S3135
    );
notg_495: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IN_out_6,
        out1 => S3136
    );
notg_496: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IMM1_out_7,
        out1 => S3137
    );
notg_497: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IN_out_7,
        out1 => S3138
    );
notg_498: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IMM1_out_8,
        out1 => S3139
    );
notg_499: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IN_out_8,
        out1 => S3140
    );
notg_500: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IMM1_out_9,
        out1 => S3141
    );
notg_501: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IN_out_9,
        out1 => S3142
    );
notg_502: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IMM1_out_10,
        out1 => S3143
    );
notg_503: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IN_out_10,
        out1 => S3144
    );
notg_504: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IMM1_out_11,
        out1 => S3145
    );
notg_505: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IN_out_11,
        out1 => S3146
    );
notg_506: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IMM1_out_12,
        out1 => S3147
    );
notg_507: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IN_out_12,
        out1 => S3148
    );
notg_508: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IMM1_out_13,
        out1 => S3149
    );
notg_509: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IN_out_13,
        out1 => S3150
    );
notg_510: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IMM1_out_14,
        out1 => S3151
    );
notg_511: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IN_out_14,
        out1 => S3152
    );
notg_512: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IMM1_out_15,
        out1 => S3153
    );
notg_513: ENTITY WORK.notg
    PORT MAP (
        in1 => DP_IN_out_15,
        out1 => S3154
    );
notg_514: ENTITY WORK.notg
    PORT MAP (
        in1 => 'z',
        out1 => S3155
    );
nand_n_1685: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3275,
        in1(1) => S3273,
        out1 => S3156
    );
nand_n_1686: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_ldIR,
        in1(1) => DP_INC_1_in_0,
        out1 => S3157
    );
nand_n_1687: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3271,
        in1(1) => 'z',
        out1 => S3158
    );
nand_n_1688: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3158,
        in1(1) => S3157,
        out1 => S3159
    );
nor_n_984: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3159,
        in1(1) => S3156,
        out1 => S3160
    );
nand_n_1689: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_selIN_ADR,
        in1(1) => S3274,
        out1 => S3161
    );
nor_n_985: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => CU_selIN_ADR,
        in1(1) => S3273,
        out1 => S3162
    );
nand_n_1690: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3162,
        in1(1) => S3272,
        out1 => S3163
    );
nand_n_1691: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3163,
        in1(1) => S3161,
        out1 => S3164
    );
nor_n_986: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3164,
        in1(1) => S3160,
        out1 => S3117
    );
nand_n_1692: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S3271,
        out1 => S3165
    );
nand_n_1693: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_INC_1_in_1,
        in1(1) => CU_ldIR,
        out1 => S3166
    );
nand_n_1694: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3166,
        in1(1) => S3165,
        out1 => S3167
    );
nor_n_987: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3167,
        in1(1) => S3156,
        out1 => S3168
    );
nand_n_1695: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3277,
        in1(1) => CU_selIN_ADR,
        out1 => S3169
    );
nand_n_1696: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3162,
        in1(1) => S3276,
        out1 => S3170
    );
nand_n_1697: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3170,
        in1(1) => S3169,
        out1 => S3171
    );
nor_n_988: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3171,
        in1(1) => S3168,
        out1 => S3124
    );
nand_n_1698: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S3271,
        out1 => S3172
    );
nand_n_1699: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_INC_1_in_2,
        in1(1) => CU_ldIR,
        out1 => S3173
    );
nand_n_1700: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3173,
        in1(1) => S3172,
        out1 => S3174
    );
nor_n_989: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3174,
        in1(1) => S3156,
        out1 => S3175
    );
nand_n_1701: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3279,
        in1(1) => CU_selIN_ADR,
        out1 => S3176
    );
nand_n_1702: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3162,
        in1(1) => S3278,
        out1 => S3177
    );
nand_n_1703: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3177,
        in1(1) => S3176,
        out1 => S3178
    );
nor_n_990: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3178,
        in1(1) => S3175,
        out1 => S3125
    );
nand_n_1704: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S3271,
        out1 => S3179
    );
nand_n_1705: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_INC_1_in_3,
        in1(1) => CU_ldIR,
        out1 => S3180
    );
nand_n_1706: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3180,
        in1(1) => S3179,
        out1 => S3181
    );
nor_n_991: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3181,
        in1(1) => S3156,
        out1 => S3182
    );
nand_n_1707: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3281,
        in1(1) => CU_selIN_ADR,
        out1 => S3183
    );
nand_n_1708: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3162,
        in1(1) => S3280,
        out1 => S3184
    );
nand_n_1709: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3184,
        in1(1) => S3183,
        out1 => S3185
    );
nor_n_992: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3185,
        in1(1) => S3182,
        out1 => S3126
    );
nand_n_1710: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S3271,
        out1 => S3186
    );
nand_n_1711: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_INC_1_in_4,
        in1(1) => CU_ldIR,
        out1 => S3187
    );
nand_n_1712: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3187,
        in1(1) => S3186,
        out1 => S3188
    );
nor_n_993: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3188,
        in1(1) => S3156,
        out1 => S3189
    );
nand_n_1713: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3283,
        in1(1) => CU_selIN_ADR,
        out1 => S3190
    );
nand_n_1714: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3162,
        in1(1) => S3282,
        out1 => S3191
    );
nand_n_1715: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3191,
        in1(1) => S3190,
        out1 => S3192
    );
nor_n_994: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3192,
        in1(1) => S3189,
        out1 => S3127
    );
nand_n_1716: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S3271,
        out1 => S3193
    );
nand_n_1717: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_INC_1_in_5,
        in1(1) => CU_ldIR,
        out1 => S3194
    );
nand_n_1718: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3194,
        in1(1) => S3193,
        out1 => S3195
    );
nor_n_995: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3195,
        in1(1) => S3156,
        out1 => S3196
    );
nand_n_1719: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3134,
        in1(1) => CU_selIN_ADR,
        out1 => S3197
    );
nand_n_1720: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3162,
        in1(1) => S3284,
        out1 => S3198
    );
nand_n_1721: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3198,
        in1(1) => S3197,
        out1 => S3199
    );
nor_n_996: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3199,
        in1(1) => S3196,
        out1 => S3128
    );
nand_n_1722: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S3271,
        out1 => S3200
    );
nand_n_1723: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_INC_1_in_6,
        in1(1) => CU_ldIR,
        out1 => S3201
    );
nand_n_1724: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3201,
        in1(1) => S3200,
        out1 => S3202
    );
nor_n_997: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3202,
        in1(1) => S3156,
        out1 => S3203
    );
nand_n_1725: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3136,
        in1(1) => CU_selIN_ADR,
        out1 => S3204
    );
nand_n_1726: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3162,
        in1(1) => S3135,
        out1 => S3205
    );
nand_n_1727: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3205,
        in1(1) => S3204,
        out1 => S3206
    );
nor_n_998: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3206,
        in1(1) => S3203,
        out1 => S3129
    );
nand_n_1728: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S3271,
        out1 => S3207
    );
nand_n_1729: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_INC_1_in_7,
        in1(1) => CU_ldIR,
        out1 => S3208
    );
nand_n_1730: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3208,
        in1(1) => S3207,
        out1 => S3209
    );
nor_n_999: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3209,
        in1(1) => S3156,
        out1 => S3210
    );
nand_n_1731: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3138,
        in1(1) => CU_selIN_ADR,
        out1 => S3211
    );
nand_n_1732: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3162,
        in1(1) => S3137,
        out1 => S3212
    );
nand_n_1733: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3212,
        in1(1) => S3211,
        out1 => S3213
    );
nor_n_1000: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3213,
        in1(1) => S3210,
        out1 => S3130
    );
nand_n_1734: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_INC_1_in_8,
        in1(1) => CU_ldIR,
        out1 => S3214
    );
nand_n_1735: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S3271,
        out1 => S3215
    );
nand_n_1736: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3215,
        in1(1) => S3214,
        out1 => S3216
    );
nor_n_1001: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3216,
        in1(1) => S3156,
        out1 => S3217
    );
nand_n_1737: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3140,
        in1(1) => CU_selIN_ADR,
        out1 => S3218
    );
nand_n_1738: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3162,
        in1(1) => S3139,
        out1 => S3219
    );
nand_n_1739: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3219,
        in1(1) => S3218,
        out1 => S3220
    );
nor_n_1002: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3220,
        in1(1) => S3217,
        out1 => S3131
    );
nand_n_1740: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S3271,
        out1 => S3221
    );
nand_n_1741: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_INC_1_in_9,
        in1(1) => CU_ldIR,
        out1 => S3222
    );
nand_n_1742: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3222,
        in1(1) => S3221,
        out1 => S3223
    );
nor_n_1003: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3223,
        in1(1) => S3156,
        out1 => S3224
    );
nand_n_1743: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3142,
        in1(1) => CU_selIN_ADR,
        out1 => S3225
    );
nand_n_1744: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3162,
        in1(1) => S3141,
        out1 => S3226
    );
nand_n_1745: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3226,
        in1(1) => S3225,
        out1 => S3227
    );
nor_n_1004: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3227,
        in1(1) => S3224,
        out1 => S3132
    );
nand_n_1746: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_INC_1_in_10,
        in1(1) => CU_ldIR,
        out1 => S3228
    );
nand_n_1747: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S3271,
        out1 => S3229
    );
nand_n_1748: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3229,
        in1(1) => S3228,
        out1 => S3230
    );
nor_n_1005: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3230,
        in1(1) => S3156,
        out1 => S3231
    );
nand_n_1749: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3144,
        in1(1) => CU_selIN_ADR,
        out1 => S3232
    );
nand_n_1750: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3162,
        in1(1) => S3143,
        out1 => S3233
    );
nand_n_1751: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3233,
        in1(1) => S3232,
        out1 => S3234
    );
nor_n_1006: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3234,
        in1(1) => S3231,
        out1 => S3118
    );
nand_n_1752: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S3271,
        out1 => S3235
    );
nand_n_1753: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_INC_1_in_11,
        in1(1) => CU_ldIR,
        out1 => S3236
    );
nand_n_1754: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3236,
        in1(1) => S3235,
        out1 => S3237
    );
nor_n_1007: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3237,
        in1(1) => S3156,
        out1 => S3238
    );
nand_n_1755: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3146,
        in1(1) => CU_selIN_ADR,
        out1 => S3239
    );
nand_n_1756: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3162,
        in1(1) => S3145,
        out1 => S3240
    );
nand_n_1757: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3240,
        in1(1) => S3239,
        out1 => S3241
    );
nor_n_1008: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3241,
        in1(1) => S3238,
        out1 => S3119
    );
nand_n_1758: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_INC_1_in_12,
        in1(1) => CU_ldIR,
        out1 => S3242
    );
nand_n_1759: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S3271,
        out1 => S3243
    );
nand_n_1760: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3243,
        in1(1) => S3242,
        out1 => S3244
    );
nor_n_1009: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3244,
        in1(1) => S3156,
        out1 => S3245
    );
nand_n_1761: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3148,
        in1(1) => CU_selIN_ADR,
        out1 => S3246
    );
nand_n_1762: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3162,
        in1(1) => S3147,
        out1 => S3247
    );
nand_n_1763: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3247,
        in1(1) => S3246,
        out1 => S3248
    );
nor_n_1010: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3248,
        in1(1) => S3245,
        out1 => S3120
    );
nand_n_1764: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S3271,
        out1 => S3249
    );
nand_n_1765: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_INC_1_in_13,
        in1(1) => CU_ldIR,
        out1 => S3250
    );
nand_n_1766: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3250,
        in1(1) => S3249,
        out1 => S3251
    );
nor_n_1011: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3251,
        in1(1) => S3156,
        out1 => S3252
    );
nand_n_1767: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3150,
        in1(1) => CU_selIN_ADR,
        out1 => S3253
    );
nand_n_1768: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3162,
        in1(1) => S3149,
        out1 => S3254
    );
nand_n_1769: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3254,
        in1(1) => S3253,
        out1 => S3255
    );
nor_n_1012: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3255,
        in1(1) => S3252,
        out1 => S3121
    );
nand_n_1770: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_INC_1_in_14,
        in1(1) => CU_ldIR,
        out1 => S3256
    );
nand_n_1771: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S3271,
        out1 => S3257
    );
nand_n_1772: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3257,
        in1(1) => S3256,
        out1 => S3258
    );
nor_n_1013: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3258,
        in1(1) => S3156,
        out1 => S3259
    );
nand_n_1773: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3152,
        in1(1) => CU_selIN_ADR,
        out1 => S3260
    );
nand_n_1774: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3162,
        in1(1) => S3151,
        out1 => S3261
    );
nand_n_1775: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3261,
        in1(1) => S3260,
        out1 => S3262
    );
nor_n_1014: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3262,
        in1(1) => S3259,
        out1 => S3122
    );
nand_n_1776: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => 'z',
        in1(1) => S3271,
        out1 => S3263
    );
nand_n_1777: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => DP_INC_1_in_15,
        in1(1) => CU_ldIR,
        out1 => S3264
    );
nand_n_1778: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3264,
        in1(1) => S3263,
        out1 => S3265
    );
nor_n_1015: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3265,
        in1(1) => S3156,
        out1 => S3266
    );
nand_n_1779: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3154,
        in1(1) => CU_selIN_ADR,
        out1 => S3267
    );
nand_n_1780: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3162,
        in1(1) => S3153,
        out1 => S3268
    );
nand_n_1781: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3268,
        in1(1) => S3267,
        out1 => S3269
    );
nor_n_1016: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3269,
        in1(1) => S3266,
        out1 => S3123
    );
nand_n_1782: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3155,
        in1(1) => S3271,
        out1 => S3270
    );
nor_n_1017: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3270,
        in1(1) => S3156,
        out1 => S3133
    );
$_DLATCH_N__155: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S3117,
        E => S3133,
        Q => DP_addrBus_0
    );
$_DLATCH_N__156: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S3124,
        E => S3133,
        Q => DP_addrBus_1
    );
$_DLATCH_N__157: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S3125,
        E => S3133,
        Q => DP_addrBus_2
    );
$_DLATCH_N__158: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S3126,
        E => S3133,
        Q => DP_addrBus_3
    );
$_DLATCH_N__159: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S3127,
        E => S3133,
        Q => DP_addrBus_4
    );
$_DLATCH_N__160: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S3128,
        E => S3133,
        Q => DP_addrBus_5
    );
$_DLATCH_N__161: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S3129,
        E => S3133,
        Q => DP_addrBus_6
    );
$_DLATCH_N__162: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S3130,
        E => S3133,
        Q => DP_addrBus_7
    );
$_DLATCH_N__163: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S3131,
        E => S3133,
        Q => DP_addrBus_8
    );
$_DLATCH_N__164: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S3132,
        E => S3133,
        Q => DP_addrBus_9
    );
$_DLATCH_N__165: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S3118,
        E => S3133,
        Q => DP_addrBus_10
    );
$_DLATCH_N__166: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S3119,
        E => S3133,
        Q => DP_addrBus_11
    );
$_DLATCH_N__167: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S3120,
        E => S3133,
        Q => DP_addrBus_12
    );
$_DLATCH_N__168: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S3121,
        E => S3133,
        Q => DP_addrBus_13
    );
$_DLATCH_N__169: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S3122,
        E => S3133,
        Q => DP_addrBus_14
    );
$_DLATCH_N__170: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S3123,
        E => S3133,
        Q => DP_addrBus_15
    );
notg_515: ENTITY WORK.notg
    PORT MAP (
        in1 => CU_INC2,
        out1 => S3288
    );
nand_n_1783: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => CU_INC2,
        in1(1) => S36,
        out1 => S3289
    );
nand_n_1784: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3288,
        in1(1) => S4,
        out1 => S3290
    );
nand_n_1785: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3290,
        in1(1) => S3289,
        out1 => S3285
    );
nand_n_1786: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5,
        in1(1) => CU_INC2,
        out1 => S3291
    );
nand_n_1787: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S37,
        in1(1) => S3288,
        out1 => S3292
    );
nand_n_1788: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3292,
        in1(1) => S3291,
        out1 => S3286
    );
nor_n_1018: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => CU_INC1,
        in1(1) => CU_INC2,
        out1 => S3287
    );
$_DLATCH_N__171: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S3285,
        E => S3287,
        Q => DP_INC_1_inc_val_0
    );
$_DLATCH_N__172: ENTITY WORK.$_DLATCH_N_
    PORT MAP (
        D => S3286,
        E => S3287,
        Q => DP_INC_1_inc_val_1
    );
bufg_39: ENTITY WORK.bufg
    PORT MAP (
        in1 => DP_addrBus_0,
        out1 => addrBus(0)
    );
bufg_40: ENTITY WORK.bufg
    PORT MAP (
        in1 => DP_addrBus_1,
        out1 => addrBus(1)
    );
bufg_41: ENTITY WORK.bufg
    PORT MAP (
        in1 => DP_addrBus_10,
        out1 => addrBus(10)
    );
bufg_42: ENTITY WORK.bufg
    PORT MAP (
        in1 => DP_addrBus_11,
        out1 => addrBus(11)
    );
bufg_43: ENTITY WORK.bufg
    PORT MAP (
        in1 => DP_addrBus_12,
        out1 => addrBus(12)
    );
bufg_44: ENTITY WORK.bufg
    PORT MAP (
        in1 => DP_addrBus_13,
        out1 => addrBus(13)
    );
bufg_45: ENTITY WORK.bufg
    PORT MAP (
        in1 => DP_addrBus_14,
        out1 => addrBus(14)
    );
bufg_46: ENTITY WORK.bufg
    PORT MAP (
        in1 => DP_addrBus_15,
        out1 => addrBus(15)
    );
bufg_47: ENTITY WORK.bufg
    PORT MAP (
        in1 => DP_addrBus_2,
        out1 => addrBus(2)
    );
bufg_48: ENTITY WORK.bufg
    PORT MAP (
        in1 => DP_addrBus_3,
        out1 => addrBus(3)
    );
bufg_49: ENTITY WORK.bufg
    PORT MAP (
        in1 => DP_addrBus_4,
        out1 => addrBus(4)
    );
bufg_50: ENTITY WORK.bufg
    PORT MAP (
        in1 => DP_addrBus_5,
        out1 => addrBus(5)
    );
bufg_51: ENTITY WORK.bufg
    PORT MAP (
        in1 => DP_addrBus_6,
        out1 => addrBus(6)
    );
bufg_52: ENTITY WORK.bufg
    PORT MAP (
        in1 => DP_addrBus_7,
        out1 => addrBus(7)
    );
bufg_53: ENTITY WORK.bufg
    PORT MAP (
        in1 => DP_addrBus_8,
        out1 => addrBus(8)
    );
bufg_54: ENTITY WORK.bufg
    PORT MAP (
        in1 => DP_addrBus_9,
        out1 => addrBus(9)
    );
bufg_55: ENTITY WORK.bufg
    PORT MAP (
        in1 => clk,
        out1 => CU_clk
    );
bufg_56: ENTITY WORK.bufg
    PORT MAP (
        in1 => CU_readMEM,
        out1 => readMEM
    );
bufg_57: ENTITY WORK.bufg
    PORT MAP (
        in1 => rst,
        out1 => CU_rst
    );
bufg_58: ENTITY WORK.bufg
    PORT MAP (
        in1 => CU_seldataBus,
        out1 => writeMEM
    );

END ARCHITECTURE arch;
