module MAPn(clk, rst, run, pause, din, w, reg_out, dout);

wire S0;
wire S1;
wire S2;
wire S3;
wire S4;
wire S5;
wire S6;
wire S7;
wire data_out_map_0;
wire data_out_map_100;
wire data_out_map_101;
wire data_out_map_102;
wire data_out_map_103;
wire data_out_map_104;
wire data_out_map_105;
wire data_out_map_106;
wire data_out_map_107;
wire data_out_map_108;
wire data_out_map_109;
wire data_out_map_10;
wire data_out_map_110;
wire data_out_map_111;
wire data_out_map_112;
wire data_out_map_113;
wire data_out_map_114;
wire data_out_map_115;
wire data_out_map_116;
wire data_out_map_117;
wire data_out_map_118;
wire data_out_map_119;
wire data_out_map_11;
wire data_out_map_120;
wire data_out_map_121;
wire data_out_map_122;
wire data_out_map_123;
wire data_out_map_124;
wire data_out_map_125;
wire data_out_map_126;
wire data_out_map_127;
wire data_out_map_12;
wire data_out_map_13;
wire data_out_map_14;
wire data_out_map_15;
wire data_out_map_16;
wire data_out_map_17;
wire data_out_map_18;
wire data_out_map_19;
wire data_out_map_1;
wire data_out_map_20;
wire data_out_map_21;
wire data_out_map_22;
wire data_out_map_23;
wire data_out_map_24;
wire data_out_map_25;
wire data_out_map_26;
wire data_out_map_27;
wire data_out_map_28;
wire data_out_map_29;
wire data_out_map_2;
wire data_out_map_30;
wire data_out_map_31;
wire data_out_map_32;
wire data_out_map_33;
wire data_out_map_34;
wire data_out_map_35;
wire data_out_map_36;
wire data_out_map_37;
wire data_out_map_38;
wire data_out_map_39;
wire data_out_map_3;
wire data_out_map_40;
wire data_out_map_41;
wire data_out_map_42;
wire data_out_map_43;
wire data_out_map_44;
wire data_out_map_45;
wire data_out_map_46;
wire data_out_map_47;
wire data_out_map_48;
wire data_out_map_49;
wire data_out_map_4;
wire data_out_map_50;
wire data_out_map_51;
wire data_out_map_52;
wire data_out_map_53;
wire data_out_map_54;
wire data_out_map_55;
wire data_out_map_56;
wire data_out_map_57;
wire data_out_map_58;
wire data_out_map_59;
wire data_out_map_5;
wire data_out_map_60;
wire data_out_map_61;
wire data_out_map_62;
wire data_out_map_63;
wire data_out_map_64;
wire data_out_map_65;
wire data_out_map_66;
wire data_out_map_67;
wire data_out_map_68;
wire data_out_map_69;
wire data_out_map_6;
wire data_out_map_70;
wire data_out_map_71;
wire data_out_map_72;
wire data_out_map_73;
wire data_out_map_74;
wire data_out_map_75;
wire data_out_map_76;
wire data_out_map_77;
wire data_out_map_78;
wire data_out_map_79;
wire data_out_map_7;
wire data_out_map_80;
wire data_out_map_81;
wire data_out_map_82;
wire data_out_map_83;
wire data_out_map_84;
wire data_out_map_85;
wire data_out_map_86;
wire data_out_map_87;
wire data_out_map_88;
wire data_out_map_89;
wire data_out_map_8;
wire data_out_map_90;
wire data_out_map_91;
wire data_out_map_92;
wire data_out_map_93;
wire data_out_map_94;
wire data_out_map_95;
wire data_out_map_96;
wire data_out_map_97;
wire data_out_map_98;
wire data_out_map_99;
wire data_out_map_9;
wire hb0_map_ns_for:1_map_ns:4;
wire hb0_map_ns_for:2_map_ns:13;
wire hb0_map_ns_for:3_map_ns:22;
wire hb0_map_ns_for:4_map_ns:31;
input clk;
input rst;
input run;
input pause;
input [383:0] din;input [383:0] w;output reg_out;
output [31:0] dout;
BUF_X1 #() 
BUF_X1_1_ (
  .A({ clk }),
  .Z({ S0 })
);
BUF_X1 #() 
BUF_X1_2_ (
  .A({ din[0] }),
  .Z({ S1[0] })
);
BUF_X1 #() 
BUF_X1_3_ (
  .A({ din[1] }),
  .Z({ S1[1] })
);
BUF_X1 #() 
BUF_X1_4_ (
  .A({ din[10] }),
  .Z({ S1[10] })
);
BUF_X1 #() 
BUF_X1_5_ (
  .A({ din[100] }),
  .Z({ S1[100] })
);
BUF_X1 #() 
BUF_X1_6_ (
  .A({ din[101] }),
  .Z({ S1[101] })
);
BUF_X1 #() 
BUF_X1_7_ (
  .A({ din[102] }),
  .Z({ S1[102] })
);
BUF_X1 #() 
BUF_X1_8_ (
  .A({ din[103] }),
  .Z({ S1[103] })
);
BUF_X1 #() 
BUF_X1_9_ (
  .A({ din[104] }),
  .Z({ S1[104] })
);
BUF_X1 #() 
BUF_X1_10_ (
  .A({ din[105] }),
  .Z({ S1[105] })
);
BUF_X1 #() 
BUF_X1_11_ (
  .A({ din[106] }),
  .Z({ S1[106] })
);
BUF_X1 #() 
BUF_X1_12_ (
  .A({ din[107] }),
  .Z({ S1[107] })
);
BUF_X1 #() 
BUF_X1_13_ (
  .A({ din[108] }),
  .Z({ S1[108] })
);
BUF_X1 #() 
BUF_X1_14_ (
  .A({ din[109] }),
  .Z({ S1[109] })
);
BUF_X1 #() 
BUF_X1_15_ (
  .A({ din[11] }),
  .Z({ S1[11] })
);
BUF_X1 #() 
BUF_X1_16_ (
  .A({ din[110] }),
  .Z({ S1[110] })
);
BUF_X1 #() 
BUF_X1_17_ (
  .A({ din[111] }),
  .Z({ S1[111] })
);
BUF_X1 #() 
BUF_X1_18_ (
  .A({ din[112] }),
  .Z({ S1[112] })
);
BUF_X1 #() 
BUF_X1_19_ (
  .A({ din[113] }),
  .Z({ S1[113] })
);
BUF_X1 #() 
BUF_X1_20_ (
  .A({ din[114] }),
  .Z({ S1[114] })
);
BUF_X1 #() 
BUF_X1_21_ (
  .A({ din[115] }),
  .Z({ S1[115] })
);
BUF_X1 #() 
BUF_X1_22_ (
  .A({ din[116] }),
  .Z({ S1[116] })
);
BUF_X1 #() 
BUF_X1_23_ (
  .A({ din[117] }),
  .Z({ S1[117] })
);
BUF_X1 #() 
BUF_X1_24_ (
  .A({ din[118] }),
  .Z({ S1[118] })
);
BUF_X1 #() 
BUF_X1_25_ (
  .A({ din[119] }),
  .Z({ S1[119] })
);
BUF_X1 #() 
BUF_X1_26_ (
  .A({ din[12] }),
  .Z({ S1[12] })
);
BUF_X1 #() 
BUF_X1_27_ (
  .A({ din[120] }),
  .Z({ S1[120] })
);
BUF_X1 #() 
BUF_X1_28_ (
  .A({ din[121] }),
  .Z({ S1[121] })
);
BUF_X1 #() 
BUF_X1_29_ (
  .A({ din[122] }),
  .Z({ S1[122] })
);
BUF_X1 #() 
BUF_X1_30_ (
  .A({ din[123] }),
  .Z({ S1[123] })
);
BUF_X1 #() 
BUF_X1_31_ (
  .A({ din[124] }),
  .Z({ S1[124] })
);
BUF_X1 #() 
BUF_X1_32_ (
  .A({ din[125] }),
  .Z({ S1[125] })
);
BUF_X1 #() 
BUF_X1_33_ (
  .A({ din[126] }),
  .Z({ S1[126] })
);
BUF_X1 #() 
BUF_X1_34_ (
  .A({ din[127] }),
  .Z({ S1[127] })
);
BUF_X1 #() 
BUF_X1_35_ (
  .A({ din[128] }),
  .Z({ S1[128] })
);
BUF_X1 #() 
BUF_X1_36_ (
  .A({ din[129] }),
  .Z({ S1[129] })
);
BUF_X1 #() 
BUF_X1_37_ (
  .A({ din[13] }),
  .Z({ S1[13] })
);
BUF_X1 #() 
BUF_X1_38_ (
  .A({ din[130] }),
  .Z({ S1[130] })
);
BUF_X1 #() 
BUF_X1_39_ (
  .A({ din[131] }),
  .Z({ S1[131] })
);
BUF_X1 #() 
BUF_X1_40_ (
  .A({ din[132] }),
  .Z({ S1[132] })
);
BUF_X1 #() 
BUF_X1_41_ (
  .A({ din[133] }),
  .Z({ S1[133] })
);
BUF_X1 #() 
BUF_X1_42_ (
  .A({ din[134] }),
  .Z({ S1[134] })
);
BUF_X1 #() 
BUF_X1_43_ (
  .A({ din[135] }),
  .Z({ S1[135] })
);
BUF_X1 #() 
BUF_X1_44_ (
  .A({ din[136] }),
  .Z({ S1[136] })
);
BUF_X1 #() 
BUF_X1_45_ (
  .A({ din[137] }),
  .Z({ S1[137] })
);
BUF_X1 #() 
BUF_X1_46_ (
  .A({ din[138] }),
  .Z({ S1[138] })
);
BUF_X1 #() 
BUF_X1_47_ (
  .A({ din[139] }),
  .Z({ S1[139] })
);
BUF_X1 #() 
BUF_X1_48_ (
  .A({ din[14] }),
  .Z({ S1[14] })
);
BUF_X1 #() 
BUF_X1_49_ (
  .A({ din[140] }),
  .Z({ S1[140] })
);
BUF_X1 #() 
BUF_X1_50_ (
  .A({ din[141] }),
  .Z({ S1[141] })
);
BUF_X1 #() 
BUF_X1_51_ (
  .A({ din[142] }),
  .Z({ S1[142] })
);
BUF_X1 #() 
BUF_X1_52_ (
  .A({ din[143] }),
  .Z({ S1[143] })
);
BUF_X1 #() 
BUF_X1_53_ (
  .A({ din[144] }),
  .Z({ S1[144] })
);
BUF_X1 #() 
BUF_X1_54_ (
  .A({ din[145] }),
  .Z({ S1[145] })
);
BUF_X1 #() 
BUF_X1_55_ (
  .A({ din[146] }),
  .Z({ S1[146] })
);
BUF_X1 #() 
BUF_X1_56_ (
  .A({ din[147] }),
  .Z({ S1[147] })
);
BUF_X1 #() 
BUF_X1_57_ (
  .A({ din[148] }),
  .Z({ S1[148] })
);
BUF_X1 #() 
BUF_X1_58_ (
  .A({ din[149] }),
  .Z({ S1[149] })
);
BUF_X1 #() 
BUF_X1_59_ (
  .A({ din[15] }),
  .Z({ S1[15] })
);
BUF_X1 #() 
BUF_X1_60_ (
  .A({ din[150] }),
  .Z({ S1[150] })
);
BUF_X1 #() 
BUF_X1_61_ (
  .A({ din[151] }),
  .Z({ S1[151] })
);
BUF_X1 #() 
BUF_X1_62_ (
  .A({ din[152] }),
  .Z({ S1[152] })
);
BUF_X1 #() 
BUF_X1_63_ (
  .A({ din[153] }),
  .Z({ S1[153] })
);
BUF_X1 #() 
BUF_X1_64_ (
  .A({ din[154] }),
  .Z({ S1[154] })
);
BUF_X1 #() 
BUF_X1_65_ (
  .A({ din[155] }),
  .Z({ S1[155] })
);
BUF_X1 #() 
BUF_X1_66_ (
  .A({ din[156] }),
  .Z({ S1[156] })
);
BUF_X1 #() 
BUF_X1_67_ (
  .A({ din[157] }),
  .Z({ S1[157] })
);
BUF_X1 #() 
BUF_X1_68_ (
  .A({ din[158] }),
  .Z({ S1[158] })
);
BUF_X1 #() 
BUF_X1_69_ (
  .A({ din[159] }),
  .Z({ S1[159] })
);
BUF_X1 #() 
BUF_X1_70_ (
  .A({ din[16] }),
  .Z({ S1[16] })
);
BUF_X1 #() 
BUF_X1_71_ (
  .A({ din[160] }),
  .Z({ S1[160] })
);
BUF_X1 #() 
BUF_X1_72_ (
  .A({ din[161] }),
  .Z({ S1[161] })
);
BUF_X1 #() 
BUF_X1_73_ (
  .A({ din[162] }),
  .Z({ S1[162] })
);
BUF_X1 #() 
BUF_X1_74_ (
  .A({ din[163] }),
  .Z({ S1[163] })
);
BUF_X1 #() 
BUF_X1_75_ (
  .A({ din[164] }),
  .Z({ S1[164] })
);
BUF_X1 #() 
BUF_X1_76_ (
  .A({ din[165] }),
  .Z({ S1[165] })
);
BUF_X1 #() 
BUF_X1_77_ (
  .A({ din[166] }),
  .Z({ S1[166] })
);
BUF_X1 #() 
BUF_X1_78_ (
  .A({ din[167] }),
  .Z({ S1[167] })
);
BUF_X1 #() 
BUF_X1_79_ (
  .A({ din[168] }),
  .Z({ S1[168] })
);
BUF_X1 #() 
BUF_X1_80_ (
  .A({ din[169] }),
  .Z({ S1[169] })
);
BUF_X1 #() 
BUF_X1_81_ (
  .A({ din[17] }),
  .Z({ S1[17] })
);
BUF_X1 #() 
BUF_X1_82_ (
  .A({ din[170] }),
  .Z({ S1[170] })
);
BUF_X1 #() 
BUF_X1_83_ (
  .A({ din[171] }),
  .Z({ S1[171] })
);
BUF_X1 #() 
BUF_X1_84_ (
  .A({ din[172] }),
  .Z({ S1[172] })
);
BUF_X1 #() 
BUF_X1_85_ (
  .A({ din[173] }),
  .Z({ S1[173] })
);
BUF_X1 #() 
BUF_X1_86_ (
  .A({ din[174] }),
  .Z({ S1[174] })
);
BUF_X1 #() 
BUF_X1_87_ (
  .A({ din[175] }),
  .Z({ S1[175] })
);
BUF_X1 #() 
BUF_X1_88_ (
  .A({ din[176] }),
  .Z({ S1[176] })
);
BUF_X1 #() 
BUF_X1_89_ (
  .A({ din[177] }),
  .Z({ S1[177] })
);
BUF_X1 #() 
BUF_X1_90_ (
  .A({ din[178] }),
  .Z({ S1[178] })
);
BUF_X1 #() 
BUF_X1_91_ (
  .A({ din[179] }),
  .Z({ S1[179] })
);
BUF_X1 #() 
BUF_X1_92_ (
  .A({ din[18] }),
  .Z({ S1[18] })
);
BUF_X1 #() 
BUF_X1_93_ (
  .A({ din[180] }),
  .Z({ S1[180] })
);
BUF_X1 #() 
BUF_X1_94_ (
  .A({ din[181] }),
  .Z({ S1[181] })
);
BUF_X1 #() 
BUF_X1_95_ (
  .A({ din[182] }),
  .Z({ S1[182] })
);
BUF_X1 #() 
BUF_X1_96_ (
  .A({ din[183] }),
  .Z({ S1[183] })
);
BUF_X1 #() 
BUF_X1_97_ (
  .A({ din[184] }),
  .Z({ S1[184] })
);
BUF_X1 #() 
BUF_X1_98_ (
  .A({ din[185] }),
  .Z({ S1[185] })
);
BUF_X1 #() 
BUF_X1_99_ (
  .A({ din[186] }),
  .Z({ S1[186] })
);
BUF_X1 #() 
BUF_X1_100_ (
  .A({ din[187] }),
  .Z({ S1[187] })
);
BUF_X1 #() 
BUF_X1_101_ (
  .A({ din[188] }),
  .Z({ S1[188] })
);
BUF_X1 #() 
BUF_X1_102_ (
  .A({ din[189] }),
  .Z({ S1[189] })
);
BUF_X1 #() 
BUF_X1_103_ (
  .A({ din[19] }),
  .Z({ S1[19] })
);
BUF_X1 #() 
BUF_X1_104_ (
  .A({ din[190] }),
  .Z({ S1[190] })
);
BUF_X1 #() 
BUF_X1_105_ (
  .A({ din[191] }),
  .Z({ S1[191] })
);
BUF_X1 #() 
BUF_X1_106_ (
  .A({ din[192] }),
  .Z({ S1[192] })
);
BUF_X1 #() 
BUF_X1_107_ (
  .A({ din[193] }),
  .Z({ S1[193] })
);
BUF_X1 #() 
BUF_X1_108_ (
  .A({ din[194] }),
  .Z({ S1[194] })
);
BUF_X1 #() 
BUF_X1_109_ (
  .A({ din[195] }),
  .Z({ S1[195] })
);
BUF_X1 #() 
BUF_X1_110_ (
  .A({ din[196] }),
  .Z({ S1[196] })
);
BUF_X1 #() 
BUF_X1_111_ (
  .A({ din[197] }),
  .Z({ S1[197] })
);
BUF_X1 #() 
BUF_X1_112_ (
  .A({ din[198] }),
  .Z({ S1[198] })
);
BUF_X1 #() 
BUF_X1_113_ (
  .A({ din[199] }),
  .Z({ S1[199] })
);
BUF_X1 #() 
BUF_X1_114_ (
  .A({ din[2] }),
  .Z({ S1[2] })
);
BUF_X1 #() 
BUF_X1_115_ (
  .A({ din[20] }),
  .Z({ S1[20] })
);
BUF_X1 #() 
BUF_X1_116_ (
  .A({ din[200] }),
  .Z({ S1[200] })
);
BUF_X1 #() 
BUF_X1_117_ (
  .A({ din[201] }),
  .Z({ S1[201] })
);
BUF_X1 #() 
BUF_X1_118_ (
  .A({ din[202] }),
  .Z({ S1[202] })
);
BUF_X1 #() 
BUF_X1_119_ (
  .A({ din[203] }),
  .Z({ S1[203] })
);
BUF_X1 #() 
BUF_X1_120_ (
  .A({ din[204] }),
  .Z({ S1[204] })
);
BUF_X1 #() 
BUF_X1_121_ (
  .A({ din[205] }),
  .Z({ S1[205] })
);
BUF_X1 #() 
BUF_X1_122_ (
  .A({ din[206] }),
  .Z({ S1[206] })
);
BUF_X1 #() 
BUF_X1_123_ (
  .A({ din[207] }),
  .Z({ S1[207] })
);
BUF_X1 #() 
BUF_X1_124_ (
  .A({ din[208] }),
  .Z({ S1[208] })
);
BUF_X1 #() 
BUF_X1_125_ (
  .A({ din[209] }),
  .Z({ S1[209] })
);
BUF_X1 #() 
BUF_X1_126_ (
  .A({ din[21] }),
  .Z({ S1[21] })
);
BUF_X1 #() 
BUF_X1_127_ (
  .A({ din[210] }),
  .Z({ S1[210] })
);
BUF_X1 #() 
BUF_X1_128_ (
  .A({ din[211] }),
  .Z({ S1[211] })
);
BUF_X1 #() 
BUF_X1_129_ (
  .A({ din[212] }),
  .Z({ S1[212] })
);
BUF_X1 #() 
BUF_X1_130_ (
  .A({ din[213] }),
  .Z({ S1[213] })
);
BUF_X1 #() 
BUF_X1_131_ (
  .A({ din[214] }),
  .Z({ S1[214] })
);
BUF_X1 #() 
BUF_X1_132_ (
  .A({ din[215] }),
  .Z({ S1[215] })
);
BUF_X1 #() 
BUF_X1_133_ (
  .A({ din[216] }),
  .Z({ S1[216] })
);
BUF_X1 #() 
BUF_X1_134_ (
  .A({ din[217] }),
  .Z({ S1[217] })
);
BUF_X1 #() 
BUF_X1_135_ (
  .A({ din[218] }),
  .Z({ S1[218] })
);
BUF_X1 #() 
BUF_X1_136_ (
  .A({ din[219] }),
  .Z({ S1[219] })
);
BUF_X1 #() 
BUF_X1_137_ (
  .A({ din[22] }),
  .Z({ S1[22] })
);
BUF_X1 #() 
BUF_X1_138_ (
  .A({ din[220] }),
  .Z({ S1[220] })
);
BUF_X1 #() 
BUF_X1_139_ (
  .A({ din[221] }),
  .Z({ S1[221] })
);
BUF_X1 #() 
BUF_X1_140_ (
  .A({ din[222] }),
  .Z({ S1[222] })
);
BUF_X1 #() 
BUF_X1_141_ (
  .A({ din[223] }),
  .Z({ S1[223] })
);
BUF_X1 #() 
BUF_X1_142_ (
  .A({ din[224] }),
  .Z({ S1[224] })
);
BUF_X1 #() 
BUF_X1_143_ (
  .A({ din[225] }),
  .Z({ S1[225] })
);
BUF_X1 #() 
BUF_X1_144_ (
  .A({ din[226] }),
  .Z({ S1[226] })
);
BUF_X1 #() 
BUF_X1_145_ (
  .A({ din[227] }),
  .Z({ S1[227] })
);
BUF_X1 #() 
BUF_X1_146_ (
  .A({ din[228] }),
  .Z({ S1[228] })
);
BUF_X1 #() 
BUF_X1_147_ (
  .A({ din[229] }),
  .Z({ S1[229] })
);
BUF_X1 #() 
BUF_X1_148_ (
  .A({ din[23] }),
  .Z({ S1[23] })
);
BUF_X1 #() 
BUF_X1_149_ (
  .A({ din[230] }),
  .Z({ S1[230] })
);
BUF_X1 #() 
BUF_X1_150_ (
  .A({ din[231] }),
  .Z({ S1[231] })
);
BUF_X1 #() 
BUF_X1_151_ (
  .A({ din[232] }),
  .Z({ S1[232] })
);
BUF_X1 #() 
BUF_X1_152_ (
  .A({ din[233] }),
  .Z({ S1[233] })
);
BUF_X1 #() 
BUF_X1_153_ (
  .A({ din[234] }),
  .Z({ S1[234] })
);
BUF_X1 #() 
BUF_X1_154_ (
  .A({ din[235] }),
  .Z({ S1[235] })
);
BUF_X1 #() 
BUF_X1_155_ (
  .A({ din[236] }),
  .Z({ S1[236] })
);
BUF_X1 #() 
BUF_X1_156_ (
  .A({ din[237] }),
  .Z({ S1[237] })
);
BUF_X1 #() 
BUF_X1_157_ (
  .A({ din[238] }),
  .Z({ S1[238] })
);
BUF_X1 #() 
BUF_X1_158_ (
  .A({ din[239] }),
  .Z({ S1[239] })
);
BUF_X1 #() 
BUF_X1_159_ (
  .A({ din[24] }),
  .Z({ S1[24] })
);
BUF_X1 #() 
BUF_X1_160_ (
  .A({ din[240] }),
  .Z({ S1[240] })
);
BUF_X1 #() 
BUF_X1_161_ (
  .A({ din[241] }),
  .Z({ S1[241] })
);
BUF_X1 #() 
BUF_X1_162_ (
  .A({ din[242] }),
  .Z({ S1[242] })
);
BUF_X1 #() 
BUF_X1_163_ (
  .A({ din[243] }),
  .Z({ S1[243] })
);
BUF_X1 #() 
BUF_X1_164_ (
  .A({ din[244] }),
  .Z({ S1[244] })
);
BUF_X1 #() 
BUF_X1_165_ (
  .A({ din[245] }),
  .Z({ S1[245] })
);
BUF_X1 #() 
BUF_X1_166_ (
  .A({ din[246] }),
  .Z({ S1[246] })
);
BUF_X1 #() 
BUF_X1_167_ (
  .A({ din[247] }),
  .Z({ S1[247] })
);
BUF_X1 #() 
BUF_X1_168_ (
  .A({ din[248] }),
  .Z({ S1[248] })
);
BUF_X1 #() 
BUF_X1_169_ (
  .A({ din[249] }),
  .Z({ S1[249] })
);
BUF_X1 #() 
BUF_X1_170_ (
  .A({ din[25] }),
  .Z({ S1[25] })
);
BUF_X1 #() 
BUF_X1_171_ (
  .A({ din[250] }),
  .Z({ S1[250] })
);
BUF_X1 #() 
BUF_X1_172_ (
  .A({ din[251] }),
  .Z({ S1[251] })
);
BUF_X1 #() 
BUF_X1_173_ (
  .A({ din[252] }),
  .Z({ S1[252] })
);
BUF_X1 #() 
BUF_X1_174_ (
  .A({ din[253] }),
  .Z({ S1[253] })
);
BUF_X1 #() 
BUF_X1_175_ (
  .A({ din[254] }),
  .Z({ S1[254] })
);
BUF_X1 #() 
BUF_X1_176_ (
  .A({ din[255] }),
  .Z({ S1[255] })
);
BUF_X1 #() 
BUF_X1_177_ (
  .A({ din[256] }),
  .Z({ S1[256] })
);
BUF_X1 #() 
BUF_X1_178_ (
  .A({ din[257] }),
  .Z({ S1[257] })
);
BUF_X1 #() 
BUF_X1_179_ (
  .A({ din[258] }),
  .Z({ S1[258] })
);
BUF_X1 #() 
BUF_X1_180_ (
  .A({ din[259] }),
  .Z({ S1[259] })
);
BUF_X1 #() 
BUF_X1_181_ (
  .A({ din[26] }),
  .Z({ S1[26] })
);
BUF_X1 #() 
BUF_X1_182_ (
  .A({ din[260] }),
  .Z({ S1[260] })
);
BUF_X1 #() 
BUF_X1_183_ (
  .A({ din[261] }),
  .Z({ S1[261] })
);
BUF_X1 #() 
BUF_X1_184_ (
  .A({ din[262] }),
  .Z({ S1[262] })
);
BUF_X1 #() 
BUF_X1_185_ (
  .A({ din[263] }),
  .Z({ S1[263] })
);
BUF_X1 #() 
BUF_X1_186_ (
  .A({ din[264] }),
  .Z({ S1[264] })
);
BUF_X1 #() 
BUF_X1_187_ (
  .A({ din[265] }),
  .Z({ S1[265] })
);
BUF_X1 #() 
BUF_X1_188_ (
  .A({ din[266] }),
  .Z({ S1[266] })
);
BUF_X1 #() 
BUF_X1_189_ (
  .A({ din[267] }),
  .Z({ S1[267] })
);
BUF_X1 #() 
BUF_X1_190_ (
  .A({ din[268] }),
  .Z({ S1[268] })
);
BUF_X1 #() 
BUF_X1_191_ (
  .A({ din[269] }),
  .Z({ S1[269] })
);
BUF_X1 #() 
BUF_X1_192_ (
  .A({ din[27] }),
  .Z({ S1[27] })
);
BUF_X1 #() 
BUF_X1_193_ (
  .A({ din[270] }),
  .Z({ S1[270] })
);
BUF_X1 #() 
BUF_X1_194_ (
  .A({ din[271] }),
  .Z({ S1[271] })
);
BUF_X1 #() 
BUF_X1_195_ (
  .A({ din[272] }),
  .Z({ S1[272] })
);
BUF_X1 #() 
BUF_X1_196_ (
  .A({ din[273] }),
  .Z({ S1[273] })
);
BUF_X1 #() 
BUF_X1_197_ (
  .A({ din[274] }),
  .Z({ S1[274] })
);
BUF_X1 #() 
BUF_X1_198_ (
  .A({ din[275] }),
  .Z({ S1[275] })
);
BUF_X1 #() 
BUF_X1_199_ (
  .A({ din[276] }),
  .Z({ S1[276] })
);
BUF_X1 #() 
BUF_X1_200_ (
  .A({ din[277] }),
  .Z({ S1[277] })
);
BUF_X1 #() 
BUF_X1_201_ (
  .A({ din[278] }),
  .Z({ S1[278] })
);
BUF_X1 #() 
BUF_X1_202_ (
  .A({ din[279] }),
  .Z({ S1[279] })
);
BUF_X1 #() 
BUF_X1_203_ (
  .A({ din[28] }),
  .Z({ S1[28] })
);
BUF_X1 #() 
BUF_X1_204_ (
  .A({ din[280] }),
  .Z({ S1[280] })
);
BUF_X1 #() 
BUF_X1_205_ (
  .A({ din[281] }),
  .Z({ S1[281] })
);
BUF_X1 #() 
BUF_X1_206_ (
  .A({ din[282] }),
  .Z({ S1[282] })
);
BUF_X1 #() 
BUF_X1_207_ (
  .A({ din[283] }),
  .Z({ S1[283] })
);
BUF_X1 #() 
BUF_X1_208_ (
  .A({ din[284] }),
  .Z({ S1[284] })
);
BUF_X1 #() 
BUF_X1_209_ (
  .A({ din[285] }),
  .Z({ S1[285] })
);
BUF_X1 #() 
BUF_X1_210_ (
  .A({ din[286] }),
  .Z({ S1[286] })
);
BUF_X1 #() 
BUF_X1_211_ (
  .A({ din[287] }),
  .Z({ S1[287] })
);
BUF_X1 #() 
BUF_X1_212_ (
  .A({ din[288] }),
  .Z({ S1[288] })
);
BUF_X1 #() 
BUF_X1_213_ (
  .A({ din[289] }),
  .Z({ S1[289] })
);
BUF_X1 #() 
BUF_X1_214_ (
  .A({ din[29] }),
  .Z({ S1[29] })
);
BUF_X1 #() 
BUF_X1_215_ (
  .A({ din[290] }),
  .Z({ S1[290] })
);
BUF_X1 #() 
BUF_X1_216_ (
  .A({ din[291] }),
  .Z({ S1[291] })
);
BUF_X1 #() 
BUF_X1_217_ (
  .A({ din[292] }),
  .Z({ S1[292] })
);
BUF_X1 #() 
BUF_X1_218_ (
  .A({ din[293] }),
  .Z({ S1[293] })
);
BUF_X1 #() 
BUF_X1_219_ (
  .A({ din[294] }),
  .Z({ S1[294] })
);
BUF_X1 #() 
BUF_X1_220_ (
  .A({ din[295] }),
  .Z({ S1[295] })
);
BUF_X1 #() 
BUF_X1_221_ (
  .A({ din[296] }),
  .Z({ S1[296] })
);
BUF_X1 #() 
BUF_X1_222_ (
  .A({ din[297] }),
  .Z({ S1[297] })
);
BUF_X1 #() 
BUF_X1_223_ (
  .A({ din[298] }),
  .Z({ S1[298] })
);
BUF_X1 #() 
BUF_X1_224_ (
  .A({ din[299] }),
  .Z({ S1[299] })
);
BUF_X1 #() 
BUF_X1_225_ (
  .A({ din[3] }),
  .Z({ S1[3] })
);
BUF_X1 #() 
BUF_X1_226_ (
  .A({ din[30] }),
  .Z({ S1[30] })
);
BUF_X1 #() 
BUF_X1_227_ (
  .A({ din[300] }),
  .Z({ S1[300] })
);
BUF_X1 #() 
BUF_X1_228_ (
  .A({ din[301] }),
  .Z({ S1[301] })
);
BUF_X1 #() 
BUF_X1_229_ (
  .A({ din[302] }),
  .Z({ S1[302] })
);
BUF_X1 #() 
BUF_X1_230_ (
  .A({ din[303] }),
  .Z({ S1[303] })
);
BUF_X1 #() 
BUF_X1_231_ (
  .A({ din[304] }),
  .Z({ S1[304] })
);
BUF_X1 #() 
BUF_X1_232_ (
  .A({ din[305] }),
  .Z({ S1[305] })
);
BUF_X1 #() 
BUF_X1_233_ (
  .A({ din[306] }),
  .Z({ S1[306] })
);
BUF_X1 #() 
BUF_X1_234_ (
  .A({ din[307] }),
  .Z({ S1[307] })
);
BUF_X1 #() 
BUF_X1_235_ (
  .A({ din[308] }),
  .Z({ S1[308] })
);
BUF_X1 #() 
BUF_X1_236_ (
  .A({ din[309] }),
  .Z({ S1[309] })
);
BUF_X1 #() 
BUF_X1_237_ (
  .A({ din[31] }),
  .Z({ S1[31] })
);
BUF_X1 #() 
BUF_X1_238_ (
  .A({ din[310] }),
  .Z({ S1[310] })
);
BUF_X1 #() 
BUF_X1_239_ (
  .A({ din[311] }),
  .Z({ S1[311] })
);
BUF_X1 #() 
BUF_X1_240_ (
  .A({ din[312] }),
  .Z({ S1[312] })
);
BUF_X1 #() 
BUF_X1_241_ (
  .A({ din[313] }),
  .Z({ S1[313] })
);
BUF_X1 #() 
BUF_X1_242_ (
  .A({ din[314] }),
  .Z({ S1[314] })
);
BUF_X1 #() 
BUF_X1_243_ (
  .A({ din[315] }),
  .Z({ S1[315] })
);
BUF_X1 #() 
BUF_X1_244_ (
  .A({ din[316] }),
  .Z({ S1[316] })
);
BUF_X1 #() 
BUF_X1_245_ (
  .A({ din[317] }),
  .Z({ S1[317] })
);
BUF_X1 #() 
BUF_X1_246_ (
  .A({ din[318] }),
  .Z({ S1[318] })
);
BUF_X1 #() 
BUF_X1_247_ (
  .A({ din[319] }),
  .Z({ S1[319] })
);
BUF_X1 #() 
BUF_X1_248_ (
  .A({ din[32] }),
  .Z({ S1[32] })
);
BUF_X1 #() 
BUF_X1_249_ (
  .A({ din[320] }),
  .Z({ S1[320] })
);
BUF_X1 #() 
BUF_X1_250_ (
  .A({ din[321] }),
  .Z({ S1[321] })
);
BUF_X1 #() 
BUF_X1_251_ (
  .A({ din[322] }),
  .Z({ S1[322] })
);
BUF_X1 #() 
BUF_X1_252_ (
  .A({ din[323] }),
  .Z({ S1[323] })
);
BUF_X1 #() 
BUF_X1_253_ (
  .A({ din[324] }),
  .Z({ S1[324] })
);
BUF_X1 #() 
BUF_X1_254_ (
  .A({ din[325] }),
  .Z({ S1[325] })
);
BUF_X1 #() 
BUF_X1_255_ (
  .A({ din[326] }),
  .Z({ S1[326] })
);
BUF_X1 #() 
BUF_X1_256_ (
  .A({ din[327] }),
  .Z({ S1[327] })
);
BUF_X1 #() 
BUF_X1_257_ (
  .A({ din[328] }),
  .Z({ S1[328] })
);
BUF_X1 #() 
BUF_X1_258_ (
  .A({ din[329] }),
  .Z({ S1[329] })
);
BUF_X1 #() 
BUF_X1_259_ (
  .A({ din[33] }),
  .Z({ S1[33] })
);
BUF_X1 #() 
BUF_X1_260_ (
  .A({ din[330] }),
  .Z({ S1[330] })
);
BUF_X1 #() 
BUF_X1_261_ (
  .A({ din[331] }),
  .Z({ S1[331] })
);
BUF_X1 #() 
BUF_X1_262_ (
  .A({ din[332] }),
  .Z({ S1[332] })
);
BUF_X1 #() 
BUF_X1_263_ (
  .A({ din[333] }),
  .Z({ S1[333] })
);
BUF_X1 #() 
BUF_X1_264_ (
  .A({ din[334] }),
  .Z({ S1[334] })
);
BUF_X1 #() 
BUF_X1_265_ (
  .A({ din[335] }),
  .Z({ S1[335] })
);
BUF_X1 #() 
BUF_X1_266_ (
  .A({ din[336] }),
  .Z({ S1[336] })
);
BUF_X1 #() 
BUF_X1_267_ (
  .A({ din[337] }),
  .Z({ S1[337] })
);
BUF_X1 #() 
BUF_X1_268_ (
  .A({ din[338] }),
  .Z({ S1[338] })
);
BUF_X1 #() 
BUF_X1_269_ (
  .A({ din[339] }),
  .Z({ S1[339] })
);
BUF_X1 #() 
BUF_X1_270_ (
  .A({ din[34] }),
  .Z({ S1[34] })
);
BUF_X1 #() 
BUF_X1_271_ (
  .A({ din[340] }),
  .Z({ S1[340] })
);
BUF_X1 #() 
BUF_X1_272_ (
  .A({ din[341] }),
  .Z({ S1[341] })
);
BUF_X1 #() 
BUF_X1_273_ (
  .A({ din[342] }),
  .Z({ S1[342] })
);
BUF_X1 #() 
BUF_X1_274_ (
  .A({ din[343] }),
  .Z({ S1[343] })
);
BUF_X1 #() 
BUF_X1_275_ (
  .A({ din[344] }),
  .Z({ S1[344] })
);
BUF_X1 #() 
BUF_X1_276_ (
  .A({ din[345] }),
  .Z({ S1[345] })
);
BUF_X1 #() 
BUF_X1_277_ (
  .A({ din[346] }),
  .Z({ S1[346] })
);
BUF_X1 #() 
BUF_X1_278_ (
  .A({ din[347] }),
  .Z({ S1[347] })
);
BUF_X1 #() 
BUF_X1_279_ (
  .A({ din[348] }),
  .Z({ S1[348] })
);
BUF_X1 #() 
BUF_X1_280_ (
  .A({ din[349] }),
  .Z({ S1[349] })
);
BUF_X1 #() 
BUF_X1_281_ (
  .A({ din[35] }),
  .Z({ S1[35] })
);
BUF_X1 #() 
BUF_X1_282_ (
  .A({ din[350] }),
  .Z({ S1[350] })
);
BUF_X1 #() 
BUF_X1_283_ (
  .A({ din[351] }),
  .Z({ S1[351] })
);
BUF_X1 #() 
BUF_X1_284_ (
  .A({ din[352] }),
  .Z({ S1[352] })
);
BUF_X1 #() 
BUF_X1_285_ (
  .A({ din[353] }),
  .Z({ S1[353] })
);
BUF_X1 #() 
BUF_X1_286_ (
  .A({ din[354] }),
  .Z({ S1[354] })
);
BUF_X1 #() 
BUF_X1_287_ (
  .A({ din[355] }),
  .Z({ S1[355] })
);
BUF_X1 #() 
BUF_X1_288_ (
  .A({ din[356] }),
  .Z({ S1[356] })
);
BUF_X1 #() 
BUF_X1_289_ (
  .A({ din[357] }),
  .Z({ S1[357] })
);
BUF_X1 #() 
BUF_X1_290_ (
  .A({ din[358] }),
  .Z({ S1[358] })
);
BUF_X1 #() 
BUF_X1_291_ (
  .A({ din[359] }),
  .Z({ S1[359] })
);
BUF_X1 #() 
BUF_X1_292_ (
  .A({ din[36] }),
  .Z({ S1[36] })
);
BUF_X1 #() 
BUF_X1_293_ (
  .A({ din[360] }),
  .Z({ S1[360] })
);
BUF_X1 #() 
BUF_X1_294_ (
  .A({ din[361] }),
  .Z({ S1[361] })
);
BUF_X1 #() 
BUF_X1_295_ (
  .A({ din[362] }),
  .Z({ S1[362] })
);
BUF_X1 #() 
BUF_X1_296_ (
  .A({ din[363] }),
  .Z({ S1[363] })
);
BUF_X1 #() 
BUF_X1_297_ (
  .A({ din[364] }),
  .Z({ S1[364] })
);
BUF_X1 #() 
BUF_X1_298_ (
  .A({ din[365] }),
  .Z({ S1[365] })
);
BUF_X1 #() 
BUF_X1_299_ (
  .A({ din[366] }),
  .Z({ S1[366] })
);
BUF_X1 #() 
BUF_X1_300_ (
  .A({ din[367] }),
  .Z({ S1[367] })
);
BUF_X1 #() 
BUF_X1_301_ (
  .A({ din[368] }),
  .Z({ S1[368] })
);
BUF_X1 #() 
BUF_X1_302_ (
  .A({ din[369] }),
  .Z({ S1[369] })
);
BUF_X1 #() 
BUF_X1_303_ (
  .A({ din[37] }),
  .Z({ S1[37] })
);
BUF_X1 #() 
BUF_X1_304_ (
  .A({ din[370] }),
  .Z({ S1[370] })
);
BUF_X1 #() 
BUF_X1_305_ (
  .A({ din[371] }),
  .Z({ S1[371] })
);
BUF_X1 #() 
BUF_X1_306_ (
  .A({ din[372] }),
  .Z({ S1[372] })
);
BUF_X1 #() 
BUF_X1_307_ (
  .A({ din[373] }),
  .Z({ S1[373] })
);
BUF_X1 #() 
BUF_X1_308_ (
  .A({ din[374] }),
  .Z({ S1[374] })
);
BUF_X1 #() 
BUF_X1_309_ (
  .A({ din[375] }),
  .Z({ S1[375] })
);
BUF_X1 #() 
BUF_X1_310_ (
  .A({ din[376] }),
  .Z({ S1[376] })
);
BUF_X1 #() 
BUF_X1_311_ (
  .A({ din[377] }),
  .Z({ S1[377] })
);
BUF_X1 #() 
BUF_X1_312_ (
  .A({ din[378] }),
  .Z({ S1[378] })
);
BUF_X1 #() 
BUF_X1_313_ (
  .A({ din[379] }),
  .Z({ S1[379] })
);
BUF_X1 #() 
BUF_X1_314_ (
  .A({ din[38] }),
  .Z({ S1[38] })
);
BUF_X1 #() 
BUF_X1_315_ (
  .A({ din[380] }),
  .Z({ S1[380] })
);
BUF_X1 #() 
BUF_X1_316_ (
  .A({ din[381] }),
  .Z({ S1[381] })
);
BUF_X1 #() 
BUF_X1_317_ (
  .A({ din[382] }),
  .Z({ S1[382] })
);
BUF_X1 #() 
BUF_X1_318_ (
  .A({ din[383] }),
  .Z({ S1[383] })
);
BUF_X1 #() 
BUF_X1_319_ (
  .A({ din[39] }),
  .Z({ S1[39] })
);
BUF_X1 #() 
BUF_X1_320_ (
  .A({ din[4] }),
  .Z({ S1[4] })
);
BUF_X1 #() 
BUF_X1_321_ (
  .A({ din[40] }),
  .Z({ S1[40] })
);
BUF_X1 #() 
BUF_X1_322_ (
  .A({ din[41] }),
  .Z({ S1[41] })
);
BUF_X1 #() 
BUF_X1_323_ (
  .A({ din[42] }),
  .Z({ S1[42] })
);
BUF_X1 #() 
BUF_X1_324_ (
  .A({ din[43] }),
  .Z({ S1[43] })
);
BUF_X1 #() 
BUF_X1_325_ (
  .A({ din[44] }),
  .Z({ S1[44] })
);
BUF_X1 #() 
BUF_X1_326_ (
  .A({ din[45] }),
  .Z({ S1[45] })
);
BUF_X1 #() 
BUF_X1_327_ (
  .A({ din[46] }),
  .Z({ S1[46] })
);
BUF_X1 #() 
BUF_X1_328_ (
  .A({ din[47] }),
  .Z({ S1[47] })
);
BUF_X1 #() 
BUF_X1_329_ (
  .A({ din[48] }),
  .Z({ S1[48] })
);
BUF_X1 #() 
BUF_X1_330_ (
  .A({ din[49] }),
  .Z({ S1[49] })
);
BUF_X1 #() 
BUF_X1_331_ (
  .A({ din[5] }),
  .Z({ S1[5] })
);
BUF_X1 #() 
BUF_X1_332_ (
  .A({ din[50] }),
  .Z({ S1[50] })
);
BUF_X1 #() 
BUF_X1_333_ (
  .A({ din[51] }),
  .Z({ S1[51] })
);
BUF_X1 #() 
BUF_X1_334_ (
  .A({ din[52] }),
  .Z({ S1[52] })
);
BUF_X1 #() 
BUF_X1_335_ (
  .A({ din[53] }),
  .Z({ S1[53] })
);
BUF_X1 #() 
BUF_X1_336_ (
  .A({ din[54] }),
  .Z({ S1[54] })
);
BUF_X1 #() 
BUF_X1_337_ (
  .A({ din[55] }),
  .Z({ S1[55] })
);
BUF_X1 #() 
BUF_X1_338_ (
  .A({ din[56] }),
  .Z({ S1[56] })
);
BUF_X1 #() 
BUF_X1_339_ (
  .A({ din[57] }),
  .Z({ S1[57] })
);
BUF_X1 #() 
BUF_X1_340_ (
  .A({ din[58] }),
  .Z({ S1[58] })
);
BUF_X1 #() 
BUF_X1_341_ (
  .A({ din[59] }),
  .Z({ S1[59] })
);
BUF_X1 #() 
BUF_X1_342_ (
  .A({ din[6] }),
  .Z({ S1[6] })
);
BUF_X1 #() 
BUF_X1_343_ (
  .A({ din[60] }),
  .Z({ S1[60] })
);
BUF_X1 #() 
BUF_X1_344_ (
  .A({ din[61] }),
  .Z({ S1[61] })
);
BUF_X1 #() 
BUF_X1_345_ (
  .A({ din[62] }),
  .Z({ S1[62] })
);
BUF_X1 #() 
BUF_X1_346_ (
  .A({ din[63] }),
  .Z({ S1[63] })
);
BUF_X1 #() 
BUF_X1_347_ (
  .A({ din[64] }),
  .Z({ S1[64] })
);
BUF_X1 #() 
BUF_X1_348_ (
  .A({ din[65] }),
  .Z({ S1[65] })
);
BUF_X1 #() 
BUF_X1_349_ (
  .A({ din[66] }),
  .Z({ S1[66] })
);
BUF_X1 #() 
BUF_X1_350_ (
  .A({ din[67] }),
  .Z({ S1[67] })
);
BUF_X1 #() 
BUF_X1_351_ (
  .A({ din[68] }),
  .Z({ S1[68] })
);
BUF_X1 #() 
BUF_X1_352_ (
  .A({ din[69] }),
  .Z({ S1[69] })
);
BUF_X1 #() 
BUF_X1_353_ (
  .A({ din[7] }),
  .Z({ S1[7] })
);
BUF_X1 #() 
BUF_X1_354_ (
  .A({ din[70] }),
  .Z({ S1[70] })
);
BUF_X1 #() 
BUF_X1_355_ (
  .A({ din[71] }),
  .Z({ S1[71] })
);
BUF_X1 #() 
BUF_X1_356_ (
  .A({ din[72] }),
  .Z({ S1[72] })
);
BUF_X1 #() 
BUF_X1_357_ (
  .A({ din[73] }),
  .Z({ S1[73] })
);
BUF_X1 #() 
BUF_X1_358_ (
  .A({ din[74] }),
  .Z({ S1[74] })
);
BUF_X1 #() 
BUF_X1_359_ (
  .A({ din[75] }),
  .Z({ S1[75] })
);
BUF_X1 #() 
BUF_X1_360_ (
  .A({ din[76] }),
  .Z({ S1[76] })
);
BUF_X1 #() 
BUF_X1_361_ (
  .A({ din[77] }),
  .Z({ S1[77] })
);
BUF_X1 #() 
BUF_X1_362_ (
  .A({ din[78] }),
  .Z({ S1[78] })
);
BUF_X1 #() 
BUF_X1_363_ (
  .A({ din[79] }),
  .Z({ S1[79] })
);
BUF_X1 #() 
BUF_X1_364_ (
  .A({ din[8] }),
  .Z({ S1[8] })
);
BUF_X1 #() 
BUF_X1_365_ (
  .A({ din[80] }),
  .Z({ S1[80] })
);
BUF_X1 #() 
BUF_X1_366_ (
  .A({ din[81] }),
  .Z({ S1[81] })
);
BUF_X1 #() 
BUF_X1_367_ (
  .A({ din[82] }),
  .Z({ S1[82] })
);
BUF_X1 #() 
BUF_X1_368_ (
  .A({ din[83] }),
  .Z({ S1[83] })
);
BUF_X1 #() 
BUF_X1_369_ (
  .A({ din[84] }),
  .Z({ S1[84] })
);
BUF_X1 #() 
BUF_X1_370_ (
  .A({ din[85] }),
  .Z({ S1[85] })
);
BUF_X1 #() 
BUF_X1_371_ (
  .A({ din[86] }),
  .Z({ S1[86] })
);
BUF_X1 #() 
BUF_X1_372_ (
  .A({ din[87] }),
  .Z({ S1[87] })
);
BUF_X1 #() 
BUF_X1_373_ (
  .A({ din[88] }),
  .Z({ S1[88] })
);
BUF_X1 #() 
BUF_X1_374_ (
  .A({ din[89] }),
  .Z({ S1[89] })
);
BUF_X1 #() 
BUF_X1_375_ (
  .A({ din[9] }),
  .Z({ S1[9] })
);
BUF_X1 #() 
BUF_X1_376_ (
  .A({ din[90] }),
  .Z({ S1[90] })
);
BUF_X1 #() 
BUF_X1_377_ (
  .A({ din[91] }),
  .Z({ S1[91] })
);
BUF_X1 #() 
BUF_X1_378_ (
  .A({ din[92] }),
  .Z({ S1[92] })
);
BUF_X1 #() 
BUF_X1_379_ (
  .A({ din[93] }),
  .Z({ S1[93] })
);
BUF_X1 #() 
BUF_X1_380_ (
  .A({ din[94] }),
  .Z({ S1[94] })
);
BUF_X1 #() 
BUF_X1_381_ (
  .A({ din[95] }),
  .Z({ S1[95] })
);
BUF_X1 #() 
BUF_X1_382_ (
  .A({ din[96] }),
  .Z({ S1[96] })
);
BUF_X1 #() 
BUF_X1_383_ (
  .A({ din[97] }),
  .Z({ S1[97] })
);
BUF_X1 #() 
BUF_X1_384_ (
  .A({ din[98] }),
  .Z({ S1[98] })
);
BUF_X1 #() 
BUF_X1_385_ (
  .A({ din[99] }),
  .Z({ S1[99] })
);
BUF_X1 #() 
BUF_X1_386_ (
  .A({ S2[0] }),
  .Z({ dout[0] })
);
BUF_X1 #() 
BUF_X1_387_ (
  .A({ S2[1] }),
  .Z({ dout[1] })
);
BUF_X1 #() 
BUF_X1_388_ (
  .A({ S2[10] }),
  .Z({ dout[10] })
);
BUF_X1 #() 
BUF_X1_389_ (
  .A({ S2[11] }),
  .Z({ dout[11] })
);
BUF_X1 #() 
BUF_X1_390_ (
  .A({ S2[12] }),
  .Z({ dout[12] })
);
BUF_X1 #() 
BUF_X1_391_ (
  .A({ S2[13] }),
  .Z({ dout[13] })
);
BUF_X1 #() 
BUF_X1_392_ (
  .A({ S2[14] }),
  .Z({ dout[14] })
);
BUF_X1 #() 
BUF_X1_393_ (
  .A({ S2[15] }),
  .Z({ dout[15] })
);
BUF_X1 #() 
BUF_X1_394_ (
  .A({ S2[16] }),
  .Z({ dout[16] })
);
BUF_X1 #() 
BUF_X1_395_ (
  .A({ S2[17] }),
  .Z({ dout[17] })
);
BUF_X1 #() 
BUF_X1_396_ (
  .A({ S2[18] }),
  .Z({ dout[18] })
);
BUF_X1 #() 
BUF_X1_397_ (
  .A({ S2[19] }),
  .Z({ dout[19] })
);
BUF_X1 #() 
BUF_X1_398_ (
  .A({ S2[2] }),
  .Z({ dout[2] })
);
BUF_X1 #() 
BUF_X1_399_ (
  .A({ S2[20] }),
  .Z({ dout[20] })
);
BUF_X1 #() 
BUF_X1_400_ (
  .A({ S2[21] }),
  .Z({ dout[21] })
);
BUF_X1 #() 
BUF_X1_401_ (
  .A({ S2[22] }),
  .Z({ dout[22] })
);
BUF_X1 #() 
BUF_X1_402_ (
  .A({ S2[23] }),
  .Z({ dout[23] })
);
BUF_X1 #() 
BUF_X1_403_ (
  .A({ S2[24] }),
  .Z({ dout[24] })
);
BUF_X1 #() 
BUF_X1_404_ (
  .A({ S2[25] }),
  .Z({ dout[25] })
);
BUF_X1 #() 
BUF_X1_405_ (
  .A({ S2[26] }),
  .Z({ dout[26] })
);
BUF_X1 #() 
BUF_X1_406_ (
  .A({ S2[27] }),
  .Z({ dout[27] })
);
BUF_X1 #() 
BUF_X1_407_ (
  .A({ S2[28] }),
  .Z({ dout[28] })
);
BUF_X1 #() 
BUF_X1_408_ (
  .A({ S2[29] }),
  .Z({ dout[29] })
);
BUF_X1 #() 
BUF_X1_409_ (
  .A({ S2[3] }),
  .Z({ dout[3] })
);
BUF_X1 #() 
BUF_X1_410_ (
  .A({ S2[30] }),
  .Z({ dout[30] })
);
BUF_X1 #() 
BUF_X1_411_ (
  .A({ S2[31] }),
  .Z({ dout[31] })
);
BUF_X1 #() 
BUF_X1_412_ (
  .A({ S2[4] }),
  .Z({ dout[4] })
);
BUF_X1 #() 
BUF_X1_413_ (
  .A({ S2[5] }),
  .Z({ dout[5] })
);
BUF_X1 #() 
BUF_X1_414_ (
  .A({ S2[6] }),
  .Z({ dout[6] })
);
BUF_X1 #() 
BUF_X1_415_ (
  .A({ S2[7] }),
  .Z({ dout[7] })
);
BUF_X1 #() 
BUF_X1_416_ (
  .A({ S2[8] }),
  .Z({ dout[8] })
);
BUF_X1 #() 
BUF_X1_417_ (
  .A({ S2[9] }),
  .Z({ dout[9] })
);
BUF_X1 #() 
BUF_X1_418_ (
  .A({ pause }),
  .Z({ S3 })
);
BUF_X1 #() 
BUF_X1_419_ (
  .A({ S4 }),
  .Z({ reg_out })
);
BUF_X1 #() 
BUF_X1_420_ (
  .A({ rst }),
  .Z({ S5 })
);
BUF_X1 #() 
BUF_X1_421_ (
  .A({ run }),
  .Z({ S6 })
);
BUF_X1 #() 
BUF_X1_422_ (
  .A({ w[0] }),
  .Z({ S7[0] })
);
BUF_X1 #() 
BUF_X1_423_ (
  .A({ w[1] }),
  .Z({ S7[1] })
);
BUF_X1 #() 
BUF_X1_424_ (
  .A({ w[10] }),
  .Z({ S7[10] })
);
BUF_X1 #() 
BUF_X1_425_ (
  .A({ w[100] }),
  .Z({ S7[100] })
);
BUF_X1 #() 
BUF_X1_426_ (
  .A({ w[101] }),
  .Z({ S7[101] })
);
BUF_X1 #() 
BUF_X1_427_ (
  .A({ w[102] }),
  .Z({ S7[102] })
);
BUF_X1 #() 
BUF_X1_428_ (
  .A({ w[103] }),
  .Z({ S7[103] })
);
BUF_X1 #() 
BUF_X1_429_ (
  .A({ w[104] }),
  .Z({ S7[104] })
);
BUF_X1 #() 
BUF_X1_430_ (
  .A({ w[105] }),
  .Z({ S7[105] })
);
BUF_X1 #() 
BUF_X1_431_ (
  .A({ w[106] }),
  .Z({ S7[106] })
);
BUF_X1 #() 
BUF_X1_432_ (
  .A({ w[107] }),
  .Z({ S7[107] })
);
BUF_X1 #() 
BUF_X1_433_ (
  .A({ w[108] }),
  .Z({ S7[108] })
);
BUF_X1 #() 
BUF_X1_434_ (
  .A({ w[109] }),
  .Z({ S7[109] })
);
BUF_X1 #() 
BUF_X1_435_ (
  .A({ w[11] }),
  .Z({ S7[11] })
);
BUF_X1 #() 
BUF_X1_436_ (
  .A({ w[110] }),
  .Z({ S7[110] })
);
BUF_X1 #() 
BUF_X1_437_ (
  .A({ w[111] }),
  .Z({ S7[111] })
);
BUF_X1 #() 
BUF_X1_438_ (
  .A({ w[112] }),
  .Z({ S7[112] })
);
BUF_X1 #() 
BUF_X1_439_ (
  .A({ w[113] }),
  .Z({ S7[113] })
);
BUF_X1 #() 
BUF_X1_440_ (
  .A({ w[114] }),
  .Z({ S7[114] })
);
BUF_X1 #() 
BUF_X1_441_ (
  .A({ w[115] }),
  .Z({ S7[115] })
);
BUF_X1 #() 
BUF_X1_442_ (
  .A({ w[116] }),
  .Z({ S7[116] })
);
BUF_X1 #() 
BUF_X1_443_ (
  .A({ w[117] }),
  .Z({ S7[117] })
);
BUF_X1 #() 
BUF_X1_444_ (
  .A({ w[118] }),
  .Z({ S7[118] })
);
BUF_X1 #() 
BUF_X1_445_ (
  .A({ w[119] }),
  .Z({ S7[119] })
);
BUF_X1 #() 
BUF_X1_446_ (
  .A({ w[12] }),
  .Z({ S7[12] })
);
BUF_X1 #() 
BUF_X1_447_ (
  .A({ w[120] }),
  .Z({ S7[120] })
);
BUF_X1 #() 
BUF_X1_448_ (
  .A({ w[121] }),
  .Z({ S7[121] })
);
BUF_X1 #() 
BUF_X1_449_ (
  .A({ w[122] }),
  .Z({ S7[122] })
);
BUF_X1 #() 
BUF_X1_450_ (
  .A({ w[123] }),
  .Z({ S7[123] })
);
BUF_X1 #() 
BUF_X1_451_ (
  .A({ w[124] }),
  .Z({ S7[124] })
);
BUF_X1 #() 
BUF_X1_452_ (
  .A({ w[125] }),
  .Z({ S7[125] })
);
BUF_X1 #() 
BUF_X1_453_ (
  .A({ w[126] }),
  .Z({ S7[126] })
);
BUF_X1 #() 
BUF_X1_454_ (
  .A({ w[127] }),
  .Z({ S7[127] })
);
BUF_X1 #() 
BUF_X1_455_ (
  .A({ w[128] }),
  .Z({ S7[128] })
);
BUF_X1 #() 
BUF_X1_456_ (
  .A({ w[129] }),
  .Z({ S7[129] })
);
BUF_X1 #() 
BUF_X1_457_ (
  .A({ w[13] }),
  .Z({ S7[13] })
);
BUF_X1 #() 
BUF_X1_458_ (
  .A({ w[130] }),
  .Z({ S7[130] })
);
BUF_X1 #() 
BUF_X1_459_ (
  .A({ w[131] }),
  .Z({ S7[131] })
);
BUF_X1 #() 
BUF_X1_460_ (
  .A({ w[132] }),
  .Z({ S7[132] })
);
BUF_X1 #() 
BUF_X1_461_ (
  .A({ w[133] }),
  .Z({ S7[133] })
);
BUF_X1 #() 
BUF_X1_462_ (
  .A({ w[134] }),
  .Z({ S7[134] })
);
BUF_X1 #() 
BUF_X1_463_ (
  .A({ w[135] }),
  .Z({ S7[135] })
);
BUF_X1 #() 
BUF_X1_464_ (
  .A({ w[136] }),
  .Z({ S7[136] })
);
BUF_X1 #() 
BUF_X1_465_ (
  .A({ w[137] }),
  .Z({ S7[137] })
);
BUF_X1 #() 
BUF_X1_466_ (
  .A({ w[138] }),
  .Z({ S7[138] })
);
BUF_X1 #() 
BUF_X1_467_ (
  .A({ w[139] }),
  .Z({ S7[139] })
);
BUF_X1 #() 
BUF_X1_468_ (
  .A({ w[14] }),
  .Z({ S7[14] })
);
BUF_X1 #() 
BUF_X1_469_ (
  .A({ w[140] }),
  .Z({ S7[140] })
);
BUF_X1 #() 
BUF_X1_470_ (
  .A({ w[141] }),
  .Z({ S7[141] })
);
BUF_X1 #() 
BUF_X1_471_ (
  .A({ w[142] }),
  .Z({ S7[142] })
);
BUF_X1 #() 
BUF_X1_472_ (
  .A({ w[143] }),
  .Z({ S7[143] })
);
BUF_X1 #() 
BUF_X1_473_ (
  .A({ w[144] }),
  .Z({ S7[144] })
);
BUF_X1 #() 
BUF_X1_474_ (
  .A({ w[145] }),
  .Z({ S7[145] })
);
BUF_X1 #() 
BUF_X1_475_ (
  .A({ w[146] }),
  .Z({ S7[146] })
);
BUF_X1 #() 
BUF_X1_476_ (
  .A({ w[147] }),
  .Z({ S7[147] })
);
BUF_X1 #() 
BUF_X1_477_ (
  .A({ w[148] }),
  .Z({ S7[148] })
);
BUF_X1 #() 
BUF_X1_478_ (
  .A({ w[149] }),
  .Z({ S7[149] })
);
BUF_X1 #() 
BUF_X1_479_ (
  .A({ w[15] }),
  .Z({ S7[15] })
);
BUF_X1 #() 
BUF_X1_480_ (
  .A({ w[150] }),
  .Z({ S7[150] })
);
BUF_X1 #() 
BUF_X1_481_ (
  .A({ w[151] }),
  .Z({ S7[151] })
);
BUF_X1 #() 
BUF_X1_482_ (
  .A({ w[152] }),
  .Z({ S7[152] })
);
BUF_X1 #() 
BUF_X1_483_ (
  .A({ w[153] }),
  .Z({ S7[153] })
);
BUF_X1 #() 
BUF_X1_484_ (
  .A({ w[154] }),
  .Z({ S7[154] })
);
BUF_X1 #() 
BUF_X1_485_ (
  .A({ w[155] }),
  .Z({ S7[155] })
);
BUF_X1 #() 
BUF_X1_486_ (
  .A({ w[156] }),
  .Z({ S7[156] })
);
BUF_X1 #() 
BUF_X1_487_ (
  .A({ w[157] }),
  .Z({ S7[157] })
);
BUF_X1 #() 
BUF_X1_488_ (
  .A({ w[158] }),
  .Z({ S7[158] })
);
BUF_X1 #() 
BUF_X1_489_ (
  .A({ w[159] }),
  .Z({ S7[159] })
);
BUF_X1 #() 
BUF_X1_490_ (
  .A({ w[16] }),
  .Z({ S7[16] })
);
BUF_X1 #() 
BUF_X1_491_ (
  .A({ w[160] }),
  .Z({ S7[160] })
);
BUF_X1 #() 
BUF_X1_492_ (
  .A({ w[161] }),
  .Z({ S7[161] })
);
BUF_X1 #() 
BUF_X1_493_ (
  .A({ w[162] }),
  .Z({ S7[162] })
);
BUF_X1 #() 
BUF_X1_494_ (
  .A({ w[163] }),
  .Z({ S7[163] })
);
BUF_X1 #() 
BUF_X1_495_ (
  .A({ w[164] }),
  .Z({ S7[164] })
);
BUF_X1 #() 
BUF_X1_496_ (
  .A({ w[165] }),
  .Z({ S7[165] })
);
BUF_X1 #() 
BUF_X1_497_ (
  .A({ w[166] }),
  .Z({ S7[166] })
);
BUF_X1 #() 
BUF_X1_498_ (
  .A({ w[167] }),
  .Z({ S7[167] })
);
BUF_X1 #() 
BUF_X1_499_ (
  .A({ w[168] }),
  .Z({ S7[168] })
);
BUF_X1 #() 
BUF_X1_500_ (
  .A({ w[169] }),
  .Z({ S7[169] })
);
BUF_X1 #() 
BUF_X1_501_ (
  .A({ w[17] }),
  .Z({ S7[17] })
);
BUF_X1 #() 
BUF_X1_502_ (
  .A({ w[170] }),
  .Z({ S7[170] })
);
BUF_X1 #() 
BUF_X1_503_ (
  .A({ w[171] }),
  .Z({ S7[171] })
);
BUF_X1 #() 
BUF_X1_504_ (
  .A({ w[172] }),
  .Z({ S7[172] })
);
BUF_X1 #() 
BUF_X1_505_ (
  .A({ w[173] }),
  .Z({ S7[173] })
);
BUF_X1 #() 
BUF_X1_506_ (
  .A({ w[174] }),
  .Z({ S7[174] })
);
BUF_X1 #() 
BUF_X1_507_ (
  .A({ w[175] }),
  .Z({ S7[175] })
);
BUF_X1 #() 
BUF_X1_508_ (
  .A({ w[176] }),
  .Z({ S7[176] })
);
BUF_X1 #() 
BUF_X1_509_ (
  .A({ w[177] }),
  .Z({ S7[177] })
);
BUF_X1 #() 
BUF_X1_510_ (
  .A({ w[178] }),
  .Z({ S7[178] })
);
BUF_X1 #() 
BUF_X1_511_ (
  .A({ w[179] }),
  .Z({ S7[179] })
);
BUF_X1 #() 
BUF_X1_512_ (
  .A({ w[18] }),
  .Z({ S7[18] })
);
BUF_X1 #() 
BUF_X1_513_ (
  .A({ w[180] }),
  .Z({ S7[180] })
);
BUF_X1 #() 
BUF_X1_514_ (
  .A({ w[181] }),
  .Z({ S7[181] })
);
BUF_X1 #() 
BUF_X1_515_ (
  .A({ w[182] }),
  .Z({ S7[182] })
);
BUF_X1 #() 
BUF_X1_516_ (
  .A({ w[183] }),
  .Z({ S7[183] })
);
BUF_X1 #() 
BUF_X1_517_ (
  .A({ w[184] }),
  .Z({ S7[184] })
);
BUF_X1 #() 
BUF_X1_518_ (
  .A({ w[185] }),
  .Z({ S7[185] })
);
BUF_X1 #() 
BUF_X1_519_ (
  .A({ w[186] }),
  .Z({ S7[186] })
);
BUF_X1 #() 
BUF_X1_520_ (
  .A({ w[187] }),
  .Z({ S7[187] })
);
BUF_X1 #() 
BUF_X1_521_ (
  .A({ w[188] }),
  .Z({ S7[188] })
);
BUF_X1 #() 
BUF_X1_522_ (
  .A({ w[189] }),
  .Z({ S7[189] })
);
BUF_X1 #() 
BUF_X1_523_ (
  .A({ w[19] }),
  .Z({ S7[19] })
);
BUF_X1 #() 
BUF_X1_524_ (
  .A({ w[190] }),
  .Z({ S7[190] })
);
BUF_X1 #() 
BUF_X1_525_ (
  .A({ w[191] }),
  .Z({ S7[191] })
);
BUF_X1 #() 
BUF_X1_526_ (
  .A({ w[192] }),
  .Z({ S7[192] })
);
BUF_X1 #() 
BUF_X1_527_ (
  .A({ w[193] }),
  .Z({ S7[193] })
);
BUF_X1 #() 
BUF_X1_528_ (
  .A({ w[194] }),
  .Z({ S7[194] })
);
BUF_X1 #() 
BUF_X1_529_ (
  .A({ w[195] }),
  .Z({ S7[195] })
);
BUF_X1 #() 
BUF_X1_530_ (
  .A({ w[196] }),
  .Z({ S7[196] })
);
BUF_X1 #() 
BUF_X1_531_ (
  .A({ w[197] }),
  .Z({ S7[197] })
);
BUF_X1 #() 
BUF_X1_532_ (
  .A({ w[198] }),
  .Z({ S7[198] })
);
BUF_X1 #() 
BUF_X1_533_ (
  .A({ w[199] }),
  .Z({ S7[199] })
);
BUF_X1 #() 
BUF_X1_534_ (
  .A({ w[2] }),
  .Z({ S7[2] })
);
BUF_X1 #() 
BUF_X1_535_ (
  .A({ w[20] }),
  .Z({ S7[20] })
);
BUF_X1 #() 
BUF_X1_536_ (
  .A({ w[200] }),
  .Z({ S7[200] })
);
BUF_X1 #() 
BUF_X1_537_ (
  .A({ w[201] }),
  .Z({ S7[201] })
);
BUF_X1 #() 
BUF_X1_538_ (
  .A({ w[202] }),
  .Z({ S7[202] })
);
BUF_X1 #() 
BUF_X1_539_ (
  .A({ w[203] }),
  .Z({ S7[203] })
);
BUF_X1 #() 
BUF_X1_540_ (
  .A({ w[204] }),
  .Z({ S7[204] })
);
BUF_X1 #() 
BUF_X1_541_ (
  .A({ w[205] }),
  .Z({ S7[205] })
);
BUF_X1 #() 
BUF_X1_542_ (
  .A({ w[206] }),
  .Z({ S7[206] })
);
BUF_X1 #() 
BUF_X1_543_ (
  .A({ w[207] }),
  .Z({ S7[207] })
);
BUF_X1 #() 
BUF_X1_544_ (
  .A({ w[208] }),
  .Z({ S7[208] })
);
BUF_X1 #() 
BUF_X1_545_ (
  .A({ w[209] }),
  .Z({ S7[209] })
);
BUF_X1 #() 
BUF_X1_546_ (
  .A({ w[21] }),
  .Z({ S7[21] })
);
BUF_X1 #() 
BUF_X1_547_ (
  .A({ w[210] }),
  .Z({ S7[210] })
);
BUF_X1 #() 
BUF_X1_548_ (
  .A({ w[211] }),
  .Z({ S7[211] })
);
BUF_X1 #() 
BUF_X1_549_ (
  .A({ w[212] }),
  .Z({ S7[212] })
);
BUF_X1 #() 
BUF_X1_550_ (
  .A({ w[213] }),
  .Z({ S7[213] })
);
BUF_X1 #() 
BUF_X1_551_ (
  .A({ w[214] }),
  .Z({ S7[214] })
);
BUF_X1 #() 
BUF_X1_552_ (
  .A({ w[215] }),
  .Z({ S7[215] })
);
BUF_X1 #() 
BUF_X1_553_ (
  .A({ w[216] }),
  .Z({ S7[216] })
);
BUF_X1 #() 
BUF_X1_554_ (
  .A({ w[217] }),
  .Z({ S7[217] })
);
BUF_X1 #() 
BUF_X1_555_ (
  .A({ w[218] }),
  .Z({ S7[218] })
);
BUF_X1 #() 
BUF_X1_556_ (
  .A({ w[219] }),
  .Z({ S7[219] })
);
BUF_X1 #() 
BUF_X1_557_ (
  .A({ w[22] }),
  .Z({ S7[22] })
);
BUF_X1 #() 
BUF_X1_558_ (
  .A({ w[220] }),
  .Z({ S7[220] })
);
BUF_X1 #() 
BUF_X1_559_ (
  .A({ w[221] }),
  .Z({ S7[221] })
);
BUF_X1 #() 
BUF_X1_560_ (
  .A({ w[222] }),
  .Z({ S7[222] })
);
BUF_X1 #() 
BUF_X1_561_ (
  .A({ w[223] }),
  .Z({ S7[223] })
);
BUF_X1 #() 
BUF_X1_562_ (
  .A({ w[224] }),
  .Z({ S7[224] })
);
BUF_X1 #() 
BUF_X1_563_ (
  .A({ w[225] }),
  .Z({ S7[225] })
);
BUF_X1 #() 
BUF_X1_564_ (
  .A({ w[226] }),
  .Z({ S7[226] })
);
BUF_X1 #() 
BUF_X1_565_ (
  .A({ w[227] }),
  .Z({ S7[227] })
);
BUF_X1 #() 
BUF_X1_566_ (
  .A({ w[228] }),
  .Z({ S7[228] })
);
BUF_X1 #() 
BUF_X1_567_ (
  .A({ w[229] }),
  .Z({ S7[229] })
);
BUF_X1 #() 
BUF_X1_568_ (
  .A({ w[23] }),
  .Z({ S7[23] })
);
BUF_X1 #() 
BUF_X1_569_ (
  .A({ w[230] }),
  .Z({ S7[230] })
);
BUF_X1 #() 
BUF_X1_570_ (
  .A({ w[231] }),
  .Z({ S7[231] })
);
BUF_X1 #() 
BUF_X1_571_ (
  .A({ w[232] }),
  .Z({ S7[232] })
);
BUF_X1 #() 
BUF_X1_572_ (
  .A({ w[233] }),
  .Z({ S7[233] })
);
BUF_X1 #() 
BUF_X1_573_ (
  .A({ w[234] }),
  .Z({ S7[234] })
);
BUF_X1 #() 
BUF_X1_574_ (
  .A({ w[235] }),
  .Z({ S7[235] })
);
BUF_X1 #() 
BUF_X1_575_ (
  .A({ w[236] }),
  .Z({ S7[236] })
);
BUF_X1 #() 
BUF_X1_576_ (
  .A({ w[237] }),
  .Z({ S7[237] })
);
BUF_X1 #() 
BUF_X1_577_ (
  .A({ w[238] }),
  .Z({ S7[238] })
);
BUF_X1 #() 
BUF_X1_578_ (
  .A({ w[239] }),
  .Z({ S7[239] })
);
BUF_X1 #() 
BUF_X1_579_ (
  .A({ w[24] }),
  .Z({ S7[24] })
);
BUF_X1 #() 
BUF_X1_580_ (
  .A({ w[240] }),
  .Z({ S7[240] })
);
BUF_X1 #() 
BUF_X1_581_ (
  .A({ w[241] }),
  .Z({ S7[241] })
);
BUF_X1 #() 
BUF_X1_582_ (
  .A({ w[242] }),
  .Z({ S7[242] })
);
BUF_X1 #() 
BUF_X1_583_ (
  .A({ w[243] }),
  .Z({ S7[243] })
);
BUF_X1 #() 
BUF_X1_584_ (
  .A({ w[244] }),
  .Z({ S7[244] })
);
BUF_X1 #() 
BUF_X1_585_ (
  .A({ w[245] }),
  .Z({ S7[245] })
);
BUF_X1 #() 
BUF_X1_586_ (
  .A({ w[246] }),
  .Z({ S7[246] })
);
BUF_X1 #() 
BUF_X1_587_ (
  .A({ w[247] }),
  .Z({ S7[247] })
);
BUF_X1 #() 
BUF_X1_588_ (
  .A({ w[248] }),
  .Z({ S7[248] })
);
BUF_X1 #() 
BUF_X1_589_ (
  .A({ w[249] }),
  .Z({ S7[249] })
);
BUF_X1 #() 
BUF_X1_590_ (
  .A({ w[25] }),
  .Z({ S7[25] })
);
BUF_X1 #() 
BUF_X1_591_ (
  .A({ w[250] }),
  .Z({ S7[250] })
);
BUF_X1 #() 
BUF_X1_592_ (
  .A({ w[251] }),
  .Z({ S7[251] })
);
BUF_X1 #() 
BUF_X1_593_ (
  .A({ w[252] }),
  .Z({ S7[252] })
);
BUF_X1 #() 
BUF_X1_594_ (
  .A({ w[253] }),
  .Z({ S7[253] })
);
BUF_X1 #() 
BUF_X1_595_ (
  .A({ w[254] }),
  .Z({ S7[254] })
);
BUF_X1 #() 
BUF_X1_596_ (
  .A({ w[255] }),
  .Z({ S7[255] })
);
BUF_X1 #() 
BUF_X1_597_ (
  .A({ w[256] }),
  .Z({ S7[256] })
);
BUF_X1 #() 
BUF_X1_598_ (
  .A({ w[257] }),
  .Z({ S7[257] })
);
BUF_X1 #() 
BUF_X1_599_ (
  .A({ w[258] }),
  .Z({ S7[258] })
);
BUF_X1 #() 
BUF_X1_600_ (
  .A({ w[259] }),
  .Z({ S7[259] })
);
BUF_X1 #() 
BUF_X1_601_ (
  .A({ w[26] }),
  .Z({ S7[26] })
);
BUF_X1 #() 
BUF_X1_602_ (
  .A({ w[260] }),
  .Z({ S7[260] })
);
BUF_X1 #() 
BUF_X1_603_ (
  .A({ w[261] }),
  .Z({ S7[261] })
);
BUF_X1 #() 
BUF_X1_604_ (
  .A({ w[262] }),
  .Z({ S7[262] })
);
BUF_X1 #() 
BUF_X1_605_ (
  .A({ w[263] }),
  .Z({ S7[263] })
);
BUF_X1 #() 
BUF_X1_606_ (
  .A({ w[264] }),
  .Z({ S7[264] })
);
BUF_X1 #() 
BUF_X1_607_ (
  .A({ w[265] }),
  .Z({ S7[265] })
);
BUF_X1 #() 
BUF_X1_608_ (
  .A({ w[266] }),
  .Z({ S7[266] })
);
BUF_X1 #() 
BUF_X1_609_ (
  .A({ w[267] }),
  .Z({ S7[267] })
);
BUF_X1 #() 
BUF_X1_610_ (
  .A({ w[268] }),
  .Z({ S7[268] })
);
BUF_X1 #() 
BUF_X1_611_ (
  .A({ w[269] }),
  .Z({ S7[269] })
);
BUF_X1 #() 
BUF_X1_612_ (
  .A({ w[27] }),
  .Z({ S7[27] })
);
BUF_X1 #() 
BUF_X1_613_ (
  .A({ w[270] }),
  .Z({ S7[270] })
);
BUF_X1 #() 
BUF_X1_614_ (
  .A({ w[271] }),
  .Z({ S7[271] })
);
BUF_X1 #() 
BUF_X1_615_ (
  .A({ w[272] }),
  .Z({ S7[272] })
);
BUF_X1 #() 
BUF_X1_616_ (
  .A({ w[273] }),
  .Z({ S7[273] })
);
BUF_X1 #() 
BUF_X1_617_ (
  .A({ w[274] }),
  .Z({ S7[274] })
);
BUF_X1 #() 
BUF_X1_618_ (
  .A({ w[275] }),
  .Z({ S7[275] })
);
BUF_X1 #() 
BUF_X1_619_ (
  .A({ w[276] }),
  .Z({ S7[276] })
);
BUF_X1 #() 
BUF_X1_620_ (
  .A({ w[277] }),
  .Z({ S7[277] })
);
BUF_X1 #() 
BUF_X1_621_ (
  .A({ w[278] }),
  .Z({ S7[278] })
);
BUF_X1 #() 
BUF_X1_622_ (
  .A({ w[279] }),
  .Z({ S7[279] })
);
BUF_X1 #() 
BUF_X1_623_ (
  .A({ w[28] }),
  .Z({ S7[28] })
);
BUF_X1 #() 
BUF_X1_624_ (
  .A({ w[280] }),
  .Z({ S7[280] })
);
BUF_X1 #() 
BUF_X1_625_ (
  .A({ w[281] }),
  .Z({ S7[281] })
);
BUF_X1 #() 
BUF_X1_626_ (
  .A({ w[282] }),
  .Z({ S7[282] })
);
BUF_X1 #() 
BUF_X1_627_ (
  .A({ w[283] }),
  .Z({ S7[283] })
);
BUF_X1 #() 
BUF_X1_628_ (
  .A({ w[284] }),
  .Z({ S7[284] })
);
BUF_X1 #() 
BUF_X1_629_ (
  .A({ w[285] }),
  .Z({ S7[285] })
);
BUF_X1 #() 
BUF_X1_630_ (
  .A({ w[286] }),
  .Z({ S7[286] })
);
BUF_X1 #() 
BUF_X1_631_ (
  .A({ w[287] }),
  .Z({ S7[287] })
);
BUF_X1 #() 
BUF_X1_632_ (
  .A({ w[288] }),
  .Z({ S7[288] })
);
BUF_X1 #() 
BUF_X1_633_ (
  .A({ w[289] }),
  .Z({ S7[289] })
);
BUF_X1 #() 
BUF_X1_634_ (
  .A({ w[29] }),
  .Z({ S7[29] })
);
BUF_X1 #() 
BUF_X1_635_ (
  .A({ w[290] }),
  .Z({ S7[290] })
);
BUF_X1 #() 
BUF_X1_636_ (
  .A({ w[291] }),
  .Z({ S7[291] })
);
BUF_X1 #() 
BUF_X1_637_ (
  .A({ w[292] }),
  .Z({ S7[292] })
);
BUF_X1 #() 
BUF_X1_638_ (
  .A({ w[293] }),
  .Z({ S7[293] })
);
BUF_X1 #() 
BUF_X1_639_ (
  .A({ w[294] }),
  .Z({ S7[294] })
);
BUF_X1 #() 
BUF_X1_640_ (
  .A({ w[295] }),
  .Z({ S7[295] })
);
BUF_X1 #() 
BUF_X1_641_ (
  .A({ w[296] }),
  .Z({ S7[296] })
);
BUF_X1 #() 
BUF_X1_642_ (
  .A({ w[297] }),
  .Z({ S7[297] })
);
BUF_X1 #() 
BUF_X1_643_ (
  .A({ w[298] }),
  .Z({ S7[298] })
);
BUF_X1 #() 
BUF_X1_644_ (
  .A({ w[299] }),
  .Z({ S7[299] })
);
BUF_X1 #() 
BUF_X1_645_ (
  .A({ w[3] }),
  .Z({ S7[3] })
);
BUF_X1 #() 
BUF_X1_646_ (
  .A({ w[30] }),
  .Z({ S7[30] })
);
BUF_X1 #() 
BUF_X1_647_ (
  .A({ w[300] }),
  .Z({ S7[300] })
);
BUF_X1 #() 
BUF_X1_648_ (
  .A({ w[301] }),
  .Z({ S7[301] })
);
BUF_X1 #() 
BUF_X1_649_ (
  .A({ w[302] }),
  .Z({ S7[302] })
);
BUF_X1 #() 
BUF_X1_650_ (
  .A({ w[303] }),
  .Z({ S7[303] })
);
BUF_X1 #() 
BUF_X1_651_ (
  .A({ w[304] }),
  .Z({ S7[304] })
);
BUF_X1 #() 
BUF_X1_652_ (
  .A({ w[305] }),
  .Z({ S7[305] })
);
BUF_X1 #() 
BUF_X1_653_ (
  .A({ w[306] }),
  .Z({ S7[306] })
);
BUF_X1 #() 
BUF_X1_654_ (
  .A({ w[307] }),
  .Z({ S7[307] })
);
BUF_X1 #() 
BUF_X1_655_ (
  .A({ w[308] }),
  .Z({ S7[308] })
);
BUF_X1 #() 
BUF_X1_656_ (
  .A({ w[309] }),
  .Z({ S7[309] })
);
BUF_X1 #() 
BUF_X1_657_ (
  .A({ w[31] }),
  .Z({ S7[31] })
);
BUF_X1 #() 
BUF_X1_658_ (
  .A({ w[310] }),
  .Z({ S7[310] })
);
BUF_X1 #() 
BUF_X1_659_ (
  .A({ w[311] }),
  .Z({ S7[311] })
);
BUF_X1 #() 
BUF_X1_660_ (
  .A({ w[312] }),
  .Z({ S7[312] })
);
BUF_X1 #() 
BUF_X1_661_ (
  .A({ w[313] }),
  .Z({ S7[313] })
);
BUF_X1 #() 
BUF_X1_662_ (
  .A({ w[314] }),
  .Z({ S7[314] })
);
BUF_X1 #() 
BUF_X1_663_ (
  .A({ w[315] }),
  .Z({ S7[315] })
);
BUF_X1 #() 
BUF_X1_664_ (
  .A({ w[316] }),
  .Z({ S7[316] })
);
BUF_X1 #() 
BUF_X1_665_ (
  .A({ w[317] }),
  .Z({ S7[317] })
);
BUF_X1 #() 
BUF_X1_666_ (
  .A({ w[318] }),
  .Z({ S7[318] })
);
BUF_X1 #() 
BUF_X1_667_ (
  .A({ w[319] }),
  .Z({ S7[319] })
);
BUF_X1 #() 
BUF_X1_668_ (
  .A({ w[32] }),
  .Z({ S7[32] })
);
BUF_X1 #() 
BUF_X1_669_ (
  .A({ w[320] }),
  .Z({ S7[320] })
);
BUF_X1 #() 
BUF_X1_670_ (
  .A({ w[321] }),
  .Z({ S7[321] })
);
BUF_X1 #() 
BUF_X1_671_ (
  .A({ w[322] }),
  .Z({ S7[322] })
);
BUF_X1 #() 
BUF_X1_672_ (
  .A({ w[323] }),
  .Z({ S7[323] })
);
BUF_X1 #() 
BUF_X1_673_ (
  .A({ w[324] }),
  .Z({ S7[324] })
);
BUF_X1 #() 
BUF_X1_674_ (
  .A({ w[325] }),
  .Z({ S7[325] })
);
BUF_X1 #() 
BUF_X1_675_ (
  .A({ w[326] }),
  .Z({ S7[326] })
);
BUF_X1 #() 
BUF_X1_676_ (
  .A({ w[327] }),
  .Z({ S7[327] })
);
BUF_X1 #() 
BUF_X1_677_ (
  .A({ w[328] }),
  .Z({ S7[328] })
);
BUF_X1 #() 
BUF_X1_678_ (
  .A({ w[329] }),
  .Z({ S7[329] })
);
BUF_X1 #() 
BUF_X1_679_ (
  .A({ w[33] }),
  .Z({ S7[33] })
);
BUF_X1 #() 
BUF_X1_680_ (
  .A({ w[330] }),
  .Z({ S7[330] })
);
BUF_X1 #() 
BUF_X1_681_ (
  .A({ w[331] }),
  .Z({ S7[331] })
);
BUF_X1 #() 
BUF_X1_682_ (
  .A({ w[332] }),
  .Z({ S7[332] })
);
BUF_X1 #() 
BUF_X1_683_ (
  .A({ w[333] }),
  .Z({ S7[333] })
);
BUF_X1 #() 
BUF_X1_684_ (
  .A({ w[334] }),
  .Z({ S7[334] })
);
BUF_X1 #() 
BUF_X1_685_ (
  .A({ w[335] }),
  .Z({ S7[335] })
);
BUF_X1 #() 
BUF_X1_686_ (
  .A({ w[336] }),
  .Z({ S7[336] })
);
BUF_X1 #() 
BUF_X1_687_ (
  .A({ w[337] }),
  .Z({ S7[337] })
);
BUF_X1 #() 
BUF_X1_688_ (
  .A({ w[338] }),
  .Z({ S7[338] })
);
BUF_X1 #() 
BUF_X1_689_ (
  .A({ w[339] }),
  .Z({ S7[339] })
);
BUF_X1 #() 
BUF_X1_690_ (
  .A({ w[34] }),
  .Z({ S7[34] })
);
BUF_X1 #() 
BUF_X1_691_ (
  .A({ w[340] }),
  .Z({ S7[340] })
);
BUF_X1 #() 
BUF_X1_692_ (
  .A({ w[341] }),
  .Z({ S7[341] })
);
BUF_X1 #() 
BUF_X1_693_ (
  .A({ w[342] }),
  .Z({ S7[342] })
);
BUF_X1 #() 
BUF_X1_694_ (
  .A({ w[343] }),
  .Z({ S7[343] })
);
BUF_X1 #() 
BUF_X1_695_ (
  .A({ w[344] }),
  .Z({ S7[344] })
);
BUF_X1 #() 
BUF_X1_696_ (
  .A({ w[345] }),
  .Z({ S7[345] })
);
BUF_X1 #() 
BUF_X1_697_ (
  .A({ w[346] }),
  .Z({ S7[346] })
);
BUF_X1 #() 
BUF_X1_698_ (
  .A({ w[347] }),
  .Z({ S7[347] })
);
BUF_X1 #() 
BUF_X1_699_ (
  .A({ w[348] }),
  .Z({ S7[348] })
);
BUF_X1 #() 
BUF_X1_700_ (
  .A({ w[349] }),
  .Z({ S7[349] })
);
BUF_X1 #() 
BUF_X1_701_ (
  .A({ w[35] }),
  .Z({ S7[35] })
);
BUF_X1 #() 
BUF_X1_702_ (
  .A({ w[350] }),
  .Z({ S7[350] })
);
BUF_X1 #() 
BUF_X1_703_ (
  .A({ w[351] }),
  .Z({ S7[351] })
);
BUF_X1 #() 
BUF_X1_704_ (
  .A({ w[352] }),
  .Z({ S7[352] })
);
BUF_X1 #() 
BUF_X1_705_ (
  .A({ w[353] }),
  .Z({ S7[353] })
);
BUF_X1 #() 
BUF_X1_706_ (
  .A({ w[354] }),
  .Z({ S7[354] })
);
BUF_X1 #() 
BUF_X1_707_ (
  .A({ w[355] }),
  .Z({ S7[355] })
);
BUF_X1 #() 
BUF_X1_708_ (
  .A({ w[356] }),
  .Z({ S7[356] })
);
BUF_X1 #() 
BUF_X1_709_ (
  .A({ w[357] }),
  .Z({ S7[357] })
);
BUF_X1 #() 
BUF_X1_710_ (
  .A({ w[358] }),
  .Z({ S7[358] })
);
BUF_X1 #() 
BUF_X1_711_ (
  .A({ w[359] }),
  .Z({ S7[359] })
);
BUF_X1 #() 
BUF_X1_712_ (
  .A({ w[36] }),
  .Z({ S7[36] })
);
BUF_X1 #() 
BUF_X1_713_ (
  .A({ w[360] }),
  .Z({ S7[360] })
);
BUF_X1 #() 
BUF_X1_714_ (
  .A({ w[361] }),
  .Z({ S7[361] })
);
BUF_X1 #() 
BUF_X1_715_ (
  .A({ w[362] }),
  .Z({ S7[362] })
);
BUF_X1 #() 
BUF_X1_716_ (
  .A({ w[363] }),
  .Z({ S7[363] })
);
BUF_X1 #() 
BUF_X1_717_ (
  .A({ w[364] }),
  .Z({ S7[364] })
);
BUF_X1 #() 
BUF_X1_718_ (
  .A({ w[365] }),
  .Z({ S7[365] })
);
BUF_X1 #() 
BUF_X1_719_ (
  .A({ w[366] }),
  .Z({ S7[366] })
);
BUF_X1 #() 
BUF_X1_720_ (
  .A({ w[367] }),
  .Z({ S7[367] })
);
BUF_X1 #() 
BUF_X1_721_ (
  .A({ w[368] }),
  .Z({ S7[368] })
);
BUF_X1 #() 
BUF_X1_722_ (
  .A({ w[369] }),
  .Z({ S7[369] })
);
BUF_X1 #() 
BUF_X1_723_ (
  .A({ w[37] }),
  .Z({ S7[37] })
);
BUF_X1 #() 
BUF_X1_724_ (
  .A({ w[370] }),
  .Z({ S7[370] })
);
BUF_X1 #() 
BUF_X1_725_ (
  .A({ w[371] }),
  .Z({ S7[371] })
);
BUF_X1 #() 
BUF_X1_726_ (
  .A({ w[372] }),
  .Z({ S7[372] })
);
BUF_X1 #() 
BUF_X1_727_ (
  .A({ w[373] }),
  .Z({ S7[373] })
);
BUF_X1 #() 
BUF_X1_728_ (
  .A({ w[374] }),
  .Z({ S7[374] })
);
BUF_X1 #() 
BUF_X1_729_ (
  .A({ w[375] }),
  .Z({ S7[375] })
);
BUF_X1 #() 
BUF_X1_730_ (
  .A({ w[376] }),
  .Z({ S7[376] })
);
BUF_X1 #() 
BUF_X1_731_ (
  .A({ w[377] }),
  .Z({ S7[377] })
);
BUF_X1 #() 
BUF_X1_732_ (
  .A({ w[378] }),
  .Z({ S7[378] })
);
BUF_X1 #() 
BUF_X1_733_ (
  .A({ w[379] }),
  .Z({ S7[379] })
);
BUF_X1 #() 
BUF_X1_734_ (
  .A({ w[38] }),
  .Z({ S7[38] })
);
BUF_X1 #() 
BUF_X1_735_ (
  .A({ w[380] }),
  .Z({ S7[380] })
);
BUF_X1 #() 
BUF_X1_736_ (
  .A({ w[381] }),
  .Z({ S7[381] })
);
BUF_X1 #() 
BUF_X1_737_ (
  .A({ w[382] }),
  .Z({ S7[382] })
);
BUF_X1 #() 
BUF_X1_738_ (
  .A({ w[383] }),
  .Z({ S7[383] })
);
BUF_X1 #() 
BUF_X1_739_ (
  .A({ w[39] }),
  .Z({ S7[39] })
);
BUF_X1 #() 
BUF_X1_740_ (
  .A({ w[4] }),
  .Z({ S7[4] })
);
BUF_X1 #() 
BUF_X1_741_ (
  .A({ w[40] }),
  .Z({ S7[40] })
);
BUF_X1 #() 
BUF_X1_742_ (
  .A({ w[41] }),
  .Z({ S7[41] })
);
BUF_X1 #() 
BUF_X1_743_ (
  .A({ w[42] }),
  .Z({ S7[42] })
);
BUF_X1 #() 
BUF_X1_744_ (
  .A({ w[43] }),
  .Z({ S7[43] })
);
BUF_X1 #() 
BUF_X1_745_ (
  .A({ w[44] }),
  .Z({ S7[44] })
);
BUF_X1 #() 
BUF_X1_746_ (
  .A({ w[45] }),
  .Z({ S7[45] })
);
BUF_X1 #() 
BUF_X1_747_ (
  .A({ w[46] }),
  .Z({ S7[46] })
);
BUF_X1 #() 
BUF_X1_748_ (
  .A({ w[47] }),
  .Z({ S7[47] })
);
BUF_X1 #() 
BUF_X1_749_ (
  .A({ w[48] }),
  .Z({ S7[48] })
);
BUF_X1 #() 
BUF_X1_750_ (
  .A({ w[49] }),
  .Z({ S7[49] })
);
BUF_X1 #() 
BUF_X1_751_ (
  .A({ w[5] }),
  .Z({ S7[5] })
);
BUF_X1 #() 
BUF_X1_752_ (
  .A({ w[50] }),
  .Z({ S7[50] })
);
BUF_X1 #() 
BUF_X1_753_ (
  .A({ w[51] }),
  .Z({ S7[51] })
);
BUF_X1 #() 
BUF_X1_754_ (
  .A({ w[52] }),
  .Z({ S7[52] })
);
BUF_X1 #() 
BUF_X1_755_ (
  .A({ w[53] }),
  .Z({ S7[53] })
);
BUF_X1 #() 
BUF_X1_756_ (
  .A({ w[54] }),
  .Z({ S7[54] })
);
BUF_X1 #() 
BUF_X1_757_ (
  .A({ w[55] }),
  .Z({ S7[55] })
);
BUF_X1 #() 
BUF_X1_758_ (
  .A({ w[56] }),
  .Z({ S7[56] })
);
BUF_X1 #() 
BUF_X1_759_ (
  .A({ w[57] }),
  .Z({ S7[57] })
);
BUF_X1 #() 
BUF_X1_760_ (
  .A({ w[58] }),
  .Z({ S7[58] })
);
BUF_X1 #() 
BUF_X1_761_ (
  .A({ w[59] }),
  .Z({ S7[59] })
);
BUF_X1 #() 
BUF_X1_762_ (
  .A({ w[6] }),
  .Z({ S7[6] })
);
BUF_X1 #() 
BUF_X1_763_ (
  .A({ w[60] }),
  .Z({ S7[60] })
);
BUF_X1 #() 
BUF_X1_764_ (
  .A({ w[61] }),
  .Z({ S7[61] })
);
BUF_X1 #() 
BUF_X1_765_ (
  .A({ w[62] }),
  .Z({ S7[62] })
);
BUF_X1 #() 
BUF_X1_766_ (
  .A({ w[63] }),
  .Z({ S7[63] })
);
BUF_X1 #() 
BUF_X1_767_ (
  .A({ w[64] }),
  .Z({ S7[64] })
);
BUF_X1 #() 
BUF_X1_768_ (
  .A({ w[65] }),
  .Z({ S7[65] })
);
BUF_X1 #() 
BUF_X1_769_ (
  .A({ w[66] }),
  .Z({ S7[66] })
);
BUF_X1 #() 
BUF_X1_770_ (
  .A({ w[67] }),
  .Z({ S7[67] })
);
BUF_X1 #() 
BUF_X1_771_ (
  .A({ w[68] }),
  .Z({ S7[68] })
);
BUF_X1 #() 
BUF_X1_772_ (
  .A({ w[69] }),
  .Z({ S7[69] })
);
BUF_X1 #() 
BUF_X1_773_ (
  .A({ w[7] }),
  .Z({ S7[7] })
);
BUF_X1 #() 
BUF_X1_774_ (
  .A({ w[70] }),
  .Z({ S7[70] })
);
BUF_X1 #() 
BUF_X1_775_ (
  .A({ w[71] }),
  .Z({ S7[71] })
);
BUF_X1 #() 
BUF_X1_776_ (
  .A({ w[72] }),
  .Z({ S7[72] })
);
BUF_X1 #() 
BUF_X1_777_ (
  .A({ w[73] }),
  .Z({ S7[73] })
);
BUF_X1 #() 
BUF_X1_778_ (
  .A({ w[74] }),
  .Z({ S7[74] })
);
BUF_X1 #() 
BUF_X1_779_ (
  .A({ w[75] }),
  .Z({ S7[75] })
);
BUF_X1 #() 
BUF_X1_780_ (
  .A({ w[76] }),
  .Z({ S7[76] })
);
BUF_X1 #() 
BUF_X1_781_ (
  .A({ w[77] }),
  .Z({ S7[77] })
);
BUF_X1 #() 
BUF_X1_782_ (
  .A({ w[78] }),
  .Z({ S7[78] })
);
BUF_X1 #() 
BUF_X1_783_ (
  .A({ w[79] }),
  .Z({ S7[79] })
);
BUF_X1 #() 
BUF_X1_784_ (
  .A({ w[8] }),
  .Z({ S7[8] })
);
BUF_X1 #() 
BUF_X1_785_ (
  .A({ w[80] }),
  .Z({ S7[80] })
);
BUF_X1 #() 
BUF_X1_786_ (
  .A({ w[81] }),
  .Z({ S7[81] })
);
BUF_X1 #() 
BUF_X1_787_ (
  .A({ w[82] }),
  .Z({ S7[82] })
);
BUF_X1 #() 
BUF_X1_788_ (
  .A({ w[83] }),
  .Z({ S7[83] })
);
BUF_X1 #() 
BUF_X1_789_ (
  .A({ w[84] }),
  .Z({ S7[84] })
);
BUF_X1 #() 
BUF_X1_790_ (
  .A({ w[85] }),
  .Z({ S7[85] })
);
BUF_X1 #() 
BUF_X1_791_ (
  .A({ w[86] }),
  .Z({ S7[86] })
);
BUF_X1 #() 
BUF_X1_792_ (
  .A({ w[87] }),
  .Z({ S7[87] })
);
BUF_X1 #() 
BUF_X1_793_ (
  .A({ w[88] }),
  .Z({ S7[88] })
);
BUF_X1 #() 
BUF_X1_794_ (
  .A({ w[89] }),
  .Z({ S7[89] })
);
BUF_X1 #() 
BUF_X1_795_ (
  .A({ w[9] }),
  .Z({ S7[9] })
);
BUF_X1 #() 
BUF_X1_796_ (
  .A({ w[90] }),
  .Z({ S7[90] })
);
BUF_X1 #() 
BUF_X1_797_ (
  .A({ w[91] }),
  .Z({ S7[91] })
);
BUF_X1 #() 
BUF_X1_798_ (
  .A({ w[92] }),
  .Z({ S7[92] })
);
BUF_X1 #() 
BUF_X1_799_ (
  .A({ w[93] }),
  .Z({ S7[93] })
);
BUF_X1 #() 
BUF_X1_800_ (
  .A({ w[94] }),
  .Z({ S7[94] })
);
BUF_X1 #() 
BUF_X1_801_ (
  .A({ w[95] }),
  .Z({ S7[95] })
);
BUF_X1 #() 
BUF_X1_802_ (
  .A({ w[96] }),
  .Z({ S7[96] })
);
BUF_X1 #() 
BUF_X1_803_ (
  .A({ w[97] }),
  .Z({ S7[97] })
);
BUF_X1 #() 
BUF_X1_804_ (
  .A({ w[98] }),
  .Z({ S7[98] })
);
BUF_X1 #() 
BUF_X1_805_ (
  .A({ w[99] }),
  .Z({ S7[99] })
);
convergence_accumulator_plate_4 #() 
convergence_accumulator_plate_4_1_ (
  .clk({ S0 }),
  .din({ data_out_map_0, data_out_map_1, data_out_map_2, data_out_map_3, data_out_map_4, data_out_map_5, data_out_map_6, data_out_map_7, data_out_map_8, data_out_map_9, data_out_map_10, data_out_map_11, data_out_map_12, data_out_map_13, data_out_map_14, data_out_map_15, data_out_map_16, data_out_map_17, data_out_map_18, data_out_map_19, data_out_map_20, data_out_map_21, data_out_map_22, data_out_map_23, data_out_map_24, data_out_map_25, data_out_map_26, data_out_map_27, data_out_map_28, data_out_map_29, data_out_map_30, data_out_map_31, data_out_map_32, data_out_map_33, data_out_map_34, data_out_map_35, data_out_map_36, data_out_map_37, data_out_map_38, data_out_map_39, data_out_map_40, data_out_map_41, data_out_map_42, data_out_map_43, data_out_map_44, data_out_map_45, data_out_map_46, data_out_map_47, data_out_map_48, data_out_map_49, data_out_map_50, data_out_map_51, data_out_map_52, data_out_map_53, data_out_map_54, data_out_map_55, data_out_map_56, data_out_map_57, data_out_map_58, data_out_map_59, data_out_map_60, data_out_map_61, data_out_map_62, data_out_map_63, data_out_map_64, data_out_map_65, data_out_map_66, data_out_map_67, data_out_map_68, data_out_map_69, data_out_map_70, data_out_map_71, data_out_map_72, data_out_map_73, data_out_map_74, data_out_map_75, data_out_map_76, data_out_map_77, data_out_map_78, data_out_map_79, data_out_map_80, data_out_map_81, data_out_map_82, data_out_map_83, data_out_map_84, data_out_map_85, data_out_map_86, data_out_map_87, data_out_map_88, data_out_map_89, data_out_map_90, data_out_map_91, data_out_map_92, data_out_map_93, data_out_map_94, data_out_map_95, data_out_map_96, data_out_map_97, data_out_map_98, data_out_map_99, data_out_map_100, data_out_map_101, data_out_map_102, data_out_map_103, data_out_map_104, data_out_map_105, data_out_map_106, data_out_map_107, data_out_map_108, data_out_map_109, data_out_map_110, data_out_map_111, data_out_map_112, data_out_map_113, data_out_map_114, data_out_map_115, data_out_map_116, data_out_map_117, data_out_map_118, data_out_map_119, data_out_map_120, data_out_map_121, data_out_map_122, data_out_map_123, data_out_map_124, data_out_map_125, data_out_map_126, data_out_map_127 }),
  .dout({ S2[0], S2[1], S2[2], S2[3], S2[4], S2[5], S2[6], S2[7], S2[8], S2[9], S2[10], S2[11], S2[12], S2[13], S2[14], S2[15], S2[16], S2[17], S2[18], S2[19], S2[20], S2[21], S2[22], S2[23], S2[24], S2[25], S2[26], S2[27], S2[28], S2[29], S2[30], S2[31] }),
  .reg_out({ S4 }),
  .rst({ S5 }),
  .run({ hb0_map_ns_for:1_map_ns:4 })
);
mapn_1_6_1_1_1_1_1_12 #() 
mapn_1_6_1_1_1_1_1_12_1_ (
  .clk({ S0 }),
  .din({ S1[0], S1[1], S1[2], S1[3], S1[4], S1[5], S1[6], S1[7], S1[8], S1[9], S1[10], S1[11], S1[12], S1[13], S1[14], S1[15], S1[16], S1[17], S1[18], S1[19], S1[20], S1[21], S1[22], S1[23], S1[24], S1[25], S1[26], S1[27], S1[28], S1[29], S1[30], S1[31], S1[32], S1[33], S1[34], S1[35], S1[36], S1[37], S1[38], S1[39], S1[40], S1[41], S1[42], S1[43], S1[44], S1[45], S1[46], S1[47], S1[48], S1[49], S1[50], S1[51], S1[52], S1[53], S1[54], S1[55], S1[56], S1[57], S1[58], S1[59], S1[60], S1[61], S1[62], S1[63], S1[64], S1[65], S1[66], S1[67], S1[68], S1[69], S1[70], S1[71], S1[72], S1[73], S1[74], S1[75], S1[76], S1[77], S1[78], S1[79], S1[80], S1[81], S1[82], S1[83], S1[84], S1[85], S1[86], S1[87], S1[88], S1[89], S1[90], S1[91], S1[92], S1[93], S1[94], S1[95] }),
  .dout({ data_out_map_0, data_out_map_1, data_out_map_2, data_out_map_3, data_out_map_4, data_out_map_5, data_out_map_6, data_out_map_7, data_out_map_8, data_out_map_9, data_out_map_10, data_out_map_11, data_out_map_12, data_out_map_13, data_out_map_14, data_out_map_15, data_out_map_16, data_out_map_17, data_out_map_18, data_out_map_19, data_out_map_20, data_out_map_21, data_out_map_22, data_out_map_23, data_out_map_24, data_out_map_25, data_out_map_26, data_out_map_27, data_out_map_28, data_out_map_29, data_out_map_30, data_out_map_31 }),
  .pause({ S3 }),
  .reg_out({ hb0_map_ns_for:1_map_ns:4 }),
  .rst({ S5 }),
  .run({ S6 }),
  .w({ S7[0], S7[1], S7[2], S7[3], S7[4], S7[5], S7[6], S7[7], S7[8], S7[9], S7[10], S7[11], S7[12], S7[13], S7[14], S7[15], S7[16], S7[17], S7[18], S7[19], S7[20], S7[21], S7[22], S7[23], S7[24], S7[25], S7[26], S7[27], S7[28], S7[29], S7[30], S7[31], S7[32], S7[33], S7[34], S7[35], S7[36], S7[37], S7[38], S7[39], S7[40], S7[41], S7[42], S7[43], S7[44], S7[45], S7[46], S7[47], S7[48], S7[49], S7[50], S7[51], S7[52], S7[53], S7[54], S7[55], S7[56], S7[57], S7[58], S7[59], S7[60], S7[61], S7[62], S7[63], S7[64], S7[65], S7[66], S7[67], S7[68], S7[69], S7[70], S7[71], S7[72], S7[73], S7[74], S7[75], S7[76], S7[77], S7[78], S7[79], S7[80], S7[81], S7[82], S7[83], S7[84], S7[85], S7[86], S7[87], S7[88], S7[89], S7[90], S7[91], S7[92], S7[93], S7[94], S7[95] })
);
mapn_1_6_1_1_1_1_1_12 #() 
mapn_1_6_1_1_1_1_1_12_2_ (
  .clk({ S0 }),
  .din({ S1[96], S1[97], S1[98], S1[99], S1[100], S1[101], S1[102], S1[103], S1[104], S1[105], S1[106], S1[107], S1[108], S1[109], S1[110], S1[111], S1[112], S1[113], S1[114], S1[115], S1[116], S1[117], S1[118], S1[119], S1[120], S1[121], S1[122], S1[123], S1[124], S1[125], S1[126], S1[127], S1[128], S1[129], S1[130], S1[131], S1[132], S1[133], S1[134], S1[135], S1[136], S1[137], S1[138], S1[139], S1[140], S1[141], S1[142], S1[143], S1[144], S1[145], S1[146], S1[147], S1[148], S1[149], S1[150], S1[151], S1[152], S1[153], S1[154], S1[155], S1[156], S1[157], S1[158], S1[159], S1[160], S1[161], S1[162], S1[163], S1[164], S1[165], S1[166], S1[167], S1[168], S1[169], S1[170], S1[171], S1[172], S1[173], S1[174], S1[175], S1[176], S1[177], S1[178], S1[179], S1[180], S1[181], S1[182], S1[183], S1[184], S1[185], S1[186], S1[187], S1[188], S1[189], S1[190], S1[191] }),
  .dout({ data_out_map_32, data_out_map_33, data_out_map_34, data_out_map_35, data_out_map_36, data_out_map_37, data_out_map_38, data_out_map_39, data_out_map_40, data_out_map_41, data_out_map_42, data_out_map_43, data_out_map_44, data_out_map_45, data_out_map_46, data_out_map_47, data_out_map_48, data_out_map_49, data_out_map_50, data_out_map_51, data_out_map_52, data_out_map_53, data_out_map_54, data_out_map_55, data_out_map_56, data_out_map_57, data_out_map_58, data_out_map_59, data_out_map_60, data_out_map_61, data_out_map_62, data_out_map_63 }),
  .pause({ S3 }),
  .reg_out({ hb0_map_ns_for:2_map_ns:13 }),
  .rst({ S5 }),
  .run({ S6 }),
  .w({ S7[96], S7[97], S7[98], S7[99], S7[100], S7[101], S7[102], S7[103], S7[104], S7[105], S7[106], S7[107], S7[108], S7[109], S7[110], S7[111], S7[112], S7[113], S7[114], S7[115], S7[116], S7[117], S7[118], S7[119], S7[120], S7[121], S7[122], S7[123], S7[124], S7[125], S7[126], S7[127], S7[128], S7[129], S7[130], S7[131], S7[132], S7[133], S7[134], S7[135], S7[136], S7[137], S7[138], S7[139], S7[140], S7[141], S7[142], S7[143], S7[144], S7[145], S7[146], S7[147], S7[148], S7[149], S7[150], S7[151], S7[152], S7[153], S7[154], S7[155], S7[156], S7[157], S7[158], S7[159], S7[160], S7[161], S7[162], S7[163], S7[164], S7[165], S7[166], S7[167], S7[168], S7[169], S7[170], S7[171], S7[172], S7[173], S7[174], S7[175], S7[176], S7[177], S7[178], S7[179], S7[180], S7[181], S7[182], S7[183], S7[184], S7[185], S7[186], S7[187], S7[188], S7[189], S7[190], S7[191] })
);
mapn_1_6_1_1_1_1_1_12 #() 
mapn_1_6_1_1_1_1_1_12_3_ (
  .clk({ S0 }),
  .din({ S1[192], S1[193], S1[194], S1[195], S1[196], S1[197], S1[198], S1[199], S1[200], S1[201], S1[202], S1[203], S1[204], S1[205], S1[206], S1[207], S1[208], S1[209], S1[210], S1[211], S1[212], S1[213], S1[214], S1[215], S1[216], S1[217], S1[218], S1[219], S1[220], S1[221], S1[222], S1[223], S1[224], S1[225], S1[226], S1[227], S1[228], S1[229], S1[230], S1[231], S1[232], S1[233], S1[234], S1[235], S1[236], S1[237], S1[238], S1[239], S1[240], S1[241], S1[242], S1[243], S1[244], S1[245], S1[246], S1[247], S1[248], S1[249], S1[250], S1[251], S1[252], S1[253], S1[254], S1[255], S1[256], S1[257], S1[258], S1[259], S1[260], S1[261], S1[262], S1[263], S1[264], S1[265], S1[266], S1[267], S1[268], S1[269], S1[270], S1[271], S1[272], S1[273], S1[274], S1[275], S1[276], S1[277], S1[278], S1[279], S1[280], S1[281], S1[282], S1[283], S1[284], S1[285], S1[286], S1[287] }),
  .dout({ data_out_map_64, data_out_map_65, data_out_map_66, data_out_map_67, data_out_map_68, data_out_map_69, data_out_map_70, data_out_map_71, data_out_map_72, data_out_map_73, data_out_map_74, data_out_map_75, data_out_map_76, data_out_map_77, data_out_map_78, data_out_map_79, data_out_map_80, data_out_map_81, data_out_map_82, data_out_map_83, data_out_map_84, data_out_map_85, data_out_map_86, data_out_map_87, data_out_map_88, data_out_map_89, data_out_map_90, data_out_map_91, data_out_map_92, data_out_map_93, data_out_map_94, data_out_map_95 }),
  .pause({ S3 }),
  .reg_out({ hb0_map_ns_for:3_map_ns:22 }),
  .rst({ S5 }),
  .run({ S6 }),
  .w({ S7[192], S7[193], S7[194], S7[195], S7[196], S7[197], S7[198], S7[199], S7[200], S7[201], S7[202], S7[203], S7[204], S7[205], S7[206], S7[207], S7[208], S7[209], S7[210], S7[211], S7[212], S7[213], S7[214], S7[215], S7[216], S7[217], S7[218], S7[219], S7[220], S7[221], S7[222], S7[223], S7[224], S7[225], S7[226], S7[227], S7[228], S7[229], S7[230], S7[231], S7[232], S7[233], S7[234], S7[235], S7[236], S7[237], S7[238], S7[239], S7[240], S7[241], S7[242], S7[243], S7[244], S7[245], S7[246], S7[247], S7[248], S7[249], S7[250], S7[251], S7[252], S7[253], S7[254], S7[255], S7[256], S7[257], S7[258], S7[259], S7[260], S7[261], S7[262], S7[263], S7[264], S7[265], S7[266], S7[267], S7[268], S7[269], S7[270], S7[271], S7[272], S7[273], S7[274], S7[275], S7[276], S7[277], S7[278], S7[279], S7[280], S7[281], S7[282], S7[283], S7[284], S7[285], S7[286], S7[287] })
);
mapn_1_6_1_1_1_1_1_12 #() 
mapn_1_6_1_1_1_1_1_12_4_ (
  .clk({ S0 }),
  .din({ S1[288], S1[289], S1[290], S1[291], S1[292], S1[293], S1[294], S1[295], S1[296], S1[297], S1[298], S1[299], S1[300], S1[301], S1[302], S1[303], S1[304], S1[305], S1[306], S1[307], S1[308], S1[309], S1[310], S1[311], S1[312], S1[313], S1[314], S1[315], S1[316], S1[317], S1[318], S1[319], S1[320], S1[321], S1[322], S1[323], S1[324], S1[325], S1[326], S1[327], S1[328], S1[329], S1[330], S1[331], S1[332], S1[333], S1[334], S1[335], S1[336], S1[337], S1[338], S1[339], S1[340], S1[341], S1[342], S1[343], S1[344], S1[345], S1[346], S1[347], S1[348], S1[349], S1[350], S1[351], S1[352], S1[353], S1[354], S1[355], S1[356], S1[357], S1[358], S1[359], S1[360], S1[361], S1[362], S1[363], S1[364], S1[365], S1[366], S1[367], S1[368], S1[369], S1[370], S1[371], S1[372], S1[373], S1[374], S1[375], S1[376], S1[377], S1[378], S1[379], S1[380], S1[381], S1[382], S1[383] }),
  .dout({ data_out_map_96, data_out_map_97, data_out_map_98, data_out_map_99, data_out_map_100, data_out_map_101, data_out_map_102, data_out_map_103, data_out_map_104, data_out_map_105, data_out_map_106, data_out_map_107, data_out_map_108, data_out_map_109, data_out_map_110, data_out_map_111, data_out_map_112, data_out_map_113, data_out_map_114, data_out_map_115, data_out_map_116, data_out_map_117, data_out_map_118, data_out_map_119, data_out_map_120, data_out_map_121, data_out_map_122, data_out_map_123, data_out_map_124, data_out_map_125, data_out_map_126, data_out_map_127 }),
  .pause({ S3 }),
  .reg_out({ hb0_map_ns_for:4_map_ns:31 }),
  .rst({ S5 }),
  .run({ S6 }),
  .w({ S7[288], S7[289], S7[290], S7[291], S7[292], S7[293], S7[294], S7[295], S7[296], S7[297], S7[298], S7[299], S7[300], S7[301], S7[302], S7[303], S7[304], S7[305], S7[306], S7[307], S7[308], S7[309], S7[310], S7[311], S7[312], S7[313], S7[314], S7[315], S7[316], S7[317], S7[318], S7[319], S7[320], S7[321], S7[322], S7[323], S7[324], S7[325], S7[326], S7[327], S7[328], S7[329], S7[330], S7[331], S7[332], S7[333], S7[334], S7[335], S7[336], S7[337], S7[338], S7[339], S7[340], S7[341], S7[342], S7[343], S7[344], S7[345], S7[346], S7[347], S7[348], S7[349], S7[350], S7[351], S7[352], S7[353], S7[354], S7[355], S7[356], S7[357], S7[358], S7[359], S7[360], S7[361], S7[362], S7[363], S7[364], S7[365], S7[366], S7[367], S7[368], S7[369], S7[370], S7[371], S7[372], S7[373], S7[374], S7[375], S7[376], S7[377], S7[378], S7[379], S7[380], S7[381], S7[382], S7[383] })
);

endmodule