module PUNEH_Top_Module(clk, rst, writeMEM, readMEM, dataBus, addrBus);

wire S0;
wire S1;
wire S2;
wire S3;
wire S4;
wire S5;
wire S6;
wire S7;
wire S8;
wire S9;
wire S10;
wire S11;
wire S12;
wire S13;
wire S14;
wire S15;
wire S16;
wire S17;
wire S18;
wire S19;
wire S20;
wire S21;
wire S22;
wire S23;
wire S24;
wire S25;
wire S26;
wire S27;
wire S28;
wire S29;
wire S30;
wire S31;
wire S32;
wire S33;
wire S34;
wire S35;
wire S36;
wire S37;
wire S38;
wire S39;
wire S40;
wire S41;
wire S42;
wire S43;
wire S44;
wire S45;
wire S46;
wire S47;
wire S48;
wire S49;
wire S50;
wire S51;
wire S52;
wire S53;
wire S54;
wire S55;
wire S56;
wire S57;
wire S58;
wire S59;
wire S60;
wire S61;
wire S62;
wire S63;
wire S64;
wire S65;
wire S66;
wire S67;
wire S68;
wire S69;
wire S70;
wire S71;
wire S72;
wire S73;
wire S74;
wire S75;
wire S76;
wire S77;
wire S78;
wire S79;
wire S80;
wire S81;
wire S82;
wire S83;
wire S84;
wire S85;
wire S86;
wire S87;
wire S88;
wire S89;
wire S90;
wire S91;
wire S92;
wire S93;
wire S94;
wire S95;
wire S96;
wire S97;
wire S98;
wire S99;
wire S100;
wire S101;
wire S102;
wire S103;
wire S104;
wire S105;
wire S106;
wire S107;
wire S108;
wire S109;
wire S110;
wire S111;
wire S112;
wire S113;
wire S114;
wire S115;
wire S116;
wire S117;
wire S118;
wire S119;
wire S120;
wire S121;
wire S122;
wire S123;
wire S124;
wire S125;
wire S126;
wire S127;
wire S128;
wire S129;
wire S130;
wire S131;
wire S132;
wire S133;
wire S134;
wire S135;
wire S136;
wire S137;
wire S138;
wire S139;
wire S140;
wire S141;
wire S142;
wire S143;
wire S144;
wire S145;
wire S146;
wire S147;
wire S148;
wire S149;
wire S150;
wire S151;
wire S152;
wire S153;
wire S154;
wire S155;
wire S156;
wire S157;
wire S158;
wire S159;
wire S160;
wire S161;
wire S162;
wire S163;
wire S164;
wire S165;
wire S166;
wire S167;
wire S168;
wire S169;
wire S170;
wire S171;
wire S172;
wire S173;
wire S174;
wire S175;
wire S176;
wire S177;
wire S178;
wire S179;
wire S180;
wire S181;
wire S182;
wire S183;
wire S184;
wire S185;
wire S186;
wire S187;
wire S188;
wire S189;
wire S190;
wire S191;
wire S192;
wire S193;
wire S194;
wire S195;
wire S196;
wire S197;
wire S198;
wire S199;
wire S200;
wire S201;
wire S202;
wire S203;
wire S204;
wire S205;
wire S206;
wire S207;
wire S208;
wire S209;
wire S210;
wire S211;
wire S212;
wire S213;
wire S214;
wire S215;
wire S216;
wire S217;
wire S218;
wire S219;
wire S220;
wire S221;
wire S222;
wire S223;
wire S224;
wire S225;
wire S226;
wire S227;
wire S228;
wire S229;
wire S230;
wire S231;
wire S232;
wire S233;
wire S234;
wire S235;
wire S236;
wire S237;
wire S238;
wire S239;
wire S240;
wire S241;
wire S242;
wire S243;
wire S244;
wire S245;
wire S246;
wire S247;
wire S248;
wire S249;
wire S250;
wire S251;
wire S252;
wire S253;
wire S254;
wire S255;
wire S256;
wire S257;
wire S258;
wire S259;
wire S260;
wire S261;
wire S262;
wire S263;
wire S264;
wire S265;
wire S266;
wire S267;
wire S268;
wire S269;
wire S270;
wire S271;
wire S272;
wire S273;
wire S274;
wire S275;
wire S276;
wire S277;
wire S278;
wire S279;
wire S280;
wire S281;
wire S282;
wire S283;
wire S284;
wire S285;
wire S286;
wire S287;
wire S288;
wire S289;
wire S290;
wire S291;
wire S292;
wire S293;
wire S294;
wire S295;
wire S296;
wire S297;
wire S298;
wire S299;
wire S300;
wire S301;
wire S302;
wire S303;
wire S304;
wire S305;
wire S306;
wire S307;
wire S308;
wire S309;
wire S310;
wire S311;
wire S312;
wire S313;
wire S314;
wire S315;
wire S316;
wire S317;
wire S318;
wire S319;
wire S320;
wire S321;
wire S322;
wire S323;
wire S324;
wire S325;
wire S326;
wire S327;
wire S328;
wire S329;
wire S330;
wire S331;
wire S332;
wire S333;
wire S334;
wire S335;
wire S336;
wire S337;
wire S338;
wire S339;
wire S340;
wire S341;
wire S342;
wire S343;
wire S344;
wire S345;
wire S346;
wire S347;
wire S348;
wire S349;
wire S350;
wire S351;
wire S352;
wire S353;
wire S354;
wire S355;
wire S356;
wire S357;
wire S358;
wire S359;
wire S360;
wire S361;
wire S362;
wire S363;
wire S364;
wire S365;
wire S366;
wire S367;
wire S368;
wire S369;
wire S370;
wire S371;
wire S372;
wire S373;
wire S374;
wire S375;
wire S376;
wire S377;
wire S378;
wire S379;
wire S380;
wire S381;
wire S382;
wire S383;
wire S384;
wire S385;
wire S386;
wire S387;
wire S388;
wire S389;
wire S390;
wire S391;
wire S392;
wire S393;
wire S394;
wire S395;
wire S396;
wire S397;
wire S398;
wire S399;
wire S400;
wire S401;
wire S402;
wire S403;
wire S404;
wire S405;
wire S406;
wire S407;
wire S408;
wire S409;
wire S410;
wire S411;
wire S412;
wire S413;
wire S414;
wire S415;
wire S416;
wire S417;
wire S418;
wire S419;
wire S420;
wire S421;
wire S422;
wire S423;
wire S424;
wire S425;
wire S426;
wire S427;
wire S428;
wire S429;
wire S430;
wire S431;
wire S432;
wire S433;
wire S434;
wire S435;
wire S436;
wire S437;
wire S438;
wire S439;
wire S440;
wire S441;
wire S442;
wire S443;
wire S444;
wire S445;
wire S446;
wire S447;
wire S448;
wire S449;
wire S450;
wire S451;
wire S452;
wire S453;
wire S454;
wire S455;
wire S456;
wire S457;
wire S458;
wire S459;
wire S460;
wire S461;
wire S462;
wire S463;
wire S464;
wire S465;
wire S466;
wire S467;
wire S468;
wire S469;
wire S470;
wire S471;
wire S472;
wire S473;
wire S474;
wire S475;
wire S476;
wire S477;
wire S478;
wire S479;
wire S480;
wire S481;
wire S482;
wire S483;
wire S484;
wire S485;
wire S486;
wire S487;
wire S488;
wire S489;
wire S490;
wire S491;
wire S492;
wire S493;
wire S494;
wire S495;
wire S496;
wire S497;
wire S498;
wire S499;
wire S500;
wire S501;
wire S502;
wire S503;
wire S504;
wire S505;
wire S506;
wire S507;
wire S508;
wire S509;
wire S510;
wire S511;
wire S512;
wire S513;
wire S514;
wire S515;
wire S516;
wire S517;
wire S518;
wire S519;
wire S520;
wire S521;
wire S522;
wire S523;
wire S524;
wire S525;
wire S526;
wire S527;
wire S528;
wire S529;
wire S530;
wire S531;
wire S532;
wire S533;
wire S534;
wire S535;
wire S536;
wire S537;
wire S538;
wire S539;
wire S540;
wire S541;
wire S542;
wire S543;
wire S544;
wire S545;
wire S546;
wire S547;
wire S548;
wire S549;
wire S550;
wire S551;
wire S552;
wire S553;
wire S554;
wire S555;
wire S556;
wire S557;
wire S558;
wire S559;
wire S560;
wire S561;
wire S562;
wire S563;
wire S564;
wire S565;
wire S566;
wire S567;
wire S568;
wire S569;
wire S570;
wire S571;
wire S572;
wire S573;
wire S574;
wire S575;
wire S576;
wire S577;
wire S578;
wire S579;
wire S580;
wire S581;
wire S582;
wire S583;
wire S584;
wire S585;
wire S586;
wire S587;
wire S588;
wire S589;
wire S590;
wire S591;
wire S592;
wire S593;
wire S594;
wire S595;
wire S596;
wire S597;
wire S598;
wire S599;
wire S600;
wire S601;
wire S602;
wire S603;
wire S604;
wire S605;
wire S606;
wire S607;
wire S608;
wire S609;
wire S610;
wire S611;
wire S612;
wire S613;
wire S614;
wire S615;
wire S616;
wire S617;
wire S618;
wire S619;
wire S620;
wire S621;
wire S622;
wire S623;
wire S624;
wire S625;
wire S626;
wire S627;
wire S628;
wire S629;
wire S630;
wire S631;
wire S632;
wire S633;
wire S634;
wire S635;
wire S636;
wire S637;
wire S638;
wire S639;
wire S640;
wire S641;
wire S642;
wire S643;
wire S644;
wire S645;
wire S646;
wire S647;
wire S648;
wire S649;
wire S650;
wire S651;
wire S652;
wire S653;
wire S654;
wire S655;
wire S656;
wire S657;
wire S658;
wire S659;
wire S660;
wire S661;
wire S662;
wire S663;
wire S664;
wire S665;
wire S666;
wire S667;
wire S668;
wire S669;
wire S670;
wire S671;
wire S672;
wire S673;
wire S674;
wire S675;
wire S676;
wire S677;
wire S678;
wire S679;
wire S680;
wire S681;
wire S682;
wire S683;
wire S684;
wire S685;
wire S686;
wire S687;
wire S688;
wire S689;
wire S690;
wire S691;
wire S692;
wire S693;
wire S694;
wire S695;
wire S696;
wire S697;
wire S698;
wire S699;
wire S700;
wire S701;
wire S702;
wire S703;
wire S704;
wire S705;
wire S706;
wire S707;
wire S708;
wire S709;
wire S710;
wire S711;
wire S712;
wire S713;
wire S714;
wire S715;
wire S716;
wire S717;
wire S718;
wire S719;
wire S720;
wire S721;
wire S722;
wire S723;
wire S724;
wire S725;
wire S726;
wire S727;
wire S728;
wire S729;
wire S730;
wire S731;
wire S732;
wire S733;
wire S734;
wire S735;
wire S736;
wire S737;
wire S738;
wire S739;
wire S740;
wire S741;
wire S742;
wire S743;
wire S744;
wire S745;
wire S746;
wire S747;
wire S748;
wire S749;
wire S750;
wire S751;
wire S752;
wire S753;
wire S754;
wire S755;
wire S756;
wire S757;
wire S758;
wire S759;
wire S760;
wire S761;
wire S762;
wire S763;
wire S764;
wire S765;
wire S766;
wire S767;
wire S768;
wire S769;
wire S770;
wire S771;
wire S772;
wire S773;
wire S774;
wire S775;
wire S776;
wire S777;
wire S778;
wire S779;
wire S780;
wire S781;
wire S782;
wire S783;
wire S784;
wire S785;
wire S786;
wire S787;
wire S788;
wire S789;
wire S790;
wire S791;
wire S792;
wire S793;
wire S794;
wire S795;
wire S796;
wire S797;
wire S798;
wire S799;
wire S800;
wire S801;
wire S802;
wire S803;
wire S804;
wire S805;
wire S806;
wire S807;
wire S808;
wire S809;
wire S810;
wire S811;
wire S812;
wire S813;
wire S814;
wire S815;
wire S816;
wire S817;
wire S818;
wire S819;
wire S820;
wire S821;
wire S822;
wire S823;
wire S824;
wire S825;
wire S826;
wire S827;
wire S828;
wire S829;
wire S830;
wire S831;
wire S832;
wire S833;
wire S834;
wire S835;
wire S836;
wire S837;
wire S838;
wire S839;
wire S840;
wire S841;
wire S842;
wire S843;
wire S844;
wire S845;
wire S846;
wire S847;
wire S848;
wire S849;
wire S850;
wire S851;
wire S852;
wire S853;
wire S854;
wire S855;
wire S856;
wire S857;
wire S858;
wire S859;
wire S860;
wire S861;
wire S862;
wire S863;
wire S864;
wire S865;
wire S866;
wire S867;
wire S868;
wire S869;
wire S870;
wire S871;
wire S872;
wire S873;
wire S874;
wire S875;
wire S876;
wire S877;
wire S878;
wire S879;
wire S880;
wire S881;
wire S882;
wire S883;
wire S884;
wire S885;
wire S886;
wire S887;
wire S888;
wire S889;
wire S890;
wire S891;
wire S892;
wire S893;
wire S894;
wire S895;
wire S896;
wire S897;
wire S898;
wire S899;
wire S900;
wire S901;
wire S902;
wire S903;
wire S904;
wire S905;
wire S906;
wire S907;
wire S908;
wire S909;
wire S910;
wire S911;
wire S912;
wire S913;
wire S914;
wire S915;
wire S916;
wire S917;
wire S918;
wire S919;
wire S920;
wire S921;
wire S922;
wire S923;
wire S924;
wire S925;
wire S926;
wire S927;
wire S928;
wire S929;
wire S930;
wire S931;
wire S932;
wire S933;
wire S934;
wire S935;
wire S936;
wire S937;
wire S938;
wire S939;
wire S940;
wire S941;
wire S942;
wire S943;
wire S944;
wire S945;
wire S946;
wire S947;
wire S948;
wire S949;
wire S950;
wire S951;
wire S952;
wire S953;
wire S954;
wire S955;
wire S956;
wire S957;
wire S958;
wire S959;
wire S960;
wire S961;
wire S962;
wire S963;
wire S964;
wire S965;
wire S966;
wire S967;
wire S968;
wire S969;
wire S970;
wire S971;
wire S972;
wire S973;
wire S974;
wire S975;
wire S976;
wire S977;
wire S978;
wire S979;
wire S980;
wire S981;
wire S982;
wire S983;
wire S984;
wire S985;
wire S986;
wire S987;
wire S988;
wire S989;
wire S990;
wire S991;
wire S992;
wire S993;
wire S994;
wire S995;
wire S996;
wire S997;
wire S998;
wire S999;
wire S1000;
wire S1001;
wire S1002;
wire S1003;
wire S1004;
wire S1005;
wire S1006;
wire S1007;
wire S1008;
wire S1009;
wire S1010;
wire S1011;
wire S1012;
wire S1013;
wire S1014;
wire S1015;
wire S1016;
wire S1017;
wire S1018;
wire S1019;
wire S1020;
wire S1021;
wire S1022;
wire S1023;
wire S1024;
wire S1025;
wire S1026;
wire S1027;
wire S1028;
wire S1029;
wire S1030;
wire S1031;
wire S1032;
wire S1033;
wire S1034;
wire S1035;
wire S1036;
wire S1037;
wire S1038;
wire S1039;
wire S1040;
wire S1041;
wire S1042;
wire S1043;
wire S1044;
wire S1045;
wire S1046;
wire S1047;
wire S1048;
wire S1049;
wire S1050;
wire S1051;
wire S1052;
wire S1053;
wire S1054;
wire S1055;
wire S1056;
wire S1057;
wire S1058;
wire S1059;
wire S1060;
wire S1061;
wire S1062;
wire S1063;
wire S1064;
wire S1065;
wire S1066;
wire S1067;
wire S1068;
wire S1069;
wire S1070;
wire S1071;
wire S1072;
wire S1073;
wire S1074;
wire S1075;
wire S1076;
wire S1077;
wire S1078;
wire S1079;
wire S1080;
wire S1081;
wire S1082;
wire S1083;
wire S1084;
wire S1085;
wire S1086;
wire S1087;
wire S1088;
wire S1089;
wire S1090;
wire S1091;
wire S1092;
wire S1093;
wire S1094;
wire S1095;
wire S1096;
wire S1097;
wire S1098;
wire S1099;
wire S1100;
wire S1101;
wire S1102;
wire S1103;
wire S1104;
wire S1105;
wire S1106;
wire S1107;
wire S1108;
wire S1109;
wire S1110;
wire S1111;
wire S1112;
wire S1113;
wire S1114;
wire S1115;
wire S1116;
wire S1117;
wire S1118;
wire S1119;
wire S1120;
wire S1121;
wire S1122;
wire S1123;
wire S1124;
wire S1125;
wire S1126;
wire S1127;
wire S1128;
wire S1129;
wire S1130;
wire S1131;
wire S1132;
wire S1133;
wire S1134;
wire S1135;
wire S1136;
wire S1137;
wire S1138;
wire S1139;
wire S1140;
wire S1141;
wire S1142;
wire S1143;
wire S1144;
wire S1145;
wire S1146;
wire S1147;
wire S1148;
wire S1149;
wire S1150;
wire S1151;
wire S1152;
wire S1153;
wire S1154;
wire S1155;
wire S1156;
wire S1157;
wire S1158;
wire S1159;
wire S1160;
wire S1161;
wire S1162;
wire S1163;
wire S1164;
wire S1165;
wire S1166;
wire S1167;
wire S1168;
wire S1169;
wire S1170;
wire S1171;
wire S1172;
wire S1173;
wire S1174;
wire S1175;
wire S1176;
wire S1177;
wire S1178;
wire S1179;
wire S1180;
wire S1181;
wire S1182;
wire S1183;
wire S1184;
wire S1185;
wire S1186;
wire S1187;
wire S1188;
wire S1189;
wire S1190;
wire S1191;
wire S1192;
wire S1193;
wire S1194;
wire S1195;
wire S1196;
wire S1197;
wire S1198;
wire S1199;
wire S1200;
wire S1201;
wire S1202;
wire S1203;
wire S1204;
wire S1205;
wire S1206;
wire S1207;
wire S1208;
wire S1209;
wire S1210;
wire S1211;
wire S1212;
wire S1213;
wire S1214;
wire S1215;
wire S1216;
wire S1217;
wire S1218;
wire S1219;
wire S1220;
wire S1221;
wire S1222;
wire S1223;
wire S1224;
wire S1225;
wire S1226;
wire S1227;
wire S1228;
wire S1229;
wire S1230;
wire S1231;
wire S1232;
wire S1233;
wire S1234;
wire S1235;
wire S1236;
wire S1237;
wire S1238;
wire S1239;
wire S1240;
wire S1241;
wire S1242;
wire S1243;
wire S1244;
wire S1245;
wire S1246;
wire S1247;
wire S1248;
wire S1249;
wire S1250;
wire S1251;
wire S1252;
wire S1253;
wire S1254;
wire S1255;
wire S1256;
wire S1257;
wire S1258;
wire S1259;
wire S1260;
wire S1261;
wire S1262;
wire S1263;
wire S1264;
wire S1265;
wire S1266;
wire S1267;
wire S1268;
wire S1269;
wire S1270;
wire S1271;
wire S1272;
wire S1273;
wire S1274;
wire S1275;
wire S1276;
wire S1277;
wire S1278;
wire S1279;
wire S1280;
wire S1281;
wire S1282;
wire S1283;
wire S1284;
wire S1285;
wire S1286;
wire S1287;
wire S1288;
wire S1289;
wire S1290;
wire S1291;
wire S1292;
wire S1293;
wire S1294;
wire S1295;
wire S1296;
wire S1297;
wire S1298;
wire S1299;
wire S1300;
wire S1301;
wire S1302;
wire S1303;
wire S1304;
wire S1305;
wire S1306;
wire S1307;
wire S1308;
wire S1309;
wire S1310;
wire S1311;
wire S1312;
wire S1313;
wire S1314;
wire S1315;
wire S1316;
wire S1317;
wire S1318;
wire S1319;
wire S1320;
wire S1321;
wire S1322;
wire S1323;
wire S1324;
wire S1325;
wire S1326;
wire S1327;
wire S1328;
wire S1329;
wire S1330;
wire S1331;
wire S1332;
wire S1333;
wire S1334;
wire S1335;
wire S1336;
wire S1337;
wire S1338;
wire S1339;
wire S1340;
wire S1341;
wire S1342;
wire S1343;
wire S1344;
wire S1345;
wire S1346;
wire S1347;
wire S1348;
wire S1349;
wire S1350;
wire S1351;
wire S1352;
wire S1353;
wire S1354;
wire S1355;
wire S1356;
wire S1357;
wire S1358;
wire S1359;
wire S1360;
wire S1361;
wire S1362;
wire S1363;
wire S1364;
wire S1365;
wire S1366;
wire S1367;
wire S1368;
wire S1369;
wire S1370;
wire S1371;
wire S1372;
wire S1373;
wire S1374;
wire S1375;
wire S1376;
wire S1377;
wire S1378;
wire S1379;
wire S1380;
wire S1381;
wire S1382;
wire S1383;
wire S1384;
wire S1385;
wire S1386;
wire S1387;
wire S1388;
wire S1389;
wire S1390;
wire S1391;
wire S1392;
wire S1393;
wire S1394;
wire S1395;
wire S1396;
wire S1397;
wire S1398;
wire S1399;
wire S1400;
wire S1401;
wire S1402;
wire S1403;
wire S1404;
wire S1405;
wire S1406;
wire S1407;
wire S1408;
wire S1409;
wire S1410;
wire S1411;
wire S1412;
wire S1413;
wire S1414;
wire S1415;
wire S1416;
wire S1417;
wire S1418;
wire S1419;
wire S1420;
wire S1421;
wire S1422;
wire S1423;
wire S1424;
wire S1425;
wire S1426;
wire S1427;
wire S1428;
wire S1429;
wire S1430;
wire S1431;
wire S1432;
wire S1433;
wire S1434;
wire S1435;
wire S1436;
wire S1437;
wire S1438;
wire S1439;
wire S1440;
wire S1441;
wire S1442;
wire S1443;
wire S1444;
wire S1445;
wire S1446;
wire S1447;
wire S1448;
wire S1449;
wire S1450;
wire S1451;
wire S1452;
wire S1453;
wire S1454;
wire S1455;
wire S1456;
wire S1457;
wire S1458;
wire S1459;
wire S1460;
wire S1461;
wire S1462;
wire S1463;
wire S1464;
wire S1465;
wire S1466;
wire S1467;
wire S1468;
wire S1469;
wire S1470;
wire S1471;
wire S1472;
wire S1473;
wire S1474;
wire S1475;
wire S1476;
wire S1477;
wire S1478;
wire S1479;
wire S1480;
wire S1481;
wire S1482;
wire S1483;
wire S1484;
wire S1485;
wire S1486;
wire S1487;
wire S1488;
wire S1489;
wire S1490;
wire S1491;
wire S1492;
wire S1493;
wire S1494;
wire S1495;
wire S1496;
wire S1497;
wire S1498;
wire S1499;
wire S1500;
wire S1501;
wire S1502;
wire S1503;
wire S1504;
wire S1505;
wire S1506;
wire S1507;
wire S1508;
wire S1509;
wire S1510;
wire S1511;
wire S1512;
wire S1513;
wire S1514;
wire S1515;
wire S1516;
wire S1517;
wire S1518;
wire S1519;
wire S1520;
wire S1521;
wire S1522;
wire S1523;
wire S1524;
wire S1525;
wire S1526;
wire S1527;
wire S1528;
wire S1529;
wire S1530;
wire S1531;
wire S1532;
wire S1533;
wire S1534;
wire S1535;
wire S1536;
wire S1537;
wire S1538;
wire S1539;
wire S1540;
wire S1541;
wire S1542;
wire S1543;
wire S1544;
wire S1545;
wire S1546;
wire S1547;
wire S1548;
wire S1549;
wire S1550;
wire S1551;
wire S1552;
wire S1553;
wire S1554;
wire S1555;
wire S1556;
wire S1557;
wire S1558;
wire S1559;
wire S1560;
wire S1561;
wire S1562;
wire S1563;
wire S1564;
wire S1565;
wire S1566;
wire S1567;
wire S1568;
wire S1569;
wire S1570;
wire S1571;
wire S1572;
wire S1573;
wire S1574;
wire S1575;
wire S1576;
wire S1577;
wire S1578;
wire S1579;
wire S1580;
wire S1581;
wire S1582;
wire S1583;
wire S1584;
wire S1585;
wire S1586;
wire S1587;
wire S1588;
wire S1589;
wire S1590;
wire S1591;
wire S1592;
wire S1593;
wire S1594;
wire S1595;
wire S1596;
wire S1597;
wire S1598;
wire S1599;
wire S1600;
wire S1601;
wire S1602;
wire S1603;
wire S1604;
wire S1605;
wire S1606;
wire S1607;
wire S1608;
wire S1609;
wire S1610;
wire S1611;
wire S1612;
wire S1613;
wire S1614;
wire S1615;
wire S1616;
wire S1617;
wire S1618;
wire S1619;
wire S1620;
wire S1621;
wire S1622;
wire S1623;
wire S1624;
wire S1625;
wire S1626;
wire S1627;
wire S1628;
wire S1629;
wire S1630;
wire S1631;
wire S1632;
wire S1633;
wire S1634;
wire S1635;
wire S1636;
wire S1637;
wire S1638;
wire S1639;
wire S1640;
wire S1641;
wire S1642;
wire S1643;
wire S1644;
wire S1645;
wire S1646;
wire S1647;
wire S1648;
wire S1649;
wire S1650;
wire S1651;
wire S1652;
wire S1653;
wire S1654;
wire S1655;
wire S1656;
wire S1657;
wire S1658;
wire S1659;
wire S1660;
wire S1661;
wire S1662;
wire S1663;
wire S1664;
wire S1665;
wire S1666;
wire S1667;
wire S1668;
wire S1669;
wire S1670;
wire S1671;
wire S1672;
wire S1673;
wire S1674;
wire S1675;
wire S1676;
wire S1677;
wire S1678;
wire S1679;
wire S1680;
wire S1681;
wire S1682;
wire S1683;
wire S1684;
wire S1685;
wire S1686;
wire S1687;
wire S1688;
wire S1689;
wire S1690;
wire S1691;
wire S1692;
wire S1693;
wire S1694;
wire S1695;
wire S1696;
wire S1697;
wire S1698;
wire S1699;
wire S1700;
wire S1701;
wire S1702;
wire S1703;
wire S1704;
wire S1705;
wire S1706;
wire S1707;
wire S1708;
wire S1709;
wire S1710;
wire S1711;
wire S1712;
wire S1713;
wire S1714;
wire S1715;
wire S1716;
wire S1717;
wire S1718;
wire S1719;
wire S1720;
wire S1721;
wire S1722;
wire S1723;
wire S1724;
wire S1725;
wire S1726;
wire S1727;
wire S1728;
wire S1729;
wire S1730;
wire S1731;
wire S1732;
wire S1733;
wire S1734;
wire S1735;
wire S1736;
wire S1737;
wire S1738;
wire S1739;
wire S1740;
wire S1741;
wire S1742;
wire S1743;
wire S1744;
wire S1745;
wire S1746;
wire S1747;
wire S1748;
wire S1749;
wire S1750;
wire S1751;
wire S1752;
wire S1753;
wire S1754;
wire S1755;
wire S1756;
wire S1757;
wire S1758;
wire S1759;
wire S1760;
wire S1761;
wire S1762;
wire S1763;
wire S1764;
wire S1765;
wire S1766;
wire S1767;
wire S1768;
wire S1769;
wire S1770;
wire S1771;
wire S1772;
wire S1773;
wire S1774;
wire S1775;
wire S1776;
wire S1777;
wire S1778;
wire S1779;
wire S1780;
wire S1781;
wire S1782;
wire S1783;
wire S1784;
wire S1785;
wire S1786;
wire S1787;
wire S1788;
wire S1789;
wire S1790;
wire S1791;
wire S1792;
wire S1793;
wire S1794;
wire S1795;
wire S1796;
wire S1797;
wire S1798;
wire S1799;
wire S1800;
wire S1801;
wire S1802;
wire S1803;
wire S1804;
wire S1805;
wire S1806;
wire S1807;
wire S1808;
wire S1809;
wire S1810;
wire S1811;
wire S1812;
wire S1813;
wire S1814;
wire S1815;
wire S1816;
wire S1817;
wire S1818;
wire S1819;
wire S1820;
wire S1821;
wire S1822;
wire S1823;
wire S1824;
wire S1825;
wire S1826;
wire S1827;
wire S1828;
wire S1829;
wire S1830;
wire S1831;
wire S1832;
wire S1833;
wire S1834;
wire S1835;
wire S1836;
wire S1837;
wire S1838;
wire S1839;
wire S1840;
wire S1841;
wire S1842;
wire S1843;
wire S1844;
wire S1845;
wire S1846;
wire S1847;
wire S1848;
wire S1849;
wire S1850;
wire S1851;
wire S1852;
wire S1853;
wire S1854;
wire S1855;
wire S1856;
wire S1857;
wire S1858;
wire S1859;
wire S1860;
wire S1861;
wire S1862;
wire S1863;
wire S1864;
wire S1865;
wire S1866;
wire S1867;
wire S1868;
wire S1869;
wire S1870;
wire S1871;
wire S1872;
wire S1873;
wire S1874;
wire S1875;
wire S1876;
wire S1877;
wire S1878;
wire S1879;
wire S1880;
wire S1881;
wire S1882;
wire S1883;
wire S1884;
wire S1885;
wire S1886;
wire S1887;
wire S1888;
wire S1889;
wire S1890;
wire S1891;
wire S1892;
wire S1893;
wire S1894;
wire S1895;
wire S1896;
wire S1897;
wire S1898;
wire S1899;
wire S1900;
wire S1901;
wire S1902;
wire S1903;
wire S1904;
wire S1905;
wire S1906;
wire S1907;
wire S1908;
wire S1909;
wire S1910;
wire S1911;
wire S1912;
wire S1913;
wire S1914;
wire S1915;
wire S1916;
wire S1917;
wire S1918;
wire S1919;
wire S1920;
wire S1921;
wire S1922;
wire S1923;
wire S1924;
wire S1925;
wire S1926;
wire S1927;
wire S1928;
wire S1929;
wire S1930;
wire S1931;
wire S1932;
wire S1933;
wire S1934;
wire S1935;
wire S1936;
wire S1937;
wire S1938;
wire S1939;
wire S1940;
wire S1941;
wire S1942;
wire S1943;
wire S1944;
wire S1945;
wire S1946;
wire S1947;
wire S1948;
wire S1949;
wire S1950;
wire S1951;
wire S1952;
wire S1953;
wire S1954;
wire S1955;
wire S1956;
wire S1957;
wire S1958;
wire S1959;
wire S1960;
wire S1961;
wire S1962;
wire S1963;
wire S1964;
wire S1965;
wire S1966;
wire S1967;
wire S1968;
wire S1969;
wire S1970;
wire S1971;
wire S1972;
wire S1973;
wire S1974;
wire S1975;
wire S1976;
wire S1977;
wire S1978;
wire S1979;
wire S1980;
wire S1981;
wire S1982;
wire S1983;
wire S1984;
wire S1985;
wire S1986;
wire S1987;
wire S1988;
wire S1989;
wire S1990;
wire S1991;
wire S1992;
wire S1993;
wire S1994;
wire S1995;
wire S1996;
wire S1997;
wire S1998;
wire S1999;
wire S2000;
wire S2001;
wire S2002;
wire S2003;
wire S2004;
wire S2005;
wire S2006;
wire S2007;
wire S2008;
wire S2009;
wire S2010;
wire S2011;
wire S2012;
wire S2013;
wire S2014;
wire S2015;
wire S2016;
wire S2017;
wire S2018;
wire S2019;
wire S2020;
wire S2021;
wire S2022;
wire S2023;
wire S2024;
wire S2025;
wire S2026;
wire S2027;
wire S2028;
wire S2029;
wire S2030;
wire S2031;
wire S2032;
wire S2033;
wire S2034;
wire S2035;
wire S2036;
wire S2037;
wire S2038;
wire S2039;
wire S2040;
wire S2041;
wire S2042;
wire S2043;
wire S2044;
wire S2045;
wire S2046;
wire S2047;
wire S2048;
wire S2049;
wire S2050;
wire S2051;
wire S2052;
wire S2053;
wire S2054;
wire S2055;
wire S2056;
wire S2057;
wire S2058;
wire S2059;
wire S2060;
wire S2061;
wire S2062;
wire S2063;
wire S2064;
wire S2065;
wire S2066;
wire S2067;
wire S2068;
wire S2069;
wire S2070;
wire S2071;
wire S2072;
wire S2073;
wire S2074;
wire S2075;
wire S2076;
wire S2077;
wire S2078;
wire S2079;
wire S2080;
wire S2081;
wire S2082;
wire S2083;
wire S2084;
wire S2085;
wire S2086;
wire S2087;
wire S2088;
wire S2089;
wire S2090;
wire S2091;
wire S2092;
wire S2093;
wire S2094;
wire S2095;
wire S2096;
wire S2097;
wire S2098;
wire S2099;
wire S2100;
wire S2101;
wire S2102;
wire S2103;
wire S2104;
wire S2105;
wire S2106;
wire S2107;
wire S2108;
wire S2109;
wire S2110;
wire S2111;
wire S2112;
wire S2113;
wire S2114;
wire S2115;
wire S2116;
wire S2117;
wire S2118;
wire S2119;
wire S2120;
wire S2121;
wire S2122;
wire S2123;
wire S2124;
wire S2125;
wire S2126;
wire S2127;
wire S2128;
wire S2129;
wire S2130;
wire S2131;
wire S2132;
wire S2133;
wire S2134;
wire S2135;
wire S2136;
wire S2137;
wire S2138;
wire S2139;
wire S2140;
wire S2141;
wire S2142;
wire S2143;
wire S2144;
wire S2145;
wire S2146;
wire S2147;
wire S2148;
wire S2149;
wire S2150;
wire S2151;
wire S2152;
wire S2153;
wire S2154;
wire S2155;
wire S2156;
wire S2157;
wire S2158;
wire S2159;
wire S2160;
wire S2161;
wire S2162;
wire S2163;
wire S2164;
wire S2165;
wire S2166;
wire S2167;
wire S2168;
wire S2169;
wire S2170;
wire S2171;
wire S2172;
wire S2173;
wire S2174;
wire S2175;
wire S2176;
wire S2177;
wire S2178;
wire S2179;
wire S2180;
wire S2181;
wire S2182;
wire S2183;
wire S2184;
wire S2185;
wire S2186;
wire S2187;
wire S2188;
wire S2189;
wire S2190;
wire S2191;
wire S2192;
wire S2193;
wire S2194;
wire S2195;
wire S2196;
wire S2197;
wire S2198;
wire S2199;
wire S2200;
wire S2201;
wire S2202;
wire S2203;
wire S2204;
wire S2205;
wire S2206;
wire S2207;
wire S2208;
wire S2209;
wire S2210;
wire S2211;
wire S2212;
wire S2213;
wire S2214;
wire S2215;
wire S2216;
wire S2217;
wire S2218;
wire S2219;
wire S2220;
wire S2221;
wire S2222;
wire S2223;
wire S2224;
wire S2225;
wire S2226;
wire S2227;
wire S2228;
wire S2229;
wire S2230;
wire S2231;
wire S2232;
wire S2233;
wire S2234;
wire S2235;
wire S2236;
wire S2237;
wire S2238;
wire S2239;
wire S2240;
wire S2241;
wire S2242;
wire S2243;
wire S2244;
wire S2245;
wire S2246;
wire S2247;
wire S2248;
wire S2249;
wire S2250;
wire S2251;
wire S2252;
wire S2253;
wire S2254;
wire S2255;
wire S2256;
wire S2257;
wire S2258;
wire S2259;
wire S2260;
wire S2261;
wire S2262;
wire S2263;
wire S2264;
wire S2265;
wire S2266;
wire S2267;
wire S2268;
wire S2269;
wire S2270;
wire S2271;
wire S2272;
wire S2273;
wire S2274;
wire S2275;
wire S2276;
wire S2277;
wire S2278;
wire S2279;
wire S2280;
wire S2281;
wire S2282;
wire S2283;
wire S2284;
wire S2285;
wire S2286;
wire S2287;
wire S2288;
wire S2289;
wire S2290;
wire S2291;
wire S2292;
wire S2293;
wire S2294;
wire S2295;
wire S2296;
wire S2297;
wire S2298;
wire S2299;
wire S2300;
wire S2301;
wire S2302;
wire S2303;
wire S2304;
wire S2305;
wire S2306;
wire S2307;
wire S2308;
wire S2309;
wire S2310;
wire S2311;
wire S2312;
wire S2313;
wire S2314;
wire S2315;
wire S2316;
wire S2317;
wire S2318;
wire S2319;
wire S2320;
wire S2321;
wire S2322;
wire S2323;
wire S2324;
wire S2325;
wire S2326;
wire S2327;
wire S2328;
wire S2329;
wire S2330;
wire S2331;
wire S2332;
wire S2333;
wire S2334;
wire S2335;
wire S2336;
wire S2337;
wire S2338;
wire S2339;
wire S2340;
wire S2341;
wire S2342;
wire S2343;
wire S2344;
wire S2345;
wire S2346;
wire S2347;
wire S2348;
wire S2349;
wire S2350;
wire S2351;
wire S2352;
wire S2353;
wire S2354;
wire S2355;
wire S2356;
wire S2357;
wire S2358;
wire S2359;
wire S2360;
wire S2361;
wire S2362;
wire S2363;
wire S2364;
wire S2365;
wire S2366;
wire S2367;
wire S2368;
wire S2369;
wire S2370;
wire S2371;
wire S2372;
wire S2373;
wire S2374;
wire S2375;
wire S2376;
wire S2377;
wire S2378;
wire S2379;
wire S2380;
wire S2381;
wire S2382;
wire S2383;
wire S2384;
wire S2385;
wire S2386;
wire S2387;
wire S2388;
wire S2389;
wire S2390;
wire S2391;
wire S2392;
wire S2393;
wire S2394;
wire S2395;
wire S2396;
wire S2397;
wire S2398;
wire S2399;
wire S2400;
wire S2401;
wire S2402;
wire S2403;
wire S2404;
wire S2405;
wire S2406;
wire S2407;
wire S2408;
wire S2409;
wire S2410;
wire S2411;
wire S2412;
wire S2413;
wire S2414;
wire S2415;
wire S2416;
wire S2417;
wire S2418;
wire S2419;
wire S2420;
wire S2421;
wire S2422;
wire S2423;
wire S2424;
wire S2425;
wire S2426;
wire S2427;
wire S2428;
wire S2429;
wire S2430;
wire S2431;
wire S2432;
wire S2433;
wire S2434;
wire S2435;
wire S2436;
wire S2437;
wire S2438;
wire S2439;
wire S2440;
wire S2441;
wire S2442;
wire S2443;
wire S2444;
wire S2445;
wire S2446;
wire S2447;
wire S2448;
wire S2449;
wire S2450;
wire S2451;
wire S2452;
wire S2453;
wire S2454;
wire S2455;
wire S2456;
wire S2457;
wire S2458;
wire S2459;
wire S2460;
wire S2461;
wire S2462;
wire S2463;
wire S2464;
wire S2465;
wire S2466;
wire S2467;
wire S2468;
wire S2469;
wire S2470;
wire S2471;
wire S2472;
wire S2473;
wire S2474;
wire S2475;
wire S2476;
wire S2477;
wire S2478;
wire S2479;
wire S2480;
wire S2481;
wire S2482;
wire S2483;
wire S2484;
wire S2485;
wire S2486;
wire S2487;
wire S2488;
wire S2489;
wire S2490;
wire S2491;
wire S2492;
wire S2493;
wire S2494;
wire S2495;
wire S2496;
wire S2497;
wire S2498;
wire S2499;
wire S2500;
wire S2501;
wire S2502;
wire S2503;
wire S2504;
wire S2505;
wire S2506;
wire S2507;
wire S2508;
wire S2509;
wire S2510;
wire S2511;
wire S2512;
wire S2513;
wire S2514;
wire S2515;
wire S2516;
wire S2517;
wire S2518;
wire S2519;
wire S2520;
wire S2521;
wire S2522;
wire S2523;
wire S2524;
wire S2525;
wire S2526;
wire S2527;
wire S2528;
wire S2529;
wire S2530;
wire S2531;
wire S2532;
wire S2533;
wire S2534;
wire S2535;
wire S2536;
wire S2537;
wire S2538;
wire S2539;
wire S2540;
wire S2541;
wire S2542;
wire S2543;
wire S2544;
wire S2545;
wire S2546;
wire S2547;
wire S2548;
wire S2549;
wire S2550;
wire S2551;
wire S2552;
wire S2553;
wire S2554;
wire S2555;
wire S2556;
wire S2557;
wire S2558;
wire S2559;
wire S2560;
wire S2561;
wire S2562;
wire S2563;
wire S2564;
wire S2565;
wire S2566;
wire S2567;
wire S2568;
wire S2569;
wire S2570;
wire S2571;
wire S2572;
wire S2573;
wire S2574;
wire S2575;
wire S2576;
wire S2577;
wire S2578;
wire S2579;
wire S2580;
wire S2581;
wire S2582;
wire S2583;
wire S2584;
wire S2585;
wire S2586;
wire S2587;
wire S2588;
wire S2589;
wire S2590;
wire S2591;
wire S2592;
wire S2593;
wire S2594;
wire S2595;
wire S2596;
wire S2597;
wire S2598;
wire S2599;
wire S2600;
wire S2601;
wire S2602;
wire S2603;
wire S2604;
wire S2605;
wire S2606;
wire S2607;
wire S2608;
wire S2609;
wire S2610;
wire S2611;
wire S2612;
wire S2613;
wire S2614;
wire S2615;
wire S2616;
wire S2617;
wire S2618;
wire S2619;
wire S2620;
wire S2621;
wire S2622;
wire S2623;
wire S2624;
wire S2625;
wire S2626;
wire S2627;
wire S2628;
wire S2629;
wire S2630;
wire S2631;
wire S2632;
wire S2633;
wire S2634;
wire S2635;
wire S2636;
wire S2637;
wire S2638;
wire S2639;
wire S2640;
wire S2641;
wire S2642;
wire S2643;
wire S2644;
wire S2645;
wire S2646;
wire S2647;
wire S2648;
wire S2649;
wire S2650;
wire S2651;
wire S2652;
wire S2653;
wire S2654;
wire S2655;
wire S2656;
wire S2657;
wire S2658;
wire S2659;
wire S2660;
wire S2661;
wire S2662;
wire S2663;
wire S2664;
wire S2665;
wire S2666;
wire S2667;
wire S2668;
wire S2669;
wire S2670;
wire S2671;
wire S2672;
wire S2673;
wire S2674;
wire S2675;
wire S2676;
wire S2677;
wire S2678;
wire S2679;
wire S2680;
wire S2681;
wire S2682;
wire S2683;
wire S2684;
wire S2685;
wire S2686;
wire S2687;
wire S2688;
wire S2689;
wire S2690;
wire S2691;
wire S2692;
wire S2693;
wire S2694;
wire S2695;
wire S2696;
wire S2697;
wire S2698;
wire S2699;
wire S2700;
wire S2701;
wire S2702;
wire S2703;
wire S2704;
wire S2705;
wire S2706;
wire S2707;
wire S2708;
wire S2709;
wire S2710;
wire S2711;
wire S2712;
wire S2713;
wire S2714;
wire S2715;
wire S2716;
wire S2717;
wire S2718;
wire S2719;
wire S2720;
wire S2721;
wire S2722;
wire S2723;
wire S2724;
wire S2725;
wire S2726;
wire S2727;
wire S2728;
wire S2729;
wire S2730;
wire S2731;
wire S2732;
wire S2733;
wire S2734;
wire S2735;
wire S2736;
wire S2737;
wire S2738;
wire S2739;
wire S2740;
wire S2741;
wire S2742;
wire S2743;
wire S2744;
wire S2745;
wire S2746;
wire S2747;
wire S2748;
wire S2749;
wire S2750;
wire S2751;
wire S2752;
wire S2753;
wire S2754;
wire S2755;
wire S2756;
wire S2757;
wire S2758;
wire S2759;
wire S2760;
wire S2761;
wire S2762;
wire S2763;
wire S2764;
wire S2765;
wire S2766;
wire S2767;
wire S2768;
wire S2769;
wire S2770;
wire S2771;
wire S2772;
wire S2773;
wire S2774;
wire S2775;
wire S2776;
wire S2777;
wire S2778;
wire S2779;
wire S2780;
wire S2781;
wire S2782;
wire S2783;
wire S2784;
wire S2785;
wire S2786;
wire S2787;
wire S2788;
wire S2789;
wire S2790;
wire S2791;
wire S2792;
wire S2793;
wire S2794;
wire S2795;
wire S2796;
wire S2797;
wire S2798;
wire S2799;
wire S2800;
wire S2801;
wire S2802;
wire S2803;
wire S2804;
wire S2805;
wire S2806;
wire S2807;
wire S2808;
wire S2809;
wire S2810;
wire S2811;
wire S2812;
wire S2813;
wire S2814;
wire S2815;
wire S2816;
wire S2817;
wire S2818;
wire S2819;
wire S2820;
wire S2821;
wire S2822;
wire S2823;
wire S2824;
wire S2825;
wire S2826;
wire S2827;
wire S2828;
wire S2829;
wire S2830;
wire S2831;
wire S2832;
wire S2833;
wire S2834;
wire S2835;
wire S2836;
wire S2837;
wire S2838;
wire S2839;
wire S2840;
wire S2841;
wire S2842;
wire S2843;
wire S2844;
wire S2845;
wire S2846;
wire S2847;
wire S2848;
wire S2849;
wire S2850;
wire S2851;
wire S2852;
wire S2853;
wire S2854;
wire S2855;
wire S2856;
wire S2857;
wire S2858;
wire S2859;
wire S2860;
wire S2861;
wire S2862;
wire S2863;
wire S2864;
wire S2865;
wire S2866;
wire S2867;
wire S2868;
wire S2869;
wire S2870;
wire S2871;
wire S2872;
wire S2873;
wire S2874;
wire S2875;
wire S2876;
wire S2877;
wire S2878;
wire S2879;
wire S2880;
wire S2881;
wire S2882;
wire S2883;
wire S2884;
wire S2885;
wire S2886;
wire S2887;
wire S2888;
wire S2889;
wire S2890;
wire S2891;
wire S2892;
wire S2893;
wire S2894;
wire S2895;
wire S2896;
wire S2897;
wire S2898;
wire S2899;
wire S2900;
wire S2901;
wire S2902;
wire S2903;
wire S2904;
wire S2905;
wire S2906;
wire S2907;
wire S2908;
wire S2909;
wire S2910;
wire S2911;
wire S2912;
wire S2913;
wire S2914;
wire S2915;
wire S2916;
wire S2917;
wire S2918;
wire S2919;
wire S2920;
wire S2921;
wire S2922;
wire S2923;
wire S2924;
wire S2925;
wire S2926;
wire S2927;
wire S2928;
wire S2929;
wire S2930;
wire S2931;
wire S2932;
wire S2933;
wire S2934;
wire S2935;
wire S2936;
wire S2937;
wire S2938;
wire S2939;
wire S2940;
wire S2941;
wire S2942;
wire S2943;
wire S2944;
wire S2945;
wire S2946;
wire S2947;
wire S2948;
wire S2949;
wire S2950;
wire S2951;
wire S2952;
wire S2953;
wire S2954;
wire S2955;
wire S2956;
wire S2957;
wire S2958;
wire S2959;
wire S2960;
wire S2961;
wire S2962;
wire S2963;
wire S2964;
wire S2965;
wire S2966;
wire S2967;
wire S2968;
wire S2969;
wire S2970;
wire S2971;
wire S2972;
wire S2973;
wire S2974;
wire S2975;
wire S2976;
wire S2977;
wire S2978;
wire S2979;
wire S2980;
wire S2981;
wire S2982;
wire S2983;
wire S2984;
wire S2985;
wire S2986;
wire S2987;
wire S2988;
wire S2989;
wire S2990;
wire S2991;
wire S2992;
wire S2993;
wire S2994;
wire S2995;
wire S2996;
wire S2997;
wire S2998;
wire S2999;
wire S3000;
wire S3001;
wire S3002;
wire S3003;
wire S3004;
wire S3005;
wire S3006;
wire S3007;
wire S3008;
wire S3009;
wire S3010;
wire S3011;
wire S3012;
wire S3013;
wire S3014;
wire S3015;
wire S3016;
wire S3017;
wire S3018;
wire S3019;
wire S3020;
wire S3021;
wire S3022;
wire S3023;
wire S3024;
wire S3025;
wire S3026;
wire S3027;
wire S3028;
wire S3029;
wire S3030;
wire S3031;
wire S3032;
wire S3033;
wire S3034;
wire S3035;
wire S3036;
wire S3037;
wire S3038;
wire S3039;
wire S3040;
wire S3041;
wire S3042;
wire S3043;
wire S3044;
wire S3045;
wire S3046;
wire S3047;
wire S3048;
wire S3049;
wire S3050;
wire S3051;
wire S3052;
wire S3053;
wire S3054;
wire S3055;
wire S3056;
wire S3057;
wire S3058;
wire S3059;
wire S3060;
wire S3061;
wire S3062;
wire S3063;
wire S3064;
wire S3065;
wire S3066;
wire S3067;
wire S3068;
wire S3069;
wire S3070;
wire S3071;
wire S3072;
wire S3073;
wire S3074;
wire S3075;
wire S3076;
wire S3077;
wire S3078;
wire S3079;
wire S3080;
wire S3081;
wire S3082;
wire S3083;
wire S3084;
wire S3085;
wire S3086;
wire S3087;
wire S3088;
wire S3089;
wire S3090;
wire S3091;
wire S3092;
wire S3093;
wire S3094;
wire S3095;
wire S3096;
wire S3097;
wire S3098;
wire S3099;
wire S3100;
wire S3101;
wire CU_ADD;
wire CU_AND;
wire CU_INC1;
wire CU_INC2;
wire CU_LSB0E;
wire CU_MUL;
wire CU_NOT;
wire CU_SE12bits;
wire CU_SE4bits;
wire CU_SHF_0;
wire CU_SHF_1;
wire CU_clk;
wire CU_conOF;
wire CU_enSKP;
wire CU_inst_0;
wire CU_inst_10;
wire CU_inst_11;
wire CU_inst_12;
wire CU_inst_13;
wire CU_inst_14;
wire CU_inst_15;
wire CU_inst_1;
wire CU_inst_2;
wire CU_inst_3;
wire CU_inst_4;
wire CU_inst_5;
wire CU_inst_6;
wire CU_inst_7;
wire CU_inst_8;
wire CU_inst_9;
wire CU_ldAC;
wire CU_ldIN;
wire CU_ldIR;
wire CU_ldOF;
wire CU_ldPC;
wire CU_ldSR_0;
wire CU_ldSR_1;
wire CU_ldSR_2;
wire CU_ldSR_3;
wire CU_nstate_0;
wire CU_nstate_1;
wire CU_pstate_0;
wire CU_pstate_1;
wire CU_readMEM;
wire CU_rst;
wire CU_sel1_ARU;
wire CU_selAC_MEM;
wire CU_selARU_AC;
wire CU_selARU_SR;
wire CU_selIMM_AC;
wire CU_selIMM_LGU;
wire CU_selIMM_OF;
wire CU_selIMM_PC;
wire CU_selINC_IN;
wire CU_selINC_PC;
wire CU_selIN_ADR;
wire CU_selIN_MEM;
wire CU_selIR_ADR;
wire CU_selLGU_AC;
wire CU_selLGU_SR;
wire CU_selMEM_AC;
wire CU_selMEM_IN;
wire CU_selMEM_LGU;
wire CU_selMEM_PC;
wire CU_selPC_MEM;
wire CU_selPC_OF;
wire CU_selSET_SR;
wire CU_seldataBus;
wire CU_zeroAC;
wire DP_AC_din_0;
wire DP_AC_din_10;
wire DP_AC_din_11;
wire DP_AC_din_12;
wire DP_AC_din_13;
wire DP_AC_din_14;
wire DP_AC_din_15;
wire DP_AC_din_1;
wire DP_AC_din_2;
wire DP_AC_din_3;
wire DP_AC_din_4;
wire DP_AC_din_5;
wire DP_AC_din_6;
wire DP_AC_din_7;
wire DP_AC_din_8;
wire DP_AC_din_9;
wire DP_AC_dout_0;
wire DP_AC_dout_10;
wire DP_AC_dout_11;
wire DP_AC_dout_12;
wire DP_AC_dout_13;
wire DP_AC_dout_14;
wire DP_AC_dout_15;
wire DP_AC_dout_1;
wire DP_AC_dout_2;
wire DP_AC_dout_3;
wire DP_AC_dout_4;
wire DP_AC_dout_5;
wire DP_AC_dout_6;
wire DP_AC_dout_7;
wire DP_AC_dout_8;
wire DP_AC_dout_9;
wire DP_ARU1_C;
wire DP_ARU1_N;
wire DP_ARU1_V;
wire DP_ARU1_Z;
wire DP_ARU1_in1_0;
wire DP_ARU1_in1_10;
wire DP_ARU1_in1_11;
wire DP_ARU1_in1_12;
wire DP_ARU1_in1_13;
wire DP_ARU1_in1_14;
wire DP_ARU1_in1_15;
wire DP_ARU1_in1_1;
wire DP_ARU1_in1_2;
wire DP_ARU1_in1_3;
wire DP_ARU1_in1_4;
wire DP_ARU1_in1_5;
wire DP_ARU1_in1_6;
wire DP_ARU1_in1_7;
wire DP_ARU1_in1_8;
wire DP_ARU1_in1_9;
wire DP_ARU1_out_0;
wire DP_ARU1_out_10;
wire DP_ARU1_out_11;
wire DP_ARU1_out_12;
wire DP_ARU1_out_13;
wire DP_ARU1_out_14;
wire DP_ARU1_out_1;
wire DP_ARU1_out_2;
wire DP_ARU1_out_3;
wire DP_ARU1_out_4;
wire DP_ARU1_out_5;
wire DP_ARU1_out_6;
wire DP_ARU1_out_7;
wire DP_ARU1_out_8;
wire DP_ARU1_out_9;
wire DP_IMM1_in1_0;
wire DP_IMM1_in1_1;
wire DP_IMM1_in1_2;
wire DP_IMM1_in1_3;
wire DP_IMM1_out_0;
wire DP_IMM1_out_10;
wire DP_IMM1_out_11;
wire DP_IMM1_out_12;
wire DP_IMM1_out_13;
wire DP_IMM1_out_14;
wire DP_IMM1_out_15;
wire DP_IMM1_out_1;
wire DP_IMM1_out_2;
wire DP_IMM1_out_3;
wire DP_IMM1_out_4;
wire DP_IMM1_out_5;
wire DP_IMM1_out_6;
wire DP_IMM1_out_7;
wire DP_IMM1_out_8;
wire DP_IMM1_out_9;
wire DP_IN_din_0;
wire DP_IN_din_10;
wire DP_IN_din_11;
wire DP_IN_din_12;
wire DP_IN_din_13;
wire DP_IN_din_14;
wire DP_IN_din_15;
wire DP_IN_din_1;
wire DP_IN_din_2;
wire DP_IN_din_3;
wire DP_IN_din_4;
wire DP_IN_din_5;
wire DP_IN_din_6;
wire DP_IN_din_7;
wire DP_IN_din_8;
wire DP_IN_din_9;
wire DP_IN_dout_0;
wire DP_IN_dout_10;
wire DP_IN_dout_11;
wire DP_IN_dout_12;
wire DP_IN_dout_13;
wire DP_IN_dout_14;
wire DP_IN_dout_15;
wire DP_IN_dout_1;
wire DP_IN_dout_2;
wire DP_IN_dout_3;
wire DP_IN_dout_4;
wire DP_IN_dout_5;
wire DP_IN_dout_6;
wire DP_IN_dout_7;
wire DP_IN_dout_8;
wire DP_IN_dout_9;
wire DP_INC2_out_0;
wire DP_INC2_out_10;
wire DP_INC2_out_11;
wire DP_INC2_out_12;
wire DP_INC2_out_13;
wire DP_INC2_out_14;
wire DP_INC2_out_15;
wire DP_INC2_out_1;
wire DP_INC2_out_2;
wire DP_INC2_out_3;
wire DP_INC2_out_4;
wire DP_INC2_out_5;
wire DP_INC2_out_6;
wire DP_INC2_out_7;
wire DP_INC2_out_8;
wire DP_INC2_out_9;
wire DP_INC_1_in_0;
wire DP_INC_1_in_10;
wire DP_INC_1_in_11;
wire DP_INC_1_in_12;
wire DP_INC_1_in_13;
wire DP_INC_1_in_14;
wire DP_INC_1_in_15;
wire DP_INC_1_in_1;
wire DP_INC_1_in_2;
wire DP_INC_1_in_3;
wire DP_INC_1_in_4;
wire DP_INC_1_in_5;
wire DP_INC_1_in_6;
wire DP_INC_1_in_7;
wire DP_INC_1_in_8;
wire DP_INC_1_in_9;
wire DP_INC_1_inc_value_0;
wire DP_INC_1_inc_value_1;
wire DP_INC_1_out_0;
wire DP_INC_1_out_10;
wire DP_INC_1_out_11;
wire DP_INC_1_out_12;
wire DP_INC_1_out_13;
wire DP_INC_1_out_14;
wire DP_INC_1_out_15;
wire DP_INC_1_out_1;
wire DP_INC_1_out_2;
wire DP_INC_1_out_3;
wire DP_INC_1_out_4;
wire DP_INC_1_out_5;
wire DP_INC_1_out_6;
wire DP_INC_1_out_7;
wire DP_INC_1_out_8;
wire DP_INC_1_out_9;
wire DP_LGU1_N;
wire DP_LGU1_Z;
wire DP_LGU1_in1_0;
wire DP_LGU1_in1_10;
wire DP_LGU1_in1_11;
wire DP_LGU1_in1_12;
wire DP_LGU1_in1_13;
wire DP_LGU1_in1_14;
wire DP_LGU1_in1_15;
wire DP_LGU1_in1_1;
wire DP_LGU1_in1_2;
wire DP_LGU1_in1_3;
wire DP_LGU1_in1_4;
wire DP_LGU1_in1_5;
wire DP_LGU1_in1_6;
wire DP_LGU1_in1_7;
wire DP_LGU1_in1_8;
wire DP_LGU1_in1_9;
wire DP_LGU1_out_0;
wire DP_LGU1_out_10;
wire DP_LGU1_out_11;
wire DP_LGU1_out_12;
wire DP_LGU1_out_13;
wire DP_LGU1_out_14;
wire DP_LGU1_out_1;
wire DP_LGU1_out_2;
wire DP_LGU1_out_3;
wire DP_LGU1_out_4;
wire DP_LGU1_out_5;
wire DP_LGU1_out_6;
wire DP_LGU1_out_7;
wire DP_LGU1_out_8;
wire DP_LGU1_out_9;
wire DP_OF_din_0;
wire DP_OF_din_1;
wire DP_OF_din_2;
wire DP_OF_din_3;
wire DP_PC_din_0;
wire DP_PC_din_10;
wire DP_PC_din_11;
wire DP_PC_din_12;
wire DP_PC_din_13;
wire DP_PC_din_14;
wire DP_PC_din_15;
wire DP_PC_din_1;
wire DP_PC_din_2;
wire DP_PC_din_3;
wire DP_PC_din_4;
wire DP_PC_din_5;
wire DP_PC_din_6;
wire DP_PC_din_7;
wire DP_PC_din_8;
wire DP_PC_din_9;
wire DP_SR_C_din;
wire DP_SR_C_dout;
wire DP_SR_N_din;
wire DP_SR_N_dout;
wire DP_SR_V_din;
wire DP_SR_V_dout;
wire DP_SR_Z_din;
wire DP_SR_Z_dout;
wire DP_addrBus_0;
wire DP_addrBus_10;
wire DP_addrBus_11;
wire DP_addrBus_12;
wire DP_addrBus_13;
wire DP_addrBus_14;
wire DP_addrBus_15;
wire DP_addrBus_1;
wire DP_addrBus_2;
wire DP_addrBus_3;
wire DP_addrBus_4;
wire DP_addrBus_5;
wire DP_addrBus_6;
wire DP_addrBus_7;
wire DP_addrBus_8;
wire DP_addrBus_9;
input clk;
input rst;
output writeMEM;
output readMEM;
output [15:0] addrBus;
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_1_ (
  .in1({ 1'b1 }),
  .out1({ S0 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_2_ (
  .in1({ 1'b1 }),
  .out1({ S1 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_3_ (
  .in1({ 1'b1 }),
  .out1({ S2 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_4_ (
  .in1({ 1'b1 }),
  .out1({ S3 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_5_ (
  .in1({ 1'b1 }),
  .out1({ S4 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_6_ (
  .in1({ 1'b1 }),
  .out1({ S5 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_7_ (
  .in1({ 1'b0 }),
  .out1({ S6 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_8_ (
  .in1({ 1'b0 }),
  .out1({ S7 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_9_ (
  .in1({ 1'b0 }),
  .out1({ S8 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_10_ (
  .in1({ 1'b0 }),
  .out1({ S9 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_11_ (
  .in1({ 1'b0 }),
  .out1({ S10 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_12_ (
  .in1({ 1'b0 }),
  .out1({ S11 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_13_ (
  .in1({ 1'b0 }),
  .out1({ S12 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_14_ (
  .in1({ 1'b0 }),
  .out1({ S13 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_15_ (
  .in1({ 1'b0 }),
  .out1({ S14 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_16_ (
  .in1({ 1'b0 }),
  .out1({ S15 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_17_ (
  .in1({ 1'b0 }),
  .out1({ S16 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_18_ (
  .in1({ 1'b0 }),
  .out1({ S17 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_19_ (
  .in1({ 1'b0 }),
  .out1({ S18 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_20_ (
  .in1({ 1'b0 }),
  .out1({ S19 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_21_ (
  .in1({ 1'b0 }),
  .out1({ S20 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_22_ (
  .in1({ 1'b0 }),
  .out1({ S21 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_23_ (
  .in1({ 1'b0 }),
  .out1({ S22 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_24_ (
  .in1({ 1'b0 }),
  .out1({ S23 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_25_ (
  .in1({ 1'b0 }),
  .out1({ S24 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_26_ (
  .in1({ 1'b0 }),
  .out1({ S25 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_27_ (
  .in1({ 1'b0 }),
  .out1({ S26 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_28_ (
  .in1({ 1'b0 }),
  .out1({ S27 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_29_ (
  .in1({ 1'b0 }),
  .out1({ S28 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_30_ (
  .in1({ 1'b0 }),
  .out1({ S29 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_31_ (
  .in1({ 1'b0 }),
  .out1({ S30 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_32_ (
  .in1({ 1'b0 }),
  .out1({ S31 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_33_ (
  .in1({ 1'b0 }),
  .out1({ S32 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_34_ (
  .in1({ 1'b0 }),
  .out1({ S33 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_35_ (
  .in1({ 1'b0 }),
  .out1({ S34 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_36_ (
  .in1({ 1'b0 }),
  .out1({ S35 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_37_ (
  .in1({ 1'b0 }),
  .out1({ S36 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_38_ (
  .in1({ 1'b0 }),
  .out1({ S37 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_1_ (
  .in1({ CU_pstate_1 }),
  .out1({ S207 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_2_ (
  .in1({ CU_pstate_0 }),
  .out1({ S208 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_3_ (
  .in1({ CU_inst_9 }),
  .out1({ S209 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_4_ (
  .in1({ CU_inst_8 }),
  .out1({ S210 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_5_ (
  .in1({ CU_inst_10 }),
  .out1({ S211 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_6_ (
  .in1({ CU_inst_13 }),
  .out1({ S212 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_7_ (
  .in1({ CU_inst_12 }),
  .out1({ S213 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_8_ (
  .in1({ CU_inst_14 }),
  .out1({ S214 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_9_ (
  .in1({ CU_inst_15 }),
  .out1({ S215 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_10_ (
  .in1({ CU_inst_5 }),
  .out1({ S216 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_11_ (
  .in1({ CU_inst_6 }),
  .out1({ S217 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_12_ (
  .in1({ CU_inst_7 }),
  .out1({ S218 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_13_ (
  .in1({ CU_enSKP }),
  .out1({ S219 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1_ (
  .in1({ CU_pstate_0, CU_pstate_1 }),
  .out1({ CU_ldIR })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_14_ (
  .in1({ CU_ldIR }),
  .out1({ S220 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_2_ (
  .in1({ S208, CU_pstate_1 }),
  .out1({ S221 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1_ (
  .in1({ CU_pstate_0, S207 }),
  .out1({ S222 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_3_ (
  .in1({ S215, S214 }),
  .out1({ S223 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_2_ (
  .in1({ CU_inst_15, CU_inst_14 }),
  .out1({ S224 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_3_ (
  .in1({ CU_inst_12, CU_inst_13 }),
  .out1({ S225 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_15_ (
  .in1({ S225 }),
  .out1({ S226 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_4_ (
  .in1({ S225, S224 }),
  .out1({ S227 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_4_ (
  .in1({ S226, S223 }),
  .out1({ S228 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_5_ (
  .in1({ S228, S222 }),
  .out1({ S229 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_5_ (
  .in1({ S227, S221 }),
  .out1({ S230 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_6_ (
  .in1({ S211, CU_inst_11 }),
  .out1({ S231 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_7_ (
  .in1({ CU_inst_8, CU_inst_9 }),
  .out1({ S232 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_6_ (
  .in1({ S232, S231 }),
  .out1({ S233 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_8_ (
  .in1({ S233, S230 }),
  .out1({ CU_SHF_0 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_9_ (
  .in1({ CU_inst_10, CU_inst_11 }),
  .out1({ S234 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_16_ (
  .in1({ S234 }),
  .out1({ S235 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_7_ (
  .in1({ S234, CU_inst_9 }),
  .out1({ S236 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_17_ (
  .in1({ S236 }),
  .out1({ S237 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_8_ (
  .in1({ S237, CU_inst_8 }),
  .out1({ S238 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_10_ (
  .in1({ S238, S230 }),
  .out1({ CU_SHF_1 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_11_ (
  .in1({ CU_inst_15, CU_inst_14 }),
  .out1({ S38 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_9_ (
  .in1({ S215, S214 }),
  .out1({ S39 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_12_ (
  .in1({ CU_pstate_0, S207 }),
  .out1({ S40 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_10_ (
  .in1({ S208, CU_pstate_1 }),
  .out1({ S41 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_13_ (
  .in1({ CU_inst_12, S212 }),
  .out1({ S42 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_11_ (
  .in1({ S213, CU_inst_13 }),
  .out1({ S43 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_14_ (
  .in1({ S43, S41 }),
  .out1({ S44 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_12_ (
  .in1({ S42, S40 }),
  .out1({ S45 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_13_ (
  .in1({ CU_inst_12, S212 }),
  .out1({ S46 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_15_ (
  .in1({ S46, S222 }),
  .out1({ S47 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_18_ (
  .in1({ S47 }),
  .out1({ S48 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_16_ (
  .in1({ S47, S44 }),
  .out1({ S49 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_14_ (
  .in1({ S44, S38 }),
  .out1({ S50 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_17_ (
  .in1({ S49, S39 }),
  .out1({ CU_selMEM_AC })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_18_ (
  .in1({ S45, CU_inst_14 }),
  .out1({ S51 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_19_ (
  .in1({ S51 }),
  .out1({ S52 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_19_ (
  .in1({ S215, CU_inst_14 }),
  .out1({ S53 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_15_ (
  .in1({ CU_inst_15, S214 }),
  .out1({ S54 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_20_ (
  .in1({ S54, S45 }),
  .out1({ S55 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_16_ (
  .in1({ S53, S44 }),
  .out1({ S56 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_21_ (
  .in1({ S54, CU_inst_13 }),
  .out1({ S57 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_20_ (
  .in1({ S57 }),
  .out1({ S58 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_22_ (
  .in1({ S58, S222 }),
  .out1({ S59 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_23_ (
  .in1({ S59, S55 }),
  .out1({ S60 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_24_ (
  .in1({ CU_inst_8, S209 }),
  .out1({ S61 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_17_ (
  .in1({ S61, S231 }),
  .out1({ S62 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_25_ (
  .in1({ S62, S228 }),
  .out1({ S63 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_21_ (
  .in1({ S63 }),
  .out1({ S64 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_26_ (
  .in1({ S64, S222 }),
  .out1({ CU_selSET_SR })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_18_ (
  .in1({ CU_selSET_SR, CU_inst_4 }),
  .out1({ S65 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_19_ (
  .in1({ S65, S60 }),
  .out1({ CU_ldSR_0 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_20_ (
  .in1({ CU_selSET_SR, CU_inst_5 }),
  .out1({ S66 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_21_ (
  .in1({ S66, S60 }),
  .out1({ CU_ldSR_1 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_22_ (
  .in1({ S63, CU_inst_6 }),
  .out1({ S67 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_22_ (
  .in1({ S67 }),
  .out1({ S68 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_27_ (
  .in1({ S210, CU_inst_9 }),
  .out1({ S69 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_23_ (
  .in1({ CU_inst_8, S209 }),
  .out1({ S70 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_28_ (
  .in1({ S70, S235 }),
  .out1({ S71 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_24_ (
  .in1({ S69, S234 }),
  .out1({ S72 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_25_ (
  .in1({ S218, CU_inst_6 }),
  .out1({ S73 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_29_ (
  .in1({ S72, S217 }),
  .out1({ S74 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_30_ (
  .in1({ CU_inst_7, S216 }),
  .out1({ S75 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_26_ (
  .in1({ S75, S74 }),
  .out1({ S76 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_31_ (
  .in1({ S73, S72 }),
  .out1({ S77 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_27_ (
  .in1({ S77, S227 }),
  .out1({ S78 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_32_ (
  .in1({ S68, S57 }),
  .out1({ S79 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_28_ (
  .in1({ S79, S78 }),
  .out1({ S80 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_29_ (
  .in1({ S80, S221 }),
  .out1({ S81 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_33_ (
  .in1({ CU_inst_15, S214 }),
  .out1({ S82 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_30_ (
  .in1({ S215, CU_inst_14 }),
  .out1({ S83 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_31_ (
  .in1({ CU_inst_14, CU_inst_13 }),
  .out1({ S84 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_34_ (
  .in1({ S84, CU_inst_15 }),
  .out1({ S85 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_32_ (
  .in1({ S82, CU_inst_13 }),
  .out1({ S86 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_35_ (
  .in1({ S86, S222 }),
  .out1({ CU_AND })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_36_ (
  .in1({ CU_AND, S55 }),
  .out1({ S87 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_33_ (
  .in1({ S87, S81 }),
  .out1({ CU_ldSR_2 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_34_ (
  .in1({ S53, S43 }),
  .out1({ S88 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_37_ (
  .in1({ S88, S222 }),
  .out1({ S89 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_23_ (
  .in1({ S89 }),
  .out1({ S90 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_35_ (
  .in1({ S90, S56 }),
  .out1({ CU_selARU_SR })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_36_ (
  .in1({ S63, CU_inst_7 }),
  .out1({ S91 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_37_ (
  .in1({ S91, S88 }),
  .out1({ S92 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_38_ (
  .in1({ S92, S85 }),
  .out1({ S93 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_38_ (
  .in1({ S93, S78 }),
  .out1({ S94 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_39_ (
  .in1({ S94, S221 }),
  .out1({ S95 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_40_ (
  .in1({ S95, S56 }),
  .out1({ CU_ldSR_3 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_41_ (
  .in1({ S83, S43 }),
  .out1({ S96 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_42_ (
  .in1({ S96, S84 }),
  .out1({ S97 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_39_ (
  .in1({ S224, CU_inst_12 }),
  .out1({ S98 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_43_ (
  .in1({ S223, S213 }),
  .out1({ S99 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_44_ (
  .in1({ S42, S223 }),
  .out1({ S100 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_24_ (
  .in1({ S100 }),
  .out1({ S101 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_45_ (
  .in1({ S100, S97 }),
  .out1({ S102 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_25_ (
  .in1({ S102 }),
  .out1({ S103 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_40_ (
  .in1({ S103, S41 }),
  .out1({ S104 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_46_ (
  .in1({ S102, S40 }),
  .out1({ S105 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_47_ (
  .in1({ S97, S221 }),
  .out1({ S106 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_26_ (
  .in1({ S106 }),
  .out1({ S107 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_48_ (
  .in1({ S106, S105 }),
  .out1({ CU_ldPC })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_41_ (
  .in1({ S224, CU_inst_13 }),
  .out1({ S108 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_27_ (
  .in1({ S108 }),
  .out1({ S109 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_42_ (
  .in1({ S39, S213 }),
  .out1({ S110 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_49_ (
  .in1({ S43, S38 }),
  .out1({ S111 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_50_ (
  .in1({ S111, S100 }),
  .out1({ S112 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_28_ (
  .in1({ S112 }),
  .out1({ S113 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_43_ (
  .in1({ S108, S106 }),
  .out1({ S114 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_29_ (
  .in1({ S114 }),
  .out1({ S115 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_44_ (
  .in1({ S115, S112 }),
  .out1({ S116 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_51_ (
  .in1({ S114, S113 }),
  .out1({ S117 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_45_ (
  .in1({ CU_inst_6, CU_inst_5 }),
  .out1({ S118 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_30_ (
  .in1({ S118 }),
  .out1({ S119 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_46_ (
  .in1({ S119, S218 }),
  .out1({ S120 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_52_ (
  .in1({ S118, CU_inst_7 }),
  .out1({ S121 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_47_ (
  .in1({ S121, S72 }),
  .out1({ S122 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_53_ (
  .in1({ S120, S71 }),
  .out1({ S123 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_54_ (
  .in1({ S123, S227 }),
  .out1({ S124 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_55_ (
  .in1({ S124, S86 }),
  .out1({ S125 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_48_ (
  .in1({ S125, S117 }),
  .out1({ S126 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_49_ (
  .in1({ S126, S55 }),
  .out1({ S127 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_31_ (
  .in1({ S127 }),
  .out1({ CU_selARU_AC })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_50_ (
  .in1({ S54, S225 }),
  .out1({ S128 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_32_ (
  .in1({ S128 }),
  .out1({ S129 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_51_ (
  .in1({ S128, S127 }),
  .out1({ CU_ADD })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_56_ (
  .in1({ S236, S233 }),
  .out1({ S130 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_52_ (
  .in1({ S130, S228 }),
  .out1({ S131 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_57_ (
  .in1({ S131, S76 }),
  .out1({ S132 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_33_ (
  .in1({ S132 }),
  .out1({ S133 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_53_ (
  .in1({ S132, S122 }),
  .out1({ S134 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_54_ (
  .in1({ S39, S225 }),
  .out1({ S135 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_55_ (
  .in1({ S135, S101 }),
  .out1({ S136 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_58_ (
  .in1({ S136, S109 }),
  .out1({ S137 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_56_ (
  .in1({ S137, S134 }),
  .out1({ S138 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_59_ (
  .in1({ S138, S107 }),
  .out1({ S139 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_60_ (
  .in1({ S139, S52 }),
  .out1({ CU_ldAC })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_57_ (
  .in1({ CU_inst_12, CU_inst_13 }),
  .out1({ S140 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_58_ (
  .in1({ S83, S41 }),
  .out1({ S141 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_61_ (
  .in1({ S141, S140 }),
  .out1({ S142 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_62_ (
  .in1({ S135, S221 }),
  .out1({ S143 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_63_ (
  .in1({ S143, S142 }),
  .out1({ CU_selAC_MEM })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_59_ (
  .in1({ S100, S222 }),
  .out1({ CU_selPC_MEM })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_34_ (
  .in1({ CU_selPC_MEM }),
  .out1({ S144 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_60_ (
  .in1({ S83, S46 }),
  .out1({ S145 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_64_ (
  .in1({ S145, S40 }),
  .out1({ S146 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_35_ (
  .in1({ S146 }),
  .out1({ S147 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_61_ (
  .in1({ S147, CU_selAC_MEM }),
  .out1({ S148 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_65_ (
  .in1({ S148, S144 }),
  .out1({ CU_seldataBus })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_62_ (
  .in1({ S223, S222 }),
  .out1({ S149 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_66_ (
  .in1({ S149, S111 }),
  .out1({ S150 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_63_ (
  .in1({ S85, S57 }),
  .out1({ S151 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_64_ (
  .in1({ S151, CU_inst_12 }),
  .out1({ S152 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_67_ (
  .in1({ S111, S224 }),
  .out1({ S153 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_36_ (
  .in1({ S153 }),
  .out1({ S154 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_65_ (
  .in1({ S152, S106 }),
  .out1({ S155 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_66_ (
  .in1({ S99, CU_inst_13 }),
  .out1({ S156 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_68_ (
  .in1({ S155, S154 }),
  .out1({ S157 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_69_ (
  .in1({ S157, S56 }),
  .out1({ CU_selMEM_LGU })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_70_ (
  .in1({ S75, S217 }),
  .out1({ S158 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_67_ (
  .in1({ S158, S72 }),
  .out1({ S159 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_71_ (
  .in1({ S159, S227 }),
  .out1({ S160 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_72_ (
  .in1({ S71, S227 }),
  .out1({ S161 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_68_ (
  .in1({ S161, S158 }),
  .out1({ S162 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_69_ (
  .in1({ S162, S98 }),
  .out1({ S163 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_70_ (
  .in1({ S46, S224 }),
  .out1({ S164 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_73_ (
  .in1({ S108, CU_inst_12 }),
  .out1({ S165 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_71_ (
  .in1({ S164, S106 }),
  .out1({ S166 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_74_ (
  .in1({ S166, S163 }),
  .out1({ S167 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_75_ (
  .in1({ S167, S105 }),
  .out1({ CU_selINC_PC })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_76_ (
  .in1({ S211, CU_inst_11 }),
  .out1({ S168 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_72_ (
  .in1({ S168, S219 }),
  .out1({ S169 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_77_ (
  .in1({ S169, S69 }),
  .out1({ S170 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_78_ (
  .in1({ S170, S227 }),
  .out1({ S171 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_73_ (
  .in1({ S171, S159 }),
  .out1({ S172 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_79_ (
  .in1({ S129, S113 }),
  .out1({ S173 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_74_ (
  .in1({ S173, S172 }),
  .out1({ S174 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_75_ (
  .in1({ S174, S222 }),
  .out1({ S175 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_76_ (
  .in1({ S175, CU_AND }),
  .out1({ S176 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_77_ (
  .in1({ S104, S59 }),
  .out1({ S177 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_80_ (
  .in1({ S177, S176 }),
  .out1({ CU_INC1 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_81_ (
  .in1({ S140, S38 }),
  .out1({ S178 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_82_ (
  .in1({ S228, S221 }),
  .out1({ S179 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_78_ (
  .in1({ S179, S152 }),
  .out1({ S180 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_83_ (
  .in1({ S180, S178 }),
  .out1({ S181 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_79_ (
  .in1({ S181, S156 }),
  .out1({ S182 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_37_ (
  .in1({ S182 }),
  .out1({ S183 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_84_ (
  .in1({ S183, S146 }),
  .out1({ CU_selIR_ADR })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_85_ (
  .in1({ S182, S136 }),
  .out1({ S184 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_80_ (
  .in1({ S51, CU_ldIR }),
  .out1({ S185 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_86_ (
  .in1({ S185, S184 }),
  .out1({ CU_readMEM })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_81_ (
  .in1({ S220, CU_rst }),
  .out1({ CU_nstate_0 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_82_ (
  .in1({ S103, S222 }),
  .out1({ CU_nstate_1 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_87_ (
  .in1({ S181, S146 }),
  .out1({ CU_conOF })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_88_ (
  .in1({ S116, S88 }),
  .out1({ S186 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_83_ (
  .in1({ S77, S228 }),
  .out1({ S187 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_84_ (
  .in1({ S187, S186 }),
  .out1({ CU_selLGU_SR })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_85_ (
  .in1({ S170, S230 }),
  .out1({ CU_INC2 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_86_ (
  .in1({ S83, S48 }),
  .out1({ CU_selINC_IN })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_87_ (
  .in1({ S129, S222 }),
  .out1({ CU_MUL })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_88_ (
  .in1({ S76, S230 }),
  .out1({ CU_NOT })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_89_ (
  .in1({ S160, S222 }),
  .out1({ CU_LSB0E })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_89_ (
  .in1({ S86, S54 }),
  .out1({ S188 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_90_ (
  .in1({ S188, CU_inst_12 }),
  .out1({ S189 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_91_ (
  .in1({ S189, S109 }),
  .out1({ S190 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_90_ (
  .in1({ S179, S110 }),
  .out1({ S191 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_92_ (
  .in1({ S191, S103 }),
  .out1({ S192 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_91_ (
  .in1({ S192, S190 }),
  .out1({ CU_SE4bits })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_93_ (
  .in1({ S234, S232 }),
  .out1({ S193 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_38_ (
  .in1({ S193 }),
  .out1({ S194 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_94_ (
  .in1({ S194, S229 }),
  .out1({ S195 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_39_ (
  .in1({ S195 }),
  .out1({ CU_selIMM_OF })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_95_ (
  .in1({ S130, S229 }),
  .out1({ S196 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_96_ (
  .in1({ S196, S195 }),
  .out1({ CU_SE12bits })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_92_ (
  .in1({ S186, S133 }),
  .out1({ CU_selLGU_AC })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_93_ (
  .in1({ S178, S222 }),
  .out1({ CU_selIMM_AC })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_97_ (
  .in1({ S142, S50 }),
  .out1({ CU_selIN_ADR })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_98_ (
  .in1({ S146, S56 }),
  .out1({ CU_selIN_MEM })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_94_ (
  .in1({ S163, S222 }),
  .out1({ CU_selIMM_PC })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_95_ (
  .in1({ S165, S222 }),
  .out1({ CU_selMEM_PC })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_96_ (
  .in1({ S123, S230 }),
  .out1({ CU_sel1_ARU })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_97_ (
  .in1({ S131, S112 }),
  .out1({ S197 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_99_ (
  .in1({ S197, S107 }),
  .out1({ S198 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_98_ (
  .in1({ S198, S190 }),
  .out1({ CU_selIMM_LGU })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_99_ (
  .in1({ S140, S83 }),
  .out1({ S199 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_40_ (
  .in1({ S199 }),
  .out1({ S200 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_100_ (
  .in1({ S200, S88 }),
  .out1({ S201 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_100_ (
  .in1({ S201, S150 }),
  .out1({ CU_selMEM_IN })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_101_ (
  .in1({ S118, S218 }),
  .out1({ S202 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_101_ (
  .in1({ S202, S72 }),
  .out1({ S203 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_102_ (
  .in1({ S203, S229 }),
  .out1({ S204 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_41_ (
  .in1({ S204 }),
  .out1({ CU_selPC_OF })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_102_ (
  .in1({ S230, CU_inst_5 }),
  .out1({ S205 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_103_ (
  .in1({ S205, S77 }),
  .out1({ S206 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_42_ (
  .in1({ S206 }),
  .out1({ CU_zeroAC })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_103_ (
  .in1({ S97, S222 }),
  .out1({ CU_ldIN })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_104_ (
  .in1({ S204, S195 }),
  .out1({ CU_ldOF })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_1_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ CU_nstate_0 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_pstate_0 }),
  .Si({ S3100 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_2_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ CU_nstate_1 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_pstate_1 }),
  .Si({ S3101 }),
  .global_reset({ 1'b0 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_43_ (
  .in1({ DP_SR_V_dout }),
  .out1({ S239 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_44_ (
  .in1({ DP_SR_C_dout }),
  .out1({ S240 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_45_ (
  .in1({ DP_SR_N_dout }),
  .out1({ S241 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_46_ (
  .in1({ DP_SR_Z_dout }),
  .out1({ S242 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_104_ (
  .in1({ S241, CU_inst_2 }),
  .out1({ S243 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_105_ (
  .in1({ S241, CU_inst_2 }),
  .out1({ S244 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_106_ (
  .in1({ S244, CU_inst_6 }),
  .out1({ S245 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_105_ (
  .in1({ S245, S243 }),
  .out1({ S246 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_106_ (
  .in1({ S242, CU_inst_3 }),
  .out1({ S247 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_107_ (
  .in1({ S242, CU_inst_3 }),
  .out1({ S248 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_108_ (
  .in1({ S248, CU_inst_7 }),
  .out1({ S249 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_107_ (
  .in1({ S249, S247 }),
  .out1({ S250 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_108_ (
  .in1({ S250, S246 }),
  .out1({ S251 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_109_ (
  .in1({ S239, CU_inst_0 }),
  .out1({ S252 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_109_ (
  .in1({ S239, CU_inst_0 }),
  .out1({ S253 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_110_ (
  .in1({ S253, CU_inst_4 }),
  .out1({ S254 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_110_ (
  .in1({ S254, S252 }),
  .out1({ S255 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_111_ (
  .in1({ S240, CU_inst_1 }),
  .out1({ S256 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_111_ (
  .in1({ S240, CU_inst_1 }),
  .out1({ S257 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_112_ (
  .in1({ S257, CU_inst_5 }),
  .out1({ S258 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_112_ (
  .in1({ S258, S256 }),
  .out1({ S259 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_113_ (
  .in1({ S259, S255 }),
  .out1({ S260 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_113_ (
  .in1({ S260, S251 }),
  .out1({ CU_enSKP })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_47_ (
  .in1({ CU_ldAC }),
  .out1({ S278 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_114_ (
  .in1({ CU_ldAC, CU_zeroAC }),
  .out1({ S279 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_114_ (
  .in1({ S279, DP_AC_dout_0 }),
  .out1({ S280 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_115_ (
  .in1({ S278, CU_zeroAC }),
  .out1({ S281 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_115_ (
  .in1({ S281, DP_AC_din_0 }),
  .out1({ S282 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_116_ (
  .in1({ S282, S280 }),
  .out1({ S261 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_117_ (
  .in1({ S279, DP_AC_dout_1 }),
  .out1({ S283 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_118_ (
  .in1({ S281, DP_AC_din_1 }),
  .out1({ S284 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_119_ (
  .in1({ S284, S283 }),
  .out1({ S262 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_120_ (
  .in1({ S279, DP_AC_dout_2 }),
  .out1({ S285 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_121_ (
  .in1({ S281, DP_AC_din_2 }),
  .out1({ S286 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_122_ (
  .in1({ S286, S285 }),
  .out1({ S263 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_123_ (
  .in1({ S279, DP_AC_dout_3 }),
  .out1({ S287 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_124_ (
  .in1({ S281, DP_AC_din_3 }),
  .out1({ S288 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_125_ (
  .in1({ S288, S287 }),
  .out1({ S264 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_126_ (
  .in1({ S279, DP_AC_dout_4 }),
  .out1({ S289 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_127_ (
  .in1({ S281, DP_AC_din_4 }),
  .out1({ S290 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_128_ (
  .in1({ S290, S289 }),
  .out1({ S265 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_129_ (
  .in1({ S279, DP_AC_dout_5 }),
  .out1({ S291 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_130_ (
  .in1({ S281, DP_AC_din_5 }),
  .out1({ S292 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_131_ (
  .in1({ S292, S291 }),
  .out1({ S266 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_132_ (
  .in1({ S279, DP_AC_dout_6 }),
  .out1({ S293 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_133_ (
  .in1({ S281, DP_AC_din_6 }),
  .out1({ S294 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_134_ (
  .in1({ S294, S293 }),
  .out1({ S267 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_135_ (
  .in1({ S279, DP_AC_dout_7 }),
  .out1({ S295 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_136_ (
  .in1({ S281, DP_AC_din_7 }),
  .out1({ S296 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_137_ (
  .in1({ S296, S295 }),
  .out1({ S268 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_138_ (
  .in1({ S279, DP_AC_dout_8 }),
  .out1({ S297 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_139_ (
  .in1({ S281, DP_AC_din_8 }),
  .out1({ S298 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_140_ (
  .in1({ S298, S297 }),
  .out1({ S269 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_141_ (
  .in1({ S279, DP_AC_dout_9 }),
  .out1({ S299 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_142_ (
  .in1({ S281, DP_AC_din_9 }),
  .out1({ S300 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_143_ (
  .in1({ S300, S299 }),
  .out1({ S270 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_144_ (
  .in1({ S279, DP_AC_dout_10 }),
  .out1({ S301 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_145_ (
  .in1({ S281, DP_AC_din_10 }),
  .out1({ S302 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_146_ (
  .in1({ S302, S301 }),
  .out1({ S271 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_147_ (
  .in1({ S279, DP_AC_dout_11 }),
  .out1({ S303 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_148_ (
  .in1({ S281, DP_AC_din_11 }),
  .out1({ S304 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_149_ (
  .in1({ S304, S303 }),
  .out1({ S272 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_150_ (
  .in1({ S279, DP_AC_dout_12 }),
  .out1({ S305 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_151_ (
  .in1({ S281, DP_AC_din_12 }),
  .out1({ S306 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_152_ (
  .in1({ S306, S305 }),
  .out1({ S273 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_153_ (
  .in1({ S279, DP_AC_dout_13 }),
  .out1({ S307 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_154_ (
  .in1({ S281, DP_AC_din_13 }),
  .out1({ S308 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_155_ (
  .in1({ S308, S307 }),
  .out1({ S274 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_156_ (
  .in1({ S279, DP_AC_dout_14 }),
  .out1({ S309 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_157_ (
  .in1({ S281, DP_AC_din_14 }),
  .out1({ S310 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_158_ (
  .in1({ S310, S309 }),
  .out1({ S275 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_159_ (
  .in1({ S279, DP_AC_dout_15 }),
  .out1({ S311 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_160_ (
  .in1({ S281, DP_AC_din_15 }),
  .out1({ S277 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_161_ (
  .in1({ S277, S311 }),
  .out1({ S276 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_3_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S261 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_dout_0 }),
  .Si({ S3042 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_4_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S262 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_dout_1 }),
  .Si({ S3041 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_5_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S263 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_dout_2 }),
  .Si({ S3040 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_6_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S264 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_dout_3 }),
  .Si({ S3039 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_7_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S265 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_dout_4 }),
  .Si({ S3038 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_8_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S266 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_dout_5 }),
  .Si({ S3037 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_9_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S267 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_dout_6 }),
  .Si({ S3036 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_10_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S268 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_dout_7 }),
  .Si({ S3035 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_11_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S269 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_dout_8 }),
  .Si({ S3034 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_12_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S270 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_dout_9 }),
  .Si({ S3033 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_13_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S271 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_dout_10 }),
  .Si({ S3032 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_14_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S272 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_dout_11 }),
  .Si({ S3031 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_15_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S273 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_dout_12 }),
  .Si({ S3030 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_16_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S274 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_dout_13 }),
  .Si({ S3029 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_17_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S275 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_dout_14 }),
  .Si({ S3028 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_18_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S276 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_dout_15 }),
  .Si({ S3091 }),
  .global_reset({ 1'b0 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_48_ (
  .in1({ DP_AC_dout_0 }),
  .out1({ S773 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_49_ (
  .in1({ DP_ARU1_in1_0 }),
  .out1({ S784 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_50_ (
  .in1({ CU_ADD }),
  .out1({ S795 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_51_ (
  .in1({ DP_AC_dout_1 }),
  .out1({ S806 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_52_ (
  .in1({ DP_ARU1_in1_1 }),
  .out1({ S817 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_53_ (
  .in1({ DP_AC_dout_2 }),
  .out1({ S828 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_54_ (
  .in1({ DP_ARU1_in1_2 }),
  .out1({ S839 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_55_ (
  .in1({ DP_AC_dout_3 }),
  .out1({ S850 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_56_ (
  .in1({ DP_ARU1_in1_3 }),
  .out1({ S861 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_57_ (
  .in1({ DP_AC_dout_4 }),
  .out1({ S871 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_58_ (
  .in1({ DP_ARU1_in1_4 }),
  .out1({ S882 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_59_ (
  .in1({ DP_AC_dout_5 }),
  .out1({ S893 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_60_ (
  .in1({ DP_ARU1_in1_5 }),
  .out1({ S904 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_61_ (
  .in1({ DP_AC_dout_6 }),
  .out1({ S915 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_62_ (
  .in1({ DP_ARU1_in1_6 }),
  .out1({ S926 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_63_ (
  .in1({ DP_AC_dout_7 }),
  .out1({ S937 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_64_ (
  .in1({ DP_ARU1_in1_7 }),
  .out1({ S948 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_65_ (
  .in1({ DP_AC_dout_8 }),
  .out1({ S959 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_66_ (
  .in1({ DP_ARU1_in1_8 }),
  .out1({ S969 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_67_ (
  .in1({ DP_AC_dout_9 }),
  .out1({ S980 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_68_ (
  .in1({ DP_ARU1_in1_9 }),
  .out1({ S991 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_69_ (
  .in1({ DP_AC_dout_11 }),
  .out1({ S1002 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_70_ (
  .in1({ DP_ARU1_in1_11 }),
  .out1({ S1013 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_71_ (
  .in1({ DP_AC_dout_14 }),
  .out1({ S1024 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_72_ (
  .in1({ DP_ARU1_in1_14 }),
  .out1({ S1035 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_73_ (
  .in1({ DP_AC_dout_15 }),
  .out1({ S1046 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_74_ (
  .in1({ DP_ARU1_in1_15 }),
  .out1({ S1056 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_116_ (
  .in1({ DP_ARU1_in1_0, DP_AC_dout_0 }),
  .out1({ S1067 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_117_ (
  .in1({ S784, S773 }),
  .out1({ S1078 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_162_ (
  .in1({ DP_ARU1_in1_0, DP_AC_dout_0 }),
  .out1({ S1089 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_118_ (
  .in1({ S1089, S795 }),
  .out1({ S1100 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_119_ (
  .in1({ S1067, S795 }),
  .out1({ S1111 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_120_ (
  .in1({ S1111, S1078 }),
  .out1({ S1122 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_121_ (
  .in1({ S1122, S1100 }),
  .out1({ DP_ARU1_out_0 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_122_ (
  .in1({ S817, S806 }),
  .out1({ S1142 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_163_ (
  .in1({ DP_ARU1_in1_1, DP_AC_dout_1 }),
  .out1({ S1153 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_123_ (
  .in1({ DP_ARU1_in1_1, DP_AC_dout_1 }),
  .out1({ S1164 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_124_ (
  .in1({ S1164, S1142 }),
  .out1({ S1175 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_75_ (
  .in1({ S1175 }),
  .out1({ S1186 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_125_ (
  .in1({ S1186, S1089 }),
  .out1({ S1196 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_164_ (
  .in1({ S1175, S1078 }),
  .out1({ S1207 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_126_ (
  .in1({ S1175, S1078 }),
  .out1({ S1218 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_127_ (
  .in1({ S817, S773 }),
  .out1({ S1229 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_128_ (
  .in1({ S806, S784 }),
  .out1({ S1239 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_129_ (
  .in1({ S1153, S1089 }),
  .out1({ S1250 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_165_ (
  .in1({ S1142, S1078 }),
  .out1({ S1261 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_130_ (
  .in1({ S1239, S1229 }),
  .out1({ S1271 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_131_ (
  .in1({ S1271, S1250 }),
  .out1({ S322 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_166_ (
  .in1({ S322, S795 }),
  .out1({ S332 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_132_ (
  .in1({ S1218, S795 }),
  .out1({ S341 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_167_ (
  .in1({ S341, S1207 }),
  .out1({ S343 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_168_ (
  .in1({ S343, S332 }),
  .out1({ DP_ARU1_out_1 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_133_ (
  .in1({ S1196, S1142 }),
  .out1({ S344 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_169_ (
  .in1({ S1207, S1153 }),
  .out1({ S345 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_134_ (
  .in1({ S839, S828 }),
  .out1({ S346 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_170_ (
  .in1({ DP_ARU1_in1_2, DP_AC_dout_2 }),
  .out1({ S347 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_135_ (
  .in1({ DP_ARU1_in1_2, DP_AC_dout_2 }),
  .out1({ S348 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_76_ (
  .in1({ S348 }),
  .out1({ S349 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_136_ (
  .in1({ S348, S346 }),
  .out1({ S350 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_171_ (
  .in1({ S349, S347 }),
  .out1({ S351 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_172_ (
  .in1({ S351, S344 }),
  .out1({ S352 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_173_ (
  .in1({ S350, S345 }),
  .out1({ S353 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_174_ (
  .in1({ S353, S352 }),
  .out1({ S354 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_175_ (
  .in1({ S354, CU_ADD }),
  .out1({ S355 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_176_ (
  .in1({ DP_ARU1_in1_2, DP_AC_dout_0 }),
  .out1({ S356 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_177_ (
  .in1({ DP_AC_dout_2, DP_ARU1_in1_0 }),
  .out1({ S357 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_178_ (
  .in1({ DP_AC_dout_2, DP_ARU1_in1_1 }),
  .out1({ S358 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_77_ (
  .in1({ S358 }),
  .out1({ S359 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_137_ (
  .in1({ S357, S1153 }),
  .out1({ S360 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_78_ (
  .in1({ S360 }),
  .out1({ S361 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_179_ (
  .in1({ S357, S1153 }),
  .out1({ S362 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_180_ (
  .in1({ S362, S361 }),
  .out1({ S363 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_138_ (
  .in1({ S363, S356 }),
  .out1({ S364 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_79_ (
  .in1({ S364 }),
  .out1({ S365 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_181_ (
  .in1({ S363, S356 }),
  .out1({ S366 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_80_ (
  .in1({ S366 }),
  .out1({ S367 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_139_ (
  .in1({ S367, S364 }),
  .out1({ S368 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_182_ (
  .in1({ S366, S365 }),
  .out1({ S369 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_140_ (
  .in1({ S368, S1250 }),
  .out1({ S370 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_141_ (
  .in1({ S369, S1261 }),
  .out1({ S371 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_142_ (
  .in1({ S371, S370 }),
  .out1({ S372 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_143_ (
  .in1({ S372, CU_ADD }),
  .out1({ S373 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_81_ (
  .in1({ S373 }),
  .out1({ S374 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_183_ (
  .in1({ S374, S355 }),
  .out1({ S375 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_82_ (
  .in1({ S375 }),
  .out1({ DP_ARU1_out_2 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_184_ (
  .in1({ S353, S347 }),
  .out1({ S376 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_144_ (
  .in1({ S861, S850 }),
  .out1({ S377 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_185_ (
  .in1({ DP_ARU1_in1_3, DP_AC_dout_3 }),
  .out1({ S378 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_145_ (
  .in1({ DP_ARU1_in1_3, DP_AC_dout_3 }),
  .out1({ S379 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_146_ (
  .in1({ S379, S377 }),
  .out1({ S380 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_186_ (
  .in1({ S380, S376 }),
  .out1({ S381 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_83_ (
  .in1({ S381 }),
  .out1({ S382 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_147_ (
  .in1({ S380, S376 }),
  .out1({ S383 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_148_ (
  .in1({ S383, S382 }),
  .out1({ S384 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_187_ (
  .in1({ S384, CU_ADD }),
  .out1({ S385 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_188_ (
  .in1({ DP_ARU1_in1_3, DP_AC_dout_0 }),
  .out1({ S386 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_84_ (
  .in1({ S386 }),
  .out1({ S387 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_149_ (
  .in1({ S364, S360 }),
  .out1({ S388 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_189_ (
  .in1({ DP_ARU1_in1_2, DP_AC_dout_1 }),
  .out1({ S389 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_85_ (
  .in1({ S389 }),
  .out1({ S390 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_190_ (
  .in1({ DP_AC_dout_3, DP_ARU1_in1_0 }),
  .out1({ S391 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_86_ (
  .in1({ S391 }),
  .out1({ S392 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_191_ (
  .in1({ DP_AC_dout_3, DP_ARU1_in1_1 }),
  .out1({ S393 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_150_ (
  .in1({ S391, S358 }),
  .out1({ S394 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_192_ (
  .in1({ S392, S359 }),
  .out1({ S395 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_193_ (
  .in1({ S391, S358 }),
  .out1({ S396 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_87_ (
  .in1({ S396 }),
  .out1({ S397 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_151_ (
  .in1({ S397, S394 }),
  .out1({ S398 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_194_ (
  .in1({ S396, S395 }),
  .out1({ S399 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_152_ (
  .in1({ S399, S389 }),
  .out1({ S400 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_195_ (
  .in1({ S398, S390 }),
  .out1({ S401 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_196_ (
  .in1({ S399, S389 }),
  .out1({ S402 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_197_ (
  .in1({ S402, S401 }),
  .out1({ S403 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_153_ (
  .in1({ S403, S388 }),
  .out1({ S404 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_88_ (
  .in1({ S404 }),
  .out1({ S405 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_198_ (
  .in1({ S403, S388 }),
  .out1({ S406 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_199_ (
  .in1({ S406, S405 }),
  .out1({ S407 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_154_ (
  .in1({ S407, S386 }),
  .out1({ S408 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_200_ (
  .in1({ S407, S386 }),
  .out1({ S409 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_89_ (
  .in1({ S409 }),
  .out1({ S410 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_155_ (
  .in1({ S410, S408 }),
  .out1({ S411 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_201_ (
  .in1({ S411, S371 }),
  .out1({ S412 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_156_ (
  .in1({ S411, S371 }),
  .out1({ S413 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_157_ (
  .in1({ S413, CU_ADD }),
  .out1({ S414 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_202_ (
  .in1({ S414, S412 }),
  .out1({ S415 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_203_ (
  .in1({ S415, S385 }),
  .out1({ DP_ARU1_out_3 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_158_ (
  .in1({ S882, S871 }),
  .out1({ S416 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_204_ (
  .in1({ DP_ARU1_in1_4, DP_AC_dout_4 }),
  .out1({ S417 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_159_ (
  .in1({ DP_ARU1_in1_4, DP_AC_dout_4 }),
  .out1({ S418 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_160_ (
  .in1({ S418, S416 }),
  .out1({ S419 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_161_ (
  .in1({ S377, S376 }),
  .out1({ S420 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_162_ (
  .in1({ S420, S379 }),
  .out1({ S421 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_205_ (
  .in1({ S421, S419 }),
  .out1({ S422 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_90_ (
  .in1({ S422 }),
  .out1({ S423 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_163_ (
  .in1({ S421, S419 }),
  .out1({ S424 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_164_ (
  .in1({ S424, S423 }),
  .out1({ S425 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_165_ (
  .in1({ S408, S404 }),
  .out1({ S426 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_206_ (
  .in1({ DP_ARU1_in1_4, DP_AC_dout_0 }),
  .out1({ S427 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_207_ (
  .in1({ DP_ARU1_in1_3, DP_AC_dout_1 }),
  .out1({ S428 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_208_ (
  .in1({ DP_ARU1_in1_4, DP_AC_dout_1 }),
  .out1({ S429 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_91_ (
  .in1({ S429 }),
  .out1({ S430 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_166_ (
  .in1({ S429, S386 }),
  .out1({ S431 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_209_ (
  .in1({ S430, S387 }),
  .out1({ S432 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_210_ (
  .in1({ S428, S427 }),
  .out1({ S433 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_211_ (
  .in1({ S433, S432 }),
  .out1({ S434 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_92_ (
  .in1({ S434 }),
  .out1({ S435 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_167_ (
  .in1({ S400, S394 }),
  .out1({ S436 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_212_ (
  .in1({ S401, S395 }),
  .out1({ S437 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_213_ (
  .in1({ DP_AC_dout_4, DP_ARU1_in1_0 }),
  .out1({ S438 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_214_ (
  .in1({ S438, S393 }),
  .out1({ S439 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_93_ (
  .in1({ S439 }),
  .out1({ S440 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_215_ (
  .in1({ DP_AC_dout_4, DP_ARU1_in1_1 }),
  .out1({ S441 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_94_ (
  .in1({ S441 }),
  .out1({ S442 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_168_ (
  .in1({ S438, S393 }),
  .out1({ S443 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_216_ (
  .in1({ S442, S392 }),
  .out1({ S444 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_169_ (
  .in1({ S443, S440 }),
  .out1({ S445 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_217_ (
  .in1({ S444, S439 }),
  .out1({ S446 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_170_ (
  .in1({ S446, S347 }),
  .out1({ S447 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_218_ (
  .in1({ S445, S346 }),
  .out1({ S448 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_171_ (
  .in1({ S445, S346 }),
  .out1({ S449 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_219_ (
  .in1({ S446, S347 }),
  .out1({ S450 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_172_ (
  .in1({ S449, S447 }),
  .out1({ S451 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_220_ (
  .in1({ S450, S448 }),
  .out1({ S452 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_173_ (
  .in1({ S452, S436 }),
  .out1({ S453 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_221_ (
  .in1({ S451, S437 }),
  .out1({ S454 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_174_ (
  .in1({ S451, S437 }),
  .out1({ S455 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_222_ (
  .in1({ S452, S436 }),
  .out1({ S456 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_175_ (
  .in1({ S455, S453 }),
  .out1({ S457 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_223_ (
  .in1({ S456, S454 }),
  .out1({ S458 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_176_ (
  .in1({ S458, S434 }),
  .out1({ S459 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_224_ (
  .in1({ S457, S435 }),
  .out1({ S460 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_225_ (
  .in1({ S458, S434 }),
  .out1({ S461 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_226_ (
  .in1({ S461, S460 }),
  .out1({ S462 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_227_ (
  .in1({ S462, S426 }),
  .out1({ S463 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_177_ (
  .in1({ S462, S426 }),
  .out1({ S464 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_95_ (
  .in1({ S464 }),
  .out1({ S465 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_228_ (
  .in1({ S465, S463 }),
  .out1({ S466 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_229_ (
  .in1({ S466, S412 }),
  .out1({ S467 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_178_ (
  .in1({ S466, S412 }),
  .out1({ S468 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_96_ (
  .in1({ S468 }),
  .out1({ S469 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_179_ (
  .in1({ S468, CU_ADD }),
  .out1({ S470 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_230_ (
  .in1({ S470, S467 }),
  .out1({ S471 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_231_ (
  .in1({ S425, CU_ADD }),
  .out1({ S472 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_232_ (
  .in1({ S472, S471 }),
  .out1({ DP_ARU1_out_4 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_97_ (
  .in1({ DP_ARU1_out_4 }),
  .out1({ S473 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_233_ (
  .in1({ S422, S417 }),
  .out1({ S474 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_180_ (
  .in1({ S904, S893 }),
  .out1({ S475 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_234_ (
  .in1({ DP_ARU1_in1_5, DP_AC_dout_5 }),
  .out1({ S476 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_181_ (
  .in1({ DP_ARU1_in1_5, DP_AC_dout_5 }),
  .out1({ S477 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_182_ (
  .in1({ S477, S475 }),
  .out1({ S478 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_183_ (
  .in1({ S478, S474 }),
  .out1({ S479 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_235_ (
  .in1({ S478, S474 }),
  .out1({ S480 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_98_ (
  .in1({ S480 }),
  .out1({ S481 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_184_ (
  .in1({ S481, S479 }),
  .out1({ S482 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_185_ (
  .in1({ S482, S795 }),
  .out1({ S483 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_186_ (
  .in1({ S459, S453 }),
  .out1({ S484 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_236_ (
  .in1({ S460, S454 }),
  .out1({ S485 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_237_ (
  .in1({ DP_ARU1_in1_5, DP_AC_dout_0 }),
  .out1({ S486 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_238_ (
  .in1({ DP_ARU1_in1_3, DP_AC_dout_2 }),
  .out1({ S487 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_239_ (
  .in1({ DP_ARU1_in1_4, DP_AC_dout_2 }),
  .out1({ S488 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_187_ (
  .in1({ S487, S429 }),
  .out1({ S489 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_99_ (
  .in1({ S489 }),
  .out1({ S490 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_240_ (
  .in1({ S487, S429 }),
  .out1({ S491 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_241_ (
  .in1({ S491, S490 }),
  .out1({ S492 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_188_ (
  .in1({ S492, S486 }),
  .out1({ S493 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_100_ (
  .in1({ S493 }),
  .out1({ S494 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_242_ (
  .in1({ S492, S486 }),
  .out1({ S495 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_101_ (
  .in1({ S495 }),
  .out1({ S496 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_189_ (
  .in1({ S496, S493 }),
  .out1({ S497 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_243_ (
  .in1({ S495, S494 }),
  .out1({ S498 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_190_ (
  .in1({ S447, S443 }),
  .out1({ S499 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_244_ (
  .in1({ S448, S444 }),
  .out1({ S500 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_245_ (
  .in1({ DP_AC_dout_3, DP_ARU1_in1_2 }),
  .out1({ S501 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_102_ (
  .in1({ S501 }),
  .out1({ S502 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_246_ (
  .in1({ DP_AC_dout_5, DP_ARU1_in1_0 }),
  .out1({ S503 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_103_ (
  .in1({ S503 }),
  .out1({ S504 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_247_ (
  .in1({ DP_AC_dout_5, DP_ARU1_in1_1 }),
  .out1({ S505 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_191_ (
  .in1({ S503, S441 }),
  .out1({ S506 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_248_ (
  .in1({ S504, S442 }),
  .out1({ S507 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_249_ (
  .in1({ S503, S441 }),
  .out1({ S508 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_104_ (
  .in1({ S508 }),
  .out1({ S509 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_192_ (
  .in1({ S509, S506 }),
  .out1({ S510 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_250_ (
  .in1({ S508, S507 }),
  .out1({ S511 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_193_ (
  .in1({ S511, S501 }),
  .out1({ S512 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_251_ (
  .in1({ S510, S502 }),
  .out1({ S513 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_194_ (
  .in1({ S510, S502 }),
  .out1({ S514 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_252_ (
  .in1({ S511, S501 }),
  .out1({ S515 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_195_ (
  .in1({ S514, S512 }),
  .out1({ S516 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_253_ (
  .in1({ S515, S513 }),
  .out1({ S517 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_196_ (
  .in1({ S517, S499 }),
  .out1({ S518 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_254_ (
  .in1({ S516, S500 }),
  .out1({ S519 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_197_ (
  .in1({ S516, S500 }),
  .out1({ S520 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_255_ (
  .in1({ S517, S499 }),
  .out1({ S521 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_198_ (
  .in1({ S520, S518 }),
  .out1({ S522 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_256_ (
  .in1({ S521, S519 }),
  .out1({ S523 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_199_ (
  .in1({ S523, S498 }),
  .out1({ S524 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_257_ (
  .in1({ S522, S497 }),
  .out1({ S525 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_200_ (
  .in1({ S522, S497 }),
  .out1({ S526 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_258_ (
  .in1({ S523, S498 }),
  .out1({ S527 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_201_ (
  .in1({ S526, S524 }),
  .out1({ S528 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_259_ (
  .in1({ S527, S525 }),
  .out1({ S529 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_202_ (
  .in1({ S529, S484 }),
  .out1({ S530 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_260_ (
  .in1({ S528, S485 }),
  .out1({ S531 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_203_ (
  .in1({ S528, S485 }),
  .out1({ S532 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_261_ (
  .in1({ S529, S484 }),
  .out1({ S533 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_204_ (
  .in1({ S532, S530 }),
  .out1({ S534 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_262_ (
  .in1({ S533, S531 }),
  .out1({ S535 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_205_ (
  .in1({ S535, S432 }),
  .out1({ S536 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_263_ (
  .in1({ S534, S431 }),
  .out1({ S537 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_206_ (
  .in1({ S534, S431 }),
  .out1({ S538 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_264_ (
  .in1({ S535, S432 }),
  .out1({ S539 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_207_ (
  .in1({ S538, S536 }),
  .out1({ S540 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_265_ (
  .in1({ S539, S537 }),
  .out1({ S541 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_208_ (
  .in1({ S541, S465 }),
  .out1({ S542 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_266_ (
  .in1({ S540, S464 }),
  .out1({ S543 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_209_ (
  .in1({ S540, S464 }),
  .out1({ S544 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_210_ (
  .in1({ S544, S542 }),
  .out1({ S545 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_105_ (
  .in1({ S545 }),
  .out1({ S546 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_211_ (
  .in1({ S545, S468 }),
  .out1({ S547 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_212_ (
  .in1({ S546, S469 }),
  .out1({ S548 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_267_ (
  .in1({ S545, S468 }),
  .out1({ S549 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_213_ (
  .in1({ S548, S547 }),
  .out1({ S550 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_214_ (
  .in1({ S550, CU_ADD }),
  .out1({ S551 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_215_ (
  .in1({ S551, S483 }),
  .out1({ DP_ARU1_out_5 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_268_ (
  .in1({ S480, S476 }),
  .out1({ S552 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_216_ (
  .in1({ S926, S915 }),
  .out1({ S553 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_269_ (
  .in1({ DP_ARU1_in1_6, DP_AC_dout_6 }),
  .out1({ S554 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_217_ (
  .in1({ DP_ARU1_in1_6, DP_AC_dout_6 }),
  .out1({ S555 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_218_ (
  .in1({ S555, S553 }),
  .out1({ S556 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_219_ (
  .in1({ S556, S552 }),
  .out1({ S557 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_270_ (
  .in1({ S556, S552 }),
  .out1({ S558 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_220_ (
  .in1({ S536, S530 }),
  .out1({ S559 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_271_ (
  .in1({ S537, S531 }),
  .out1({ S560 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_272_ (
  .in1({ DP_ARU1_in1_6, DP_AC_dout_0 }),
  .out1({ S561 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_106_ (
  .in1({ S561 }),
  .out1({ S562 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_221_ (
  .in1({ S493, S489 }),
  .out1({ S563 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_107_ (
  .in1({ S563 }),
  .out1({ S564 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_273_ (
  .in1({ S563, S561 }),
  .out1({ S565 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_108_ (
  .in1({ S565 }),
  .out1({ S566 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_222_ (
  .in1({ S563, S561 }),
  .out1({ S567 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_274_ (
  .in1({ S564, S562 }),
  .out1({ S568 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_223_ (
  .in1({ S567, S566 }),
  .out1({ S569 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_275_ (
  .in1({ S568, S565 }),
  .out1({ S570 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_224_ (
  .in1({ S524, S518 }),
  .out1({ S571 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_276_ (
  .in1({ S525, S519 }),
  .out1({ S572 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_277_ (
  .in1({ DP_ARU1_in1_5, DP_AC_dout_1 }),
  .out1({ S573 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_278_ (
  .in1({ DP_ARU1_in1_4, DP_AC_dout_3 }),
  .out1({ S574 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_225_ (
  .in1({ S488, S378 }),
  .out1({ S575 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_109_ (
  .in1({ S575 }),
  .out1({ S576 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_279_ (
  .in1({ S488, S378 }),
  .out1({ S577 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_280_ (
  .in1({ S577, S576 }),
  .out1({ S578 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_226_ (
  .in1({ S578, S573 }),
  .out1({ S579 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_110_ (
  .in1({ S579 }),
  .out1({ S580 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_281_ (
  .in1({ S578, S573 }),
  .out1({ S581 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_111_ (
  .in1({ S581 }),
  .out1({ S582 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_227_ (
  .in1({ S582, S579 }),
  .out1({ S583 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_282_ (
  .in1({ S581, S580 }),
  .out1({ S584 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_228_ (
  .in1({ S512, S506 }),
  .out1({ S585 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_283_ (
  .in1({ S513, S507 }),
  .out1({ S586 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_284_ (
  .in1({ DP_AC_dout_4, DP_ARU1_in1_2 }),
  .out1({ S587 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_112_ (
  .in1({ S587 }),
  .out1({ S588 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_285_ (
  .in1({ DP_AC_dout_6, DP_ARU1_in1_0 }),
  .out1({ S589 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_229_ (
  .in1({ S915, S817 }),
  .out1({ S590 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_286_ (
  .in1({ DP_AC_dout_6, DP_ARU1_in1_1 }),
  .out1({ S591 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_230_ (
  .in1({ S591, S503 }),
  .out1({ S592 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_287_ (
  .in1({ S590, S504 }),
  .out1({ S593 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_288_ (
  .in1({ S589, S505 }),
  .out1({ S594 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_113_ (
  .in1({ S594 }),
  .out1({ S595 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_231_ (
  .in1({ S595, S592 }),
  .out1({ S596 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_289_ (
  .in1({ S594, S593 }),
  .out1({ S597 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_232_ (
  .in1({ S597, S587 }),
  .out1({ S598 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_290_ (
  .in1({ S596, S588 }),
  .out1({ S599 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_233_ (
  .in1({ S596, S588 }),
  .out1({ S600 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_291_ (
  .in1({ S597, S587 }),
  .out1({ S601 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_234_ (
  .in1({ S600, S598 }),
  .out1({ S602 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_292_ (
  .in1({ S601, S599 }),
  .out1({ S603 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_235_ (
  .in1({ S603, S585 }),
  .out1({ S604 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_293_ (
  .in1({ S602, S586 }),
  .out1({ S605 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_236_ (
  .in1({ S602, S586 }),
  .out1({ S606 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_294_ (
  .in1({ S603, S585 }),
  .out1({ S607 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_237_ (
  .in1({ S606, S604 }),
  .out1({ S608 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_295_ (
  .in1({ S607, S605 }),
  .out1({ S609 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_238_ (
  .in1({ S609, S584 }),
  .out1({ S610 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_296_ (
  .in1({ S608, S583 }),
  .out1({ S611 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_239_ (
  .in1({ S608, S583 }),
  .out1({ S612 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_297_ (
  .in1({ S609, S584 }),
  .out1({ S613 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_240_ (
  .in1({ S612, S610 }),
  .out1({ S614 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_298_ (
  .in1({ S613, S611 }),
  .out1({ S615 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_241_ (
  .in1({ S615, S571 }),
  .out1({ S616 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_299_ (
  .in1({ S614, S572 }),
  .out1({ S617 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_242_ (
  .in1({ S614, S572 }),
  .out1({ S618 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_300_ (
  .in1({ S615, S571 }),
  .out1({ S619 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_243_ (
  .in1({ S618, S616 }),
  .out1({ S620 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_301_ (
  .in1({ S619, S617 }),
  .out1({ S621 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_244_ (
  .in1({ S621, S570 }),
  .out1({ S622 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_302_ (
  .in1({ S620, S569 }),
  .out1({ S623 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_245_ (
  .in1({ S620, S569 }),
  .out1({ S624 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_303_ (
  .in1({ S621, S570 }),
  .out1({ S625 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_246_ (
  .in1({ S624, S622 }),
  .out1({ S626 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_304_ (
  .in1({ S625, S623 }),
  .out1({ S627 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_247_ (
  .in1({ S627, S559 }),
  .out1({ S628 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_305_ (
  .in1({ S626, S560 }),
  .out1({ S629 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_248_ (
  .in1({ S626, S560 }),
  .out1({ S630 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_306_ (
  .in1({ S627, S559 }),
  .out1({ S631 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_249_ (
  .in1({ S630, S628 }),
  .out1({ S632 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_307_ (
  .in1({ S631, S629 }),
  .out1({ S633 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_250_ (
  .in1({ S632, S542 }),
  .out1({ S634 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_308_ (
  .in1({ S633, S543 }),
  .out1({ S635 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_251_ (
  .in1({ S633, S543 }),
  .out1({ S636 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_309_ (
  .in1({ S632, S542 }),
  .out1({ S637 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_252_ (
  .in1({ S636, S634 }),
  .out1({ S638 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_310_ (
  .in1({ S637, S635 }),
  .out1({ S639 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_253_ (
  .in1({ S638, S548 }),
  .out1({ S640 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_114_ (
  .in1({ S640 }),
  .out1({ S641 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_254_ (
  .in1({ S639, S549 }),
  .out1({ S642 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_311_ (
  .in1({ S638, S548 }),
  .out1({ S643 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_312_ (
  .in1({ S643, S641 }),
  .out1({ S644 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_255_ (
  .in1({ S557, S795 }),
  .out1({ S645 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_313_ (
  .in1({ S645, S558 }),
  .out1({ S646 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_115_ (
  .in1({ S646 }),
  .out1({ S647 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_256_ (
  .in1({ S644, CU_ADD }),
  .out1({ S648 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_257_ (
  .in1({ S648, S647 }),
  .out1({ S649 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_116_ (
  .in1({ S649 }),
  .out1({ DP_ARU1_out_6 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_314_ (
  .in1({ S558, S554 }),
  .out1({ S650 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_117_ (
  .in1({ S650 }),
  .out1({ S651 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_258_ (
  .in1({ S948, S937 }),
  .out1({ S652 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_315_ (
  .in1({ DP_ARU1_in1_7, DP_AC_dout_7 }),
  .out1({ S653 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_259_ (
  .in1({ DP_ARU1_in1_7, DP_AC_dout_7 }),
  .out1({ S654 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_260_ (
  .in1({ S654, S652 }),
  .out1({ S655 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_261_ (
  .in1({ S655, S651 }),
  .out1({ S656 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_316_ (
  .in1({ S655, S651 }),
  .out1({ S657 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_262_ (
  .in1({ S642, S636 }),
  .out1({ S658 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_317_ (
  .in1({ S643, S637 }),
  .out1({ S659 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_263_ (
  .in1({ S622, S616 }),
  .out1({ S660 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_318_ (
  .in1({ S623, S617 }),
  .out1({ S661 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_319_ (
  .in1({ DP_ARU1_in1_7, DP_AC_dout_0 }),
  .out1({ S662 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_320_ (
  .in1({ DP_ARU1_in1_6, DP_AC_dout_1 }),
  .out1({ S663 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_264_ (
  .in1({ S579, S575 }),
  .out1({ S664 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_265_ (
  .in1({ S664, S663 }),
  .out1({ S665 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_118_ (
  .in1({ S665 }),
  .out1({ S666 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_321_ (
  .in1({ S664, S663 }),
  .out1({ S667 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_322_ (
  .in1({ S667, S666 }),
  .out1({ S668 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_266_ (
  .in1({ S668, S662 }),
  .out1({ S669 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_119_ (
  .in1({ S669 }),
  .out1({ S670 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_323_ (
  .in1({ S668, S662 }),
  .out1({ S671 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_120_ (
  .in1({ S671 }),
  .out1({ S672 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_267_ (
  .in1({ S672, S669 }),
  .out1({ S673 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_324_ (
  .in1({ S671, S670 }),
  .out1({ S674 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_268_ (
  .in1({ S610, S604 }),
  .out1({ S675 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_325_ (
  .in1({ S611, S605 }),
  .out1({ S676 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_326_ (
  .in1({ DP_ARU1_in1_5, DP_AC_dout_2 }),
  .out1({ S677 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_327_ (
  .in1({ DP_AC_dout_4, DP_ARU1_in1_3 }),
  .out1({ S678 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_269_ (
  .in1({ S417, S378 }),
  .out1({ S679 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_121_ (
  .in1({ S679 }),
  .out1({ S680 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_328_ (
  .in1({ S678, S574 }),
  .out1({ S681 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_329_ (
  .in1({ S681, S680 }),
  .out1({ S682 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_270_ (
  .in1({ S682, S677 }),
  .out1({ S683 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_122_ (
  .in1({ S683 }),
  .out1({ S684 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_330_ (
  .in1({ S682, S677 }),
  .out1({ S685 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_123_ (
  .in1({ S685 }),
  .out1({ S686 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_271_ (
  .in1({ S686, S683 }),
  .out1({ S687 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_331_ (
  .in1({ S685, S684 }),
  .out1({ S688 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_272_ (
  .in1({ S598, S592 }),
  .out1({ S689 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_332_ (
  .in1({ S599, S593 }),
  .out1({ S690 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_333_ (
  .in1({ DP_AC_dout_5, DP_ARU1_in1_2 }),
  .out1({ S691 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_124_ (
  .in1({ S691 }),
  .out1({ S692 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_334_ (
  .in1({ DP_AC_dout_7, DP_ARU1_in1_0 }),
  .out1({ S693 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_335_ (
  .in1({ DP_AC_dout_7, DP_ARU1_in1_1 }),
  .out1({ S694 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_273_ (
  .in1({ S694, S589 }),
  .out1({ S695 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_125_ (
  .in1({ S695 }),
  .out1({ S696 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_336_ (
  .in1({ S693, S591 }),
  .out1({ S697 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_126_ (
  .in1({ S697 }),
  .out1({ S698 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_274_ (
  .in1({ S698, S695 }),
  .out1({ S699 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_337_ (
  .in1({ S697, S696 }),
  .out1({ S700 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_275_ (
  .in1({ S700, S691 }),
  .out1({ S701 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_338_ (
  .in1({ S699, S692 }),
  .out1({ S702 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_276_ (
  .in1({ S699, S692 }),
  .out1({ S703 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_339_ (
  .in1({ S700, S691 }),
  .out1({ S704 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_277_ (
  .in1({ S703, S701 }),
  .out1({ S705 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_340_ (
  .in1({ S704, S702 }),
  .out1({ S706 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_278_ (
  .in1({ S706, S689 }),
  .out1({ S707 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_341_ (
  .in1({ S705, S690 }),
  .out1({ S708 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_279_ (
  .in1({ S705, S690 }),
  .out1({ S709 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_342_ (
  .in1({ S706, S689 }),
  .out1({ S710 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_280_ (
  .in1({ S709, S707 }),
  .out1({ S711 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_343_ (
  .in1({ S710, S708 }),
  .out1({ S712 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_281_ (
  .in1({ S712, S688 }),
  .out1({ S713 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_344_ (
  .in1({ S711, S687 }),
  .out1({ S714 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_282_ (
  .in1({ S711, S687 }),
  .out1({ S715 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_345_ (
  .in1({ S712, S688 }),
  .out1({ S716 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_283_ (
  .in1({ S715, S713 }),
  .out1({ S717 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_346_ (
  .in1({ S716, S714 }),
  .out1({ S718 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_284_ (
  .in1({ S718, S675 }),
  .out1({ S719 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_347_ (
  .in1({ S717, S676 }),
  .out1({ S720 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_285_ (
  .in1({ S717, S676 }),
  .out1({ S721 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_348_ (
  .in1({ S718, S675 }),
  .out1({ S722 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_286_ (
  .in1({ S721, S719 }),
  .out1({ S723 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_349_ (
  .in1({ S722, S720 }),
  .out1({ S724 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_287_ (
  .in1({ S724, S674 }),
  .out1({ S725 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_350_ (
  .in1({ S723, S673 }),
  .out1({ S726 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_288_ (
  .in1({ S723, S673 }),
  .out1({ S727 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_351_ (
  .in1({ S724, S674 }),
  .out1({ S728 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_289_ (
  .in1({ S727, S725 }),
  .out1({ S729 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_352_ (
  .in1({ S728, S726 }),
  .out1({ S730 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_290_ (
  .in1({ S730, S660 }),
  .out1({ S731 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_353_ (
  .in1({ S729, S661 }),
  .out1({ S732 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_291_ (
  .in1({ S729, S661 }),
  .out1({ S733 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_354_ (
  .in1({ S730, S660 }),
  .out1({ S734 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_292_ (
  .in1({ S733, S731 }),
  .out1({ S735 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_355_ (
  .in1({ S734, S732 }),
  .out1({ S736 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_293_ (
  .in1({ S736, S568 }),
  .out1({ S737 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_356_ (
  .in1({ S735, S567 }),
  .out1({ S738 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_294_ (
  .in1({ S735, S567 }),
  .out1({ S739 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_357_ (
  .in1({ S736, S568 }),
  .out1({ S740 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_295_ (
  .in1({ S739, S737 }),
  .out1({ S741 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_358_ (
  .in1({ S740, S738 }),
  .out1({ S742 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_296_ (
  .in1({ S741, S628 }),
  .out1({ S743 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_359_ (
  .in1({ S742, S629 }),
  .out1({ S744 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_297_ (
  .in1({ S742, S629 }),
  .out1({ S745 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_360_ (
  .in1({ S741, S628 }),
  .out1({ S746 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_298_ (
  .in1({ S745, S743 }),
  .out1({ S747 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_361_ (
  .in1({ S746, S744 }),
  .out1({ S748 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_299_ (
  .in1({ S748, S658 }),
  .out1({ S749 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_362_ (
  .in1({ S747, S659 }),
  .out1({ S750 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_300_ (
  .in1({ S747, S659 }),
  .out1({ S751 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_301_ (
  .in1({ S751, S749 }),
  .out1({ S752 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_302_ (
  .in1({ S752, CU_ADD }),
  .out1({ S753 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_363_ (
  .in1({ S657, CU_ADD }),
  .out1({ S754 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_303_ (
  .in1({ S754, S656 }),
  .out1({ S755 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_304_ (
  .in1({ S755, S753 }),
  .out1({ DP_ARU1_out_7 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_305_ (
  .in1({ S969, S959 }),
  .out1({ S756 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_364_ (
  .in1({ DP_ARU1_in1_8, DP_AC_dout_8 }),
  .out1({ S757 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_306_ (
  .in1({ DP_ARU1_in1_8, DP_AC_dout_8 }),
  .out1({ S758 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_307_ (
  .in1({ S758, S756 }),
  .out1({ S759 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_127_ (
  .in1({ S759 }),
  .out1({ S760 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_308_ (
  .in1({ S652, S650 }),
  .out1({ S761 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_309_ (
  .in1({ S761, S654 }),
  .out1({ S762 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_128_ (
  .in1({ S762 }),
  .out1({ S763 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_310_ (
  .in1({ S763, S760 }),
  .out1({ S764 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_365_ (
  .in1({ S762, S759 }),
  .out1({ S765 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_311_ (
  .in1({ S762, S759 }),
  .out1({ S766 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_312_ (
  .in1({ S766, S764 }),
  .out1({ S767 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_313_ (
  .in1({ S749, S745 }),
  .out1({ S768 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_366_ (
  .in1({ S750, S746 }),
  .out1({ S769 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_314_ (
  .in1({ S737, S731 }),
  .out1({ S770 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_367_ (
  .in1({ S738, S732 }),
  .out1({ S771 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_315_ (
  .in1({ S669, S665 }),
  .out1({ S772 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_316_ (
  .in1({ S725, S719 }),
  .out1({ S774 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_129_ (
  .in1({ S774 }),
  .out1({ S775 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_368_ (
  .in1({ DP_ARU1_in1_7, DP_AC_dout_1 }),
  .out1({ S776 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_369_ (
  .in1({ DP_ARU1_in1_6, DP_AC_dout_2 }),
  .out1({ S777 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_317_ (
  .in1({ S683, S679 }),
  .out1({ S778 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_370_ (
  .in1({ S778, S777 }),
  .out1({ S779 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_318_ (
  .in1({ S778, S777 }),
  .out1({ S780 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_130_ (
  .in1({ S780 }),
  .out1({ S781 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_371_ (
  .in1({ S781, S779 }),
  .out1({ S782 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_372_ (
  .in1({ S782, S776 }),
  .out1({ S783 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_131_ (
  .in1({ S783 }),
  .out1({ S785 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_319_ (
  .in1({ S782, S776 }),
  .out1({ S786 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_132_ (
  .in1({ S786 }),
  .out1({ S787 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_320_ (
  .in1({ S786, S785 }),
  .out1({ S788 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_373_ (
  .in1({ S787, S783 }),
  .out1({ S789 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_321_ (
  .in1({ S713, S707 }),
  .out1({ S790 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_374_ (
  .in1({ S714, S708 }),
  .out1({ S791 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_375_ (
  .in1({ DP_ARU1_in1_5, DP_AC_dout_3 }),
  .out1({ S792 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_376_ (
  .in1({ DP_AC_dout_5, DP_ARU1_in1_3 }),
  .out1({ S793 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_377_ (
  .in1({ DP_AC_dout_5, DP_ARU1_in1_4 }),
  .out1({ S794 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_322_ (
  .in1({ S793, S417 }),
  .out1({ S796 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_133_ (
  .in1({ S796 }),
  .out1({ S797 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_378_ (
  .in1({ S793, S417 }),
  .out1({ S798 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_379_ (
  .in1({ S798, S797 }),
  .out1({ S799 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_323_ (
  .in1({ S799, S792 }),
  .out1({ S800 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_134_ (
  .in1({ S800 }),
  .out1({ S801 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_380_ (
  .in1({ S799, S792 }),
  .out1({ S802 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_135_ (
  .in1({ S802 }),
  .out1({ S803 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_324_ (
  .in1({ S803, S800 }),
  .out1({ S804 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_381_ (
  .in1({ S802, S801 }),
  .out1({ S805 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_325_ (
  .in1({ S701, S695 }),
  .out1({ S807 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_136_ (
  .in1({ S807 }),
  .out1({ S808 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_382_ (
  .in1({ DP_AC_dout_6, DP_ARU1_in1_2 }),
  .out1({ S809 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_383_ (
  .in1({ S809, S694 }),
  .out1({ S810 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_326_ (
  .in1({ S937, S839 }),
  .out1({ S811 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_384_ (
  .in1({ DP_AC_dout_7, DP_ARU1_in1_2 }),
  .out1({ S812 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_327_ (
  .in1({ S812, S591 }),
  .out1({ S813 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_385_ (
  .in1({ S811, S590 }),
  .out1({ S814 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_386_ (
  .in1({ S814, S810 }),
  .out1({ S815 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_137_ (
  .in1({ S815 }),
  .out1({ S816 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_328_ (
  .in1({ S815, S807 }),
  .out1({ S818 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_387_ (
  .in1({ S816, S808 }),
  .out1({ S819 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_388_ (
  .in1({ S815, S807 }),
  .out1({ S820 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_138_ (
  .in1({ S820 }),
  .out1({ S821 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_329_ (
  .in1({ S821, S818 }),
  .out1({ S822 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_389_ (
  .in1({ S820, S819 }),
  .out1({ S823 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_330_ (
  .in1({ S823, S805 }),
  .out1({ S824 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_390_ (
  .in1({ S822, S804 }),
  .out1({ S825 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_331_ (
  .in1({ S822, S804 }),
  .out1({ S826 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_391_ (
  .in1({ S823, S805 }),
  .out1({ S827 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_332_ (
  .in1({ S826, S824 }),
  .out1({ S829 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_392_ (
  .in1({ S827, S825 }),
  .out1({ S830 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_333_ (
  .in1({ S830, S790 }),
  .out1({ S831 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_393_ (
  .in1({ S829, S791 }),
  .out1({ S832 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_334_ (
  .in1({ S829, S791 }),
  .out1({ S833 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_394_ (
  .in1({ S830, S790 }),
  .out1({ S834 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_335_ (
  .in1({ S833, S831 }),
  .out1({ S835 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_395_ (
  .in1({ S834, S832 }),
  .out1({ S836 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_336_ (
  .in1({ S836, S789 }),
  .out1({ S837 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_396_ (
  .in1({ S835, S788 }),
  .out1({ S838 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_337_ (
  .in1({ S835, S788 }),
  .out1({ S840 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_397_ (
  .in1({ S836, S789 }),
  .out1({ S841 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_338_ (
  .in1({ S840, S837 }),
  .out1({ S842 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_398_ (
  .in1({ S841, S838 }),
  .out1({ S843 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_339_ (
  .in1({ S843, S774 }),
  .out1({ S844 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_399_ (
  .in1({ S842, S775 }),
  .out1({ S845 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_400_ (
  .in1({ S843, S774 }),
  .out1({ S846 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_401_ (
  .in1({ S846, S845 }),
  .out1({ S847 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_340_ (
  .in1({ S847, S772 }),
  .out1({ S848 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_139_ (
  .in1({ S848 }),
  .out1({ S849 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_402_ (
  .in1({ S847, S772 }),
  .out1({ S851 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_140_ (
  .in1({ S851 }),
  .out1({ S852 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_341_ (
  .in1({ S852, S848 }),
  .out1({ S853 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_403_ (
  .in1({ S851, S849 }),
  .out1({ S854 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_342_ (
  .in1({ S853, S771 }),
  .out1({ S855 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_404_ (
  .in1({ S854, S770 }),
  .out1({ S856 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_343_ (
  .in1({ S854, S770 }),
  .out1({ S857 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_405_ (
  .in1({ S853, S771 }),
  .out1({ S858 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_344_ (
  .in1({ S857, S855 }),
  .out1({ S859 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_406_ (
  .in1({ S858, S856 }),
  .out1({ S860 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_407_ (
  .in1({ S860, S768 }),
  .out1({ S862 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_345_ (
  .in1({ S860, S768 }),
  .out1({ S863 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_408_ (
  .in1({ S859, S769 }),
  .out1({ S864 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_409_ (
  .in1({ S864, S862 }),
  .out1({ S865 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_346_ (
  .in1({ S865, CU_ADD }),
  .out1({ S866 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_410_ (
  .in1({ S767, CU_ADD }),
  .out1({ S867 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_141_ (
  .in1({ S867 }),
  .out1({ S868 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_347_ (
  .in1({ S868, S866 }),
  .out1({ S869 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_142_ (
  .in1({ S869 }),
  .out1({ DP_ARU1_out_8 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_348_ (
  .in1({ S764, S756 }),
  .out1({ S870 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_411_ (
  .in1({ S765, S757 }),
  .out1({ S872 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_349_ (
  .in1({ S991, S980 }),
  .out1({ S873 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_412_ (
  .in1({ DP_ARU1_in1_9, DP_AC_dout_9 }),
  .out1({ S874 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_350_ (
  .in1({ DP_ARU1_in1_9, DP_AC_dout_9 }),
  .out1({ S875 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_413_ (
  .in1({ S991, S980 }),
  .out1({ S876 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_351_ (
  .in1({ S875, S873 }),
  .out1({ S877 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_414_ (
  .in1({ S876, S874 }),
  .out1({ S878 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_415_ (
  .in1({ S878, S872 }),
  .out1({ S879 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_416_ (
  .in1({ S877, S870 }),
  .out1({ S880 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_417_ (
  .in1({ S880, S879 }),
  .out1({ S881 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_352_ (
  .in1({ S863, S857 }),
  .out1({ S883 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_418_ (
  .in1({ S864, S858 }),
  .out1({ S884 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_353_ (
  .in1({ S848, S844 }),
  .out1({ S885 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_143_ (
  .in1({ S885 }),
  .out1({ S886 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_354_ (
  .in1({ S786, S780 }),
  .out1({ S887 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_144_ (
  .in1({ S887 }),
  .out1({ S888 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_355_ (
  .in1({ S837, S831 }),
  .out1({ S889 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_419_ (
  .in1({ S838, S832 }),
  .out1({ S890 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_420_ (
  .in1({ DP_ARU1_in1_7, DP_AC_dout_2 }),
  .out1({ S891 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_421_ (
  .in1({ DP_ARU1_in1_6, DP_AC_dout_3 }),
  .out1({ S892 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_356_ (
  .in1({ S800, S796 }),
  .out1({ S894 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_422_ (
  .in1({ S894, S892 }),
  .out1({ S895 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_357_ (
  .in1({ S894, S892 }),
  .out1({ S896 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_145_ (
  .in1({ S896 }),
  .out1({ S897 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_423_ (
  .in1({ S897, S895 }),
  .out1({ S898 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_424_ (
  .in1({ S898, S891 }),
  .out1({ S899 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_146_ (
  .in1({ S899 }),
  .out1({ S900 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_358_ (
  .in1({ S898, S891 }),
  .out1({ S901 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_147_ (
  .in1({ S901 }),
  .out1({ S902 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_359_ (
  .in1({ S901, S900 }),
  .out1({ S903 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_425_ (
  .in1({ S902, S899 }),
  .out1({ S905 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_360_ (
  .in1({ S824, S818 }),
  .out1({ S906 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_426_ (
  .in1({ S825, S819 }),
  .out1({ S907 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_427_ (
  .in1({ DP_ARU1_in1_5, DP_AC_dout_4 }),
  .out1({ S908 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_428_ (
  .in1({ DP_AC_dout_6, DP_ARU1_in1_3 }),
  .out1({ S909 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_429_ (
  .in1({ DP_AC_dout_6, DP_ARU1_in1_4 }),
  .out1({ S910 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_148_ (
  .in1({ S910 }),
  .out1({ S911 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_361_ (
  .in1({ S910, S793 }),
  .out1({ S912 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_149_ (
  .in1({ S912 }),
  .out1({ S913 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_430_ (
  .in1({ S909, S794 }),
  .out1({ S914 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_431_ (
  .in1({ S914, S913 }),
  .out1({ S916 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_362_ (
  .in1({ S916, S908 }),
  .out1({ S917 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_150_ (
  .in1({ S917 }),
  .out1({ S918 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_432_ (
  .in1({ S916, S908 }),
  .out1({ S919 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_151_ (
  .in1({ S919 }),
  .out1({ S920 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_363_ (
  .in1({ S920, S917 }),
  .out1({ S921 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_433_ (
  .in1({ S919, S918 }),
  .out1({ S922 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_364_ (
  .in1({ S812, S590 }),
  .out1({ S923 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_434_ (
  .in1({ S811, S591 }),
  .out1({ S924 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_365_ (
  .in1({ S924, S922 }),
  .out1({ S925 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_435_ (
  .in1({ S923, S921 }),
  .out1({ S927 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_366_ (
  .in1({ S923, S921 }),
  .out1({ S928 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_436_ (
  .in1({ S924, S922 }),
  .out1({ S929 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_367_ (
  .in1({ S928, S925 }),
  .out1({ S930 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_437_ (
  .in1({ S929, S927 }),
  .out1({ S931 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_368_ (
  .in1({ S931, S906 }),
  .out1({ S932 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_438_ (
  .in1({ S930, S907 }),
  .out1({ S933 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_369_ (
  .in1({ S930, S907 }),
  .out1({ S934 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_439_ (
  .in1({ S931, S906 }),
  .out1({ S935 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_370_ (
  .in1({ S934, S932 }),
  .out1({ S936 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_440_ (
  .in1({ S935, S933 }),
  .out1({ S938 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_371_ (
  .in1({ S938, S905 }),
  .out1({ S939 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_441_ (
  .in1({ S936, S903 }),
  .out1({ S940 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_372_ (
  .in1({ S936, S903 }),
  .out1({ S941 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_442_ (
  .in1({ S938, S905 }),
  .out1({ S942 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_373_ (
  .in1({ S941, S939 }),
  .out1({ S943 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_443_ (
  .in1({ S942, S940 }),
  .out1({ S944 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_374_ (
  .in1({ S944, S889 }),
  .out1({ S945 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_444_ (
  .in1({ S943, S890 }),
  .out1({ S946 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_445_ (
  .in1({ S944, S889 }),
  .out1({ S947 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_446_ (
  .in1({ S947, S946 }),
  .out1({ S949 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_152_ (
  .in1({ S949 }),
  .out1({ S950 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_447_ (
  .in1({ S950, S888 }),
  .out1({ S951 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_153_ (
  .in1({ S951 }),
  .out1({ S952 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_448_ (
  .in1({ S949, S887 }),
  .out1({ S953 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_449_ (
  .in1({ S953, S951 }),
  .out1({ S954 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_154_ (
  .in1({ S954 }),
  .out1({ S955 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_450_ (
  .in1({ S955, S886 }),
  .out1({ S956 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_155_ (
  .in1({ S956 }),
  .out1({ S957 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_451_ (
  .in1({ S954, S885 }),
  .out1({ S958 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_452_ (
  .in1({ S958, S956 }),
  .out1({ S960 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_156_ (
  .in1({ S960 }),
  .out1({ S961 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_375_ (
  .in1({ S961, S884 }),
  .out1({ S962 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_376_ (
  .in1({ S960, S883 }),
  .out1({ S963 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_453_ (
  .in1({ S961, S884 }),
  .out1({ S964 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_377_ (
  .in1({ S963, S962 }),
  .out1({ S965 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_378_ (
  .in1({ S965, CU_ADD }),
  .out1({ S966 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_379_ (
  .in1({ S881, S795 }),
  .out1({ S967 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_380_ (
  .in1({ S967, S966 }),
  .out1({ DP_ARU1_out_9 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_454_ (
  .in1({ DP_ARU1_in1_10, DP_AC_dout_10 }),
  .out1({ S968 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_381_ (
  .in1({ DP_ARU1_in1_10, DP_AC_dout_10 }),
  .out1({ S970 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_157_ (
  .in1({ S970 }),
  .out1({ S971 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_455_ (
  .in1({ S971, S968 }),
  .out1({ S972 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_158_ (
  .in1({ S972 }),
  .out1({ S973 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_382_ (
  .in1({ S873, S872 }),
  .out1({ S974 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_456_ (
  .in1({ S874, S870 }),
  .out1({ S975 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_383_ (
  .in1({ S974, S875 }),
  .out1({ S976 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_457_ (
  .in1({ S975, S876 }),
  .out1({ S977 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_458_ (
  .in1({ S976, S973 }),
  .out1({ S978 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_459_ (
  .in1({ S977, S972 }),
  .out1({ S979 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_460_ (
  .in1({ S979, S978 }),
  .out1({ S981 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_461_ (
  .in1({ S981, CU_ADD }),
  .out1({ S982 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_384_ (
  .in1({ S963, S957 }),
  .out1({ S983 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_462_ (
  .in1({ S964, S956 }),
  .out1({ S984 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_385_ (
  .in1({ S952, S945 }),
  .out1({ S985 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_159_ (
  .in1({ S985 }),
  .out1({ S986 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_386_ (
  .in1({ S901, S896 }),
  .out1({ S987 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_387_ (
  .in1({ S939, S932 }),
  .out1({ S988 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_463_ (
  .in1({ DP_ARU1_in1_7, DP_AC_dout_3 }),
  .out1({ S989 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_464_ (
  .in1({ DP_ARU1_in1_6, DP_AC_dout_4 }),
  .out1({ S990 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_388_ (
  .in1({ S917, S912 }),
  .out1({ S992 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_465_ (
  .in1({ S992, S990 }),
  .out1({ S993 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_389_ (
  .in1({ S992, S990 }),
  .out1({ S994 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_160_ (
  .in1({ S994 }),
  .out1({ S995 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_466_ (
  .in1({ S995, S993 }),
  .out1({ S996 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_467_ (
  .in1({ S996, S989 }),
  .out1({ S997 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_161_ (
  .in1({ S997 }),
  .out1({ S998 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_390_ (
  .in1({ S996, S989 }),
  .out1({ S999 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_162_ (
  .in1({ S999 }),
  .out1({ S1000 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_391_ (
  .in1({ S999, S998 }),
  .out1({ S1001 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_468_ (
  .in1({ S1000, S997 }),
  .out1({ S1003 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_392_ (
  .in1({ S925, S813 }),
  .out1({ S1004 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_469_ (
  .in1({ S927, S814 }),
  .out1({ S1005 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_470_ (
  .in1({ DP_AC_dout_7, DP_ARU1_in1_3 }),
  .out1({ S1006 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_471_ (
  .in1({ DP_AC_dout_7, DP_ARU1_in1_4 }),
  .out1({ S1007 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_393_ (
  .in1({ S1007, S909 }),
  .out1({ S1008 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_163_ (
  .in1({ S1008 }),
  .out1({ S1009 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_472_ (
  .in1({ S1006, S910 }),
  .out1({ S1010 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_164_ (
  .in1({ S1010 }),
  .out1({ S1011 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_394_ (
  .in1({ S1011, S1008 }),
  .out1({ S1012 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_473_ (
  .in1({ S1010, S1009 }),
  .out1({ S1014 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_395_ (
  .in1({ S1014, S476 }),
  .out1({ S1015 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_165_ (
  .in1({ S1015 }),
  .out1({ S1016 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_396_ (
  .in1({ S1012, S475 }),
  .out1({ S1017 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_474_ (
  .in1({ S1014, S476 }),
  .out1({ S1018 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_397_ (
  .in1({ S1017, S1015 }),
  .out1({ S1019 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_475_ (
  .in1({ S1018, S1016 }),
  .out1({ S1020 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_398_ (
  .in1({ S1020, S1004 }),
  .out1({ S1021 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_476_ (
  .in1({ S1019, S1005 }),
  .out1({ S1022 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_399_ (
  .in1({ S1019, S1005 }),
  .out1({ S1023 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_477_ (
  .in1({ S1020, S1004 }),
  .out1({ S1025 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_400_ (
  .in1({ S1023, S1021 }),
  .out1({ S1026 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_478_ (
  .in1({ S1025, S1022 }),
  .out1({ S1027 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_401_ (
  .in1({ S1027, S1003 }),
  .out1({ S1028 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_479_ (
  .in1({ S1026, S1001 }),
  .out1({ S1029 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_480_ (
  .in1({ S1027, S1003 }),
  .out1({ S1030 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_481_ (
  .in1({ S1030, S1029 }),
  .out1({ S1031 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_402_ (
  .in1({ S1031, S988 }),
  .out1({ S1032 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_166_ (
  .in1({ S1032 }),
  .out1({ S1033 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_482_ (
  .in1({ S1031, S988 }),
  .out1({ S1034 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_483_ (
  .in1({ S1034, S1033 }),
  .out1({ S1036 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_403_ (
  .in1({ S1036, S987 }),
  .out1({ S1037 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_167_ (
  .in1({ S1037 }),
  .out1({ S1038 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_484_ (
  .in1({ S1036, S987 }),
  .out1({ S1039 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_485_ (
  .in1({ S1039, S1038 }),
  .out1({ S1040 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_168_ (
  .in1({ S1040 }),
  .out1({ S1041 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_486_ (
  .in1({ S1040, S985 }),
  .out1({ S1042 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_487_ (
  .in1({ S1041, S986 }),
  .out1({ S1043 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_169_ (
  .in1({ S1043 }),
  .out1({ S1044 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_488_ (
  .in1({ S1043, S1042 }),
  .out1({ S1045 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_170_ (
  .in1({ S1045 }),
  .out1({ S1047 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_404_ (
  .in1({ S1047, S984 }),
  .out1({ S1048 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_405_ (
  .in1({ S1045, S983 }),
  .out1({ S1049 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_489_ (
  .in1({ S1047, S984 }),
  .out1({ S1050 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_406_ (
  .in1({ S1049, S1048 }),
  .out1({ S1051 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_407_ (
  .in1({ S1051, CU_ADD }),
  .out1({ S1052 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_171_ (
  .in1({ S1052 }),
  .out1({ S1053 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_490_ (
  .in1({ S1053, S982 }),
  .out1({ S1054 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_172_ (
  .in1({ S1054 }),
  .out1({ DP_ARU1_out_10 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_491_ (
  .in1({ S978, S968 }),
  .out1({ S1055 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_173_ (
  .in1({ S1055 }),
  .out1({ S1057 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_408_ (
  .in1({ S1013, S1002 }),
  .out1({ S1058 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_492_ (
  .in1({ DP_ARU1_in1_11, DP_AC_dout_11 }),
  .out1({ S1059 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_409_ (
  .in1({ DP_ARU1_in1_11, DP_AC_dout_11 }),
  .out1({ S1060 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_174_ (
  .in1({ S1060 }),
  .out1({ S1061 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_410_ (
  .in1({ S1060, S1058 }),
  .out1({ S1062 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_493_ (
  .in1({ S1061, S1059 }),
  .out1({ S1063 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_494_ (
  .in1({ S1063, S1055 }),
  .out1({ S1064 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_495_ (
  .in1({ S1062, S1057 }),
  .out1({ S1065 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_496_ (
  .in1({ S1065, S1064 }),
  .out1({ S1066 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_411_ (
  .in1({ S1049, S1044 }),
  .out1({ S1068 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_497_ (
  .in1({ S1050, S1043 }),
  .out1({ S1069 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_412_ (
  .in1({ S1037, S1032 }),
  .out1({ S1070 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_175_ (
  .in1({ S1070 }),
  .out1({ S1071 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_413_ (
  .in1({ S999, S994 }),
  .out1({ S1072 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_176_ (
  .in1({ S1072 }),
  .out1({ S1073 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_414_ (
  .in1({ S1028, S1021 }),
  .out1({ S1074 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_177_ (
  .in1({ S1074 }),
  .out1({ S1075 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_498_ (
  .in1({ DP_ARU1_in1_7, DP_AC_dout_4 }),
  .out1({ S1076 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_499_ (
  .in1({ DP_ARU1_in1_6, DP_AC_dout_5 }),
  .out1({ S1077 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_415_ (
  .in1({ S1015, S1008 }),
  .out1({ S1079 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_500_ (
  .in1({ S1079, S1077 }),
  .out1({ S1080 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_416_ (
  .in1({ S1079, S1077 }),
  .out1({ S1081 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_178_ (
  .in1({ S1081 }),
  .out1({ S1082 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_501_ (
  .in1({ S1082, S1080 }),
  .out1({ S1083 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_502_ (
  .in1({ S1083, S1076 }),
  .out1({ S1084 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_179_ (
  .in1({ S1084 }),
  .out1({ S1085 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_417_ (
  .in1({ S1083, S1076 }),
  .out1({ S1086 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_180_ (
  .in1({ S1086 }),
  .out1({ S1087 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_418_ (
  .in1({ S1086, S1085 }),
  .out1({ S1088 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_503_ (
  .in1({ S1087, S1084 }),
  .out1({ S1090 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_504_ (
  .in1({ DP_AC_dout_6, DP_ARU1_in1_5 }),
  .out1({ S1091 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_419_ (
  .in1({ S937, S904 }),
  .out1({ S1092 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_505_ (
  .in1({ DP_AC_dout_7, DP_ARU1_in1_5 }),
  .out1({ S1093 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_420_ (
  .in1({ S1093, S910 }),
  .out1({ S1094 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_506_ (
  .in1({ S1092, S911 }),
  .out1({ S1095 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_507_ (
  .in1({ S1091, S1007 }),
  .out1({ S1096 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_181_ (
  .in1({ S1096 }),
  .out1({ S1097 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_421_ (
  .in1({ S1097, S1094 }),
  .out1({ S1098 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_508_ (
  .in1({ S1096, S1095 }),
  .out1({ S1099 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_422_ (
  .in1({ S1099, S1090 }),
  .out1({ S1101 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_509_ (
  .in1({ S1098, S1088 }),
  .out1({ S1102 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_510_ (
  .in1({ S1099, S1090 }),
  .out1({ S1103 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_511_ (
  .in1({ S1103, S1102 }),
  .out1({ S1104 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_182_ (
  .in1({ S1104 }),
  .out1({ S1105 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_512_ (
  .in1({ S1105, S1075 }),
  .out1({ S1106 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_183_ (
  .in1({ S1106 }),
  .out1({ S1107 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_513_ (
  .in1({ S1104, S1074 }),
  .out1({ S1108 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_514_ (
  .in1({ S1108, S1106 }),
  .out1({ S1109 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_184_ (
  .in1({ S1109 }),
  .out1({ S1110 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_515_ (
  .in1({ S1110, S1073 }),
  .out1({ S1112 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_185_ (
  .in1({ S1112 }),
  .out1({ S1113 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_516_ (
  .in1({ S1109, S1072 }),
  .out1({ S1114 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_517_ (
  .in1({ S1114, S1112 }),
  .out1({ S1115 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_186_ (
  .in1({ S1115 }),
  .out1({ S1116 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_518_ (
  .in1({ S1115, S1070 }),
  .out1({ S1117 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_519_ (
  .in1({ S1116, S1071 }),
  .out1({ S1118 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_187_ (
  .in1({ S1118 }),
  .out1({ S1119 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_520_ (
  .in1({ S1118, S1117 }),
  .out1({ S1120 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_188_ (
  .in1({ S1120 }),
  .out1({ S1121 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_423_ (
  .in1({ S1121, S1069 }),
  .out1({ S1123 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_424_ (
  .in1({ S1120, S1068 }),
  .out1({ S1124 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_521_ (
  .in1({ S1121, S1069 }),
  .out1({ S1125 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_425_ (
  .in1({ S1124, S1123 }),
  .out1({ S1126 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_426_ (
  .in1({ S1126, CU_ADD }),
  .out1({ S1127 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_427_ (
  .in1({ S1066, S795 }),
  .out1({ S1128 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_428_ (
  .in1({ S1128, S1127 }),
  .out1({ DP_ARU1_out_11 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_522_ (
  .in1({ DP_ARU1_in1_12, DP_AC_dout_12 }),
  .out1({ S1129 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_189_ (
  .in1({ S1129 }),
  .out1({ S1130 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_429_ (
  .in1({ DP_ARU1_in1_12, DP_AC_dout_12 }),
  .out1({ S1131 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_430_ (
  .in1({ S1131, S1130 }),
  .out1({ S1132 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_431_ (
  .in1({ S1058, S1055 }),
  .out1({ S1133 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_432_ (
  .in1({ S1133, S1060 }),
  .out1({ S1134 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_523_ (
  .in1({ S1134, S1132 }),
  .out1({ S1135 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_433_ (
  .in1({ S1134, S1132 }),
  .out1({ S1136 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_434_ (
  .in1({ S1124, S1119 }),
  .out1({ S1137 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_524_ (
  .in1({ S1125, S1118 }),
  .out1({ S1138 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_435_ (
  .in1({ S1113, S1107 }),
  .out1({ S1139 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_190_ (
  .in1({ S1139 }),
  .out1({ S1140 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_436_ (
  .in1({ S1086, S1081 }),
  .out1({ S1141 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_191_ (
  .in1({ S1141 }),
  .out1({ S1143 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_525_ (
  .in1({ DP_ARU1_in1_7, DP_AC_dout_5 }),
  .out1({ S1144 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_192_ (
  .in1({ S1144 }),
  .out1({ S1145 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_526_ (
  .in1({ S1095, S554 }),
  .out1({ S1146 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_527_ (
  .in1({ S1094, DP_ARU1_in1_6 }),
  .out1({ S1147 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_193_ (
  .in1({ S1147 }),
  .out1({ S1148 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_528_ (
  .in1({ S1147, S1146 }),
  .out1({ S1149 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_194_ (
  .in1({ S1149 }),
  .out1({ S1150 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_529_ (
  .in1({ S1149, S1144 }),
  .out1({ S1151 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_195_ (
  .in1({ S1151 }),
  .out1({ S1152 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_437_ (
  .in1({ S1149, S1144 }),
  .out1({ S1154 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_530_ (
  .in1({ S1150, S1145 }),
  .out1({ S1155 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_438_ (
  .in1({ S1154, S1152 }),
  .out1({ S1156 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_531_ (
  .in1({ S1155, S1151 }),
  .out1({ S1157 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_439_ (
  .in1({ S1157, S1093 }),
  .out1({ S1158 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_532_ (
  .in1({ S1156, S1092 }),
  .out1({ S1159 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_533_ (
  .in1({ S1157, S1093 }),
  .out1({ S1160 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_534_ (
  .in1({ S1160, S1159 }),
  .out1({ S1161 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_196_ (
  .in1({ S1161 }),
  .out1({ S1162 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_535_ (
  .in1({ S1161, S1102 }),
  .out1({ S1163 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_536_ (
  .in1({ S1162, S1101 }),
  .out1({ S1165 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_197_ (
  .in1({ S1165 }),
  .out1({ S1166 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_537_ (
  .in1({ S1165, S1163 }),
  .out1({ S1167 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_198_ (
  .in1({ S1167 }),
  .out1({ S1168 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_538_ (
  .in1({ S1167, S1141 }),
  .out1({ S1169 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_440_ (
  .in1({ S1167, S1141 }),
  .out1({ S1170 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_539_ (
  .in1({ S1168, S1143 }),
  .out1({ S1171 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_540_ (
  .in1({ S1171, S1169 }),
  .out1({ S1172 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_199_ (
  .in1({ S1172 }),
  .out1({ S1173 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_541_ (
  .in1({ S1172, S1139 }),
  .out1({ S1174 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_542_ (
  .in1({ S1173, S1140 }),
  .out1({ S1176 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_200_ (
  .in1({ S1176 }),
  .out1({ S1177 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_543_ (
  .in1({ S1176, S1174 }),
  .out1({ S1178 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_201_ (
  .in1({ S1178 }),
  .out1({ S1179 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_544_ (
  .in1({ S1178, S1137 }),
  .out1({ S1180 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_441_ (
  .in1({ S1178, S1137 }),
  .out1({ S1181 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_545_ (
  .in1({ S1179, S1138 }),
  .out1({ S1182 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_546_ (
  .in1({ S1182, S1180 }),
  .out1({ S1183 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_442_ (
  .in1({ S1136, S795 }),
  .out1({ S1184 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_547_ (
  .in1({ S1184, S1135 }),
  .out1({ S1185 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_202_ (
  .in1({ S1185 }),
  .out1({ S1187 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_443_ (
  .in1({ S1183, CU_ADD }),
  .out1({ S1188 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_444_ (
  .in1({ S1188, S1187 }),
  .out1({ S1189 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_203_ (
  .in1({ S1189 }),
  .out1({ DP_ARU1_out_12 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_548_ (
  .in1({ S1135, S1129 }),
  .out1({ S1190 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_549_ (
  .in1({ DP_ARU1_in1_13, DP_AC_dout_13 }),
  .out1({ S1191 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_445_ (
  .in1({ DP_ARU1_in1_13, DP_AC_dout_13 }),
  .out1({ S1192 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_204_ (
  .in1({ S1192 }),
  .out1({ S1193 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_550_ (
  .in1({ S1193, S1191 }),
  .out1({ S1194 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_551_ (
  .in1({ S1194, S1190 }),
  .out1({ S1195 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_446_ (
  .in1({ S1194, S1190 }),
  .out1({ S1197 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_447_ (
  .in1({ S1181, S1177 }),
  .out1({ S1198 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_552_ (
  .in1({ S1182, S1176 }),
  .out1({ S1199 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_448_ (
  .in1({ S1170, S1166 }),
  .out1({ S1200 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_553_ (
  .in1({ S1171, S1165 }),
  .out1({ S1201 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_449_ (
  .in1({ S1154, S1148 }),
  .out1({ S1202 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_554_ (
  .in1({ S1155, S1147 }),
  .out1({ S1203 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_555_ (
  .in1({ DP_ARU1_in1_7, DP_AC_dout_6 }),
  .out1({ S1204 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_556_ (
  .in1({ DP_AC_dout_7, DP_ARU1_in1_6 }),
  .out1({ S1205 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_450_ (
  .in1({ S653, S554 }),
  .out1({ S1206 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_205_ (
  .in1({ S1206 }),
  .out1({ S1208 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_557_ (
  .in1({ S1205, S1204 }),
  .out1({ S1209 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_206_ (
  .in1({ S1209 }),
  .out1({ S1210 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_451_ (
  .in1({ S1210, S1206 }),
  .out1({ S1211 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_558_ (
  .in1({ S1209, S1208 }),
  .out1({ S1212 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_452_ (
  .in1({ S1211, S1158 }),
  .out1({ S1213 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_559_ (
  .in1({ S1212, S1159 }),
  .out1({ S1214 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_560_ (
  .in1({ S1211, S1158 }),
  .out1({ S1215 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_207_ (
  .in1({ S1215 }),
  .out1({ S1216 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_453_ (
  .in1({ S1216, S1213 }),
  .out1({ S1217 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_561_ (
  .in1({ S1215, S1214 }),
  .out1({ S1219 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_454_ (
  .in1({ S1217, S1203 }),
  .out1({ S1220 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_562_ (
  .in1({ S1219, S1202 }),
  .out1({ S1221 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_563_ (
  .in1({ S1217, S1203 }),
  .out1({ S1222 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_208_ (
  .in1({ S1222 }),
  .out1({ S1223 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_455_ (
  .in1({ S1223, S1220 }),
  .out1({ S1224 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_564_ (
  .in1({ S1222, S1221 }),
  .out1({ S1225 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_456_ (
  .in1({ S1224, S1201 }),
  .out1({ S1226 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_457_ (
  .in1({ S1225, S1200 }),
  .out1({ S1227 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_458_ (
  .in1({ S1227, S1226 }),
  .out1({ S1228 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_459_ (
  .in1({ S1228, S1198 }),
  .out1({ S1230 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_565_ (
  .in1({ S1228, S1198 }),
  .out1({ S1231 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_566_ (
  .in1({ S1195, CU_ADD }),
  .out1({ S1232 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_460_ (
  .in1({ S1232, S1197 }),
  .out1({ S1233 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_567_ (
  .in1({ S1231, S795 }),
  .out1({ S1234 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_461_ (
  .in1({ S1234, S1230 }),
  .out1({ S1235 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_462_ (
  .in1({ S1235, S1233 }),
  .out1({ DP_ARU1_out_13 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_463_ (
  .in1({ S1035, S1024 }),
  .out1({ S1236 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_464_ (
  .in1({ DP_ARU1_in1_14, DP_AC_dout_14 }),
  .out1({ S1237 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_465_ (
  .in1({ S1237, S1236 }),
  .out1({ S1238 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_209_ (
  .in1({ S1238 }),
  .out1({ S1240 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_568_ (
  .in1({ S1193, S1190 }),
  .out1({ S1241 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_569_ (
  .in1({ S1241, S1191 }),
  .out1({ S1242 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_210_ (
  .in1({ S1242 }),
  .out1({ S1243 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_466_ (
  .in1({ S1243, S1240 }),
  .out1({ S1244 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_467_ (
  .in1({ S1242, S1238 }),
  .out1({ S1245 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_468_ (
  .in1({ S1245, S1244 }),
  .out1({ S1246 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_469_ (
  .in1({ S1246, S795 }),
  .out1({ S1247 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_570_ (
  .in1({ S1222, S1215 }),
  .out1({ S1248 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_211_ (
  .in1({ S1248 }),
  .out1({ S1249 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_470_ (
  .in1({ S653, S553 }),
  .out1({ S1251 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_571_ (
  .in1({ S652, S554 }),
  .out1({ S1252 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_471_ (
  .in1({ S1251, S1248 }),
  .out1({ S1253 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_472_ (
  .in1({ S1252, S1249 }),
  .out1({ S1254 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_473_ (
  .in1({ S1254, S1253 }),
  .out1({ S1255 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_212_ (
  .in1({ S1255 }),
  .out1({ S1256 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_474_ (
  .in1({ S1226, S1198 }),
  .out1({ S1257 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_475_ (
  .in1({ S1227, S1199 }),
  .out1({ S1258 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_476_ (
  .in1({ S1257, S1227 }),
  .out1({ S1259 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_477_ (
  .in1({ S1258, S1226 }),
  .out1({ S1260 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_478_ (
  .in1({ S1260, S1255 }),
  .out1({ S1262 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_479_ (
  .in1({ S1259, S1256 }),
  .out1({ S1263 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_572_ (
  .in1({ S1260, S1255 }),
  .out1({ S1264 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_480_ (
  .in1({ S1263, S1262 }),
  .out1({ S1265 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_481_ (
  .in1({ S1265, CU_ADD }),
  .out1({ S1266 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_482_ (
  .in1({ S1266, S1247 }),
  .out1({ DP_ARU1_out_14 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_483_ (
  .in1({ S1206, CU_ADD }),
  .out1({ S1267 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_213_ (
  .in1({ S1267 }),
  .out1({ S1268 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_484_ (
  .in1({ S1268, S1254 }),
  .out1({ S1269 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_573_ (
  .in1({ S1269, S1264 }),
  .out1({ S1270 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_485_ (
  .in1({ S1056, S1046 }),
  .out1({ S312 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_574_ (
  .in1({ DP_ARU1_in1_15, DP_AC_dout_15 }),
  .out1({ S313 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_486_ (
  .in1({ DP_ARU1_in1_15, DP_AC_dout_15 }),
  .out1({ S314 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_487_ (
  .in1({ S314, S312 }),
  .out1({ S315 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_488_ (
  .in1({ S1244, S1236 }),
  .out1({ S316 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_575_ (
  .in1({ S316, S315 }),
  .out1({ S317 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_489_ (
  .in1({ S316, S315 }),
  .out1({ S318 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_490_ (
  .in1({ S318, S795 }),
  .out1({ S319 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_576_ (
  .in1({ S319, S317 }),
  .out1({ S320 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_577_ (
  .in1({ S320, S1270 }),
  .out1({ S321 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_214_ (
  .in1({ S321 }),
  .out1({ DP_ARU1_N })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_491_ (
  .in1({ DP_ARU1_out_1, DP_ARU1_out_0 }),
  .out1({ S323 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_578_ (
  .in1({ S323, S375 }),
  .out1({ S324 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_492_ (
  .in1({ S324, DP_ARU1_out_3 }),
  .out1({ S325 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_579_ (
  .in1({ S325, S473 }),
  .out1({ S326 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_493_ (
  .in1({ S326, DP_ARU1_out_5 }),
  .out1({ S327 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_580_ (
  .in1({ S327, S649 }),
  .out1({ S328 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_494_ (
  .in1({ S328, DP_ARU1_out_7 }),
  .out1({ S329 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_581_ (
  .in1({ S329, S869 }),
  .out1({ S330 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_495_ (
  .in1({ S330, DP_ARU1_out_9 }),
  .out1({ S331 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_582_ (
  .in1({ S331, S1054 }),
  .out1({ S333 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_496_ (
  .in1({ S333, DP_ARU1_out_11 }),
  .out1({ S334 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_583_ (
  .in1({ S334, S1189 }),
  .out1({ S335 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_497_ (
  .in1({ S335, DP_ARU1_out_13 }),
  .out1({ S336 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_584_ (
  .in1({ S336, S321 }),
  .out1({ S337 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_498_ (
  .in1({ S337, DP_ARU1_out_14 }),
  .out1({ DP_ARU1_Z })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_585_ (
  .in1({ DP_ARU1_N, S314 }),
  .out1({ S338 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_586_ (
  .in1({ S321, S312 }),
  .out1({ S339 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_587_ (
  .in1({ S339, S338 }),
  .out1({ DP_ARU1_V })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_588_ (
  .in1({ S316, S313 }),
  .out1({ S340 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_589_ (
  .in1({ S340, CU_ADD }),
  .out1({ S342 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_499_ (
  .in1({ S342, S314 }),
  .out1({ DP_ARU1_C })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_215_ (
  .in1({ CU_inst_0 }),
  .out1({ S1272 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_216_ (
  .in1({ CU_SE12bits }),
  .out1({ S1273 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_217_ (
  .in1({ CU_conOF }),
  .out1({ S1274 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_218_ (
  .in1({ CU_inst_1 }),
  .out1({ S1275 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_219_ (
  .in1({ CU_inst_2 }),
  .out1({ S1276 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_220_ (
  .in1({ CU_inst_3 }),
  .out1({ S1277 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_500_ (
  .in1({ CU_SE12bits, CU_SE4bits }),
  .out1({ S1278 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_221_ (
  .in1({ S1278 }),
  .out1({ S1279 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_501_ (
  .in1({ S1279, CU_conOF }),
  .out1({ S1280 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_502_ (
  .in1({ S1280, S1272 }),
  .out1({ DP_IMM1_out_0 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_503_ (
  .in1({ S1280, S1275 }),
  .out1({ DP_IMM1_out_1 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_504_ (
  .in1({ S1280, S1276 }),
  .out1({ DP_IMM1_out_2 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_505_ (
  .in1({ S1280, S1277 }),
  .out1({ DP_IMM1_out_3 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_590_ (
  .in1({ S1273, CU_SE4bits }),
  .out1({ S1281 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_591_ (
  .in1({ S1281, S1274 }),
  .out1({ S1282 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_592_ (
  .in1({ S1282, CU_inst_4 }),
  .out1({ S1283 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_506_ (
  .in1({ CU_conOF, S1273 }),
  .out1({ S1284 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_593_ (
  .in1({ CU_inst_3, CU_SE12bits }),
  .out1({ S1285 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_507_ (
  .in1({ S1285, CU_conOF }),
  .out1({ S1286 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_594_ (
  .in1({ S1284, CU_inst_3 }),
  .out1({ S1287 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_595_ (
  .in1({ S1287, S1283 }),
  .out1({ DP_IMM1_out_4 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_596_ (
  .in1({ S1282, CU_inst_5 }),
  .out1({ S1288 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_597_ (
  .in1({ S1288, S1287 }),
  .out1({ DP_IMM1_out_5 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_598_ (
  .in1({ S1282, CU_inst_6 }),
  .out1({ S1289 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_599_ (
  .in1({ S1289, S1287 }),
  .out1({ DP_IMM1_out_6 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_600_ (
  .in1({ S1282, CU_inst_7 }),
  .out1({ S1290 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_601_ (
  .in1({ S1290, S1287 }),
  .out1({ DP_IMM1_out_7 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_602_ (
  .in1({ S1282, CU_inst_8 }),
  .out1({ S1291 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_603_ (
  .in1({ S1291, S1287 }),
  .out1({ DP_IMM1_out_8 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_604_ (
  .in1({ S1282, CU_inst_9 }),
  .out1({ S1292 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_605_ (
  .in1({ S1292, S1287 }),
  .out1({ DP_IMM1_out_9 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_606_ (
  .in1({ S1282, CU_inst_10 }),
  .out1({ S1293 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_607_ (
  .in1({ S1293, S1287 }),
  .out1({ DP_IMM1_out_10 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_608_ (
  .in1({ S1282, CU_inst_11 }),
  .out1({ S1294 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_609_ (
  .in1({ S1294, S1287 }),
  .out1({ DP_IMM1_out_11 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_610_ (
  .in1({ S1278, CU_LSB0E }),
  .out1({ S1295 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_611_ (
  .in1({ S1295, S1274 }),
  .out1({ S1296 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_612_ (
  .in1({ S1296, DP_IMM1_in1_0 }),
  .out1({ S1297 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_613_ (
  .in1({ CU_inst_11, S1274 }),
  .out1({ S1298 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_508_ (
  .in1({ S1298, S1281 }),
  .out1({ S1299 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_509_ (
  .in1({ S1299, S1286 }),
  .out1({ S1300 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_614_ (
  .in1({ S1300, S1297 }),
  .out1({ DP_IMM1_out_12 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_615_ (
  .in1({ S1296, DP_IMM1_in1_1 }),
  .out1({ S1301 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_616_ (
  .in1({ S1301, S1300 }),
  .out1({ DP_IMM1_out_13 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_617_ (
  .in1({ S1296, DP_IMM1_in1_2 }),
  .out1({ S1302 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_618_ (
  .in1({ S1302, S1300 }),
  .out1({ DP_IMM1_out_14 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_619_ (
  .in1({ S1296, DP_IMM1_in1_3 }),
  .out1({ S1303 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_620_ (
  .in1({ S1303, S1300 }),
  .out1({ DP_IMM1_out_15 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_222_ (
  .in1({ CU_ldIN }),
  .out1({ S1321 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_510_ (
  .in1({ CU_ldIN, S6 }),
  .out1({ S1322 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_621_ (
  .in1({ S1322, DP_IN_dout_0 }),
  .out1({ S1323 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_511_ (
  .in1({ S1321, S7 }),
  .out1({ S1324 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_622_ (
  .in1({ S1324, DP_IN_din_0 }),
  .out1({ S1325 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_623_ (
  .in1({ S1325, S1323 }),
  .out1({ S1304 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_624_ (
  .in1({ S1322, DP_IN_dout_1 }),
  .out1({ S1326 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_625_ (
  .in1({ S1324, DP_IN_din_1 }),
  .out1({ S1327 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_626_ (
  .in1({ S1327, S1326 }),
  .out1({ S1305 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_627_ (
  .in1({ S1322, DP_IN_dout_2 }),
  .out1({ S1328 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_628_ (
  .in1({ S1324, DP_IN_din_2 }),
  .out1({ S1329 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_629_ (
  .in1({ S1329, S1328 }),
  .out1({ S1306 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_630_ (
  .in1({ S1322, DP_IN_dout_3 }),
  .out1({ S1330 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_631_ (
  .in1({ S1324, DP_IN_din_3 }),
  .out1({ S1331 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_632_ (
  .in1({ S1331, S1330 }),
  .out1({ S1307 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_633_ (
  .in1({ S1322, DP_IN_dout_4 }),
  .out1({ S1332 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_634_ (
  .in1({ S1324, DP_IN_din_4 }),
  .out1({ S1333 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_635_ (
  .in1({ S1333, S1332 }),
  .out1({ S1308 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_636_ (
  .in1({ S1322, DP_IN_dout_5 }),
  .out1({ S1334 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_637_ (
  .in1({ S1324, DP_IN_din_5 }),
  .out1({ S1335 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_638_ (
  .in1({ S1335, S1334 }),
  .out1({ S1309 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_639_ (
  .in1({ S1322, DP_IN_dout_6 }),
  .out1({ S1336 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_640_ (
  .in1({ S1324, DP_IN_din_6 }),
  .out1({ S1337 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_641_ (
  .in1({ S1337, S1336 }),
  .out1({ S1310 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_642_ (
  .in1({ S1322, DP_IN_dout_7 }),
  .out1({ S1338 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_643_ (
  .in1({ S1324, DP_IN_din_7 }),
  .out1({ S1339 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_644_ (
  .in1({ S1339, S1338 }),
  .out1({ S1311 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_645_ (
  .in1({ S1322, DP_IN_dout_8 }),
  .out1({ S1340 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_646_ (
  .in1({ S1324, DP_IN_din_8 }),
  .out1({ S1341 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_647_ (
  .in1({ S1341, S1340 }),
  .out1({ S1312 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_648_ (
  .in1({ S1322, DP_IN_dout_9 }),
  .out1({ S1342 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_649_ (
  .in1({ S1324, DP_IN_din_9 }),
  .out1({ S1343 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_650_ (
  .in1({ S1343, S1342 }),
  .out1({ S1313 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_651_ (
  .in1({ S1322, DP_IN_dout_10 }),
  .out1({ S1344 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_652_ (
  .in1({ S1324, DP_IN_din_10 }),
  .out1({ S1345 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_653_ (
  .in1({ S1345, S1344 }),
  .out1({ S1314 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_654_ (
  .in1({ S1322, DP_IN_dout_11 }),
  .out1({ S1346 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_655_ (
  .in1({ S1324, DP_IN_din_11 }),
  .out1({ S1347 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_656_ (
  .in1({ S1347, S1346 }),
  .out1({ S1315 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_657_ (
  .in1({ S1322, DP_IN_dout_12 }),
  .out1({ S1348 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_658_ (
  .in1({ S1324, DP_IN_din_12 }),
  .out1({ S1349 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_659_ (
  .in1({ S1349, S1348 }),
  .out1({ S1316 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_660_ (
  .in1({ S1322, DP_IN_dout_13 }),
  .out1({ S1350 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_661_ (
  .in1({ S1324, DP_IN_din_13 }),
  .out1({ S1351 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_662_ (
  .in1({ S1351, S1350 }),
  .out1({ S1317 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_663_ (
  .in1({ S1322, DP_IN_dout_14 }),
  .out1({ S1352 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_664_ (
  .in1({ S1324, DP_IN_din_14 }),
  .out1({ S1353 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_665_ (
  .in1({ S1353, S1352 }),
  .out1({ S1318 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_666_ (
  .in1({ S1322, DP_IN_dout_15 }),
  .out1({ S1354 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_667_ (
  .in1({ S1324, DP_IN_din_15 }),
  .out1({ S1320 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_668_ (
  .in1({ S1320, S1354 }),
  .out1({ S1319 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_19_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1304 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_dout_0 }),
  .Si({ S3057 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_20_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1305 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_dout_1 }),
  .Si({ S3056 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_21_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1306 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_dout_2 }),
  .Si({ S3055 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_22_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1307 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_dout_3 }),
  .Si({ S3054 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_23_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1308 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_dout_4 }),
  .Si({ S3053 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_24_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1309 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_dout_5 }),
  .Si({ S3052 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_25_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1310 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_dout_6 }),
  .Si({ S3051 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_26_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1311 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_dout_7 }),
  .Si({ S3050 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_27_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1312 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_dout_8 }),
  .Si({ S3049 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_28_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1313 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_dout_9 }),
  .Si({ S3048 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_29_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1314 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_dout_10 }),
  .Si({ S3047 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_30_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1315 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_dout_11 }),
  .Si({ S3046 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_31_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1316 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_dout_12 }),
  .Si({ S3045 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_32_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1317 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_dout_13 }),
  .Si({ S3044 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_33_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1318 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_dout_14 }),
  .Si({ S3043 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_34_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1319 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_dout_15 }),
  .Si({ S3092 }),
  .global_reset({ 1'b0 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_223_ (
  .in1({ DP_INC_1_in_0 }),
  .out1({ S1372 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_224_ (
  .in1({ DP_INC_1_inc_value_0 }),
  .out1({ S1373 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_225_ (
  .in1({ DP_INC_1_in_1 }),
  .out1({ S1374 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_226_ (
  .in1({ DP_INC_1_inc_value_1 }),
  .out1({ S1375 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_227_ (
  .in1({ DP_INC_1_in_2 }),
  .out1({ S1376 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_228_ (
  .in1({ DP_INC_1_in_3 }),
  .out1({ S1377 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_229_ (
  .in1({ DP_INC_1_in_4 }),
  .out1({ S1378 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_230_ (
  .in1({ DP_INC_1_in_5 }),
  .out1({ S1379 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_231_ (
  .in1({ DP_INC_1_in_6 }),
  .out1({ S1380 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_232_ (
  .in1({ DP_INC_1_in_7 }),
  .out1({ S1381 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_233_ (
  .in1({ DP_INC_1_in_8 }),
  .out1({ S1382 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_234_ (
  .in1({ DP_INC_1_in_9 }),
  .out1({ S1383 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_235_ (
  .in1({ DP_INC_1_in_10 }),
  .out1({ S1384 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_236_ (
  .in1({ DP_INC_1_in_11 }),
  .out1({ S1385 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_237_ (
  .in1({ DP_INC_1_in_12 }),
  .out1({ S1386 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_238_ (
  .in1({ DP_INC_1_in_13 }),
  .out1({ S1387 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_239_ (
  .in1({ DP_INC_1_in_14 }),
  .out1({ S1388 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_240_ (
  .in1({ DP_INC_1_in_15 }),
  .out1({ S1389 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_512_ (
  .in1({ S1373, S1372 }),
  .out1({ S1390 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_669_ (
  .in1({ DP_INC_1_inc_value_0, DP_INC_1_in_0 }),
  .out1({ S1391 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_513_ (
  .in1({ DP_INC_1_inc_value_0, DP_INC_1_in_0 }),
  .out1({ S1392 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_514_ (
  .in1({ S1392, S1390 }),
  .out1({ DP_INC_1_out_0 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_515_ (
  .in1({ S1375, S1374 }),
  .out1({ S1393 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_670_ (
  .in1({ DP_INC_1_inc_value_1, DP_INC_1_in_1 }),
  .out1({ S1394 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_516_ (
  .in1({ DP_INC_1_inc_value_1, DP_INC_1_in_1 }),
  .out1({ S1395 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_241_ (
  .in1({ S1395 }),
  .out1({ S1396 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_517_ (
  .in1({ S1395, S1393 }),
  .out1({ S1397 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_671_ (
  .in1({ S1396, S1394 }),
  .out1({ S1398 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_518_ (
  .in1({ S1398, S1391 }),
  .out1({ S1399 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_672_ (
  .in1({ S1397, S1390 }),
  .out1({ S1400 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_519_ (
  .in1({ S1397, S1390 }),
  .out1({ S1401 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_520_ (
  .in1({ S1401, S1399 }),
  .out1({ DP_INC_1_out_1 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_521_ (
  .in1({ S1399, S1393 }),
  .out1({ S1402 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_673_ (
  .in1({ S1400, S1394 }),
  .out1({ S1403 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_522_ (
  .in1({ S1402, S1376 }),
  .out1({ S1404 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_674_ (
  .in1({ S1403, DP_INC_1_in_2 }),
  .out1({ S1405 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_523_ (
  .in1({ S1403, DP_INC_1_in_2 }),
  .out1({ S1406 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_524_ (
  .in1({ S1406, S1404 }),
  .out1({ DP_INC_1_out_2 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_525_ (
  .in1({ S1405, S1377 }),
  .out1({ S1407 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_675_ (
  .in1({ S1404, DP_INC_1_in_3 }),
  .out1({ S1408 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_526_ (
  .in1({ S1404, DP_INC_1_in_3 }),
  .out1({ S1409 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_527_ (
  .in1({ S1409, S1407 }),
  .out1({ DP_INC_1_out_3 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_528_ (
  .in1({ S1408, S1378 }),
  .out1({ S1410 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_676_ (
  .in1({ S1407, DP_INC_1_in_4 }),
  .out1({ S1411 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_529_ (
  .in1({ S1407, DP_INC_1_in_4 }),
  .out1({ S1412 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_530_ (
  .in1({ S1412, S1410 }),
  .out1({ DP_INC_1_out_4 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_531_ (
  .in1({ S1411, S1379 }),
  .out1({ S1413 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_677_ (
  .in1({ S1410, DP_INC_1_in_5 }),
  .out1({ S1414 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_532_ (
  .in1({ S1410, DP_INC_1_in_5 }),
  .out1({ S1415 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_533_ (
  .in1({ S1415, S1413 }),
  .out1({ DP_INC_1_out_5 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_534_ (
  .in1({ S1414, S1380 }),
  .out1({ S1416 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_678_ (
  .in1({ S1413, DP_INC_1_in_6 }),
  .out1({ S1417 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_535_ (
  .in1({ S1413, DP_INC_1_in_6 }),
  .out1({ S1418 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_536_ (
  .in1({ S1418, S1416 }),
  .out1({ DP_INC_1_out_6 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_537_ (
  .in1({ S1417, S1381 }),
  .out1({ S1419 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_679_ (
  .in1({ S1416, DP_INC_1_in_7 }),
  .out1({ S1420 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_538_ (
  .in1({ S1416, DP_INC_1_in_7 }),
  .out1({ S1421 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_539_ (
  .in1({ S1421, S1419 }),
  .out1({ DP_INC_1_out_7 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_540_ (
  .in1({ S1420, S1382 }),
  .out1({ S1422 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_680_ (
  .in1({ S1419, DP_INC_1_in_8 }),
  .out1({ S1423 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_541_ (
  .in1({ S1419, DP_INC_1_in_8 }),
  .out1({ S1424 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_542_ (
  .in1({ S1424, S1422 }),
  .out1({ DP_INC_1_out_8 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_543_ (
  .in1({ S1423, S1383 }),
  .out1({ S1425 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_681_ (
  .in1({ S1422, DP_INC_1_in_9 }),
  .out1({ S1426 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_544_ (
  .in1({ S1422, DP_INC_1_in_9 }),
  .out1({ S1427 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_545_ (
  .in1({ S1427, S1425 }),
  .out1({ DP_INC_1_out_9 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_546_ (
  .in1({ S1426, S1384 }),
  .out1({ S1355 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_682_ (
  .in1({ S1425, DP_INC_1_in_10 }),
  .out1({ S1356 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_547_ (
  .in1({ S1425, DP_INC_1_in_10 }),
  .out1({ S1357 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_548_ (
  .in1({ S1357, S1355 }),
  .out1({ DP_INC_1_out_10 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_549_ (
  .in1({ S1356, S1385 }),
  .out1({ S1358 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_683_ (
  .in1({ S1355, DP_INC_1_in_11 }),
  .out1({ S1359 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_550_ (
  .in1({ S1355, DP_INC_1_in_11 }),
  .out1({ S1360 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_551_ (
  .in1({ S1360, S1358 }),
  .out1({ DP_INC_1_out_11 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_552_ (
  .in1({ S1359, S1386 }),
  .out1({ S1361 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_684_ (
  .in1({ S1358, DP_INC_1_in_12 }),
  .out1({ S1362 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_553_ (
  .in1({ S1358, DP_INC_1_in_12 }),
  .out1({ S1363 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_554_ (
  .in1({ S1363, S1361 }),
  .out1({ DP_INC_1_out_12 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_555_ (
  .in1({ S1362, S1387 }),
  .out1({ S1364 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_685_ (
  .in1({ S1361, DP_INC_1_in_13 }),
  .out1({ S1365 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_556_ (
  .in1({ S1361, DP_INC_1_in_13 }),
  .out1({ S1366 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_557_ (
  .in1({ S1366, S1364 }),
  .out1({ DP_INC_1_out_13 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_558_ (
  .in1({ S1365, S1388 }),
  .out1({ S1367 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_686_ (
  .in1({ S1364, DP_INC_1_in_14 }),
  .out1({ S1368 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_559_ (
  .in1({ S1364, DP_INC_1_in_14 }),
  .out1({ S1369 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_560_ (
  .in1({ S1369, S1367 }),
  .out1({ DP_INC_1_out_14 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_561_ (
  .in1({ S1367, DP_INC_1_in_15 }),
  .out1({ S1370 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_562_ (
  .in1({ S1368, S1389 }),
  .out1({ S1371 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_563_ (
  .in1({ S1371, S1370 }),
  .out1({ DP_INC_1_out_15 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_242_ (
  .in1({ dataBus[0] }),
  .out1({ S1445 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_243_ (
  .in1({ S0 }),
  .out1({ S1446 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_244_ (
  .in1({ dataBus[1] }),
  .out1({ S1447 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_245_ (
  .in1({ S8 }),
  .out1({ S1448 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_246_ (
  .in1({ dataBus[2] }),
  .out1({ S1449 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_247_ (
  .in1({ dataBus[3] }),
  .out1({ S1450 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_248_ (
  .in1({ dataBus[4] }),
  .out1({ S1451 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_249_ (
  .in1({ dataBus[5] }),
  .out1({ S1452 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_250_ (
  .in1({ dataBus[6] }),
  .out1({ S1453 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_251_ (
  .in1({ dataBus[7] }),
  .out1({ S1454 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_252_ (
  .in1({ dataBus[8] }),
  .out1({ S1455 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_253_ (
  .in1({ dataBus[9] }),
  .out1({ S1456 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_254_ (
  .in1({ dataBus[10] }),
  .out1({ S1457 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_255_ (
  .in1({ dataBus[11] }),
  .out1({ S1458 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_256_ (
  .in1({ dataBus[12] }),
  .out1({ S1459 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_257_ (
  .in1({ dataBus[13] }),
  .out1({ S1460 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_258_ (
  .in1({ dataBus[14] }),
  .out1({ S1461 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_259_ (
  .in1({ dataBus[15] }),
  .out1({ S1462 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_564_ (
  .in1({ S1446, S1445 }),
  .out1({ S1463 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_687_ (
  .in1({ S1, dataBus[0] }),
  .out1({ S1464 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_565_ (
  .in1({ S2, dataBus[0] }),
  .out1({ S1465 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_566_ (
  .in1({ S1465, S1463 }),
  .out1({ DP_INC2_out_0 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_567_ (
  .in1({ S1448, S1447 }),
  .out1({ S1466 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_688_ (
  .in1({ S9, dataBus[1] }),
  .out1({ S1467 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_568_ (
  .in1({ S10, dataBus[1] }),
  .out1({ S1468 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_260_ (
  .in1({ S1468 }),
  .out1({ S1469 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_569_ (
  .in1({ S1468, S1466 }),
  .out1({ S1470 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_689_ (
  .in1({ S1469, S1467 }),
  .out1({ S1471 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_570_ (
  .in1({ S1471, S1464 }),
  .out1({ S1472 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_690_ (
  .in1({ S1470, S1463 }),
  .out1({ S1473 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_571_ (
  .in1({ S1470, S1463 }),
  .out1({ S1474 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_572_ (
  .in1({ S1474, S1472 }),
  .out1({ DP_INC2_out_1 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_573_ (
  .in1({ S1472, S1466 }),
  .out1({ S1475 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_691_ (
  .in1({ S1473, S1467 }),
  .out1({ S1476 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_574_ (
  .in1({ S1475, S1449 }),
  .out1({ S1477 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_692_ (
  .in1({ S1476, dataBus[2] }),
  .out1({ S1478 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_575_ (
  .in1({ S1476, dataBus[2] }),
  .out1({ S1479 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_576_ (
  .in1({ S1479, S1477 }),
  .out1({ DP_INC2_out_2 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_577_ (
  .in1({ S1478, S1450 }),
  .out1({ S1480 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_693_ (
  .in1({ S1477, dataBus[3] }),
  .out1({ S1481 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_578_ (
  .in1({ S1477, dataBus[3] }),
  .out1({ S1482 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_579_ (
  .in1({ S1482, S1480 }),
  .out1({ DP_INC2_out_3 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_580_ (
  .in1({ S1481, S1451 }),
  .out1({ S1483 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_694_ (
  .in1({ S1480, dataBus[4] }),
  .out1({ S1484 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_581_ (
  .in1({ S1480, dataBus[4] }),
  .out1({ S1485 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_582_ (
  .in1({ S1485, S1483 }),
  .out1({ DP_INC2_out_4 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_583_ (
  .in1({ S1484, S1452 }),
  .out1({ S1486 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_695_ (
  .in1({ S1483, dataBus[5] }),
  .out1({ S1487 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_584_ (
  .in1({ S1483, dataBus[5] }),
  .out1({ S1488 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_585_ (
  .in1({ S1488, S1486 }),
  .out1({ DP_INC2_out_5 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_586_ (
  .in1({ S1487, S1453 }),
  .out1({ S1489 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_696_ (
  .in1({ S1486, dataBus[6] }),
  .out1({ S1490 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_587_ (
  .in1({ S1486, dataBus[6] }),
  .out1({ S1491 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_588_ (
  .in1({ S1491, S1489 }),
  .out1({ DP_INC2_out_6 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_589_ (
  .in1({ S1490, S1454 }),
  .out1({ S1492 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_697_ (
  .in1({ S1489, dataBus[7] }),
  .out1({ S1493 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_590_ (
  .in1({ S1489, dataBus[7] }),
  .out1({ S1494 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_591_ (
  .in1({ S1494, S1492 }),
  .out1({ DP_INC2_out_7 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_592_ (
  .in1({ S1493, S1455 }),
  .out1({ S1495 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_698_ (
  .in1({ S1492, dataBus[8] }),
  .out1({ S1496 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_593_ (
  .in1({ S1492, dataBus[8] }),
  .out1({ S1497 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_594_ (
  .in1({ S1497, S1495 }),
  .out1({ DP_INC2_out_8 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_595_ (
  .in1({ S1496, S1456 }),
  .out1({ S1498 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_699_ (
  .in1({ S1495, dataBus[9] }),
  .out1({ S1499 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_596_ (
  .in1({ S1495, dataBus[9] }),
  .out1({ S1500 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_597_ (
  .in1({ S1500, S1498 }),
  .out1({ DP_INC2_out_9 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_598_ (
  .in1({ S1499, S1457 }),
  .out1({ S1428 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_700_ (
  .in1({ S1498, dataBus[10] }),
  .out1({ S1429 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_599_ (
  .in1({ S1498, dataBus[10] }),
  .out1({ S1430 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_600_ (
  .in1({ S1430, S1428 }),
  .out1({ DP_INC2_out_10 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_601_ (
  .in1({ S1429, S1458 }),
  .out1({ S1431 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_701_ (
  .in1({ S1428, dataBus[11] }),
  .out1({ S1432 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_602_ (
  .in1({ S1428, dataBus[11] }),
  .out1({ S1433 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_603_ (
  .in1({ S1433, S1431 }),
  .out1({ DP_INC2_out_11 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_604_ (
  .in1({ S1432, S1459 }),
  .out1({ S1434 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_702_ (
  .in1({ S1431, dataBus[12] }),
  .out1({ S1435 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_605_ (
  .in1({ S1431, dataBus[12] }),
  .out1({ S1436 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_606_ (
  .in1({ S1436, S1434 }),
  .out1({ DP_INC2_out_12 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_607_ (
  .in1({ S1435, S1460 }),
  .out1({ S1437 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_703_ (
  .in1({ S1434, dataBus[13] }),
  .out1({ S1438 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_608_ (
  .in1({ S1434, dataBus[13] }),
  .out1({ S1439 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_609_ (
  .in1({ S1439, S1437 }),
  .out1({ DP_INC2_out_13 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_610_ (
  .in1({ S1438, S1461 }),
  .out1({ S1440 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_704_ (
  .in1({ S1437, dataBus[14] }),
  .out1({ S1441 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_611_ (
  .in1({ S1437, dataBus[14] }),
  .out1({ S1442 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_612_ (
  .in1({ S1442, S1440 }),
  .out1({ DP_INC2_out_14 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_613_ (
  .in1({ S1440, dataBus[15] }),
  .out1({ S1443 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_614_ (
  .in1({ S1441, S1462 }),
  .out1({ S1444 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_615_ (
  .in1({ S1444, S1443 }),
  .out1({ DP_INC2_out_15 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_261_ (
  .in1({ CU_ldIR }),
  .out1({ S1518 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_616_ (
  .in1({ CU_ldIR, S11 }),
  .out1({ S1519 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_705_ (
  .in1({ S1519, CU_inst_0 }),
  .out1({ S1520 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_617_ (
  .in1({ S1518, S12 }),
  .out1({ S1521 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_706_ (
  .in1({ S1521, dataBus[0] }),
  .out1({ S1522 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_707_ (
  .in1({ S1522, S1520 }),
  .out1({ S1501 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_708_ (
  .in1({ S1519, CU_inst_1 }),
  .out1({ S1523 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_709_ (
  .in1({ S1521, dataBus[1] }),
  .out1({ S1524 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_710_ (
  .in1({ S1524, S1523 }),
  .out1({ S1502 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_711_ (
  .in1({ S1519, CU_inst_2 }),
  .out1({ S1525 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_712_ (
  .in1({ S1521, dataBus[2] }),
  .out1({ S1526 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_713_ (
  .in1({ S1526, S1525 }),
  .out1({ S1503 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_714_ (
  .in1({ S1519, CU_inst_3 }),
  .out1({ S1527 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_715_ (
  .in1({ S1521, dataBus[3] }),
  .out1({ S1528 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_716_ (
  .in1({ S1528, S1527 }),
  .out1({ S1504 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_717_ (
  .in1({ S1519, CU_inst_4 }),
  .out1({ S1529 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_718_ (
  .in1({ S1521, dataBus[4] }),
  .out1({ S1530 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_719_ (
  .in1({ S1530, S1529 }),
  .out1({ S1505 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_720_ (
  .in1({ S1519, CU_inst_5 }),
  .out1({ S1531 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_721_ (
  .in1({ S1521, dataBus[5] }),
  .out1({ S1532 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_722_ (
  .in1({ S1532, S1531 }),
  .out1({ S1506 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_723_ (
  .in1({ S1519, CU_inst_6 }),
  .out1({ S1533 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_724_ (
  .in1({ S1521, dataBus[6] }),
  .out1({ S1534 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_725_ (
  .in1({ S1534, S1533 }),
  .out1({ S1507 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_726_ (
  .in1({ S1519, CU_inst_7 }),
  .out1({ S1535 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_727_ (
  .in1({ S1521, dataBus[7] }),
  .out1({ S1536 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_728_ (
  .in1({ S1536, S1535 }),
  .out1({ S1508 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_729_ (
  .in1({ S1519, CU_inst_8 }),
  .out1({ S1537 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_730_ (
  .in1({ S1521, dataBus[8] }),
  .out1({ S1538 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_731_ (
  .in1({ S1538, S1537 }),
  .out1({ S1509 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_732_ (
  .in1({ S1519, CU_inst_9 }),
  .out1({ S1539 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_733_ (
  .in1({ S1521, dataBus[9] }),
  .out1({ S1540 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_734_ (
  .in1({ S1540, S1539 }),
  .out1({ S1510 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_735_ (
  .in1({ S1519, CU_inst_10 }),
  .out1({ S1541 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_736_ (
  .in1({ S1521, dataBus[10] }),
  .out1({ S1542 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_737_ (
  .in1({ S1542, S1541 }),
  .out1({ S1511 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_738_ (
  .in1({ S1519, CU_inst_11 }),
  .out1({ S1543 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_739_ (
  .in1({ S1521, dataBus[11] }),
  .out1({ S1544 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_740_ (
  .in1({ S1544, S1543 }),
  .out1({ S1512 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_741_ (
  .in1({ S1519, CU_inst_12 }),
  .out1({ S1545 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_742_ (
  .in1({ S1521, dataBus[12] }),
  .out1({ S1546 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_743_ (
  .in1({ S1546, S1545 }),
  .out1({ S1513 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_744_ (
  .in1({ S1519, CU_inst_13 }),
  .out1({ S1547 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_745_ (
  .in1({ S1521, dataBus[13] }),
  .out1({ S1548 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_746_ (
  .in1({ S1548, S1547 }),
  .out1({ S1514 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_747_ (
  .in1({ S1519, CU_inst_14 }),
  .out1({ S1549 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_748_ (
  .in1({ S1521, dataBus[14] }),
  .out1({ S1550 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_749_ (
  .in1({ S1550, S1549 }),
  .out1({ S1515 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_750_ (
  .in1({ S1519, CU_inst_15 }),
  .out1({ S1551 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_751_ (
  .in1({ S1521, dataBus[15] }),
  .out1({ S1517 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_752_ (
  .in1({ S1517, S1551 }),
  .out1({ S1516 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_35_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1501 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_0 }),
  .Si({ S3072 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_36_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1502 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_1 }),
  .Si({ S3071 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_37_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1503 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_2 }),
  .Si({ S3070 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_38_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1504 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_3 }),
  .Si({ S3069 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_39_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1505 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_4 }),
  .Si({ S3068 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_40_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1506 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_5 }),
  .Si({ S3067 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_41_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1507 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_6 }),
  .Si({ S3066 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_42_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1508 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_7 }),
  .Si({ S3065 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_43_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1509 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_8 }),
  .Si({ S3064 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_44_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1510 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_9 }),
  .Si({ S3063 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_45_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1511 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_10 }),
  .Si({ S3062 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_46_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1512 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_11 }),
  .Si({ S3061 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_47_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1513 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_12 }),
  .Si({ S3060 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_48_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1514 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_13 }),
  .Si({ S3059 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_49_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1515 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_14 }),
  .Si({ S3058 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_50_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1516 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_15 }),
  .Si({ S3093 }),
  .global_reset({ 1'b0 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_262_ (
  .in1({ DP_AC_dout_0 }),
  .out1({ S1991 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_263_ (
  .in1({ DP_LGU1_in1_1 }),
  .out1({ S2001 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_264_ (
  .in1({ DP_LGU1_in1_0 }),
  .out1({ S2012 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_265_ (
  .in1({ DP_AC_dout_5 }),
  .out1({ S2023 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_266_ (
  .in1({ DP_LGU1_in1_2 }),
  .out1({ S2033 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_267_ (
  .in1({ DP_AC_dout_11 }),
  .out1({ S2044 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_268_ (
  .in1({ DP_AC_dout_15 }),
  .out1({ S2054 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_269_ (
  .in1({ DP_LGU1_in1_3 }),
  .out1({ S2065 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_270_ (
  .in1({ CU_SHF_1 }),
  .out1({ S2075 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_271_ (
  .in1({ CU_SHF_0 }),
  .out1({ S2086 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_272_ (
  .in1({ CU_NOT }),
  .out1({ S2096 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_273_ (
  .in1({ CU_AND }),
  .out1({ S2105 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_274_ (
  .in1({ DP_LGU1_in1_4 }),
  .out1({ S2106 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_275_ (
  .in1({ DP_LGU1_in1_5 }),
  .out1({ S2107 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_276_ (
  .in1({ DP_LGU1_in1_6 }),
  .out1({ S2108 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_277_ (
  .in1({ DP_LGU1_in1_8 }),
  .out1({ S2109 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_278_ (
  .in1({ DP_LGU1_in1_9 }),
  .out1({ S2110 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_279_ (
  .in1({ DP_LGU1_in1_12 }),
  .out1({ S2111 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_280_ (
  .in1({ DP_LGU1_in1_13 }),
  .out1({ S2112 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_753_ (
  .in1({ DP_LGU1_in1_0, DP_AC_dout_0 }),
  .out1({ S2113 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_754_ (
  .in1({ S2113, CU_AND }),
  .out1({ S2114 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_618_ (
  .in1({ CU_SHF_1, DP_LGU1_in1_3 }),
  .out1({ S2115 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_281_ (
  .in1({ S2115 }),
  .out1({ S2116 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_755_ (
  .in1({ DP_AC_dout_2, S2012 }),
  .out1({ S2117 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_756_ (
  .in1({ DP_AC_dout_3, DP_LGU1_in1_0 }),
  .out1({ S2118 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_757_ (
  .in1({ S2118, S2117 }),
  .out1({ S2119 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_758_ (
  .in1({ DP_LGU1_in1_0, DP_AC_dout_1 }),
  .out1({ S2120 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_282_ (
  .in1({ S2120 }),
  .out1({ S2121 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_619_ (
  .in1({ DP_LGU1_in1_0, S1991 }),
  .out1({ S2122 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_759_ (
  .in1({ S2012, DP_AC_dout_0 }),
  .out1({ S2123 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_760_ (
  .in1({ S2119, DP_LGU1_in1_1 }),
  .out1({ S2124 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_620_ (
  .in1({ S2123, DP_LGU1_in1_1 }),
  .out1({ S2125 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_761_ (
  .in1({ S2122, S2001 }),
  .out1({ S2126 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_621_ (
  .in1({ S2122, S2121 }),
  .out1({ S2127 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_622_ (
  .in1({ S2127, DP_LGU1_in1_1 }),
  .out1({ S2128 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_623_ (
  .in1({ S2128, DP_LGU1_in1_2 }),
  .out1({ S2129 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_762_ (
  .in1({ S2129, S2124 }),
  .out1({ S2130 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_763_ (
  .in1({ DP_AC_dout_4, S2012 }),
  .out1({ S2131 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_764_ (
  .in1({ DP_AC_dout_5, DP_LGU1_in1_0 }),
  .out1({ S2132 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_765_ (
  .in1({ S2132, S2131 }),
  .out1({ S2133 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_766_ (
  .in1({ S2133, S2001 }),
  .out1({ S2134 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_767_ (
  .in1({ DP_AC_dout_6, S2012 }),
  .out1({ S2135 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_768_ (
  .in1({ DP_AC_dout_7, DP_LGU1_in1_0 }),
  .out1({ S2136 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_769_ (
  .in1({ S2136, S2135 }),
  .out1({ S2137 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_283_ (
  .in1({ S2137 }),
  .out1({ S2138 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_770_ (
  .in1({ S2137, DP_LGU1_in1_1 }),
  .out1({ S2139 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_771_ (
  .in1({ S2139, S2134 }),
  .out1({ S1552 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_284_ (
  .in1({ S1552 }),
  .out1({ S1553 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_772_ (
  .in1({ S1553, DP_LGU1_in1_2 }),
  .out1({ S1554 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_773_ (
  .in1({ S1554, S2130 }),
  .out1({ S1555 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_774_ (
  .in1({ S1555, S2115 }),
  .out1({ S1556 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_624_ (
  .in1({ CU_SHF_1, S2065 }),
  .out1({ S1557 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_775_ (
  .in1({ S2075, DP_LGU1_in1_3 }),
  .out1({ S1558 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_776_ (
  .in1({ DP_AC_dout_8, S2012 }),
  .out1({ S1559 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_777_ (
  .in1({ DP_AC_dout_9, DP_LGU1_in1_0 }),
  .out1({ S1560 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_778_ (
  .in1({ S1560, S1559 }),
  .out1({ S1561 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_779_ (
  .in1({ S1561, S2001 }),
  .out1({ S1562 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_780_ (
  .in1({ DP_AC_dout_10, S2012 }),
  .out1({ S1563 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_781_ (
  .in1({ DP_AC_dout_11, DP_LGU1_in1_0 }),
  .out1({ S1564 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_782_ (
  .in1({ S1564, S1563 }),
  .out1({ S1565 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_783_ (
  .in1({ S1565, DP_LGU1_in1_1 }),
  .out1({ S1566 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_784_ (
  .in1({ S1566, S1562 }),
  .out1({ S1567 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_285_ (
  .in1({ S1567 }),
  .out1({ S1568 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_785_ (
  .in1({ S1567, S2033 }),
  .out1({ S1569 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_786_ (
  .in1({ DP_AC_dout_12, S2012 }),
  .out1({ S1570 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_787_ (
  .in1({ DP_AC_dout_13, DP_LGU1_in1_0 }),
  .out1({ S1571 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_788_ (
  .in1({ S1571, S1570 }),
  .out1({ S1572 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_789_ (
  .in1({ S1572, S2001 }),
  .out1({ S1573 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_790_ (
  .in1({ DP_AC_dout_14, S2012 }),
  .out1({ S1574 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_791_ (
  .in1({ DP_AC_dout_15, DP_LGU1_in1_0 }),
  .out1({ S1575 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_792_ (
  .in1({ S1575, S1574 }),
  .out1({ S1576 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_286_ (
  .in1({ S1576 }),
  .out1({ S1577 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_793_ (
  .in1({ S1576, DP_LGU1_in1_1 }),
  .out1({ S1578 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_794_ (
  .in1({ S1578, S1573 }),
  .out1({ S1579 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_795_ (
  .in1({ S1579, DP_LGU1_in1_2 }),
  .out1({ S1580 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_796_ (
  .in1({ S1580, S1569 }),
  .out1({ S1581 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_625_ (
  .in1({ S1581, S1558 }),
  .out1({ S1582 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_797_ (
  .in1({ S2126, CU_SHF_1 }),
  .out1({ S1583 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_626_ (
  .in1({ S2075, S2033 }),
  .out1({ S1584 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_798_ (
  .in1({ CU_SHF_1, DP_LGU1_in1_2 }),
  .out1({ S1585 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_799_ (
  .in1({ CU_SHF_1, DP_LGU1_in1_3 }),
  .out1({ S1586 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_800_ (
  .in1({ S1586, S2096 }),
  .out1({ S1587 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_627_ (
  .in1({ S1587, S1584 }),
  .out1({ S1588 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_801_ (
  .in1({ S1588, S1583 }),
  .out1({ S1589 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_628_ (
  .in1({ S1589, S1582 }),
  .out1({ S1590 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_802_ (
  .in1({ S1590, S1556 }),
  .out1({ S1591 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_629_ (
  .in1({ S2096, DP_AC_dout_0 }),
  .out1({ S1592 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_630_ (
  .in1({ S1592, CU_AND }),
  .out1({ S1593 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_803_ (
  .in1({ S1593, S1591 }),
  .out1({ S1594 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_804_ (
  .in1({ S1594, S2114 }),
  .out1({ S1595 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_287_ (
  .in1({ S1595 }),
  .out1({ DP_LGU1_out_0 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_805_ (
  .in1({ DP_AC_dout_9, S2012 }),
  .out1({ S1596 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_806_ (
  .in1({ DP_AC_dout_10, DP_LGU1_in1_0 }),
  .out1({ S1597 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_288_ (
  .in1({ S1597 }),
  .out1({ S1598 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_807_ (
  .in1({ S1597, S1596 }),
  .out1({ S1599 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_631_ (
  .in1({ S2044, DP_LGU1_in1_0 }),
  .out1({ S1600 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_808_ (
  .in1({ DP_AC_dout_11, S2012 }),
  .out1({ S1601 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_809_ (
  .in1({ DP_AC_dout_12, DP_LGU1_in1_0 }),
  .out1({ S1602 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_289_ (
  .in1({ S1602 }),
  .out1({ S1603 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_632_ (
  .in1({ S1603, S1600 }),
  .out1({ S1604 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_810_ (
  .in1({ S1602, S1601 }),
  .out1({ S1605 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_633_ (
  .in1({ S1605, S2001 }),
  .out1({ S1606 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_811_ (
  .in1({ S1604, DP_LGU1_in1_1 }),
  .out1({ S1607 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_634_ (
  .in1({ S1599, DP_LGU1_in1_1 }),
  .out1({ S1608 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_290_ (
  .in1({ S1608 }),
  .out1({ S1609 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_812_ (
  .in1({ S1609, S1607 }),
  .out1({ S1610 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_635_ (
  .in1({ S1608, S1606 }),
  .out1({ S1611 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_813_ (
  .in1({ S1611, S2033 }),
  .out1({ S1612 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_814_ (
  .in1({ S1612, DP_LGU1_in1_3 }),
  .out1({ S1613 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_815_ (
  .in1({ DP_AC_dout_13, S2012 }),
  .out1({ S1614 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_816_ (
  .in1({ DP_AC_dout_14, DP_LGU1_in1_0 }),
  .out1({ S1615 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_817_ (
  .in1({ S1615, S1614 }),
  .out1({ S1616 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_818_ (
  .in1({ S1616, S2001 }),
  .out1({ S1617 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_819_ (
  .in1({ DP_AC_dout_15, S2012 }),
  .out1({ S1618 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_291_ (
  .in1({ S1618 }),
  .out1({ S1619 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_820_ (
  .in1({ S1619, DP_LGU1_in1_1 }),
  .out1({ S1620 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_821_ (
  .in1({ S1620, S1617 }),
  .out1({ S1621 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_292_ (
  .in1({ S1621 }),
  .out1({ S1622 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_636_ (
  .in1({ S1622, S2033 }),
  .out1({ S1623 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_822_ (
  .in1({ S1621, DP_LGU1_in1_2 }),
  .out1({ S1624 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_823_ (
  .in1({ DP_AC_dout_15, DP_LGU1_in1_1 }),
  .out1({ S1625 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_824_ (
  .in1({ S1625, S1617 }),
  .out1({ S1626 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_825_ (
  .in1({ S1626, DP_LGU1_in1_2 }),
  .out1({ S1627 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_826_ (
  .in1({ S1623, CU_SHF_0 }),
  .out1({ S1628 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_637_ (
  .in1({ S1627, CU_SHF_0 }),
  .out1({ S1629 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_638_ (
  .in1({ S1629, S1613 }),
  .out1({ S1630 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_827_ (
  .in1({ S1630, S1628 }),
  .out1({ S1631 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_639_ (
  .in1({ S2023, DP_LGU1_in1_0 }),
  .out1({ S1632 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_828_ (
  .in1({ DP_AC_dout_5, S2012 }),
  .out1({ S1633 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_829_ (
  .in1({ DP_AC_dout_6, DP_LGU1_in1_0 }),
  .out1({ S1634 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_293_ (
  .in1({ S1634 }),
  .out1({ S1635 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_640_ (
  .in1({ S1635, S1632 }),
  .out1({ S1636 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_641_ (
  .in1({ S1636, DP_LGU1_in1_1 }),
  .out1({ S1637 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_830_ (
  .in1({ DP_AC_dout_7, S2012 }),
  .out1({ S1638 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_831_ (
  .in1({ DP_AC_dout_8, DP_LGU1_in1_0 }),
  .out1({ S1639 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_832_ (
  .in1({ S1639, S1638 }),
  .out1({ S1640 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_833_ (
  .in1({ S1640, DP_LGU1_in1_1 }),
  .out1({ S1641 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_294_ (
  .in1({ S1641 }),
  .out1({ S1642 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_642_ (
  .in1({ S1642, S1637 }),
  .out1({ S1643 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_643_ (
  .in1({ S1643, S2033 }),
  .out1({ S1644 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_834_ (
  .in1({ S2012, DP_AC_dout_1 }),
  .out1({ S1645 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_835_ (
  .in1({ DP_AC_dout_2, DP_LGU1_in1_0 }),
  .out1({ S1646 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_836_ (
  .in1({ S1646, S1645 }),
  .out1({ S1647 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_837_ (
  .in1({ S1647, S2001 }),
  .out1({ S1648 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_838_ (
  .in1({ DP_AC_dout_3, S2012 }),
  .out1({ S1649 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_839_ (
  .in1({ DP_AC_dout_4, DP_LGU1_in1_0 }),
  .out1({ S1650 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_840_ (
  .in1({ S1650, S1649 }),
  .out1({ S1651 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_841_ (
  .in1({ S1651, DP_LGU1_in1_1 }),
  .out1({ S1652 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_842_ (
  .in1({ S1652, S1648 }),
  .out1({ S1653 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_843_ (
  .in1({ S1653, S2033 }),
  .out1({ S1654 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_844_ (
  .in1({ S1654, S2115 }),
  .out1({ S1655 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_644_ (
  .in1({ S1655, S1644 }),
  .out1({ S1656 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_845_ (
  .in1({ S1645, S2113 }),
  .out1({ S1657 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_295_ (
  .in1({ S1657 }),
  .out1({ S1658 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_645_ (
  .in1({ S1658, DP_LGU1_in1_1 }),
  .out1({ S1659 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_846_ (
  .in1({ S1657, S2001 }),
  .out1({ S1660 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_646_ (
  .in1({ DP_LGU1_in1_3, DP_LGU1_in1_2 }),
  .out1({ S1661 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_296_ (
  .in1({ S1661 }),
  .out1({ S1662 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_847_ (
  .in1({ S1661, S1659 }),
  .out1({ S1663 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_848_ (
  .in1({ S1663, CU_SHF_1 }),
  .out1({ S1664 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_297_ (
  .in1({ S1664 }),
  .out1({ S1665 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_647_ (
  .in1({ S1665, S1656 }),
  .out1({ S1666 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_849_ (
  .in1({ S1666, S1631 }),
  .out1({ S1667 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_850_ (
  .in1({ S1667, S2096 }),
  .out1({ S1668 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_851_ (
  .in1({ CU_NOT, DP_AC_dout_1 }),
  .out1({ S1669 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_298_ (
  .in1({ S1669 }),
  .out1({ S1670 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_648_ (
  .in1({ S1670, CU_AND }),
  .out1({ S1671 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_852_ (
  .in1({ S1671, S1668 }),
  .out1({ S1672 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_649_ (
  .in1({ S2105, S2001 }),
  .out1({ S1673 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_853_ (
  .in1({ S1673, DP_AC_dout_1 }),
  .out1({ S1674 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_854_ (
  .in1({ S1674, S1672 }),
  .out1({ DP_LGU1_out_1 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_855_ (
  .in1({ S2119, S2001 }),
  .out1({ S1675 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_856_ (
  .in1({ S2133, DP_LGU1_in1_1 }),
  .out1({ S1676 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_857_ (
  .in1({ S1676, S1675 }),
  .out1({ S1677 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_650_ (
  .in1({ S2138, DP_LGU1_in1_1 }),
  .out1({ S1678 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_858_ (
  .in1({ S1561, DP_LGU1_in1_1 }),
  .out1({ S1679 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_299_ (
  .in1({ S1679 }),
  .out1({ S1680 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_651_ (
  .in1({ S1680, S1678 }),
  .out1({ S1681 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_652_ (
  .in1({ S1677, DP_LGU1_in1_2 }),
  .out1({ S1682 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_859_ (
  .in1({ S1681, DP_LGU1_in1_2 }),
  .out1({ S1683 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_860_ (
  .in1({ S1683, S2075 }),
  .out1({ S1684 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_653_ (
  .in1({ S1684, S1682 }),
  .out1({ S1685 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_654_ (
  .in1({ S2075, DP_LGU1_in1_2 }),
  .out1({ S1686 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_861_ (
  .in1({ CU_SHF_1, S2033 }),
  .out1({ S1687 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_862_ (
  .in1({ S2120, S2117 }),
  .out1({ S1688 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_655_ (
  .in1({ S2122, S2001 }),
  .out1({ S1689 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_863_ (
  .in1({ S2123, DP_LGU1_in1_1 }),
  .out1({ S1690 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_656_ (
  .in1({ S1688, DP_LGU1_in1_1 }),
  .out1({ S1691 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_300_ (
  .in1({ S1691 }),
  .out1({ S1692 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_864_ (
  .in1({ S1692, S1690 }),
  .out1({ S1693 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_657_ (
  .in1({ S1691, S1689 }),
  .out1({ S1694 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_865_ (
  .in1({ S1694, S1686 }),
  .out1({ S1695 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_866_ (
  .in1({ S1695, S1558 }),
  .out1({ S1696 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_658_ (
  .in1({ S1696, S1685 }),
  .out1({ S1697 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_659_ (
  .in1({ CU_SHF_0, CU_SHF_1 }),
  .out1({ S1698 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_867_ (
  .in1({ S2086, S2075 }),
  .out1({ S1699 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_868_ (
  .in1({ S1565, S2001 }),
  .out1({ S1700 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_869_ (
  .in1({ S1572, DP_LGU1_in1_1 }),
  .out1({ S1701 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_870_ (
  .in1({ S1701, S1700 }),
  .out1({ S1702 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_871_ (
  .in1({ S1702, S2033 }),
  .out1({ S1703 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_660_ (
  .in1({ S1577, DP_LGU1_in1_1 }),
  .out1({ S1704 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_872_ (
  .in1({ S1576, S2001 }),
  .out1({ S1705 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_873_ (
  .in1({ S1705, S1625 }),
  .out1({ S1706 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_874_ (
  .in1({ S1706, DP_LGU1_in1_2 }),
  .out1({ S1707 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_875_ (
  .in1({ S1707, S1703 }),
  .out1({ S1708 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_876_ (
  .in1({ S1708, S1698 }),
  .out1({ S1709 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_661_ (
  .in1({ S2086, CU_SHF_1 }),
  .out1({ S1710 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_877_ (
  .in1({ CU_SHF_0, S2075 }),
  .out1({ S1711 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_878_ (
  .in1({ S1704, DP_LGU1_in1_2 }),
  .out1({ S1712 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_879_ (
  .in1({ S1712, S1703 }),
  .out1({ S1713 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_301_ (
  .in1({ S1713 }),
  .out1({ S1714 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_662_ (
  .in1({ S1714, S1711 }),
  .out1({ S1715 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_880_ (
  .in1({ S1713, S1710 }),
  .out1({ S1716 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_881_ (
  .in1({ S1709, DP_LGU1_in1_3 }),
  .out1({ S1717 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_663_ (
  .in1({ S1717, S1715 }),
  .out1({ S1718 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_664_ (
  .in1({ S1718, S1697 }),
  .out1({ S1719 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_665_ (
  .in1({ S1719, CU_NOT }),
  .out1({ S1720 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_882_ (
  .in1({ CU_NOT, DP_AC_dout_2 }),
  .out1({ S1721 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_883_ (
  .in1({ S1721, S2105 }),
  .out1({ S1722 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_666_ (
  .in1({ S1722, S1720 }),
  .out1({ S1723 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_884_ (
  .in1({ DP_LGU1_in1_2, DP_AC_dout_2 }),
  .out1({ S1724 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_667_ (
  .in1({ S1724, S2105 }),
  .out1({ S1725 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_668_ (
  .in1({ S1725, S1723 }),
  .out1({ S1726 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_302_ (
  .in1({ S1726 }),
  .out1({ DP_LGU1_out_2 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_669_ (
  .in1({ S1604, DP_LGU1_in1_1 }),
  .out1({ S1727 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_885_ (
  .in1({ S1605, S2001 }),
  .out1({ S1728 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_886_ (
  .in1({ S1616, DP_LGU1_in1_1 }),
  .out1({ S1729 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_303_ (
  .in1({ S1729 }),
  .out1({ S1730 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_670_ (
  .in1({ S1730, S1727 }),
  .out1({ S1731 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_887_ (
  .in1({ S1729, S1728 }),
  .out1({ S1732 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_671_ (
  .in1({ S1731, DP_LGU1_in1_2 }),
  .out1({ S1733 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_888_ (
  .in1({ S1732, S2033 }),
  .out1({ S1734 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_672_ (
  .in1({ S1618, DP_LGU1_in1_1 }),
  .out1({ S1735 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_889_ (
  .in1({ S1735, DP_LGU1_in1_2 }),
  .out1({ S1736 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_304_ (
  .in1({ S1736 }),
  .out1({ S1737 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_673_ (
  .in1({ S1737, S1733 }),
  .out1({ S1738 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_674_ (
  .in1({ S1738, S1711 }),
  .out1({ S1739 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_890_ (
  .in1({ DP_AC_dout_15, DP_LGU1_in1_2 }),
  .out1({ S1740 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_891_ (
  .in1({ S1740, S1734 }),
  .out1({ S1741 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_892_ (
  .in1({ S1741, S1698 }),
  .out1({ S1742 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_893_ (
  .in1({ S1742, DP_LGU1_in1_3 }),
  .out1({ S1743 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_675_ (
  .in1({ S1743, S1739 }),
  .out1({ S1744 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_894_ (
  .in1({ S1640, S2001 }),
  .out1({ S1745 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_895_ (
  .in1({ S1599, DP_LGU1_in1_1 }),
  .out1({ S1746 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_896_ (
  .in1({ S1746, S1745 }),
  .out1({ S1747 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_676_ (
  .in1({ S1747, S2033 }),
  .out1({ S1748 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_897_ (
  .in1({ S1651, S2001 }),
  .out1({ S1749 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_677_ (
  .in1({ S1636, S2001 }),
  .out1({ S1750 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_678_ (
  .in1({ S1750, DP_LGU1_in1_2 }),
  .out1({ S1751 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_898_ (
  .in1({ S1751, S1749 }),
  .out1({ S1752 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_899_ (
  .in1({ S1752, S2075 }),
  .out1({ S1753 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_679_ (
  .in1({ S1753, S1748 }),
  .out1({ S1754 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_900_ (
  .in1({ S1649, S1646 }),
  .out1({ S1755 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_901_ (
  .in1({ S1755, S2001 }),
  .out1({ S1756 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_902_ (
  .in1({ S1657, DP_LGU1_in1_1 }),
  .out1({ S1757 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_903_ (
  .in1({ S1757, S1756 }),
  .out1({ S1758 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_305_ (
  .in1({ S1758 }),
  .out1({ S1759 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_904_ (
  .in1({ S1758, S1686 }),
  .out1({ S1760 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_905_ (
  .in1({ S1760, S1558 }),
  .out1({ S1761 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_680_ (
  .in1({ S1761, S1754 }),
  .out1({ S1762 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_681_ (
  .in1({ S1762, S1744 }),
  .out1({ S1763 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_682_ (
  .in1({ S1763, CU_NOT }),
  .out1({ S1764 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_906_ (
  .in1({ CU_NOT, DP_AC_dout_3 }),
  .out1({ S1765 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_907_ (
  .in1({ S1765, S2105 }),
  .out1({ S1766 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_683_ (
  .in1({ S1766, S1764 }),
  .out1({ S1767 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_908_ (
  .in1({ DP_LGU1_in1_3, DP_AC_dout_3 }),
  .out1({ S1768 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_684_ (
  .in1({ S1768, S2105 }),
  .out1({ S1769 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_685_ (
  .in1({ S1769, S1767 }),
  .out1({ S1770 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_306_ (
  .in1({ S1770 }),
  .out1({ DP_LGU1_out_3 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_909_ (
  .in1({ S1579, S2033 }),
  .out1({ S1771 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_686_ (
  .in1({ S1740, CU_SHF_0 }),
  .out1({ S1772 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_307_ (
  .in1({ S1772 }),
  .out1({ S1773 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_910_ (
  .in1({ S1773, S1771 }),
  .out1({ S1774 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_911_ (
  .in1({ S1774, S1557 }),
  .out1({ S1775 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_912_ (
  .in1({ S1775, S2096 }),
  .out1({ S1776 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_913_ (
  .in1({ S2131, S2118 }),
  .out1({ S1777 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_914_ (
  .in1({ S1777, S2001 }),
  .out1({ S1778 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_915_ (
  .in1({ S1688, DP_LGU1_in1_1 }),
  .out1({ S1779 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_916_ (
  .in1({ S1779, S1778 }),
  .out1({ S1780 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_687_ (
  .in1({ S2125, S2033 }),
  .out1({ S1781 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_917_ (
  .in1({ S2126, DP_LGU1_in1_2 }),
  .out1({ S1782 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_688_ (
  .in1({ S1780, DP_LGU1_in1_2 }),
  .out1({ S1783 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_308_ (
  .in1({ S1783 }),
  .out1({ S1784 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_918_ (
  .in1({ S1784, S1782 }),
  .out1({ S1785 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_689_ (
  .in1({ S1783, S1781 }),
  .out1({ S1786 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_690_ (
  .in1({ S2075, DP_LGU1_in1_3 }),
  .out1({ S1787 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_919_ (
  .in1({ S1787, S1786 }),
  .out1({ S1788 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_920_ (
  .in1({ S1568, DP_LGU1_in1_2 }),
  .out1({ S1789 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_691_ (
  .in1({ S1552, DP_LGU1_in1_2 }),
  .out1({ S1790 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_692_ (
  .in1({ S1790, S2116 }),
  .out1({ S1791 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_921_ (
  .in1({ S1791, S1789 }),
  .out1({ S1792 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_922_ (
  .in1({ S1792, S1788 }),
  .out1({ S1793 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_923_ (
  .in1({ S1771, S1740 }),
  .out1({ S1794 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_693_ (
  .in1({ S1793, S1776 }),
  .out1({ S1795 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_924_ (
  .in1({ CU_NOT, DP_AC_dout_4 }),
  .out1({ S1796 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_925_ (
  .in1({ S1796, S2105 }),
  .out1({ S1797 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_694_ (
  .in1({ S1797, S1795 }),
  .out1({ S1798 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_926_ (
  .in1({ CU_AND, DP_AC_dout_4 }),
  .out1({ S1799 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_695_ (
  .in1({ S1799, S2106 }),
  .out1({ S1800 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_696_ (
  .in1({ S1800, S1798 }),
  .out1({ S1801 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_309_ (
  .in1({ S1801 }),
  .out1({ DP_LGU1_out_4 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_927_ (
  .in1({ CU_AND, DP_AC_dout_5 }),
  .out1({ S1802 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_697_ (
  .in1({ S1802, S2107 }),
  .out1({ S1803 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_698_ (
  .in1({ S1711, DP_LGU1_in1_2 }),
  .out1({ S1804 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_310_ (
  .in1({ S1804 }),
  .out1({ S1805 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_928_ (
  .in1({ S1804, S1621 }),
  .out1({ S1806 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_929_ (
  .in1({ S1626, S2033 }),
  .out1({ S1807 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_930_ (
  .in1({ S1807, S1740 }),
  .out1({ S1808 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_931_ (
  .in1({ S1808, S1698 }),
  .out1({ S1809 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_932_ (
  .in1({ S1809, S1806 }),
  .out1({ S1810 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_699_ (
  .in1({ S1810, S2065 }),
  .out1({ S1811 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_933_ (
  .in1({ S1610, DP_LGU1_in1_2 }),
  .out1({ S1812 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_934_ (
  .in1({ S1643, S2033 }),
  .out1({ S1813 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_935_ (
  .in1({ S1813, S1812 }),
  .out1({ S1814 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_700_ (
  .in1({ S1814, CU_SHF_1 }),
  .out1({ S1815 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_936_ (
  .in1({ S1650, S1633 }),
  .out1({ S1816 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_311_ (
  .in1({ S1816 }),
  .out1({ S1817 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_701_ (
  .in1({ S1817, DP_LGU1_in1_1 }),
  .out1({ S1818 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_937_ (
  .in1({ S1755, DP_LGU1_in1_1 }),
  .out1({ S1819 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_312_ (
  .in1({ S1819 }),
  .out1({ S1820 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_702_ (
  .in1({ S1820, S1818 }),
  .out1({ S1821 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_313_ (
  .in1({ S1821 }),
  .out1({ S1822 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_703_ (
  .in1({ S1821, S1687 }),
  .out1({ S1823 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_938_ (
  .in1({ S1822, S1686 }),
  .out1({ S1824 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_704_ (
  .in1({ S1660, S1585 }),
  .out1({ S1825 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_939_ (
  .in1({ S1659, S1584 }),
  .out1({ S1826 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_705_ (
  .in1({ S1825, S1823 }),
  .out1({ S1827 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_940_ (
  .in1({ S1826, S1824 }),
  .out1({ S1828 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_941_ (
  .in1({ S1827, S1558 }),
  .out1({ S1829 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_706_ (
  .in1({ S1829, S1815 }),
  .out1({ S1830 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_707_ (
  .in1({ S1830, S1811 }),
  .out1({ S1831 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_708_ (
  .in1({ S1831, CU_NOT }),
  .out1({ S1832 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_942_ (
  .in1({ CU_NOT, DP_AC_dout_5 }),
  .out1({ S1833 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_943_ (
  .in1({ S1833, S2105 }),
  .out1({ S1834 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_709_ (
  .in1({ S1834, S1832 }),
  .out1({ S1835 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_710_ (
  .in1({ S1835, S1803 }),
  .out1({ S1836 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_314_ (
  .in1({ S1836 }),
  .out1({ DP_LGU1_out_5 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_944_ (
  .in1({ CU_AND, DP_AC_dout_6 }),
  .out1({ S1837 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_711_ (
  .in1({ S1837, S2108 }),
  .out1({ S1838 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_712_ (
  .in1({ S1805, S1705 }),
  .out1({ S1839 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_945_ (
  .in1({ S1804, S1704 }),
  .out1({ S1840 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_946_ (
  .in1({ S1706, S2033 }),
  .out1({ S1841 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_947_ (
  .in1({ S1841, S1740 }),
  .out1({ S1842 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_948_ (
  .in1({ S1842, S1698 }),
  .out1({ S1843 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_315_ (
  .in1({ S1843 }),
  .out1({ S1844 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_713_ (
  .in1({ S1844, S1839 }),
  .out1({ S1845 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_949_ (
  .in1({ S1843, S1840 }),
  .out1({ S1846 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_714_ (
  .in1({ S1846, S2065 }),
  .out1({ S1847 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_715_ (
  .in1({ S1681, DP_LGU1_in1_2 }),
  .out1({ S1848 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_950_ (
  .in1({ S1702, DP_LGU1_in1_2 }),
  .out1({ S1849 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_316_ (
  .in1({ S1849 }),
  .out1({ S1850 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_716_ (
  .in1({ S1850, S1848 }),
  .out1({ S1851 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_717_ (
  .in1({ S1851, CU_SHF_1 }),
  .out1({ S1852 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_951_ (
  .in1({ S2135, S2132 }),
  .out1({ S1853 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_317_ (
  .in1({ S1853 }),
  .out1({ S1854 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_718_ (
  .in1({ S1854, DP_LGU1_in1_1 }),
  .out1({ S1855 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_952_ (
  .in1({ S1777, DP_LGU1_in1_1 }),
  .out1({ S1856 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_318_ (
  .in1({ S1856 }),
  .out1({ S1857 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_719_ (
  .in1({ S1857, S1855 }),
  .out1({ S1858 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_720_ (
  .in1({ S1858, S1687 }),
  .out1({ S1859 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_721_ (
  .in1({ S1693, S1585 }),
  .out1({ S1860 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_722_ (
  .in1({ S1860, S1859 }),
  .out1({ S1861 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_953_ (
  .in1({ S1861, S1558 }),
  .out1({ S1862 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_723_ (
  .in1({ S1862, S1852 }),
  .out1({ S1863 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_724_ (
  .in1({ S1863, S1847 }),
  .out1({ S1864 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_725_ (
  .in1({ S1864, CU_NOT }),
  .out1({ S1865 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_954_ (
  .in1({ CU_NOT, DP_AC_dout_6 }),
  .out1({ S1866 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_955_ (
  .in1({ S1866, S2105 }),
  .out1({ S1867 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_726_ (
  .in1({ S1867, S1865 }),
  .out1({ S1868 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_727_ (
  .in1({ S1868, S1838 }),
  .out1({ S1869 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_319_ (
  .in1({ S1869 }),
  .out1({ DP_LGU1_out_6 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_956_ (
  .in1({ CU_AND, DP_AC_dout_7 }),
  .out1({ S1870 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_320_ (
  .in1({ S1870 }),
  .out1({ S1871 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_957_ (
  .in1({ S1871, DP_LGU1_in1_7 }),
  .out1({ S1872 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_728_ (
  .in1({ S1732, S2033 }),
  .out1({ S1873 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_729_ (
  .in1({ S1747, DP_LGU1_in1_2 }),
  .out1({ S1874 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_730_ (
  .in1({ S1874, S1873 }),
  .out1({ S1875 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_958_ (
  .in1({ S1875, S2075 }),
  .out1({ S1876 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_959_ (
  .in1({ S1638, S1634 }),
  .out1({ S1877 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_321_ (
  .in1({ S1877 }),
  .out1({ S1878 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_731_ (
  .in1({ S1878, DP_LGU1_in1_1 }),
  .out1({ S1879 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_960_ (
  .in1({ S1877, S2001 }),
  .out1({ S1880 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_961_ (
  .in1({ S1816, DP_LGU1_in1_1 }),
  .out1({ S1881 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_322_ (
  .in1({ S1881 }),
  .out1({ S1882 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_732_ (
  .in1({ S1882, S1879 }),
  .out1({ S1883 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_962_ (
  .in1({ S1881, S1880 }),
  .out1({ S1884 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_733_ (
  .in1({ S1883, S1687 }),
  .out1({ S1885 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_963_ (
  .in1({ S1884, S1686 }),
  .out1({ S1886 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_734_ (
  .in1({ S1759, S1585 }),
  .out1({ S1887 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_964_ (
  .in1({ S1758, S1584 }),
  .out1({ S1888 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_735_ (
  .in1({ S1887, S1885 }),
  .out1({ S1889 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_965_ (
  .in1({ S1888, S1886 }),
  .out1({ S1890 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_736_ (
  .in1({ S1890, DP_LGU1_in1_3 }),
  .out1({ S1891 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_966_ (
  .in1({ S1891, S1876 }),
  .out1({ S1892 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_967_ (
  .in1({ S1804, S1735 }),
  .out1({ S1893 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_323_ (
  .in1({ S1893 }),
  .out1({ S1894 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_737_ (
  .in1({ S1699, S2054 }),
  .out1({ S1895 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_968_ (
  .in1({ S1698, DP_AC_dout_15 }),
  .out1({ S1896 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_738_ (
  .in1({ S1895, S1894 }),
  .out1({ S1897 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_969_ (
  .in1({ S1897, DP_LGU1_in1_3 }),
  .out1({ S1898 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_970_ (
  .in1({ S1898, S1892 }),
  .out1({ S1899 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_971_ (
  .in1({ S1899, S2096 }),
  .out1({ S1900 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_972_ (
  .in1({ CU_NOT, DP_AC_dout_7 }),
  .out1({ S1901 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_324_ (
  .in1({ S1901 }),
  .out1({ S1902 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_739_ (
  .in1({ S1902, CU_AND }),
  .out1({ S1903 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_973_ (
  .in1({ S1903, S1900 }),
  .out1({ S1904 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_974_ (
  .in1({ S1904, S1872 }),
  .out1({ DP_LGU1_out_7 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_740_ (
  .in1({ DP_LGU1_in1_3, S2033 }),
  .out1({ S1905 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_741_ (
  .in1({ S1687, S2126 }),
  .out1({ S1906 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_742_ (
  .in1({ S1906, S1787 }),
  .out1({ S1907 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_975_ (
  .in1({ S1559, S2136 }),
  .out1({ S1908 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_976_ (
  .in1({ S1908, S2001 }),
  .out1({ S1909 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_977_ (
  .in1({ S1853, DP_LGU1_in1_1 }),
  .out1({ S1910 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_978_ (
  .in1({ S1910, S1909 }),
  .out1({ S1911 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_979_ (
  .in1({ S1911, S2033 }),
  .out1({ S1912 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_980_ (
  .in1({ S1780, DP_LGU1_in1_2 }),
  .out1({ S1913 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_981_ (
  .in1({ S1913, S1912 }),
  .out1({ S1914 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_743_ (
  .in1({ S1914, DP_LGU1_in1_3 }),
  .out1({ S1915 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_744_ (
  .in1({ S1915, S1907 }),
  .out1({ S1916 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_982_ (
  .in1({ S1581, S2115 }),
  .out1({ S1917 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_745_ (
  .in1({ S1896, S2065 }),
  .out1({ S1918 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_746_ (
  .in1({ S1918, CU_NOT }),
  .out1({ S1919 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_325_ (
  .in1({ S1919 }),
  .out1({ S1920 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_983_ (
  .in1({ S1919, S1917 }),
  .out1({ S1921 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_747_ (
  .in1({ S1921, S1916 }),
  .out1({ S1922 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_984_ (
  .in1({ CU_NOT, DP_AC_dout_8 }),
  .out1({ S1923 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_985_ (
  .in1({ S1923, S2105 }),
  .out1({ S1924 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_748_ (
  .in1({ S1924, S1922 }),
  .out1({ S1925 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_986_ (
  .in1({ CU_AND, DP_AC_dout_8 }),
  .out1({ S1926 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_749_ (
  .in1({ S1926, S2109 }),
  .out1({ S1927 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_750_ (
  .in1({ S1927, S1925 }),
  .out1({ S1928 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_326_ (
  .in1({ S1928 }),
  .out1({ DP_LGU1_out_8 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_987_ (
  .in1({ CU_AND, DP_AC_dout_9 }),
  .out1({ S1929 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_751_ (
  .in1({ S1929, S2110 }),
  .out1({ S1930 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_988_ (
  .in1({ S1627, S1612 }),
  .out1({ S1931 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_752_ (
  .in1({ S1699, DP_LGU1_in1_3 }),
  .out1({ S1932 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_989_ (
  .in1({ S1932, S1931 }),
  .out1({ S1933 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_990_ (
  .in1({ S1933, S1919 }),
  .out1({ S1934 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_991_ (
  .in1({ S1905, S1821 }),
  .out1({ S1935 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_753_ (
  .in1({ S1687, S1660 }),
  .out1({ S1936 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_754_ (
  .in1({ S1936, S1787 }),
  .out1({ S1937 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_992_ (
  .in1({ S1639, S1596 }),
  .out1({ S1938 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_993_ (
  .in1({ S1938, S2001 }),
  .out1({ S1939 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_994_ (
  .in1({ S1877, DP_LGU1_in1_1 }),
  .out1({ S1940 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_995_ (
  .in1({ S1940, S1939 }),
  .out1({ S1941 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_755_ (
  .in1({ S1941, S1662 }),
  .out1({ S1942 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_756_ (
  .in1({ S1942, S1937 }),
  .out1({ S1943 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_996_ (
  .in1({ S1943, S1935 }),
  .out1({ S1944 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_997_ (
  .in1({ S1624, S1612 }),
  .out1({ S1945 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_757_ (
  .in1({ S2116, S2086 }),
  .out1({ S1946 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_998_ (
  .in1({ S2115, CU_SHF_0 }),
  .out1({ S1947 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_999_ (
  .in1({ S1946, S1945 }),
  .out1({ S1948 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1000_ (
  .in1({ S1948, S1944 }),
  .out1({ S1949 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_758_ (
  .in1({ S1949, S1934 }),
  .out1({ S1950 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1001_ (
  .in1({ CU_NOT, DP_AC_dout_9 }),
  .out1({ S1951 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1002_ (
  .in1({ S1951, S2105 }),
  .out1({ S1952 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_759_ (
  .in1({ S1952, S1950 }),
  .out1({ S1953 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_760_ (
  .in1({ S1953, S1930 }),
  .out1({ S1954 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_327_ (
  .in1({ S1954 }),
  .out1({ DP_LGU1_out_9 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1003_ (
  .in1({ S1695, DP_LGU1_in1_3 }),
  .out1({ S1955 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1004_ (
  .in1({ S1563, S1560 }),
  .out1({ S1956 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1005_ (
  .in1({ S1956, S2001 }),
  .out1({ S1957 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1006_ (
  .in1({ S1908, DP_LGU1_in1_1 }),
  .out1({ S1958 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1007_ (
  .in1({ S1958, S1957 }),
  .out1({ S1959 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1008_ (
  .in1({ S1959, S1686 }),
  .out1({ S1960 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_761_ (
  .in1({ S1858, S1585 }),
  .out1({ S1961 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1009_ (
  .in1({ S1960, S1586 }),
  .out1({ S1962 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_762_ (
  .in1({ S1962, S1961 }),
  .out1({ S1963 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1010_ (
  .in1({ S1963, S1716 }),
  .out1({ S1964 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1011_ (
  .in1({ S1964, S1955 }),
  .out1({ S1965 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_763_ (
  .in1({ S1709, DP_LGU1_in1_3 }),
  .out1({ S1966 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_764_ (
  .in1({ S1966, S1920 }),
  .out1({ S1967 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1012_ (
  .in1({ S1967, S1965 }),
  .out1({ S1968 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1013_ (
  .in1({ CU_NOT, DP_AC_dout_10 }),
  .out1({ S1969 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_328_ (
  .in1({ S1969 }),
  .out1({ S1970 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_765_ (
  .in1({ S1970, CU_AND }),
  .out1({ S1971 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1014_ (
  .in1({ S1971, S1968 }),
  .out1({ S1972 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1015_ (
  .in1({ CU_AND, DP_AC_dout_10 }),
  .out1({ S1973 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_329_ (
  .in1({ S1973 }),
  .out1({ S1974 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1016_ (
  .in1({ S1974, DP_LGU1_in1_10 }),
  .out1({ S1975 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1017_ (
  .in1({ S1975, S1972 }),
  .out1({ DP_LGU1_out_10 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1018_ (
  .in1({ S1760, DP_LGU1_in1_3 }),
  .out1({ S1976 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_766_ (
  .in1({ S1600, S1598 }),
  .out1({ S1977 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_767_ (
  .in1({ S1977, DP_LGU1_in1_1 }),
  .out1({ S1978 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1019_ (
  .in1({ S1938, DP_LGU1_in1_1 }),
  .out1({ S1979 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_330_ (
  .in1({ S1979 }),
  .out1({ S1980 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_768_ (
  .in1({ S1980, S1978 }),
  .out1({ S1981 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_769_ (
  .in1({ S1981, S1687 }),
  .out1({ S1982 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_770_ (
  .in1({ S1982, DP_LGU1_in1_3 }),
  .out1({ S1983 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1020_ (
  .in1({ S1983, S1742 }),
  .out1({ S1984 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1021_ (
  .in1({ S1984, S1558 }),
  .out1({ S1985 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_771_ (
  .in1({ S1883, S1585 }),
  .out1({ S1986 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_772_ (
  .in1({ S1986, S1739 }),
  .out1({ S1987 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1022_ (
  .in1({ S1987, S1985 }),
  .out1({ S1988 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1023_ (
  .in1({ S1988, S1976 }),
  .out1({ S1989 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1024_ (
  .in1({ S1989, S1919 }),
  .out1({ S1990 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1025_ (
  .in1({ CU_NOT, DP_AC_dout_11 }),
  .out1({ S1992 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_331_ (
  .in1({ S1992 }),
  .out1({ S1993 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_773_ (
  .in1({ S1993, CU_AND }),
  .out1({ S1994 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1026_ (
  .in1({ S1994, S1990 }),
  .out1({ S1995 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1027_ (
  .in1({ CU_AND, DP_AC_dout_11 }),
  .out1({ S1996 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_332_ (
  .in1({ S1996 }),
  .out1({ S1997 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1028_ (
  .in1({ S1997, DP_LGU1_in1_11 }),
  .out1({ S1998 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1029_ (
  .in1({ S1998, S1995 }),
  .out1({ DP_LGU1_out_11 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_774_ (
  .in1({ S1947, S1771 }),
  .out1({ S1999 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1030_ (
  .in1({ S1570, S1564 }),
  .out1({ S2000 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_333_ (
  .in1({ S2000 }),
  .out1({ S2002 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_775_ (
  .in1({ S1956, S2001 }),
  .out1({ S2003 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_776_ (
  .in1({ S2000, DP_LGU1_in1_1 }),
  .out1({ S2004 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_777_ (
  .in1({ S2004, S2003 }),
  .out1({ S2005 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1031_ (
  .in1({ S2005, S2033 }),
  .out1({ S2006 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1032_ (
  .in1({ S1911, DP_LGU1_in1_2 }),
  .out1({ S2007 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1033_ (
  .in1({ S2007, S2006 }),
  .out1({ S2008 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_778_ (
  .in1({ S2008, DP_LGU1_in1_3 }),
  .out1({ S2009 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1034_ (
  .in1({ S1785, DP_LGU1_in1_3 }),
  .out1({ S2010 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1035_ (
  .in1({ S2010, S1711 }),
  .out1({ S2011 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_779_ (
  .in1({ S2011, S2009 }),
  .out1({ S2013 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_780_ (
  .in1({ S2013, S1999 }),
  .out1({ S2014 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_781_ (
  .in1({ S2014, S1698 }),
  .out1({ S2015 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1036_ (
  .in1({ S1932, S1794 }),
  .out1({ S2016 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1037_ (
  .in1({ S2016, S1919 }),
  .out1({ S2017 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_782_ (
  .in1({ S2017, S2015 }),
  .out1({ S2018 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1038_ (
  .in1({ CU_NOT, DP_AC_dout_12 }),
  .out1({ S2019 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1039_ (
  .in1({ S2019, S2105 }),
  .out1({ S2020 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_783_ (
  .in1({ S2020, S2018 }),
  .out1({ S2021 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1040_ (
  .in1({ CU_AND, DP_AC_dout_12 }),
  .out1({ S2022 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_784_ (
  .in1({ S2022, S2111 }),
  .out1({ S2024 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_785_ (
  .in1({ S2024, S2021 }),
  .out1({ S2025 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_334_ (
  .in1({ S2025 }),
  .out1({ DP_LGU1_out_12 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1041_ (
  .in1({ S1941, S1584 }),
  .out1({ S2026 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1042_ (
  .in1({ S1614, S1602 }),
  .out1({ S2027 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_786_ (
  .in1({ S2027, DP_LGU1_in1_1 }),
  .out1({ S2028 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1043_ (
  .in1({ S1977, DP_LGU1_in1_1 }),
  .out1({ S2029 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_787_ (
  .in1({ S2028, S1687 }),
  .out1({ S2030 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1044_ (
  .in1({ S2030, S2029 }),
  .out1({ S2031 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1045_ (
  .in1({ S2031, S2026 }),
  .out1({ S2032 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_788_ (
  .in1({ S2032, S1810 }),
  .out1({ S2034 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_789_ (
  .in1({ S2034, DP_LGU1_in1_3 }),
  .out1({ S2035 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1046_ (
  .in1({ S1828, DP_LGU1_in1_3 }),
  .out1({ S2036 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1047_ (
  .in1({ S2036, S1919 }),
  .out1({ S2037 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_790_ (
  .in1({ S2037, S2035 }),
  .out1({ S2038 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1048_ (
  .in1({ CU_NOT, DP_AC_dout_13 }),
  .out1({ S2039 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1049_ (
  .in1({ S2039, S2105 }),
  .out1({ S2040 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_791_ (
  .in1({ S2040, S2038 }),
  .out1({ S2041 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1050_ (
  .in1({ CU_AND, DP_AC_dout_13 }),
  .out1({ S2042 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_792_ (
  .in1({ S2042, S2112 }),
  .out1({ S2043 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_793_ (
  .in1({ S2043, S2041 }),
  .out1({ S2045 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_335_ (
  .in1({ S2045 }),
  .out1({ DP_LGU1_out_13 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1051_ (
  .in1({ CU_AND, DP_AC_dout_14 }),
  .out1({ S2046 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_336_ (
  .in1({ S2046 }),
  .out1({ S2047 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1052_ (
  .in1({ S2047, DP_LGU1_in1_14 }),
  .out1({ S2048 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1053_ (
  .in1({ S2002, DP_LGU1_in1_1 }),
  .out1({ S2049 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1054_ (
  .in1({ S1574, S1571 }),
  .out1({ S2050 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_794_ (
  .in1({ S2050, DP_LGU1_in1_1 }),
  .out1({ S2051 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1055_ (
  .in1({ S2049, S1686 }),
  .out1({ S2052 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_795_ (
  .in1({ S2052, S2051 }),
  .out1({ S2053 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1056_ (
  .in1({ S1959, S1584 }),
  .out1({ S2055 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1057_ (
  .in1({ S2055, S2065 }),
  .out1({ S2056 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_796_ (
  .in1({ S2056, S2053 }),
  .out1({ S2057 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1058_ (
  .in1({ S2057, S1845 }),
  .out1({ S2058 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1059_ (
  .in1({ S1861, DP_LGU1_in1_3 }),
  .out1({ S2059 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1060_ (
  .in1({ S2059, S2058 }),
  .out1({ S2060 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1061_ (
  .in1({ S2060, S1919 }),
  .out1({ S2061 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1062_ (
  .in1({ CU_NOT, DP_AC_dout_14 }),
  .out1({ S2062 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_337_ (
  .in1({ S2062 }),
  .out1({ S2063 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_797_ (
  .in1({ S2063, CU_AND }),
  .out1({ S2064 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1063_ (
  .in1({ S2064, S2061 }),
  .out1({ S2066 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1064_ (
  .in1({ S2066, S2048 }),
  .out1({ DP_LGU1_out_14 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1065_ (
  .in1({ S1618, S1615 }),
  .out1({ S2067 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1066_ (
  .in1({ S2067, S2001 }),
  .out1({ S2068 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1067_ (
  .in1({ S2027, DP_LGU1_in1_1 }),
  .out1({ S2069 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1068_ (
  .in1({ S2069, S2068 }),
  .out1({ S2070 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1069_ (
  .in1({ S2070, S1686 }),
  .out1({ S2071 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_798_ (
  .in1({ S1981, S1585 }),
  .out1({ S2072 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1070_ (
  .in1({ S1897, S1586 }),
  .out1({ S2073 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_799_ (
  .in1({ S2073, S2072 }),
  .out1({ S2074 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1071_ (
  .in1({ S2074, S2071 }),
  .out1({ S2076 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1072_ (
  .in1({ S1896, DP_LGU1_in1_3 }),
  .out1({ S2077 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_338_ (
  .in1({ S2077 }),
  .out1({ S2078 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1073_ (
  .in1({ S2078, S1889 }),
  .out1({ S2079 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1074_ (
  .in1({ S2079, S2076 }),
  .out1({ S2080 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1075_ (
  .in1({ S2080, S2096 }),
  .out1({ S2081 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1076_ (
  .in1({ CU_NOT, DP_AC_dout_15 }),
  .out1({ S2082 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_339_ (
  .in1({ S2082 }),
  .out1({ S2083 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_800_ (
  .in1({ S2083, CU_AND }),
  .out1({ S2084 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1077_ (
  .in1({ S2084, S2081 }),
  .out1({ S2085 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1078_ (
  .in1({ CU_AND, DP_AC_dout_15 }),
  .out1({ S2087 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_340_ (
  .in1({ S2087 }),
  .out1({ S2088 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1079_ (
  .in1({ S2088, DP_LGU1_in1_15 }),
  .out1({ S2089 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1080_ (
  .in1({ S2089, S2085 }),
  .out1({ DP_LGU1_N })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1081_ (
  .in1({ S1801, S1595 }),
  .out1({ S2090 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_801_ (
  .in1({ S2090, DP_LGU1_out_1 }),
  .out1({ S2091 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_802_ (
  .in1({ DP_LGU1_out_10, DP_LGU1_out_7 }),
  .out1({ S2092 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1082_ (
  .in1({ S2092, S2091 }),
  .out1({ S2093 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_803_ (
  .in1({ S2093, DP_LGU1_out_11 }),
  .out1({ S2094 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1083_ (
  .in1({ S2094, S2025 }),
  .out1({ S2095 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1084_ (
  .in1({ S2045, S1869 }),
  .out1({ S2097 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_804_ (
  .in1({ S2097, DP_LGU1_out_14 }),
  .out1({ S2098 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1085_ (
  .in1({ S1954, S1928 }),
  .out1({ S2099 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_805_ (
  .in1({ S2099, DP_LGU1_N }),
  .out1({ S2100 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1086_ (
  .in1({ S2100, S1726 }),
  .out1({ S2101 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1087_ (
  .in1({ S1836, S1770 }),
  .out1({ S2102 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_806_ (
  .in1({ S2102, S2101 }),
  .out1({ S2103 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1088_ (
  .in1({ S2103, S2098 }),
  .out1({ S2104 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_807_ (
  .in1({ S2104, S2095 }),
  .out1({ DP_LGU1_Z })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_341_ (
  .in1({ CU_ldOF }),
  .out1({ S2144 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_808_ (
  .in1({ CU_ldOF, S13 }),
  .out1({ S2145 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1089_ (
  .in1({ S2145, DP_IMM1_in1_0 }),
  .out1({ S2146 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_809_ (
  .in1({ S2144, S14 }),
  .out1({ S2147 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1090_ (
  .in1({ S2147, DP_OF_din_0 }),
  .out1({ S2148 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1091_ (
  .in1({ S2148, S2146 }),
  .out1({ S2140 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1092_ (
  .in1({ S2145, DP_IMM1_in1_1 }),
  .out1({ S2149 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1093_ (
  .in1({ S2147, DP_OF_din_1 }),
  .out1({ S2150 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1094_ (
  .in1({ S2150, S2149 }),
  .out1({ S2141 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1095_ (
  .in1({ S2145, DP_IMM1_in1_2 }),
  .out1({ S2151 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1096_ (
  .in1({ S2147, DP_OF_din_2 }),
  .out1({ S2152 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1097_ (
  .in1({ S2152, S2151 }),
  .out1({ S2142 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1098_ (
  .in1({ S2145, DP_IMM1_in1_3 }),
  .out1({ S2153 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1099_ (
  .in1({ S2147, DP_OF_din_3 }),
  .out1({ S2154 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1100_ (
  .in1({ S2154, S2153 }),
  .out1({ S2143 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_51_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2140 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IMM1_in1_0 }),
  .Si({ S3075 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_52_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2141 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IMM1_in1_1 }),
  .Si({ S3074 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_53_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2142 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IMM1_in1_2 }),
  .Si({ S3073 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_54_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2143 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IMM1_in1_3 }),
  .Si({ S3094 }),
  .global_reset({ 1'b0 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_342_ (
  .in1({ CU_ldPC }),
  .out1({ S2172 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_810_ (
  .in1({ CU_ldPC, S15 }),
  .out1({ S2173 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1101_ (
  .in1({ S2173, DP_INC_1_in_0 }),
  .out1({ S2174 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_811_ (
  .in1({ S2172, S16 }),
  .out1({ S2175 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1102_ (
  .in1({ S2175, DP_PC_din_0 }),
  .out1({ S2176 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1103_ (
  .in1({ S2176, S2174 }),
  .out1({ S2155 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1104_ (
  .in1({ S2173, DP_INC_1_in_1 }),
  .out1({ S2177 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1105_ (
  .in1({ S2175, DP_PC_din_1 }),
  .out1({ S2178 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1106_ (
  .in1({ S2178, S2177 }),
  .out1({ S2156 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1107_ (
  .in1({ S2173, DP_INC_1_in_2 }),
  .out1({ S2179 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1108_ (
  .in1({ S2175, DP_PC_din_2 }),
  .out1({ S2180 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1109_ (
  .in1({ S2180, S2179 }),
  .out1({ S2157 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1110_ (
  .in1({ S2173, DP_INC_1_in_3 }),
  .out1({ S2181 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1111_ (
  .in1({ S2175, DP_PC_din_3 }),
  .out1({ S2182 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1112_ (
  .in1({ S2182, S2181 }),
  .out1({ S2158 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1113_ (
  .in1({ S2173, DP_INC_1_in_4 }),
  .out1({ S2183 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1114_ (
  .in1({ S2175, DP_PC_din_4 }),
  .out1({ S2184 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1115_ (
  .in1({ S2184, S2183 }),
  .out1({ S2159 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1116_ (
  .in1({ S2173, DP_INC_1_in_5 }),
  .out1({ S2185 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1117_ (
  .in1({ S2175, DP_PC_din_5 }),
  .out1({ S2186 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1118_ (
  .in1({ S2186, S2185 }),
  .out1({ S2160 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1119_ (
  .in1({ S2173, DP_INC_1_in_6 }),
  .out1({ S2187 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1120_ (
  .in1({ S2175, DP_PC_din_6 }),
  .out1({ S2188 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1121_ (
  .in1({ S2188, S2187 }),
  .out1({ S2161 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1122_ (
  .in1({ S2173, DP_INC_1_in_7 }),
  .out1({ S2189 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1123_ (
  .in1({ S2175, DP_PC_din_7 }),
  .out1({ S2190 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1124_ (
  .in1({ S2190, S2189 }),
  .out1({ S2162 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1125_ (
  .in1({ S2173, DP_INC_1_in_8 }),
  .out1({ S2191 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1126_ (
  .in1({ S2175, DP_PC_din_8 }),
  .out1({ S2192 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1127_ (
  .in1({ S2192, S2191 }),
  .out1({ S2163 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1128_ (
  .in1({ S2173, DP_INC_1_in_9 }),
  .out1({ S2193 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1129_ (
  .in1({ S2175, DP_PC_din_9 }),
  .out1({ S2194 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1130_ (
  .in1({ S2194, S2193 }),
  .out1({ S2164 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1131_ (
  .in1({ S2173, DP_INC_1_in_10 }),
  .out1({ S2195 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1132_ (
  .in1({ S2175, DP_PC_din_10 }),
  .out1({ S2196 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1133_ (
  .in1({ S2196, S2195 }),
  .out1({ S2165 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1134_ (
  .in1({ S2173, DP_INC_1_in_11 }),
  .out1({ S2197 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1135_ (
  .in1({ S2175, DP_PC_din_11 }),
  .out1({ S2198 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1136_ (
  .in1({ S2198, S2197 }),
  .out1({ S2166 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1137_ (
  .in1({ S2173, DP_INC_1_in_12 }),
  .out1({ S2199 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1138_ (
  .in1({ S2175, DP_PC_din_12 }),
  .out1({ S2200 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1139_ (
  .in1({ S2200, S2199 }),
  .out1({ S2167 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1140_ (
  .in1({ S2173, DP_INC_1_in_13 }),
  .out1({ S2201 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1141_ (
  .in1({ S2175, DP_PC_din_13 }),
  .out1({ S2202 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1142_ (
  .in1({ S2202, S2201 }),
  .out1({ S2168 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1143_ (
  .in1({ S2173, DP_INC_1_in_14 }),
  .out1({ S2203 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1144_ (
  .in1({ S2175, DP_PC_din_14 }),
  .out1({ S2204 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1145_ (
  .in1({ S2204, S2203 }),
  .out1({ S2169 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1146_ (
  .in1({ S2173, DP_INC_1_in_15 }),
  .out1({ S2205 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1147_ (
  .in1({ S2175, DP_PC_din_15 }),
  .out1({ S2171 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1148_ (
  .in1({ S2171, S2205 }),
  .out1({ S2170 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_55_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2155 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_0 }),
  .Si({ S3090 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_56_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2156 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_1 }),
  .Si({ S3089 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_57_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2157 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_2 }),
  .Si({ S3088 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_58_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2158 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_3 }),
  .Si({ S3087 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_59_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2159 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_4 }),
  .Si({ S3086 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_60_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2160 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_5 }),
  .Si({ S3085 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_61_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2161 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_6 }),
  .Si({ S3084 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_62_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2162 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_7 }),
  .Si({ S3083 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_63_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2163 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_8 }),
  .Si({ S3082 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_64_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2164 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_9 }),
  .Si({ S3081 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_65_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2165 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_10 }),
  .Si({ S3080 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_66_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2166 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_11 }),
  .Si({ S3079 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_67_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2167 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_12 }),
  .Si({ S3078 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_68_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2168 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_13 }),
  .Si({ S3077 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_69_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2169 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_14 }),
  .Si({ S3076 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_70_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2170 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_15 }),
  .Si({ S3095 }),
  .global_reset({ 1'b0 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_343_ (
  .in1({ DP_SR_C_dout }),
  .out1({ S2208 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1149_ (
  .in1({ DP_SR_C_din, CU_ldSR_1 }),
  .out1({ S2209 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_344_ (
  .in1({ S2209 }),
  .out1({ S2210 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_812_ (
  .in1({ S2208, CU_ldSR_1 }),
  .out1({ S2211 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_813_ (
  .in1({ S2211, S2210 }),
  .out1({ S2207 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_814_ (
  .in1({ S2207, S17 }),
  .out1({ S2206 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_71_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2206 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_SR_C_dout }),
  .Si({ S3096 }),
  .global_reset({ 1'b0 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_345_ (
  .in1({ DP_SR_N_dout }),
  .out1({ S2214 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1150_ (
  .in1({ DP_SR_N_din, CU_ldSR_2 }),
  .out1({ S2215 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_346_ (
  .in1({ S2215 }),
  .out1({ S2216 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_815_ (
  .in1({ S2214, CU_ldSR_2 }),
  .out1({ S2217 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_816_ (
  .in1({ S2217, S2216 }),
  .out1({ S2213 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_817_ (
  .in1({ S2213, S18 }),
  .out1({ S2212 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_72_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2212 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_SR_N_dout }),
  .Si({ S3097 }),
  .global_reset({ 1'b0 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_347_ (
  .in1({ DP_SR_V_dout }),
  .out1({ S2220 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1151_ (
  .in1({ DP_SR_V_din, CU_ldSR_0 }),
  .out1({ S2221 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_348_ (
  .in1({ S2221 }),
  .out1({ S2222 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_818_ (
  .in1({ S2220, CU_ldSR_0 }),
  .out1({ S2223 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_819_ (
  .in1({ S2223, S2222 }),
  .out1({ S2219 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_820_ (
  .in1({ S2219, S19 }),
  .out1({ S2218 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_73_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2218 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_SR_V_dout }),
  .Si({ S3098 }),
  .global_reset({ 1'b0 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_349_ (
  .in1({ DP_SR_Z_dout }),
  .out1({ S2226 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1152_ (
  .in1({ DP_SR_Z_din, CU_ldSR_3 }),
  .out1({ S2227 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_350_ (
  .in1({ S2227 }),
  .out1({ S2228 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_821_ (
  .in1({ S2226, CU_ldSR_3 }),
  .out1({ S2229 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_822_ (
  .in1({ S2229, S2228 }),
  .out1({ S2225 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_823_ (
  .in1({ S2225, S20 }),
  .out1({ S2224 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_74_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2224 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_SR_Z_dout }),
  .Si({ S3099 }),
  .global_reset({ 1'b0 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_351_ (
  .in1({ DP_LGU1_out_0 }),
  .out1({ S2375 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_352_ (
  .in1({ CU_selIMM_AC }),
  .out1({ S2376 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_353_ (
  .in1({ DP_LGU1_out_1 }),
  .out1({ S2377 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_354_ (
  .in1({ DP_LGU1_out_2 }),
  .out1({ S2378 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_355_ (
  .in1({ DP_LGU1_out_3 }),
  .out1({ S2379 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_356_ (
  .in1({ DP_LGU1_out_4 }),
  .out1({ S2380 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_357_ (
  .in1({ DP_LGU1_out_5 }),
  .out1({ S2381 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_358_ (
  .in1({ DP_LGU1_out_6 }),
  .out1({ S2382 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_359_ (
  .in1({ DP_LGU1_out_7 }),
  .out1({ S2383 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_360_ (
  .in1({ DP_LGU1_out_8 }),
  .out1({ S2384 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_361_ (
  .in1({ DP_LGU1_out_9 }),
  .out1({ S2385 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_362_ (
  .in1({ DP_LGU1_out_10 }),
  .out1({ S2386 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_363_ (
  .in1({ DP_LGU1_out_11 }),
  .out1({ S2387 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_364_ (
  .in1({ DP_LGU1_out_12 }),
  .out1({ S2388 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_365_ (
  .in1({ DP_LGU1_out_13 }),
  .out1({ S2389 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_366_ (
  .in1({ DP_LGU1_out_14 }),
  .out1({ S2390 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_367_ (
  .in1({ DP_LGU1_N }),
  .out1({ S2230 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_824_ (
  .in1({ S2376, DP_IMM1_out_0 }),
  .out1({ S2231 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1153_ (
  .in1({ CU_selARU_AC, DP_ARU1_out_0 }),
  .out1({ S2232 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_368_ (
  .in1({ S2232 }),
  .out1({ S2233 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_825_ (
  .in1({ CU_selARU_AC, S2375 }),
  .out1({ S2234 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_826_ (
  .in1({ S2234, S2233 }),
  .out1({ S2235 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_827_ (
  .in1({ S2235, CU_selMEM_AC }),
  .out1({ S2236 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1154_ (
  .in1({ CU_selMEM_AC, dataBus[0] }),
  .out1({ S2237 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1155_ (
  .in1({ S2237, S2376 }),
  .out1({ S2238 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_828_ (
  .in1({ S2238, S2236 }),
  .out1({ S2239 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_829_ (
  .in1({ S2239, S2231 }),
  .out1({ DP_AC_din_0 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_830_ (
  .in1({ DP_IMM1_out_1, S2376 }),
  .out1({ S2240 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1156_ (
  .in1({ DP_ARU1_out_1, CU_selARU_AC }),
  .out1({ S2241 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_369_ (
  .in1({ S2241 }),
  .out1({ S2242 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_831_ (
  .in1({ S2377, CU_selARU_AC }),
  .out1({ S2243 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_832_ (
  .in1({ S2243, S2242 }),
  .out1({ S2244 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_833_ (
  .in1({ S2244, CU_selMEM_AC }),
  .out1({ S2245 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1157_ (
  .in1({ dataBus[1], CU_selMEM_AC }),
  .out1({ S2246 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1158_ (
  .in1({ S2246, S2376 }),
  .out1({ S2247 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_834_ (
  .in1({ S2247, S2245 }),
  .out1({ S2248 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_835_ (
  .in1({ S2248, S2240 }),
  .out1({ DP_AC_din_1 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_836_ (
  .in1({ DP_IMM1_out_2, S2376 }),
  .out1({ S2249 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1159_ (
  .in1({ DP_ARU1_out_2, CU_selARU_AC }),
  .out1({ S2250 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_370_ (
  .in1({ S2250 }),
  .out1({ S2251 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_837_ (
  .in1({ S2378, CU_selARU_AC }),
  .out1({ S2252 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_838_ (
  .in1({ S2252, S2251 }),
  .out1({ S2253 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_839_ (
  .in1({ S2253, CU_selMEM_AC }),
  .out1({ S2254 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1160_ (
  .in1({ dataBus[2], CU_selMEM_AC }),
  .out1({ S2255 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1161_ (
  .in1({ S2255, S2376 }),
  .out1({ S2256 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_840_ (
  .in1({ S2256, S2254 }),
  .out1({ S2257 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_841_ (
  .in1({ S2257, S2249 }),
  .out1({ DP_AC_din_2 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_842_ (
  .in1({ DP_IMM1_out_3, S2376 }),
  .out1({ S2258 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1162_ (
  .in1({ DP_ARU1_out_3, CU_selARU_AC }),
  .out1({ S2259 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_371_ (
  .in1({ S2259 }),
  .out1({ S2260 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_843_ (
  .in1({ S2379, CU_selARU_AC }),
  .out1({ S2261 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_844_ (
  .in1({ S2261, S2260 }),
  .out1({ S2262 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_845_ (
  .in1({ S2262, CU_selMEM_AC }),
  .out1({ S2263 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1163_ (
  .in1({ dataBus[3], CU_selMEM_AC }),
  .out1({ S2264 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1164_ (
  .in1({ S2264, S2376 }),
  .out1({ S2265 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_846_ (
  .in1({ S2265, S2263 }),
  .out1({ S2266 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_847_ (
  .in1({ S2266, S2258 }),
  .out1({ DP_AC_din_3 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_848_ (
  .in1({ DP_IMM1_out_4, S2376 }),
  .out1({ S2267 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1165_ (
  .in1({ DP_ARU1_out_4, CU_selARU_AC }),
  .out1({ S2268 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_372_ (
  .in1({ S2268 }),
  .out1({ S2269 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_849_ (
  .in1({ S2380, CU_selARU_AC }),
  .out1({ S2270 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_850_ (
  .in1({ S2270, S2269 }),
  .out1({ S2271 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_851_ (
  .in1({ S2271, CU_selMEM_AC }),
  .out1({ S2272 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1166_ (
  .in1({ dataBus[4], CU_selMEM_AC }),
  .out1({ S2273 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1167_ (
  .in1({ S2273, S2376 }),
  .out1({ S2274 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_852_ (
  .in1({ S2274, S2272 }),
  .out1({ S2275 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_853_ (
  .in1({ S2275, S2267 }),
  .out1({ DP_AC_din_4 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_854_ (
  .in1({ DP_IMM1_out_5, S2376 }),
  .out1({ S2276 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1168_ (
  .in1({ DP_ARU1_out_5, CU_selARU_AC }),
  .out1({ S2277 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_373_ (
  .in1({ S2277 }),
  .out1({ S2278 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_855_ (
  .in1({ S2381, CU_selARU_AC }),
  .out1({ S2279 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_856_ (
  .in1({ S2279, S2278 }),
  .out1({ S2280 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_857_ (
  .in1({ S2280, CU_selMEM_AC }),
  .out1({ S2281 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1169_ (
  .in1({ dataBus[5], CU_selMEM_AC }),
  .out1({ S2282 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1170_ (
  .in1({ S2282, S2376 }),
  .out1({ S2283 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_858_ (
  .in1({ S2283, S2281 }),
  .out1({ S2284 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_859_ (
  .in1({ S2284, S2276 }),
  .out1({ DP_AC_din_5 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_860_ (
  .in1({ DP_IMM1_out_6, S2376 }),
  .out1({ S2285 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1171_ (
  .in1({ DP_ARU1_out_6, CU_selARU_AC }),
  .out1({ S2286 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_374_ (
  .in1({ S2286 }),
  .out1({ S2287 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_861_ (
  .in1({ S2382, CU_selARU_AC }),
  .out1({ S2288 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_862_ (
  .in1({ S2288, S2287 }),
  .out1({ S2289 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_863_ (
  .in1({ S2289, CU_selMEM_AC }),
  .out1({ S2290 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1172_ (
  .in1({ dataBus[6], CU_selMEM_AC }),
  .out1({ S2291 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1173_ (
  .in1({ S2291, S2376 }),
  .out1({ S2292 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_864_ (
  .in1({ S2292, S2290 }),
  .out1({ S2293 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_865_ (
  .in1({ S2293, S2285 }),
  .out1({ DP_AC_din_6 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_866_ (
  .in1({ DP_IMM1_out_7, S2376 }),
  .out1({ S2294 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1174_ (
  .in1({ DP_ARU1_out_7, CU_selARU_AC }),
  .out1({ S2295 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_375_ (
  .in1({ S2295 }),
  .out1({ S2296 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_867_ (
  .in1({ S2383, CU_selARU_AC }),
  .out1({ S2297 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_868_ (
  .in1({ S2297, S2296 }),
  .out1({ S2298 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_869_ (
  .in1({ S2298, CU_selMEM_AC }),
  .out1({ S2299 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1175_ (
  .in1({ dataBus[7], CU_selMEM_AC }),
  .out1({ S2300 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1176_ (
  .in1({ S2300, S2376 }),
  .out1({ S2301 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_870_ (
  .in1({ S2301, S2299 }),
  .out1({ S2302 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_871_ (
  .in1({ S2302, S2294 }),
  .out1({ DP_AC_din_7 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_872_ (
  .in1({ DP_IMM1_out_8, S2376 }),
  .out1({ S2303 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1177_ (
  .in1({ DP_ARU1_out_8, CU_selARU_AC }),
  .out1({ S2304 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_376_ (
  .in1({ S2304 }),
  .out1({ S2305 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_873_ (
  .in1({ S2384, CU_selARU_AC }),
  .out1({ S2306 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_874_ (
  .in1({ S2306, S2305 }),
  .out1({ S2307 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_875_ (
  .in1({ S2307, CU_selMEM_AC }),
  .out1({ S2308 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1178_ (
  .in1({ dataBus[8], CU_selMEM_AC }),
  .out1({ S2309 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1179_ (
  .in1({ S2309, S2376 }),
  .out1({ S2310 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_876_ (
  .in1({ S2310, S2308 }),
  .out1({ S2311 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_877_ (
  .in1({ S2311, S2303 }),
  .out1({ DP_AC_din_8 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_878_ (
  .in1({ DP_IMM1_out_9, S2376 }),
  .out1({ S2312 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1180_ (
  .in1({ DP_ARU1_out_9, CU_selARU_AC }),
  .out1({ S2313 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_377_ (
  .in1({ S2313 }),
  .out1({ S2314 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_879_ (
  .in1({ S2385, CU_selARU_AC }),
  .out1({ S2315 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_880_ (
  .in1({ S2315, S2314 }),
  .out1({ S2316 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_881_ (
  .in1({ S2316, CU_selMEM_AC }),
  .out1({ S2317 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1181_ (
  .in1({ dataBus[9], CU_selMEM_AC }),
  .out1({ S2318 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1182_ (
  .in1({ S2318, S2376 }),
  .out1({ S2319 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_882_ (
  .in1({ S2319, S2317 }),
  .out1({ S2320 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_883_ (
  .in1({ S2320, S2312 }),
  .out1({ DP_AC_din_9 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_884_ (
  .in1({ DP_IMM1_out_10, S2376 }),
  .out1({ S2321 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1183_ (
  .in1({ DP_ARU1_out_10, CU_selARU_AC }),
  .out1({ S2322 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_378_ (
  .in1({ S2322 }),
  .out1({ S2323 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_885_ (
  .in1({ S2386, CU_selARU_AC }),
  .out1({ S2324 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_886_ (
  .in1({ S2324, S2323 }),
  .out1({ S2325 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_887_ (
  .in1({ S2325, CU_selMEM_AC }),
  .out1({ S2326 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1184_ (
  .in1({ dataBus[10], CU_selMEM_AC }),
  .out1({ S2327 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1185_ (
  .in1({ S2327, S2376 }),
  .out1({ S2328 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_888_ (
  .in1({ S2328, S2326 }),
  .out1({ S2329 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_889_ (
  .in1({ S2329, S2321 }),
  .out1({ DP_AC_din_10 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_890_ (
  .in1({ DP_IMM1_out_11, S2376 }),
  .out1({ S2330 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1186_ (
  .in1({ DP_ARU1_out_11, CU_selARU_AC }),
  .out1({ S2331 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_379_ (
  .in1({ S2331 }),
  .out1({ S2332 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_891_ (
  .in1({ S2387, CU_selARU_AC }),
  .out1({ S2333 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_892_ (
  .in1({ S2333, S2332 }),
  .out1({ S2334 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_893_ (
  .in1({ S2334, CU_selMEM_AC }),
  .out1({ S2335 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1187_ (
  .in1({ dataBus[11], CU_selMEM_AC }),
  .out1({ S2336 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1188_ (
  .in1({ S2336, S2376 }),
  .out1({ S2337 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_894_ (
  .in1({ S2337, S2335 }),
  .out1({ S2338 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_895_ (
  .in1({ S2338, S2330 }),
  .out1({ DP_AC_din_11 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_896_ (
  .in1({ DP_IMM1_out_12, S2376 }),
  .out1({ S2339 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1189_ (
  .in1({ DP_ARU1_out_12, CU_selARU_AC }),
  .out1({ S2340 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_380_ (
  .in1({ S2340 }),
  .out1({ S2341 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_897_ (
  .in1({ S2388, CU_selARU_AC }),
  .out1({ S2342 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_898_ (
  .in1({ S2342, S2341 }),
  .out1({ S2343 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_899_ (
  .in1({ S2343, CU_selMEM_AC }),
  .out1({ S2344 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1190_ (
  .in1({ dataBus[12], CU_selMEM_AC }),
  .out1({ S2345 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1191_ (
  .in1({ S2345, S2376 }),
  .out1({ S2346 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_900_ (
  .in1({ S2346, S2344 }),
  .out1({ S2347 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_901_ (
  .in1({ S2347, S2339 }),
  .out1({ DP_AC_din_12 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_902_ (
  .in1({ DP_IMM1_out_13, S2376 }),
  .out1({ S2348 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1192_ (
  .in1({ DP_ARU1_out_13, CU_selARU_AC }),
  .out1({ S2349 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_381_ (
  .in1({ S2349 }),
  .out1({ S2350 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_903_ (
  .in1({ S2389, CU_selARU_AC }),
  .out1({ S2351 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_904_ (
  .in1({ S2351, S2350 }),
  .out1({ S2352 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_905_ (
  .in1({ S2352, CU_selMEM_AC }),
  .out1({ S2353 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1193_ (
  .in1({ dataBus[13], CU_selMEM_AC }),
  .out1({ S2354 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1194_ (
  .in1({ S2354, S2376 }),
  .out1({ S2355 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_906_ (
  .in1({ S2355, S2353 }),
  .out1({ S2356 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_907_ (
  .in1({ S2356, S2348 }),
  .out1({ DP_AC_din_13 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_908_ (
  .in1({ DP_IMM1_out_14, S2376 }),
  .out1({ S2357 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1195_ (
  .in1({ DP_ARU1_out_14, CU_selARU_AC }),
  .out1({ S2358 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_382_ (
  .in1({ S2358 }),
  .out1({ S2359 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_909_ (
  .in1({ S2390, CU_selARU_AC }),
  .out1({ S2360 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_910_ (
  .in1({ S2360, S2359 }),
  .out1({ S2361 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_911_ (
  .in1({ S2361, CU_selMEM_AC }),
  .out1({ S2362 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1196_ (
  .in1({ dataBus[14], CU_selMEM_AC }),
  .out1({ S2363 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1197_ (
  .in1({ S2363, S2376 }),
  .out1({ S2364 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_912_ (
  .in1({ S2364, S2362 }),
  .out1({ S2365 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_913_ (
  .in1({ S2365, S2357 }),
  .out1({ DP_AC_din_14 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_914_ (
  .in1({ DP_IMM1_out_15, S2376 }),
  .out1({ S2366 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1198_ (
  .in1({ DP_ARU1_N, CU_selARU_AC }),
  .out1({ S2367 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_383_ (
  .in1({ S2367 }),
  .out1({ S2368 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_915_ (
  .in1({ S2230, CU_selARU_AC }),
  .out1({ S2369 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_916_ (
  .in1({ S2369, S2368 }),
  .out1({ S2370 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_917_ (
  .in1({ S2370, CU_selMEM_AC }),
  .out1({ S2371 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1199_ (
  .in1({ dataBus[15], CU_selMEM_AC }),
  .out1({ S2372 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1200_ (
  .in1({ S2372, S2376 }),
  .out1({ S2373 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_918_ (
  .in1({ S2373, S2371 }),
  .out1({ S2374 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_919_ (
  .in1({ S2374, S2366 }),
  .out1({ DP_AC_din_15 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_384_ (
  .in1({ 1'bz }),
  .out1({ S2391 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_385_ (
  .in1({ CU_selSET_SR }),
  .out1({ S2392 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_386_ (
  .in1({ 1'bz }),
  .out1({ S2393 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_387_ (
  .in1({ 1'bz }),
  .out1({ S2394 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_388_ (
  .in1({ 1'bz }),
  .out1({ S2395 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_920_ (
  .in1({ S2392, CU_inst_0 }),
  .out1({ S2396 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1201_ (
  .in1({ CU_selARU_SR, DP_ARU1_V }),
  .out1({ S2397 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_389_ (
  .in1({ S2397 }),
  .out1({ S2398 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_921_ (
  .in1({ CU_selARU_SR, S2391 }),
  .out1({ S2399 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_922_ (
  .in1({ S2399, S2398 }),
  .out1({ S2400 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_923_ (
  .in1({ S2400, CU_selLGU_SR }),
  .out1({ S2401 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1202_ (
  .in1({ CU_selLGU_SR, 1'bz }),
  .out1({ S2402 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1203_ (
  .in1({ S2402, S2392 }),
  .out1({ S2403 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_924_ (
  .in1({ S2403, S2401 }),
  .out1({ S2404 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_925_ (
  .in1({ S2404, S2396 }),
  .out1({ DP_SR_V_din })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_926_ (
  .in1({ CU_inst_1, S2392 }),
  .out1({ S2405 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1204_ (
  .in1({ DP_ARU1_C, CU_selARU_SR }),
  .out1({ S2406 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_390_ (
  .in1({ S2406 }),
  .out1({ S2407 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_927_ (
  .in1({ S2393, CU_selARU_SR }),
  .out1({ S2408 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_928_ (
  .in1({ S2408, S2407 }),
  .out1({ S2409 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_929_ (
  .in1({ S2409, CU_selLGU_SR }),
  .out1({ S2410 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1205_ (
  .in1({ 1'bz, CU_selLGU_SR }),
  .out1({ S2411 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1206_ (
  .in1({ S2411, S2392 }),
  .out1({ S2412 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_930_ (
  .in1({ S2412, S2410 }),
  .out1({ S2413 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_931_ (
  .in1({ S2413, S2405 }),
  .out1({ DP_SR_C_din })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_932_ (
  .in1({ CU_inst_2, S2392 }),
  .out1({ S2414 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1207_ (
  .in1({ DP_ARU1_N, CU_selARU_SR }),
  .out1({ S2415 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_391_ (
  .in1({ S2415 }),
  .out1({ S2416 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_933_ (
  .in1({ S2394, CU_selARU_SR }),
  .out1({ S2417 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_934_ (
  .in1({ S2417, S2416 }),
  .out1({ S2418 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_935_ (
  .in1({ S2418, CU_selLGU_SR }),
  .out1({ S2419 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1208_ (
  .in1({ DP_LGU1_N, CU_selLGU_SR }),
  .out1({ S2420 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1209_ (
  .in1({ S2420, S2392 }),
  .out1({ S2421 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_936_ (
  .in1({ S2421, S2419 }),
  .out1({ S2422 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_937_ (
  .in1({ S2422, S2414 }),
  .out1({ DP_SR_N_din })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_938_ (
  .in1({ CU_inst_3, S2392 }),
  .out1({ S2423 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1210_ (
  .in1({ DP_ARU1_Z, CU_selARU_SR }),
  .out1({ S2424 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_392_ (
  .in1({ S2424 }),
  .out1({ S2425 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_939_ (
  .in1({ S2395, CU_selARU_SR }),
  .out1({ S2426 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_940_ (
  .in1({ S2426, S2425 }),
  .out1({ S2427 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_941_ (
  .in1({ S2427, CU_selLGU_SR }),
  .out1({ S2428 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1211_ (
  .in1({ DP_LGU1_Z, CU_selLGU_SR }),
  .out1({ S2429 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1212_ (
  .in1({ S2429, S2392 }),
  .out1({ S2430 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_942_ (
  .in1({ S2430, S2428 }),
  .out1({ S2431 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_943_ (
  .in1({ S2431, S2423 }),
  .out1({ DP_SR_Z_din })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_393_ (
  .in1({ 1'bz }),
  .out1({ S2577 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_394_ (
  .in1({ CU_selINC_PC }),
  .out1({ S2578 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_395_ (
  .in1({ 1'bz }),
  .out1({ S2579 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_396_ (
  .in1({ 1'bz }),
  .out1({ S2580 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_397_ (
  .in1({ 1'bz }),
  .out1({ S2581 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_398_ (
  .in1({ 1'bz }),
  .out1({ S2582 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_399_ (
  .in1({ 1'bz }),
  .out1({ S2583 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_400_ (
  .in1({ 1'bz }),
  .out1({ S2584 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_401_ (
  .in1({ 1'bz }),
  .out1({ S2585 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_402_ (
  .in1({ 1'bz }),
  .out1({ S2586 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_403_ (
  .in1({ 1'bz }),
  .out1({ S2587 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_404_ (
  .in1({ 1'bz }),
  .out1({ S2588 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_405_ (
  .in1({ 1'bz }),
  .out1({ S2589 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_406_ (
  .in1({ 1'bz }),
  .out1({ S2590 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_407_ (
  .in1({ 1'bz }),
  .out1({ S2591 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_408_ (
  .in1({ 1'bz }),
  .out1({ S2592 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_409_ (
  .in1({ 1'bz }),
  .out1({ S2432 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_944_ (
  .in1({ S2578, DP_INC_1_out_0 }),
  .out1({ S2433 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1213_ (
  .in1({ CU_selIMM_PC, DP_IMM1_out_0 }),
  .out1({ S2434 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_410_ (
  .in1({ S2434 }),
  .out1({ S2435 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_945_ (
  .in1({ CU_selIMM_PC, S2577 }),
  .out1({ S2436 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_946_ (
  .in1({ S2436, S2435 }),
  .out1({ S2437 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_947_ (
  .in1({ S2437, CU_selMEM_PC }),
  .out1({ S2438 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1214_ (
  .in1({ CU_selMEM_PC, dataBus[0] }),
  .out1({ S2439 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1215_ (
  .in1({ S2439, S2578 }),
  .out1({ S2440 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_948_ (
  .in1({ S2440, S2438 }),
  .out1({ S2441 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_949_ (
  .in1({ S2441, S2433 }),
  .out1({ DP_PC_din_0 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_950_ (
  .in1({ DP_INC_1_out_1, S2578 }),
  .out1({ S2442 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1216_ (
  .in1({ DP_IMM1_out_1, CU_selIMM_PC }),
  .out1({ S2443 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_411_ (
  .in1({ S2443 }),
  .out1({ S2444 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_951_ (
  .in1({ S2579, CU_selIMM_PC }),
  .out1({ S2445 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_952_ (
  .in1({ S2445, S2444 }),
  .out1({ S2446 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_953_ (
  .in1({ S2446, CU_selMEM_PC }),
  .out1({ S2447 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1217_ (
  .in1({ dataBus[1], CU_selMEM_PC }),
  .out1({ S2448 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1218_ (
  .in1({ S2448, S2578 }),
  .out1({ S2449 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_954_ (
  .in1({ S2449, S2447 }),
  .out1({ S2450 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_955_ (
  .in1({ S2450, S2442 }),
  .out1({ DP_PC_din_1 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_956_ (
  .in1({ DP_INC_1_out_2, S2578 }),
  .out1({ S2451 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1219_ (
  .in1({ DP_IMM1_out_2, CU_selIMM_PC }),
  .out1({ S2452 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_412_ (
  .in1({ S2452 }),
  .out1({ S2453 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_957_ (
  .in1({ S2580, CU_selIMM_PC }),
  .out1({ S2454 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_958_ (
  .in1({ S2454, S2453 }),
  .out1({ S2455 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_959_ (
  .in1({ S2455, CU_selMEM_PC }),
  .out1({ S2456 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1220_ (
  .in1({ dataBus[2], CU_selMEM_PC }),
  .out1({ S2457 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1221_ (
  .in1({ S2457, S2578 }),
  .out1({ S2458 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_960_ (
  .in1({ S2458, S2456 }),
  .out1({ S2459 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_961_ (
  .in1({ S2459, S2451 }),
  .out1({ DP_PC_din_2 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_962_ (
  .in1({ DP_INC_1_out_3, S2578 }),
  .out1({ S2460 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1222_ (
  .in1({ DP_IMM1_out_3, CU_selIMM_PC }),
  .out1({ S2461 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_413_ (
  .in1({ S2461 }),
  .out1({ S2462 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_963_ (
  .in1({ S2581, CU_selIMM_PC }),
  .out1({ S2463 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_964_ (
  .in1({ S2463, S2462 }),
  .out1({ S2464 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_965_ (
  .in1({ S2464, CU_selMEM_PC }),
  .out1({ S2465 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1223_ (
  .in1({ dataBus[3], CU_selMEM_PC }),
  .out1({ S2466 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1224_ (
  .in1({ S2466, S2578 }),
  .out1({ S2467 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_966_ (
  .in1({ S2467, S2465 }),
  .out1({ S2468 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_967_ (
  .in1({ S2468, S2460 }),
  .out1({ DP_PC_din_3 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_968_ (
  .in1({ DP_INC_1_out_4, S2578 }),
  .out1({ S2469 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1225_ (
  .in1({ DP_IMM1_out_4, CU_selIMM_PC }),
  .out1({ S2470 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_414_ (
  .in1({ S2470 }),
  .out1({ S2471 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_969_ (
  .in1({ S2582, CU_selIMM_PC }),
  .out1({ S2472 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_970_ (
  .in1({ S2472, S2471 }),
  .out1({ S2473 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_971_ (
  .in1({ S2473, CU_selMEM_PC }),
  .out1({ S2474 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1226_ (
  .in1({ dataBus[4], CU_selMEM_PC }),
  .out1({ S2475 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1227_ (
  .in1({ S2475, S2578 }),
  .out1({ S2476 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_972_ (
  .in1({ S2476, S2474 }),
  .out1({ S2477 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_973_ (
  .in1({ S2477, S2469 }),
  .out1({ DP_PC_din_4 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_974_ (
  .in1({ DP_INC_1_out_5, S2578 }),
  .out1({ S2478 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1228_ (
  .in1({ DP_IMM1_out_5, CU_selIMM_PC }),
  .out1({ S2479 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_415_ (
  .in1({ S2479 }),
  .out1({ S2480 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_975_ (
  .in1({ S2583, CU_selIMM_PC }),
  .out1({ S2481 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_976_ (
  .in1({ S2481, S2480 }),
  .out1({ S2482 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_977_ (
  .in1({ S2482, CU_selMEM_PC }),
  .out1({ S2483 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1229_ (
  .in1({ dataBus[5], CU_selMEM_PC }),
  .out1({ S2484 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1230_ (
  .in1({ S2484, S2578 }),
  .out1({ S2485 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_978_ (
  .in1({ S2485, S2483 }),
  .out1({ S2486 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_979_ (
  .in1({ S2486, S2478 }),
  .out1({ DP_PC_din_5 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_980_ (
  .in1({ DP_INC_1_out_6, S2578 }),
  .out1({ S2487 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1231_ (
  .in1({ DP_IMM1_out_6, CU_selIMM_PC }),
  .out1({ S2488 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_416_ (
  .in1({ S2488 }),
  .out1({ S2489 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_981_ (
  .in1({ S2584, CU_selIMM_PC }),
  .out1({ S2490 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_982_ (
  .in1({ S2490, S2489 }),
  .out1({ S2491 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_983_ (
  .in1({ S2491, CU_selMEM_PC }),
  .out1({ S2492 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1232_ (
  .in1({ dataBus[6], CU_selMEM_PC }),
  .out1({ S2493 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1233_ (
  .in1({ S2493, S2578 }),
  .out1({ S2494 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_984_ (
  .in1({ S2494, S2492 }),
  .out1({ S2495 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_985_ (
  .in1({ S2495, S2487 }),
  .out1({ DP_PC_din_6 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_986_ (
  .in1({ DP_INC_1_out_7, S2578 }),
  .out1({ S2496 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1234_ (
  .in1({ DP_IMM1_out_7, CU_selIMM_PC }),
  .out1({ S2497 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_417_ (
  .in1({ S2497 }),
  .out1({ S2498 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_987_ (
  .in1({ S2585, CU_selIMM_PC }),
  .out1({ S2499 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_988_ (
  .in1({ S2499, S2498 }),
  .out1({ S2500 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_989_ (
  .in1({ S2500, CU_selMEM_PC }),
  .out1({ S2501 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1235_ (
  .in1({ dataBus[7], CU_selMEM_PC }),
  .out1({ S2502 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1236_ (
  .in1({ S2502, S2578 }),
  .out1({ S2503 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_990_ (
  .in1({ S2503, S2501 }),
  .out1({ S2504 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_991_ (
  .in1({ S2504, S2496 }),
  .out1({ DP_PC_din_7 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_992_ (
  .in1({ DP_INC_1_out_8, S2578 }),
  .out1({ S2505 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1237_ (
  .in1({ DP_IMM1_out_8, CU_selIMM_PC }),
  .out1({ S2506 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_418_ (
  .in1({ S2506 }),
  .out1({ S2507 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_993_ (
  .in1({ S2586, CU_selIMM_PC }),
  .out1({ S2508 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_994_ (
  .in1({ S2508, S2507 }),
  .out1({ S2509 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_995_ (
  .in1({ S2509, CU_selMEM_PC }),
  .out1({ S2510 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1238_ (
  .in1({ dataBus[8], CU_selMEM_PC }),
  .out1({ S2511 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1239_ (
  .in1({ S2511, S2578 }),
  .out1({ S2512 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_996_ (
  .in1({ S2512, S2510 }),
  .out1({ S2513 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_997_ (
  .in1({ S2513, S2505 }),
  .out1({ DP_PC_din_8 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_998_ (
  .in1({ DP_INC_1_out_9, S2578 }),
  .out1({ S2514 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1240_ (
  .in1({ DP_IMM1_out_9, CU_selIMM_PC }),
  .out1({ S2515 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_419_ (
  .in1({ S2515 }),
  .out1({ S2516 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_999_ (
  .in1({ S2587, CU_selIMM_PC }),
  .out1({ S2517 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1000_ (
  .in1({ S2517, S2516 }),
  .out1({ S2518 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1001_ (
  .in1({ S2518, CU_selMEM_PC }),
  .out1({ S2519 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1241_ (
  .in1({ dataBus[9], CU_selMEM_PC }),
  .out1({ S2520 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1242_ (
  .in1({ S2520, S2578 }),
  .out1({ S2521 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1002_ (
  .in1({ S2521, S2519 }),
  .out1({ S2522 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1003_ (
  .in1({ S2522, S2514 }),
  .out1({ DP_PC_din_9 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1004_ (
  .in1({ DP_INC_1_out_10, S2578 }),
  .out1({ S2523 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1243_ (
  .in1({ DP_IMM1_out_10, CU_selIMM_PC }),
  .out1({ S2524 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_420_ (
  .in1({ S2524 }),
  .out1({ S2525 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1005_ (
  .in1({ S2588, CU_selIMM_PC }),
  .out1({ S2526 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1006_ (
  .in1({ S2526, S2525 }),
  .out1({ S2527 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1007_ (
  .in1({ S2527, CU_selMEM_PC }),
  .out1({ S2528 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1244_ (
  .in1({ dataBus[10], CU_selMEM_PC }),
  .out1({ S2529 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1245_ (
  .in1({ S2529, S2578 }),
  .out1({ S2530 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1008_ (
  .in1({ S2530, S2528 }),
  .out1({ S2531 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1009_ (
  .in1({ S2531, S2523 }),
  .out1({ DP_PC_din_10 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1010_ (
  .in1({ DP_INC_1_out_11, S2578 }),
  .out1({ S2532 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1246_ (
  .in1({ DP_IMM1_out_11, CU_selIMM_PC }),
  .out1({ S2533 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_421_ (
  .in1({ S2533 }),
  .out1({ S2534 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1011_ (
  .in1({ S2589, CU_selIMM_PC }),
  .out1({ S2535 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1012_ (
  .in1({ S2535, S2534 }),
  .out1({ S2536 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1013_ (
  .in1({ S2536, CU_selMEM_PC }),
  .out1({ S2537 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1247_ (
  .in1({ dataBus[11], CU_selMEM_PC }),
  .out1({ S2538 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1248_ (
  .in1({ S2538, S2578 }),
  .out1({ S2539 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1014_ (
  .in1({ S2539, S2537 }),
  .out1({ S2540 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1015_ (
  .in1({ S2540, S2532 }),
  .out1({ DP_PC_din_11 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1016_ (
  .in1({ DP_INC_1_out_12, S2578 }),
  .out1({ S2541 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1249_ (
  .in1({ DP_IMM1_out_12, CU_selIMM_PC }),
  .out1({ S2542 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_422_ (
  .in1({ S2542 }),
  .out1({ S2543 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1017_ (
  .in1({ S2590, CU_selIMM_PC }),
  .out1({ S2544 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1018_ (
  .in1({ S2544, S2543 }),
  .out1({ S2545 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1019_ (
  .in1({ S2545, CU_selMEM_PC }),
  .out1({ S2546 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1250_ (
  .in1({ dataBus[12], CU_selMEM_PC }),
  .out1({ S2547 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1251_ (
  .in1({ S2547, S2578 }),
  .out1({ S2548 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1020_ (
  .in1({ S2548, S2546 }),
  .out1({ S2549 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1021_ (
  .in1({ S2549, S2541 }),
  .out1({ DP_PC_din_12 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1022_ (
  .in1({ DP_INC_1_out_13, S2578 }),
  .out1({ S2550 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1252_ (
  .in1({ DP_IMM1_out_13, CU_selIMM_PC }),
  .out1({ S2551 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_423_ (
  .in1({ S2551 }),
  .out1({ S2552 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1023_ (
  .in1({ S2591, CU_selIMM_PC }),
  .out1({ S2553 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1024_ (
  .in1({ S2553, S2552 }),
  .out1({ S2554 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1025_ (
  .in1({ S2554, CU_selMEM_PC }),
  .out1({ S2555 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1253_ (
  .in1({ dataBus[13], CU_selMEM_PC }),
  .out1({ S2556 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1254_ (
  .in1({ S2556, S2578 }),
  .out1({ S2557 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1026_ (
  .in1({ S2557, S2555 }),
  .out1({ S2558 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1027_ (
  .in1({ S2558, S2550 }),
  .out1({ DP_PC_din_13 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1028_ (
  .in1({ DP_INC_1_out_14, S2578 }),
  .out1({ S2559 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1255_ (
  .in1({ DP_IMM1_out_14, CU_selIMM_PC }),
  .out1({ S2560 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_424_ (
  .in1({ S2560 }),
  .out1({ S2561 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1029_ (
  .in1({ S2592, CU_selIMM_PC }),
  .out1({ S2562 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1030_ (
  .in1({ S2562, S2561 }),
  .out1({ S2563 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1031_ (
  .in1({ S2563, CU_selMEM_PC }),
  .out1({ S2564 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1256_ (
  .in1({ dataBus[14], CU_selMEM_PC }),
  .out1({ S2565 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1257_ (
  .in1({ S2565, S2578 }),
  .out1({ S2566 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1032_ (
  .in1({ S2566, S2564 }),
  .out1({ S2567 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1033_ (
  .in1({ S2567, S2559 }),
  .out1({ DP_PC_din_14 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1034_ (
  .in1({ DP_INC_1_out_15, S2578 }),
  .out1({ S2568 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1258_ (
  .in1({ DP_IMM1_out_15, CU_selIMM_PC }),
  .out1({ S2569 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_425_ (
  .in1({ S2569 }),
  .out1({ S2570 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1035_ (
  .in1({ S2432, CU_selIMM_PC }),
  .out1({ S2571 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1036_ (
  .in1({ S2571, S2570 }),
  .out1({ S2572 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1037_ (
  .in1({ S2572, CU_selMEM_PC }),
  .out1({ S2573 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1259_ (
  .in1({ dataBus[15], CU_selMEM_PC }),
  .out1({ S2574 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1260_ (
  .in1({ S2574, S2578 }),
  .out1({ S2575 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1038_ (
  .in1({ S2575, S2573 }),
  .out1({ S2576 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1039_ (
  .in1({ S2576, S2568 }),
  .out1({ DP_PC_din_15 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_426_ (
  .in1({ CU_selINC_IN }),
  .out1({ S2593 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1261_ (
  .in1({ CU_selINC_IN, DP_INC2_out_0 }),
  .out1({ S2594 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1262_ (
  .in1({ S2593, dataBus[0] }),
  .out1({ S2595 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1263_ (
  .in1({ S2595, S2594 }),
  .out1({ DP_IN_din_0 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1264_ (
  .in1({ DP_INC2_out_1, CU_selINC_IN }),
  .out1({ S2596 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1265_ (
  .in1({ dataBus[1], S2593 }),
  .out1({ S2597 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1266_ (
  .in1({ S2597, S2596 }),
  .out1({ DP_IN_din_1 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1267_ (
  .in1({ DP_INC2_out_2, CU_selINC_IN }),
  .out1({ S2598 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1268_ (
  .in1({ dataBus[2], S2593 }),
  .out1({ S2599 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1269_ (
  .in1({ S2599, S2598 }),
  .out1({ DP_IN_din_2 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1270_ (
  .in1({ DP_INC2_out_3, CU_selINC_IN }),
  .out1({ S2600 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1271_ (
  .in1({ dataBus[3], S2593 }),
  .out1({ S2601 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1272_ (
  .in1({ S2601, S2600 }),
  .out1({ DP_IN_din_3 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1273_ (
  .in1({ DP_INC2_out_4, CU_selINC_IN }),
  .out1({ S2602 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1274_ (
  .in1({ dataBus[4], S2593 }),
  .out1({ S2603 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1275_ (
  .in1({ S2603, S2602 }),
  .out1({ DP_IN_din_4 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1276_ (
  .in1({ DP_INC2_out_5, CU_selINC_IN }),
  .out1({ S2604 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1277_ (
  .in1({ dataBus[5], S2593 }),
  .out1({ S2605 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1278_ (
  .in1({ S2605, S2604 }),
  .out1({ DP_IN_din_5 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1279_ (
  .in1({ DP_INC2_out_6, CU_selINC_IN }),
  .out1({ S2606 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1280_ (
  .in1({ dataBus[6], S2593 }),
  .out1({ S2607 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1281_ (
  .in1({ S2607, S2606 }),
  .out1({ DP_IN_din_6 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1282_ (
  .in1({ DP_INC2_out_7, CU_selINC_IN }),
  .out1({ S2608 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1283_ (
  .in1({ dataBus[7], S2593 }),
  .out1({ S2609 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1284_ (
  .in1({ S2609, S2608 }),
  .out1({ DP_IN_din_7 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1285_ (
  .in1({ DP_INC2_out_8, CU_selINC_IN }),
  .out1({ S2610 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1286_ (
  .in1({ dataBus[8], S2593 }),
  .out1({ S2611 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1287_ (
  .in1({ S2611, S2610 }),
  .out1({ DP_IN_din_8 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1288_ (
  .in1({ DP_INC2_out_9, CU_selINC_IN }),
  .out1({ S2612 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1289_ (
  .in1({ dataBus[9], S2593 }),
  .out1({ S2613 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1290_ (
  .in1({ S2613, S2612 }),
  .out1({ DP_IN_din_9 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1291_ (
  .in1({ DP_INC2_out_10, CU_selINC_IN }),
  .out1({ S2614 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1292_ (
  .in1({ dataBus[10], S2593 }),
  .out1({ S2615 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1293_ (
  .in1({ S2615, S2614 }),
  .out1({ DP_IN_din_10 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1294_ (
  .in1({ DP_INC2_out_11, CU_selINC_IN }),
  .out1({ S2616 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1295_ (
  .in1({ dataBus[11], S2593 }),
  .out1({ S2617 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1296_ (
  .in1({ S2617, S2616 }),
  .out1({ DP_IN_din_11 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1297_ (
  .in1({ DP_INC2_out_12, CU_selINC_IN }),
  .out1({ S2618 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1298_ (
  .in1({ dataBus[12], S2593 }),
  .out1({ S2619 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1299_ (
  .in1({ S2619, S2618 }),
  .out1({ DP_IN_din_12 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1300_ (
  .in1({ DP_INC2_out_13, CU_selINC_IN }),
  .out1({ S2620 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1301_ (
  .in1({ dataBus[13], S2593 }),
  .out1({ S2621 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1302_ (
  .in1({ S2621, S2620 }),
  .out1({ DP_IN_din_13 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1303_ (
  .in1({ DP_INC2_out_14, CU_selINC_IN }),
  .out1({ S2622 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1304_ (
  .in1({ dataBus[14], S2593 }),
  .out1({ S2623 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1305_ (
  .in1({ S2623, S2622 }),
  .out1({ DP_IN_din_14 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1306_ (
  .in1({ DP_INC2_out_15, CU_selINC_IN }),
  .out1({ S2624 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1307_ (
  .in1({ dataBus[15], S2593 }),
  .out1({ S2625 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1308_ (
  .in1({ S2625, S2624 }),
  .out1({ DP_IN_din_15 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_427_ (
  .in1({ 1'bz }),
  .out1({ S2771 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_428_ (
  .in1({ CU_selIN_MEM }),
  .out1({ S2772 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_429_ (
  .in1({ 1'bz }),
  .out1({ S2773 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_430_ (
  .in1({ 1'bz }),
  .out1({ S2774 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_431_ (
  .in1({ 1'bz }),
  .out1({ S2775 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_432_ (
  .in1({ 1'bz }),
  .out1({ S2776 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_433_ (
  .in1({ 1'bz }),
  .out1({ S2777 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_434_ (
  .in1({ 1'bz }),
  .out1({ S2778 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_435_ (
  .in1({ 1'bz }),
  .out1({ S2779 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_436_ (
  .in1({ 1'bz }),
  .out1({ S2780 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_437_ (
  .in1({ 1'bz }),
  .out1({ S2781 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_438_ (
  .in1({ 1'bz }),
  .out1({ S2782 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_439_ (
  .in1({ 1'bz }),
  .out1({ S2783 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_440_ (
  .in1({ 1'bz }),
  .out1({ S2784 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_441_ (
  .in1({ 1'bz }),
  .out1({ S2785 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_442_ (
  .in1({ 1'bz }),
  .out1({ S2786 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_443_ (
  .in1({ 1'bz }),
  .out1({ S2626 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1040_ (
  .in1({ S2772, DP_IN_dout_0 }),
  .out1({ S2627 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1309_ (
  .in1({ CU_selAC_MEM, DP_AC_dout_0 }),
  .out1({ S2628 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_444_ (
  .in1({ S2628 }),
  .out1({ S2629 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1041_ (
  .in1({ CU_selAC_MEM, S2771 }),
  .out1({ S2630 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1042_ (
  .in1({ S2630, S2629 }),
  .out1({ S2631 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1043_ (
  .in1({ S2631, CU_selPC_MEM }),
  .out1({ S2632 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1310_ (
  .in1({ CU_selPC_MEM, DP_INC_1_out_0 }),
  .out1({ S2633 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1311_ (
  .in1({ S2633, S2772 }),
  .out1({ S2634 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1044_ (
  .in1({ S2634, S2632 }),
  .out1({ S2635 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1045_ (
  .in1({ S2635, S2627 }),
  .out1({ dataBus[0] })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1046_ (
  .in1({ DP_IN_dout_1, S2772 }),
  .out1({ S2636 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1312_ (
  .in1({ DP_AC_dout_1, CU_selAC_MEM }),
  .out1({ S2637 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_445_ (
  .in1({ S2637 }),
  .out1({ S2638 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1047_ (
  .in1({ S2773, CU_selAC_MEM }),
  .out1({ S2639 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1048_ (
  .in1({ S2639, S2638 }),
  .out1({ S2640 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1049_ (
  .in1({ S2640, CU_selPC_MEM }),
  .out1({ S2641 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1313_ (
  .in1({ DP_INC_1_out_1, CU_selPC_MEM }),
  .out1({ S2642 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1314_ (
  .in1({ S2642, S2772 }),
  .out1({ S2643 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1050_ (
  .in1({ S2643, S2641 }),
  .out1({ S2644 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1051_ (
  .in1({ S2644, S2636 }),
  .out1({ dataBus[1] })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1052_ (
  .in1({ DP_IN_dout_2, S2772 }),
  .out1({ S2645 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1315_ (
  .in1({ DP_AC_dout_2, CU_selAC_MEM }),
  .out1({ S2646 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_446_ (
  .in1({ S2646 }),
  .out1({ S2647 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1053_ (
  .in1({ S2774, CU_selAC_MEM }),
  .out1({ S2648 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1054_ (
  .in1({ S2648, S2647 }),
  .out1({ S2649 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1055_ (
  .in1({ S2649, CU_selPC_MEM }),
  .out1({ S2650 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1316_ (
  .in1({ DP_INC_1_out_2, CU_selPC_MEM }),
  .out1({ S2651 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1317_ (
  .in1({ S2651, S2772 }),
  .out1({ S2652 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1056_ (
  .in1({ S2652, S2650 }),
  .out1({ S2653 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1057_ (
  .in1({ S2653, S2645 }),
  .out1({ dataBus[2] })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1058_ (
  .in1({ DP_IN_dout_3, S2772 }),
  .out1({ S2654 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1318_ (
  .in1({ DP_AC_dout_3, CU_selAC_MEM }),
  .out1({ S2655 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_447_ (
  .in1({ S2655 }),
  .out1({ S2656 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1059_ (
  .in1({ S2775, CU_selAC_MEM }),
  .out1({ S2657 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1060_ (
  .in1({ S2657, S2656 }),
  .out1({ S2658 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1061_ (
  .in1({ S2658, CU_selPC_MEM }),
  .out1({ S2659 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1319_ (
  .in1({ DP_INC_1_out_3, CU_selPC_MEM }),
  .out1({ S2660 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1320_ (
  .in1({ S2660, S2772 }),
  .out1({ S2661 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1062_ (
  .in1({ S2661, S2659 }),
  .out1({ S2662 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1063_ (
  .in1({ S2662, S2654 }),
  .out1({ dataBus[3] })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1064_ (
  .in1({ DP_IN_dout_4, S2772 }),
  .out1({ S2663 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1321_ (
  .in1({ DP_AC_dout_4, CU_selAC_MEM }),
  .out1({ S2664 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_448_ (
  .in1({ S2664 }),
  .out1({ S2665 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1065_ (
  .in1({ S2776, CU_selAC_MEM }),
  .out1({ S2666 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1066_ (
  .in1({ S2666, S2665 }),
  .out1({ S2667 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1067_ (
  .in1({ S2667, CU_selPC_MEM }),
  .out1({ S2668 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1322_ (
  .in1({ DP_INC_1_out_4, CU_selPC_MEM }),
  .out1({ S2669 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1323_ (
  .in1({ S2669, S2772 }),
  .out1({ S2670 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1068_ (
  .in1({ S2670, S2668 }),
  .out1({ S2671 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1069_ (
  .in1({ S2671, S2663 }),
  .out1({ dataBus[4] })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1070_ (
  .in1({ DP_IN_dout_5, S2772 }),
  .out1({ S2672 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1324_ (
  .in1({ DP_AC_dout_5, CU_selAC_MEM }),
  .out1({ S2673 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_449_ (
  .in1({ S2673 }),
  .out1({ S2674 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1071_ (
  .in1({ S2777, CU_selAC_MEM }),
  .out1({ S2675 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1072_ (
  .in1({ S2675, S2674 }),
  .out1({ S2676 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1073_ (
  .in1({ S2676, CU_selPC_MEM }),
  .out1({ S2677 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1325_ (
  .in1({ DP_INC_1_out_5, CU_selPC_MEM }),
  .out1({ S2678 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1326_ (
  .in1({ S2678, S2772 }),
  .out1({ S2679 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1074_ (
  .in1({ S2679, S2677 }),
  .out1({ S2680 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1075_ (
  .in1({ S2680, S2672 }),
  .out1({ dataBus[5] })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1076_ (
  .in1({ DP_IN_dout_6, S2772 }),
  .out1({ S2681 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1327_ (
  .in1({ DP_AC_dout_6, CU_selAC_MEM }),
  .out1({ S2682 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_450_ (
  .in1({ S2682 }),
  .out1({ S2683 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1077_ (
  .in1({ S2778, CU_selAC_MEM }),
  .out1({ S2684 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1078_ (
  .in1({ S2684, S2683 }),
  .out1({ S2685 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1079_ (
  .in1({ S2685, CU_selPC_MEM }),
  .out1({ S2686 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1328_ (
  .in1({ DP_INC_1_out_6, CU_selPC_MEM }),
  .out1({ S2687 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1329_ (
  .in1({ S2687, S2772 }),
  .out1({ S2688 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1080_ (
  .in1({ S2688, S2686 }),
  .out1({ S2689 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1081_ (
  .in1({ S2689, S2681 }),
  .out1({ dataBus[6] })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1082_ (
  .in1({ DP_IN_dout_7, S2772 }),
  .out1({ S2690 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1330_ (
  .in1({ DP_AC_dout_7, CU_selAC_MEM }),
  .out1({ S2691 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_451_ (
  .in1({ S2691 }),
  .out1({ S2692 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1083_ (
  .in1({ S2779, CU_selAC_MEM }),
  .out1({ S2693 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1084_ (
  .in1({ S2693, S2692 }),
  .out1({ S2694 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1085_ (
  .in1({ S2694, CU_selPC_MEM }),
  .out1({ S2695 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1331_ (
  .in1({ DP_INC_1_out_7, CU_selPC_MEM }),
  .out1({ S2696 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1332_ (
  .in1({ S2696, S2772 }),
  .out1({ S2697 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1086_ (
  .in1({ S2697, S2695 }),
  .out1({ S2698 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1087_ (
  .in1({ S2698, S2690 }),
  .out1({ dataBus[7] })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1088_ (
  .in1({ DP_IN_dout_8, S2772 }),
  .out1({ S2699 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1333_ (
  .in1({ DP_AC_dout_8, CU_selAC_MEM }),
  .out1({ S2700 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_452_ (
  .in1({ S2700 }),
  .out1({ S2701 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1089_ (
  .in1({ S2780, CU_selAC_MEM }),
  .out1({ S2702 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1090_ (
  .in1({ S2702, S2701 }),
  .out1({ S2703 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1091_ (
  .in1({ S2703, CU_selPC_MEM }),
  .out1({ S2704 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1334_ (
  .in1({ DP_INC_1_out_8, CU_selPC_MEM }),
  .out1({ S2705 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1335_ (
  .in1({ S2705, S2772 }),
  .out1({ S2706 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1092_ (
  .in1({ S2706, S2704 }),
  .out1({ S2707 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1093_ (
  .in1({ S2707, S2699 }),
  .out1({ dataBus[8] })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1094_ (
  .in1({ DP_IN_dout_9, S2772 }),
  .out1({ S2708 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1336_ (
  .in1({ DP_AC_dout_9, CU_selAC_MEM }),
  .out1({ S2709 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_453_ (
  .in1({ S2709 }),
  .out1({ S2710 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1095_ (
  .in1({ S2781, CU_selAC_MEM }),
  .out1({ S2711 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1096_ (
  .in1({ S2711, S2710 }),
  .out1({ S2712 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1097_ (
  .in1({ S2712, CU_selPC_MEM }),
  .out1({ S2713 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1337_ (
  .in1({ DP_INC_1_out_9, CU_selPC_MEM }),
  .out1({ S2714 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1338_ (
  .in1({ S2714, S2772 }),
  .out1({ S2715 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1098_ (
  .in1({ S2715, S2713 }),
  .out1({ S2716 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1099_ (
  .in1({ S2716, S2708 }),
  .out1({ dataBus[9] })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1100_ (
  .in1({ DP_IN_dout_10, S2772 }),
  .out1({ S2717 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1339_ (
  .in1({ DP_AC_dout_10, CU_selAC_MEM }),
  .out1({ S2718 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_454_ (
  .in1({ S2718 }),
  .out1({ S2719 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1101_ (
  .in1({ S2782, CU_selAC_MEM }),
  .out1({ S2720 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1102_ (
  .in1({ S2720, S2719 }),
  .out1({ S2721 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1103_ (
  .in1({ S2721, CU_selPC_MEM }),
  .out1({ S2722 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1340_ (
  .in1({ DP_INC_1_out_10, CU_selPC_MEM }),
  .out1({ S2723 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1341_ (
  .in1({ S2723, S2772 }),
  .out1({ S2724 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1104_ (
  .in1({ S2724, S2722 }),
  .out1({ S2725 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1105_ (
  .in1({ S2725, S2717 }),
  .out1({ dataBus[10] })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1106_ (
  .in1({ DP_IN_dout_11, S2772 }),
  .out1({ S2726 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1342_ (
  .in1({ DP_AC_dout_11, CU_selAC_MEM }),
  .out1({ S2727 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_455_ (
  .in1({ S2727 }),
  .out1({ S2728 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1107_ (
  .in1({ S2783, CU_selAC_MEM }),
  .out1({ S2729 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1108_ (
  .in1({ S2729, S2728 }),
  .out1({ S2730 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1109_ (
  .in1({ S2730, CU_selPC_MEM }),
  .out1({ S2731 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1343_ (
  .in1({ DP_INC_1_out_11, CU_selPC_MEM }),
  .out1({ S2732 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1344_ (
  .in1({ S2732, S2772 }),
  .out1({ S2733 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1110_ (
  .in1({ S2733, S2731 }),
  .out1({ S2734 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1111_ (
  .in1({ S2734, S2726 }),
  .out1({ dataBus[11] })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1112_ (
  .in1({ DP_IN_dout_12, S2772 }),
  .out1({ S2735 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1345_ (
  .in1({ DP_AC_dout_12, CU_selAC_MEM }),
  .out1({ S2736 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_456_ (
  .in1({ S2736 }),
  .out1({ S2737 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1113_ (
  .in1({ S2784, CU_selAC_MEM }),
  .out1({ S2738 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1114_ (
  .in1({ S2738, S2737 }),
  .out1({ S2739 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1115_ (
  .in1({ S2739, CU_selPC_MEM }),
  .out1({ S2740 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1346_ (
  .in1({ DP_INC_1_out_12, CU_selPC_MEM }),
  .out1({ S2741 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1347_ (
  .in1({ S2741, S2772 }),
  .out1({ S2742 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1116_ (
  .in1({ S2742, S2740 }),
  .out1({ S2743 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1117_ (
  .in1({ S2743, S2735 }),
  .out1({ dataBus[12] })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1118_ (
  .in1({ DP_IN_dout_13, S2772 }),
  .out1({ S2744 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1348_ (
  .in1({ DP_AC_dout_13, CU_selAC_MEM }),
  .out1({ S2745 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_457_ (
  .in1({ S2745 }),
  .out1({ S2746 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1119_ (
  .in1({ S2785, CU_selAC_MEM }),
  .out1({ S2747 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1120_ (
  .in1({ S2747, S2746 }),
  .out1({ S2748 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1121_ (
  .in1({ S2748, CU_selPC_MEM }),
  .out1({ S2749 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1349_ (
  .in1({ DP_INC_1_out_13, CU_selPC_MEM }),
  .out1({ S2750 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1350_ (
  .in1({ S2750, S2772 }),
  .out1({ S2751 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1122_ (
  .in1({ S2751, S2749 }),
  .out1({ S2752 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1123_ (
  .in1({ S2752, S2744 }),
  .out1({ dataBus[13] })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1124_ (
  .in1({ DP_IN_dout_14, S2772 }),
  .out1({ S2753 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1351_ (
  .in1({ DP_AC_dout_14, CU_selAC_MEM }),
  .out1({ S2754 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_458_ (
  .in1({ S2754 }),
  .out1({ S2755 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1125_ (
  .in1({ S2786, CU_selAC_MEM }),
  .out1({ S2756 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1126_ (
  .in1({ S2756, S2755 }),
  .out1({ S2757 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1127_ (
  .in1({ S2757, CU_selPC_MEM }),
  .out1({ S2758 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1352_ (
  .in1({ DP_INC_1_out_14, CU_selPC_MEM }),
  .out1({ S2759 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1353_ (
  .in1({ S2759, S2772 }),
  .out1({ S2760 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1128_ (
  .in1({ S2760, S2758 }),
  .out1({ S2761 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1129_ (
  .in1({ S2761, S2753 }),
  .out1({ dataBus[14] })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1130_ (
  .in1({ DP_IN_dout_15, S2772 }),
  .out1({ S2762 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1354_ (
  .in1({ DP_AC_dout_15, CU_selAC_MEM }),
  .out1({ S2763 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_459_ (
  .in1({ S2763 }),
  .out1({ S2764 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1131_ (
  .in1({ S2626, CU_selAC_MEM }),
  .out1({ S2765 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1132_ (
  .in1({ S2765, S2764 }),
  .out1({ S2766 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1133_ (
  .in1({ S2766, CU_selPC_MEM }),
  .out1({ S2767 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1355_ (
  .in1({ DP_INC_1_out_15, CU_selPC_MEM }),
  .out1({ S2768 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1356_ (
  .in1({ S2768, S2772 }),
  .out1({ S2769 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1134_ (
  .in1({ S2769, S2767 }),
  .out1({ S2770 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1135_ (
  .in1({ S2770, S2762 }),
  .out1({ dataBus[15] })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_460_ (
  .in1({ 1'bz }),
  .out1({ S2932 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_461_ (
  .in1({ CU_selIN_ADR }),
  .out1({ S2933 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_462_ (
  .in1({ 1'bz }),
  .out1({ S2934 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_463_ (
  .in1({ 1'bz }),
  .out1({ S2935 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_464_ (
  .in1({ 1'bz }),
  .out1({ S2936 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_465_ (
  .in1({ 1'bz }),
  .out1({ S2937 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_466_ (
  .in1({ 1'bz }),
  .out1({ S2938 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_467_ (
  .in1({ 1'bz }),
  .out1({ S2939 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_468_ (
  .in1({ 1'bz }),
  .out1({ S2940 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_469_ (
  .in1({ 1'bz }),
  .out1({ S2941 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_470_ (
  .in1({ 1'bz }),
  .out1({ S2942 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_471_ (
  .in1({ 1'bz }),
  .out1({ S2943 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_472_ (
  .in1({ 1'bz }),
  .out1({ S2944 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_473_ (
  .in1({ 1'bz }),
  .out1({ S2945 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_474_ (
  .in1({ 1'bz }),
  .out1({ S2946 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_475_ (
  .in1({ 1'bz }),
  .out1({ S2947 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_476_ (
  .in1({ 1'bz }),
  .out1({ S2787 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1136_ (
  .in1({ S2933, DP_IN_dout_0 }),
  .out1({ S2788 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1357_ (
  .in1({ CU_ldIR, DP_INC_1_in_0 }),
  .out1({ S2789 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_477_ (
  .in1({ S2789 }),
  .out1({ S2790 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1137_ (
  .in1({ CU_ldIR, S2932 }),
  .out1({ S2791 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1138_ (
  .in1({ S2791, S2790 }),
  .out1({ S2792 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1139_ (
  .in1({ S2792, CU_selIR_ADR }),
  .out1({ S2793 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1358_ (
  .in1({ CU_selIR_ADR, DP_IMM1_out_0 }),
  .out1({ S2794 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1359_ (
  .in1({ S2794, S2933 }),
  .out1({ S2795 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1140_ (
  .in1({ S2795, S2793 }),
  .out1({ S2796 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1141_ (
  .in1({ S2796, S2788 }),
  .out1({ DP_addrBus_0 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1142_ (
  .in1({ DP_IN_dout_1, S2933 }),
  .out1({ S2797 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1360_ (
  .in1({ DP_INC_1_in_1, CU_ldIR }),
  .out1({ S2798 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_478_ (
  .in1({ S2798 }),
  .out1({ S2799 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1143_ (
  .in1({ S2934, CU_ldIR }),
  .out1({ S2800 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1144_ (
  .in1({ S2800, S2799 }),
  .out1({ S2801 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1145_ (
  .in1({ S2801, CU_selIR_ADR }),
  .out1({ S2802 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1361_ (
  .in1({ DP_IMM1_out_1, CU_selIR_ADR }),
  .out1({ S2803 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1362_ (
  .in1({ S2803, S2933 }),
  .out1({ S2804 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1146_ (
  .in1({ S2804, S2802 }),
  .out1({ S2805 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1147_ (
  .in1({ S2805, S2797 }),
  .out1({ DP_addrBus_1 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1148_ (
  .in1({ DP_IN_dout_2, S2933 }),
  .out1({ S2806 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1363_ (
  .in1({ DP_INC_1_in_2, CU_ldIR }),
  .out1({ S2807 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_479_ (
  .in1({ S2807 }),
  .out1({ S2808 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1149_ (
  .in1({ S2935, CU_ldIR }),
  .out1({ S2809 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1150_ (
  .in1({ S2809, S2808 }),
  .out1({ S2810 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1151_ (
  .in1({ S2810, CU_selIR_ADR }),
  .out1({ S2811 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1364_ (
  .in1({ DP_IMM1_out_2, CU_selIR_ADR }),
  .out1({ S2812 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1365_ (
  .in1({ S2812, S2933 }),
  .out1({ S2813 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1152_ (
  .in1({ S2813, S2811 }),
  .out1({ S2814 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1153_ (
  .in1({ S2814, S2806 }),
  .out1({ DP_addrBus_2 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1154_ (
  .in1({ DP_IN_dout_3, S2933 }),
  .out1({ S2815 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1366_ (
  .in1({ DP_INC_1_in_3, CU_ldIR }),
  .out1({ S2816 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_480_ (
  .in1({ S2816 }),
  .out1({ S2817 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1155_ (
  .in1({ S2936, CU_ldIR }),
  .out1({ S2818 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1156_ (
  .in1({ S2818, S2817 }),
  .out1({ S2819 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1157_ (
  .in1({ S2819, CU_selIR_ADR }),
  .out1({ S2820 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1367_ (
  .in1({ DP_IMM1_out_3, CU_selIR_ADR }),
  .out1({ S2821 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1368_ (
  .in1({ S2821, S2933 }),
  .out1({ S2822 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1158_ (
  .in1({ S2822, S2820 }),
  .out1({ S2823 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1159_ (
  .in1({ S2823, S2815 }),
  .out1({ DP_addrBus_3 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1160_ (
  .in1({ DP_IN_dout_4, S2933 }),
  .out1({ S2824 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1369_ (
  .in1({ DP_INC_1_in_4, CU_ldIR }),
  .out1({ S2825 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_481_ (
  .in1({ S2825 }),
  .out1({ S2826 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1161_ (
  .in1({ S2937, CU_ldIR }),
  .out1({ S2827 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1162_ (
  .in1({ S2827, S2826 }),
  .out1({ S2828 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1163_ (
  .in1({ S2828, CU_selIR_ADR }),
  .out1({ S2829 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1370_ (
  .in1({ DP_IMM1_out_4, CU_selIR_ADR }),
  .out1({ S2830 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1371_ (
  .in1({ S2830, S2933 }),
  .out1({ S2831 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1164_ (
  .in1({ S2831, S2829 }),
  .out1({ S2832 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1165_ (
  .in1({ S2832, S2824 }),
  .out1({ DP_addrBus_4 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1166_ (
  .in1({ DP_IN_dout_5, S2933 }),
  .out1({ S2833 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1372_ (
  .in1({ DP_INC_1_in_5, CU_ldIR }),
  .out1({ S2834 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_482_ (
  .in1({ S2834 }),
  .out1({ S2835 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1167_ (
  .in1({ S2938, CU_ldIR }),
  .out1({ S2836 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1168_ (
  .in1({ S2836, S2835 }),
  .out1({ S2837 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1169_ (
  .in1({ S2837, CU_selIR_ADR }),
  .out1({ S2838 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1373_ (
  .in1({ DP_IMM1_out_5, CU_selIR_ADR }),
  .out1({ S2839 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1374_ (
  .in1({ S2839, S2933 }),
  .out1({ S2840 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1170_ (
  .in1({ S2840, S2838 }),
  .out1({ S2841 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1171_ (
  .in1({ S2841, S2833 }),
  .out1({ DP_addrBus_5 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1172_ (
  .in1({ DP_IN_dout_6, S2933 }),
  .out1({ S2842 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1375_ (
  .in1({ DP_INC_1_in_6, CU_ldIR }),
  .out1({ S2843 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_483_ (
  .in1({ S2843 }),
  .out1({ S2844 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1173_ (
  .in1({ S2939, CU_ldIR }),
  .out1({ S2845 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1174_ (
  .in1({ S2845, S2844 }),
  .out1({ S2846 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1175_ (
  .in1({ S2846, CU_selIR_ADR }),
  .out1({ S2847 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1376_ (
  .in1({ DP_IMM1_out_6, CU_selIR_ADR }),
  .out1({ S2848 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1377_ (
  .in1({ S2848, S2933 }),
  .out1({ S2849 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1176_ (
  .in1({ S2849, S2847 }),
  .out1({ S2850 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1177_ (
  .in1({ S2850, S2842 }),
  .out1({ DP_addrBus_6 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1178_ (
  .in1({ DP_IN_dout_7, S2933 }),
  .out1({ S2851 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1378_ (
  .in1({ DP_INC_1_in_7, CU_ldIR }),
  .out1({ S2852 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_484_ (
  .in1({ S2852 }),
  .out1({ S2853 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1179_ (
  .in1({ S2940, CU_ldIR }),
  .out1({ S2854 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1180_ (
  .in1({ S2854, S2853 }),
  .out1({ S2855 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1181_ (
  .in1({ S2855, CU_selIR_ADR }),
  .out1({ S2856 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1379_ (
  .in1({ DP_IMM1_out_7, CU_selIR_ADR }),
  .out1({ S2857 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1380_ (
  .in1({ S2857, S2933 }),
  .out1({ S2858 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1182_ (
  .in1({ S2858, S2856 }),
  .out1({ S2859 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1183_ (
  .in1({ S2859, S2851 }),
  .out1({ DP_addrBus_7 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1184_ (
  .in1({ DP_IN_dout_8, S2933 }),
  .out1({ S2860 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1381_ (
  .in1({ DP_INC_1_in_8, CU_ldIR }),
  .out1({ S2861 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_485_ (
  .in1({ S2861 }),
  .out1({ S2862 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1185_ (
  .in1({ S2941, CU_ldIR }),
  .out1({ S2863 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1186_ (
  .in1({ S2863, S2862 }),
  .out1({ S2864 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1187_ (
  .in1({ S2864, CU_selIR_ADR }),
  .out1({ S2865 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1382_ (
  .in1({ DP_IMM1_out_8, CU_selIR_ADR }),
  .out1({ S2866 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1383_ (
  .in1({ S2866, S2933 }),
  .out1({ S2867 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1188_ (
  .in1({ S2867, S2865 }),
  .out1({ S2868 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1189_ (
  .in1({ S2868, S2860 }),
  .out1({ DP_addrBus_8 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1190_ (
  .in1({ DP_IN_dout_9, S2933 }),
  .out1({ S2869 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1384_ (
  .in1({ DP_INC_1_in_9, CU_ldIR }),
  .out1({ S2870 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_486_ (
  .in1({ S2870 }),
  .out1({ S2871 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1191_ (
  .in1({ S2942, CU_ldIR }),
  .out1({ S2872 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1192_ (
  .in1({ S2872, S2871 }),
  .out1({ S2873 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1193_ (
  .in1({ S2873, CU_selIR_ADR }),
  .out1({ S2874 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1385_ (
  .in1({ DP_IMM1_out_9, CU_selIR_ADR }),
  .out1({ S2875 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1386_ (
  .in1({ S2875, S2933 }),
  .out1({ S2876 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1194_ (
  .in1({ S2876, S2874 }),
  .out1({ S2877 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1195_ (
  .in1({ S2877, S2869 }),
  .out1({ DP_addrBus_9 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1196_ (
  .in1({ DP_IN_dout_10, S2933 }),
  .out1({ S2878 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1387_ (
  .in1({ DP_INC_1_in_10, CU_ldIR }),
  .out1({ S2879 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_487_ (
  .in1({ S2879 }),
  .out1({ S2880 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1197_ (
  .in1({ S2943, CU_ldIR }),
  .out1({ S2881 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1198_ (
  .in1({ S2881, S2880 }),
  .out1({ S2882 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1199_ (
  .in1({ S2882, CU_selIR_ADR }),
  .out1({ S2883 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1388_ (
  .in1({ DP_IMM1_out_10, CU_selIR_ADR }),
  .out1({ S2884 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1389_ (
  .in1({ S2884, S2933 }),
  .out1({ S2885 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1200_ (
  .in1({ S2885, S2883 }),
  .out1({ S2886 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1201_ (
  .in1({ S2886, S2878 }),
  .out1({ DP_addrBus_10 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1202_ (
  .in1({ DP_IN_dout_11, S2933 }),
  .out1({ S2887 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1390_ (
  .in1({ DP_INC_1_in_11, CU_ldIR }),
  .out1({ S2888 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_488_ (
  .in1({ S2888 }),
  .out1({ S2889 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1203_ (
  .in1({ S2944, CU_ldIR }),
  .out1({ S2890 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1204_ (
  .in1({ S2890, S2889 }),
  .out1({ S2891 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1205_ (
  .in1({ S2891, CU_selIR_ADR }),
  .out1({ S2892 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1391_ (
  .in1({ DP_IMM1_out_11, CU_selIR_ADR }),
  .out1({ S2893 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1392_ (
  .in1({ S2893, S2933 }),
  .out1({ S2894 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1206_ (
  .in1({ S2894, S2892 }),
  .out1({ S2895 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1207_ (
  .in1({ S2895, S2887 }),
  .out1({ DP_addrBus_11 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1208_ (
  .in1({ DP_IN_dout_12, S2933 }),
  .out1({ S2896 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1393_ (
  .in1({ DP_INC_1_in_12, CU_ldIR }),
  .out1({ S2897 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_489_ (
  .in1({ S2897 }),
  .out1({ S2898 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1209_ (
  .in1({ S2945, CU_ldIR }),
  .out1({ S2899 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1210_ (
  .in1({ S2899, S2898 }),
  .out1({ S2900 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1211_ (
  .in1({ S2900, CU_selIR_ADR }),
  .out1({ S2901 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1394_ (
  .in1({ DP_IMM1_out_12, CU_selIR_ADR }),
  .out1({ S2902 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1395_ (
  .in1({ S2902, S2933 }),
  .out1({ S2903 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1212_ (
  .in1({ S2903, S2901 }),
  .out1({ S2904 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1213_ (
  .in1({ S2904, S2896 }),
  .out1({ DP_addrBus_12 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1214_ (
  .in1({ DP_IN_dout_13, S2933 }),
  .out1({ S2905 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1396_ (
  .in1({ DP_INC_1_in_13, CU_ldIR }),
  .out1({ S2906 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_490_ (
  .in1({ S2906 }),
  .out1({ S2907 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1215_ (
  .in1({ S2946, CU_ldIR }),
  .out1({ S2908 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1216_ (
  .in1({ S2908, S2907 }),
  .out1({ S2909 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1217_ (
  .in1({ S2909, CU_selIR_ADR }),
  .out1({ S2910 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1397_ (
  .in1({ DP_IMM1_out_13, CU_selIR_ADR }),
  .out1({ S2911 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1398_ (
  .in1({ S2911, S2933 }),
  .out1({ S2912 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1218_ (
  .in1({ S2912, S2910 }),
  .out1({ S2913 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1219_ (
  .in1({ S2913, S2905 }),
  .out1({ DP_addrBus_13 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1220_ (
  .in1({ DP_IN_dout_14, S2933 }),
  .out1({ S2914 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1399_ (
  .in1({ DP_INC_1_in_14, CU_ldIR }),
  .out1({ S2915 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_491_ (
  .in1({ S2915 }),
  .out1({ S2916 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1221_ (
  .in1({ S2947, CU_ldIR }),
  .out1({ S2917 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1222_ (
  .in1({ S2917, S2916 }),
  .out1({ S2918 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1223_ (
  .in1({ S2918, CU_selIR_ADR }),
  .out1({ S2919 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1400_ (
  .in1({ DP_IMM1_out_14, CU_selIR_ADR }),
  .out1({ S2920 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1401_ (
  .in1({ S2920, S2933 }),
  .out1({ S2921 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1224_ (
  .in1({ S2921, S2919 }),
  .out1({ S2922 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1225_ (
  .in1({ S2922, S2914 }),
  .out1({ DP_addrBus_14 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1226_ (
  .in1({ DP_IN_dout_15, S2933 }),
  .out1({ S2923 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1402_ (
  .in1({ DP_INC_1_in_15, CU_ldIR }),
  .out1({ S2924 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_492_ (
  .in1({ S2924 }),
  .out1({ S2925 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1227_ (
  .in1({ S2787, CU_ldIR }),
  .out1({ S2926 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1228_ (
  .in1({ S2926, S2925 }),
  .out1({ S2927 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1229_ (
  .in1({ S2927, CU_selIR_ADR }),
  .out1({ S2928 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1403_ (
  .in1({ DP_IMM1_out_15, CU_selIR_ADR }),
  .out1({ S2929 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1404_ (
  .in1({ S2929, S2933 }),
  .out1({ S2930 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1230_ (
  .in1({ S2930, S2928 }),
  .out1({ S2931 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1231_ (
  .in1({ S2931, S2923 }),
  .out1({ DP_addrBus_15 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_493_ (
  .in1({ CU_selIMM_LGU }),
  .out1({ S2948 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1405_ (
  .in1({ CU_selIMM_LGU, DP_IMM1_out_0 }),
  .out1({ S2949 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1406_ (
  .in1({ S2948, dataBus[0] }),
  .out1({ S2950 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1407_ (
  .in1({ S2950, S2949 }),
  .out1({ DP_LGU1_in1_0 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1408_ (
  .in1({ DP_IMM1_out_1, CU_selIMM_LGU }),
  .out1({ S2951 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1409_ (
  .in1({ dataBus[1], S2948 }),
  .out1({ S2952 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1410_ (
  .in1({ S2952, S2951 }),
  .out1({ DP_LGU1_in1_1 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1411_ (
  .in1({ DP_IMM1_out_2, CU_selIMM_LGU }),
  .out1({ S2953 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1412_ (
  .in1({ dataBus[2], S2948 }),
  .out1({ S2954 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1413_ (
  .in1({ S2954, S2953 }),
  .out1({ DP_LGU1_in1_2 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1414_ (
  .in1({ DP_IMM1_out_3, CU_selIMM_LGU }),
  .out1({ S2955 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1415_ (
  .in1({ dataBus[3], S2948 }),
  .out1({ S2956 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1416_ (
  .in1({ S2956, S2955 }),
  .out1({ DP_LGU1_in1_3 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1417_ (
  .in1({ DP_IMM1_out_4, CU_selIMM_LGU }),
  .out1({ S2957 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1418_ (
  .in1({ dataBus[4], S2948 }),
  .out1({ S2958 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1419_ (
  .in1({ S2958, S2957 }),
  .out1({ DP_LGU1_in1_4 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1420_ (
  .in1({ DP_IMM1_out_5, CU_selIMM_LGU }),
  .out1({ S2959 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1421_ (
  .in1({ dataBus[5], S2948 }),
  .out1({ S2960 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1422_ (
  .in1({ S2960, S2959 }),
  .out1({ DP_LGU1_in1_5 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1423_ (
  .in1({ DP_IMM1_out_6, CU_selIMM_LGU }),
  .out1({ S2961 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1424_ (
  .in1({ dataBus[6], S2948 }),
  .out1({ S2962 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1425_ (
  .in1({ S2962, S2961 }),
  .out1({ DP_LGU1_in1_6 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1426_ (
  .in1({ DP_IMM1_out_7, CU_selIMM_LGU }),
  .out1({ S2963 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1427_ (
  .in1({ dataBus[7], S2948 }),
  .out1({ S2964 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1428_ (
  .in1({ S2964, S2963 }),
  .out1({ DP_LGU1_in1_7 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1429_ (
  .in1({ DP_IMM1_out_8, CU_selIMM_LGU }),
  .out1({ S2965 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1430_ (
  .in1({ dataBus[8], S2948 }),
  .out1({ S2966 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1431_ (
  .in1({ S2966, S2965 }),
  .out1({ DP_LGU1_in1_8 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1432_ (
  .in1({ DP_IMM1_out_9, CU_selIMM_LGU }),
  .out1({ S2967 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1433_ (
  .in1({ dataBus[9], S2948 }),
  .out1({ S2968 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1434_ (
  .in1({ S2968, S2967 }),
  .out1({ DP_LGU1_in1_9 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1435_ (
  .in1({ DP_IMM1_out_10, CU_selIMM_LGU }),
  .out1({ S2969 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1436_ (
  .in1({ dataBus[10], S2948 }),
  .out1({ S2970 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1437_ (
  .in1({ S2970, S2969 }),
  .out1({ DP_LGU1_in1_10 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1438_ (
  .in1({ DP_IMM1_out_11, CU_selIMM_LGU }),
  .out1({ S2971 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1439_ (
  .in1({ dataBus[11], S2948 }),
  .out1({ S2972 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1440_ (
  .in1({ S2972, S2971 }),
  .out1({ DP_LGU1_in1_11 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1441_ (
  .in1({ DP_IMM1_out_12, CU_selIMM_LGU }),
  .out1({ S2973 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1442_ (
  .in1({ dataBus[12], S2948 }),
  .out1({ S2974 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1443_ (
  .in1({ S2974, S2973 }),
  .out1({ DP_LGU1_in1_12 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1444_ (
  .in1({ DP_IMM1_out_13, CU_selIMM_LGU }),
  .out1({ S2975 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1445_ (
  .in1({ dataBus[13], S2948 }),
  .out1({ S2976 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1446_ (
  .in1({ S2976, S2975 }),
  .out1({ DP_LGU1_in1_13 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1447_ (
  .in1({ DP_IMM1_out_14, CU_selIMM_LGU }),
  .out1({ S2977 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1448_ (
  .in1({ dataBus[14], S2948 }),
  .out1({ S2978 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1449_ (
  .in1({ S2978, S2977 }),
  .out1({ DP_LGU1_in1_14 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1450_ (
  .in1({ DP_IMM1_out_15, CU_selIMM_LGU }),
  .out1({ S2979 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1451_ (
  .in1({ dataBus[15], S2948 }),
  .out1({ S2980 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1452_ (
  .in1({ S2980, S2979 }),
  .out1({ DP_LGU1_in1_15 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_494_ (
  .in1({ CU_sel1_ARU }),
  .out1({ S2981 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1453_ (
  .in1({ CU_sel1_ARU, S3 }),
  .out1({ S2982 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1454_ (
  .in1({ S2981, DP_LGU1_in1_0 }),
  .out1({ S2983 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1455_ (
  .in1({ S2983, S2982 }),
  .out1({ DP_ARU1_in1_0 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1456_ (
  .in1({ S21, CU_sel1_ARU }),
  .out1({ S2984 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1457_ (
  .in1({ DP_LGU1_in1_1, S2981 }),
  .out1({ S2985 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1458_ (
  .in1({ S2985, S2984 }),
  .out1({ DP_ARU1_in1_1 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1459_ (
  .in1({ S22, CU_sel1_ARU }),
  .out1({ S2986 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1460_ (
  .in1({ DP_LGU1_in1_2, S2981 }),
  .out1({ S2987 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1461_ (
  .in1({ S2987, S2986 }),
  .out1({ DP_ARU1_in1_2 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1462_ (
  .in1({ S23, CU_sel1_ARU }),
  .out1({ S2988 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1463_ (
  .in1({ DP_LGU1_in1_3, S2981 }),
  .out1({ S2989 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1464_ (
  .in1({ S2989, S2988 }),
  .out1({ DP_ARU1_in1_3 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1465_ (
  .in1({ S24, CU_sel1_ARU }),
  .out1({ S2990 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1466_ (
  .in1({ DP_LGU1_in1_4, S2981 }),
  .out1({ S2991 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1467_ (
  .in1({ S2991, S2990 }),
  .out1({ DP_ARU1_in1_4 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1468_ (
  .in1({ S25, CU_sel1_ARU }),
  .out1({ S2992 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1469_ (
  .in1({ DP_LGU1_in1_5, S2981 }),
  .out1({ S2993 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1470_ (
  .in1({ S2993, S2992 }),
  .out1({ DP_ARU1_in1_5 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1471_ (
  .in1({ S26, CU_sel1_ARU }),
  .out1({ S2994 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1472_ (
  .in1({ DP_LGU1_in1_6, S2981 }),
  .out1({ S2995 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1473_ (
  .in1({ S2995, S2994 }),
  .out1({ DP_ARU1_in1_6 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1474_ (
  .in1({ S27, CU_sel1_ARU }),
  .out1({ S2996 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1475_ (
  .in1({ DP_LGU1_in1_7, S2981 }),
  .out1({ S2997 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1476_ (
  .in1({ S2997, S2996 }),
  .out1({ DP_ARU1_in1_7 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1477_ (
  .in1({ S28, CU_sel1_ARU }),
  .out1({ S2998 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1478_ (
  .in1({ DP_LGU1_in1_8, S2981 }),
  .out1({ S2999 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1479_ (
  .in1({ S2999, S2998 }),
  .out1({ DP_ARU1_in1_8 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1480_ (
  .in1({ S29, CU_sel1_ARU }),
  .out1({ S3000 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1481_ (
  .in1({ DP_LGU1_in1_9, S2981 }),
  .out1({ S3001 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1482_ (
  .in1({ S3001, S3000 }),
  .out1({ DP_ARU1_in1_9 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1483_ (
  .in1({ S30, CU_sel1_ARU }),
  .out1({ S3002 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1484_ (
  .in1({ DP_LGU1_in1_10, S2981 }),
  .out1({ S3003 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1485_ (
  .in1({ S3003, S3002 }),
  .out1({ DP_ARU1_in1_10 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1486_ (
  .in1({ S31, CU_sel1_ARU }),
  .out1({ S3004 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1487_ (
  .in1({ DP_LGU1_in1_11, S2981 }),
  .out1({ S3005 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1488_ (
  .in1({ S3005, S3004 }),
  .out1({ DP_ARU1_in1_11 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1489_ (
  .in1({ S32, CU_sel1_ARU }),
  .out1({ S3006 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1490_ (
  .in1({ DP_LGU1_in1_12, S2981 }),
  .out1({ S3007 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1491_ (
  .in1({ S3007, S3006 }),
  .out1({ DP_ARU1_in1_12 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1492_ (
  .in1({ S33, CU_sel1_ARU }),
  .out1({ S3008 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1493_ (
  .in1({ DP_LGU1_in1_13, S2981 }),
  .out1({ S3009 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1494_ (
  .in1({ S3009, S3008 }),
  .out1({ DP_ARU1_in1_13 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1495_ (
  .in1({ S34, CU_sel1_ARU }),
  .out1({ S3010 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1496_ (
  .in1({ DP_LGU1_in1_14, S2981 }),
  .out1({ S3011 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1497_ (
  .in1({ S3011, S3010 }),
  .out1({ DP_ARU1_in1_14 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1498_ (
  .in1({ S35, CU_sel1_ARU }),
  .out1({ S3012 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1499_ (
  .in1({ DP_LGU1_in1_15, S2981 }),
  .out1({ S3013 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1500_ (
  .in1({ S3013, S3012 }),
  .out1({ DP_ARU1_in1_15 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_495_ (
  .in1({ CU_selPC_OF }),
  .out1({ S3014 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1501_ (
  .in1({ CU_selPC_OF, DP_INC_1_in_12 }),
  .out1({ S3015 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1502_ (
  .in1({ S3014, DP_IMM1_out_0 }),
  .out1({ S3016 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1503_ (
  .in1({ S3016, S3015 }),
  .out1({ DP_OF_din_0 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1504_ (
  .in1({ DP_INC_1_in_13, CU_selPC_OF }),
  .out1({ S3017 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1505_ (
  .in1({ DP_IMM1_out_1, S3014 }),
  .out1({ S3018 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1506_ (
  .in1({ S3018, S3017 }),
  .out1({ DP_OF_din_1 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1507_ (
  .in1({ DP_INC_1_in_14, CU_selPC_OF }),
  .out1({ S3019 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1508_ (
  .in1({ DP_IMM1_out_2, S3014 }),
  .out1({ S3020 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1509_ (
  .in1({ S3020, S3019 }),
  .out1({ DP_OF_din_2 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1510_ (
  .in1({ DP_INC_1_in_15, CU_selPC_OF }),
  .out1({ S3021 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1511_ (
  .in1({ DP_IMM1_out_3, S3014 }),
  .out1({ S3022 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1512_ (
  .in1({ S3022, S3021 }),
  .out1({ DP_OF_din_3 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_496_ (
  .in1({ CU_INC2 }),
  .out1({ S3026 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1513_ (
  .in1({ CU_INC2, S36 }),
  .out1({ S3027 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1514_ (
  .in1({ S3026, S4 }),
  .out1({ S3023 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1515_ (
  .in1({ S3023, S3027 }),
  .out1({ DP_INC_1_inc_value_0 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1516_ (
  .in1({ S5, CU_INC2 }),
  .out1({ S3024 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1517_ (
  .in1({ S37, S3026 }),
  .out1({ S3025 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1518_ (
  .in1({ S3025, S3024 }),
  .out1({ DP_INC_1_inc_value_1 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_39_ (
  .in1({ DP_addrBus_0 }),
  .out1({ addrBus[0] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_40_ (
  .in1({ DP_addrBus_1 }),
  .out1({ addrBus[1] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_41_ (
  .in1({ DP_addrBus_10 }),
  .out1({ addrBus[10] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_42_ (
  .in1({ DP_addrBus_11 }),
  .out1({ addrBus[11] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_43_ (
  .in1({ DP_addrBus_12 }),
  .out1({ addrBus[12] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_44_ (
  .in1({ DP_addrBus_13 }),
  .out1({ addrBus[13] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_45_ (
  .in1({ DP_addrBus_14 }),
  .out1({ addrBus[14] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_46_ (
  .in1({ DP_addrBus_15 }),
  .out1({ addrBus[15] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_47_ (
  .in1({ DP_addrBus_2 }),
  .out1({ addrBus[2] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_48_ (
  .in1({ DP_addrBus_3 }),
  .out1({ addrBus[3] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_49_ (
  .in1({ DP_addrBus_4 }),
  .out1({ addrBus[4] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_50_ (
  .in1({ DP_addrBus_5 }),
  .out1({ addrBus[5] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_51_ (
  .in1({ DP_addrBus_6 }),
  .out1({ addrBus[6] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_52_ (
  .in1({ DP_addrBus_7 }),
  .out1({ addrBus[7] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_53_ (
  .in1({ DP_addrBus_8 }),
  .out1({ addrBus[8] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_54_ (
  .in1({ DP_addrBus_9 }),
  .out1({ addrBus[9] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_55_ (
  .in1({ clk }),
  .out1({ CU_clk })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_56_ (
  .in1({ CU_readMEM }),
  .out1({ readMEM })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_57_ (
  .in1({ rst }),
  .out1({ CU_rst })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_58_ (
  .in1({ CU_seldataBus }),
  .out1({ writeMEM })
);

endmodule