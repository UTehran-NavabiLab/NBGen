module AES(enable, in, key128, expected128, decrypted128, encrypted128, e128, d128);

wire S0;
wire S1;
wire S2;
wire S3;
wire S4;
wire S5;
wire S6;
wire S7;
wire S8;
wire S9;
wire S10;
wire S11;
wire S12;
wire S13;
wire S14;
wire S15;
wire S16;
wire S17;
wire S18;
wire S19;
wire S20;
wire S21;
wire S22;
wire S23;
wire S24;
wire S25;
wire S26;
wire S27;
wire S28;
wire S29;
wire S30;
wire S31;
wire S32;
wire S33;
wire S34;
wire S35;
wire S36;
wire S37;
wire S38;
wire S39;
wire S40;
wire S41;
wire S42;
wire S43;
wire S44;
wire S45;
wire S46;
wire S47;
wire S48;
wire S49;
wire S50;
wire S51;
wire S52;
wire S53;
wire S54;
wire S55;
wire S56;
wire S57;
wire S58;
wire S59;
wire S60;
wire S61;
wire S62;
wire S63;
wire S64;
wire S65;
wire S66;
wire S67;
wire S68;
wire S69;
wire S70;
wire S71;
wire S72;
wire S73;
wire S74;
wire S75;
wire S76;
wire S77;
wire S78;
wire S79;
wire S80;
wire S81;
wire S82;
wire S83;
wire S84;
wire S85;
wire S86;
wire S87;
wire S88;
wire S89;
wire S90;
wire S91;
wire S92;
wire S93;
wire S94;
wire S95;
wire S96;
wire S97;
wire S98;
wire S99;
wire S100;
wire S101;
wire S102;
wire S103;
wire S104;
wire S105;
wire S106;
wire S107;
wire S108;
wire S109;
wire S110;
wire S111;
wire S112;
wire S113;
wire S114;
wire S115;
wire S116;
wire S117;
wire S118;
wire S119;
wire S120;
wire S121;
wire S122;
wire S123;
wire S124;
wire S125;
wire S126;
wire S127;
wire S128;
wire S129;
wire S130;
wire S131;
wire S132;
wire S133;
wire S134;
wire S135;
wire S136;
wire S137;
wire S138;
wire S139;
wire S140;
wire S141;
wire S142;
wire S143;
wire S144;
wire S145;
wire S146;
wire S147;
wire S148;
wire S149;
wire S150;
wire S151;
wire S152;
wire S153;
wire S154;
wire S155;
wire S156;
wire S157;
wire S158;
wire S159;
wire S160;
wire S161;
wire S162;
wire S163;
wire S164;
wire S165;
wire S166;
wire S167;
wire S168;
wire S169;
wire S170;
wire S171;
wire S172;
wire S173;
wire S174;
wire S175;
wire S176;
wire S177;
wire S178;
wire S179;
wire S180;
wire S181;
wire S182;
wire S183;
wire S184;
wire S185;
wire S186;
wire S187;
wire S188;
wire S189;
wire S190;
wire S191;
wire S192;
wire S193;
wire S194;
wire S195;
wire S196;
wire S197;
wire S198;
wire S199;
wire S200;
wire S201;
wire S202;
wire S203;
wire S204;
wire S205;
wire S206;
wire S207;
wire S208;
wire S209;
wire S210;
wire S211;
wire S212;
wire S213;
wire S214;
wire S215;
wire S216;
wire S217;
wire S218;
wire S219;
wire S220;
wire S221;
wire S222;
wire S223;
wire S224;
wire S225;
wire S226;
wire S227;
wire S228;
wire S229;
wire S230;
wire S231;
wire S232;
wire S233;
wire S234;
wire S235;
wire S236;
wire S237;
wire S238;
wire S239;
wire S240;
wire S241;
wire S242;
wire S243;
wire S244;
wire S245;
wire S246;
wire S247;
wire S248;
wire S249;
wire S250;
wire S251;
wire S252;
wire S253;
wire S254;
wire S255;
wire S256;
wire S257;
wire S258;
wire S259;
wire S260;
wire S261;
wire S262;
wire S263;
wire S264;
wire S265;
wire S266;
wire S267;
wire S268;
wire S269;
wire S270;
wire S271;
wire S272;
wire S273;
wire S274;
wire S275;
wire S276;
wire S277;
wire S278;
wire S279;
wire S280;
wire S281;
wire S282;
wire S283;
wire S284;
wire S285;
wire S286;
wire S287;
wire S288;
wire S289;
wire S290;
wire S291;
wire S292;
wire S293;
wire S294;
wire S295;
wire S296;
wire S297;
wire S298;
wire S299;
wire S300;
wire S301;
wire S302;
wire S303;
wire S304;
wire S305;
wire S306;
wire S307;
wire S308;
wire S309;
wire S310;
wire S311;
wire S312;
wire S313;
wire S314;
wire S315;
wire S316;
wire S317;
wire S318;
wire S319;
wire S320;
wire S321;
wire S322;
wire S323;
wire S324;
wire S325;
wire S326;
wire S327;
wire S328;
wire S329;
wire S330;
wire S331;
wire S332;
wire S333;
wire S334;
wire S335;
wire S336;
wire S337;
wire S338;
wire S339;
wire S340;
wire S341;
wire S342;
wire S343;
wire S344;
wire S345;
wire S346;
wire S347;
wire S348;
wire S349;
wire S350;
wire S351;
wire S352;
wire S353;
wire S354;
wire S355;
wire S356;
wire S357;
wire S358;
wire S359;
wire S360;
wire S361;
wire S362;
wire S363;
wire S364;
wire S365;
wire S366;
wire S367;
wire S368;
wire S369;
wire S370;
wire S371;
wire S372;
wire S373;
wire S374;
wire S375;
wire S376;
wire S377;
wire S378;
wire S379;
wire S380;
wire S381;
wire S382;
wire S383;
wire S384;
wire S385;
wire S386;
wire S387;
wire S388;
wire S389;
wire S390;
wire S391;
wire S392;
wire S393;
wire S394;
wire S395;
wire S396;
wire S397;
wire S398;
wire S399;
wire S400;
wire S401;
wire S402;
wire S403;
wire S404;
wire S405;
wire S406;
wire S407;
wire S408;
wire S409;
wire S410;
wire S411;
wire S412;
wire S413;
wire S414;
wire S415;
wire S416;
wire S417;
wire S418;
wire S419;
wire S420;
wire S421;
wire S422;
wire S423;
wire S424;
wire S425;
wire S426;
wire S427;
wire S428;
wire S429;
wire S430;
wire S431;
wire S432;
wire S433;
wire S434;
wire S435;
wire S436;
wire S437;
wire S438;
wire S439;
wire S440;
wire S441;
wire S442;
wire S443;
wire S444;
wire S445;
wire S446;
wire S447;
wire S448;
wire S449;
wire S450;
wire S451;
wire S452;
wire S453;
wire S454;
wire S455;
wire S456;
wire S457;
wire S458;
wire S459;
wire S460;
wire S461;
wire S462;
wire S463;
wire S464;
wire S465;
wire S466;
wire S467;
wire S468;
wire S469;
wire S470;
wire S471;
wire S472;
wire S473;
wire S474;
wire S475;
wire S476;
wire S477;
wire S478;
wire S479;
wire S480;
wire S481;
wire S482;
wire S483;
wire S484;
wire S485;
wire S486;
wire S487;
wire S488;
wire S489;
wire S490;
wire S491;
wire S492;
wire S493;
wire S494;
wire S495;
wire S496;
wire S497;
wire S498;
wire S499;
wire S500;
wire S501;
wire S502;
wire S503;
wire S504;
wire S505;
wire S506;
wire S507;
wire S508;
wire S509;
wire S510;
wire S511;
wire S512;
wire S513;
wire S514;
wire S515;
wire S516;
wire S517;
wire S518;
wire S519;
wire S520;
wire S521;
wire S522;
wire S523;
wire S524;
wire S525;
wire S526;
wire S527;
wire S528;
wire S529;
wire S530;
wire S531;
wire S532;
wire S533;
wire S534;
wire S535;
wire S536;
wire S537;
wire S538;
wire S539;
wire S540;
wire S541;
wire S542;
wire S543;
wire S544;
wire S545;
wire S546;
wire S547;
wire S548;
wire S549;
wire S550;
wire S551;
wire S552;
wire S553;
wire S554;
wire S555;
wire S556;
wire S557;
wire S558;
wire S559;
wire S560;
wire S561;
wire S562;
wire S563;
wire S564;
wire S565;
wire S566;
wire S567;
wire S568;
wire S569;
wire S570;
wire S571;
wire S572;
wire S573;
wire S574;
wire S575;
wire S576;
wire S577;
wire S578;
wire S579;
wire S580;
wire S581;
wire S582;
wire S583;
wire S584;
wire S585;
wire S586;
wire S587;
wire S588;
wire S589;
wire S590;
wire S591;
wire S592;
wire S593;
wire S594;
wire S595;
wire S596;
wire S597;
wire S598;
wire S599;
wire S600;
wire S601;
wire S602;
wire S603;
wire S604;
wire S605;
wire S606;
wire S607;
wire S608;
wire S609;
wire S610;
wire S611;
wire S612;
wire S613;
wire S614;
wire S615;
wire S616;
wire S617;
wire S618;
wire S619;
wire S620;
wire S621;
wire S622;
wire S623;
wire S624;
wire S625;
wire S626;
wire S627;
wire S628;
wire S629;
wire S630;
wire S631;
wire S632;
wire S633;
wire S634;
wire S635;
wire S636;
wire S637;
wire S638;
wire S639;
wire S640;
wire S641;
wire S642;
wire S643;
wire S644;
wire S645;
wire S646;
wire S647;
wire S648;
wire S649;
wire S650;
wire S651;
wire S652;
wire S653;
wire S654;
wire S655;
wire S656;
wire S657;
wire S658;
wire S659;
wire S660;
wire S661;
wire S662;
wire S663;
wire S664;
wire S665;
wire S666;
wire S667;
wire S668;
wire S669;
wire S670;
wire S671;
wire S672;
wire S673;
wire S674;
wire S675;
wire S676;
wire S677;
wire S678;
wire S679;
wire S680;
wire S681;
wire S682;
wire S683;
wire S684;
wire S685;
wire S686;
wire S687;
wire S688;
wire S689;
wire S690;
wire S691;
wire S692;
wire S693;
wire S694;
wire S695;
wire S696;
wire S697;
wire S698;
wire S699;
wire S700;
wire S701;
wire S702;
wire S703;
wire S704;
wire S705;
wire S706;
wire S707;
wire S708;
wire S709;
wire S710;
wire S711;
wire S712;
wire S713;
wire S714;
wire S715;
wire S716;
wire S717;
wire S718;
wire S719;
wire S720;
wire S721;
wire S722;
wire S723;
wire S724;
wire S725;
wire S726;
wire S727;
wire S728;
wire S729;
wire S730;
wire S731;
wire S732;
wire S733;
wire S734;
wire S735;
wire S736;
wire S737;
wire S738;
wire S739;
wire S740;
wire S741;
wire S742;
wire S743;
wire S744;
wire S745;
wire S746;
wire S747;
wire S748;
wire S749;
wire S750;
wire S751;
wire S752;
wire S753;
wire S754;
wire S755;
wire S756;
wire S757;
wire S758;
wire S759;
wire S760;
wire S761;
wire S762;
wire S763;
wire S764;
wire S765;
wire S766;
wire S767;
wire S768;
wire S769;
wire S770;
wire S771;
wire S772;
wire S773;
wire S774;
wire S775;
wire S776;
wire S777;
wire S778;
wire S779;
wire S780;
wire S781;
wire S782;
wire S783;
wire S784;
wire S785;
wire S786;
wire S787;
wire S788;
wire S789;
wire S790;
wire S791;
wire S792;
wire S793;
input enable;
input [127:0] in;input [127:0] key128;input [127:0] expected128;output [127:0] decrypted128;output [127:0] encrypted128;output e128;
output d128;

XNOR2_X1 #() 
XNOR2_X1_1_ (
  .A({ S791[72] }),
  .B({ S790[72] }),
  .ZN({ S303 })
);
XNOR2_X1 #() 
XNOR2_X1_2_ (
  .A({ S791[98] }),
  .B({ S790[98] }),
  .ZN({ S304 })
);
XNOR2_X1 #() 
XNOR2_X1_3_ (
  .A({ S791[100] }),
  .B({ S790[100] }),
  .ZN({ S305 })
);
NAND3_X1 #() 
NAND3_X1_1_ (
  .A1({ S303 }),
  .A2({ S304 }),
  .A3({ S305 }),
  .ZN({ S306 })
);
XNOR2_X1 #() 
XNOR2_X1_4_ (
  .A({ S791[96] }),
  .B({ S790[96] }),
  .ZN({ S307 })
);
INV_X1 #() 
INV_X1_1_ (
  .A({ S790[34] }),
  .ZN({ S308 })
);
INV_X1 #() 
INV_X1_2_ (
  .A({ S789 }),
  .ZN({ S309 })
);
AOI21_X1 #() 
AOI21_X1_1_ (
  .A({ S309 }),
  .B1({ S308 }),
  .B2({ S791[34] }),
  .ZN({ S310 })
);
XNOR2_X1 #() 
XNOR2_X1_5_ (
  .A({ S791[26] }),
  .B({ S790[26] }),
  .ZN({ S311 })
);
XNOR2_X1 #() 
XNOR2_X1_6_ (
  .A({ S791[28] }),
  .B({ S790[28] }),
  .ZN({ S312 })
);
NAND4_X1 #() 
NAND4_X1_1_ (
  .A1({ S311 }),
  .A2({ S312 }),
  .A3({ S307 }),
  .A4({ S310 }),
  .ZN({ S313 })
);
INV_X1 #() 
INV_X1_3_ (
  .A({ S791[56] }),
  .ZN({ S314 })
);
INV_X1 #() 
INV_X1_4_ (
  .A({ S790[66] }),
  .ZN({ S315 })
);
AOI22_X1 #() 
AOI22_X1_1_ (
  .A1({ S314 }),
  .A2({ S790[56] }),
  .B1({ S315 }),
  .B2({ S791[66] }),
  .ZN({ S316 })
);
XNOR2_X1 #() 
XNOR2_X1_7_ (
  .A({ S791[36] }),
  .B({ S790[36] }),
  .ZN({ S317 })
);
INV_X1 #() 
INV_X1_5_ (
  .A({ S791[34] }),
  .ZN({ S318 })
);
INV_X1 #() 
INV_X1_6_ (
  .A({ S790[54] }),
  .ZN({ S319 })
);
AOI22_X1 #() 
AOI22_X1_2_ (
  .A1({ S318 }),
  .A2({ S790[34] }),
  .B1({ S319 }),
  .B2({ S791[54] }),
  .ZN({ S320 })
);
INV_X1 #() 
INV_X1_7_ (
  .A({ S791[54] }),
  .ZN({ S321 })
);
INV_X1 #() 
INV_X1_8_ (
  .A({ S790[56] }),
  .ZN({ S322 })
);
AOI22_X1 #() 
AOI22_X1_3_ (
  .A1({ S321 }),
  .A2({ S790[54] }),
  .B1({ S322 }),
  .B2({ S791[56] }),
  .ZN({ S323 })
);
NAND4_X1 #() 
NAND4_X1_2_ (
  .A1({ S323 }),
  .A2({ S320 }),
  .A3({ S317 }),
  .A4({ S316 }),
  .ZN({ S324 })
);
NOR3_X1 #() 
NOR3_X1_1_ (
  .A1({ S324 }),
  .A2({ S313 }),
  .A3({ S306 }),
  .ZN({ S325 })
);
INV_X1 #() 
INV_X1_9_ (
  .A({ S790[60] }),
  .ZN({ S326 })
);
INV_X1 #() 
INV_X1_10_ (
  .A({ S791[64] }),
  .ZN({ S327 })
);
AOI22_X1 #() 
AOI22_X1_4_ (
  .A1({ S327 }),
  .A2({ S790[64] }),
  .B1({ S326 }),
  .B2({ S791[60] }),
  .ZN({ S328 })
);
INV_X1 #() 
INV_X1_11_ (
  .A({ S790[58] }),
  .ZN({ S329 })
);
INV_X1 #() 
INV_X1_12_ (
  .A({ S791[60] }),
  .ZN({ S330 })
);
AOI22_X1 #() 
AOI22_X1_5_ (
  .A1({ S330 }),
  .A2({ S790[60] }),
  .B1({ S329 }),
  .B2({ S791[58] }),
  .ZN({ S331 })
);
INV_X1 #() 
INV_X1_13_ (
  .A({ S790[74] }),
  .ZN({ S332 })
);
INV_X1 #() 
INV_X1_14_ (
  .A({ S791[76] }),
  .ZN({ S333 })
);
AOI22_X1 #() 
AOI22_X1_6_ (
  .A1({ S333 }),
  .A2({ S790[76] }),
  .B1({ S332 }),
  .B2({ S791[74] }),
  .ZN({ S334 })
);
INV_X1 #() 
INV_X1_15_ (
  .A({ S790[64] }),
  .ZN({ S335 })
);
INV_X1 #() 
INV_X1_16_ (
  .A({ S791[74] }),
  .ZN({ S336 })
);
AOI22_X1 #() 
AOI22_X1_7_ (
  .A1({ S336 }),
  .A2({ S790[74] }),
  .B1({ S335 }),
  .B2({ S791[64] }),
  .ZN({ S337 })
);
AND4_X1 #() 
AND4_X1_1_ (
  .A1({ S328 }),
  .A2({ S334 }),
  .A3({ S337 }),
  .A4({ S331 }),
  .ZN({ S338 })
);
INV_X1 #() 
INV_X1_17_ (
  .A({ S791[82] }),
  .ZN({ S339 })
);
NAND2_X1 #() 
NAND2_X1_1_ (
  .A1({ S339 }),
  .A2({ S790[82] }),
  .ZN({ S340 })
);
INV_X1 #() 
INV_X1_18_ (
  .A({ S790[8] }),
  .ZN({ S341 })
);
NAND2_X1 #() 
NAND2_X1_2_ (
  .A1({ S341 }),
  .A2({ S791[8] }),
  .ZN({ S342 })
);
INV_X1 #() 
INV_X1_19_ (
  .A({ S791[8] }),
  .ZN({ S343 })
);
NAND2_X1 #() 
NAND2_X1_3_ (
  .A1({ S343 }),
  .A2({ S790[8] }),
  .ZN({ S344 })
);
INV_X1 #() 
INV_X1_20_ (
  .A({ S790[12] }),
  .ZN({ S345 })
);
NAND2_X1 #() 
NAND2_X1_4_ (
  .A1({ S345 }),
  .A2({ S791[12] }),
  .ZN({ S346 })
);
NAND4_X1 #() 
NAND4_X1_3_ (
  .A1({ S344 }),
  .A2({ S346 }),
  .A3({ S340 }),
  .A4({ S342 }),
  .ZN({ S347 })
);
INV_X1 #() 
INV_X1_21_ (
  .A({ S791[58] }),
  .ZN({ S348 })
);
NAND2_X1 #() 
NAND2_X1_5_ (
  .A1({ S348 }),
  .A2({ S790[58] }),
  .ZN({ S349 })
);
INV_X1 #() 
INV_X1_22_ (
  .A({ S790[62] }),
  .ZN({ S350 })
);
NAND2_X1 #() 
NAND2_X1_6_ (
  .A1({ S350 }),
  .A2({ S791[62] }),
  .ZN({ S351 })
);
INV_X1 #() 
INV_X1_23_ (
  .A({ S791[62] }),
  .ZN({ S352 })
);
NAND2_X1 #() 
NAND2_X1_7_ (
  .A1({ S352 }),
  .A2({ S790[62] }),
  .ZN({ S353 })
);
INV_X1 #() 
INV_X1_24_ (
  .A({ S790[82] }),
  .ZN({ S354 })
);
NAND2_X1 #() 
NAND2_X1_8_ (
  .A1({ S354 }),
  .A2({ S791[82] }),
  .ZN({ S355 })
);
NAND4_X1 #() 
NAND4_X1_4_ (
  .A1({ S353 }),
  .A2({ S355 }),
  .A3({ S349 }),
  .A4({ S351 }),
  .ZN({ S356 })
);
NOR2_X1 #() 
NOR2_X1_1_ (
  .A1({ S347 }),
  .A2({ S356 }),
  .ZN({ S357 })
);
INV_X1 #() 
INV_X1_25_ (
  .A({ S791[32] }),
  .ZN({ S358 })
);
NAND2_X1 #() 
NAND2_X1_9_ (
  .A1({ S358 }),
  .A2({ S790[32] }),
  .ZN({ S359 })
);
INV_X1 #() 
INV_X1_26_ (
  .A({ S790[22] }),
  .ZN({ S360 })
);
NAND2_X1 #() 
NAND2_X1_10_ (
  .A1({ S360 }),
  .A2({ S791[22] }),
  .ZN({ S361 })
);
INV_X1 #() 
INV_X1_27_ (
  .A({ S791[22] }),
  .ZN({ S362 })
);
NAND2_X1 #() 
NAND2_X1_11_ (
  .A1({ S362 }),
  .A2({ S790[22] }),
  .ZN({ S363 })
);
INV_X1 #() 
INV_X1_28_ (
  .A({ S790[80] }),
  .ZN({ S364 })
);
NAND2_X1 #() 
NAND2_X1_12_ (
  .A1({ S364 }),
  .A2({ S791[80] }),
  .ZN({ S365 })
);
NAND4_X1 #() 
NAND4_X1_5_ (
  .A1({ S363 }),
  .A2({ S365 }),
  .A3({ S359 }),
  .A4({ S361 }),
  .ZN({ S366 })
);
INV_X1 #() 
INV_X1_29_ (
  .A({ S790[32] }),
  .ZN({ S367 })
);
NAND2_X1 #() 
NAND2_X1_13_ (
  .A1({ S367 }),
  .A2({ S791[32] }),
  .ZN({ S368 })
);
INV_X1 #() 
INV_X1_30_ (
  .A({ S791[66] }),
  .ZN({ S369 })
);
NAND2_X1 #() 
NAND2_X1_14_ (
  .A1({ S369 }),
  .A2({ S790[66] }),
  .ZN({ S370 })
);
AND2_X1 #() 
AND2_X1_1_ (
  .A1({ S790[68] }),
  .A2({ S791[68] }),
  .ZN({ S371 })
);
NOR2_X1 #() 
NOR2_X1_2_ (
  .A1({ S791[68] }),
  .A2({ S790[68] }),
  .ZN({ S372 })
);
OAI211_X1 #() 
OAI211_X1_1_ (
  .A({ S370 }),
  .B({ S368 }),
  .C1({ S371 }),
  .C2({ S372 }),
  .ZN({ S373 })
);
NOR2_X1 #() 
NOR2_X1_3_ (
  .A1({ S366 }),
  .A2({ S373 }),
  .ZN({ S374 })
);
INV_X1 #() 
INV_X1_31_ (
  .A({ S791[70] }),
  .ZN({ S375 })
);
NAND2_X1 #() 
NAND2_X1_15_ (
  .A1({ S375 }),
  .A2({ S790[70] }),
  .ZN({ S376 })
);
INV_X1 #() 
INV_X1_32_ (
  .A({ S790[84] }),
  .ZN({ S377 })
);
NAND2_X1 #() 
NAND2_X1_16_ (
  .A1({ S377 }),
  .A2({ S791[84] }),
  .ZN({ S378 })
);
INV_X1 #() 
INV_X1_33_ (
  .A({ S791[84] }),
  .ZN({ S379 })
);
NAND2_X1 #() 
NAND2_X1_17_ (
  .A1({ S379 }),
  .A2({ S790[84] }),
  .ZN({ S380 })
);
INV_X1 #() 
INV_X1_34_ (
  .A({ S790[76] }),
  .ZN({ S381 })
);
NAND2_X1 #() 
NAND2_X1_18_ (
  .A1({ S381 }),
  .A2({ S791[76] }),
  .ZN({ S382 })
);
NAND4_X1 #() 
NAND4_X1_6_ (
  .A1({ S380 }),
  .A2({ S382 }),
  .A3({ S376 }),
  .A4({ S378 }),
  .ZN({ S383 })
);
INV_X1 #() 
INV_X1_35_ (
  .A({ S791[80] }),
  .ZN({ S384 })
);
NAND2_X1 #() 
NAND2_X1_19_ (
  .A1({ S384 }),
  .A2({ S790[80] }),
  .ZN({ S385 })
);
INV_X1 #() 
INV_X1_36_ (
  .A({ S790[78] }),
  .ZN({ S386 })
);
NAND2_X1 #() 
NAND2_X1_20_ (
  .A1({ S386 }),
  .A2({ S791[78] }),
  .ZN({ S387 })
);
INV_X1 #() 
INV_X1_37_ (
  .A({ S791[78] }),
  .ZN({ S388 })
);
NAND2_X1 #() 
NAND2_X1_21_ (
  .A1({ S388 }),
  .A2({ S790[78] }),
  .ZN({ S389 })
);
INV_X1 #() 
INV_X1_38_ (
  .A({ S790[70] }),
  .ZN({ S390 })
);
NAND2_X1 #() 
NAND2_X1_22_ (
  .A1({ S390 }),
  .A2({ S791[70] }),
  .ZN({ S391 })
);
NAND4_X1 #() 
NAND4_X1_7_ (
  .A1({ S389 }),
  .A2({ S391 }),
  .A3({ S385 }),
  .A4({ S387 }),
  .ZN({ S392 })
);
NOR2_X1 #() 
NOR2_X1_4_ (
  .A1({ S383 }),
  .A2({ S392 }),
  .ZN({ S393 })
);
AND4_X1 #() 
AND4_X1_2_ (
  .A1({ S338 }),
  .A2({ S393 }),
  .A3({ S357 }),
  .A4({ S374 }),
  .ZN({ S394 })
);
INV_X1 #() 
INV_X1_39_ (
  .A({ S790[59] }),
  .ZN({ S395 })
);
INV_X1 #() 
INV_X1_40_ (
  .A({ S791[75] }),
  .ZN({ S396 })
);
OAI22_X1 #() 
OAI22_X1_1_ (
  .A1({ S395 }),
  .A2({ S791[59] }),
  .B1({ S396 }),
  .B2({ S790[75] }),
  .ZN({ S397 })
);
INV_X1 #() 
INV_X1_41_ (
  .A({ S791[63] }),
  .ZN({ S398 })
);
AND2_X1 #() 
AND2_X1_2_ (
  .A1({ S398 }),
  .A2({ S790[63] }),
  .ZN({ S399 })
);
NOR2_X1 #() 
NOR2_X1_5_ (
  .A1({ S398 }),
  .A2({ S790[63] }),
  .ZN({ S400 })
);
NOR3_X1 #() 
NOR3_X1_2_ (
  .A1({ S397 }),
  .A2({ S399 }),
  .A3({ S400 }),
  .ZN({ S401 })
);
INV_X1 #() 
INV_X1_42_ (
  .A({ S791[73] }),
  .ZN({ S402 })
);
INV_X1 #() 
INV_X1_43_ (
  .A({ S790[83] }),
  .ZN({ S403 })
);
AOI22_X1 #() 
AOI22_X1_8_ (
  .A1({ S402 }),
  .A2({ S790[73] }),
  .B1({ S403 }),
  .B2({ S791[83] }),
  .ZN({ S404 })
);
INV_X1 #() 
INV_X1_44_ (
  .A({ S791[69] }),
  .ZN({ S405 })
);
AOI22_X1 #() 
AOI22_X1_9_ (
  .A1({ S790[69] }),
  .A2({ S405 }),
  .B1({ S396 }),
  .B2({ S790[75] }),
  .ZN({ S406 })
);
AND2_X1 #() 
AND2_X1_3_ (
  .A1({ S406 }),
  .A2({ S404 }),
  .ZN({ S407 })
);
INV_X1 #() 
INV_X1_45_ (
  .A({ S790[57] }),
  .ZN({ S408 })
);
INV_X1 #() 
INV_X1_46_ (
  .A({ S791[65] }),
  .ZN({ S409 })
);
OAI22_X1 #() 
OAI22_X1_2_ (
  .A1({ S408 }),
  .A2({ S791[57] }),
  .B1({ S409 }),
  .B2({ S790[65] }),
  .ZN({ S410 })
);
INV_X1 #() 
INV_X1_47_ (
  .A({ S791[61] }),
  .ZN({ S411 })
);
OAI22_X1 #() 
OAI22_X1_3_ (
  .A1({ S411 }),
  .A2({ S790[61] }),
  .B1({ S403 }),
  .B2({ S791[83] }),
  .ZN({ S412 })
);
NOR2_X1 #() 
NOR2_X1_6_ (
  .A1({ S410 }),
  .A2({ S412 }),
  .ZN({ S413 })
);
INV_X1 #() 
INV_X1_48_ (
  .A({ S790[71] }),
  .ZN({ S414 })
);
INV_X1 #() 
INV_X1_49_ (
  .A({ S790[77] }),
  .ZN({ S415 })
);
AOI22_X1 #() 
AOI22_X1_10_ (
  .A1({ S791[77] }),
  .A2({ S415 }),
  .B1({ S414 }),
  .B2({ S791[71] }),
  .ZN({ S416 })
);
INV_X1 #() 
INV_X1_50_ (
  .A({ S791[31] }),
  .ZN({ S417 })
);
AOI22_X1 #() 
AOI22_X1_11_ (
  .A1({ S790[31] }),
  .A2({ S417 }),
  .B1({ S411 }),
  .B2({ S790[61] }),
  .ZN({ S418 })
);
AND2_X1 #() 
AND2_X1_4_ (
  .A1({ S418 }),
  .A2({ S416 }),
  .ZN({ S419 })
);
NAND4_X1 #() 
NAND4_X1_8_ (
  .A1({ S419 }),
  .A2({ S407 }),
  .A3({ S401 }),
  .A4({ S413 }),
  .ZN({ S420 })
);
INV_X1 #() 
INV_X1_51_ (
  .A({ S791[42] }),
  .ZN({ S421 })
);
INV_X1 #() 
INV_X1_52_ (
  .A({ S790[46] }),
  .ZN({ S422 })
);
OAI22_X1 #() 
OAI22_X1_4_ (
  .A1({ S421 }),
  .A2({ S790[42] }),
  .B1({ S422 }),
  .B2({ S791[46] }),
  .ZN({ S423 })
);
INV_X1 #() 
INV_X1_53_ (
  .A({ S791[40] }),
  .ZN({ S424 })
);
INV_X1 #() 
INV_X1_54_ (
  .A({ S790[42] }),
  .ZN({ S425 })
);
OAI22_X1 #() 
OAI22_X1_5_ (
  .A1({ S424 }),
  .A2({ S790[40] }),
  .B1({ S425 }),
  .B2({ S791[42] }),
  .ZN({ S426 })
);
NOR2_X1 #() 
NOR2_X1_7_ (
  .A1({ S423 }),
  .A2({ S426 }),
  .ZN({ S427 })
);
INV_X1 #() 
INV_X1_55_ (
  .A({ S791[10] }),
  .ZN({ S428 })
);
OAI22_X1 #() 
OAI22_X1_6_ (
  .A1({ S428 }),
  .A2({ S790[10] }),
  .B1({ S345 }),
  .B2({ S791[12] }),
  .ZN({ S429 })
);
INV_X1 #() 
INV_X1_56_ (
  .A({ S790[10] }),
  .ZN({ S430 })
);
INV_X1 #() 
INV_X1_57_ (
  .A({ S791[46] }),
  .ZN({ S431 })
);
OAI22_X1 #() 
OAI22_X1_7_ (
  .A1({ S430 }),
  .A2({ S791[10] }),
  .B1({ S431 }),
  .B2({ S790[46] }),
  .ZN({ S432 })
);
NOR2_X1 #() 
NOR2_X1_8_ (
  .A1({ S429 }),
  .A2({ S432 }),
  .ZN({ S433 })
);
INV_X1 #() 
INV_X1_58_ (
  .A({ S791[6] }),
  .ZN({ S434 })
);
AOI22_X1 #() 
AOI22_X1_12_ (
  .A1({ S434 }),
  .A2({ S790[6] }),
  .B1({ S395 }),
  .B2({ S791[59] }),
  .ZN({ S435 })
);
INV_X1 #() 
INV_X1_59_ (
  .A({ S790[41] }),
  .ZN({ S436 })
);
INV_X1 #() 
INV_X1_60_ (
  .A({ S791[81] }),
  .ZN({ S437 })
);
AOI22_X1 #() 
AOI22_X1_13_ (
  .A1({ S437 }),
  .A2({ S790[81] }),
  .B1({ S436 }),
  .B2({ S791[41] }),
  .ZN({ S438 })
);
AND2_X1 #() 
AND2_X1_5_ (
  .A1({ S438 }),
  .A2({ S435 }),
  .ZN({ S439 })
);
INV_X1 #() 
INV_X1_61_ (
  .A({ S790[40] }),
  .ZN({ S440 })
);
INV_X1 #() 
INV_X1_62_ (
  .A({ S791[44] }),
  .ZN({ S441 })
);
OAI22_X1 #() 
OAI22_X1_8_ (
  .A1({ S440 }),
  .A2({ S791[40] }),
  .B1({ S441 }),
  .B2({ S790[44] }),
  .ZN({ S442 })
);
INV_X1 #() 
INV_X1_63_ (
  .A({ S790[44] }),
  .ZN({ S443 })
);
OAI22_X1 #() 
OAI22_X1_9_ (
  .A1({ S434 }),
  .A2({ S790[6] }),
  .B1({ S443 }),
  .B2({ S791[44] }),
  .ZN({ S444 })
);
NOR2_X1 #() 
NOR2_X1_9_ (
  .A1({ S442 }),
  .A2({ S444 }),
  .ZN({ S445 })
);
NAND4_X1 #() 
NAND4_X1_9_ (
  .A1({ S439 }),
  .A2({ S445 }),
  .A3({ S427 }),
  .A4({ S433 }),
  .ZN({ S446 })
);
NOR2_X1 #() 
NOR2_X1_10_ (
  .A1({ S420 }),
  .A2({ S446 }),
  .ZN({ S447 })
);
NAND3_X1 #() 
NAND3_X1_2_ (
  .A1({ S447 }),
  .A2({ S394 }),
  .A3({ S325 }),
  .ZN({ S448 })
);
INV_X1 #() 
INV_X1_64_ (
  .A({ S790[127] }),
  .ZN({ S449 })
);
INV_X1 #() 
INV_X1_65_ (
  .A({ S791[125] }),
  .ZN({ S450 })
);
AOI22_X1 #() 
AOI22_X1_14_ (
  .A1({ S450 }),
  .A2({ S790[125] }),
  .B1({ S449 }),
  .B2({ S791[127] }),
  .ZN({ S451 })
);
OAI21_X1 #() 
OAI21_X1_1_ (
  .A({ S451 }),
  .B1({ S791[127] }),
  .B2({ S449 }),
  .ZN({ S452 })
);
INV_X1 #() 
INV_X1_66_ (
  .A({ S791[122] }),
  .ZN({ S453 })
);
INV_X1 #() 
INV_X1_67_ (
  .A({ S791[126] }),
  .ZN({ S454 })
);
NAND2_X1 #() 
NAND2_X1_23_ (
  .A1({ S454 }),
  .A2({ S790[126] }),
  .ZN({ S455 })
);
INV_X1 #() 
INV_X1_68_ (
  .A({ S791[123] }),
  .ZN({ S456 })
);
AOI22_X1 #() 
AOI22_X1_15_ (
  .A1({ S790[122] }),
  .A2({ S453 }),
  .B1({ S456 }),
  .B2({ S790[123] }),
  .ZN({ S457 })
);
OAI211_X1 #() 
OAI211_X1_2_ (
  .A({ S457 }),
  .B({ S455 }),
  .C1({ S790[122] }),
  .C2({ S453 }),
  .ZN({ S458 })
);
INV_X1 #() 
INV_X1_69_ (
  .A({ S791[117] }),
  .ZN({ S459 })
);
INV_X1 #() 
INV_X1_70_ (
  .A({ S790[109] }),
  .ZN({ S460 })
);
AOI22_X1 #() 
AOI22_X1_16_ (
  .A1({ S459 }),
  .A2({ S790[117] }),
  .B1({ S460 }),
  .B2({ S791[109] }),
  .ZN({ S461 })
);
OAI221_X1 #() 
OAI221_X1_1_ (
  .A({ S461 }),
  .B1({ S454 }),
  .B2({ S790[126] }),
  .C1({ S790[117] }),
  .C2({ S459 }),
  .ZN({ S462 })
);
NOR3_X1 #() 
NOR3_X1_3_ (
  .A1({ S462 }),
  .A2({ S458 }),
  .A3({ S452 }),
  .ZN({ S463 })
);
INV_X1 #() 
INV_X1_71_ (
  .A({ S791[16] }),
  .ZN({ S464 })
);
INV_X1 #() 
INV_X1_72_ (
  .A({ S790[18] }),
  .ZN({ S465 })
);
OAI22_X1 #() 
OAI22_X1_10_ (
  .A1({ S464 }),
  .A2({ S790[16] }),
  .B1({ S465 }),
  .B2({ S791[18] }),
  .ZN({ S466 })
);
INV_X1 #() 
INV_X1_73_ (
  .A({ S791[14] }),
  .ZN({ S467 })
);
INV_X1 #() 
INV_X1_74_ (
  .A({ S790[16] }),
  .ZN({ S468 })
);
OAI22_X1 #() 
OAI22_X1_11_ (
  .A1({ S467 }),
  .A2({ S790[14] }),
  .B1({ S468 }),
  .B2({ S791[16] }),
  .ZN({ S469 })
);
INV_X1 #() 
INV_X1_75_ (
  .A({ S790[106] }),
  .ZN({ S470 })
);
INV_X1 #() 
INV_X1_76_ (
  .A({ S791[124] }),
  .ZN({ S471 })
);
AOI22_X1 #() 
AOI22_X1_17_ (
  .A1({ S471 }),
  .A2({ S790[124] }),
  .B1({ S470 }),
  .B2({ S791[106] }),
  .ZN({ S472 })
);
INV_X1 #() 
INV_X1_77_ (
  .A({ S791[106] }),
  .ZN({ S473 })
);
AOI22_X1 #() 
AOI22_X1_18_ (
  .A1({ S473 }),
  .A2({ S790[106] }),
  .B1({ S465 }),
  .B2({ S791[18] }),
  .ZN({ S474 })
);
NAND2_X1 #() 
NAND2_X1_24_ (
  .A1({ S472 }),
  .A2({ S474 }),
  .ZN({ S475 })
);
INV_X1 #() 
INV_X1_78_ (
  .A({ S791[115] }),
  .ZN({ S476 })
);
INV_X1 #() 
INV_X1_79_ (
  .A({ S790[121] }),
  .ZN({ S477 })
);
AOI22_X1 #() 
AOI22_X1_19_ (
  .A1({ S476 }),
  .A2({ S790[115] }),
  .B1({ S477 }),
  .B2({ S791[121] }),
  .ZN({ S478 })
);
INV_X1 #() 
INV_X1_80_ (
  .A({ S791[105] }),
  .ZN({ S479 })
);
INV_X1 #() 
INV_X1_81_ (
  .A({ S791[113] }),
  .ZN({ S480 })
);
AOI22_X1 #() 
AOI22_X1_20_ (
  .A1({ S790[105] }),
  .A2({ S479 }),
  .B1({ S480 }),
  .B2({ S790[113] }),
  .ZN({ S481 })
);
INV_X1 #() 
INV_X1_82_ (
  .A({ S790[4] }),
  .ZN({ S482 })
);
AOI22_X1 #() 
AOI22_X1_21_ (
  .A1({ S467 }),
  .A2({ S790[14] }),
  .B1({ S482 }),
  .B2({ S791[4] }),
  .ZN({ S483 })
);
INV_X1 #() 
INV_X1_83_ (
  .A({ S791[4] }),
  .ZN({ S484 })
);
INV_X1 #() 
INV_X1_84_ (
  .A({ S790[115] }),
  .ZN({ S485 })
);
AOI22_X1 #() 
AOI22_X1_22_ (
  .A1({ S484 }),
  .A2({ S790[4] }),
  .B1({ S485 }),
  .B2({ S791[115] }),
  .ZN({ S486 })
);
NAND4_X1 #() 
NAND4_X1_10_ (
  .A1({ S483 }),
  .A2({ S486 }),
  .A3({ S478 }),
  .A4({ S481 }),
  .ZN({ S487 })
);
NOR4_X1 #() 
NOR4_X1_1_ (
  .A1({ S487 }),
  .A2({ S475 }),
  .A3({ S469 }),
  .A4({ S466 }),
  .ZN({ S488 })
);
INV_X1 #() 
INV_X1_85_ (
  .A({ S790[37] }),
  .ZN({ S489 })
);
INV_X1 #() 
INV_X1_86_ (
  .A({ S791[77] }),
  .ZN({ S490 })
);
AOI22_X1 #() 
AOI22_X1_23_ (
  .A1({ S490 }),
  .A2({ S790[77] }),
  .B1({ S489 }),
  .B2({ S791[37] }),
  .ZN({ S491 })
);
INV_X1 #() 
INV_X1_87_ (
  .A({ S791[53] }),
  .ZN({ S492 })
);
INV_X1 #() 
INV_X1_88_ (
  .A({ S790[81] }),
  .ZN({ S493 })
);
AOI22_X1 #() 
AOI22_X1_24_ (
  .A1({ S492 }),
  .A2({ S790[53] }),
  .B1({ S493 }),
  .B2({ S791[81] }),
  .ZN({ S494 })
);
INV_X1 #() 
INV_X1_89_ (
  .A({ S791[91] }),
  .ZN({ S495 })
);
INV_X1 #() 
INV_X1_90_ (
  .A({ S790[93] }),
  .ZN({ S496 })
);
AOI22_X1 #() 
AOI22_X1_25_ (
  .A1({ S495 }),
  .A2({ S790[91] }),
  .B1({ S496 }),
  .B2({ S791[93] }),
  .ZN({ S497 })
);
INV_X1 #() 
INV_X1_91_ (
  .A({ S791[33] }),
  .ZN({ S498 })
);
INV_X1 #() 
INV_X1_92_ (
  .A({ S791[87] }),
  .ZN({ S499 })
);
AOI22_X1 #() 
AOI22_X1_26_ (
  .A1({ S790[33] }),
  .A2({ S498 }),
  .B1({ S499 }),
  .B2({ S790[87] }),
  .ZN({ S500 })
);
NAND4_X1 #() 
NAND4_X1_11_ (
  .A1({ S497 }),
  .A2({ S500 }),
  .A3({ S491 }),
  .A4({ S494 }),
  .ZN({ S501 })
);
INV_X1 #() 
INV_X1_93_ (
  .A({ S791[110] }),
  .ZN({ S502 })
);
INV_X1 #() 
INV_X1_94_ (
  .A({ S790[116] }),
  .ZN({ S503 })
);
OAI22_X1 #() 
OAI22_X1_12_ (
  .A1({ S502 }),
  .A2({ S790[110] }),
  .B1({ S503 }),
  .B2({ S791[116] }),
  .ZN({ S504 })
);
INV_X1 #() 
INV_X1_95_ (
  .A({ S790[110] }),
  .ZN({ S505 })
);
OAI22_X1 #() 
OAI22_X1_13_ (
  .A1({ S505 }),
  .A2({ S791[110] }),
  .B1({ S471 }),
  .B2({ S790[124] }),
  .ZN({ S506 })
);
INV_X1 #() 
INV_X1_96_ (
  .A({ S791[55] }),
  .ZN({ S507 })
);
AOI22_X1 #() 
AOI22_X1_27_ (
  .A1({ S507 }),
  .A2({ S790[55] }),
  .B1({ S408 }),
  .B2({ S791[57] }),
  .ZN({ S508 })
);
INV_X1 #() 
INV_X1_97_ (
  .A({ S790[67] }),
  .ZN({ S509 })
);
AOI22_X1 #() 
AOI22_X1_28_ (
  .A1({ S791[116] }),
  .A2({ S503 }),
  .B1({ S509 }),
  .B2({ S791[67] }),
  .ZN({ S510 })
);
NAND2_X1 #() 
NAND2_X1_25_ (
  .A1({ S508 }),
  .A2({ S510 }),
  .ZN({ S511 })
);
NOR4_X1 #() 
NOR4_X1_2_ (
  .A1({ S501 }),
  .A2({ S511 }),
  .A3({ S506 }),
  .A4({ S504 }),
  .ZN({ S512 })
);
NAND3_X1 #() 
NAND3_X1_3_ (
  .A1({ S488 }),
  .A2({ S512 }),
  .A3({ S463 }),
  .ZN({ S513 })
);
INV_X1 #() 
INV_X1_98_ (
  .A({ S790[94] }),
  .ZN({ S514 })
);
NAND2_X1 #() 
NAND2_X1_26_ (
  .A1({ S514 }),
  .A2({ S791[94] }),
  .ZN({ S515 })
);
INV_X1 #() 
INV_X1_99_ (
  .A({ S791[24] }),
  .ZN({ S516 })
);
NAND2_X1 #() 
NAND2_X1_27_ (
  .A1({ S516 }),
  .A2({ S790[24] }),
  .ZN({ S517 })
);
INV_X1 #() 
INV_X1_100_ (
  .A({ S790[24] }),
  .ZN({ S518 })
);
NAND2_X1 #() 
NAND2_X1_28_ (
  .A1({ S518 }),
  .A2({ S791[24] }),
  .ZN({ S519 })
);
INV_X1 #() 
INV_X1_101_ (
  .A({ S790[33] }),
  .ZN({ S520 })
);
NAND2_X1 #() 
NAND2_X1_29_ (
  .A1({ S520 }),
  .A2({ S791[33] }),
  .ZN({ S521 })
);
NAND4_X1 #() 
NAND4_X1_12_ (
  .A1({ S519 }),
  .A2({ S521 }),
  .A3({ S515 }),
  .A4({ S517 }),
  .ZN({ S522 })
);
INV_X1 #() 
INV_X1_102_ (
  .A({ S791[90] }),
  .ZN({ S523 })
);
NAND2_X1 #() 
NAND2_X1_30_ (
  .A1({ S523 }),
  .A2({ S790[90] }),
  .ZN({ S524 })
);
INV_X1 #() 
INV_X1_103_ (
  .A({ S791[94] }),
  .ZN({ S525 })
);
NAND2_X1 #() 
NAND2_X1_31_ (
  .A1({ S525 }),
  .A2({ S790[94] }),
  .ZN({ S526 })
);
INV_X1 #() 
INV_X1_104_ (
  .A({ S790[88] }),
  .ZN({ S527 })
);
NAND2_X1 #() 
NAND2_X1_32_ (
  .A1({ S527 }),
  .A2({ S791[88] }),
  .ZN({ S528 })
);
INV_X1 #() 
INV_X1_105_ (
  .A({ S791[92] }),
  .ZN({ S529 })
);
NAND2_X1 #() 
NAND2_X1_33_ (
  .A1({ S529 }),
  .A2({ S790[92] }),
  .ZN({ S530 })
);
NAND4_X1 #() 
NAND4_X1_13_ (
  .A1({ S528 }),
  .A2({ S530 }),
  .A3({ S524 }),
  .A4({ S526 }),
  .ZN({ S531 })
);
NOR2_X1 #() 
NOR2_X1_11_ (
  .A1({ S522 }),
  .A2({ S531 }),
  .ZN({ S532 })
);
INV_X1 #() 
INV_X1_106_ (
  .A({ S791[27] }),
  .ZN({ S533 })
);
INV_X1 #() 
INV_X1_107_ (
  .A({ S790[29] }),
  .ZN({ S534 })
);
AOI22_X1 #() 
AOI22_X1_29_ (
  .A1({ S533 }),
  .A2({ S790[27] }),
  .B1({ S534 }),
  .B2({ S791[29] }),
  .ZN({ S535 })
);
INV_X1 #() 
INV_X1_108_ (
  .A({ S791[51] }),
  .ZN({ S536 })
);
INV_X1 #() 
INV_X1_109_ (
  .A({ S791[95] }),
  .ZN({ S537 })
);
AOI22_X1 #() 
AOI22_X1_30_ (
  .A1({ S790[51] }),
  .A2({ S536 }),
  .B1({ S537 }),
  .B2({ S790[95] }),
  .ZN({ S538 })
);
INV_X1 #() 
INV_X1_110_ (
  .A({ S791[21] }),
  .ZN({ S539 })
);
INV_X1 #() 
INV_X1_111_ (
  .A({ S791[25] }),
  .ZN({ S540 })
);
AOI22_X1 #() 
AOI22_X1_31_ (
  .A1({ S790[21] }),
  .A2({ S539 }),
  .B1({ S540 }),
  .B2({ S790[25] }),
  .ZN({ S541 })
);
INV_X1 #() 
INV_X1_112_ (
  .A({ S790[23] }),
  .ZN({ S542 })
);
INV_X1 #() 
INV_X1_113_ (
  .A({ S790[27] }),
  .ZN({ S543 })
);
AOI22_X1 #() 
AOI22_X1_32_ (
  .A1({ S791[27] }),
  .A2({ S543 }),
  .B1({ S542 }),
  .B2({ S791[23] }),
  .ZN({ S544 })
);
AND4_X1 #() 
AND4_X1_3_ (
  .A1({ S535 }),
  .A2({ S541 }),
  .A3({ S544 }),
  .A4({ S538 }),
  .ZN({ S545 })
);
INV_X1 #() 
INV_X1_114_ (
  .A({ S790[92] }),
  .ZN({ S546 })
);
NAND2_X1 #() 
NAND2_X1_34_ (
  .A1({ S546 }),
  .A2({ S791[92] }),
  .ZN({ S547 })
);
INV_X1 #() 
INV_X1_115_ (
  .A({ S791[52] }),
  .ZN({ S548 })
);
NAND2_X1 #() 
NAND2_X1_35_ (
  .A1({ S548 }),
  .A2({ S790[52] }),
  .ZN({ S549 })
);
INV_X1 #() 
INV_X1_116_ (
  .A({ S790[50] }),
  .ZN({ S550 })
);
NAND2_X1 #() 
NAND2_X1_36_ (
  .A1({ S550 }),
  .A2({ S791[50] }),
  .ZN({ S551 })
);
INV_X1 #() 
INV_X1_117_ (
  .A({ S790[48] }),
  .ZN({ S552 })
);
NAND2_X1 #() 
NAND2_X1_37_ (
  .A1({ S552 }),
  .A2({ S791[48] }),
  .ZN({ S553 })
);
NAND4_X1 #() 
NAND4_X1_14_ (
  .A1({ S551 }),
  .A2({ S553 }),
  .A3({ S547 }),
  .A4({ S549 }),
  .ZN({ S554 })
);
INV_X1 #() 
INV_X1_118_ (
  .A({ S791[120] }),
  .ZN({ S555 })
);
NAND2_X1 #() 
NAND2_X1_38_ (
  .A1({ S555 }),
  .A2({ S790[120] }),
  .ZN({ S556 })
);
INV_X1 #() 
INV_X1_119_ (
  .A({ S790[118] }),
  .ZN({ S557 })
);
NAND2_X1 #() 
NAND2_X1_39_ (
  .A1({ S557 }),
  .A2({ S791[118] }),
  .ZN({ S558 })
);
INV_X1 #() 
INV_X1_120_ (
  .A({ S791[118] }),
  .ZN({ S559 })
);
NAND2_X1 #() 
NAND2_X1_40_ (
  .A1({ S559 }),
  .A2({ S790[118] }),
  .ZN({ S560 })
);
INV_X1 #() 
INV_X1_121_ (
  .A({ S791[88] }),
  .ZN({ S561 })
);
NAND2_X1 #() 
NAND2_X1_41_ (
  .A1({ S561 }),
  .A2({ S790[88] }),
  .ZN({ S562 })
);
NAND4_X1 #() 
NAND4_X1_15_ (
  .A1({ S560 }),
  .A2({ S562 }),
  .A3({ S556 }),
  .A4({ S558 }),
  .ZN({ S563 })
);
NOR2_X1 #() 
NOR2_X1_12_ (
  .A1({ S554 }),
  .A2({ S563 }),
  .ZN({ S564 })
);
AND2_X1 #() 
AND2_X1_6_ (
  .A1({ S790[86] }),
  .A2({ S791[86] }),
  .ZN({ S565 })
);
NOR2_X1 #() 
NOR2_X1_13_ (
  .A1({ S791[86] }),
  .A2({ S790[86] }),
  .ZN({ S566 })
);
INV_X1 #() 
INV_X1_122_ (
  .A({ S790[30] }),
  .ZN({ S567 })
);
NAND2_X1 #() 
NAND2_X1_42_ (
  .A1({ S567 }),
  .A2({ S791[30] }),
  .ZN({ S568 })
);
INV_X1 #() 
INV_X1_123_ (
  .A({ S790[90] }),
  .ZN({ S569 })
);
NAND2_X1 #() 
NAND2_X1_43_ (
  .A1({ S569 }),
  .A2({ S791[90] }),
  .ZN({ S570 })
);
OAI211_X1 #() 
OAI211_X1_3_ (
  .A({ S570 }),
  .B({ S568 }),
  .C1({ S565 }),
  .C2({ S566 }),
  .ZN({ S571 })
);
INV_X1 #() 
INV_X1_124_ (
  .A({ S791[48] }),
  .ZN({ S572 })
);
NAND2_X1 #() 
NAND2_X1_44_ (
  .A1({ S572 }),
  .A2({ S790[48] }),
  .ZN({ S573 })
);
INV_X1 #() 
INV_X1_125_ (
  .A({ S791[30] }),
  .ZN({ S574 })
);
NAND2_X1 #() 
NAND2_X1_45_ (
  .A1({ S574 }),
  .A2({ S790[30] }),
  .ZN({ S575 })
);
INV_X1 #() 
INV_X1_126_ (
  .A({ S790[52] }),
  .ZN({ S576 })
);
NAND2_X1 #() 
NAND2_X1_46_ (
  .A1({ S576 }),
  .A2({ S791[52] }),
  .ZN({ S577 })
);
INV_X1 #() 
INV_X1_127_ (
  .A({ S791[50] }),
  .ZN({ S578 })
);
NAND2_X1 #() 
NAND2_X1_47_ (
  .A1({ S578 }),
  .A2({ S790[50] }),
  .ZN({ S579 })
);
NAND4_X1 #() 
NAND4_X1_16_ (
  .A1({ S577 }),
  .A2({ S579 }),
  .A3({ S573 }),
  .A4({ S575 }),
  .ZN({ S580 })
);
NOR2_X1 #() 
NOR2_X1_14_ (
  .A1({ S580 }),
  .A2({ S571 }),
  .ZN({ S581 })
);
AND4_X1 #() 
AND4_X1_4_ (
  .A1({ S545 }),
  .A2({ S532 }),
  .A3({ S564 }),
  .A4({ S581 }),
  .ZN({ S582 })
);
INV_X1 #() 
INV_X1_128_ (
  .A({ S790[15] }),
  .ZN({ S583 })
);
INV_X1 #() 
INV_X1_129_ (
  .A({ S791[19] }),
  .ZN({ S584 })
);
AOI22_X1 #() 
AOI22_X1_33_ (
  .A1({ S584 }),
  .A2({ S790[19] }),
  .B1({ S583 }),
  .B2({ S791[15] }),
  .ZN({ S585 })
);
INV_X1 #() 
INV_X1_130_ (
  .A({ S791[7] }),
  .ZN({ S586 })
);
INV_X1 #() 
INV_X1_131_ (
  .A({ S791[49] }),
  .ZN({ S587 })
);
AOI22_X1 #() 
AOI22_X1_34_ (
  .A1({ S790[7] }),
  .A2({ S586 }),
  .B1({ S587 }),
  .B2({ S790[49] }),
  .ZN({ S588 })
);
AND2_X1 #() 
AND2_X1_7_ (
  .A1({ S588 }),
  .A2({ S585 }),
  .ZN({ S589 })
);
XOR2_X1 #() 
XOR2_X1_1_ (
  .A({ S791[1] }),
  .B({ S790[1] }),
  .Z({ S590 })
);
INV_X1 #() 
INV_X1_132_ (
  .A({ S790[111] }),
  .ZN({ S591 })
);
OAI22_X1 #() 
OAI22_X1_14_ (
  .A1({ S591 }),
  .A2({ S791[111] }),
  .B1({ S480 }),
  .B2({ S790[113] }),
  .ZN({ S592 })
);
NOR2_X1 #() 
NOR2_X1_15_ (
  .A1({ S590 }),
  .A2({ S592 }),
  .ZN({ S593 })
);
INV_X1 #() 
INV_X1_133_ (
  .A({ S790[87] }),
  .ZN({ S594 })
);
INV_X1 #() 
INV_X1_134_ (
  .A({ S790[97] }),
  .ZN({ S595 })
);
AOI22_X1 #() 
AOI22_X1_35_ (
  .A1({ S791[97] }),
  .A2({ S595 }),
  .B1({ S594 }),
  .B2({ S791[87] }),
  .ZN({ S596 })
);
INV_X1 #() 
INV_X1_135_ (
  .A({ S791[89] }),
  .ZN({ S597 })
);
INV_X1 #() 
INV_X1_136_ (
  .A({ S790[101] }),
  .ZN({ S598 })
);
AOI22_X1 #() 
AOI22_X1_36_ (
  .A1({ S597 }),
  .A2({ S790[89] }),
  .B1({ S598 }),
  .B2({ S791[101] }),
  .ZN({ S599 })
);
AND2_X1 #() 
AND2_X1_8_ (
  .A1({ S599 }),
  .A2({ S596 }),
  .ZN({ S600 })
);
INV_X1 #() 
INV_X1_137_ (
  .A({ S790[11] }),
  .ZN({ S601 })
);
INV_X1 #() 
INV_X1_138_ (
  .A({ S790[45] }),
  .ZN({ S602 })
);
OAI22_X1 #() 
OAI22_X1_15_ (
  .A1({ S791[11] }),
  .A2({ S601 }),
  .B1({ S602 }),
  .B2({ S791[45] }),
  .ZN({ S603 })
);
OAI22_X1 #() 
OAI22_X1_16_ (
  .A1({ S492 }),
  .A2({ S790[53] }),
  .B1({ S595 }),
  .B2({ S791[97] }),
  .ZN({ S604 })
);
NOR2_X1 #() 
NOR2_X1_16_ (
  .A1({ S603 }),
  .A2({ S604 }),
  .ZN({ S605 })
);
NAND4_X1 #() 
NAND4_X1_17_ (
  .A1({ S593 }),
  .A2({ S589 }),
  .A3({ S600 }),
  .A4({ S605 }),
  .ZN({ S606 })
);
INV_X1 #() 
INV_X1_139_ (
  .A({ S791[9] }),
  .ZN({ S607 })
);
NAND2_X1 #() 
NAND2_X1_48_ (
  .A1({ S607 }),
  .A2({ S790[9] }),
  .ZN({ S608 })
);
OR2_X1 #() 
OR2_X1_1_ (
  .A1({ S607 }),
  .A2({ S790[9] }),
  .ZN({ S609 })
);
INV_X1 #() 
INV_X1_140_ (
  .A({ S791[13] }),
  .ZN({ S610 })
);
INV_X1 #() 
INV_X1_141_ (
  .A({ S790[17] }),
  .ZN({ S611 })
);
AOI22_X1 #() 
AOI22_X1_37_ (
  .A1({ S610 }),
  .A2({ S790[13] }),
  .B1({ S611 }),
  .B2({ S791[17] }),
  .ZN({ S612 })
);
AND3_X1 #() 
AND3_X1_1_ (
  .A1({ S612 }),
  .A2({ S609 }),
  .A3({ S608 }),
  .ZN({ S613 })
);
INV_X1 #() 
INV_X1_142_ (
  .A({ S791[11] }),
  .ZN({ S614 })
);
OAI22_X1 #() 
OAI22_X1_17_ (
  .A1({ S790[7] }),
  .A2({ S586 }),
  .B1({ S614 }),
  .B2({ S790[11] }),
  .ZN({ S615 })
);
OAI22_X1 #() 
OAI22_X1_18_ (
  .A1({ S790[13] }),
  .A2({ S610 }),
  .B1({ S536 }),
  .B2({ S790[51] }),
  .ZN({ S616 })
);
NOR2_X1 #() 
NOR2_X1_17_ (
  .A1({ S615 }),
  .A2({ S616 }),
  .ZN({ S617 })
);
OAI22_X1 #() 
OAI22_X1_19_ (
  .A1({ S542 }),
  .A2({ S791[23] }),
  .B1({ S417 }),
  .B2({ S790[31] }),
  .ZN({ S618 })
);
INV_X1 #() 
INV_X1_143_ (
  .A({ S791[3] }),
  .ZN({ S619 })
);
INV_X1 #() 
INV_X1_144_ (
  .A({ S791[5] }),
  .ZN({ S620 })
);
OAI22_X1 #() 
OAI22_X1_20_ (
  .A1({ S790[3] }),
  .A2({ S619 }),
  .B1({ S620 }),
  .B2({ S790[5] }),
  .ZN({ S621 })
);
NOR2_X1 #() 
NOR2_X1_18_ (
  .A1({ S618 }),
  .A2({ S621 }),
  .ZN({ S622 })
);
INV_X1 #() 
INV_X1_145_ (
  .A({ S791[45] }),
  .ZN({ S623 })
);
OAI22_X1 #() 
OAI22_X1_21_ (
  .A1({ S436 }),
  .A2({ S791[41] }),
  .B1({ S623 }),
  .B2({ S790[45] }),
  .ZN({ S624 })
);
INV_X1 #() 
INV_X1_146_ (
  .A({ S790[47] }),
  .ZN({ S625 })
);
OAI22_X1 #() 
OAI22_X1_22_ (
  .A1({ S540 }),
  .A2({ S790[25] }),
  .B1({ S625 }),
  .B2({ S791[47] }),
  .ZN({ S626 })
);
NOR2_X1 #() 
NOR2_X1_19_ (
  .A1({ S624 }),
  .A2({ S626 }),
  .ZN({ S627 })
);
NAND4_X1 #() 
NAND4_X1_18_ (
  .A1({ S613 }),
  .A2({ S617 }),
  .A3({ S622 }),
  .A4({ S627 }),
  .ZN({ S628 })
);
NOR2_X1 #() 
NOR2_X1_20_ (
  .A1({ S606 }),
  .A2({ S628 }),
  .ZN({ S629 })
);
INV_X1 #() 
INV_X1_147_ (
  .A({ S791[99] }),
  .ZN({ S630 })
);
OAI22_X1 #() 
OAI22_X1_23_ (
  .A1({ S790[95] }),
  .A2({ S537 }),
  .B1({ S630 }),
  .B2({ S790[99] }),
  .ZN({ S631 })
);
INV_X1 #() 
INV_X1_148_ (
  .A({ S790[85] }),
  .ZN({ S632 })
);
INV_X1 #() 
INV_X1_149_ (
  .A({ S790[99] }),
  .ZN({ S633 })
);
OAI22_X1 #() 
OAI22_X1_24_ (
  .A1({ S791[85] }),
  .A2({ S632 }),
  .B1({ S633 }),
  .B2({ S791[99] }),
  .ZN({ S634 })
);
NOR2_X1 #() 
NOR2_X1_21_ (
  .A1({ S631 }),
  .A2({ S634 }),
  .ZN({ S635 })
);
INV_X1 #() 
INV_X1_150_ (
  .A({ S790[103] }),
  .ZN({ S636 })
);
OAI22_X1 #() 
OAI22_X1_25_ (
  .A1({ S636 }),
  .A2({ S791[103] }),
  .B1({ S479 }),
  .B2({ S790[105] }),
  .ZN({ S637 })
);
OAI22_X1 #() 
OAI22_X1_26_ (
  .A1({ S611 }),
  .A2({ S791[17] }),
  .B1({ S539 }),
  .B2({ S790[21] }),
  .ZN({ S638 })
);
NOR2_X1 #() 
NOR2_X1_22_ (
  .A1({ S637 }),
  .A2({ S638 }),
  .ZN({ S639 })
);
INV_X1 #() 
INV_X1_151_ (
  .A({ S791[79] }),
  .ZN({ S640 })
);
OAI22_X1 #() 
OAI22_X1_27_ (
  .A1({ S790[55] }),
  .A2({ S507 }),
  .B1({ S640 }),
  .B2({ S790[79] }),
  .ZN({ S641 })
);
INV_X1 #() 
INV_X1_152_ (
  .A({ S790[79] }),
  .ZN({ S642 })
);
OAI22_X1 #() 
OAI22_X1_28_ (
  .A1({ S791[71] }),
  .A2({ S414 }),
  .B1({ S642 }),
  .B2({ S791[79] }),
  .ZN({ S643 })
);
NOR2_X1 #() 
NOR2_X1_23_ (
  .A1({ S641 }),
  .A2({ S643 }),
  .ZN({ S644 })
);
OAI22_X1 #() 
OAI22_X1_29_ (
  .A1({ S509 }),
  .A2({ S791[67] }),
  .B1({ S495 }),
  .B2({ S790[91] }),
  .ZN({ S645 })
);
OAI22_X1 #() 
OAI22_X1_30_ (
  .A1({ S597 }),
  .A2({ S790[89] }),
  .B1({ S496 }),
  .B2({ S791[93] }),
  .ZN({ S646 })
);
NOR2_X1 #() 
NOR2_X1_24_ (
  .A1({ S645 }),
  .A2({ S646 }),
  .ZN({ S647 })
);
NAND4_X1 #() 
NAND4_X1_19_ (
  .A1({ S644 }),
  .A2({ S647 }),
  .A3({ S635 }),
  .A4({ S639 }),
  .ZN({ S648 })
);
INV_X1 #() 
INV_X1_153_ (
  .A({ S791[43] }),
  .ZN({ S649 })
);
OAI22_X1 #() 
OAI22_X1_31_ (
  .A1({ S790[43] }),
  .A2({ S649 }),
  .B1({ S587 }),
  .B2({ S790[49] }),
  .ZN({ S650 })
);
INV_X1 #() 
INV_X1_154_ (
  .A({ S790[43] }),
  .ZN({ S651 })
);
OAI22_X1 #() 
OAI22_X1_32_ (
  .A1({ S791[37] }),
  .A2({ S489 }),
  .B1({ S651 }),
  .B2({ S791[43] }),
  .ZN({ S652 })
);
NOR2_X1 #() 
NOR2_X1_25_ (
  .A1({ S650 }),
  .A2({ S652 }),
  .ZN({ S653 })
);
NAND2_X1 #() 
NAND2_X1_49_ (
  .A1({ S632 }),
  .A2({ S791[85] }),
  .ZN({ S654 })
);
NAND2_X1 #() 
NAND2_X1_50_ (
  .A1({ S625 }),
  .A2({ S791[47] }),
  .ZN({ S655 })
);
INV_X1 #() 
INV_X1_155_ (
  .A({ S791[39] }),
  .ZN({ S656 })
);
NAND2_X1 #() 
NAND2_X1_51_ (
  .A1({ S656 }),
  .A2({ S790[39] }),
  .ZN({ S657 })
);
NAND2_X1 #() 
NAND2_X1_52_ (
  .A1({ S620 }),
  .A2({ S790[5] }),
  .ZN({ S658 })
);
AND4_X1 #() 
AND4_X1_5_ (
  .A1({ S654 }),
  .A2({ S657 }),
  .A3({ S658 }),
  .A4({ S655 }),
  .ZN({ S659 })
);
INV_X1 #() 
INV_X1_156_ (
  .A({ S790[3] }),
  .ZN({ S660 })
);
OAI22_X1 #() 
OAI22_X1_33_ (
  .A1({ S660 }),
  .A2({ S791[3] }),
  .B1({ S584 }),
  .B2({ S790[19] }),
  .ZN({ S661 })
);
INV_X1 #() 
INV_X1_157_ (
  .A({ S790[0] }),
  .ZN({ S662 })
);
AND2_X1 #() 
AND2_X1_9_ (
  .A1({ S662 }),
  .A2({ S791[0] }),
  .ZN({ S663 })
);
NOR2_X1 #() 
NOR2_X1_26_ (
  .A1({ S662 }),
  .A2({ S791[0] }),
  .ZN({ S664 })
);
NOR3_X1 #() 
NOR3_X1_4_ (
  .A1({ S661 }),
  .A2({ S663 }),
  .A3({ S664 }),
  .ZN({ S665 })
);
OAI22_X1 #() 
OAI22_X1_34_ (
  .A1({ S583 }),
  .A2({ S791[15] }),
  .B1({ S656 }),
  .B2({ S790[39] }),
  .ZN({ S666 })
);
INV_X1 #() 
INV_X1_158_ (
  .A({ S791[35] }),
  .ZN({ S667 })
);
OAI22_X1 #() 
OAI22_X1_35_ (
  .A1({ S534 }),
  .A2({ S791[29] }),
  .B1({ S667 }),
  .B2({ S790[35] }),
  .ZN({ S668 })
);
NOR2_X1 #() 
NOR2_X1_27_ (
  .A1({ S666 }),
  .A2({ S668 }),
  .ZN({ S669 })
);
NAND4_X1 #() 
NAND4_X1_20_ (
  .A1({ S665 }),
  .A2({ S669 }),
  .A3({ S659 }),
  .A4({ S653 }),
  .ZN({ S670 })
);
NOR2_X1 #() 
NOR2_X1_28_ (
  .A1({ S648 }),
  .A2({ S670 }),
  .ZN({ S671 })
);
INV_X1 #() 
INV_X1_159_ (
  .A({ S791[103] }),
  .ZN({ S672 })
);
OAI22_X1 #() 
OAI22_X1_36_ (
  .A1({ S598 }),
  .A2({ S791[101] }),
  .B1({ S672 }),
  .B2({ S790[103] }),
  .ZN({ S673 })
);
INV_X1 #() 
INV_X1_160_ (
  .A({ S791[111] }),
  .ZN({ S674 })
);
OAI22_X1 #() 
OAI22_X1_37_ (
  .A1({ S460 }),
  .A2({ S791[109] }),
  .B1({ S674 }),
  .B2({ S790[111] }),
  .ZN({ S675 })
);
NOR2_X1 #() 
NOR2_X1_29_ (
  .A1({ S673 }),
  .A2({ S675 }),
  .ZN({ S676 })
);
NAND2_X1 #() 
NAND2_X1_53_ (
  .A1({ S791[112] }),
  .A2({ S790[112] }),
  .ZN({ S677 })
);
OR2_X1 #() 
OR2_X1_2_ (
  .A1({ S791[112] }),
  .A2({ S790[112] }),
  .ZN({ S678 })
);
NAND2_X1 #() 
NAND2_X1_54_ (
  .A1({ S791[2] }),
  .A2({ S790[2] }),
  .ZN({ S679 })
);
OR2_X1 #() 
OR2_X1_3_ (
  .A1({ S791[2] }),
  .A2({ S790[2] }),
  .ZN({ S680 })
);
AOI22_X1 #() 
AOI22_X1_38_ (
  .A1({ S679 }),
  .A2({ S680 }),
  .B1({ S678 }),
  .B2({ S677 }),
  .ZN({ S681 })
);
OAI22_X1 #() 
OAI22_X1_38_ (
  .A1({ S477 }),
  .A2({ S791[121] }),
  .B1({ S456 }),
  .B2({ S790[123] }),
  .ZN({ S682 })
);
OAI22_X1 #() 
OAI22_X1_39_ (
  .A1({ S790[120] }),
  .A2({ S555 }),
  .B1({ S450 }),
  .B2({ S790[125] }),
  .ZN({ S683 })
);
NOR2_X1 #() 
NOR2_X1_30_ (
  .A1({ S682 }),
  .A2({ S683 }),
  .ZN({ S684 })
);
INV_X1 #() 
INV_X1_161_ (
  .A({ S790[107] }),
  .ZN({ S685 })
);
NAND2_X1 #() 
NAND2_X1_55_ (
  .A1({ S685 }),
  .A2({ S791[107] }),
  .ZN({ S686 })
);
INV_X1 #() 
INV_X1_162_ (
  .A({ S791[107] }),
  .ZN({ S687 })
);
NAND2_X1 #() 
NAND2_X1_56_ (
  .A1({ S687 }),
  .A2({ S790[107] }),
  .ZN({ S688 })
);
INV_X1 #() 
INV_X1_163_ (
  .A({ S790[119] }),
  .ZN({ S689 })
);
NAND2_X1 #() 
NAND2_X1_57_ (
  .A1({ S689 }),
  .A2({ S791[119] }),
  .ZN({ S690 })
);
INV_X1 #() 
INV_X1_164_ (
  .A({ S791[119] }),
  .ZN({ S691 })
);
NAND2_X1 #() 
NAND2_X1_58_ (
  .A1({ S691 }),
  .A2({ S790[119] }),
  .ZN({ S692 })
);
AND4_X1 #() 
AND4_X1_6_ (
  .A1({ S686 }),
  .A2({ S690 }),
  .A3({ S692 }),
  .A4({ S688 }),
  .ZN({ S693 })
);
NAND4_X1 #() 
NAND4_X1_21_ (
  .A1({ S684 }),
  .A2({ S693 }),
  .A3({ S676 }),
  .A4({ S681 }),
  .ZN({ S694 })
);
NAND2_X1 #() 
NAND2_X1_59_ (
  .A1({ S791[114] }),
  .A2({ S790[114] }),
  .ZN({ S695 })
);
OR2_X1 #() 
OR2_X1_4_ (
  .A1({ S791[114] }),
  .A2({ S790[114] }),
  .ZN({ S696 })
);
NAND2_X1 #() 
NAND2_X1_60_ (
  .A1({ S791[104] }),
  .A2({ S790[104] }),
  .ZN({ S697 })
);
OR2_X1 #() 
OR2_X1_5_ (
  .A1({ S791[104] }),
  .A2({ S790[104] }),
  .ZN({ S698 })
);
AOI22_X1 #() 
AOI22_X1_39_ (
  .A1({ S697 }),
  .A2({ S698 }),
  .B1({ S696 }),
  .B2({ S695 }),
  .ZN({ S699 })
);
INV_X1 #() 
INV_X1_165_ (
  .A({ S790[35] }),
  .ZN({ S700 })
);
OAI22_X1 #() 
OAI22_X1_40_ (
  .A1({ S700 }),
  .A2({ S791[35] }),
  .B1({ S402 }),
  .B2({ S790[73] }),
  .ZN({ S701 })
);
INV_X1 #() 
INV_X1_166_ (
  .A({ S790[65] }),
  .ZN({ S702 })
);
OAI22_X1 #() 
OAI22_X1_41_ (
  .A1({ S702 }),
  .A2({ S791[65] }),
  .B1({ S405 }),
  .B2({ S790[69] }),
  .ZN({ S703 })
);
NOR2_X1 #() 
NOR2_X1_31_ (
  .A1({ S701 }),
  .A2({ S703 }),
  .ZN({ S704 })
);
NAND2_X1 #() 
NAND2_X1_61_ (
  .A1({ S791[38] }),
  .A2({ S790[38] }),
  .ZN({ S705 })
);
OR2_X1 #() 
OR2_X1_6_ (
  .A1({ S791[38] }),
  .A2({ S790[38] }),
  .ZN({ S706 })
);
NAND2_X1 #() 
NAND2_X1_62_ (
  .A1({ S791[20] }),
  .A2({ S790[20] }),
  .ZN({ S707 })
);
OR2_X1 #() 
OR2_X1_7_ (
  .A1({ S791[20] }),
  .A2({ S790[20] }),
  .ZN({ S708 })
);
AOI22_X1 #() 
AOI22_X1_40_ (
  .A1({ S707 }),
  .A2({ S708 }),
  .B1({ S706 }),
  .B2({ S705 }),
  .ZN({ S709 })
);
NAND2_X1 #() 
NAND2_X1_63_ (
  .A1({ S791[108] }),
  .A2({ S790[108] }),
  .ZN({ S710 })
);
OR2_X1 #() 
OR2_X1_8_ (
  .A1({ S791[108] }),
  .A2({ S790[108] }),
  .ZN({ S711 })
);
NAND2_X1 #() 
NAND2_X1_64_ (
  .A1({ S791[102] }),
  .A2({ S790[102] }),
  .ZN({ S712 })
);
OR2_X1 #() 
OR2_X1_9_ (
  .A1({ S791[102] }),
  .A2({ S790[102] }),
  .ZN({ S713 })
);
AOI22_X1 #() 
AOI22_X1_41_ (
  .A1({ S712 }),
  .A2({ S713 }),
  .B1({ S711 }),
  .B2({ S710 }),
  .ZN({ S714 })
);
NAND4_X1 #() 
NAND4_X1_22_ (
  .A1({ S704 }),
  .A2({ S699 }),
  .A3({ S709 }),
  .A4({ S714 }),
  .ZN({ S715 })
);
NOR2_X1 #() 
NOR2_X1_32_ (
  .A1({ S694 }),
  .A2({ S715 }),
  .ZN({ S716 })
);
NAND4_X1 #() 
NAND4_X1_23_ (
  .A1({ S629 }),
  .A2({ S671 }),
  .A3({ S582 }),
  .A4({ S716 }),
  .ZN({ S717 })
);
NOR3_X1 #() 
NOR3_X1_5_ (
  .A1({ S717 }),
  .A2({ S448 }),
  .A3({ S513 }),
  .ZN({ S788 })
);
XNOR2_X1 #() 
XNOR2_X1_8_ (
  .A({ S792[72] }),
  .B({ S787[72] }),
  .ZN({ S718 })
);
XNOR2_X1 #() 
XNOR2_X1_9_ (
  .A({ S792[18] }),
  .B({ S787[18] }),
  .ZN({ S719 })
);
XNOR2_X1 #() 
XNOR2_X1_10_ (
  .A({ S792[20] }),
  .B({ S787[20] }),
  .ZN({ S720 })
);
NAND3_X1 #() 
NAND3_X1_4_ (
  .A1({ S718 }),
  .A2({ S719 }),
  .A3({ S720 }),
  .ZN({ S721 })
);
XNOR2_X1 #() 
XNOR2_X1_11_ (
  .A({ S792[70] }),
  .B({ S787[70] }),
  .ZN({ S722 })
);
XNOR2_X1 #() 
XNOR2_X1_12_ (
  .A({ S792[16] }),
  .B({ S787[16] }),
  .ZN({ S723 })
);
XNOR2_X1 #() 
XNOR2_X1_13_ (
  .A({ S792[30] }),
  .B({ S787[30] }),
  .ZN({ S724 })
);
XNOR2_X1 #() 
XNOR2_X1_14_ (
  .A({ S792[36] }),
  .B({ S787[36] }),
  .ZN({ S725 })
);
NAND4_X1 #() 
NAND4_X1_24_ (
  .A1({ S724 }),
  .A2({ S725 }),
  .A3({ S722 }),
  .A4({ S723 }),
  .ZN({ S726 })
);
INV_X1 #() 
INV_X1_167_ (
  .A({ S792[56] }),
  .ZN({ S727 })
);
INV_X1 #() 
INV_X1_168_ (
  .A({ S787[60] }),
  .ZN({ S728 })
);
AOI22_X1 #() 
AOI22_X1_42_ (
  .A1({ S727 }),
  .A2({ S787[56] }),
  .B1({ S728 }),
  .B2({ S792[60] }),
  .ZN({ S729 })
);
INV_X1 #() 
INV_X1_169_ (
  .A({ S792[60] }),
  .ZN({ S730 })
);
INV_X1 #() 
INV_X1_170_ (
  .A({ S787[66] }),
  .ZN({ S731 })
);
AOI22_X1 #() 
AOI22_X1_43_ (
  .A1({ S730 }),
  .A2({ S787[60] }),
  .B1({ S731 }),
  .B2({ S792[66] }),
  .ZN({ S732 })
);
INV_X1 #() 
INV_X1_171_ (
  .A({ S787[76] }),
  .ZN({ S733 })
);
AOI21_X1 #() 
AOI21_X1_2_ (
  .A({ S309 }),
  .B1({ S792[76] }),
  .B2({ S733 }),
  .ZN({ S734 })
);
INV_X1 #() 
INV_X1_172_ (
  .A({ S787[56] }),
  .ZN({ S735 })
);
INV_X1 #() 
INV_X1_173_ (
  .A({ S792[76] }),
  .ZN({ S736 })
);
AOI22_X1 #() 
AOI22_X1_44_ (
  .A1({ S736 }),
  .A2({ S787[76] }),
  .B1({ S735 }),
  .B2({ S792[56] }),
  .ZN({ S737 })
);
NAND4_X1 #() 
NAND4_X1_25_ (
  .A1({ S737 }),
  .A2({ S732 }),
  .A3({ S729 }),
  .A4({ S734 }),
  .ZN({ S738 })
);
NOR3_X1 #() 
NOR3_X1_6_ (
  .A1({ S726 }),
  .A2({ S738 }),
  .A3({ S721 }),
  .ZN({ S739 })
);
INV_X1 #() 
INV_X1_174_ (
  .A({ S792[88] }),
  .ZN({ S740 })
);
INV_X1 #() 
INV_X1_175_ (
  .A({ S787[92] }),
  .ZN({ S741 })
);
AOI22_X1 #() 
AOI22_X1_45_ (
  .A1({ S740 }),
  .A2({ S787[88] }),
  .B1({ S741 }),
  .B2({ S792[92] }),
  .ZN({ S742 })
);
INV_X1 #() 
INV_X1_176_ (
  .A({ S792[22] }),
  .ZN({ S743 })
);
INV_X1 #() 
INV_X1_177_ (
  .A({ S787[40] }),
  .ZN({ S744 })
);
AOI22_X1 #() 
AOI22_X1_46_ (
  .A1({ S743 }),
  .A2({ S787[22] }),
  .B1({ S744 }),
  .B2({ S792[40] }),
  .ZN({ S745 })
);
INV_X1 #() 
INV_X1_178_ (
  .A({ S792[86] }),
  .ZN({ S746 })
);
INV_X1 #() 
INV_X1_179_ (
  .A({ S787[98] }),
  .ZN({ S747 })
);
AOI22_X1 #() 
AOI22_X1_47_ (
  .A1({ S746 }),
  .A2({ S787[86] }),
  .B1({ S747 }),
  .B2({ S792[98] }),
  .ZN({ S748 })
);
INV_X1 #() 
INV_X1_180_ (
  .A({ S787[88] }),
  .ZN({ S749 })
);
INV_X1 #() 
INV_X1_181_ (
  .A({ S792[98] }),
  .ZN({ S750 })
);
AOI22_X1 #() 
AOI22_X1_48_ (
  .A1({ S750 }),
  .A2({ S787[98] }),
  .B1({ S749 }),
  .B2({ S792[88] }),
  .ZN({ S751 })
);
AND4_X1 #() 
AND4_X1_7_ (
  .A1({ S742 }),
  .A2({ S748 }),
  .A3({ S751 }),
  .A4({ S745 }),
  .ZN({ S752 })
);
INV_X1 #() 
INV_X1_182_ (
  .A({ S792[94] }),
  .ZN({ S753 })
);
INV_X1 #() 
INV_X1_183_ (
  .A({ S787[100] }),
  .ZN({ S754 })
);
AOI22_X1 #() 
AOI22_X1_49_ (
  .A1({ S753 }),
  .A2({ S787[94] }),
  .B1({ S754 }),
  .B2({ S792[100] }),
  .ZN({ S755 })
);
INV_X1 #() 
INV_X1_184_ (
  .A({ S792[92] }),
  .ZN({ S756 })
);
INV_X1 #() 
INV_X1_185_ (
  .A({ S792[100] }),
  .ZN({ S757 })
);
AOI22_X1 #() 
AOI22_X1_50_ (
  .A1({ S787[92] }),
  .A2({ S756 }),
  .B1({ S757 }),
  .B2({ S787[100] }),
  .ZN({ S758 })
);
INV_X1 #() 
INV_X1_186_ (
  .A({ S792[40] }),
  .ZN({ S759 })
);
INV_X1 #() 
INV_X1_187_ (
  .A({ S787[96] }),
  .ZN({ S760 })
);
AOI22_X1 #() 
AOI22_X1_51_ (
  .A1({ S759 }),
  .A2({ S787[40] }),
  .B1({ S760 }),
  .B2({ S792[96] }),
  .ZN({ S761 })
);
INV_X1 #() 
INV_X1_188_ (
  .A({ S787[94] }),
  .ZN({ S762 })
);
INV_X1 #() 
INV_X1_189_ (
  .A({ S792[96] }),
  .ZN({ S763 })
);
AOI22_X1 #() 
AOI22_X1_52_ (
  .A1({ S763 }),
  .A2({ S787[96] }),
  .B1({ S762 }),
  .B2({ S792[94] }),
  .ZN({ S764 })
);
AND4_X1 #() 
AND4_X1_8_ (
  .A1({ S755 }),
  .A2({ S761 }),
  .A3({ S764 }),
  .A4({ S758 }),
  .ZN({ S765 })
);
AND2_X1 #() 
AND2_X1_10_ (
  .A1({ S787[68] }),
  .A2({ S792[68] }),
  .ZN({ S766 })
);
NOR2_X1 #() 
NOR2_X1_33_ (
  .A1({ S792[68] }),
  .A2({ S787[68] }),
  .ZN({ S767 })
);
INV_X1 #() 
INV_X1_190_ (
  .A({ S792[74] }),
  .ZN({ S768 })
);
NAND2_X1 #() 
NAND2_X1_65_ (
  .A1({ S768 }),
  .A2({ S787[74] }),
  .ZN({ S769 })
);
INV_X1 #() 
INV_X1_191_ (
  .A({ S787[34] }),
  .ZN({ S770 })
);
NAND2_X1 #() 
NAND2_X1_66_ (
  .A1({ S770 }),
  .A2({ S792[34] }),
  .ZN({ S771 })
);
OAI211_X1 #() 
OAI211_X1_4_ (
  .A({ S771 }),
  .B({ S769 }),
  .C1({ S766 }),
  .C2({ S767 }),
  .ZN({ S772 })
);
AND2_X1 #() 
AND2_X1_11_ (
  .A1({ S787[80] }),
  .A2({ S792[80] }),
  .ZN({ S773 })
);
NOR2_X1 #() 
NOR2_X1_34_ (
  .A1({ S792[80] }),
  .A2({ S787[80] }),
  .ZN({ S774 })
);
INV_X1 #() 
INV_X1_192_ (
  .A({ S787[74] }),
  .ZN({ S775 })
);
NAND2_X1 #() 
NAND2_X1_67_ (
  .A1({ S775 }),
  .A2({ S792[74] }),
  .ZN({ S776 })
);
INV_X1 #() 
INV_X1_193_ (
  .A({ S792[66] }),
  .ZN({ S777 })
);
NAND2_X1 #() 
NAND2_X1_68_ (
  .A1({ S777 }),
  .A2({ S787[66] }),
  .ZN({ S778 })
);
OAI211_X1 #() 
OAI211_X1_5_ (
  .A({ S778 }),
  .B({ S776 }),
  .C1({ S773 }),
  .C2({ S774 }),
  .ZN({ S779 })
);
NOR2_X1 #() 
NOR2_X1_35_ (
  .A1({ S772 }),
  .A2({ S779 }),
  .ZN({ S780 })
);
INV_X1 #() 
INV_X1_194_ (
  .A({ S787[82] }),
  .ZN({ S781 })
);
INV_X1 #() 
INV_X1_195_ (
  .A({ S792[84] }),
  .ZN({ S782 })
);
AOI22_X1 #() 
AOI22_X1_53_ (
  .A1({ S782 }),
  .A2({ S787[84] }),
  .B1({ S781 }),
  .B2({ S792[82] }),
  .ZN({ S783 })
);
INV_X1 #() 
INV_X1_196_ (
  .A({ S792[82] }),
  .ZN({ S784 })
);
INV_X1 #() 
INV_X1_197_ (
  .A({ S787[86] }),
  .ZN({ S785 })
);
AOI22_X1 #() 
AOI22_X1_54_ (
  .A1({ S784 }),
  .A2({ S787[82] }),
  .B1({ S785 }),
  .B2({ S792[86] }),
  .ZN({ S0 })
);
INV_X1 #() 
INV_X1_198_ (
  .A({ S792[34] }),
  .ZN({ S1 })
);
INV_X1 #() 
INV_X1_199_ (
  .A({ S787[58] }),
  .ZN({ S2 })
);
AOI22_X1 #() 
AOI22_X1_55_ (
  .A1({ S1 }),
  .A2({ S787[34] }),
  .B1({ S2 }),
  .B2({ S792[58] }),
  .ZN({ S3 })
);
INV_X1 #() 
INV_X1_200_ (
  .A({ S792[58] }),
  .ZN({ S4 })
);
INV_X1 #() 
INV_X1_201_ (
  .A({ S787[84] }),
  .ZN({ S5 })
);
AOI22_X1 #() 
AOI22_X1_56_ (
  .A1({ S4 }),
  .A2({ S787[58] }),
  .B1({ S5 }),
  .B2({ S792[84] }),
  .ZN({ S6 })
);
AND4_X1 #() 
AND4_X1_9_ (
  .A1({ S783 }),
  .A2({ S3 }),
  .A3({ S6 }),
  .A4({ S0 }),
  .ZN({ S7 })
);
AND4_X1 #() 
AND4_X1_10_ (
  .A1({ S752 }),
  .A2({ S7 }),
  .A3({ S765 }),
  .A4({ S780 }),
  .ZN({ S8 })
);
INV_X1 #() 
INV_X1_202_ (
  .A({ S787[57] }),
  .ZN({ S9 })
);
NAND2_X1 #() 
NAND2_X1_69_ (
  .A1({ S9 }),
  .A2({ S792[57] }),
  .ZN({ S10 })
);
INV_X1 #() 
INV_X1_203_ (
  .A({ S787[73] }),
  .ZN({ S11 })
);
NAND2_X1 #() 
NAND2_X1_70_ (
  .A1({ S11 }),
  .A2({ S792[73] }),
  .ZN({ S12 })
);
INV_X1 #() 
INV_X1_204_ (
  .A({ S792[79] }),
  .ZN({ S13 })
);
NAND2_X1 #() 
NAND2_X1_71_ (
  .A1({ S13 }),
  .A2({ S787[79] }),
  .ZN({ S14 })
);
INV_X1 #() 
INV_X1_205_ (
  .A({ S792[71] }),
  .ZN({ S15 })
);
NAND2_X1 #() 
NAND2_X1_72_ (
  .A1({ S15 }),
  .A2({ S787[71] }),
  .ZN({ S16 })
);
NAND4_X1 #() 
NAND4_X1_26_ (
  .A1({ S14 }),
  .A2({ S16 }),
  .A3({ S10 }),
  .A4({ S12 }),
  .ZN({ S17 })
);
INV_X1 #() 
INV_X1_206_ (
  .A({ S787[63] }),
  .ZN({ S18 })
);
NAND2_X1 #() 
NAND2_X1_73_ (
  .A1({ S18 }),
  .A2({ S792[63] }),
  .ZN({ S19 })
);
INV_X1 #() 
INV_X1_207_ (
  .A({ S792[63] }),
  .ZN({ S20 })
);
NAND2_X1 #() 
NAND2_X1_74_ (
  .A1({ S20 }),
  .A2({ S787[63] }),
  .ZN({ S21 })
);
INV_X1 #() 
INV_X1_208_ (
  .A({ S792[61] }),
  .ZN({ S22 })
);
NAND2_X1 #() 
NAND2_X1_75_ (
  .A1({ S22 }),
  .A2({ S787[61] }),
  .ZN({ S23 })
);
INV_X1 #() 
INV_X1_209_ (
  .A({ S787[65] }),
  .ZN({ S24 })
);
NAND2_X1 #() 
NAND2_X1_76_ (
  .A1({ S24 }),
  .A2({ S792[65] }),
  .ZN({ S25 })
);
NAND4_X1 #() 
NAND4_X1_27_ (
  .A1({ S23 }),
  .A2({ S25 }),
  .A3({ S19 }),
  .A4({ S21 }),
  .ZN({ S26 })
);
NOR2_X1 #() 
NOR2_X1_36_ (
  .A1({ S17 }),
  .A2({ S26 }),
  .ZN({ S27 })
);
INV_X1 #() 
INV_X1_210_ (
  .A({ S787[1] }),
  .ZN({ S28 })
);
INV_X1 #() 
INV_X1_211_ (
  .A({ S787[15] }),
  .ZN({ S29 })
);
AOI22_X1 #() 
AOI22_X1_57_ (
  .A1({ S792[15] }),
  .A2({ S29 }),
  .B1({ S28 }),
  .B2({ S792[1] }),
  .ZN({ S30 })
);
XNOR2_X1 #() 
XNOR2_X1_15_ (
  .A({ S792[0] }),
  .B({ S787[0] }),
  .ZN({ S31 })
);
INV_X1 #() 
INV_X1_212_ (
  .A({ S792[69] }),
  .ZN({ S32 })
);
INV_X1 #() 
INV_X1_213_ (
  .A({ S787[81] }),
  .ZN({ S33 })
);
AOI22_X1 #() 
AOI22_X1_58_ (
  .A1({ S32 }),
  .A2({ S787[69] }),
  .B1({ S33 }),
  .B2({ S792[81] }),
  .ZN({ S34 })
);
INV_X1 #() 
INV_X1_214_ (
  .A({ S792[13] }),
  .ZN({ S35 })
);
INV_X1 #() 
INV_X1_215_ (
  .A({ S787[21] }),
  .ZN({ S36 })
);
AOI22_X1 #() 
AOI22_X1_59_ (
  .A1({ S35 }),
  .A2({ S787[13] }),
  .B1({ S36 }),
  .B2({ S792[21] }),
  .ZN({ S37 })
);
AND4_X1 #() 
AND4_X1_11_ (
  .A1({ S30 }),
  .A2({ S37 }),
  .A3({ S31 }),
  .A4({ S34 }),
  .ZN({ S38 })
);
INV_X1 #() 
INV_X1_216_ (
  .A({ S792[2] }),
  .ZN({ S39 })
);
NAND2_X1 #() 
NAND2_X1_77_ (
  .A1({ S39 }),
  .A2({ S787[2] }),
  .ZN({ S40 })
);
INV_X1 #() 
INV_X1_217_ (
  .A({ S792[42] }),
  .ZN({ S41 })
);
NAND2_X1 #() 
NAND2_X1_78_ (
  .A1({ S41 }),
  .A2({ S787[42] }),
  .ZN({ S42 })
);
AND2_X1 #() 
AND2_X1_12_ (
  .A1({ S787[4] }),
  .A2({ S792[4] }),
  .ZN({ S43 })
);
NOR2_X1 #() 
NOR2_X1_37_ (
  .A1({ S792[4] }),
  .A2({ S787[4] }),
  .ZN({ S44 })
);
OAI211_X1 #() 
OAI211_X1_6_ (
  .A({ S42 }),
  .B({ S40 }),
  .C1({ S43 }),
  .C2({ S44 }),
  .ZN({ S45 })
);
AND2_X1 #() 
AND2_X1_13_ (
  .A1({ S787[90] }),
  .A2({ S792[90] }),
  .ZN({ S46 })
);
NOR2_X1 #() 
NOR2_X1_38_ (
  .A1({ S792[90] }),
  .A2({ S787[90] }),
  .ZN({ S47 })
);
INV_X1 #() 
INV_X1_218_ (
  .A({ S787[42] }),
  .ZN({ S48 })
);
NAND2_X1 #() 
NAND2_X1_79_ (
  .A1({ S48 }),
  .A2({ S792[42] }),
  .ZN({ S49 })
);
INV_X1 #() 
INV_X1_219_ (
  .A({ S787[2] }),
  .ZN({ S50 })
);
NAND2_X1 #() 
NAND2_X1_80_ (
  .A1({ S50 }),
  .A2({ S792[2] }),
  .ZN({ S51 })
);
OAI211_X1 #() 
OAI211_X1_7_ (
  .A({ S51 }),
  .B({ S49 }),
  .C1({ S46 }),
  .C2({ S47 }),
  .ZN({ S52 })
);
NOR2_X1 #() 
NOR2_X1_39_ (
  .A1({ S45 }),
  .A2({ S52 }),
  .ZN({ S53 })
);
AND2_X1 #() 
AND2_X1_14_ (
  .A1({ S787[44] }),
  .A2({ S792[44] }),
  .ZN({ S54 })
);
NOR2_X1 #() 
NOR2_X1_40_ (
  .A1({ S792[44] }),
  .A2({ S787[44] }),
  .ZN({ S55 })
);
INV_X1 #() 
INV_X1_220_ (
  .A({ S787[22] }),
  .ZN({ S56 })
);
NAND2_X1 #() 
NAND2_X1_81_ (
  .A1({ S56 }),
  .A2({ S792[22] }),
  .ZN({ S57 })
);
INV_X1 #() 
INV_X1_221_ (
  .A({ S792[55] }),
  .ZN({ S58 })
);
NAND2_X1 #() 
NAND2_X1_82_ (
  .A1({ S58 }),
  .A2({ S787[55] }),
  .ZN({ S59 })
);
OAI211_X1 #() 
OAI211_X1_8_ (
  .A({ S59 }),
  .B({ S57 }),
  .C1({ S54 }),
  .C2({ S55 }),
  .ZN({ S60 })
);
INV_X1 #() 
INV_X1_222_ (
  .A({ S787[32] }),
  .ZN({ S61 })
);
NAND2_X1 #() 
NAND2_X1_83_ (
  .A1({ S61 }),
  .A2({ S792[32] }),
  .ZN({ S62 })
);
INV_X1 #() 
INV_X1_223_ (
  .A({ S792[32] }),
  .ZN({ S63 })
);
NAND2_X1 #() 
NAND2_X1_84_ (
  .A1({ S63 }),
  .A2({ S787[32] }),
  .ZN({ S64 })
);
AND2_X1 #() 
AND2_X1_15_ (
  .A1({ S787[46] }),
  .A2({ S792[46] }),
  .ZN({ S65 })
);
NOR2_X1 #() 
NOR2_X1_41_ (
  .A1({ S792[46] }),
  .A2({ S787[46] }),
  .ZN({ S66 })
);
OAI211_X1 #() 
OAI211_X1_9_ (
  .A({ S64 }),
  .B({ S62 }),
  .C1({ S65 }),
  .C2({ S66 }),
  .ZN({ S67 })
);
NOR2_X1 #() 
NOR2_X1_42_ (
  .A1({ S60 }),
  .A2({ S67 }),
  .ZN({ S68 })
);
AND4_X1 #() 
AND4_X1_12_ (
  .A1({ S38 }),
  .A2({ S27 }),
  .A3({ S53 }),
  .A4({ S68 }),
  .ZN({ S69 })
);
NAND3_X1 #() 
NAND3_X1_5_ (
  .A1({ S8 }),
  .A2({ S739 }),
  .A3({ S69 }),
  .ZN({ S70 })
);
INV_X1 #() 
INV_X1_224_ (
  .A({ S787[39] }),
  .ZN({ S71 })
);
INV_X1 #() 
INV_X1_225_ (
  .A({ S787[5] }),
  .ZN({ S72 })
);
NAND2_X1 #() 
NAND2_X1_85_ (
  .A1({ S72 }),
  .A2({ S792[5] }),
  .ZN({ S73 })
);
OAI221_X1 #() 
OAI221_X1_2_ (
  .A({ S73 }),
  .B1({ S792[39] }),
  .B2({ S71 }),
  .C1({ S29 }),
  .C2({ S792[15] }),
  .ZN({ S74 })
);
INV_X1 #() 
INV_X1_226_ (
  .A({ S792[122] }),
  .ZN({ S75 })
);
NAND2_X1 #() 
NAND2_X1_86_ (
  .A1({ S75 }),
  .A2({ S787[122] }),
  .ZN({ S76 })
);
INV_X1 #() 
INV_X1_227_ (
  .A({ S787[35] }),
  .ZN({ S77 })
);
INV_X1 #() 
INV_X1_228_ (
  .A({ S787[41] }),
  .ZN({ S78 })
);
AOI22_X1 #() 
AOI22_X1_60_ (
  .A1({ S792[41] }),
  .A2({ S78 }),
  .B1({ S77 }),
  .B2({ S792[35] }),
  .ZN({ S79 })
);
OAI211_X1 #() 
OAI211_X1_10_ (
  .A({ S79 }),
  .B({ S76 }),
  .C1({ S787[71] }),
  .C2({ S15 }),
  .ZN({ S80 })
);
INV_X1 #() 
INV_X1_229_ (
  .A({ S787[124] }),
  .ZN({ S81 })
);
INV_X1 #() 
INV_X1_230_ (
  .A({ S787[125] }),
  .ZN({ S82 })
);
AOI22_X1 #() 
AOI22_X1_61_ (
  .A1({ S792[125] }),
  .A2({ S82 }),
  .B1({ S81 }),
  .B2({ S792[124] }),
  .ZN({ S83 })
);
OAI221_X1 #() 
OAI221_X1_3_ (
  .A({ S83 }),
  .B1({ S792[124] }),
  .B2({ S81 }),
  .C1({ S787[122] }),
  .C2({ S75 }),
  .ZN({ S84 })
);
NOR3_X1 #() 
NOR3_X1_7_ (
  .A1({ S84 }),
  .A2({ S80 }),
  .A3({ S74 }),
  .ZN({ S85 })
);
XNOR2_X1 #() 
XNOR2_X1_16_ (
  .A({ S792[48] }),
  .B({ S787[48] }),
  .ZN({ S86 })
);
INV_X1 #() 
INV_X1_231_ (
  .A({ S792[113] }),
  .ZN({ S87 })
);
INV_X1 #() 
INV_X1_232_ (
  .A({ S787[117] }),
  .ZN({ S88 })
);
AOI22_X1 #() 
AOI22_X1_62_ (
  .A1({ S87 }),
  .A2({ S787[113] }),
  .B1({ S88 }),
  .B2({ S792[117] }),
  .ZN({ S89 })
);
XNOR2_X1 #() 
XNOR2_X1_17_ (
  .A({ S792[24] }),
  .B({ S787[24] }),
  .ZN({ S90 })
);
XNOR2_X1 #() 
XNOR2_X1_18_ (
  .A({ S792[50] }),
  .B({ S787[50] }),
  .ZN({ S91 })
);
NAND4_X1 #() 
NAND4_X1_28_ (
  .A1({ S90 }),
  .A2({ S91 }),
  .A3({ S86 }),
  .A4({ S89 }),
  .ZN({ S92 })
);
XNOR2_X1 #() 
XNOR2_X1_19_ (
  .A({ S792[107] }),
  .B({ S787[107] }),
  .ZN({ S93 })
);
INV_X1 #() 
INV_X1_233_ (
  .A({ S787[119] }),
  .ZN({ S94 })
);
INV_X1 #() 
INV_X1_234_ (
  .A({ S792[123] }),
  .ZN({ S95 })
);
AOI22_X1 #() 
AOI22_X1_63_ (
  .A1({ S95 }),
  .A2({ S787[123] }),
  .B1({ S94 }),
  .B2({ S792[119] }),
  .ZN({ S96 })
);
XNOR2_X1 #() 
XNOR2_X1_20_ (
  .A({ S792[115] }),
  .B({ S787[115] }),
  .ZN({ S97 })
);
INV_X1 #() 
INV_X1_235_ (
  .A({ S792[125] }),
  .ZN({ S98 })
);
INV_X1 #() 
INV_X1_236_ (
  .A({ S792[127] }),
  .ZN({ S99 })
);
AOI22_X1 #() 
AOI22_X1_64_ (
  .A1({ S787[125] }),
  .A2({ S98 }),
  .B1({ S99 }),
  .B2({ S787[127] }),
  .ZN({ S100 })
);
NAND4_X1 #() 
NAND4_X1_29_ (
  .A1({ S97 }),
  .A2({ S100 }),
  .A3({ S93 }),
  .A4({ S96 }),
  .ZN({ S101 })
);
NOR2_X1 #() 
NOR2_X1_43_ (
  .A1({ S92 }),
  .A2({ S101 }),
  .ZN({ S102 })
);
INV_X1 #() 
INV_X1_237_ (
  .A({ S787[93] }),
  .ZN({ S103 })
);
INV_X1 #() 
INV_X1_238_ (
  .A({ S792[97] }),
  .ZN({ S104 })
);
AOI22_X1 #() 
AOI22_X1_65_ (
  .A1({ S104 }),
  .A2({ S787[97] }),
  .B1({ S103 }),
  .B2({ S792[93] }),
  .ZN({ S105 })
);
XNOR2_X1 #() 
XNOR2_X1_21_ (
  .A({ S792[116] }),
  .B({ S787[116] }),
  .ZN({ S106 })
);
XNOR2_X1 #() 
XNOR2_X1_22_ (
  .A({ S792[89] }),
  .B({ S787[89] }),
  .ZN({ S107 })
);
INV_X1 #() 
INV_X1_239_ (
  .A({ S792[59] }),
  .ZN({ S108 })
);
INV_X1 #() 
INV_X1_240_ (
  .A({ S787[61] }),
  .ZN({ S109 })
);
AOI22_X1 #() 
AOI22_X1_66_ (
  .A1({ S108 }),
  .A2({ S787[59] }),
  .B1({ S109 }),
  .B2({ S792[61] }),
  .ZN({ S110 })
);
NAND4_X1 #() 
NAND4_X1_30_ (
  .A1({ S110 }),
  .A2({ S107 }),
  .A3({ S106 }),
  .A4({ S105 }),
  .ZN({ S111 })
);
XNOR2_X1 #() 
XNOR2_X1_23_ (
  .A({ S792[106] }),
  .B({ S787[106] }),
  .ZN({ S112 })
);
XNOR2_X1 #() 
XNOR2_X1_24_ (
  .A({ S792[52] }),
  .B({ S787[52] }),
  .ZN({ S113 })
);
XNOR2_X1 #() 
XNOR2_X1_25_ (
  .A({ S792[110] }),
  .B({ S787[110] }),
  .ZN({ S114 })
);
XNOR2_X1 #() 
XNOR2_X1_26_ (
  .A({ S792[126] }),
  .B({ S787[126] }),
  .ZN({ S115 })
);
NAND4_X1 #() 
NAND4_X1_31_ (
  .A1({ S114 }),
  .A2({ S115 }),
  .A3({ S112 }),
  .A4({ S113 }),
  .ZN({ S116 })
);
NOR2_X1 #() 
NOR2_X1_44_ (
  .A1({ S116 }),
  .A2({ S111 }),
  .ZN({ S117 })
);
NAND3_X1 #() 
NAND3_X1_6_ (
  .A1({ S85 }),
  .A2({ S102 }),
  .A3({ S117 }),
  .ZN({ S118 })
);
NAND2_X1 #() 
NAND2_X1_87_ (
  .A1({ S792[78] }),
  .A2({ S787[78] }),
  .ZN({ S119 })
);
OR2_X1 #() 
OR2_X1_10_ (
  .A1({ S792[78] }),
  .A2({ S787[78] }),
  .ZN({ S120 })
);
NAND2_X1 #() 
NAND2_X1_88_ (
  .A1({ S792[6] }),
  .A2({ S787[6] }),
  .ZN({ S121 })
);
OR2_X1 #() 
OR2_X1_11_ (
  .A1({ S792[6] }),
  .A2({ S787[6] }),
  .ZN({ S122 })
);
AOI22_X1 #() 
AOI22_X1_67_ (
  .A1({ S121 }),
  .A2({ S122 }),
  .B1({ S120 }),
  .B2({ S119 }),
  .ZN({ S123 })
);
NAND2_X1 #() 
NAND2_X1_89_ (
  .A1({ S792[54] }),
  .A2({ S787[54] }),
  .ZN({ S124 })
);
OR2_X1 #() 
OR2_X1_12_ (
  .A1({ S792[54] }),
  .A2({ S787[54] }),
  .ZN({ S125 })
);
NAND2_X1 #() 
NAND2_X1_90_ (
  .A1({ S792[10] }),
  .A2({ S787[10] }),
  .ZN({ S126 })
);
OR2_X1 #() 
OR2_X1_13_ (
  .A1({ S792[10] }),
  .A2({ S787[10] }),
  .ZN({ S127 })
);
AOI22_X1 #() 
AOI22_X1_68_ (
  .A1({ S126 }),
  .A2({ S127 }),
  .B1({ S125 }),
  .B2({ S124 }),
  .ZN({ S128 })
);
INV_X1 #() 
INV_X1_241_ (
  .A({ S787[64] }),
  .ZN({ S129 })
);
NOR2_X1 #() 
NOR2_X1_45_ (
  .A1({ S129 }),
  .A2({ S792[64] }),
  .ZN({ S130 })
);
AND2_X1 #() 
AND2_X1_16_ (
  .A1({ S129 }),
  .A2({ S792[64] }),
  .ZN({ S131 })
);
INV_X1 #() 
INV_X1_242_ (
  .A({ S787[31] }),
  .ZN({ S132 })
);
INV_X1 #() 
INV_X1_243_ (
  .A({ S787[51] }),
  .ZN({ S133 })
);
OAI22_X1 #() 
OAI22_X1_42_ (
  .A1({ S792[31] }),
  .A2({ S132 }),
  .B1({ S133 }),
  .B2({ S792[51] }),
  .ZN({ S134 })
);
NOR3_X1 #() 
NOR3_X1_8_ (
  .A1({ S134 }),
  .A2({ S131 }),
  .A3({ S130 }),
  .ZN({ S135 })
);
INV_X1 #() 
INV_X1_244_ (
  .A({ S792[12] }),
  .ZN({ S136 })
);
INV_X1 #() 
INV_X1_245_ (
  .A({ S787[14] }),
  .ZN({ S137 })
);
OAI22_X1 #() 
OAI22_X1_43_ (
  .A1({ S136 }),
  .A2({ S787[12] }),
  .B1({ S137 }),
  .B2({ S792[14] }),
  .ZN({ S138 })
);
INV_X1 #() 
INV_X1_246_ (
  .A({ S787[8] }),
  .ZN({ S139 })
);
INV_X1 #() 
INV_X1_247_ (
  .A({ S792[14] }),
  .ZN({ S140 })
);
OAI22_X1 #() 
OAI22_X1_44_ (
  .A1({ S139 }),
  .A2({ S792[8] }),
  .B1({ S140 }),
  .B2({ S787[14] }),
  .ZN({ S141 })
);
NOR2_X1 #() 
NOR2_X1_46_ (
  .A1({ S138 }),
  .A2({ S141 }),
  .ZN({ S142 })
);
NAND4_X1 #() 
NAND4_X1_32_ (
  .A1({ S135 }),
  .A2({ S142 }),
  .A3({ S123 }),
  .A4({ S128 }),
  .ZN({ S143 })
);
OAI22_X1 #() 
OAI22_X1_45_ (
  .A1({ S88 }),
  .A2({ S792[117] }),
  .B1({ S99 }),
  .B2({ S787[127] }),
  .ZN({ S144 })
);
INV_X1 #() 
INV_X1_248_ (
  .A({ S787[121] }),
  .ZN({ S145 })
);
OAI22_X1 #() 
OAI22_X1_46_ (
  .A1({ S145 }),
  .A2({ S792[121] }),
  .B1({ S95 }),
  .B2({ S787[123] }),
  .ZN({ S146 })
);
NOR2_X1 #() 
NOR2_X1_47_ (
  .A1({ S144 }),
  .A2({ S146 }),
  .ZN({ S147 })
);
INV_X1 #() 
INV_X1_249_ (
  .A({ S792[119] }),
  .ZN({ S148 })
);
AOI22_X1 #() 
AOI22_X1_69_ (
  .A1({ S148 }),
  .A2({ S787[119] }),
  .B1({ S145 }),
  .B2({ S792[121] }),
  .ZN({ S149 })
);
INV_X1 #() 
INV_X1_250_ (
  .A({ S792[101] }),
  .ZN({ S150 })
);
INV_X1 #() 
INV_X1_251_ (
  .A({ S787[111] }),
  .ZN({ S151 })
);
AOI22_X1 #() 
AOI22_X1_70_ (
  .A1({ S150 }),
  .A2({ S787[101] }),
  .B1({ S151 }),
  .B2({ S792[111] }),
  .ZN({ S152 })
);
AND2_X1 #() 
AND2_X1_17_ (
  .A1({ S152 }),
  .A2({ S149 }),
  .ZN({ S153 })
);
INV_X1 #() 
INV_X1_252_ (
  .A({ S792[8] }),
  .ZN({ S154 })
);
INV_X1 #() 
INV_X1_253_ (
  .A({ S787[12] }),
  .ZN({ S155 })
);
OAI22_X1 #() 
OAI22_X1_47_ (
  .A1({ S154 }),
  .A2({ S787[8] }),
  .B1({ S155 }),
  .B2({ S792[12] }),
  .ZN({ S156 })
);
AND2_X1 #() 
AND2_X1_18_ (
  .A1({ S787[62] }),
  .A2({ S792[62] }),
  .ZN({ S157 })
);
NOR2_X1 #() 
NOR2_X1_48_ (
  .A1({ S792[62] }),
  .A2({ S787[62] }),
  .ZN({ S158 })
);
NOR2_X1 #() 
NOR2_X1_49_ (
  .A1({ S157 }),
  .A2({ S158 }),
  .ZN({ S159 })
);
NOR2_X1 #() 
NOR2_X1_50_ (
  .A1({ S159 }),
  .A2({ S156 }),
  .ZN({ S160 })
);
NAND2_X1 #() 
NAND2_X1_91_ (
  .A1({ S792[120] }),
  .A2({ S787[120] }),
  .ZN({ S161 })
);
OR2_X1 #() 
OR2_X1_14_ (
  .A1({ S792[120] }),
  .A2({ S787[120] }),
  .ZN({ S162 })
);
NAND2_X1 #() 
NAND2_X1_92_ (
  .A1({ S792[118] }),
  .A2({ S787[118] }),
  .ZN({ S163 })
);
OR2_X1 #() 
OR2_X1_15_ (
  .A1({ S792[118] }),
  .A2({ S787[118] }),
  .ZN({ S164 })
);
AOI22_X1 #() 
AOI22_X1_71_ (
  .A1({ S163 }),
  .A2({ S164 }),
  .B1({ S162 }),
  .B2({ S161 }),
  .ZN({ S165 })
);
NAND4_X1 #() 
NAND4_X1_33_ (
  .A1({ S153 }),
  .A2({ S147 }),
  .A3({ S160 }),
  .A4({ S165 }),
  .ZN({ S166 })
);
NOR2_X1 #() 
NOR2_X1_51_ (
  .A1({ S166 }),
  .A2({ S143 }),
  .ZN({ S167 })
);
INV_X1 #() 
INV_X1_254_ (
  .A({ S787[29] }),
  .ZN({ S168 })
);
INV_X1 #() 
INV_X1_255_ (
  .A({ S792[31] }),
  .ZN({ S169 })
);
OAI22_X1 #() 
OAI22_X1_48_ (
  .A1({ S168 }),
  .A2({ S792[29] }),
  .B1({ S169 }),
  .B2({ S787[31] }),
  .ZN({ S170 })
);
OAI22_X1 #() 
OAI22_X1_49_ (
  .A1({ S787[13] }),
  .A2({ S35 }),
  .B1({ S104 }),
  .B2({ S787[97] }),
  .ZN({ S171 })
);
NOR2_X1 #() 
NOR2_X1_52_ (
  .A1({ S170 }),
  .A2({ S171 }),
  .ZN({ S172 })
);
INV_X1 #() 
INV_X1_256_ (
  .A({ S792[37] }),
  .ZN({ S173 })
);
AOI22_X1 #() 
AOI22_X1_72_ (
  .A1({ S173 }),
  .A2({ S787[37] }),
  .B1({ S71 }),
  .B2({ S792[39] }),
  .ZN({ S174 })
);
INV_X1 #() 
INV_X1_257_ (
  .A({ S792[43] }),
  .ZN({ S175 })
);
INV_X1 #() 
INV_X1_258_ (
  .A({ S787[45] }),
  .ZN({ S176 })
);
AOI22_X1 #() 
AOI22_X1_73_ (
  .A1({ S175 }),
  .A2({ S787[43] }),
  .B1({ S176 }),
  .B2({ S792[45] }),
  .ZN({ S177 })
);
AND2_X1 #() 
AND2_X1_19_ (
  .A1({ S177 }),
  .A2({ S174 }),
  .ZN({ S178 })
);
XNOR2_X1 #() 
XNOR2_X1_27_ (
  .A({ S792[11] }),
  .B({ S787[11] }),
  .ZN({ S179 })
);
INV_X1 #() 
INV_X1_259_ (
  .A({ S792[87] }),
  .ZN({ S180 })
);
INV_X1 #() 
INV_X1_260_ (
  .A({ S787[99] }),
  .ZN({ S181 })
);
AOI22_X1 #() 
AOI22_X1_74_ (
  .A1({ S180 }),
  .A2({ S787[87] }),
  .B1({ S181 }),
  .B2({ S792[99] }),
  .ZN({ S182 })
);
AND2_X1 #() 
AND2_X1_20_ (
  .A1({ S179 }),
  .A2({ S182 }),
  .ZN({ S183 })
);
INV_X1 #() 
INV_X1_261_ (
  .A({ S792[9] }),
  .ZN({ S184 })
);
INV_X1 #() 
INV_X1_262_ (
  .A({ S792[93] }),
  .ZN({ S185 })
);
AOI22_X1 #() 
AOI22_X1_75_ (
  .A1({ S787[9] }),
  .A2({ S184 }),
  .B1({ S185 }),
  .B2({ S787[93] }),
  .ZN({ S186 })
);
INV_X1 #() 
INV_X1_263_ (
  .A({ S792[17] }),
  .ZN({ S187 })
);
INV_X1 #() 
INV_X1_264_ (
  .A({ S787[19] }),
  .ZN({ S188 })
);
AOI22_X1 #() 
AOI22_X1_76_ (
  .A1({ S187 }),
  .A2({ S787[17] }),
  .B1({ S188 }),
  .B2({ S792[19] }),
  .ZN({ S189 })
);
AND2_X1 #() 
AND2_X1_21_ (
  .A1({ S189 }),
  .A2({ S186 }),
  .ZN({ S190 })
);
NAND4_X1 #() 
NAND4_X1_34_ (
  .A1({ S190 }),
  .A2({ S183 }),
  .A3({ S178 }),
  .A4({ S172 }),
  .ZN({ S191 })
);
INV_X1 #() 
INV_X1_265_ (
  .A({ S787[77] }),
  .ZN({ S192 })
);
AND2_X1 #() 
AND2_X1_22_ (
  .A1({ S192 }),
  .A2({ S792[77] }),
  .ZN({ S193 })
);
NOR2_X1 #() 
NOR2_X1_53_ (
  .A1({ S192 }),
  .A2({ S792[77] }),
  .ZN({ S194 })
);
OAI22_X1 #() 
OAI22_X1_50_ (
  .A1({ S77 }),
  .A2({ S792[35] }),
  .B1({ S173 }),
  .B2({ S787[37] }),
  .ZN({ S195 })
);
NOR3_X1 #() 
NOR3_X1_9_ (
  .A1({ S195 }),
  .A2({ S193 }),
  .A3({ S194 }),
  .ZN({ S196 })
);
INV_X1 #() 
INV_X1_266_ (
  .A({ S787[3] }),
  .ZN({ S197 })
);
OAI22_X1 #() 
OAI22_X1_51_ (
  .A1({ S792[1] }),
  .A2({ S28 }),
  .B1({ S197 }),
  .B2({ S792[3] }),
  .ZN({ S198 })
);
OAI22_X1 #() 
OAI22_X1_52_ (
  .A1({ S9 }),
  .A2({ S792[57] }),
  .B1({ S108 }),
  .B2({ S787[59] }),
  .ZN({ S199 })
);
NOR2_X1 #() 
NOR2_X1_54_ (
  .A1({ S198 }),
  .A2({ S199 }),
  .ZN({ S200 })
);
INV_X1 #() 
INV_X1_267_ (
  .A({ S792[47] }),
  .ZN({ S201 })
);
OAI22_X1 #() 
OAI22_X1_53_ (
  .A1({ S787[17] }),
  .A2({ S187 }),
  .B1({ S201 }),
  .B2({ S787[47] }),
  .ZN({ S202 })
);
OAI22_X1 #() 
OAI22_X1_54_ (
  .A1({ S151 }),
  .A2({ S792[111] }),
  .B1({ S87 }),
  .B2({ S787[113] }),
  .ZN({ S203 })
);
NOR2_X1 #() 
NOR2_X1_55_ (
  .A1({ S202 }),
  .A2({ S203 }),
  .ZN({ S204 })
);
INV_X1 #() 
INV_X1_268_ (
  .A({ S792[85] }),
  .ZN({ S205 })
);
OAI22_X1 #() 
OAI22_X1_55_ (
  .A1({ S33 }),
  .A2({ S792[81] }),
  .B1({ S205 }),
  .B2({ S787[85] }),
  .ZN({ S206 })
);
INV_X1 #() 
INV_X1_269_ (
  .A({ S792[23] }),
  .ZN({ S207 })
);
INV_X1 #() 
INV_X1_270_ (
  .A({ S792[27] }),
  .ZN({ S208 })
);
OAI22_X1 #() 
OAI22_X1_56_ (
  .A1({ S787[23] }),
  .A2({ S207 }),
  .B1({ S208 }),
  .B2({ S787[27] }),
  .ZN({ S209 })
);
NOR2_X1 #() 
NOR2_X1_56_ (
  .A1({ S206 }),
  .A2({ S209 }),
  .ZN({ S210 })
);
NAND4_X1 #() 
NAND4_X1_35_ (
  .A1({ S196 }),
  .A2({ S200 }),
  .A3({ S204 }),
  .A4({ S210 }),
  .ZN({ S211 })
);
NOR2_X1 #() 
NOR2_X1_57_ (
  .A1({ S191 }),
  .A2({ S211 }),
  .ZN({ S212 })
);
INV_X1 #() 
INV_X1_271_ (
  .A({ S787[103] }),
  .ZN({ S213 })
);
INV_X1 #() 
INV_X1_272_ (
  .A({ S792[105] }),
  .ZN({ S214 })
);
OAI22_X1 #() 
OAI22_X1_57_ (
  .A1({ S213 }),
  .A2({ S792[103] }),
  .B1({ S214 }),
  .B2({ S787[105] }),
  .ZN({ S215 })
);
OAI22_X1 #() 
OAI22_X1_58_ (
  .A1({ S78 }),
  .A2({ S792[41] }),
  .B1({ S175 }),
  .B2({ S787[43] }),
  .ZN({ S216 })
);
NOR2_X1 #() 
NOR2_X1_58_ (
  .A1({ S215 }),
  .A2({ S216 }),
  .ZN({ S217 })
);
INV_X1 #() 
INV_X1_273_ (
  .A({ S787[53] }),
  .ZN({ S218 })
);
OAI22_X1 #() 
OAI22_X1_59_ (
  .A1({ S218 }),
  .A2({ S792[53] }),
  .B1({ S58 }),
  .B2({ S787[55] }),
  .ZN({ S219 })
);
INV_X1 #() 
INV_X1_274_ (
  .A({ S787[83] }),
  .ZN({ S220 })
);
AND2_X1 #() 
AND2_X1_23_ (
  .A1({ S220 }),
  .A2({ S792[83] }),
  .ZN({ S221 })
);
NOR2_X1 #() 
NOR2_X1_59_ (
  .A1({ S220 }),
  .A2({ S792[83] }),
  .ZN({ S222 })
);
NOR3_X1 #() 
NOR3_X1_10_ (
  .A1({ S219 }),
  .A2({ S221 }),
  .A3({ S222 }),
  .ZN({ S223 })
);
OAI22_X1 #() 
OAI22_X1_60_ (
  .A1({ S72 }),
  .A2({ S792[5] }),
  .B1({ S184 }),
  .B2({ S787[9] }),
  .ZN({ S224 })
);
XOR2_X1 #() 
XOR2_X1_2_ (
  .A({ S792[7] }),
  .B({ S787[7] }),
  .Z({ S225 })
);
NOR2_X1 #() 
NOR2_X1_60_ (
  .A1({ S225 }),
  .A2({ S224 }),
  .ZN({ S226 })
);
INV_X1 #() 
INV_X1_275_ (
  .A({ S787[49] }),
  .ZN({ S227 })
);
NAND2_X1 #() 
NAND2_X1_93_ (
  .A1({ S227 }),
  .A2({ S792[49] }),
  .ZN({ S228 })
);
NAND2_X1 #() 
NAND2_X1_94_ (
  .A1({ S201 }),
  .A2({ S787[47] }),
  .ZN({ S229 })
);
INV_X1 #() 
INV_X1_276_ (
  .A({ S787[25] }),
  .ZN({ S230 })
);
NAND2_X1 #() 
NAND2_X1_95_ (
  .A1({ S230 }),
  .A2({ S792[25] }),
  .ZN({ S231 })
);
NAND2_X1 #() 
NAND2_X1_96_ (
  .A1({ S207 }),
  .A2({ S787[23] }),
  .ZN({ S232 })
);
AND4_X1 #() 
AND4_X1_13_ (
  .A1({ S228 }),
  .A2({ S231 }),
  .A3({ S232 }),
  .A4({ S229 }),
  .ZN({ S233 })
);
NAND4_X1 #() 
NAND4_X1_36_ (
  .A1({ S226 }),
  .A2({ S223 }),
  .A3({ S217 }),
  .A4({ S233 }),
  .ZN({ S234 })
);
INV_X1 #() 
INV_X1_277_ (
  .A({ S792[29] }),
  .ZN({ S235 })
);
OAI22_X1 #() 
OAI22_X1_61_ (
  .A1({ S235 }),
  .A2({ S787[29] }),
  .B1({ S176 }),
  .B2({ S792[45] }),
  .ZN({ S236 })
);
OAI22_X1 #() 
OAI22_X1_62_ (
  .A1({ S792[21] }),
  .A2({ S36 }),
  .B1({ S227 }),
  .B2({ S792[49] }),
  .ZN({ S237 })
);
NOR2_X1 #() 
NOR2_X1_61_ (
  .A1({ S236 }),
  .A2({ S237 }),
  .ZN({ S238 })
);
INV_X1 #() 
INV_X1_278_ (
  .A({ S792[3] }),
  .ZN({ S239 })
);
OAI22_X1 #() 
OAI22_X1_63_ (
  .A1({ S239 }),
  .A2({ S787[3] }),
  .B1({ S188 }),
  .B2({ S792[19] }),
  .ZN({ S240 })
);
INV_X1 #() 
INV_X1_279_ (
  .A({ S787[27] }),
  .ZN({ S241 })
);
INV_X1 #() 
INV_X1_280_ (
  .A({ S787[33] }),
  .ZN({ S242 })
);
OAI22_X1 #() 
OAI22_X1_64_ (
  .A1({ S792[27] }),
  .A2({ S241 }),
  .B1({ S242 }),
  .B2({ S792[33] }),
  .ZN({ S243 })
);
NOR2_X1 #() 
NOR2_X1_62_ (
  .A1({ S240 }),
  .A2({ S243 }),
  .ZN({ S244 })
);
OAI22_X1 #() 
OAI22_X1_65_ (
  .A1({ S11 }),
  .A2({ S792[73] }),
  .B1({ S13 }),
  .B2({ S787[79] }),
  .ZN({ S245 })
);
INV_X1 #() 
INV_X1_281_ (
  .A({ S787[75] }),
  .ZN({ S246 })
);
AND2_X1 #() 
AND2_X1_24_ (
  .A1({ S246 }),
  .A2({ S792[75] }),
  .ZN({ S247 })
);
NOR2_X1 #() 
NOR2_X1_63_ (
  .A1({ S246 }),
  .A2({ S792[75] }),
  .ZN({ S248 })
);
NOR3_X1 #() 
NOR3_X1_11_ (
  .A1({ S245 }),
  .A2({ S247 }),
  .A3({ S248 }),
  .ZN({ S249 })
);
INV_X1 #() 
INV_X1_282_ (
  .A({ S792[33] }),
  .ZN({ S250 })
);
OAI22_X1 #() 
OAI22_X1_66_ (
  .A1({ S230 }),
  .A2({ S792[25] }),
  .B1({ S250 }),
  .B2({ S787[33] }),
  .ZN({ S251 })
);
INV_X1 #() 
INV_X1_283_ (
  .A({ S792[51] }),
  .ZN({ S252 })
);
INV_X1 #() 
INV_X1_284_ (
  .A({ S792[53] }),
  .ZN({ S253 })
);
OAI22_X1 #() 
OAI22_X1_67_ (
  .A1({ S787[51] }),
  .A2({ S252 }),
  .B1({ S253 }),
  .B2({ S787[53] }),
  .ZN({ S254 })
);
NOR2_X1 #() 
NOR2_X1_64_ (
  .A1({ S251 }),
  .A2({ S254 }),
  .ZN({ S255 })
);
NAND4_X1 #() 
NAND4_X1_37_ (
  .A1({ S249 }),
  .A2({ S255 }),
  .A3({ S238 }),
  .A4({ S244 }),
  .ZN({ S256 })
);
NOR2_X1 #() 
NOR2_X1_65_ (
  .A1({ S234 }),
  .A2({ S256 }),
  .ZN({ S257 })
);
NAND2_X1 #() 
NAND2_X1_97_ (
  .A1({ S792[28] }),
  .A2({ S787[28] }),
  .ZN({ S258 })
);
OR2_X1 #() 
OR2_X1_16_ (
  .A1({ S792[28] }),
  .A2({ S787[28] }),
  .ZN({ S259 })
);
NAND2_X1 #() 
NAND2_X1_98_ (
  .A1({ S792[26] }),
  .A2({ S787[26] }),
  .ZN({ S260 })
);
OR2_X1 #() 
OR2_X1_17_ (
  .A1({ S792[26] }),
  .A2({ S787[26] }),
  .ZN({ S261 })
);
AOI22_X1 #() 
AOI22_X1_77_ (
  .A1({ S260 }),
  .A2({ S261 }),
  .B1({ S259 }),
  .B2({ S258 }),
  .ZN({ S262 })
);
NAND2_X1 #() 
NAND2_X1_99_ (
  .A1({ S792[108] }),
  .A2({ S787[108] }),
  .ZN({ S263 })
);
OR2_X1 #() 
OR2_X1_18_ (
  .A1({ S792[108] }),
  .A2({ S787[108] }),
  .ZN({ S264 })
);
NAND2_X1 #() 
NAND2_X1_100_ (
  .A1({ S792[102] }),
  .A2({ S787[102] }),
  .ZN({ S265 })
);
OR2_X1 #() 
OR2_X1_19_ (
  .A1({ S792[102] }),
  .A2({ S787[102] }),
  .ZN({ S266 })
);
AOI22_X1 #() 
AOI22_X1_78_ (
  .A1({ S265 }),
  .A2({ S266 }),
  .B1({ S264 }),
  .B2({ S263 }),
  .ZN({ S267 })
);
INV_X1 #() 
INV_X1_285_ (
  .A({ S792[103] }),
  .ZN({ S268 })
);
INV_X1 #() 
INV_X1_286_ (
  .A({ S792[109] }),
  .ZN({ S269 })
);
OAI22_X1 #() 
OAI22_X1_68_ (
  .A1({ S787[103] }),
  .A2({ S268 }),
  .B1({ S269 }),
  .B2({ S787[109] }),
  .ZN({ S270 })
);
INV_X1 #() 
INV_X1_287_ (
  .A({ S787[105] }),
  .ZN({ S271 })
);
INV_X1 #() 
INV_X1_288_ (
  .A({ S787[109] }),
  .ZN({ S272 })
);
OAI22_X1 #() 
OAI22_X1_69_ (
  .A1({ S792[105] }),
  .A2({ S271 }),
  .B1({ S272 }),
  .B2({ S792[109] }),
  .ZN({ S273 })
);
NOR2_X1 #() 
NOR2_X1_66_ (
  .A1({ S270 }),
  .A2({ S273 }),
  .ZN({ S274 })
);
NAND2_X1 #() 
NAND2_X1_101_ (
  .A1({ S792[112] }),
  .A2({ S787[112] }),
  .ZN({ S275 })
);
OR2_X1 #() 
OR2_X1_20_ (
  .A1({ S792[112] }),
  .A2({ S787[112] }),
  .ZN({ S276 })
);
NAND2_X1 #() 
NAND2_X1_102_ (
  .A1({ S792[38] }),
  .A2({ S787[38] }),
  .ZN({ S277 })
);
OR2_X1 #() 
OR2_X1_21_ (
  .A1({ S792[38] }),
  .A2({ S787[38] }),
  .ZN({ S278 })
);
AOI22_X1 #() 
AOI22_X1_79_ (
  .A1({ S277 }),
  .A2({ S278 }),
  .B1({ S276 }),
  .B2({ S275 }),
  .ZN({ S279 })
);
NAND4_X1 #() 
NAND4_X1_38_ (
  .A1({ S274 }),
  .A2({ S279 }),
  .A3({ S262 }),
  .A4({ S267 }),
  .ZN({ S280 })
);
INV_X1 #() 
INV_X1_289_ (
  .A({ S792[67] }),
  .ZN({ S281 })
);
OAI22_X1 #() 
OAI22_X1_70_ (
  .A1({ S24 }),
  .A2({ S792[65] }),
  .B1({ S281 }),
  .B2({ S787[67] }),
  .ZN({ S282 })
);
INV_X1 #() 
INV_X1_290_ (
  .A({ S787[67] }),
  .ZN({ S283 })
);
OAI22_X1 #() 
OAI22_X1_71_ (
  .A1({ S283 }),
  .A2({ S792[67] }),
  .B1({ S32 }),
  .B2({ S787[69] }),
  .ZN({ S284 })
);
NOR2_X1 #() 
NOR2_X1_67_ (
  .A1({ S282 }),
  .A2({ S284 }),
  .ZN({ S285 })
);
OAI22_X1 #() 
OAI22_X1_72_ (
  .A1({ S181 }),
  .A2({ S792[99] }),
  .B1({ S150 }),
  .B2({ S787[101] }),
  .ZN({ S286 })
);
INV_X1 #() 
INV_X1_291_ (
  .A({ S787[95] }),
  .ZN({ S287 })
);
AND2_X1 #() 
AND2_X1_25_ (
  .A1({ S287 }),
  .A2({ S792[95] }),
  .ZN({ S288 })
);
NOR2_X1 #() 
NOR2_X1_68_ (
  .A1({ S287 }),
  .A2({ S792[95] }),
  .ZN({ S289 })
);
NOR3_X1 #() 
NOR3_X1_12_ (
  .A1({ S286 }),
  .A2({ S288 }),
  .A3({ S289 }),
  .ZN({ S290 })
);
NAND2_X1 #() 
NAND2_X1_103_ (
  .A1({ S792[114] }),
  .A2({ S787[114] }),
  .ZN({ S291 })
);
OR2_X1 #() 
OR2_X1_22_ (
  .A1({ S792[114] }),
  .A2({ S787[114] }),
  .ZN({ S292 })
);
NAND2_X1 #() 
NAND2_X1_104_ (
  .A1({ S792[104] }),
  .A2({ S787[104] }),
  .ZN({ S293 })
);
OR2_X1 #() 
OR2_X1_23_ (
  .A1({ S792[104] }),
  .A2({ S787[104] }),
  .ZN({ S294 })
);
AOI22_X1 #() 
AOI22_X1_80_ (
  .A1({ S293 }),
  .A2({ S294 }),
  .B1({ S292 }),
  .B2({ S291 }),
  .ZN({ S295 })
);
INV_X1 #() 
INV_X1_292_ (
  .A({ S787[85] }),
  .ZN({ S296 })
);
OAI22_X1 #() 
OAI22_X1_73_ (
  .A1({ S296 }),
  .A2({ S792[85] }),
  .B1({ S180 }),
  .B2({ S787[87] }),
  .ZN({ S297 })
);
XOR2_X1 #() 
XOR2_X1_3_ (
  .A({ S792[91] }),
  .B({ S787[91] }),
  .Z({ S298 })
);
NOR2_X1 #() 
NOR2_X1_69_ (
  .A1({ S298 }),
  .A2({ S297 }),
  .ZN({ S299 })
);
NAND4_X1 #() 
NAND4_X1_39_ (
  .A1({ S299 }),
  .A2({ S290 }),
  .A3({ S295 }),
  .A4({ S285 }),
  .ZN({ S300 })
);
NOR2_X1 #() 
NOR2_X1_70_ (
  .A1({ S300 }),
  .A2({ S280 }),
  .ZN({ S301 })
);
NAND4_X1 #() 
NAND4_X1_40_ (
  .A1({ S212 }),
  .A2({ S257 }),
  .A3({ S167 }),
  .A4({ S301 }),
  .ZN({ S302 })
);
NOR3_X1 #() 
NOR3_X1_13_ (
  .A1({ S302 }),
  .A2({ S70 }),
  .A3({ S118 }),
  .ZN({ S786 })
);
BUF_X1 #() 
BUF_X1_1_ (
  .A({ S786 }),
  .Z({ d128 })
);
BUF_X1 #() 
BUF_X1_2_ (
  .A({ S787[0] }),
  .Z({ decrypted128[0] })
);
BUF_X1 #() 
BUF_X1_3_ (
  .A({ S787[1] }),
  .Z({ decrypted128[1] })
);
BUF_X1 #() 
BUF_X1_4_ (
  .A({ S787[10] }),
  .Z({ decrypted128[10] })
);
BUF_X1 #() 
BUF_X1_5_ (
  .A({ S787[100] }),
  .Z({ decrypted128[100] })
);
BUF_X1 #() 
BUF_X1_6_ (
  .A({ S787[101] }),
  .Z({ decrypted128[101] })
);
BUF_X1 #() 
BUF_X1_7_ (
  .A({ S787[102] }),
  .Z({ decrypted128[102] })
);
BUF_X1 #() 
BUF_X1_8_ (
  .A({ S787[103] }),
  .Z({ decrypted128[103] })
);
BUF_X1 #() 
BUF_X1_9_ (
  .A({ S787[104] }),
  .Z({ decrypted128[104] })
);
BUF_X1 #() 
BUF_X1_10_ (
  .A({ S787[105] }),
  .Z({ decrypted128[105] })
);
BUF_X1 #() 
BUF_X1_11_ (
  .A({ S787[106] }),
  .Z({ decrypted128[106] })
);
BUF_X1 #() 
BUF_X1_12_ (
  .A({ S787[107] }),
  .Z({ decrypted128[107] })
);
BUF_X1 #() 
BUF_X1_13_ (
  .A({ S787[108] }),
  .Z({ decrypted128[108] })
);
BUF_X1 #() 
BUF_X1_14_ (
  .A({ S787[109] }),
  .Z({ decrypted128[109] })
);
BUF_X1 #() 
BUF_X1_15_ (
  .A({ S787[11] }),
  .Z({ decrypted128[11] })
);
BUF_X1 #() 
BUF_X1_16_ (
  .A({ S787[110] }),
  .Z({ decrypted128[110] })
);
BUF_X1 #() 
BUF_X1_17_ (
  .A({ S787[111] }),
  .Z({ decrypted128[111] })
);
BUF_X1 #() 
BUF_X1_18_ (
  .A({ S787[112] }),
  .Z({ decrypted128[112] })
);
BUF_X1 #() 
BUF_X1_19_ (
  .A({ S787[113] }),
  .Z({ decrypted128[113] })
);
BUF_X1 #() 
BUF_X1_20_ (
  .A({ S787[114] }),
  .Z({ decrypted128[114] })
);
BUF_X1 #() 
BUF_X1_21_ (
  .A({ S787[115] }),
  .Z({ decrypted128[115] })
);
BUF_X1 #() 
BUF_X1_22_ (
  .A({ S787[116] }),
  .Z({ decrypted128[116] })
);
BUF_X1 #() 
BUF_X1_23_ (
  .A({ S787[117] }),
  .Z({ decrypted128[117] })
);
BUF_X1 #() 
BUF_X1_24_ (
  .A({ S787[118] }),
  .Z({ decrypted128[118] })
);
BUF_X1 #() 
BUF_X1_25_ (
  .A({ S787[119] }),
  .Z({ decrypted128[119] })
);
BUF_X1 #() 
BUF_X1_26_ (
  .A({ S787[12] }),
  .Z({ decrypted128[12] })
);
BUF_X1 #() 
BUF_X1_27_ (
  .A({ S787[120] }),
  .Z({ decrypted128[120] })
);
BUF_X1 #() 
BUF_X1_28_ (
  .A({ S787[121] }),
  .Z({ decrypted128[121] })
);
BUF_X1 #() 
BUF_X1_29_ (
  .A({ S787[122] }),
  .Z({ decrypted128[122] })
);
BUF_X1 #() 
BUF_X1_30_ (
  .A({ S787[123] }),
  .Z({ decrypted128[123] })
);
BUF_X1 #() 
BUF_X1_31_ (
  .A({ S787[124] }),
  .Z({ decrypted128[124] })
);
BUF_X1 #() 
BUF_X1_32_ (
  .A({ S787[125] }),
  .Z({ decrypted128[125] })
);
BUF_X1 #() 
BUF_X1_33_ (
  .A({ S787[126] }),
  .Z({ decrypted128[126] })
);
BUF_X1 #() 
BUF_X1_34_ (
  .A({ S787[127] }),
  .Z({ decrypted128[127] })
);
BUF_X1 #() 
BUF_X1_35_ (
  .A({ S787[13] }),
  .Z({ decrypted128[13] })
);
BUF_X1 #() 
BUF_X1_36_ (
  .A({ S787[14] }),
  .Z({ decrypted128[14] })
);
BUF_X1 #() 
BUF_X1_37_ (
  .A({ S787[15] }),
  .Z({ decrypted128[15] })
);
BUF_X1 #() 
BUF_X1_38_ (
  .A({ S787[16] }),
  .Z({ decrypted128[16] })
);
BUF_X1 #() 
BUF_X1_39_ (
  .A({ S787[17] }),
  .Z({ decrypted128[17] })
);
BUF_X1 #() 
BUF_X1_40_ (
  .A({ S787[18] }),
  .Z({ decrypted128[18] })
);
BUF_X1 #() 
BUF_X1_41_ (
  .A({ S787[19] }),
  .Z({ decrypted128[19] })
);
BUF_X1 #() 
BUF_X1_42_ (
  .A({ S787[2] }),
  .Z({ decrypted128[2] })
);
BUF_X1 #() 
BUF_X1_43_ (
  .A({ S787[20] }),
  .Z({ decrypted128[20] })
);
BUF_X1 #() 
BUF_X1_44_ (
  .A({ S787[21] }),
  .Z({ decrypted128[21] })
);
BUF_X1 #() 
BUF_X1_45_ (
  .A({ S787[22] }),
  .Z({ decrypted128[22] })
);
BUF_X1 #() 
BUF_X1_46_ (
  .A({ S787[23] }),
  .Z({ decrypted128[23] })
);
BUF_X1 #() 
BUF_X1_47_ (
  .A({ S787[24] }),
  .Z({ decrypted128[24] })
);
BUF_X1 #() 
BUF_X1_48_ (
  .A({ S787[25] }),
  .Z({ decrypted128[25] })
);
BUF_X1 #() 
BUF_X1_49_ (
  .A({ S787[26] }),
  .Z({ decrypted128[26] })
);
BUF_X1 #() 
BUF_X1_50_ (
  .A({ S787[27] }),
  .Z({ decrypted128[27] })
);
BUF_X1 #() 
BUF_X1_51_ (
  .A({ S787[28] }),
  .Z({ decrypted128[28] })
);
BUF_X1 #() 
BUF_X1_52_ (
  .A({ S787[29] }),
  .Z({ decrypted128[29] })
);
BUF_X1 #() 
BUF_X1_53_ (
  .A({ S787[3] }),
  .Z({ decrypted128[3] })
);
BUF_X1 #() 
BUF_X1_54_ (
  .A({ S787[30] }),
  .Z({ decrypted128[30] })
);
BUF_X1 #() 
BUF_X1_55_ (
  .A({ S787[31] }),
  .Z({ decrypted128[31] })
);
BUF_X1 #() 
BUF_X1_56_ (
  .A({ S787[32] }),
  .Z({ decrypted128[32] })
);
BUF_X1 #() 
BUF_X1_57_ (
  .A({ S787[33] }),
  .Z({ decrypted128[33] })
);
BUF_X1 #() 
BUF_X1_58_ (
  .A({ S787[34] }),
  .Z({ decrypted128[34] })
);
BUF_X1 #() 
BUF_X1_59_ (
  .A({ S787[35] }),
  .Z({ decrypted128[35] })
);
BUF_X1 #() 
BUF_X1_60_ (
  .A({ S787[36] }),
  .Z({ decrypted128[36] })
);
BUF_X1 #() 
BUF_X1_61_ (
  .A({ S787[37] }),
  .Z({ decrypted128[37] })
);
BUF_X1 #() 
BUF_X1_62_ (
  .A({ S787[38] }),
  .Z({ decrypted128[38] })
);
BUF_X1 #() 
BUF_X1_63_ (
  .A({ S787[39] }),
  .Z({ decrypted128[39] })
);
BUF_X1 #() 
BUF_X1_64_ (
  .A({ S787[4] }),
  .Z({ decrypted128[4] })
);
BUF_X1 #() 
BUF_X1_65_ (
  .A({ S787[40] }),
  .Z({ decrypted128[40] })
);
BUF_X1 #() 
BUF_X1_66_ (
  .A({ S787[41] }),
  .Z({ decrypted128[41] })
);
BUF_X1 #() 
BUF_X1_67_ (
  .A({ S787[42] }),
  .Z({ decrypted128[42] })
);
BUF_X1 #() 
BUF_X1_68_ (
  .A({ S787[43] }),
  .Z({ decrypted128[43] })
);
BUF_X1 #() 
BUF_X1_69_ (
  .A({ S787[44] }),
  .Z({ decrypted128[44] })
);
BUF_X1 #() 
BUF_X1_70_ (
  .A({ S787[45] }),
  .Z({ decrypted128[45] })
);
BUF_X1 #() 
BUF_X1_71_ (
  .A({ S787[46] }),
  .Z({ decrypted128[46] })
);
BUF_X1 #() 
BUF_X1_72_ (
  .A({ S787[47] }),
  .Z({ decrypted128[47] })
);
BUF_X1 #() 
BUF_X1_73_ (
  .A({ S787[48] }),
  .Z({ decrypted128[48] })
);
BUF_X1 #() 
BUF_X1_74_ (
  .A({ S787[49] }),
  .Z({ decrypted128[49] })
);
BUF_X1 #() 
BUF_X1_75_ (
  .A({ S787[5] }),
  .Z({ decrypted128[5] })
);
BUF_X1 #() 
BUF_X1_76_ (
  .A({ S787[50] }),
  .Z({ decrypted128[50] })
);
BUF_X1 #() 
BUF_X1_77_ (
  .A({ S787[51] }),
  .Z({ decrypted128[51] })
);
BUF_X1 #() 
BUF_X1_78_ (
  .A({ S787[52] }),
  .Z({ decrypted128[52] })
);
BUF_X1 #() 
BUF_X1_79_ (
  .A({ S787[53] }),
  .Z({ decrypted128[53] })
);
BUF_X1 #() 
BUF_X1_80_ (
  .A({ S787[54] }),
  .Z({ decrypted128[54] })
);
BUF_X1 #() 
BUF_X1_81_ (
  .A({ S787[55] }),
  .Z({ decrypted128[55] })
);
BUF_X1 #() 
BUF_X1_82_ (
  .A({ S787[56] }),
  .Z({ decrypted128[56] })
);
BUF_X1 #() 
BUF_X1_83_ (
  .A({ S787[57] }),
  .Z({ decrypted128[57] })
);
BUF_X1 #() 
BUF_X1_84_ (
  .A({ S787[58] }),
  .Z({ decrypted128[58] })
);
BUF_X1 #() 
BUF_X1_85_ (
  .A({ S787[59] }),
  .Z({ decrypted128[59] })
);
BUF_X1 #() 
BUF_X1_86_ (
  .A({ S787[6] }),
  .Z({ decrypted128[6] })
);
BUF_X1 #() 
BUF_X1_87_ (
  .A({ S787[60] }),
  .Z({ decrypted128[60] })
);
BUF_X1 #() 
BUF_X1_88_ (
  .A({ S787[61] }),
  .Z({ decrypted128[61] })
);
BUF_X1 #() 
BUF_X1_89_ (
  .A({ S787[62] }),
  .Z({ decrypted128[62] })
);
BUF_X1 #() 
BUF_X1_90_ (
  .A({ S787[63] }),
  .Z({ decrypted128[63] })
);
BUF_X1 #() 
BUF_X1_91_ (
  .A({ S787[64] }),
  .Z({ decrypted128[64] })
);
BUF_X1 #() 
BUF_X1_92_ (
  .A({ S787[65] }),
  .Z({ decrypted128[65] })
);
BUF_X1 #() 
BUF_X1_93_ (
  .A({ S787[66] }),
  .Z({ decrypted128[66] })
);
BUF_X1 #() 
BUF_X1_94_ (
  .A({ S787[67] }),
  .Z({ decrypted128[67] })
);
BUF_X1 #() 
BUF_X1_95_ (
  .A({ S787[68] }),
  .Z({ decrypted128[68] })
);
BUF_X1 #() 
BUF_X1_96_ (
  .A({ S787[69] }),
  .Z({ decrypted128[69] })
);
BUF_X1 #() 
BUF_X1_97_ (
  .A({ S787[7] }),
  .Z({ decrypted128[7] })
);
BUF_X1 #() 
BUF_X1_98_ (
  .A({ S787[70] }),
  .Z({ decrypted128[70] })
);
BUF_X1 #() 
BUF_X1_99_ (
  .A({ S787[71] }),
  .Z({ decrypted128[71] })
);
BUF_X1 #() 
BUF_X1_100_ (
  .A({ S787[72] }),
  .Z({ decrypted128[72] })
);
BUF_X1 #() 
BUF_X1_101_ (
  .A({ S787[73] }),
  .Z({ decrypted128[73] })
);
BUF_X1 #() 
BUF_X1_102_ (
  .A({ S787[74] }),
  .Z({ decrypted128[74] })
);
BUF_X1 #() 
BUF_X1_103_ (
  .A({ S787[75] }),
  .Z({ decrypted128[75] })
);
BUF_X1 #() 
BUF_X1_104_ (
  .A({ S787[76] }),
  .Z({ decrypted128[76] })
);
BUF_X1 #() 
BUF_X1_105_ (
  .A({ S787[77] }),
  .Z({ decrypted128[77] })
);
BUF_X1 #() 
BUF_X1_106_ (
  .A({ S787[78] }),
  .Z({ decrypted128[78] })
);
BUF_X1 #() 
BUF_X1_107_ (
  .A({ S787[79] }),
  .Z({ decrypted128[79] })
);
BUF_X1 #() 
BUF_X1_108_ (
  .A({ S787[8] }),
  .Z({ decrypted128[8] })
);
BUF_X1 #() 
BUF_X1_109_ (
  .A({ S787[80] }),
  .Z({ decrypted128[80] })
);
BUF_X1 #() 
BUF_X1_110_ (
  .A({ S787[81] }),
  .Z({ decrypted128[81] })
);
BUF_X1 #() 
BUF_X1_111_ (
  .A({ S787[82] }),
  .Z({ decrypted128[82] })
);
BUF_X1 #() 
BUF_X1_112_ (
  .A({ S787[83] }),
  .Z({ decrypted128[83] })
);
BUF_X1 #() 
BUF_X1_113_ (
  .A({ S787[84] }),
  .Z({ decrypted128[84] })
);
BUF_X1 #() 
BUF_X1_114_ (
  .A({ S787[85] }),
  .Z({ decrypted128[85] })
);
BUF_X1 #() 
BUF_X1_115_ (
  .A({ S787[86] }),
  .Z({ decrypted128[86] })
);
BUF_X1 #() 
BUF_X1_116_ (
  .A({ S787[87] }),
  .Z({ decrypted128[87] })
);
BUF_X1 #() 
BUF_X1_117_ (
  .A({ S787[88] }),
  .Z({ decrypted128[88] })
);
BUF_X1 #() 
BUF_X1_118_ (
  .A({ S787[89] }),
  .Z({ decrypted128[89] })
);
BUF_X1 #() 
BUF_X1_119_ (
  .A({ S787[9] }),
  .Z({ decrypted128[9] })
);
BUF_X1 #() 
BUF_X1_120_ (
  .A({ S787[90] }),
  .Z({ decrypted128[90] })
);
BUF_X1 #() 
BUF_X1_121_ (
  .A({ S787[91] }),
  .Z({ decrypted128[91] })
);
BUF_X1 #() 
BUF_X1_122_ (
  .A({ S787[92] }),
  .Z({ decrypted128[92] })
);
BUF_X1 #() 
BUF_X1_123_ (
  .A({ S787[93] }),
  .Z({ decrypted128[93] })
);
BUF_X1 #() 
BUF_X1_124_ (
  .A({ S787[94] }),
  .Z({ decrypted128[94] })
);
BUF_X1 #() 
BUF_X1_125_ (
  .A({ S787[95] }),
  .Z({ decrypted128[95] })
);
BUF_X1 #() 
BUF_X1_126_ (
  .A({ S787[96] }),
  .Z({ decrypted128[96] })
);
BUF_X1 #() 
BUF_X1_127_ (
  .A({ S787[97] }),
  .Z({ decrypted128[97] })
);
BUF_X1 #() 
BUF_X1_128_ (
  .A({ S787[98] }),
  .Z({ decrypted128[98] })
);
BUF_X1 #() 
BUF_X1_129_ (
  .A({ S787[99] }),
  .Z({ decrypted128[99] })
);
BUF_X1 #() 
BUF_X1_130_ (
  .A({ S788 }),
  .Z({ e128 })
);
BUF_X1 #() 
BUF_X1_131_ (
  .A({ enable }),
  .Z({ S789 })
);
BUF_X1 #() 
BUF_X1_132_ (
  .A({ S790[0] }),
  .Z({ encrypted128[0] })
);
BUF_X1 #() 
BUF_X1_133_ (
  .A({ S790[1] }),
  .Z({ encrypted128[1] })
);
BUF_X1 #() 
BUF_X1_134_ (
  .A({ S790[10] }),
  .Z({ encrypted128[10] })
);
BUF_X1 #() 
BUF_X1_135_ (
  .A({ S790[100] }),
  .Z({ encrypted128[100] })
);
BUF_X1 #() 
BUF_X1_136_ (
  .A({ S790[101] }),
  .Z({ encrypted128[101] })
);
BUF_X1 #() 
BUF_X1_137_ (
  .A({ S790[102] }),
  .Z({ encrypted128[102] })
);
BUF_X1 #() 
BUF_X1_138_ (
  .A({ S790[103] }),
  .Z({ encrypted128[103] })
);
BUF_X1 #() 
BUF_X1_139_ (
  .A({ S790[104] }),
  .Z({ encrypted128[104] })
);
BUF_X1 #() 
BUF_X1_140_ (
  .A({ S790[105] }),
  .Z({ encrypted128[105] })
);
BUF_X1 #() 
BUF_X1_141_ (
  .A({ S790[106] }),
  .Z({ encrypted128[106] })
);
BUF_X1 #() 
BUF_X1_142_ (
  .A({ S790[107] }),
  .Z({ encrypted128[107] })
);
BUF_X1 #() 
BUF_X1_143_ (
  .A({ S790[108] }),
  .Z({ encrypted128[108] })
);
BUF_X1 #() 
BUF_X1_144_ (
  .A({ S790[109] }),
  .Z({ encrypted128[109] })
);
BUF_X1 #() 
BUF_X1_145_ (
  .A({ S790[11] }),
  .Z({ encrypted128[11] })
);
BUF_X1 #() 
BUF_X1_146_ (
  .A({ S790[110] }),
  .Z({ encrypted128[110] })
);
BUF_X1 #() 
BUF_X1_147_ (
  .A({ S790[111] }),
  .Z({ encrypted128[111] })
);
BUF_X1 #() 
BUF_X1_148_ (
  .A({ S790[112] }),
  .Z({ encrypted128[112] })
);
BUF_X1 #() 
BUF_X1_149_ (
  .A({ S790[113] }),
  .Z({ encrypted128[113] })
);
BUF_X1 #() 
BUF_X1_150_ (
  .A({ S790[114] }),
  .Z({ encrypted128[114] })
);
BUF_X1 #() 
BUF_X1_151_ (
  .A({ S790[115] }),
  .Z({ encrypted128[115] })
);
BUF_X1 #() 
BUF_X1_152_ (
  .A({ S790[116] }),
  .Z({ encrypted128[116] })
);
BUF_X1 #() 
BUF_X1_153_ (
  .A({ S790[117] }),
  .Z({ encrypted128[117] })
);
BUF_X1 #() 
BUF_X1_154_ (
  .A({ S790[118] }),
  .Z({ encrypted128[118] })
);
BUF_X1 #() 
BUF_X1_155_ (
  .A({ S790[119] }),
  .Z({ encrypted128[119] })
);
BUF_X1 #() 
BUF_X1_156_ (
  .A({ S790[12] }),
  .Z({ encrypted128[12] })
);
BUF_X1 #() 
BUF_X1_157_ (
  .A({ S790[120] }),
  .Z({ encrypted128[120] })
);
BUF_X1 #() 
BUF_X1_158_ (
  .A({ S790[121] }),
  .Z({ encrypted128[121] })
);
BUF_X1 #() 
BUF_X1_159_ (
  .A({ S790[122] }),
  .Z({ encrypted128[122] })
);
BUF_X1 #() 
BUF_X1_160_ (
  .A({ S790[123] }),
  .Z({ encrypted128[123] })
);
BUF_X1 #() 
BUF_X1_161_ (
  .A({ S790[124] }),
  .Z({ encrypted128[124] })
);
BUF_X1 #() 
BUF_X1_162_ (
  .A({ S790[125] }),
  .Z({ encrypted128[125] })
);
BUF_X1 #() 
BUF_X1_163_ (
  .A({ S790[126] }),
  .Z({ encrypted128[126] })
);
BUF_X1 #() 
BUF_X1_164_ (
  .A({ S790[127] }),
  .Z({ encrypted128[127] })
);
BUF_X1 #() 
BUF_X1_165_ (
  .A({ S790[13] }),
  .Z({ encrypted128[13] })
);
BUF_X1 #() 
BUF_X1_166_ (
  .A({ S790[14] }),
  .Z({ encrypted128[14] })
);
BUF_X1 #() 
BUF_X1_167_ (
  .A({ S790[15] }),
  .Z({ encrypted128[15] })
);
BUF_X1 #() 
BUF_X1_168_ (
  .A({ S790[16] }),
  .Z({ encrypted128[16] })
);
BUF_X1 #() 
BUF_X1_169_ (
  .A({ S790[17] }),
  .Z({ encrypted128[17] })
);
BUF_X1 #() 
BUF_X1_170_ (
  .A({ S790[18] }),
  .Z({ encrypted128[18] })
);
BUF_X1 #() 
BUF_X1_171_ (
  .A({ S790[19] }),
  .Z({ encrypted128[19] })
);
BUF_X1 #() 
BUF_X1_172_ (
  .A({ S790[2] }),
  .Z({ encrypted128[2] })
);
BUF_X1 #() 
BUF_X1_173_ (
  .A({ S790[20] }),
  .Z({ encrypted128[20] })
);
BUF_X1 #() 
BUF_X1_174_ (
  .A({ S790[21] }),
  .Z({ encrypted128[21] })
);
BUF_X1 #() 
BUF_X1_175_ (
  .A({ S790[22] }),
  .Z({ encrypted128[22] })
);
BUF_X1 #() 
BUF_X1_176_ (
  .A({ S790[23] }),
  .Z({ encrypted128[23] })
);
BUF_X1 #() 
BUF_X1_177_ (
  .A({ S790[24] }),
  .Z({ encrypted128[24] })
);
BUF_X1 #() 
BUF_X1_178_ (
  .A({ S790[25] }),
  .Z({ encrypted128[25] })
);
BUF_X1 #() 
BUF_X1_179_ (
  .A({ S790[26] }),
  .Z({ encrypted128[26] })
);
BUF_X1 #() 
BUF_X1_180_ (
  .A({ S790[27] }),
  .Z({ encrypted128[27] })
);
BUF_X1 #() 
BUF_X1_181_ (
  .A({ S790[28] }),
  .Z({ encrypted128[28] })
);
BUF_X1 #() 
BUF_X1_182_ (
  .A({ S790[29] }),
  .Z({ encrypted128[29] })
);
BUF_X1 #() 
BUF_X1_183_ (
  .A({ S790[3] }),
  .Z({ encrypted128[3] })
);
BUF_X1 #() 
BUF_X1_184_ (
  .A({ S790[30] }),
  .Z({ encrypted128[30] })
);
BUF_X1 #() 
BUF_X1_185_ (
  .A({ S790[31] }),
  .Z({ encrypted128[31] })
);
BUF_X1 #() 
BUF_X1_186_ (
  .A({ S790[32] }),
  .Z({ encrypted128[32] })
);
BUF_X1 #() 
BUF_X1_187_ (
  .A({ S790[33] }),
  .Z({ encrypted128[33] })
);
BUF_X1 #() 
BUF_X1_188_ (
  .A({ S790[34] }),
  .Z({ encrypted128[34] })
);
BUF_X1 #() 
BUF_X1_189_ (
  .A({ S790[35] }),
  .Z({ encrypted128[35] })
);
BUF_X1 #() 
BUF_X1_190_ (
  .A({ S790[36] }),
  .Z({ encrypted128[36] })
);
BUF_X1 #() 
BUF_X1_191_ (
  .A({ S790[37] }),
  .Z({ encrypted128[37] })
);
BUF_X1 #() 
BUF_X1_192_ (
  .A({ S790[38] }),
  .Z({ encrypted128[38] })
);
BUF_X1 #() 
BUF_X1_193_ (
  .A({ S790[39] }),
  .Z({ encrypted128[39] })
);
BUF_X1 #() 
BUF_X1_194_ (
  .A({ S790[4] }),
  .Z({ encrypted128[4] })
);
BUF_X1 #() 
BUF_X1_195_ (
  .A({ S790[40] }),
  .Z({ encrypted128[40] })
);
BUF_X1 #() 
BUF_X1_196_ (
  .A({ S790[41] }),
  .Z({ encrypted128[41] })
);
BUF_X1 #() 
BUF_X1_197_ (
  .A({ S790[42] }),
  .Z({ encrypted128[42] })
);
BUF_X1 #() 
BUF_X1_198_ (
  .A({ S790[43] }),
  .Z({ encrypted128[43] })
);
BUF_X1 #() 
BUF_X1_199_ (
  .A({ S790[44] }),
  .Z({ encrypted128[44] })
);
BUF_X1 #() 
BUF_X1_200_ (
  .A({ S790[45] }),
  .Z({ encrypted128[45] })
);
BUF_X1 #() 
BUF_X1_201_ (
  .A({ S790[46] }),
  .Z({ encrypted128[46] })
);
BUF_X1 #() 
BUF_X1_202_ (
  .A({ S790[47] }),
  .Z({ encrypted128[47] })
);
BUF_X1 #() 
BUF_X1_203_ (
  .A({ S790[48] }),
  .Z({ encrypted128[48] })
);
BUF_X1 #() 
BUF_X1_204_ (
  .A({ S790[49] }),
  .Z({ encrypted128[49] })
);
BUF_X1 #() 
BUF_X1_205_ (
  .A({ S790[5] }),
  .Z({ encrypted128[5] })
);
BUF_X1 #() 
BUF_X1_206_ (
  .A({ S790[50] }),
  .Z({ encrypted128[50] })
);
BUF_X1 #() 
BUF_X1_207_ (
  .A({ S790[51] }),
  .Z({ encrypted128[51] })
);
BUF_X1 #() 
BUF_X1_208_ (
  .A({ S790[52] }),
  .Z({ encrypted128[52] })
);
BUF_X1 #() 
BUF_X1_209_ (
  .A({ S790[53] }),
  .Z({ encrypted128[53] })
);
BUF_X1 #() 
BUF_X1_210_ (
  .A({ S790[54] }),
  .Z({ encrypted128[54] })
);
BUF_X1 #() 
BUF_X1_211_ (
  .A({ S790[55] }),
  .Z({ encrypted128[55] })
);
BUF_X1 #() 
BUF_X1_212_ (
  .A({ S790[56] }),
  .Z({ encrypted128[56] })
);
BUF_X1 #() 
BUF_X1_213_ (
  .A({ S790[57] }),
  .Z({ encrypted128[57] })
);
BUF_X1 #() 
BUF_X1_214_ (
  .A({ S790[58] }),
  .Z({ encrypted128[58] })
);
BUF_X1 #() 
BUF_X1_215_ (
  .A({ S790[59] }),
  .Z({ encrypted128[59] })
);
BUF_X1 #() 
BUF_X1_216_ (
  .A({ S790[6] }),
  .Z({ encrypted128[6] })
);
BUF_X1 #() 
BUF_X1_217_ (
  .A({ S790[60] }),
  .Z({ encrypted128[60] })
);
BUF_X1 #() 
BUF_X1_218_ (
  .A({ S790[61] }),
  .Z({ encrypted128[61] })
);
BUF_X1 #() 
BUF_X1_219_ (
  .A({ S790[62] }),
  .Z({ encrypted128[62] })
);
BUF_X1 #() 
BUF_X1_220_ (
  .A({ S790[63] }),
  .Z({ encrypted128[63] })
);
BUF_X1 #() 
BUF_X1_221_ (
  .A({ S790[64] }),
  .Z({ encrypted128[64] })
);
BUF_X1 #() 
BUF_X1_222_ (
  .A({ S790[65] }),
  .Z({ encrypted128[65] })
);
BUF_X1 #() 
BUF_X1_223_ (
  .A({ S790[66] }),
  .Z({ encrypted128[66] })
);
BUF_X1 #() 
BUF_X1_224_ (
  .A({ S790[67] }),
  .Z({ encrypted128[67] })
);
BUF_X1 #() 
BUF_X1_225_ (
  .A({ S790[68] }),
  .Z({ encrypted128[68] })
);
BUF_X1 #() 
BUF_X1_226_ (
  .A({ S790[69] }),
  .Z({ encrypted128[69] })
);
BUF_X1 #() 
BUF_X1_227_ (
  .A({ S790[7] }),
  .Z({ encrypted128[7] })
);
BUF_X1 #() 
BUF_X1_228_ (
  .A({ S790[70] }),
  .Z({ encrypted128[70] })
);
BUF_X1 #() 
BUF_X1_229_ (
  .A({ S790[71] }),
  .Z({ encrypted128[71] })
);
BUF_X1 #() 
BUF_X1_230_ (
  .A({ S790[72] }),
  .Z({ encrypted128[72] })
);
BUF_X1 #() 
BUF_X1_231_ (
  .A({ S790[73] }),
  .Z({ encrypted128[73] })
);
BUF_X1 #() 
BUF_X1_232_ (
  .A({ S790[74] }),
  .Z({ encrypted128[74] })
);
BUF_X1 #() 
BUF_X1_233_ (
  .A({ S790[75] }),
  .Z({ encrypted128[75] })
);
BUF_X1 #() 
BUF_X1_234_ (
  .A({ S790[76] }),
  .Z({ encrypted128[76] })
);
BUF_X1 #() 
BUF_X1_235_ (
  .A({ S790[77] }),
  .Z({ encrypted128[77] })
);
BUF_X1 #() 
BUF_X1_236_ (
  .A({ S790[78] }),
  .Z({ encrypted128[78] })
);
BUF_X1 #() 
BUF_X1_237_ (
  .A({ S790[79] }),
  .Z({ encrypted128[79] })
);
BUF_X1 #() 
BUF_X1_238_ (
  .A({ S790[8] }),
  .Z({ encrypted128[8] })
);
BUF_X1 #() 
BUF_X1_239_ (
  .A({ S790[80] }),
  .Z({ encrypted128[80] })
);
BUF_X1 #() 
BUF_X1_240_ (
  .A({ S790[81] }),
  .Z({ encrypted128[81] })
);
BUF_X1 #() 
BUF_X1_241_ (
  .A({ S790[82] }),
  .Z({ encrypted128[82] })
);
BUF_X1 #() 
BUF_X1_242_ (
  .A({ S790[83] }),
  .Z({ encrypted128[83] })
);
BUF_X1 #() 
BUF_X1_243_ (
  .A({ S790[84] }),
  .Z({ encrypted128[84] })
);
BUF_X1 #() 
BUF_X1_244_ (
  .A({ S790[85] }),
  .Z({ encrypted128[85] })
);
BUF_X1 #() 
BUF_X1_245_ (
  .A({ S790[86] }),
  .Z({ encrypted128[86] })
);
BUF_X1 #() 
BUF_X1_246_ (
  .A({ S790[87] }),
  .Z({ encrypted128[87] })
);
BUF_X1 #() 
BUF_X1_247_ (
  .A({ S790[88] }),
  .Z({ encrypted128[88] })
);
BUF_X1 #() 
BUF_X1_248_ (
  .A({ S790[89] }),
  .Z({ encrypted128[89] })
);
BUF_X1 #() 
BUF_X1_249_ (
  .A({ S790[9] }),
  .Z({ encrypted128[9] })
);
BUF_X1 #() 
BUF_X1_250_ (
  .A({ S790[90] }),
  .Z({ encrypted128[90] })
);
BUF_X1 #() 
BUF_X1_251_ (
  .A({ S790[91] }),
  .Z({ encrypted128[91] })
);
BUF_X1 #() 
BUF_X1_252_ (
  .A({ S790[92] }),
  .Z({ encrypted128[92] })
);
BUF_X1 #() 
BUF_X1_253_ (
  .A({ S790[93] }),
  .Z({ encrypted128[93] })
);
BUF_X1 #() 
BUF_X1_254_ (
  .A({ S790[94] }),
  .Z({ encrypted128[94] })
);
BUF_X1 #() 
BUF_X1_255_ (
  .A({ S790[95] }),
  .Z({ encrypted128[95] })
);
BUF_X1 #() 
BUF_X1_256_ (
  .A({ S790[96] }),
  .Z({ encrypted128[96] })
);
BUF_X1 #() 
BUF_X1_257_ (
  .A({ S790[97] }),
  .Z({ encrypted128[97] })
);
BUF_X1 #() 
BUF_X1_258_ (
  .A({ S790[98] }),
  .Z({ encrypted128[98] })
);
BUF_X1 #() 
BUF_X1_259_ (
  .A({ S790[99] }),
  .Z({ encrypted128[99] })
);
BUF_X1 #() 
BUF_X1_260_ (
  .A({ expected128[0] }),
  .Z({ S791[0] })
);
BUF_X1 #() 
BUF_X1_261_ (
  .A({ expected128[1] }),
  .Z({ S791[1] })
);
BUF_X1 #() 
BUF_X1_262_ (
  .A({ expected128[10] }),
  .Z({ S791[10] })
);
BUF_X1 #() 
BUF_X1_263_ (
  .A({ expected128[100] }),
  .Z({ S791[100] })
);
BUF_X1 #() 
BUF_X1_264_ (
  .A({ expected128[101] }),
  .Z({ S791[101] })
);
BUF_X1 #() 
BUF_X1_265_ (
  .A({ expected128[102] }),
  .Z({ S791[102] })
);
BUF_X1 #() 
BUF_X1_266_ (
  .A({ expected128[103] }),
  .Z({ S791[103] })
);
BUF_X1 #() 
BUF_X1_267_ (
  .A({ expected128[104] }),
  .Z({ S791[104] })
);
BUF_X1 #() 
BUF_X1_268_ (
  .A({ expected128[105] }),
  .Z({ S791[105] })
);
BUF_X1 #() 
BUF_X1_269_ (
  .A({ expected128[106] }),
  .Z({ S791[106] })
);
BUF_X1 #() 
BUF_X1_270_ (
  .A({ expected128[107] }),
  .Z({ S791[107] })
);
BUF_X1 #() 
BUF_X1_271_ (
  .A({ expected128[108] }),
  .Z({ S791[108] })
);
BUF_X1 #() 
BUF_X1_272_ (
  .A({ expected128[109] }),
  .Z({ S791[109] })
);
BUF_X1 #() 
BUF_X1_273_ (
  .A({ expected128[11] }),
  .Z({ S791[11] })
);
BUF_X1 #() 
BUF_X1_274_ (
  .A({ expected128[110] }),
  .Z({ S791[110] })
);
BUF_X1 #() 
BUF_X1_275_ (
  .A({ expected128[111] }),
  .Z({ S791[111] })
);
BUF_X1 #() 
BUF_X1_276_ (
  .A({ expected128[112] }),
  .Z({ S791[112] })
);
BUF_X1 #() 
BUF_X1_277_ (
  .A({ expected128[113] }),
  .Z({ S791[113] })
);
BUF_X1 #() 
BUF_X1_278_ (
  .A({ expected128[114] }),
  .Z({ S791[114] })
);
BUF_X1 #() 
BUF_X1_279_ (
  .A({ expected128[115] }),
  .Z({ S791[115] })
);
BUF_X1 #() 
BUF_X1_280_ (
  .A({ expected128[116] }),
  .Z({ S791[116] })
);
BUF_X1 #() 
BUF_X1_281_ (
  .A({ expected128[117] }),
  .Z({ S791[117] })
);
BUF_X1 #() 
BUF_X1_282_ (
  .A({ expected128[118] }),
  .Z({ S791[118] })
);
BUF_X1 #() 
BUF_X1_283_ (
  .A({ expected128[119] }),
  .Z({ S791[119] })
);
BUF_X1 #() 
BUF_X1_284_ (
  .A({ expected128[12] }),
  .Z({ S791[12] })
);
BUF_X1 #() 
BUF_X1_285_ (
  .A({ expected128[120] }),
  .Z({ S791[120] })
);
BUF_X1 #() 
BUF_X1_286_ (
  .A({ expected128[121] }),
  .Z({ S791[121] })
);
BUF_X1 #() 
BUF_X1_287_ (
  .A({ expected128[122] }),
  .Z({ S791[122] })
);
BUF_X1 #() 
BUF_X1_288_ (
  .A({ expected128[123] }),
  .Z({ S791[123] })
);
BUF_X1 #() 
BUF_X1_289_ (
  .A({ expected128[124] }),
  .Z({ S791[124] })
);
BUF_X1 #() 
BUF_X1_290_ (
  .A({ expected128[125] }),
  .Z({ S791[125] })
);
BUF_X1 #() 
BUF_X1_291_ (
  .A({ expected128[126] }),
  .Z({ S791[126] })
);
BUF_X1 #() 
BUF_X1_292_ (
  .A({ expected128[127] }),
  .Z({ S791[127] })
);
BUF_X1 #() 
BUF_X1_293_ (
  .A({ expected128[13] }),
  .Z({ S791[13] })
);
BUF_X1 #() 
BUF_X1_294_ (
  .A({ expected128[14] }),
  .Z({ S791[14] })
);
BUF_X1 #() 
BUF_X1_295_ (
  .A({ expected128[15] }),
  .Z({ S791[15] })
);
BUF_X1 #() 
BUF_X1_296_ (
  .A({ expected128[16] }),
  .Z({ S791[16] })
);
BUF_X1 #() 
BUF_X1_297_ (
  .A({ expected128[17] }),
  .Z({ S791[17] })
);
BUF_X1 #() 
BUF_X1_298_ (
  .A({ expected128[18] }),
  .Z({ S791[18] })
);
BUF_X1 #() 
BUF_X1_299_ (
  .A({ expected128[19] }),
  .Z({ S791[19] })
);
BUF_X1 #() 
BUF_X1_300_ (
  .A({ expected128[2] }),
  .Z({ S791[2] })
);
BUF_X1 #() 
BUF_X1_301_ (
  .A({ expected128[20] }),
  .Z({ S791[20] })
);
BUF_X1 #() 
BUF_X1_302_ (
  .A({ expected128[21] }),
  .Z({ S791[21] })
);
BUF_X1 #() 
BUF_X1_303_ (
  .A({ expected128[22] }),
  .Z({ S791[22] })
);
BUF_X1 #() 
BUF_X1_304_ (
  .A({ expected128[23] }),
  .Z({ S791[23] })
);
BUF_X1 #() 
BUF_X1_305_ (
  .A({ expected128[24] }),
  .Z({ S791[24] })
);
BUF_X1 #() 
BUF_X1_306_ (
  .A({ expected128[25] }),
  .Z({ S791[25] })
);
BUF_X1 #() 
BUF_X1_307_ (
  .A({ expected128[26] }),
  .Z({ S791[26] })
);
BUF_X1 #() 
BUF_X1_308_ (
  .A({ expected128[27] }),
  .Z({ S791[27] })
);
BUF_X1 #() 
BUF_X1_309_ (
  .A({ expected128[28] }),
  .Z({ S791[28] })
);
BUF_X1 #() 
BUF_X1_310_ (
  .A({ expected128[29] }),
  .Z({ S791[29] })
);
BUF_X1 #() 
BUF_X1_311_ (
  .A({ expected128[3] }),
  .Z({ S791[3] })
);
BUF_X1 #() 
BUF_X1_312_ (
  .A({ expected128[30] }),
  .Z({ S791[30] })
);
BUF_X1 #() 
BUF_X1_313_ (
  .A({ expected128[31] }),
  .Z({ S791[31] })
);
BUF_X1 #() 
BUF_X1_314_ (
  .A({ expected128[32] }),
  .Z({ S791[32] })
);
BUF_X1 #() 
BUF_X1_315_ (
  .A({ expected128[33] }),
  .Z({ S791[33] })
);
BUF_X1 #() 
BUF_X1_316_ (
  .A({ expected128[34] }),
  .Z({ S791[34] })
);
BUF_X1 #() 
BUF_X1_317_ (
  .A({ expected128[35] }),
  .Z({ S791[35] })
);
BUF_X1 #() 
BUF_X1_318_ (
  .A({ expected128[36] }),
  .Z({ S791[36] })
);
BUF_X1 #() 
BUF_X1_319_ (
  .A({ expected128[37] }),
  .Z({ S791[37] })
);
BUF_X1 #() 
BUF_X1_320_ (
  .A({ expected128[38] }),
  .Z({ S791[38] })
);
BUF_X1 #() 
BUF_X1_321_ (
  .A({ expected128[39] }),
  .Z({ S791[39] })
);
BUF_X1 #() 
BUF_X1_322_ (
  .A({ expected128[4] }),
  .Z({ S791[4] })
);
BUF_X1 #() 
BUF_X1_323_ (
  .A({ expected128[40] }),
  .Z({ S791[40] })
);
BUF_X1 #() 
BUF_X1_324_ (
  .A({ expected128[41] }),
  .Z({ S791[41] })
);
BUF_X1 #() 
BUF_X1_325_ (
  .A({ expected128[42] }),
  .Z({ S791[42] })
);
BUF_X1 #() 
BUF_X1_326_ (
  .A({ expected128[43] }),
  .Z({ S791[43] })
);
BUF_X1 #() 
BUF_X1_327_ (
  .A({ expected128[44] }),
  .Z({ S791[44] })
);
BUF_X1 #() 
BUF_X1_328_ (
  .A({ expected128[45] }),
  .Z({ S791[45] })
);
BUF_X1 #() 
BUF_X1_329_ (
  .A({ expected128[46] }),
  .Z({ S791[46] })
);
BUF_X1 #() 
BUF_X1_330_ (
  .A({ expected128[47] }),
  .Z({ S791[47] })
);
BUF_X1 #() 
BUF_X1_331_ (
  .A({ expected128[48] }),
  .Z({ S791[48] })
);
BUF_X1 #() 
BUF_X1_332_ (
  .A({ expected128[49] }),
  .Z({ S791[49] })
);
BUF_X1 #() 
BUF_X1_333_ (
  .A({ expected128[5] }),
  .Z({ S791[5] })
);
BUF_X1 #() 
BUF_X1_334_ (
  .A({ expected128[50] }),
  .Z({ S791[50] })
);
BUF_X1 #() 
BUF_X1_335_ (
  .A({ expected128[51] }),
  .Z({ S791[51] })
);
BUF_X1 #() 
BUF_X1_336_ (
  .A({ expected128[52] }),
  .Z({ S791[52] })
);
BUF_X1 #() 
BUF_X1_337_ (
  .A({ expected128[53] }),
  .Z({ S791[53] })
);
BUF_X1 #() 
BUF_X1_338_ (
  .A({ expected128[54] }),
  .Z({ S791[54] })
);
BUF_X1 #() 
BUF_X1_339_ (
  .A({ expected128[55] }),
  .Z({ S791[55] })
);
BUF_X1 #() 
BUF_X1_340_ (
  .A({ expected128[56] }),
  .Z({ S791[56] })
);
BUF_X1 #() 
BUF_X1_341_ (
  .A({ expected128[57] }),
  .Z({ S791[57] })
);
BUF_X1 #() 
BUF_X1_342_ (
  .A({ expected128[58] }),
  .Z({ S791[58] })
);
BUF_X1 #() 
BUF_X1_343_ (
  .A({ expected128[59] }),
  .Z({ S791[59] })
);
BUF_X1 #() 
BUF_X1_344_ (
  .A({ expected128[6] }),
  .Z({ S791[6] })
);
BUF_X1 #() 
BUF_X1_345_ (
  .A({ expected128[60] }),
  .Z({ S791[60] })
);
BUF_X1 #() 
BUF_X1_346_ (
  .A({ expected128[61] }),
  .Z({ S791[61] })
);
BUF_X1 #() 
BUF_X1_347_ (
  .A({ expected128[62] }),
  .Z({ S791[62] })
);
BUF_X1 #() 
BUF_X1_348_ (
  .A({ expected128[63] }),
  .Z({ S791[63] })
);
BUF_X1 #() 
BUF_X1_349_ (
  .A({ expected128[64] }),
  .Z({ S791[64] })
);
BUF_X1 #() 
BUF_X1_350_ (
  .A({ expected128[65] }),
  .Z({ S791[65] })
);
BUF_X1 #() 
BUF_X1_351_ (
  .A({ expected128[66] }),
  .Z({ S791[66] })
);
BUF_X1 #() 
BUF_X1_352_ (
  .A({ expected128[67] }),
  .Z({ S791[67] })
);
BUF_X1 #() 
BUF_X1_353_ (
  .A({ expected128[68] }),
  .Z({ S791[68] })
);
BUF_X1 #() 
BUF_X1_354_ (
  .A({ expected128[69] }),
  .Z({ S791[69] })
);
BUF_X1 #() 
BUF_X1_355_ (
  .A({ expected128[7] }),
  .Z({ S791[7] })
);
BUF_X1 #() 
BUF_X1_356_ (
  .A({ expected128[70] }),
  .Z({ S791[70] })
);
BUF_X1 #() 
BUF_X1_357_ (
  .A({ expected128[71] }),
  .Z({ S791[71] })
);
BUF_X1 #() 
BUF_X1_358_ (
  .A({ expected128[72] }),
  .Z({ S791[72] })
);
BUF_X1 #() 
BUF_X1_359_ (
  .A({ expected128[73] }),
  .Z({ S791[73] })
);
BUF_X1 #() 
BUF_X1_360_ (
  .A({ expected128[74] }),
  .Z({ S791[74] })
);
BUF_X1 #() 
BUF_X1_361_ (
  .A({ expected128[75] }),
  .Z({ S791[75] })
);
BUF_X1 #() 
BUF_X1_362_ (
  .A({ expected128[76] }),
  .Z({ S791[76] })
);
BUF_X1 #() 
BUF_X1_363_ (
  .A({ expected128[77] }),
  .Z({ S791[77] })
);
BUF_X1 #() 
BUF_X1_364_ (
  .A({ expected128[78] }),
  .Z({ S791[78] })
);
BUF_X1 #() 
BUF_X1_365_ (
  .A({ expected128[79] }),
  .Z({ S791[79] })
);
BUF_X1 #() 
BUF_X1_366_ (
  .A({ expected128[8] }),
  .Z({ S791[8] })
);
BUF_X1 #() 
BUF_X1_367_ (
  .A({ expected128[80] }),
  .Z({ S791[80] })
);
BUF_X1 #() 
BUF_X1_368_ (
  .A({ expected128[81] }),
  .Z({ S791[81] })
);
BUF_X1 #() 
BUF_X1_369_ (
  .A({ expected128[82] }),
  .Z({ S791[82] })
);
BUF_X1 #() 
BUF_X1_370_ (
  .A({ expected128[83] }),
  .Z({ S791[83] })
);
BUF_X1 #() 
BUF_X1_371_ (
  .A({ expected128[84] }),
  .Z({ S791[84] })
);
BUF_X1 #() 
BUF_X1_372_ (
  .A({ expected128[85] }),
  .Z({ S791[85] })
);
BUF_X1 #() 
BUF_X1_373_ (
  .A({ expected128[86] }),
  .Z({ S791[86] })
);
BUF_X1 #() 
BUF_X1_374_ (
  .A({ expected128[87] }),
  .Z({ S791[87] })
);
BUF_X1 #() 
BUF_X1_375_ (
  .A({ expected128[88] }),
  .Z({ S791[88] })
);
BUF_X1 #() 
BUF_X1_376_ (
  .A({ expected128[89] }),
  .Z({ S791[89] })
);
BUF_X1 #() 
BUF_X1_377_ (
  .A({ expected128[9] }),
  .Z({ S791[9] })
);
BUF_X1 #() 
BUF_X1_378_ (
  .A({ expected128[90] }),
  .Z({ S791[90] })
);
BUF_X1 #() 
BUF_X1_379_ (
  .A({ expected128[91] }),
  .Z({ S791[91] })
);
BUF_X1 #() 
BUF_X1_380_ (
  .A({ expected128[92] }),
  .Z({ S791[92] })
);
BUF_X1 #() 
BUF_X1_381_ (
  .A({ expected128[93] }),
  .Z({ S791[93] })
);
BUF_X1 #() 
BUF_X1_382_ (
  .A({ expected128[94] }),
  .Z({ S791[94] })
);
BUF_X1 #() 
BUF_X1_383_ (
  .A({ expected128[95] }),
  .Z({ S791[95] })
);
BUF_X1 #() 
BUF_X1_384_ (
  .A({ expected128[96] }),
  .Z({ S791[96] })
);
BUF_X1 #() 
BUF_X1_385_ (
  .A({ expected128[97] }),
  .Z({ S791[97] })
);
BUF_X1 #() 
BUF_X1_386_ (
  .A({ expected128[98] }),
  .Z({ S791[98] })
);
BUF_X1 #() 
BUF_X1_387_ (
  .A({ expected128[99] }),
  .Z({ S791[99] })
);
BUF_X1 #() 
BUF_X1_388_ (
  .A({ in[0] }),
  .Z({ S792[0] })
);
BUF_X1 #() 
BUF_X1_389_ (
  .A({ in[1] }),
  .Z({ S792[1] })
);
BUF_X1 #() 
BUF_X1_390_ (
  .A({ in[10] }),
  .Z({ S792[10] })
);
BUF_X1 #() 
BUF_X1_391_ (
  .A({ in[100] }),
  .Z({ S792[100] })
);
BUF_X1 #() 
BUF_X1_392_ (
  .A({ in[101] }),
  .Z({ S792[101] })
);
BUF_X1 #() 
BUF_X1_393_ (
  .A({ in[102] }),
  .Z({ S792[102] })
);
BUF_X1 #() 
BUF_X1_394_ (
  .A({ in[103] }),
  .Z({ S792[103] })
);
BUF_X1 #() 
BUF_X1_395_ (
  .A({ in[104] }),
  .Z({ S792[104] })
);
BUF_X1 #() 
BUF_X1_396_ (
  .A({ in[105] }),
  .Z({ S792[105] })
);
BUF_X1 #() 
BUF_X1_397_ (
  .A({ in[106] }),
  .Z({ S792[106] })
);
BUF_X1 #() 
BUF_X1_398_ (
  .A({ in[107] }),
  .Z({ S792[107] })
);
BUF_X1 #() 
BUF_X1_399_ (
  .A({ in[108] }),
  .Z({ S792[108] })
);
BUF_X1 #() 
BUF_X1_400_ (
  .A({ in[109] }),
  .Z({ S792[109] })
);
BUF_X1 #() 
BUF_X1_401_ (
  .A({ in[11] }),
  .Z({ S792[11] })
);
BUF_X1 #() 
BUF_X1_402_ (
  .A({ in[110] }),
  .Z({ S792[110] })
);
BUF_X1 #() 
BUF_X1_403_ (
  .A({ in[111] }),
  .Z({ S792[111] })
);
BUF_X1 #() 
BUF_X1_404_ (
  .A({ in[112] }),
  .Z({ S792[112] })
);
BUF_X1 #() 
BUF_X1_405_ (
  .A({ in[113] }),
  .Z({ S792[113] })
);
BUF_X1 #() 
BUF_X1_406_ (
  .A({ in[114] }),
  .Z({ S792[114] })
);
BUF_X1 #() 
BUF_X1_407_ (
  .A({ in[115] }),
  .Z({ S792[115] })
);
BUF_X1 #() 
BUF_X1_408_ (
  .A({ in[116] }),
  .Z({ S792[116] })
);
BUF_X1 #() 
BUF_X1_409_ (
  .A({ in[117] }),
  .Z({ S792[117] })
);
BUF_X1 #() 
BUF_X1_410_ (
  .A({ in[118] }),
  .Z({ S792[118] })
);
BUF_X1 #() 
BUF_X1_411_ (
  .A({ in[119] }),
  .Z({ S792[119] })
);
BUF_X1 #() 
BUF_X1_412_ (
  .A({ in[12] }),
  .Z({ S792[12] })
);
BUF_X1 #() 
BUF_X1_413_ (
  .A({ in[120] }),
  .Z({ S792[120] })
);
BUF_X1 #() 
BUF_X1_414_ (
  .A({ in[121] }),
  .Z({ S792[121] })
);
BUF_X1 #() 
BUF_X1_415_ (
  .A({ in[122] }),
  .Z({ S792[122] })
);
BUF_X1 #() 
BUF_X1_416_ (
  .A({ in[123] }),
  .Z({ S792[123] })
);
BUF_X1 #() 
BUF_X1_417_ (
  .A({ in[124] }),
  .Z({ S792[124] })
);
BUF_X1 #() 
BUF_X1_418_ (
  .A({ in[125] }),
  .Z({ S792[125] })
);
BUF_X1 #() 
BUF_X1_419_ (
  .A({ in[126] }),
  .Z({ S792[126] })
);
BUF_X1 #() 
BUF_X1_420_ (
  .A({ in[127] }),
  .Z({ S792[127] })
);
BUF_X1 #() 
BUF_X1_421_ (
  .A({ in[13] }),
  .Z({ S792[13] })
);
BUF_X1 #() 
BUF_X1_422_ (
  .A({ in[14] }),
  .Z({ S792[14] })
);
BUF_X1 #() 
BUF_X1_423_ (
  .A({ in[15] }),
  .Z({ S792[15] })
);
BUF_X1 #() 
BUF_X1_424_ (
  .A({ in[16] }),
  .Z({ S792[16] })
);
BUF_X1 #() 
BUF_X1_425_ (
  .A({ in[17] }),
  .Z({ S792[17] })
);
BUF_X1 #() 
BUF_X1_426_ (
  .A({ in[18] }),
  .Z({ S792[18] })
);
BUF_X1 #() 
BUF_X1_427_ (
  .A({ in[19] }),
  .Z({ S792[19] })
);
BUF_X1 #() 
BUF_X1_428_ (
  .A({ in[2] }),
  .Z({ S792[2] })
);
BUF_X1 #() 
BUF_X1_429_ (
  .A({ in[20] }),
  .Z({ S792[20] })
);
BUF_X1 #() 
BUF_X1_430_ (
  .A({ in[21] }),
  .Z({ S792[21] })
);
BUF_X1 #() 
BUF_X1_431_ (
  .A({ in[22] }),
  .Z({ S792[22] })
);
BUF_X1 #() 
BUF_X1_432_ (
  .A({ in[23] }),
  .Z({ S792[23] })
);
BUF_X1 #() 
BUF_X1_433_ (
  .A({ in[24] }),
  .Z({ S792[24] })
);
BUF_X1 #() 
BUF_X1_434_ (
  .A({ in[25] }),
  .Z({ S792[25] })
);
BUF_X1 #() 
BUF_X1_435_ (
  .A({ in[26] }),
  .Z({ S792[26] })
);
BUF_X1 #() 
BUF_X1_436_ (
  .A({ in[27] }),
  .Z({ S792[27] })
);
BUF_X1 #() 
BUF_X1_437_ (
  .A({ in[28] }),
  .Z({ S792[28] })
);
BUF_X1 #() 
BUF_X1_438_ (
  .A({ in[29] }),
  .Z({ S792[29] })
);
BUF_X1 #() 
BUF_X1_439_ (
  .A({ in[3] }),
  .Z({ S792[3] })
);
BUF_X1 #() 
BUF_X1_440_ (
  .A({ in[30] }),
  .Z({ S792[30] })
);
BUF_X1 #() 
BUF_X1_441_ (
  .A({ in[31] }),
  .Z({ S792[31] })
);
BUF_X1 #() 
BUF_X1_442_ (
  .A({ in[32] }),
  .Z({ S792[32] })
);
BUF_X1 #() 
BUF_X1_443_ (
  .A({ in[33] }),
  .Z({ S792[33] })
);
BUF_X1 #() 
BUF_X1_444_ (
  .A({ in[34] }),
  .Z({ S792[34] })
);
BUF_X1 #() 
BUF_X1_445_ (
  .A({ in[35] }),
  .Z({ S792[35] })
);
BUF_X1 #() 
BUF_X1_446_ (
  .A({ in[36] }),
  .Z({ S792[36] })
);
BUF_X1 #() 
BUF_X1_447_ (
  .A({ in[37] }),
  .Z({ S792[37] })
);
BUF_X1 #() 
BUF_X1_448_ (
  .A({ in[38] }),
  .Z({ S792[38] })
);
BUF_X1 #() 
BUF_X1_449_ (
  .A({ in[39] }),
  .Z({ S792[39] })
);
BUF_X1 #() 
BUF_X1_450_ (
  .A({ in[4] }),
  .Z({ S792[4] })
);
BUF_X1 #() 
BUF_X1_451_ (
  .A({ in[40] }),
  .Z({ S792[40] })
);
BUF_X1 #() 
BUF_X1_452_ (
  .A({ in[41] }),
  .Z({ S792[41] })
);
BUF_X1 #() 
BUF_X1_453_ (
  .A({ in[42] }),
  .Z({ S792[42] })
);
BUF_X1 #() 
BUF_X1_454_ (
  .A({ in[43] }),
  .Z({ S792[43] })
);
BUF_X1 #() 
BUF_X1_455_ (
  .A({ in[44] }),
  .Z({ S792[44] })
);
BUF_X1 #() 
BUF_X1_456_ (
  .A({ in[45] }),
  .Z({ S792[45] })
);
BUF_X1 #() 
BUF_X1_457_ (
  .A({ in[46] }),
  .Z({ S792[46] })
);
BUF_X1 #() 
BUF_X1_458_ (
  .A({ in[47] }),
  .Z({ S792[47] })
);
BUF_X1 #() 
BUF_X1_459_ (
  .A({ in[48] }),
  .Z({ S792[48] })
);
BUF_X1 #() 
BUF_X1_460_ (
  .A({ in[49] }),
  .Z({ S792[49] })
);
BUF_X1 #() 
BUF_X1_461_ (
  .A({ in[5] }),
  .Z({ S792[5] })
);
BUF_X1 #() 
BUF_X1_462_ (
  .A({ in[50] }),
  .Z({ S792[50] })
);
BUF_X1 #() 
BUF_X1_463_ (
  .A({ in[51] }),
  .Z({ S792[51] })
);
BUF_X1 #() 
BUF_X1_464_ (
  .A({ in[52] }),
  .Z({ S792[52] })
);
BUF_X1 #() 
BUF_X1_465_ (
  .A({ in[53] }),
  .Z({ S792[53] })
);
BUF_X1 #() 
BUF_X1_466_ (
  .A({ in[54] }),
  .Z({ S792[54] })
);
BUF_X1 #() 
BUF_X1_467_ (
  .A({ in[55] }),
  .Z({ S792[55] })
);
BUF_X1 #() 
BUF_X1_468_ (
  .A({ in[56] }),
  .Z({ S792[56] })
);
BUF_X1 #() 
BUF_X1_469_ (
  .A({ in[57] }),
  .Z({ S792[57] })
);
BUF_X1 #() 
BUF_X1_470_ (
  .A({ in[58] }),
  .Z({ S792[58] })
);
BUF_X1 #() 
BUF_X1_471_ (
  .A({ in[59] }),
  .Z({ S792[59] })
);
BUF_X1 #() 
BUF_X1_472_ (
  .A({ in[6] }),
  .Z({ S792[6] })
);
BUF_X1 #() 
BUF_X1_473_ (
  .A({ in[60] }),
  .Z({ S792[60] })
);
BUF_X1 #() 
BUF_X1_474_ (
  .A({ in[61] }),
  .Z({ S792[61] })
);
BUF_X1 #() 
BUF_X1_475_ (
  .A({ in[62] }),
  .Z({ S792[62] })
);
BUF_X1 #() 
BUF_X1_476_ (
  .A({ in[63] }),
  .Z({ S792[63] })
);
BUF_X1 #() 
BUF_X1_477_ (
  .A({ in[64] }),
  .Z({ S792[64] })
);
BUF_X1 #() 
BUF_X1_478_ (
  .A({ in[65] }),
  .Z({ S792[65] })
);
BUF_X1 #() 
BUF_X1_479_ (
  .A({ in[66] }),
  .Z({ S792[66] })
);
BUF_X1 #() 
BUF_X1_480_ (
  .A({ in[67] }),
  .Z({ S792[67] })
);
BUF_X1 #() 
BUF_X1_481_ (
  .A({ in[68] }),
  .Z({ S792[68] })
);
BUF_X1 #() 
BUF_X1_482_ (
  .A({ in[69] }),
  .Z({ S792[69] })
);
BUF_X1 #() 
BUF_X1_483_ (
  .A({ in[7] }),
  .Z({ S792[7] })
);
BUF_X1 #() 
BUF_X1_484_ (
  .A({ in[70] }),
  .Z({ S792[70] })
);
BUF_X1 #() 
BUF_X1_485_ (
  .A({ in[71] }),
  .Z({ S792[71] })
);
BUF_X1 #() 
BUF_X1_486_ (
  .A({ in[72] }),
  .Z({ S792[72] })
);
BUF_X1 #() 
BUF_X1_487_ (
  .A({ in[73] }),
  .Z({ S792[73] })
);
BUF_X1 #() 
BUF_X1_488_ (
  .A({ in[74] }),
  .Z({ S792[74] })
);
BUF_X1 #() 
BUF_X1_489_ (
  .A({ in[75] }),
  .Z({ S792[75] })
);
BUF_X1 #() 
BUF_X1_490_ (
  .A({ in[76] }),
  .Z({ S792[76] })
);
BUF_X1 #() 
BUF_X1_491_ (
  .A({ in[77] }),
  .Z({ S792[77] })
);
BUF_X1 #() 
BUF_X1_492_ (
  .A({ in[78] }),
  .Z({ S792[78] })
);
BUF_X1 #() 
BUF_X1_493_ (
  .A({ in[79] }),
  .Z({ S792[79] })
);
BUF_X1 #() 
BUF_X1_494_ (
  .A({ in[8] }),
  .Z({ S792[8] })
);
BUF_X1 #() 
BUF_X1_495_ (
  .A({ in[80] }),
  .Z({ S792[80] })
);
BUF_X1 #() 
BUF_X1_496_ (
  .A({ in[81] }),
  .Z({ S792[81] })
);
BUF_X1 #() 
BUF_X1_497_ (
  .A({ in[82] }),
  .Z({ S792[82] })
);
BUF_X1 #() 
BUF_X1_498_ (
  .A({ in[83] }),
  .Z({ S792[83] })
);
BUF_X1 #() 
BUF_X1_499_ (
  .A({ in[84] }),
  .Z({ S792[84] })
);
BUF_X1 #() 
BUF_X1_500_ (
  .A({ in[85] }),
  .Z({ S792[85] })
);
BUF_X1 #() 
BUF_X1_501_ (
  .A({ in[86] }),
  .Z({ S792[86] })
);
BUF_X1 #() 
BUF_X1_502_ (
  .A({ in[87] }),
  .Z({ S792[87] })
);
BUF_X1 #() 
BUF_X1_503_ (
  .A({ in[88] }),
  .Z({ S792[88] })
);
BUF_X1 #() 
BUF_X1_504_ (
  .A({ in[89] }),
  .Z({ S792[89] })
);
BUF_X1 #() 
BUF_X1_505_ (
  .A({ in[9] }),
  .Z({ S792[9] })
);
BUF_X1 #() 
BUF_X1_506_ (
  .A({ in[90] }),
  .Z({ S792[90] })
);
BUF_X1 #() 
BUF_X1_507_ (
  .A({ in[91] }),
  .Z({ S792[91] })
);
BUF_X1 #() 
BUF_X1_508_ (
  .A({ in[92] }),
  .Z({ S792[92] })
);
BUF_X1 #() 
BUF_X1_509_ (
  .A({ in[93] }),
  .Z({ S792[93] })
);
BUF_X1 #() 
BUF_X1_510_ (
  .A({ in[94] }),
  .Z({ S792[94] })
);
BUF_X1 #() 
BUF_X1_511_ (
  .A({ in[95] }),
  .Z({ S792[95] })
);
BUF_X1 #() 
BUF_X1_512_ (
  .A({ in[96] }),
  .Z({ S792[96] })
);
BUF_X1 #() 
BUF_X1_513_ (
  .A({ in[97] }),
  .Z({ S792[97] })
);
BUF_X1 #() 
BUF_X1_514_ (
  .A({ in[98] }),
  .Z({ S792[98] })
);
BUF_X1 #() 
BUF_X1_515_ (
  .A({ in[99] }),
  .Z({ S792[99] })
);
BUF_X1 #() 
BUF_X1_516_ (
  .A({ key128[0] }),
  .Z({ S793[0] })
);
BUF_X1 #() 
BUF_X1_517_ (
  .A({ key128[1] }),
  .Z({ S793[1] })
);
BUF_X1 #() 
BUF_X1_518_ (
  .A({ key128[10] }),
  .Z({ S793[10] })
);
BUF_X1 #() 
BUF_X1_519_ (
  .A({ key128[100] }),
  .Z({ S793[100] })
);
BUF_X1 #() 
BUF_X1_520_ (
  .A({ key128[101] }),
  .Z({ S793[101] })
);
BUF_X1 #() 
BUF_X1_521_ (
  .A({ key128[102] }),
  .Z({ S793[102] })
);
BUF_X1 #() 
BUF_X1_522_ (
  .A({ key128[103] }),
  .Z({ S793[103] })
);
BUF_X1 #() 
BUF_X1_523_ (
  .A({ key128[104] }),
  .Z({ S793[104] })
);
BUF_X1 #() 
BUF_X1_524_ (
  .A({ key128[105] }),
  .Z({ S793[105] })
);
BUF_X1 #() 
BUF_X1_525_ (
  .A({ key128[106] }),
  .Z({ S793[106] })
);
BUF_X1 #() 
BUF_X1_526_ (
  .A({ key128[107] }),
  .Z({ S793[107] })
);
BUF_X1 #() 
BUF_X1_527_ (
  .A({ key128[108] }),
  .Z({ S793[108] })
);
BUF_X1 #() 
BUF_X1_528_ (
  .A({ key128[109] }),
  .Z({ S793[109] })
);
BUF_X1 #() 
BUF_X1_529_ (
  .A({ key128[11] }),
  .Z({ S793[11] })
);
BUF_X1 #() 
BUF_X1_530_ (
  .A({ key128[110] }),
  .Z({ S793[110] })
);
BUF_X1 #() 
BUF_X1_531_ (
  .A({ key128[111] }),
  .Z({ S793[111] })
);
BUF_X1 #() 
BUF_X1_532_ (
  .A({ key128[112] }),
  .Z({ S793[112] })
);
BUF_X1 #() 
BUF_X1_533_ (
  .A({ key128[113] }),
  .Z({ S793[113] })
);
BUF_X1 #() 
BUF_X1_534_ (
  .A({ key128[114] }),
  .Z({ S793[114] })
);
BUF_X1 #() 
BUF_X1_535_ (
  .A({ key128[115] }),
  .Z({ S793[115] })
);
BUF_X1 #() 
BUF_X1_536_ (
  .A({ key128[116] }),
  .Z({ S793[116] })
);
BUF_X1 #() 
BUF_X1_537_ (
  .A({ key128[117] }),
  .Z({ S793[117] })
);
BUF_X1 #() 
BUF_X1_538_ (
  .A({ key128[118] }),
  .Z({ S793[118] })
);
BUF_X1 #() 
BUF_X1_539_ (
  .A({ key128[119] }),
  .Z({ S793[119] })
);
BUF_X1 #() 
BUF_X1_540_ (
  .A({ key128[12] }),
  .Z({ S793[12] })
);
BUF_X1 #() 
BUF_X1_541_ (
  .A({ key128[120] }),
  .Z({ S793[120] })
);
BUF_X1 #() 
BUF_X1_542_ (
  .A({ key128[121] }),
  .Z({ S793[121] })
);
BUF_X1 #() 
BUF_X1_543_ (
  .A({ key128[122] }),
  .Z({ S793[122] })
);
BUF_X1 #() 
BUF_X1_544_ (
  .A({ key128[123] }),
  .Z({ S793[123] })
);
BUF_X1 #() 
BUF_X1_545_ (
  .A({ key128[124] }),
  .Z({ S793[124] })
);
BUF_X1 #() 
BUF_X1_546_ (
  .A({ key128[125] }),
  .Z({ S793[125] })
);
BUF_X1 #() 
BUF_X1_547_ (
  .A({ key128[126] }),
  .Z({ S793[126] })
);
BUF_X1 #() 
BUF_X1_548_ (
  .A({ key128[127] }),
  .Z({ S793[127] })
);
BUF_X1 #() 
BUF_X1_549_ (
  .A({ key128[13] }),
  .Z({ S793[13] })
);
BUF_X1 #() 
BUF_X1_550_ (
  .A({ key128[14] }),
  .Z({ S793[14] })
);
BUF_X1 #() 
BUF_X1_551_ (
  .A({ key128[15] }),
  .Z({ S793[15] })
);
BUF_X1 #() 
BUF_X1_552_ (
  .A({ key128[16] }),
  .Z({ S793[16] })
);
BUF_X1 #() 
BUF_X1_553_ (
  .A({ key128[17] }),
  .Z({ S793[17] })
);
BUF_X1 #() 
BUF_X1_554_ (
  .A({ key128[18] }),
  .Z({ S793[18] })
);
BUF_X1 #() 
BUF_X1_555_ (
  .A({ key128[19] }),
  .Z({ S793[19] })
);
BUF_X1 #() 
BUF_X1_556_ (
  .A({ key128[2] }),
  .Z({ S793[2] })
);
BUF_X1 #() 
BUF_X1_557_ (
  .A({ key128[20] }),
  .Z({ S793[20] })
);
BUF_X1 #() 
BUF_X1_558_ (
  .A({ key128[21] }),
  .Z({ S793[21] })
);
BUF_X1 #() 
BUF_X1_559_ (
  .A({ key128[22] }),
  .Z({ S793[22] })
);
BUF_X1 #() 
BUF_X1_560_ (
  .A({ key128[23] }),
  .Z({ S793[23] })
);
BUF_X1 #() 
BUF_X1_561_ (
  .A({ key128[24] }),
  .Z({ S793[24] })
);
BUF_X1 #() 
BUF_X1_562_ (
  .A({ key128[25] }),
  .Z({ S793[25] })
);
BUF_X1 #() 
BUF_X1_563_ (
  .A({ key128[26] }),
  .Z({ S793[26] })
);
BUF_X1 #() 
BUF_X1_564_ (
  .A({ key128[27] }),
  .Z({ S793[27] })
);
BUF_X1 #() 
BUF_X1_565_ (
  .A({ key128[28] }),
  .Z({ S793[28] })
);
BUF_X1 #() 
BUF_X1_566_ (
  .A({ key128[29] }),
  .Z({ S793[29] })
);
BUF_X1 #() 
BUF_X1_567_ (
  .A({ key128[3] }),
  .Z({ S793[3] })
);
BUF_X1 #() 
BUF_X1_568_ (
  .A({ key128[30] }),
  .Z({ S793[30] })
);
BUF_X1 #() 
BUF_X1_569_ (
  .A({ key128[31] }),
  .Z({ S793[31] })
);
BUF_X1 #() 
BUF_X1_570_ (
  .A({ key128[32] }),
  .Z({ S793[32] })
);
BUF_X1 #() 
BUF_X1_571_ (
  .A({ key128[33] }),
  .Z({ S793[33] })
);
BUF_X1 #() 
BUF_X1_572_ (
  .A({ key128[34] }),
  .Z({ S793[34] })
);
BUF_X1 #() 
BUF_X1_573_ (
  .A({ key128[35] }),
  .Z({ S793[35] })
);
BUF_X1 #() 
BUF_X1_574_ (
  .A({ key128[36] }),
  .Z({ S793[36] })
);
BUF_X1 #() 
BUF_X1_575_ (
  .A({ key128[37] }),
  .Z({ S793[37] })
);
BUF_X1 #() 
BUF_X1_576_ (
  .A({ key128[38] }),
  .Z({ S793[38] })
);
BUF_X1 #() 
BUF_X1_577_ (
  .A({ key128[39] }),
  .Z({ S793[39] })
);
BUF_X1 #() 
BUF_X1_578_ (
  .A({ key128[4] }),
  .Z({ S793[4] })
);
BUF_X1 #() 
BUF_X1_579_ (
  .A({ key128[40] }),
  .Z({ S793[40] })
);
BUF_X1 #() 
BUF_X1_580_ (
  .A({ key128[41] }),
  .Z({ S793[41] })
);
BUF_X1 #() 
BUF_X1_581_ (
  .A({ key128[42] }),
  .Z({ S793[42] })
);
BUF_X1 #() 
BUF_X1_582_ (
  .A({ key128[43] }),
  .Z({ S793[43] })
);
BUF_X1 #() 
BUF_X1_583_ (
  .A({ key128[44] }),
  .Z({ S793[44] })
);
BUF_X1 #() 
BUF_X1_584_ (
  .A({ key128[45] }),
  .Z({ S793[45] })
);
BUF_X1 #() 
BUF_X1_585_ (
  .A({ key128[46] }),
  .Z({ S793[46] })
);
BUF_X1 #() 
BUF_X1_586_ (
  .A({ key128[47] }),
  .Z({ S793[47] })
);
BUF_X1 #() 
BUF_X1_587_ (
  .A({ key128[48] }),
  .Z({ S793[48] })
);
BUF_X1 #() 
BUF_X1_588_ (
  .A({ key128[49] }),
  .Z({ S793[49] })
);
BUF_X1 #() 
BUF_X1_589_ (
  .A({ key128[5] }),
  .Z({ S793[5] })
);
BUF_X1 #() 
BUF_X1_590_ (
  .A({ key128[50] }),
  .Z({ S793[50] })
);
BUF_X1 #() 
BUF_X1_591_ (
  .A({ key128[51] }),
  .Z({ S793[51] })
);
BUF_X1 #() 
BUF_X1_592_ (
  .A({ key128[52] }),
  .Z({ S793[52] })
);
BUF_X1 #() 
BUF_X1_593_ (
  .A({ key128[53] }),
  .Z({ S793[53] })
);
BUF_X1 #() 
BUF_X1_594_ (
  .A({ key128[54] }),
  .Z({ S793[54] })
);
BUF_X1 #() 
BUF_X1_595_ (
  .A({ key128[55] }),
  .Z({ S793[55] })
);
BUF_X1 #() 
BUF_X1_596_ (
  .A({ key128[56] }),
  .Z({ S793[56] })
);
BUF_X1 #() 
BUF_X1_597_ (
  .A({ key128[57] }),
  .Z({ S793[57] })
);
BUF_X1 #() 
BUF_X1_598_ (
  .A({ key128[58] }),
  .Z({ S793[58] })
);
BUF_X1 #() 
BUF_X1_599_ (
  .A({ key128[59] }),
  .Z({ S793[59] })
);
BUF_X1 #() 
BUF_X1_600_ (
  .A({ key128[6] }),
  .Z({ S793[6] })
);
BUF_X1 #() 
BUF_X1_601_ (
  .A({ key128[60] }),
  .Z({ S793[60] })
);
BUF_X1 #() 
BUF_X1_602_ (
  .A({ key128[61] }),
  .Z({ S793[61] })
);
BUF_X1 #() 
BUF_X1_603_ (
  .A({ key128[62] }),
  .Z({ S793[62] })
);
BUF_X1 #() 
BUF_X1_604_ (
  .A({ key128[63] }),
  .Z({ S793[63] })
);
BUF_X1 #() 
BUF_X1_605_ (
  .A({ key128[64] }),
  .Z({ S793[64] })
);
BUF_X1 #() 
BUF_X1_606_ (
  .A({ key128[65] }),
  .Z({ S793[65] })
);
BUF_X1 #() 
BUF_X1_607_ (
  .A({ key128[66] }),
  .Z({ S793[66] })
);
BUF_X1 #() 
BUF_X1_608_ (
  .A({ key128[67] }),
  .Z({ S793[67] })
);
BUF_X1 #() 
BUF_X1_609_ (
  .A({ key128[68] }),
  .Z({ S793[68] })
);
BUF_X1 #() 
BUF_X1_610_ (
  .A({ key128[69] }),
  .Z({ S793[69] })
);
BUF_X1 #() 
BUF_X1_611_ (
  .A({ key128[7] }),
  .Z({ S793[7] })
);
BUF_X1 #() 
BUF_X1_612_ (
  .A({ key128[70] }),
  .Z({ S793[70] })
);
BUF_X1 #() 
BUF_X1_613_ (
  .A({ key128[71] }),
  .Z({ S793[71] })
);
BUF_X1 #() 
BUF_X1_614_ (
  .A({ key128[72] }),
  .Z({ S793[72] })
);
BUF_X1 #() 
BUF_X1_615_ (
  .A({ key128[73] }),
  .Z({ S793[73] })
);
BUF_X1 #() 
BUF_X1_616_ (
  .A({ key128[74] }),
  .Z({ S793[74] })
);
BUF_X1 #() 
BUF_X1_617_ (
  .A({ key128[75] }),
  .Z({ S793[75] })
);
BUF_X1 #() 
BUF_X1_618_ (
  .A({ key128[76] }),
  .Z({ S793[76] })
);
BUF_X1 #() 
BUF_X1_619_ (
  .A({ key128[77] }),
  .Z({ S793[77] })
);
BUF_X1 #() 
BUF_X1_620_ (
  .A({ key128[78] }),
  .Z({ S793[78] })
);
BUF_X1 #() 
BUF_X1_621_ (
  .A({ key128[79] }),
  .Z({ S793[79] })
);
BUF_X1 #() 
BUF_X1_622_ (
  .A({ key128[8] }),
  .Z({ S793[8] })
);
BUF_X1 #() 
BUF_X1_623_ (
  .A({ key128[80] }),
  .Z({ S793[80] })
);
BUF_X1 #() 
BUF_X1_624_ (
  .A({ key128[81] }),
  .Z({ S793[81] })
);
BUF_X1 #() 
BUF_X1_625_ (
  .A({ key128[82] }),
  .Z({ S793[82] })
);
BUF_X1 #() 
BUF_X1_626_ (
  .A({ key128[83] }),
  .Z({ S793[83] })
);
BUF_X1 #() 
BUF_X1_627_ (
  .A({ key128[84] }),
  .Z({ S793[84] })
);
BUF_X1 #() 
BUF_X1_628_ (
  .A({ key128[85] }),
  .Z({ S793[85] })
);
BUF_X1 #() 
BUF_X1_629_ (
  .A({ key128[86] }),
  .Z({ S793[86] })
);
BUF_X1 #() 
BUF_X1_630_ (
  .A({ key128[87] }),
  .Z({ S793[87] })
);
BUF_X1 #() 
BUF_X1_631_ (
  .A({ key128[88] }),
  .Z({ S793[88] })
);
BUF_X1 #() 
BUF_X1_632_ (
  .A({ key128[89] }),
  .Z({ S793[89] })
);
BUF_X1 #() 
BUF_X1_633_ (
  .A({ key128[9] }),
  .Z({ S793[9] })
);
BUF_X1 #() 
BUF_X1_634_ (
  .A({ key128[90] }),
  .Z({ S793[90] })
);
BUF_X1 #() 
BUF_X1_635_ (
  .A({ key128[91] }),
  .Z({ S793[91] })
);
BUF_X1 #() 
BUF_X1_636_ (
  .A({ key128[92] }),
  .Z({ S793[92] })
);
BUF_X1 #() 
BUF_X1_637_ (
  .A({ key128[93] }),
  .Z({ S793[93] })
);
BUF_X1 #() 
BUF_X1_638_ (
  .A({ key128[94] }),
  .Z({ S793[94] })
);
BUF_X1 #() 
BUF_X1_639_ (
  .A({ key128[95] }),
  .Z({ S793[95] })
);
BUF_X1 #() 
BUF_X1_640_ (
  .A({ key128[96] }),
  .Z({ S793[96] })
);
BUF_X1 #() 
BUF_X1_641_ (
  .A({ key128[97] }),
  .Z({ S793[97] })
);
BUF_X1 #() 
BUF_X1_642_ (
  .A({ key128[98] }),
  .Z({ S793[98] })
);
BUF_X1 #() 
BUF_X1_643_ (
  .A({ key128[99] }),
  .Z({ S793[99] })
);
AES_Encrypt #() 
AES_Encrypt_1_ (
  .in({ S792[0], S792[1], S792[2], S792[3], S792[4], S792[5], S792[6], S792[7], S792[8], S792[9], S792[10], S792[11], S792[12], S792[13], S792[14], S792[15], S792[16], S792[17], S792[18], S792[19], S792[20], S792[21], S792[22], S792[23], S792[24], S792[25], S792[26], S792[27], S792[28], S792[29], S792[30], S792[31], S792[32], S792[33], S792[34], S792[35], S792[36], S792[37], S792[38], S792[39], S792[40], S792[41], S792[42], S792[43], S792[44], S792[45], S792[46], S792[47], S792[48], S792[49], S792[50], S792[51], S792[52], S792[53], S792[54], S792[55], S792[56], S792[57], S792[58], S792[59], S792[60], S792[61], S792[62], S792[63], S792[64], S792[65], S792[66], S792[67], S792[68], S792[69], S792[70], S792[71], S792[72], S792[73], S792[74], S792[75], S792[76], S792[77], S792[78], S792[79], S792[80], S792[81], S792[82], S792[83], S792[84], S792[85], S792[86], S792[87], S792[88], S792[89], S792[90], S792[91], S792[92], S792[93], S792[94], S792[95], S792[96], S792[97], S792[98], S792[99], S792[100], S792[101], S792[102], S792[103], S792[104], S792[105], S792[106], S792[107], S792[108], S792[109], S792[110], S792[111], S792[112], S792[113], S792[114], S792[115], S792[116], S792[117], S792[118], S792[119], S792[120], S792[121], S792[122], S792[123], S792[124], S792[125], S792[126], S792[127] }),
  .key({ S793[0], S793[1], S793[2], S793[3], S793[4], S793[5], S793[6], S793[7], S793[8], S793[9], S793[10], S793[11], S793[12], S793[13], S793[14], S793[15], S793[16], S793[17], S793[18], S793[19], S793[20], S793[21], S793[22], S793[23], S793[24], S793[25], S793[26], S793[27], S793[28], S793[29], S793[30], S793[31], S793[32], S793[33], S793[34], S793[35], S793[36], S793[37], S793[38], S793[39], S793[40], S793[41], S793[42], S793[43], S793[44], S793[45], S793[46], S793[47], S793[48], S793[49], S793[50], S793[51], S793[52], S793[53], S793[54], S793[55], S793[56], S793[57], S793[58], S793[59], S793[60], S793[61], S793[62], S793[63], S793[64], S793[65], S793[66], S793[67], S793[68], S793[69], S793[70], S793[71], S793[72], S793[73], S793[74], S793[75], S793[76], S793[77], S793[78], S793[79], S793[80], S793[81], S793[82], S793[83], S793[84], S793[85], S793[86], S793[87], S793[88], S793[89], S793[90], S793[91], S793[92], S793[93], S793[94], S793[95], S793[96], S793[97], S793[98], S793[99], S793[100], S793[101], S793[102], S793[103], S793[104], S793[105], S793[106], S793[107], S793[108], S793[109], S793[110], S793[111], S793[112], S793[113], S793[114], S793[115], S793[116], S793[117], S793[118], S793[119], S793[120], S793[121], S793[122], S793[123], S793[124], S793[125], S793[126], S793[127] }),
  .out({ S790[0], S790[1], S790[2], S790[3], S790[4], S790[5], S790[6], S790[7], S790[8], S790[9], S790[10], S790[11], S790[12], S790[13], S790[14], S790[15], S790[16], S790[17], S790[18], S790[19], S790[20], S790[21], S790[22], S790[23], S790[24], S790[25], S790[26], S790[27], S790[28], S790[29], S790[30], S790[31], S790[32], S790[33], S790[34], S790[35], S790[36], S790[37], S790[38], S790[39], S790[40], S790[41], S790[42], S790[43], S790[44], S790[45], S790[46], S790[47], S790[48], S790[49], S790[50], S790[51], S790[52], S790[53], S790[54], S790[55], S790[56], S790[57], S790[58], S790[59], S790[60], S790[61], S790[62], S790[63], S790[64], S790[65], S790[66], S790[67], S790[68], S790[69], S790[70], S790[71], S790[72], S790[73], S790[74], S790[75], S790[76], S790[77], S790[78], S790[79], S790[80], S790[81], S790[82], S790[83], S790[84], S790[85], S790[86], S790[87], S790[88], S790[89], S790[90], S790[91], S790[92], S790[93], S790[94], S790[95], S790[96], S790[97], S790[98], S790[99], S790[100], S790[101], S790[102], S790[103], S790[104], S790[105], S790[106], S790[107], S790[108], S790[109], S790[110], S790[111], S790[112], S790[113], S790[114], S790[115], S790[116], S790[117], S790[118], S790[119], S790[120], S790[121], S790[122], S790[123], S790[124], S790[125], S790[126], S790[127] })
);
AES_Decrypt #() 
AES_Decrypt_1_ (
  .in({ S790[0], S790[1], S790[2], S790[3], S790[4], S790[5], S790[6], S790[7], S790[8], S790[9], S790[10], S790[11], S790[12], S790[13], S790[14], S790[15], S790[16], S790[17], S790[18], S790[19], S790[20], S790[21], S790[22], S790[23], S790[24], S790[25], S790[26], S790[27], S790[28], S790[29], S790[30], S790[31], S790[32], S790[33], S790[34], S790[35], S790[36], S790[37], S790[38], S790[39], S790[40], S790[41], S790[42], S790[43], S790[44], S790[45], S790[46], S790[47], S790[48], S790[49], S790[50], S790[51], S790[52], S790[53], S790[54], S790[55], S790[56], S790[57], S790[58], S790[59], S790[60], S790[61], S790[62], S790[63], S790[64], S790[65], S790[66], S790[67], S790[68], S790[69], S790[70], S790[71], S790[72], S790[73], S790[74], S790[75], S790[76], S790[77], S790[78], S790[79], S790[80], S790[81], S790[82], S790[83], S790[84], S790[85], S790[86], S790[87], S790[88], S790[89], S790[90], S790[91], S790[92], S790[93], S790[94], S790[95], S790[96], S790[97], S790[98], S790[99], S790[100], S790[101], S790[102], S790[103], S790[104], S790[105], S790[106], S790[107], S790[108], S790[109], S790[110], S790[111], S790[112], S790[113], S790[114], S790[115], S790[116], S790[117], S790[118], S790[119], S790[120], S790[121], S790[122], S790[123], S790[124], S790[125], S790[126], S790[127] }),
  .key({ S793[0], S793[1], S793[2], S793[3], S793[4], S793[5], S793[6], S793[7], S793[8], S793[9], S793[10], S793[11], S793[12], S793[13], S793[14], S793[15], S793[16], S793[17], S793[18], S793[19], S793[20], S793[21], S793[22], S793[23], S793[24], S793[25], S793[26], S793[27], S793[28], S793[29], S793[30], S793[31], S793[32], S793[33], S793[34], S793[35], S793[36], S793[37], S793[38], S793[39], S793[40], S793[41], S793[42], S793[43], S793[44], S793[45], S793[46], S793[47], S793[48], S793[49], S793[50], S793[51], S793[52], S793[53], S793[54], S793[55], S793[56], S793[57], S793[58], S793[59], S793[60], S793[61], S793[62], S793[63], S793[64], S793[65], S793[66], S793[67], S793[68], S793[69], S793[70], S793[71], S793[72], S793[73], S793[74], S793[75], S793[76], S793[77], S793[78], S793[79], S793[80], S793[81], S793[82], S793[83], S793[84], S793[85], S793[86], S793[87], S793[88], S793[89], S793[90], S793[91], S793[92], S793[93], S793[94], S793[95], S793[96], S793[97], S793[98], S793[99], S793[100], S793[101], S793[102], S793[103], S793[104], S793[105], S793[106], S793[107], S793[108], S793[109], S793[110], S793[111], S793[112], S793[113], S793[114], S793[115], S793[116], S793[117], S793[118], S793[119], S793[120], S793[121], S793[122], S793[123], S793[124], S793[125], S793[126], S793[127] }),
  .out({ S787[0], S787[1], S787[2], S787[3], S787[4], S787[5], S787[6], S787[7], S787[8], S787[9], S787[10], S787[11], S787[12], S787[13], S787[14], S787[15], S787[16], S787[17], S787[18], S787[19], S787[20], S787[21], S787[22], S787[23], S787[24], S787[25], S787[26], S787[27], S787[28], S787[29], S787[30], S787[31], S787[32], S787[33], S787[34], S787[35], S787[36], S787[37], S787[38], S787[39], S787[40], S787[41], S787[42], S787[43], S787[44], S787[45], S787[46], S787[47], S787[48], S787[49], S787[50], S787[51], S787[52], S787[53], S787[54], S787[55], S787[56], S787[57], S787[58], S787[59], S787[60], S787[61], S787[62], S787[63], S787[64], S787[65], S787[66], S787[67], S787[68], S787[69], S787[70], S787[71], S787[72], S787[73], S787[74], S787[75], S787[76], S787[77], S787[78], S787[79], S787[80], S787[81], S787[82], S787[83], S787[84], S787[85], S787[86], S787[87], S787[88], S787[89], S787[90], S787[91], S787[92], S787[93], S787[94], S787[95], S787[96], S787[97], S787[98], S787[99], S787[100], S787[101], S787[102], S787[103], S787[104], S787[105], S787[106], S787[107], S787[108], S787[109], S787[110], S787[111], S787[112], S787[113], S787[114], S787[115], S787[116], S787[117], S787[118], S787[119], S787[120], S787[121], S787[122], S787[123], S787[124], S787[125], S787[126], S787[127] })
);

endmodule