module c432(N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, N421, N430, N431, N432);

wire _0_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _10_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _11_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _12_;
wire _130_;
wire _131_;
wire _13_;
wire _14_;
wire _15_;
wire _16_;
wire _17_;
wire _18_;
wire _19_;
wire _1_;
wire _20_;
wire _21_;
wire _22_;
wire _23_;
wire _24_;
wire _25_;
wire _26_;
wire _27_;
wire _28_;
wire _29_;
wire _2_;
wire _30_;
wire _31_;
wire _32_;
wire _33_;
wire _34_;
wire _35_;
wire _36_;
wire _37_;
wire _38_;
wire _39_;
wire _3_;
wire _40_;
wire _41_;
wire _42_;
wire _43_;
wire _44_;
wire _45_;
wire _46_;
wire _47_;
wire _48_;
wire _49_;
wire _4_;
wire _50_;
wire _51_;
wire _52_;
wire _53_;
wire _54_;
wire _55_;
wire _56_;
wire _57_;
wire _58_;
wire _59_;
wire _5_;
wire _60_;
wire _61_;
wire _62_;
wire _63_;
wire _64_;
wire _65_;
wire _66_;
wire _67_;
wire _68_;
wire _69_;
wire _6_;
wire _70_;
wire _71_;
wire _72_;
wire _73_;
wire _74_;
wire _75_;
wire _76_;
wire _77_;
wire _78_;
wire _79_;
wire _7_;
wire _80_;
wire _81_;
wire _82_;
wire _83_;
wire _84_;
wire _85_;
wire _86_;
wire _87_;
wire _88_;
wire _89_;
wire _8_;
wire _90_;
wire _91_;
wire _92_;
wire _93_;
wire _94_;
wire _95_;
wire _96_;
wire _97_;
wire _98_;
wire _99_;
wire _9_;
input N1;
input N4;
input N8;
input N11;
input N14;
input N17;
input N21;
input N24;
input N27;
input N30;
input N34;
input N37;
input N40;
input N43;
input N47;
input N50;
input N53;
input N56;
input N60;
input N63;
input N66;
input N69;
input N73;
input N76;
input N79;
input N82;
input N86;
input N89;
input N92;
input N95;
input N99;
input N102;
input N105;
input N108;
input N112;
input N115;
output N223;
output N329;
output N370;
output N421;
output N430;
output N431;
output N432;

AND2_X1 #() 
AND2_X1_1_ (
  .A1({ _84_ }),
  .A2({ N108 }),
  .ZN({ _85_ })
);
AND2_X1 #() 
AND2_X1_2_ (
  .A1({ _126_ }),
  .A2({ N8 }),
  .ZN({ _60_ })
);
AND2_X1 #() 
AND2_X1_3_ (
  .A1({ _37_ }),
  .A2({ _40_ }),
  .ZN({ _62_ })
);
AND2_X1 #() 
AND2_X1_4_ (
  .A1({ _44_ }),
  .A2({ _45_ }),
  .ZN({ _67_ })
);
AND4_X1 #() 
AND4_X1_1_ (
  .A1({ _37_ }),
  .A2({ _40_ }),
  .A3({ _43_ }),
  .A4({ _46_ }),
  .ZN({ _47_ })
);
AND4_X1 #() 
AND4_X1_2_ (
  .A1({ _49_ }),
  .A2({ _52_ }),
  .A3({ _55_ }),
  .A4({ _58_ }),
  .ZN({ _59_ })
);
AOI211_X1 #() 
AOI211_X1_1_ (
  .A({ _7_ }),
  .B({ _60_ }),
  .C1({ _127_ }),
  .C2({ N14 }),
  .ZN({ _61_ })
);
AOI21_X1 #() 
AOI21_X1_1_ (
  .A({ _90_ }),
  .B1({ _117_ }),
  .B2({ N112 }),
  .ZN({ _123_ })
);
AOI21_X1 #() 
AOI21_X1_2_ (
  .A({ _31_ }),
  .B1({ _126_ }),
  .B2({ N34 }),
  .ZN({ _36_ })
);
AOI21_X1 #() 
AOI21_X1_3_ (
  .A({ _2_ }),
  .B1({ _126_ }),
  .B2({ N21 }),
  .ZN({ _39_ })
);
AOI21_X1 #() 
AOI21_X1_4_ (
  .A({ _119_ }),
  .B1({ _126_ }),
  .B2({ N60 }),
  .ZN({ _42_ })
);
AOI21_X1 #() 
AOI21_X1_5_ (
  .A({ _27_ }),
  .B1({ _126_ }),
  .B2({ N47 }),
  .ZN({ _45_ })
);
AOI21_X1 #() 
AOI21_X1_6_ (
  .A({ _22_ }),
  .B1({ _126_ }),
  .B2({ N99 }),
  .ZN({ _50_ })
);
AOI21_X1 #() 
AOI21_X1_7_ (
  .A({ _13_ }),
  .B1({ _126_ }),
  .B2({ N86 }),
  .ZN({ _54_ })
);
AOI21_X1 #() 
AOI21_X1_8_ (
  .A({ _18_ }),
  .B1({ _126_ }),
  .B2({ N73 }),
  .ZN({ _56_ })
);
AOI21_X1 #() 
AOI21_X1_9_ (
  .A({ _61_ }),
  .B1({ _47_ }),
  .B2({ _59_ }),
  .ZN({ _128_ })
);
AOI22_X1 #() 
AOI22_X1_1_ (
  .A1({ N56 }),
  .A2({ _71_ }),
  .B1({ _72_ }),
  .B2({ N95 }),
  .ZN({ _73_ })
);
AOI22_X1 #() 
AOI22_X1_2_ (
  .A1({ _26_ }),
  .A2({ _28_ }),
  .B1({ _30_ }),
  .B2({ _32_ }),
  .ZN({ _33_ })
);
AOI22_X1 #() 
AOI22_X1_3_ (
  .A1({ _67_ }),
  .A2({ _37_ }),
  .B1({ _38_ }),
  .B2({ _39_ }),
  .ZN({ _68_ })
);
AOI22_X1 #() 
AOI22_X1_4_ (
  .A1({ _74_ }),
  .A2({ N4 }),
  .B1({ _75_ }),
  .B2({ N43 }),
  .ZN({ _76_ })
);
AOI22_X1 #() 
AOI22_X1_5_ (
  .A1({ N17 }),
  .A2({ _77_ }),
  .B1({ _78_ }),
  .B2({ N30 }),
  .ZN({ _79_ })
);
AOI22_X1 #() 
AOI22_X1_6_ (
  .A1({ N69 }),
  .A2({ _80_ }),
  .B1({ _81_ }),
  .B2({ N82 }),
  .ZN({ _82_ })
);
AOI22_X1 #() 
AOI22_X1_7_ (
  .A1({ _93_ }),
  .A2({ _94_ }),
  .B1({ _97_ }),
  .B2({ _96_ }),
  .ZN({ _98_ })
);
AOI22_X1 #() 
AOI22_X1_8_ (
  .A1({ _100_ }),
  .A2({ _101_ }),
  .B1({ _86_ }),
  .B2({ _70_ }),
  .ZN({ _102_ })
);
AOI22_X1 #() 
AOI22_X1_9_ (
  .A1({ _104_ }),
  .A2({ _105_ }),
  .B1({ _108_ }),
  .B2({ _107_ }),
  .ZN({ _109_ })
);
AOI22_X1 #() 
AOI22_X1_10_ (
  .A1({ _111_ }),
  .A2({ _112_ }),
  .B1({ _115_ }),
  .B2({ _114_ }),
  .ZN({ _116_ })
);
AOI22_X1 #() 
AOI22_X1_11_ (
  .A1({ _17_ }),
  .A2({ _19_ }),
  .B1({ _21_ }),
  .B2({ _23_ }),
  .ZN({ _24_ })
);
BUF_X1 #() 
BUF_X1_1_ (
  .A({ _125_ }),
  .Z({ N223 })
);
BUF_X1 #() 
BUF_X1_2_ (
  .A({ _126_ }),
  .Z({ N329 })
);
BUF_X1 #() 
BUF_X1_3_ (
  .A({ _127_ }),
  .Z({ N370 })
);
BUF_X1 #() 
BUF_X1_4_ (
  .A({ _128_ }),
  .Z({ N421 })
);
BUF_X1 #() 
BUF_X1_5_ (
  .A({ _129_ }),
  .Z({ N430 })
);
BUF_X1 #() 
BUF_X1_6_ (
  .A({ _130_ }),
  .Z({ N431 })
);
BUF_X1 #() 
BUF_X1_7_ (
  .A({ _131_ }),
  .Z({ N432 })
);
INV_X1 #() 
INV_X1_1_ (
  .A({ N56 }),
  .ZN({ _69_ })
);
INV_X1 #() 
INV_X1_2_ (
  .A({ N102 }),
  .ZN({ _84_ })
);
INV_X1 #() 
INV_X1_3_ (
  .A({ _87_ }),
  .ZN({ _88_ })
);
INV_X1 #() 
INV_X1_4_ (
  .A({ N43 }),
  .ZN({ _92_ })
);
INV_X1 #() 
INV_X1_5_ (
  .A({ N82 }),
  .ZN({ _95_ })
);
INV_X1 #() 
INV_X1_6_ (
  .A({ N69 }),
  .ZN({ _99_ })
);
INV_X1 #() 
INV_X1_7_ (
  .A({ N4 }),
  .ZN({ _103_ })
);
INV_X1 #() 
INV_X1_8_ (
  .A({ N17 }),
  .ZN({ _106_ })
);
INV_X1 #() 
INV_X1_9_ (
  .A({ N95 }),
  .ZN({ _110_ })
);
INV_X1 #() 
INV_X1_10_ (
  .A({ N30 }),
  .ZN({ _113_ })
);
INV_X1 #() 
INV_X1_11_ (
  .A({ N115 }),
  .ZN({ _122_ })
);
INV_X1 #() 
INV_X1_12_ (
  .A({ N50 }),
  .ZN({ _71_ })
);
INV_X1 #() 
INV_X1_13_ (
  .A({ _0_ }),
  .ZN({ _1_ })
);
INV_X1 #() 
INV_X1_14_ (
  .A({ _5_ }),
  .ZN({ _6_ })
);
INV_X1 #() 
INV_X1_15_ (
  .A({ _11_ }),
  .ZN({ _12_ })
);
INV_X1 #() 
INV_X1_16_ (
  .A({ _118_ }),
  .ZN({ _126_ })
);
INV_X1 #() 
INV_X1_17_ (
  .A({ _47_ }),
  .ZN({ _129_ })
);
INV_X1 #() 
INV_X1_18_ (
  .A({ _58_ }),
  .ZN({ _64_ })
);
INV_X1 #() 
INV_X1_19_ (
  .A({ _89_ }),
  .ZN({ _125_ })
);
INV_X1 #() 
INV_X1_20_ (
  .A({ N89 }),
  .ZN({ _72_ })
);
INV_X1 #() 
INV_X1_21_ (
  .A({ N1 }),
  .ZN({ _74_ })
);
INV_X1 #() 
INV_X1_22_ (
  .A({ N37 }),
  .ZN({ _75_ })
);
INV_X1 #() 
INV_X1_23_ (
  .A({ N11 }),
  .ZN({ _77_ })
);
INV_X1 #() 
INV_X1_24_ (
  .A({ N24 }),
  .ZN({ _78_ })
);
INV_X1 #() 
INV_X1_25_ (
  .A({ N63 }),
  .ZN({ _80_ })
);
INV_X1 #() 
INV_X1_26_ (
  .A({ N76 }),
  .ZN({ _81_ })
);
NAND2_X1 #() 
NAND2_X1_1_ (
  .A1({ _86_ }),
  .A2({ _70_ }),
  .ZN({ _87_ })
);
NAND2_X1 #() 
NAND2_X1_2_ (
  .A1({ _101_ }),
  .A2({ _100_ }),
  .ZN({ _16_ })
);
NAND2_X1 #() 
NAND2_X1_3_ (
  .A1({ _101_ }),
  .A2({ N69 }),
  .ZN({ _18_ })
);
NAND2_X1 #() 
NAND2_X1_4_ (
  .A1({ _112_ }),
  .A2({ _111_ }),
  .ZN({ _20_ })
);
NAND2_X1 #() 
NAND2_X1_5_ (
  .A1({ _112_ }),
  .A2({ N95 }),
  .ZN({ _22_ })
);
NAND2_X1 #() 
NAND2_X1_6_ (
  .A1({ _94_ }),
  .A2({ _93_ }),
  .ZN({ _25_ })
);
NAND2_X1 #() 
NAND2_X1_7_ (
  .A1({ _94_ }),
  .A2({ N43 }),
  .ZN({ _27_ })
);
NAND2_X1 #() 
NAND2_X1_8_ (
  .A1({ _115_ }),
  .A2({ _114_ }),
  .ZN({ _29_ })
);
NAND2_X1 #() 
NAND2_X1_9_ (
  .A1({ _115_ }),
  .A2({ N30 }),
  .ZN({ _31_ })
);
NAND2_X1 #() 
NAND2_X1_10_ (
  .A1({ _35_ }),
  .A2({ _36_ }),
  .ZN({ _37_ })
);
NAND2_X1 #() 
NAND2_X1_11_ (
  .A1({ _38_ }),
  .A2({ _39_ }),
  .ZN({ _40_ })
);
NAND2_X1 #() 
NAND2_X1_12_ (
  .A1({ _86_ }),
  .A2({ N56 }),
  .ZN({ _119_ })
);
NAND2_X1 #() 
NAND2_X1_13_ (
  .A1({ _41_ }),
  .A2({ _42_ }),
  .ZN({ _43_ })
);
NAND2_X1 #() 
NAND2_X1_14_ (
  .A1({ _44_ }),
  .A2({ _45_ }),
  .ZN({ _46_ })
);
NAND2_X1 #() 
NAND2_X1_15_ (
  .A1({ _48_ }),
  .A2({ _123_ }),
  .ZN({ _49_ })
);
NAND2_X1 #() 
NAND2_X1_16_ (
  .A1({ _51_ }),
  .A2({ _50_ }),
  .ZN({ _52_ })
);
NAND2_X1 #() 
NAND2_X1_17_ (
  .A1({ _53_ }),
  .A2({ _54_ }),
  .ZN({ _55_ })
);
NAND2_X1 #() 
NAND2_X1_18_ (
  .A1({ _57_ }),
  .A2({ _56_ }),
  .ZN({ _58_ })
);
NAND2_X1 #() 
NAND2_X1_19_ (
  .A1({ _43_ }),
  .A2({ _46_ }),
  .ZN({ _63_ })
);
NAND2_X1 #() 
NAND2_X1_20_ (
  .A1({ _123_ }),
  .A2({ _122_ }),
  .ZN({ _124_ })
);
NAND2_X1 #() 
NAND2_X1_21_ (
  .A1({ _108_ }),
  .A2({ _107_ }),
  .ZN({ _0_ })
);
NAND2_X1 #() 
NAND2_X1_22_ (
  .A1({ _108_ }),
  .A2({ N17 }),
  .ZN({ _2_ })
);
NAND2_X1 #() 
NAND2_X1_23_ (
  .A1({ _105_ }),
  .A2({ _104_ }),
  .ZN({ _5_ })
);
NAND2_X1 #() 
NAND2_X1_24_ (
  .A1({ _105_ }),
  .A2({ N4 }),
  .ZN({ _7_ })
);
NAND2_X1 #() 
NAND2_X1_25_ (
  .A1({ _97_ }),
  .A2({ _96_ }),
  .ZN({ _11_ })
);
NAND2_X1 #() 
NAND2_X1_26_ (
  .A1({ _97_ }),
  .A2({ N82 }),
  .ZN({ _13_ })
);
NAND3_X1 #() 
NAND3_X1_1_ (
  .A1({ _24_ }),
  .A2({ _33_ }),
  .A3({ _15_ }),
  .ZN({ _34_ })
);
NAND3_X1 #() 
NAND3_X1_2_ (
  .A1({ _37_ }),
  .A2({ _46_ }),
  .A3({ _55_ }),
  .ZN({ _66_ })
);
NAND4_X1 #() 
NAND4_X1_1_ (
  .A1({ _73_ }),
  .A2({ _76_ }),
  .A3({ _79_ }),
  .A4({ _82_ }),
  .ZN({ _83_ })
);
NAND4_X1 #() 
NAND4_X1_2_ (
  .A1({ _98_ }),
  .A2({ _102_ }),
  .A3({ _109_ }),
  .A4({ _116_ }),
  .ZN({ _117_ })
);
NAND4_X1 #() 
NAND4_X1_3_ (
  .A1({ _121_ }),
  .A2({ _4_ }),
  .A3({ _9_ }),
  .A4({ _124_ }),
  .ZN({ _10_ })
);
NAND4_X1 #() 
NAND4_X1_4_ (
  .A1({ _64_ }),
  .A2({ _37_ }),
  .A3({ _43_ }),
  .A4({ _46_ }),
  .ZN({ _65_ })
);
NOR2_X1 #() 
NOR2_X1_1_ (
  .A1({ _69_ }),
  .A2({ N60 }),
  .ZN({ _70_ })
);
NOR2_X1 #() 
NOR2_X1_2_ (
  .A1({ _113_ }),
  .A2({ N34 }),
  .ZN({ _114_ })
);
NOR2_X1 #() 
NOR2_X1_3_ (
  .A1({ _117_ }),
  .A2({ _91_ }),
  .ZN({ _118_ })
);
NOR2_X1 #() 
NOR2_X1_4_ (
  .A1({ _119_ }),
  .A2({ N66 }),
  .ZN({ _120_ })
);
NOR2_X1 #() 
NOR2_X1_5_ (
  .A1({ _2_ }),
  .A2({ N27 }),
  .ZN({ _3_ })
);
NOR2_X1 #() 
NOR2_X1_6_ (
  .A1({ _7_ }),
  .A2({ N14 }),
  .ZN({ _8_ })
);
NOR2_X1 #() 
NOR2_X1_7_ (
  .A1({ _13_ }),
  .A2({ N92 }),
  .ZN({ _14_ })
);
NOR2_X1 #() 
NOR2_X1_8_ (
  .A1({ _18_ }),
  .A2({ N79 }),
  .ZN({ _19_ })
);
NOR2_X1 #() 
NOR2_X1_9_ (
  .A1({ _22_ }),
  .A2({ N105 }),
  .ZN({ _23_ })
);
NOR2_X1 #() 
NOR2_X1_10_ (
  .A1({ _27_ }),
  .A2({ N53 }),
  .ZN({ _28_ })
);
NOR2_X1 #() 
NOR2_X1_11_ (
  .A1({ _31_ }),
  .A2({ N40 }),
  .ZN({ _32_ })
);
NOR2_X1 #() 
NOR2_X1_12_ (
  .A1({ _83_ }),
  .A2({ _85_ }),
  .ZN({ _89_ })
);
NOR2_X1 #() 
NOR2_X1_13_ (
  .A1({ _90_ }),
  .A2({ N112 }),
  .ZN({ _91_ })
);
NOR2_X1 #() 
NOR2_X1_14_ (
  .A1({ _92_ }),
  .A2({ N47 }),
  .ZN({ _93_ })
);
NOR2_X1 #() 
NOR2_X1_15_ (
  .A1({ _95_ }),
  .A2({ N86 }),
  .ZN({ _96_ })
);
NOR2_X1 #() 
NOR2_X1_16_ (
  .A1({ _99_ }),
  .A2({ N73 }),
  .ZN({ _100_ })
);
NOR2_X1 #() 
NOR2_X1_17_ (
  .A1({ _103_ }),
  .A2({ N8 }),
  .ZN({ _104_ })
);
NOR2_X1 #() 
NOR2_X1_18_ (
  .A1({ _106_ }),
  .A2({ N21 }),
  .ZN({ _107_ })
);
NOR2_X1 #() 
NOR2_X1_19_ (
  .A1({ _110_ }),
  .A2({ N99 }),
  .ZN({ _111_ })
);
OAI211_X1 #() 
OAI211_X1_1_ (
  .A({ _65_ }),
  .B({ _62_ }),
  .C1({ _63_ }),
  .C2({ _55_ }),
  .ZN({ _130_ })
);
OAI211_X1 #() 
OAI211_X1_2_ (
  .A({ _65_ }),
  .B({ _68_ }),
  .C1({ _52_ }),
  .C2({ _66_ }),
  .ZN({ _131_ })
);
OAI21_X1 #() 
OAI21_X1_1_ (
  .A({ N50 }),
  .B1({ _83_ }),
  .B2({ _85_ }),
  .ZN({ _86_ })
);
OAI21_X1 #() 
OAI21_X1_2_ (
  .A({ _120_ }),
  .B1({ _118_ }),
  .B2({ _88_ }),
  .ZN({ _121_ })
);
OAI21_X1 #() 
OAI21_X1_3_ (
  .A({ _3_ }),
  .B1({ _118_ }),
  .B2({ _1_ }),
  .ZN({ _4_ })
);
OAI21_X1 #() 
OAI21_X1_4_ (
  .A({ _8_ }),
  .B1({ _118_ }),
  .B2({ _6_ }),
  .ZN({ _9_ })
);
OAI21_X1 #() 
OAI21_X1_5_ (
  .A({ _14_ }),
  .B1({ _118_ }),
  .B2({ _12_ }),
  .ZN({ _15_ })
);
OAI21_X1 #() 
OAI21_X1_6_ (
  .A({ _16_ }),
  .B1({ _117_ }),
  .B2({ _91_ }),
  .ZN({ _17_ })
);
OAI21_X1 #() 
OAI21_X1_7_ (
  .A({ _20_ }),
  .B1({ _117_ }),
  .B2({ _91_ }),
  .ZN({ _21_ })
);
OAI21_X1 #() 
OAI21_X1_8_ (
  .A({ _25_ }),
  .B1({ _117_ }),
  .B2({ _91_ }),
  .ZN({ _26_ })
);
OAI21_X1 #() 
OAI21_X1_9_ (
  .A({ _29_ }),
  .B1({ _117_ }),
  .B2({ _91_ }),
  .ZN({ _30_ })
);
OAI21_X1 #() 
OAI21_X1_10_ (
  .A({ N40 }),
  .B1({ _34_ }),
  .B2({ _10_ }),
  .ZN({ _35_ })
);
OAI21_X1 #() 
OAI21_X1_11_ (
  .A({ N27 }),
  .B1({ _34_ }),
  .B2({ _10_ }),
  .ZN({ _38_ })
);
OAI21_X1 #() 
OAI21_X1_12_ (
  .A({ N108 }),
  .B1({ _89_ }),
  .B2({ _84_ }),
  .ZN({ _90_ })
);
OAI21_X1 #() 
OAI21_X1_13_ (
  .A({ N66 }),
  .B1({ _34_ }),
  .B2({ _10_ }),
  .ZN({ _41_ })
);
OAI21_X1 #() 
OAI21_X1_14_ (
  .A({ N53 }),
  .B1({ _34_ }),
  .B2({ _10_ }),
  .ZN({ _44_ })
);
OAI21_X1 #() 
OAI21_X1_15_ (
  .A({ N115 }),
  .B1({ _34_ }),
  .B2({ _10_ }),
  .ZN({ _48_ })
);
OAI21_X1 #() 
OAI21_X1_16_ (
  .A({ N105 }),
  .B1({ _34_ }),
  .B2({ _10_ }),
  .ZN({ _51_ })
);
OAI21_X1 #() 
OAI21_X1_17_ (
  .A({ N92 }),
  .B1({ _34_ }),
  .B2({ _10_ }),
  .ZN({ _53_ })
);
OAI21_X1 #() 
OAI21_X1_18_ (
  .A({ N79 }),
  .B1({ _34_ }),
  .B2({ _10_ }),
  .ZN({ _57_ })
);
OAI21_X1 #() 
OAI21_X1_19_ (
  .A({ N37 }),
  .B1({ _83_ }),
  .B2({ _85_ }),
  .ZN({ _94_ })
);
OAI21_X1 #() 
OAI21_X1_20_ (
  .A({ N76 }),
  .B1({ _83_ }),
  .B2({ _85_ }),
  .ZN({ _97_ })
);
OAI21_X1 #() 
OAI21_X1_21_ (
  .A({ N63 }),
  .B1({ _83_ }),
  .B2({ _85_ }),
  .ZN({ _101_ })
);
OAI21_X1 #() 
OAI21_X1_22_ (
  .A({ N1 }),
  .B1({ _83_ }),
  .B2({ _85_ }),
  .ZN({ _105_ })
);
OAI21_X1 #() 
OAI21_X1_23_ (
  .A({ N11 }),
  .B1({ _83_ }),
  .B2({ _85_ }),
  .ZN({ _108_ })
);
OAI21_X1 #() 
OAI21_X1_24_ (
  .A({ N89 }),
  .B1({ _83_ }),
  .B2({ _85_ }),
  .ZN({ _112_ })
);
OAI21_X1 #() 
OAI21_X1_25_ (
  .A({ N24 }),
  .B1({ _83_ }),
  .B2({ _85_ }),
  .ZN({ _115_ })
);
OR2_X1 #() 
OR2_X1_1_ (
  .A1({ _34_ }),
  .A2({ _10_ }),
  .ZN({ _127_ })
);

endmodule