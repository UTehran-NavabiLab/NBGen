module TopLevel(clk, rst, writeMEM, readMEM, dataBus, addrBus);

wire S0;
wire S1;
wire S2;
wire S3;
wire S4;
wire S5;
wire S6;
wire S7;
wire S8;
wire S9;
wire S10;
wire S11;
wire S12;
wire S13;
wire S14;
wire S15;
wire S16;
wire S17;
wire S18;
wire S19;
wire S20;
wire S21;
wire S22;
wire S23;
wire S24;
wire S25;
wire S26;
wire S27;
wire S28;
wire S29;
wire S30;
wire S31;
wire S32;
wire S33;
wire S34;
wire S35;
wire S36;
wire S37;
wire S38;
wire S39;
wire S40;
wire S41;
wire S42;
wire S43;
wire S44;
wire S45;
wire S46;
wire S47;
wire S48;
wire S49;
wire S50;
wire S51;
wire S52;
wire S53;
wire S54;
wire S55;
wire S56;
wire S57;
wire S58;
wire S59;
wire S60;
wire S61;
wire S62;
wire S63;
wire S64;
wire S65;
wire S66;
wire S67;
wire S68;
wire S69;
wire S70;
wire S71;
wire S72;
wire S73;
wire S74;
wire S75;
wire S76;
wire S77;
wire S78;
wire S79;
wire S80;
wire S81;
wire S82;
wire S83;
wire S84;
wire S85;
wire S86;
wire S87;
wire S88;
wire S89;
wire S90;
wire S91;
wire S92;
wire S93;
wire S94;
wire S95;
wire S96;
wire S97;
wire S98;
wire S99;
wire S100;
wire S101;
wire S102;
wire S103;
wire S104;
wire S105;
wire S106;
wire S107;
wire S108;
wire S109;
wire S110;
wire S111;
wire S112;
wire S113;
wire S114;
wire S115;
wire S116;
wire S117;
wire S118;
wire S119;
wire S120;
wire S121;
wire S122;
wire S123;
wire S124;
wire S125;
wire S126;
wire S127;
wire S128;
wire S129;
wire S130;
wire S131;
wire S132;
wire S133;
wire S134;
wire S135;
wire S136;
wire S137;
wire S138;
wire S139;
wire S140;
wire S141;
wire S142;
wire S143;
wire S144;
wire S145;
wire S146;
wire S147;
wire S148;
wire S149;
wire S150;
wire S151;
wire S152;
wire S153;
wire S154;
wire S155;
wire S156;
wire S157;
wire S158;
wire S159;
wire S160;
wire S161;
wire S162;
wire S163;
wire S164;
wire S165;
wire S166;
wire S167;
wire S168;
wire S169;
wire S170;
wire S171;
wire S172;
wire S173;
wire S174;
wire S175;
wire S176;
wire S177;
wire S178;
wire S179;
wire S180;
wire S181;
wire S182;
wire S183;
wire S184;
wire S185;
wire S186;
wire S187;
wire S188;
wire S189;
wire S190;
wire S191;
wire S192;
wire S193;
wire S194;
wire S195;
wire S196;
wire S197;
wire S198;
wire S199;
wire S200;
wire S201;
wire S202;
wire S203;
wire S204;
wire S205;
wire S206;
wire S207;
wire S208;
wire S209;
wire S210;
wire S211;
wire S212;
wire S213;
wire S214;
wire S215;
wire S216;
wire S217;
wire S218;
wire S219;
wire S220;
wire S221;
wire S222;
wire S223;
wire S224;
wire S225;
wire S226;
wire S227;
wire S228;
wire S229;
wire S230;
wire S231;
wire S232;
wire S233;
wire S234;
wire S235;
wire S236;
wire S237;
wire S238;
wire S239;
wire S240;
wire S241;
wire S242;
wire S243;
wire S244;
wire S245;
wire S246;
wire S247;
wire S248;
wire S249;
wire S250;
wire S251;
wire S252;
wire S253;
wire S254;
wire S255;
wire S256;
wire S257;
wire S258;
wire S259;
wire S260;
wire S261;
wire S262;
wire S263;
wire S264;
wire S265;
wire S266;
wire S267;
wire S268;
wire S269;
wire S270;
wire S271;
wire S272;
wire S273;
wire S274;
wire S275;
wire S276;
wire S277;
wire S278;
wire S279;
wire S280;
wire S281;
wire S282;
wire S283;
wire S284;
wire S285;
wire S286;
wire S287;
wire S288;
wire S289;
wire S290;
wire S291;
wire S292;
wire S293;
wire S294;
wire S295;
wire S296;
wire S297;
wire S298;
wire S299;
wire S300;
wire S301;
wire S302;
wire S303;
wire S304;
wire S305;
wire S306;
wire S307;
wire S308;
wire S309;
wire S310;
wire S311;
wire S312;
wire S313;
wire S314;
wire S315;
wire S316;
wire S317;
wire S318;
wire S319;
wire S320;
wire S321;
wire S322;
wire S323;
wire S324;
wire S325;
wire S326;
wire S327;
wire S328;
wire S329;
wire S330;
wire S331;
wire S332;
wire S333;
wire S334;
wire S335;
wire S336;
wire S337;
wire S338;
wire S339;
wire S340;
wire S341;
wire S342;
wire S343;
wire S344;
wire S345;
wire S346;
wire S347;
wire S348;
wire S349;
wire S350;
wire S351;
wire S352;
wire S353;
wire S354;
wire S355;
wire S356;
wire S357;
wire S358;
wire S359;
wire S360;
wire S361;
wire S362;
wire S363;
wire S364;
wire S365;
wire S366;
wire S367;
wire S368;
wire S369;
wire S370;
wire S371;
wire S372;
wire S373;
wire S374;
wire S375;
wire S376;
wire S377;
wire S378;
wire S379;
wire S380;
wire S381;
wire S382;
wire S383;
wire S384;
wire S385;
wire S386;
wire S387;
wire S388;
wire S389;
wire S390;
wire S391;
wire S392;
wire S393;
wire S394;
wire S395;
wire S396;
wire S397;
wire S398;
wire S399;
wire S400;
wire S401;
wire S402;
wire S403;
wire S404;
wire S405;
wire S406;
wire S407;
wire S408;
wire S409;
wire S410;
wire S411;
wire S412;
wire S413;
wire S414;
wire S415;
wire S416;
wire S417;
wire S418;
wire S419;
wire S420;
wire S421;
wire S422;
wire S423;
wire S424;
wire S425;
wire S426;
wire S427;
wire S428;
wire S429;
wire S430;
wire S431;
wire S432;
wire S433;
wire S434;
wire S435;
wire S436;
wire S437;
wire S438;
wire S439;
wire S440;
wire S441;
wire S442;
wire S443;
wire S444;
wire S445;
wire S446;
wire S447;
wire S448;
wire S449;
wire S450;
wire S451;
wire S452;
wire S453;
wire S454;
wire S455;
wire S456;
wire S457;
wire S458;
wire S459;
wire S460;
wire S461;
wire S462;
wire S463;
wire S464;
wire S465;
wire S466;
wire S467;
wire S468;
wire S469;
wire S470;
wire S471;
wire S472;
wire S473;
wire S474;
wire S475;
wire S476;
wire S477;
wire S478;
wire S479;
wire S480;
wire S481;
wire S482;
wire S483;
wire S484;
wire S485;
wire S486;
wire S487;
wire S488;
wire S489;
wire S490;
wire S491;
wire S492;
wire S493;
wire S494;
wire S495;
wire S496;
wire S497;
wire S498;
wire S499;
wire S500;
wire S501;
wire S502;
wire S503;
wire S504;
wire S505;
wire S506;
wire S507;
wire S508;
wire S509;
wire S510;
wire S511;
wire S512;
wire S513;
wire S514;
wire S515;
wire S516;
wire S517;
wire S518;
wire S519;
wire S520;
wire S521;
wire S522;
wire S523;
wire S524;
wire S525;
wire S526;
wire S527;
wire S528;
wire S529;
wire S530;
wire S531;
wire S532;
wire S533;
wire S534;
wire S535;
wire S536;
wire S537;
wire S538;
wire S539;
wire S540;
wire S541;
wire S542;
wire S543;
wire S544;
wire S545;
wire S546;
wire S547;
wire S548;
wire S549;
wire S550;
wire S551;
wire S552;
wire S553;
wire S554;
wire S555;
wire S556;
wire S557;
wire S558;
wire S559;
wire S560;
wire S561;
wire S562;
wire S563;
wire S564;
wire S565;
wire S566;
wire S567;
wire S568;
wire S569;
wire S570;
wire S571;
wire S572;
wire S573;
wire S574;
wire S575;
wire S576;
wire S577;
wire S578;
wire S579;
wire S580;
wire S581;
wire S582;
wire S583;
wire S584;
wire S585;
wire S586;
wire S587;
wire S588;
wire S589;
wire S590;
wire S591;
wire S592;
wire S593;
wire S594;
wire S595;
wire S596;
wire S597;
wire S598;
wire S599;
wire S600;
wire S601;
wire S602;
wire S603;
wire S604;
wire S605;
wire S606;
wire S607;
wire S608;
wire S609;
wire S610;
wire S611;
wire S612;
wire S613;
wire S614;
wire S615;
wire S616;
wire S617;
wire S618;
wire S619;
wire S620;
wire S621;
wire S622;
wire S623;
wire S624;
wire S625;
wire S626;
wire S627;
wire S628;
wire S629;
wire S630;
wire S631;
wire S632;
wire S633;
wire S634;
wire S635;
wire S636;
wire S637;
wire S638;
wire S639;
wire S640;
wire S641;
wire S642;
wire S643;
wire S644;
wire S645;
wire S646;
wire S647;
wire S648;
wire S649;
wire S650;
wire S651;
wire S652;
wire S653;
wire S654;
wire S655;
wire S656;
wire S657;
wire S658;
wire S659;
wire S660;
wire S661;
wire S662;
wire S663;
wire S664;
wire S665;
wire S666;
wire S667;
wire S668;
wire S669;
wire S670;
wire S671;
wire S672;
wire S673;
wire S674;
wire S675;
wire S676;
wire S677;
wire S678;
wire S679;
wire S680;
wire S681;
wire S682;
wire S683;
wire S684;
wire S685;
wire S686;
wire S687;
wire S688;
wire S689;
wire S690;
wire S691;
wire S692;
wire S693;
wire S694;
wire S695;
wire S696;
wire S697;
wire S698;
wire S699;
wire S700;
wire S701;
wire S702;
wire S703;
wire S704;
wire S705;
wire S706;
wire S707;
wire S708;
wire S709;
wire S710;
wire S711;
wire S712;
wire S713;
wire S714;
wire S715;
wire S716;
wire S717;
wire S718;
wire S719;
wire S720;
wire S721;
wire S722;
wire S723;
wire S724;
wire S725;
wire S726;
wire S727;
wire S728;
wire S729;
wire S730;
wire S731;
wire S732;
wire S733;
wire S734;
wire S735;
wire S736;
wire S737;
wire S738;
wire S739;
wire S740;
wire S741;
wire S742;
wire S743;
wire S744;
wire S745;
wire S746;
wire S747;
wire S748;
wire S749;
wire S750;
wire S751;
wire S752;
wire S753;
wire S754;
wire S755;
wire S756;
wire S757;
wire S758;
wire S759;
wire S760;
wire S761;
wire S762;
wire S763;
wire S764;
wire S765;
wire S766;
wire S767;
wire S768;
wire S769;
wire S770;
wire S771;
wire S772;
wire S773;
wire S774;
wire S775;
wire S776;
wire S777;
wire S778;
wire S779;
wire S780;
wire S781;
wire S782;
wire S783;
wire S784;
wire S785;
wire S786;
wire S787;
wire S788;
wire S789;
wire S790;
wire S791;
wire S792;
wire S793;
wire S794;
wire S795;
wire S796;
wire S797;
wire S798;
wire S799;
wire S800;
wire S801;
wire S802;
wire S803;
wire S804;
wire S805;
wire S806;
wire S807;
wire S808;
wire S809;
wire S810;
wire S811;
wire S812;
wire S813;
wire S814;
wire S815;
wire S816;
wire S817;
wire S818;
wire S819;
wire S820;
wire S821;
wire S822;
wire S823;
wire S824;
wire S825;
wire S826;
wire S827;
wire S828;
wire S829;
wire S830;
wire S831;
wire S832;
wire S833;
wire S834;
wire S835;
wire S836;
wire S837;
wire S838;
wire S839;
wire S840;
wire S841;
wire S842;
wire S843;
wire S844;
wire S845;
wire S846;
wire S847;
wire S848;
wire S849;
wire S850;
wire S851;
wire S852;
wire S853;
wire S854;
wire S855;
wire S856;
wire S857;
wire S858;
wire S859;
wire S860;
wire S861;
wire S862;
wire S863;
wire S864;
wire S865;
wire S866;
wire S867;
wire S868;
wire S869;
wire S870;
wire S871;
wire S872;
wire S873;
wire S874;
wire S875;
wire S876;
wire S877;
wire S878;
wire S879;
wire S880;
wire S881;
wire S882;
wire S883;
wire S884;
wire S885;
wire S886;
wire S887;
wire S888;
wire S889;
wire S890;
wire S891;
wire S892;
wire S893;
wire S894;
wire S895;
wire S896;
wire S897;
wire S898;
wire S899;
wire S900;
wire S901;
wire S902;
wire S903;
wire S904;
wire S905;
wire S906;
wire S907;
wire S908;
wire S909;
wire S910;
wire S911;
wire S912;
wire S913;
wire S914;
wire S915;
wire S916;
wire S917;
wire S918;
wire S919;
wire S920;
wire S921;
wire S922;
wire S923;
wire S924;
wire S925;
wire S926;
wire S927;
wire S928;
wire S929;
wire S930;
wire S931;
wire S932;
wire S933;
wire S934;
wire S935;
wire S936;
wire S937;
wire S938;
wire S939;
wire S940;
wire S941;
wire S942;
wire S943;
wire S944;
wire S945;
wire S946;
wire S947;
wire S948;
wire S949;
wire S950;
wire S951;
wire S952;
wire S953;
wire S954;
wire S955;
wire S956;
wire S957;
wire S958;
wire S959;
wire S960;
wire S961;
wire S962;
wire S963;
wire S964;
wire S965;
wire S966;
wire S967;
wire S968;
wire S969;
wire S970;
wire S971;
wire S972;
wire S973;
wire S974;
wire S975;
wire S976;
wire S977;
wire S978;
wire S979;
wire S980;
wire S981;
wire S982;
wire S983;
wire S984;
wire S985;
wire S986;
wire S987;
wire S988;
wire S989;
wire S990;
wire S991;
wire S992;
wire S993;
wire S994;
wire S995;
wire S996;
wire S997;
wire S998;
wire S999;
wire S1000;
wire S1001;
wire S1002;
wire S1003;
wire S1004;
wire S1005;
wire S1006;
wire S1007;
wire S1008;
wire S1009;
wire S1010;
wire S1011;
wire S1012;
wire S1013;
wire S1014;
wire S1015;
wire S1016;
wire S1017;
wire S1018;
wire S1019;
wire S1020;
wire S1021;
wire S1022;
wire S1023;
wire S1024;
wire S1025;
wire S1026;
wire S1027;
wire S1028;
wire S1029;
wire S1030;
wire S1031;
wire S1032;
wire S1033;
wire S1034;
wire S1035;
wire S1036;
wire S1037;
wire S1038;
wire S1039;
wire S1040;
wire S1041;
wire S1042;
wire S1043;
wire S1044;
wire S1045;
wire S1046;
wire S1047;
wire S1048;
wire S1049;
wire S1050;
wire S1051;
wire S1052;
wire S1053;
wire S1054;
wire S1055;
wire S1056;
wire S1057;
wire S1058;
wire S1059;
wire S1060;
wire S1061;
wire S1062;
wire S1063;
wire S1064;
wire S1065;
wire S1066;
wire S1067;
wire S1068;
wire S1069;
wire S1070;
wire S1071;
wire S1072;
wire S1073;
wire S1074;
wire S1075;
wire S1076;
wire S1077;
wire S1078;
wire S1079;
wire S1080;
wire S1081;
wire S1082;
wire S1083;
wire S1084;
wire S1085;
wire S1086;
wire S1087;
wire S1088;
wire S1089;
wire S1090;
wire S1091;
wire S1092;
wire S1093;
wire S1094;
wire S1095;
wire S1096;
wire S1097;
wire S1098;
wire S1099;
wire S1100;
wire S1101;
wire S1102;
wire S1103;
wire S1104;
wire S1105;
wire S1106;
wire S1107;
wire S1108;
wire S1109;
wire S1110;
wire S1111;
wire S1112;
wire S1113;
wire S1114;
wire S1115;
wire S1116;
wire S1117;
wire S1118;
wire S1119;
wire S1120;
wire S1121;
wire S1122;
wire S1123;
wire S1124;
wire S1125;
wire S1126;
wire S1127;
wire S1128;
wire S1129;
wire S1130;
wire S1131;
wire S1132;
wire S1133;
wire S1134;
wire S1135;
wire S1136;
wire S1137;
wire S1138;
wire S1139;
wire S1140;
wire S1141;
wire S1142;
wire S1143;
wire S1144;
wire S1145;
wire S1146;
wire S1147;
wire S1148;
wire S1149;
wire S1150;
wire S1151;
wire S1152;
wire S1153;
wire S1154;
wire S1155;
wire S1156;
wire S1157;
wire S1158;
wire S1159;
wire S1160;
wire S1161;
wire S1162;
wire S1163;
wire S1164;
wire S1165;
wire S1166;
wire S1167;
wire S1168;
wire S1169;
wire S1170;
wire S1171;
wire S1172;
wire S1173;
wire S1174;
wire S1175;
wire S1176;
wire S1177;
wire S1178;
wire S1179;
wire S1180;
wire S1181;
wire S1182;
wire S1183;
wire S1184;
wire S1185;
wire S1186;
wire S1187;
wire S1188;
wire S1189;
wire S1190;
wire S1191;
wire S1192;
wire S1193;
wire S1194;
wire S1195;
wire S1196;
wire S1197;
wire S1198;
wire S1199;
wire S1200;
wire S1201;
wire S1202;
wire S1203;
wire S1204;
wire S1205;
wire S1206;
wire S1207;
wire S1208;
wire S1209;
wire S1210;
wire S1211;
wire S1212;
wire S1213;
wire S1214;
wire S1215;
wire S1216;
wire S1217;
wire S1218;
wire S1219;
wire S1220;
wire S1221;
wire S1222;
wire S1223;
wire S1224;
wire S1225;
wire S1226;
wire S1227;
wire S1228;
wire S1229;
wire S1230;
wire S1231;
wire S1232;
wire S1233;
wire S1234;
wire S1235;
wire S1236;
wire S1237;
wire S1238;
wire S1239;
wire S1240;
wire S1241;
wire S1242;
wire S1243;
wire S1244;
wire S1245;
wire S1246;
wire S1247;
wire S1248;
wire S1249;
wire S1250;
wire S1251;
wire S1252;
wire S1253;
wire S1254;
wire S1255;
wire S1256;
wire S1257;
wire S1258;
wire S1259;
wire S1260;
wire S1261;
wire S1262;
wire S1263;
wire S1264;
wire S1265;
wire S1266;
wire S1267;
wire S1268;
wire S1269;
wire S1270;
wire S1271;
wire S1272;
wire S1273;
wire S1274;
wire S1275;
wire S1276;
wire S1277;
wire S1278;
wire S1279;
wire S1280;
wire S1281;
wire S1282;
wire S1283;
wire S1284;
wire S1285;
wire S1286;
wire S1287;
wire S1288;
wire S1289;
wire S1290;
wire S1291;
wire S1292;
wire S1293;
wire S1294;
wire S1295;
wire S1296;
wire S1297;
wire S1298;
wire S1299;
wire S1300;
wire S1301;
wire S1302;
wire S1303;
wire S1304;
wire S1305;
wire S1306;
wire S1307;
wire S1308;
wire S1309;
wire S1310;
wire S1311;
wire S1312;
wire S1313;
wire S1314;
wire S1315;
wire S1316;
wire S1317;
wire S1318;
wire S1319;
wire S1320;
wire S1321;
wire S1322;
wire S1323;
wire S1324;
wire S1325;
wire S1326;
wire S1327;
wire S1328;
wire S1329;
wire S1330;
wire S1331;
wire S1332;
wire S1333;
wire S1334;
wire S1335;
wire S1336;
wire S1337;
wire S1338;
wire S1339;
wire S1340;
wire S1341;
wire S1342;
wire S1343;
wire S1344;
wire S1345;
wire S1346;
wire S1347;
wire S1348;
wire S1349;
wire S1350;
wire S1351;
wire S1352;
wire S1353;
wire S1354;
wire S1355;
wire S1356;
wire S1357;
wire S1358;
wire S1359;
wire S1360;
wire S1361;
wire S1362;
wire S1363;
wire S1364;
wire S1365;
wire S1366;
wire S1367;
wire S1368;
wire S1369;
wire S1370;
wire S1371;
wire S1372;
wire S1373;
wire S1374;
wire S1375;
wire S1376;
wire S1377;
wire S1378;
wire S1379;
wire S1380;
wire S1381;
wire S1382;
wire S1383;
wire S1384;
wire S1385;
wire S1386;
wire S1387;
wire S1388;
wire S1389;
wire S1390;
wire S1391;
wire S1392;
wire S1393;
wire S1394;
wire S1395;
wire S1396;
wire S1397;
wire S1398;
wire S1399;
wire S1400;
wire S1401;
wire S1402;
wire S1403;
wire S1404;
wire S1405;
wire S1406;
wire S1407;
wire S1408;
wire S1409;
wire S1410;
wire S1411;
wire S1412;
wire S1413;
wire S1414;
wire S1415;
wire S1416;
wire S1417;
wire S1418;
wire S1419;
wire S1420;
wire S1421;
wire S1422;
wire S1423;
wire S1424;
wire S1425;
wire S1426;
wire S1427;
wire S1428;
wire S1429;
wire S1430;
wire S1431;
wire S1432;
wire S1433;
wire S1434;
wire S1435;
wire S1436;
wire S1437;
wire S1438;
wire S1439;
wire S1440;
wire S1441;
wire S1442;
wire S1443;
wire S1444;
wire S1445;
wire S1446;
wire S1447;
wire S1448;
wire S1449;
wire S1450;
wire S1451;
wire S1452;
wire S1453;
wire S1454;
wire S1455;
wire S1456;
wire S1457;
wire S1458;
wire S1459;
wire S1460;
wire S1461;
wire S1462;
wire S1463;
wire S1464;
wire S1465;
wire S1466;
wire S1467;
wire S1468;
wire S1469;
wire S1470;
wire S1471;
wire S1472;
wire S1473;
wire S1474;
wire S1475;
wire S1476;
wire S1477;
wire S1478;
wire S1479;
wire S1480;
wire S1481;
wire S1482;
wire S1483;
wire S1484;
wire S1485;
wire S1486;
wire S1487;
wire S1488;
wire S1489;
wire S1490;
wire S1491;
wire S1492;
wire S1493;
wire S1494;
wire S1495;
wire S1496;
wire S1497;
wire S1498;
wire S1499;
wire S1500;
wire S1501;
wire S1502;
wire S1503;
wire S1504;
wire S1505;
wire S1506;
wire S1507;
wire S1508;
wire S1509;
wire S1510;
wire S1511;
wire S1512;
wire S1513;
wire S1514;
wire S1515;
wire S1516;
wire S1517;
wire S1518;
wire S1519;
wire S1520;
wire S1521;
wire S1522;
wire S1523;
wire S1524;
wire S1525;
wire S1526;
wire S1527;
wire S1528;
wire S1529;
wire S1530;
wire S1531;
wire S1532;
wire S1533;
wire S1534;
wire S1535;
wire S1536;
wire S1537;
wire S1538;
wire S1539;
wire S1540;
wire S1541;
wire S1542;
wire S1543;
wire S1544;
wire S1545;
wire S1546;
wire S1547;
wire S1548;
wire S1549;
wire S1550;
wire S1551;
wire S1552;
wire S1553;
wire S1554;
wire S1555;
wire S1556;
wire S1557;
wire S1558;
wire S1559;
wire S1560;
wire S1561;
wire S1562;
wire S1563;
wire S1564;
wire S1565;
wire S1566;
wire S1567;
wire S1568;
wire S1569;
wire S1570;
wire S1571;
wire S1572;
wire S1573;
wire S1574;
wire S1575;
wire S1576;
wire S1577;
wire S1578;
wire S1579;
wire S1580;
wire S1581;
wire S1582;
wire S1583;
wire S1584;
wire S1585;
wire S1586;
wire S1587;
wire S1588;
wire S1589;
wire S1590;
wire S1591;
wire S1592;
wire S1593;
wire S1594;
wire S1595;
wire S1596;
wire S1597;
wire S1598;
wire S1599;
wire S1600;
wire S1601;
wire S1602;
wire S1603;
wire S1604;
wire S1605;
wire S1606;
wire S1607;
wire S1608;
wire S1609;
wire S1610;
wire S1611;
wire S1612;
wire S1613;
wire S1614;
wire S1615;
wire S1616;
wire S1617;
wire S1618;
wire S1619;
wire S1620;
wire S1621;
wire S1622;
wire S1623;
wire S1624;
wire S1625;
wire S1626;
wire S1627;
wire S1628;
wire S1629;
wire S1630;
wire S1631;
wire S1632;
wire S1633;
wire S1634;
wire S1635;
wire S1636;
wire S1637;
wire S1638;
wire S1639;
wire S1640;
wire S1641;
wire S1642;
wire S1643;
wire S1644;
wire S1645;
wire S1646;
wire S1647;
wire S1648;
wire S1649;
wire S1650;
wire S1651;
wire S1652;
wire S1653;
wire S1654;
wire S1655;
wire S1656;
wire S1657;
wire S1658;
wire S1659;
wire S1660;
wire S1661;
wire S1662;
wire S1663;
wire S1664;
wire S1665;
wire S1666;
wire S1667;
wire S1668;
wire S1669;
wire S1670;
wire S1671;
wire S1672;
wire S1673;
wire S1674;
wire S1675;
wire S1676;
wire S1677;
wire S1678;
wire S1679;
wire S1680;
wire S1681;
wire S1682;
wire S1683;
wire S1684;
wire S1685;
wire S1686;
wire S1687;
wire S1688;
wire S1689;
wire S1690;
wire S1691;
wire S1692;
wire S1693;
wire S1694;
wire S1695;
wire S1696;
wire S1697;
wire S1698;
wire S1699;
wire S1700;
wire S1701;
wire S1702;
wire S1703;
wire S1704;
wire S1705;
wire S1706;
wire S1707;
wire S1708;
wire S1709;
wire S1710;
wire S1711;
wire S1712;
wire S1713;
wire S1714;
wire S1715;
wire S1716;
wire S1717;
wire S1718;
wire S1719;
wire S1720;
wire S1721;
wire S1722;
wire S1723;
wire S1724;
wire S1725;
wire S1726;
wire S1727;
wire S1728;
wire S1729;
wire S1730;
wire S1731;
wire S1732;
wire S1733;
wire S1734;
wire S1735;
wire S1736;
wire S1737;
wire S1738;
wire S1739;
wire S1740;
wire S1741;
wire S1742;
wire S1743;
wire S1744;
wire S1745;
wire S1746;
wire S1747;
wire S1748;
wire S1749;
wire S1750;
wire S1751;
wire S1752;
wire S1753;
wire S1754;
wire S1755;
wire S1756;
wire S1757;
wire S1758;
wire S1759;
wire S1760;
wire S1761;
wire S1762;
wire S1763;
wire S1764;
wire S1765;
wire S1766;
wire S1767;
wire S1768;
wire S1769;
wire S1770;
wire S1771;
wire S1772;
wire S1773;
wire S1774;
wire S1775;
wire S1776;
wire S1777;
wire S1778;
wire S1779;
wire S1780;
wire S1781;
wire S1782;
wire S1783;
wire S1784;
wire S1785;
wire S1786;
wire S1787;
wire S1788;
wire S1789;
wire S1790;
wire S1791;
wire S1792;
wire S1793;
wire S1794;
wire S1795;
wire S1796;
wire S1797;
wire S1798;
wire S1799;
wire S1800;
wire S1801;
wire S1802;
wire S1803;
wire S1804;
wire S1805;
wire S1806;
wire S1807;
wire S1808;
wire S1809;
wire S1810;
wire S1811;
wire S1812;
wire S1813;
wire S1814;
wire S1815;
wire S1816;
wire S1817;
wire S1818;
wire S1819;
wire S1820;
wire S1821;
wire S1822;
wire S1823;
wire S1824;
wire S1825;
wire S1826;
wire S1827;
wire S1828;
wire S1829;
wire S1830;
wire S1831;
wire S1832;
wire S1833;
wire S1834;
wire S1835;
wire S1836;
wire S1837;
wire S1838;
wire S1839;
wire S1840;
wire S1841;
wire S1842;
wire S1843;
wire S1844;
wire S1845;
wire S1846;
wire S1847;
wire S1848;
wire S1849;
wire S1850;
wire S1851;
wire S1852;
wire S1853;
wire S1854;
wire S1855;
wire S1856;
wire S1857;
wire S1858;
wire S1859;
wire S1860;
wire S1861;
wire S1862;
wire S1863;
wire S1864;
wire S1865;
wire S1866;
wire S1867;
wire S1868;
wire S1869;
wire S1870;
wire S1871;
wire S1872;
wire S1873;
wire S1874;
wire S1875;
wire S1876;
wire S1877;
wire S1878;
wire S1879;
wire S1880;
wire S1881;
wire S1882;
wire S1883;
wire S1884;
wire S1885;
wire S1886;
wire S1887;
wire S1888;
wire S1889;
wire S1890;
wire S1891;
wire S1892;
wire S1893;
wire S1894;
wire S1895;
wire S1896;
wire S1897;
wire S1898;
wire S1899;
wire S1900;
wire S1901;
wire S1902;
wire S1903;
wire S1904;
wire S1905;
wire S1906;
wire S1907;
wire S1908;
wire S1909;
wire S1910;
wire S1911;
wire S1912;
wire S1913;
wire S1914;
wire S1915;
wire S1916;
wire S1917;
wire S1918;
wire S1919;
wire S1920;
wire S1921;
wire S1922;
wire S1923;
wire S1924;
wire S1925;
wire S1926;
wire S1927;
wire S1928;
wire S1929;
wire S1930;
wire S1931;
wire S1932;
wire S1933;
wire S1934;
wire S1935;
wire S1936;
wire S1937;
wire S1938;
wire S1939;
wire S1940;
wire S1941;
wire S1942;
wire S1943;
wire S1944;
wire S1945;
wire S1946;
wire S1947;
wire S1948;
wire S1949;
wire S1950;
wire S1951;
wire S1952;
wire S1953;
wire S1954;
wire S1955;
wire S1956;
wire S1957;
wire S1958;
wire S1959;
wire S1960;
wire S1961;
wire S1962;
wire S1963;
wire S1964;
wire S1965;
wire S1966;
wire S1967;
wire S1968;
wire S1969;
wire S1970;
wire S1971;
wire S1972;
wire S1973;
wire S1974;
wire S1975;
wire S1976;
wire S1977;
wire S1978;
wire S1979;
wire S1980;
wire S1981;
wire S1982;
wire S1983;
wire S1984;
wire S1985;
wire S1986;
wire S1987;
wire S1988;
wire S1989;
wire S1990;
wire S1991;
wire S1992;
wire S1993;
wire S1994;
wire S1995;
wire S1996;
wire S1997;
wire S1998;
wire S1999;
wire S2000;
wire S2001;
wire S2002;
wire S2003;
wire S2004;
wire S2005;
wire S2006;
wire S2007;
wire S2008;
wire S2009;
wire S2010;
wire S2011;
wire S2012;
wire S2013;
wire S2014;
wire S2015;
wire S2016;
wire S2017;
wire S2018;
wire S2019;
wire S2020;
wire S2021;
wire S2022;
wire S2023;
wire S2024;
wire S2025;
wire S2026;
wire S2027;
wire S2028;
wire S2029;
wire S2030;
wire S2031;
wire S2032;
wire S2033;
wire S2034;
wire S2035;
wire S2036;
wire S2037;
wire S2038;
wire S2039;
wire S2040;
wire S2041;
wire S2042;
wire S2043;
wire S2044;
wire S2045;
wire S2046;
wire S2047;
wire S2048;
wire S2049;
wire S2050;
wire S2051;
wire S2052;
wire S2053;
wire S2054;
wire S2055;
wire S2056;
wire S2057;
wire S2058;
wire S2059;
wire S2060;
wire S2061;
wire S2062;
wire S2063;
wire S2064;
wire S2065;
wire S2066;
wire S2067;
wire S2068;
wire S2069;
wire S2070;
wire S2071;
wire S2072;
wire S2073;
wire S2074;
wire S2075;
wire S2076;
wire S2077;
wire S2078;
wire S2079;
wire S2080;
wire S2081;
wire S2082;
wire S2083;
wire S2084;
wire S2085;
wire S2086;
wire S2087;
wire S2088;
wire S2089;
wire S2090;
wire S2091;
wire S2092;
wire S2093;
wire S2094;
wire S2095;
wire S2096;
wire S2097;
wire S2098;
wire S2099;
wire S2100;
wire S2101;
wire S2102;
wire S2103;
wire S2104;
wire S2105;
wire S2106;
wire S2107;
wire S2108;
wire S2109;
wire S2110;
wire S2111;
wire S2112;
wire S2113;
wire S2114;
wire S2115;
wire S2116;
wire S2117;
wire S2118;
wire S2119;
wire S2120;
wire S2121;
wire S2122;
wire S2123;
wire S2124;
wire S2125;
wire S2126;
wire S2127;
wire S2128;
wire S2129;
wire S2130;
wire S2131;
wire S2132;
wire S2133;
wire S2134;
wire S2135;
wire S2136;
wire S2137;
wire S2138;
wire S2139;
wire S2140;
wire S2141;
wire S2142;
wire S2143;
wire S2144;
wire S2145;
wire S2146;
wire S2147;
wire S2148;
wire S2149;
wire S2150;
wire S2151;
wire S2152;
wire S2153;
wire S2154;
wire S2155;
wire S2156;
wire S2157;
wire S2158;
wire S2159;
wire S2160;
wire S2161;
wire S2162;
wire S2163;
wire S2164;
wire S2165;
wire S2166;
wire S2167;
wire S2168;
wire S2169;
wire S2170;
wire S2171;
wire S2172;
wire S2173;
wire S2174;
wire S2175;
wire S2176;
wire S2177;
wire S2178;
wire S2179;
wire S2180;
wire S2181;
wire S2182;
wire S2183;
wire S2184;
wire S2185;
wire S2186;
wire S2187;
wire S2188;
wire S2189;
wire S2190;
wire S2191;
wire S2192;
wire S2193;
wire S2194;
wire S2195;
wire S2196;
wire S2197;
wire S2198;
wire S2199;
wire S2200;
wire S2201;
wire S2202;
wire S2203;
wire S2204;
wire S2205;
wire S2206;
wire S2207;
wire S2208;
wire S2209;
wire S2210;
wire S2211;
wire S2212;
wire S2213;
wire S2214;
wire S2215;
wire S2216;
wire S2217;
wire S2218;
wire S2219;
wire S2220;
wire S2221;
wire S2222;
wire S2223;
wire S2224;
wire S2225;
wire S2226;
wire S2227;
wire S2228;
wire S2229;
wire S2230;
wire S2231;
wire S2232;
wire S2233;
wire S2234;
wire S2235;
wire S2236;
wire S2237;
wire S2238;
wire S2239;
wire S2240;
wire S2241;
wire S2242;
wire S2243;
wire S2244;
wire S2245;
wire S2246;
wire S2247;
wire S2248;
wire S2249;
wire S2250;
wire S2251;
wire S2252;
wire S2253;
wire S2254;
wire S2255;
wire S2256;
wire S2257;
wire S2258;
wire S2259;
wire S2260;
wire S2261;
wire S2262;
wire S2263;
wire S2264;
wire S2265;
wire S2266;
wire S2267;
wire S2268;
wire S2269;
wire S2270;
wire S2271;
wire S2272;
wire S2273;
wire S2274;
wire S2275;
wire S2276;
wire S2277;
wire S2278;
wire S2279;
wire S2280;
wire S2281;
wire S2282;
wire S2283;
wire S2284;
wire S2285;
wire S2286;
wire S2287;
wire S2288;
wire S2289;
wire S2290;
wire S2291;
wire S2292;
wire S2293;
wire S2294;
wire S2295;
wire S2296;
wire S2297;
wire S2298;
wire S2299;
wire S2300;
wire S2301;
wire S2302;
wire S2303;
wire S2304;
wire S2305;
wire S2306;
wire S2307;
wire S2308;
wire S2309;
wire S2310;
wire S2311;
wire S2312;
wire S2313;
wire S2314;
wire S2315;
wire S2316;
wire S2317;
wire S2318;
wire S2319;
wire S2320;
wire S2321;
wire S2322;
wire S2323;
wire S2324;
wire S2325;
wire S2326;
wire S2327;
wire S2328;
wire S2329;
wire S2330;
wire S2331;
wire S2332;
wire S2333;
wire S2334;
wire S2335;
wire S2336;
wire S2337;
wire S2338;
wire S2339;
wire S2340;
wire S2341;
wire S2342;
wire S2343;
wire S2344;
wire S2345;
wire S2346;
wire S2347;
wire S2348;
wire S2349;
wire S2350;
wire S2351;
wire S2352;
wire S2353;
wire S2354;
wire S2355;
wire S2356;
wire S2357;
wire S2358;
wire S2359;
wire S2360;
wire S2361;
wire S2362;
wire S2363;
wire S2364;
wire S2365;
wire S2366;
wire S2367;
wire S2368;
wire S2369;
wire S2370;
wire S2371;
wire S2372;
wire S2373;
wire S2374;
wire S2375;
wire S2376;
wire S2377;
wire S2378;
wire S2379;
wire S2380;
wire S2381;
wire S2382;
wire S2383;
wire S2384;
wire S2385;
wire S2386;
wire S2387;
wire S2388;
wire S2389;
wire S2390;
wire S2391;
wire S2392;
wire S2393;
wire S2394;
wire S2395;
wire S2396;
wire S2397;
wire S2398;
wire S2399;
wire S2400;
wire S2401;
wire S2402;
wire S2403;
wire S2404;
wire S2405;
wire S2406;
wire S2407;
wire S2408;
wire S2409;
wire S2410;
wire S2411;
wire S2412;
wire S2413;
wire S2414;
wire S2415;
wire S2416;
wire S2417;
wire S2418;
wire S2419;
wire S2420;
wire S2421;
wire S2422;
wire S2423;
wire S2424;
wire S2425;
wire S2426;
wire S2427;
wire S2428;
wire S2429;
wire S2430;
wire S2431;
wire S2432;
wire S2433;
wire S2434;
wire S2435;
wire S2436;
wire S2437;
wire S2438;
wire S2439;
wire S2440;
wire S2441;
wire S2442;
wire S2443;
wire S2444;
wire S2445;
wire S2446;
wire S2447;
wire S2448;
wire S2449;
wire S2450;
wire S2451;
wire S2452;
wire S2453;
wire S2454;
wire S2455;
wire S2456;
wire S2457;
wire S2458;
wire S2459;
wire S2460;
wire S2461;
wire S2462;
wire S2463;
wire S2464;
wire S2465;
wire S2466;
wire S2467;
wire S2468;
wire S2469;
wire S2470;
wire S2471;
wire S2472;
wire S2473;
wire S2474;
wire S2475;
wire S2476;
wire S2477;
wire S2478;
wire S2479;
wire S2480;
wire S2481;
wire S2482;
wire S2483;
wire S2484;
wire S2485;
wire S2486;
wire S2487;
wire S2488;
wire S2489;
wire S2490;
wire S2491;
wire S2492;
wire S2493;
wire S2494;
wire S2495;
wire S2496;
wire S2497;
wire S2498;
wire S2499;
wire S2500;
wire S2501;
wire S2502;
wire S2503;
wire S2504;
wire S2505;
wire S2506;
wire S2507;
wire S2508;
wire S2509;
wire S2510;
wire S2511;
wire S2512;
wire S2513;
wire S2514;
wire S2515;
wire S2516;
wire S2517;
wire S2518;
wire S2519;
wire S2520;
wire S2521;
wire S2522;
wire S2523;
wire S2524;
wire S2525;
wire S2526;
wire S2527;
wire S2528;
wire S2529;
wire S2530;
wire S2531;
wire S2532;
wire S2533;
wire S2534;
wire S2535;
wire S2536;
wire S2537;
wire S2538;
wire S2539;
wire S2540;
wire S2541;
wire S2542;
wire S2543;
wire S2544;
wire S2545;
wire S2546;
wire S2547;
wire S2548;
wire S2549;
wire S2550;
wire S2551;
wire S2552;
wire S2553;
wire S2554;
wire S2555;
wire S2556;
wire S2557;
wire S2558;
wire S2559;
wire S2560;
wire S2561;
wire S2562;
wire S2563;
wire S2564;
wire S2565;
wire S2566;
wire S2567;
wire S2568;
wire S2569;
wire S2570;
wire S2571;
wire S2572;
wire S2573;
wire S2574;
wire S2575;
wire S2576;
wire S2577;
wire S2578;
wire S2579;
wire S2580;
wire S2581;
wire S2582;
wire S2583;
wire S2584;
wire S2585;
wire S2586;
wire S2587;
wire S2588;
wire S2589;
wire S2590;
wire S2591;
wire S2592;
wire S2593;
wire S2594;
wire S2595;
wire S2596;
wire S2597;
wire S2598;
wire S2599;
wire S2600;
wire S2601;
wire S2602;
wire S2603;
wire S2604;
wire S2605;
wire S2606;
wire S2607;
wire S2608;
wire S2609;
wire S2610;
wire S2611;
wire S2612;
wire S2613;
wire S2614;
wire S2615;
wire S2616;
wire S2617;
wire S2618;
wire S2619;
wire S2620;
wire S2621;
wire S2622;
wire S2623;
wire S2624;
wire S2625;
wire S2626;
wire S2627;
wire S2628;
wire S2629;
wire S2630;
wire S2631;
wire S2632;
wire S2633;
wire S2634;
wire S2635;
wire S2636;
wire S2637;
wire S2638;
wire S2639;
wire S2640;
wire S2641;
wire S2642;
wire S2643;
wire S2644;
wire S2645;
wire S2646;
wire S2647;
wire S2648;
wire S2649;
wire S2650;
wire S2651;
wire S2652;
wire S2653;
wire S2654;
wire S2655;
wire S2656;
wire S2657;
wire S2658;
wire S2659;
wire S2660;
wire S2661;
wire S2662;
wire S2663;
wire S2664;
wire S2665;
wire S2666;
wire S2667;
wire S2668;
wire S2669;
wire S2670;
wire S2671;
wire S2672;
wire S2673;
wire S2674;
wire S2675;
wire S2676;
wire S2677;
wire S2678;
wire S2679;
wire S2680;
wire S2681;
wire S2682;
wire S2683;
wire S2684;
wire S2685;
wire S2686;
wire S2687;
wire S2688;
wire S2689;
wire S2690;
wire S2691;
wire S2692;
wire S2693;
wire S2694;
wire S2695;
wire S2696;
wire S2697;
wire S2698;
wire S2699;
wire S2700;
wire S2701;
wire S2702;
wire S2703;
wire S2704;
wire S2705;
wire S2706;
wire S2707;
wire S2708;
wire S2709;
wire S2710;
wire S2711;
wire S2712;
wire S2713;
wire S2714;
wire S2715;
wire S2716;
wire S2717;
wire S2718;
wire S2719;
wire S2720;
wire S2721;
wire S2722;
wire S2723;
wire S2724;
wire S2725;
wire S2726;
wire S2727;
wire S2728;
wire S2729;
wire S2730;
wire S2731;
wire S2732;
wire S2733;
wire S2734;
wire S2735;
wire S2736;
wire S2737;
wire S2738;
wire S2739;
wire S2740;
wire S2741;
wire S2742;
wire S2743;
wire S2744;
wire S2745;
wire S2746;
wire S2747;
wire S2748;
wire S2749;
wire S2750;
wire S2751;
wire S2752;
wire S2753;
wire S2754;
wire S2755;
wire S2756;
wire S2757;
wire S2758;
wire S2759;
wire S2760;
wire S2761;
wire S2762;
wire S2763;
wire S2764;
wire S2765;
wire S2766;
wire S2767;
wire S2768;
wire S2769;
wire S2770;
wire S2771;
wire S2772;
wire S2773;
wire S2774;
wire S2775;
wire S2776;
wire S2777;
wire S2778;
wire S2779;
wire S2780;
wire S2781;
wire S2782;
wire S2783;
wire S2784;
wire S2785;
wire S2786;
wire S2787;
wire S2788;
wire S2789;
wire S2790;
wire S2791;
wire S2792;
wire S2793;
wire S2794;
wire S2795;
wire S2796;
wire S2797;
wire S2798;
wire S2799;
wire S2800;
wire S2801;
wire S2802;
wire S2803;
wire S2804;
wire S2805;
wire S2806;
wire S2807;
wire S2808;
wire S2809;
wire S2810;
wire S2811;
wire S2812;
wire S2813;
wire S2814;
wire S2815;
wire S2816;
wire S2817;
wire S2818;
wire S2819;
wire S2820;
wire S2821;
wire S2822;
wire S2823;
wire S2824;
wire S2825;
wire S2826;
wire S2827;
wire S2828;
wire S2829;
wire S2830;
wire S2831;
wire S2832;
wire S2833;
wire S2834;
wire S2835;
wire S2836;
wire S2837;
wire S2838;
wire S2839;
wire S2840;
wire S2841;
wire S2842;
wire S2843;
wire S2844;
wire S2845;
wire S2846;
wire S2847;
wire S2848;
wire S2849;
wire S2850;
wire S2851;
wire S2852;
wire S2853;
wire S2854;
wire S2855;
wire S2856;
wire S2857;
wire S2858;
wire S2859;
wire S2860;
wire S2861;
wire S2862;
wire S2863;
wire S2864;
wire S2865;
wire S2866;
wire S2867;
wire S2868;
wire S2869;
wire S2870;
wire S2871;
wire S2872;
wire S2873;
wire S2874;
wire S2875;
wire S2876;
wire S2877;
wire S2878;
wire S2879;
wire S2880;
wire S2881;
wire S2882;
wire S2883;
wire S2884;
wire S2885;
wire S2886;
wire S2887;
wire S2888;
wire S2889;
wire S2890;
wire S2891;
wire S2892;
wire S2893;
wire S2894;
wire S2895;
wire S2896;
wire S2897;
wire S2898;
wire S2899;
wire S2900;
wire S2901;
wire S2902;
wire S2903;
wire S2904;
wire S2905;
wire S2906;
wire S2907;
wire S2908;
wire S2909;
wire S2910;
wire S2911;
wire S2912;
wire S2913;
wire S2914;
wire S2915;
wire S2916;
wire S2917;
wire S2918;
wire S2919;
wire S2920;
wire S2921;
wire S2922;
wire S2923;
wire S2924;
wire S2925;
wire S2926;
wire S2927;
wire S2928;
wire S2929;
wire S2930;
wire S2931;
wire S2932;
wire S2933;
wire S2934;
wire S2935;
wire S2936;
wire S2937;
wire S2938;
wire S2939;
wire S2940;
wire S2941;
wire S2942;
wire S2943;
wire S2944;
wire S2945;
wire S2946;
wire S2947;
wire S2948;
wire S2949;
wire S2950;
wire S2951;
wire S2952;
wire S2953;
wire S2954;
wire S2955;
wire S2956;
wire S2957;
wire S2958;
wire S2959;
wire S2960;
wire S2961;
wire S2962;
wire S2963;
wire S2964;
wire S2965;
wire S2966;
wire S2967;
wire S2968;
wire S2969;
wire S2970;
wire S2971;
wire S2972;
wire S2973;
wire S2974;
wire S2975;
wire S2976;
wire S2977;
wire S2978;
wire S2979;
wire S2980;
wire S2981;
wire S2982;
wire S2983;
wire S2984;
wire S2985;
wire S2986;
wire S2987;
wire S2988;
wire S2989;
wire S2990;
wire S2991;
wire S2992;
wire S2993;
wire S2994;
wire S2995;
wire S2996;
wire S2997;
wire S2998;
wire S2999;
wire S3000;
wire S3001;
wire S3002;
wire S3003;
wire S3004;
wire S3005;
wire S3006;
wire S3007;
wire S3008;
wire S3009;
wire S3010;
wire S3011;
wire S3012;
wire S3013;
wire S3014;
wire S3015;
wire S3016;
wire S3017;
wire S3018;
wire S3019;
wire S3020;
wire S3021;
wire S3022;
wire S3023;
wire S3024;
wire S3025;
wire S3026;
wire S3027;
wire S3028;
wire S3029;
wire S3030;
wire S3031;
wire S3032;
wire S3033;
wire S3034;
wire S3035;
wire S3036;
wire S3037;
wire S3038;
wire S3039;
wire S3040;
wire S3041;
wire S3042;
wire S3043;
wire S3044;
wire S3045;
wire S3046;
wire S3047;
wire S3048;
wire S3049;
wire S3050;
wire S3051;
wire S3052;
wire S3053;
wire S3054;
wire S3055;
wire S3056;
wire S3057;
wire S3058;
wire S3059;
wire S3060;
wire S3061;
wire S3062;
wire S3063;
wire S3064;
wire S3065;
wire S3066;
wire S3067;
wire S3068;
wire S3069;
wire S3070;
wire S3071;
wire S3072;
wire S3073;
wire S3074;
wire S3075;
wire S3076;
wire S3077;
wire S3078;
wire S3079;
wire S3080;
wire S3081;
wire S3082;
wire S3083;
wire S3084;
wire S3085;
wire S3086;
wire S3087;
wire S3088;
wire S3089;
wire S3090;
wire S3091;
wire S3092;
wire S3093;
wire S3094;
wire S3095;
wire S3096;
wire S3097;
wire S3098;
wire S3099;
wire S3100;
wire S3101;
wire S3102;
wire S3103;
wire S3104;
wire S3105;
wire S3106;
wire S3107;
wire S3108;
wire S3109;
wire S3110;
wire S3111;
wire S3112;
wire S3113;
wire S3114;
wire S3115;
wire S3116;
wire S3117;
wire S3118;
wire S3119;
wire S3120;
wire S3121;
wire S3122;
wire S3123;
wire S3124;
wire S3125;
wire S3126;
wire S3127;
wire S3128;
wire S3129;
wire S3130;
wire S3131;
wire S3132;
wire S3133;
wire S3134;
wire S3135;
wire S3136;
wire S3137;
wire S3138;
wire S3139;
wire S3140;
wire S3141;
wire S3142;
wire S3143;
wire S3144;
wire S3145;
wire S3146;
wire S3147;
wire S3148;
wire S3149;
wire S3150;
wire S3151;
wire S3152;
wire S3153;
wire S3154;
wire S3155;
wire S3156;
wire S3157;
wire S3158;
wire S3159;
wire S3160;
wire S3161;
wire S3162;
wire S3163;
wire S3164;
wire S3165;
wire S3166;
wire S3167;
wire S3168;
wire S3169;
wire S3170;
wire S3171;
wire S3172;
wire S3173;
wire S3174;
wire S3175;
wire S3176;
wire S3177;
wire S3178;
wire S3179;
wire S3180;
wire S3181;
wire S3182;
wire S3183;
wire S3184;
wire S3185;
wire S3186;
wire S3187;
wire S3188;
wire S3189;
wire S3190;
wire S3191;
wire S3192;
wire S3193;
wire S3194;
wire S3195;
wire S3196;
wire S3197;
wire S3198;
wire S3199;
wire S3200;
wire S3201;
wire S3202;
wire S3203;
wire S3204;
wire S3205;
wire S3206;
wire S3207;
wire S3208;
wire S3209;
wire S3210;
wire S3211;
wire S3212;
wire S3213;
wire S3214;
wire S3215;
wire S3216;
wire S3217;
wire S3218;
wire S3219;
wire S3220;
wire S3221;
wire S3222;
wire S3223;
wire S3224;
wire S3225;
wire S3226;
wire S3227;
wire S3228;
wire S3229;
wire S3230;
wire S3231;
wire S3232;
wire S3233;
wire S3234;
wire S3235;
wire S3236;
wire S3237;
wire S3238;
wire S3239;
wire S3240;
wire S3241;
wire S3242;
wire S3243;
wire S3244;
wire S3245;
wire S3246;
wire S3247;
wire S3248;
wire S3249;
wire S3250;
wire S3251;
wire S3252;
wire S3253;
wire S3254;
wire S3255;
wire S3256;
wire S3257;
wire S3258;
wire S3259;
wire S3260;
wire S3261;
wire S3262;
wire S3263;
wire S3264;
wire S3265;
wire S3266;
wire S3267;
wire S3268;
wire S3269;
wire S3270;
wire S3271;
wire S3272;
wire S3273;
wire S3274;
wire S3275;
wire S3276;
wire S3277;
wire S3278;
wire S3279;
wire S3280;
wire S3281;
wire S3282;
wire S3283;
wire S3284;
wire S3285;
wire S3286;
wire S3287;
wire S3288;
wire S3289;
wire S3290;
wire S3291;
wire S3292;
wire S3293;
wire S3294;
wire S3295;
wire S3296;
wire S3297;
wire S3298;
wire S3299;
wire S3300;
wire S3301;
wire S3302;
wire S3303;
wire S3304;
wire S3305;
wire S3306;
wire S3307;
wire S3308;
wire S3309;
wire S3310;
wire S3311;
wire S3312;
wire S3313;
wire S3314;
wire S3315;
wire S3316;
wire S3317;
wire S3318;
wire S3319;
wire S3320;
wire S3321;
wire S3322;
wire S3323;
wire S3324;
wire S3325;
wire S3326;
wire S3327;
wire S3328;
wire S3329;
wire S3330;
wire S3331;
wire S3332;
wire S3333;
wire S3334;
wire S3335;
wire S3336;
wire S3337;
wire S3338;
wire S3339;
wire S3340;
wire S3341;
wire S3342;
wire S3343;
wire S3344;
wire S3345;
wire S3346;
wire S3347;
wire S3348;
wire S3349;
wire S3350;
wire S3351;
wire S3352;
wire S3353;
wire S3354;
wire S3355;
wire S3356;
wire S3357;
wire S3358;
wire S3359;
wire S3360;
wire S3361;
wire S3362;
wire S3363;
wire S3364;
wire S3365;
wire S3366;
wire CU_ADD;
wire CU_AND;
wire CU_INC1;
wire CU_INC2;
wire CU_LSB0E;
wire CU_MUL;
wire CU_NOT;
wire CU_SE12bits;
wire CU_SE4bits;
wire CU_SHF_0;
wire CU_SHF_1;
wire CU_clk;
wire CU_conOF;
wire CU_enSKP;
wire CU_inst_0;
wire CU_inst_10;
wire CU_inst_11;
wire CU_inst_12;
wire CU_inst_13;
wire CU_inst_14;
wire CU_inst_15;
wire CU_inst_1;
wire CU_inst_2;
wire CU_inst_3;
wire CU_inst_4;
wire CU_inst_5;
wire CU_inst_6;
wire CU_inst_7;
wire CU_inst_8;
wire CU_inst_9;
wire CU_ldAC;
wire CU_ldIN;
wire CU_ldIR;
wire CU_ldOF;
wire CU_ldPC;
wire CU_ldSR_0;
wire CU_ldSR_1;
wire CU_ldSR_2;
wire CU_ldSR_3;
wire CU_nstate_0;
wire CU_nstate_1;
wire CU_pstate_0;
wire CU_pstate_1;
wire CU_readMEM;
wire CU_rst;
wire CU_sel1_ARU;
wire CU_selAC_MEM;
wire CU_selARU_AC;
wire CU_selARU_SR;
wire CU_selIMM_AC;
wire CU_selIMM_LGU;
wire CU_selIMM_OF;
wire CU_selIMM_PC;
wire CU_selINC_IN;
wire CU_selINC_PC;
wire CU_selIN_ADR;
wire CU_selIN_MEM;
wire CU_selIR_ADR;
wire CU_selLGU_AC;
wire CU_selLGU_SR;
wire CU_selMEM_AC;
wire CU_selMEM_IN;
wire CU_selMEM_LGU;
wire CU_selMEM_PC;
wire CU_selPC_MEM;
wire CU_selPC_OF;
wire CU_selSET_SR;
wire CU_seldataBus;
wire CU_zeroAC;
wire DP_AC_in_0;
wire DP_AC_in_10;
wire DP_AC_in_11;
wire DP_AC_in_12;
wire DP_AC_in_13;
wire DP_AC_in_14;
wire DP_AC_in_15;
wire DP_AC_in_1;
wire DP_AC_in_2;
wire DP_AC_in_3;
wire DP_AC_in_4;
wire DP_AC_in_5;
wire DP_AC_in_6;
wire DP_AC_in_7;
wire DP_AC_in_8;
wire DP_AC_in_9;
wire DP_AC_out_0;
wire DP_AC_out_10;
wire DP_AC_out_11;
wire DP_AC_out_12;
wire DP_AC_out_13;
wire DP_AC_out_14;
wire DP_AC_out_15;
wire DP_AC_out_1;
wire DP_AC_out_2;
wire DP_AC_out_3;
wire DP_AC_out_4;
wire DP_AC_out_5;
wire DP_AC_out_6;
wire DP_AC_out_7;
wire DP_AC_out_8;
wire DP_AC_out_9;
wire DP_ARU1_C;
wire DP_ARU1_N;
wire DP_ARU1_V;
wire DP_ARU1_Z;
wire DP_ARU1_in1_0;
wire DP_ARU1_in1_10;
wire DP_ARU1_in1_11;
wire DP_ARU1_in1_12;
wire DP_ARU1_in1_13;
wire DP_ARU1_in1_14;
wire DP_ARU1_in1_15;
wire DP_ARU1_in1_1;
wire DP_ARU1_in1_2;
wire DP_ARU1_in1_3;
wire DP_ARU1_in1_4;
wire DP_ARU1_in1_5;
wire DP_ARU1_in1_6;
wire DP_ARU1_in1_7;
wire DP_ARU1_in1_8;
wire DP_ARU1_in1_9;
wire DP_ARU1_out_0;
wire DP_ARU1_out_10;
wire DP_ARU1_out_11;
wire DP_ARU1_out_12;
wire DP_ARU1_out_13;
wire DP_ARU1_out_14;
wire DP_ARU1_out_1;
wire DP_ARU1_out_2;
wire DP_ARU1_out_3;
wire DP_ARU1_out_4;
wire DP_ARU1_out_5;
wire DP_ARU1_out_6;
wire DP_ARU1_out_7;
wire DP_ARU1_out_8;
wire DP_ARU1_out_9;
wire DP_IMM1_in1_0;
wire DP_IMM1_in1_1;
wire DP_IMM1_in1_2;
wire DP_IMM1_in1_3;
wire DP_IMM1_out_0;
wire DP_IMM1_out_10;
wire DP_IMM1_out_11;
wire DP_IMM1_out_12;
wire DP_IMM1_out_13;
wire DP_IMM1_out_14;
wire DP_IMM1_out_15;
wire DP_IMM1_out_1;
wire DP_IMM1_out_2;
wire DP_IMM1_out_3;
wire DP_IMM1_out_4;
wire DP_IMM1_out_5;
wire DP_IMM1_out_6;
wire DP_IMM1_out_7;
wire DP_IMM1_out_8;
wire DP_IMM1_out_9;
wire DP_IN_in_0;
wire DP_IN_in_10;
wire DP_IN_in_11;
wire DP_IN_in_12;
wire DP_IN_in_13;
wire DP_IN_in_14;
wire DP_IN_in_15;
wire DP_IN_in_1;
wire DP_IN_in_2;
wire DP_IN_in_3;
wire DP_IN_in_4;
wire DP_IN_in_5;
wire DP_IN_in_6;
wire DP_IN_in_7;
wire DP_IN_in_8;
wire DP_IN_in_9;
wire DP_IN_out_0;
wire DP_IN_out_10;
wire DP_IN_out_11;
wire DP_IN_out_12;
wire DP_IN_out_13;
wire DP_IN_out_14;
wire DP_IN_out_15;
wire DP_IN_out_1;
wire DP_IN_out_2;
wire DP_IN_out_3;
wire DP_IN_out_4;
wire DP_IN_out_5;
wire DP_IN_out_6;
wire DP_IN_out_7;
wire DP_IN_out_8;
wire DP_IN_out_9;
wire DP_INC2_out_0;
wire DP_INC2_out_10;
wire DP_INC2_out_11;
wire DP_INC2_out_12;
wire DP_INC2_out_13;
wire DP_INC2_out_14;
wire DP_INC2_out_15;
wire DP_INC2_out_1;
wire DP_INC2_out_2;
wire DP_INC2_out_3;
wire DP_INC2_out_4;
wire DP_INC2_out_5;
wire DP_INC2_out_6;
wire DP_INC2_out_7;
wire DP_INC2_out_8;
wire DP_INC2_out_9;
wire DP_INC_1_in_0;
wire DP_INC_1_in_10;
wire DP_INC_1_in_11;
wire DP_INC_1_in_12;
wire DP_INC_1_in_13;
wire DP_INC_1_in_14;
wire DP_INC_1_in_15;
wire DP_INC_1_in_1;
wire DP_INC_1_in_2;
wire DP_INC_1_in_3;
wire DP_INC_1_in_4;
wire DP_INC_1_in_5;
wire DP_INC_1_in_6;
wire DP_INC_1_in_7;
wire DP_INC_1_in_8;
wire DP_INC_1_in_9;
wire DP_INC_1_inc_val_0;
wire DP_INC_1_inc_val_1;
wire DP_INC_1_out_0;
wire DP_INC_1_out_10;
wire DP_INC_1_out_11;
wire DP_INC_1_out_12;
wire DP_INC_1_out_13;
wire DP_INC_1_out_14;
wire DP_INC_1_out_15;
wire DP_INC_1_out_1;
wire DP_INC_1_out_2;
wire DP_INC_1_out_3;
wire DP_INC_1_out_4;
wire DP_INC_1_out_5;
wire DP_INC_1_out_6;
wire DP_INC_1_out_7;
wire DP_INC_1_out_8;
wire DP_INC_1_out_9;
wire DP_LGU1_N;
wire DP_LGU1_Z;
wire DP_LGU1_in1_0;
wire DP_LGU1_in1_10;
wire DP_LGU1_in1_11;
wire DP_LGU1_in1_12;
wire DP_LGU1_in1_13;
wire DP_LGU1_in1_14;
wire DP_LGU1_in1_15;
wire DP_LGU1_in1_1;
wire DP_LGU1_in1_2;
wire DP_LGU1_in1_3;
wire DP_LGU1_in1_4;
wire DP_LGU1_in1_5;
wire DP_LGU1_in1_6;
wire DP_LGU1_in1_7;
wire DP_LGU1_in1_8;
wire DP_LGU1_in1_9;
wire DP_LGU1_out_0;
wire DP_LGU1_out_10;
wire DP_LGU1_out_11;
wire DP_LGU1_out_12;
wire DP_LGU1_out_13;
wire DP_LGU1_out_14;
wire DP_LGU1_out_1;
wire DP_LGU1_out_2;
wire DP_LGU1_out_3;
wire DP_LGU1_out_4;
wire DP_LGU1_out_5;
wire DP_LGU1_out_6;
wire DP_LGU1_out_7;
wire DP_LGU1_out_8;
wire DP_LGU1_out_9;
wire DP_OF_in_0;
wire DP_OF_in_1;
wire DP_OF_in_2;
wire DP_OF_in_3;
wire DP_PC_in_0;
wire DP_PC_in_10;
wire DP_PC_in_11;
wire DP_PC_in_12;
wire DP_PC_in_13;
wire DP_PC_in_14;
wire DP_PC_in_15;
wire DP_PC_in_1;
wire DP_PC_in_2;
wire DP_PC_in_3;
wire DP_PC_in_4;
wire DP_PC_in_5;
wire DP_PC_in_6;
wire DP_PC_in_7;
wire DP_PC_in_8;
wire DP_PC_in_9;
wire DP_SR_C_in;
wire DP_SR_C_out;
wire DP_SR_N_in;
wire DP_SR_N_out;
wire DP_SR_V_in;
wire DP_SR_V_out;
wire DP_SR_Z_in;
wire DP_SR_Z_out;
wire DP_addrBus_0;
wire DP_addrBus_10;
wire DP_addrBus_11;
wire DP_addrBus_12;
wire DP_addrBus_13;
wire DP_addrBus_14;
wire DP_addrBus_15;
wire DP_addrBus_1;
wire DP_addrBus_2;
wire DP_addrBus_3;
wire DP_addrBus_4;
wire DP_addrBus_5;
wire DP_addrBus_6;
wire DP_addrBus_7;
wire DP_addrBus_8;
wire DP_addrBus_9;
input clk;
input rst;
output writeMEM;
output readMEM;
output [15:0] addrBus;
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_1_ (
  .in1({ 1'b1 }),
  .out1({ S0 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_2_ (
  .in1({ 1'b1 }),
  .out1({ S1 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_3_ (
  .in1({ 1'b1 }),
  .out1({ S2 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_4_ (
  .in1({ 1'b1 }),
  .out1({ S3 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_5_ (
  .in1({ 1'b1 }),
  .out1({ S4 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_6_ (
  .in1({ 1'b1 }),
  .out1({ S5 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_7_ (
  .in1({ 1'b0 }),
  .out1({ S6 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_8_ (
  .in1({ 1'b0 }),
  .out1({ S7 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_9_ (
  .in1({ 1'b0 }),
  .out1({ S8 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_10_ (
  .in1({ 1'b0 }),
  .out1({ S9 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_11_ (
  .in1({ 1'b0 }),
  .out1({ S10 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_12_ (
  .in1({ 1'b0 }),
  .out1({ S11 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_13_ (
  .in1({ 1'b0 }),
  .out1({ S12 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_14_ (
  .in1({ 1'b0 }),
  .out1({ S13 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_15_ (
  .in1({ 1'b0 }),
  .out1({ S14 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_16_ (
  .in1({ 1'b0 }),
  .out1({ S15 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_17_ (
  .in1({ 1'b0 }),
  .out1({ S16 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_18_ (
  .in1({ 1'b0 }),
  .out1({ S17 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_19_ (
  .in1({ 1'b0 }),
  .out1({ S18 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_20_ (
  .in1({ 1'b0 }),
  .out1({ S19 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_21_ (
  .in1({ 1'b0 }),
  .out1({ S20 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_22_ (
  .in1({ 1'b0 }),
  .out1({ S21 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_23_ (
  .in1({ 1'b0 }),
  .out1({ S22 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_24_ (
  .in1({ 1'b0 }),
  .out1({ S23 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_25_ (
  .in1({ 1'b0 }),
  .out1({ S24 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_26_ (
  .in1({ 1'b0 }),
  .out1({ S25 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_27_ (
  .in1({ 1'b0 }),
  .out1({ S26 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_28_ (
  .in1({ 1'b0 }),
  .out1({ S27 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_29_ (
  .in1({ 1'b0 }),
  .out1({ S28 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_30_ (
  .in1({ 1'b0 }),
  .out1({ S29 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_31_ (
  .in1({ 1'b0 }),
  .out1({ S30 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_32_ (
  .in1({ 1'b0 }),
  .out1({ S31 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_33_ (
  .in1({ 1'b0 }),
  .out1({ S32 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_34_ (
  .in1({ 1'b0 }),
  .out1({ S33 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_35_ (
  .in1({ 1'b0 }),
  .out1({ S34 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_36_ (
  .in1({ 1'b0 }),
  .out1({ S35 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_37_ (
  .in1({ 1'b0 }),
  .out1({ S36 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_38_ (
  .in1({ 1'b0 }),
  .out1({ S37 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1_ (
  .in1({ S130, S129 }),
  .out1({ S131 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1_ (
  .in1({ S70, CU_ldIR }),
  .out1({ S132 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_2_ (
  .in1({ S132, S131 }),
  .out1({ CU_readMEM })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_2_ (
  .in1({ S129, CU_selIN_MEM }),
  .out1({ S133 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_1_ (
  .in1({ S133 }),
  .out1({ CU_conOF })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_3_ (
  .in1({ S240, CU_inst_13 }),
  .out1({ S134 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_2_ (
  .in1({ S134 }),
  .out1({ S135 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_4_ (
  .in1({ S135, CU_inst_12 }),
  .out1({ S136 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_5_ (
  .in1({ S136, S133 }),
  .out1({ CU_selIR_ADR })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_6_ (
  .in1({ CU_inst_14, S220 }),
  .out1({ S137 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_3_ (
  .in1({ S50, CU_inst_12 }),
  .out1({ S138 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_7_ (
  .in1({ S138, CU_inst_13 }),
  .out1({ S139 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_8_ (
  .in1({ S134, S120 }),
  .out1({ S140 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_9_ (
  .in1({ S134, S121 }),
  .out1({ S141 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_10_ (
  .in1({ S139, S124 }),
  .out1({ S142 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_4_ (
  .in1({ S142, S141 }),
  .out1({ S143 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_5_ (
  .in1({ S106, S74 }),
  .out1({ S144 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_6_ (
  .in1({ S144, S60 }),
  .out1({ S145 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_7_ (
  .in1({ S65, S238 }),
  .out1({ S146 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_11_ (
  .in1({ S146, S143 }),
  .out1({ S147 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_8_ (
  .in1({ S147, S145 }),
  .out1({ S148 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_9_ (
  .in1({ S148, S235 }),
  .out1({ CU_seldataBus })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_10_ (
  .in1({ S68, S230 }),
  .out1({ S149 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_12_ (
  .in1({ S92, CU_inst_1 }),
  .out1({ S150 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_3_ (
  .in1({ S150 }),
  .out1({ S151 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_11_ (
  .in1({ S150, S100 }),
  .out1({ S152 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_13_ (
  .in1({ S88, S245 }),
  .out1({ S153 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_12_ (
  .in1({ S89, S244 }),
  .out1({ S154 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_13_ (
  .in1({ S153, S152 }),
  .out1({ S155 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_14_ (
  .in1({ CU_inst_9, S224 }),
  .out1({ S156 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_15_ (
  .in1({ S44, S229 }),
  .out1({ S157 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_14_ (
  .in1({ S156, CU_enSKP }),
  .out1({ S158 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_16_ (
  .in1({ S158, S44 }),
  .out1({ S159 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_15_ (
  .in1({ S157, S156 }),
  .out1({ S160 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_16_ (
  .in1({ S88, S244 }),
  .out1({ S161 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_17_ (
  .in1({ S161, S159 }),
  .out1({ S162 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_17_ (
  .in1({ S60, CU_inst_14 }),
  .out1({ S163 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_18_ (
  .in1({ S163, S64 }),
  .out1({ S164 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_19_ (
  .in1({ S164, S49 }),
  .out1({ S165 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_18_ (
  .in1({ S165, S162 }),
  .out1({ S166 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_20_ (
  .in1({ S166, S155 }),
  .out1({ S167 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_21_ (
  .in1({ S167, S238 }),
  .out1({ S168 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_22_ (
  .in1({ S168, S149 }),
  .out1({ CU_INC1 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_23_ (
  .in1({ S113, S71 }),
  .out1({ CU_selARU_SR })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_19_ (
  .in1({ S154, S152 }),
  .out1({ S169 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_4_ (
  .in1({ S169 }),
  .out1({ S170 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_24_ (
  .in1({ S135, S238 }),
  .out1({ S171 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_20_ (
  .in1({ S171, S169 }),
  .out1({ S172 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_25_ (
  .in1({ S172, S67 }),
  .out1({ S173 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_26_ (
  .in1({ S173, S149 }),
  .out1({ CU_selINC_PC })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_27_ (
  .in1({ S149, S146 }),
  .out1({ CU_ldPC })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_28_ (
  .in1({ S84, CU_inst_2 }),
  .out1({ S174 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_21_ (
  .in1({ S174, S88 }),
  .out1({ S175 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_29_ (
  .in1({ S175, S150 }),
  .out1({ S176 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_30_ (
  .in1({ S176, S244 }),
  .out1({ S177 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_5_ (
  .in1({ S177 }),
  .out1({ S178 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_31_ (
  .in1({ S140, S67 }),
  .out1({ S179 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_22_ (
  .in1({ S179, S239 }),
  .out1({ S180 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_32_ (
  .in1({ S138, S106 }),
  .out1({ S181 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_33_ (
  .in1({ S177, S138 }),
  .out1({ S182 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_23_ (
  .in1({ S182, S107 }),
  .out1({ S183 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_34_ (
  .in1({ S183, S180 }),
  .out1({ S184 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_35_ (
  .in1({ S184, S71 }),
  .out1({ CU_selARU_AC })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_24_ (
  .in1({ S69, CU_inst_15 }),
  .out1({ S185 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_6_ (
  .in1({ S185 }),
  .out1({ S186 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_36_ (
  .in1({ S139, S238 }),
  .out1({ S187 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_37_ (
  .in1({ S187, S186 }),
  .out1({ CU_selMEM_AC })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_38_ (
  .in1({ S47, S42 }),
  .out1({ S188 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_25_ (
  .in1({ S188, S102 }),
  .out1({ S189 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_39_ (
  .in1({ S189, S178 }),
  .out1({ S190 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_40_ (
  .in1({ S134, CU_inst_12 }),
  .out1({ S191 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_41_ (
  .in1({ S191, S130 }),
  .out1({ S192 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_26_ (
  .in1({ S192, S146 }),
  .out1({ S193 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_42_ (
  .in1({ S193, S190 }),
  .out1({ S194 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_43_ (
  .in1({ S194, S69 }),
  .out1({ CU_ldAC })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_44_ (
  .in1({ S144, S122 }),
  .out1({ S195 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_45_ (
  .in1({ S195, S71 }),
  .out1({ CU_selMEM_LGU })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_46_ (
  .in1({ S73, S242 }),
  .out1({ S196 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_27_ (
  .in1({ S181, S239 }),
  .out1({ S197 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_47_ (
  .in1({ S196, S177 }),
  .out1({ S198 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_28_ (
  .in1({ S198, S179 }),
  .out1({ S199 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_48_ (
  .in1({ S199, S197 }),
  .out1({ S200 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_49_ (
  .in1({ S200, S71 }),
  .out1({ CU_ADD })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_29_ (
  .in1({ S137, S75 }),
  .out1({ S201 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_50_ (
  .in1({ S201, S180 }),
  .out1({ S202 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_51_ (
  .in1({ S98, S244 }),
  .out1({ S203 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_30_ (
  .in1({ S203, S102 }),
  .out1({ S204 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_31_ (
  .in1({ S204, S202 }),
  .out1({ CU_selLGU_SR })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_32_ (
  .in1({ S160, S40 }),
  .out1({ CU_INC2 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_33_ (
  .in1({ S63, S55 }),
  .out1({ S205 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_52_ (
  .in1({ S69, S56 }),
  .out1({ CU_selIN_ADR })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_53_ (
  .in1({ S156, S41 }),
  .out1({ S206 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_7_ (
  .in1({ S206 }),
  .out1({ CU_selIMM_OF })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_54_ (
  .in1({ S87, S238 }),
  .out1({ S207 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_34_ (
  .in1({ S207, S151 }),
  .out1({ S208 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_55_ (
  .in1({ S208, S153 }),
  .out1({ S209 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_8_ (
  .in1({ S209 }),
  .out1({ CU_selPC_OF })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_56_ (
  .in1({ S209, S206 }),
  .out1({ CU_ldOF })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_35_ (
  .in1({ S205, S239 }),
  .out1({ CU_selMEM_IN })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_36_ (
  .in1({ S123, S234 }),
  .out1({ CU_selINC_IN })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_37_ (
  .in1({ S170, S239 }),
  .out1({ CU_LSB0E })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_38_ (
  .in1({ S169, S58 }),
  .out1({ S210 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_39_ (
  .in1({ S210, S239 }),
  .out1({ CU_selIMM_PC })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_40_ (
  .in1({ S135, S123 }),
  .out1({ CU_selMEM_PC })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_57_ (
  .in1({ S189, S244 }),
  .out1({ S211 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_9_ (
  .in1({ S211 }),
  .out1({ S212 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_41_ (
  .in1({ S212, S202 }),
  .out1({ CU_selLGU_AC })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_42_ (
  .in1({ S119, S239 }),
  .out1({ CU_selIMM_AC })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_43_ (
  .in1({ S188, S245 }),
  .out1({ S213 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_44_ (
  .in1({ S137, S48 }),
  .out1({ S214 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_58_ (
  .in1({ S214, S180 }),
  .out1({ S215 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_45_ (
  .in1({ S215, S213 }),
  .out1({ CU_selIMM_LGU })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_46_ (
  .in1({ S176, S40 }),
  .out1({ CU_sel1_ARU })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_59_ (
  .in1({ S214, S240 }),
  .out1({ S216 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_47_ (
  .in1({ S216, S146 }),
  .out1({ CU_SE4bits })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_60_ (
  .in1({ S188, S39 }),
  .out1({ S217 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_61_ (
  .in1({ S217, S206 }),
  .out1({ CU_SE12bits })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_48_ (
  .in1({ S196, S239 }),
  .out1({ CU_MUL })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_10_ (
  .in1({ CU_pstate_0 }),
  .out1({ S218 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_11_ (
  .in1({ CU_pstate_1 }),
  .out1({ S219 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_12_ (
  .in1({ CU_inst_12 }),
  .out1({ S220 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_13_ (
  .in1({ CU_inst_13 }),
  .out1({ S221 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_14_ (
  .in1({ CU_inst_14 }),
  .out1({ S222 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_15_ (
  .in1({ CU_inst_15 }),
  .out1({ S223 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_16_ (
  .in1({ CU_inst_8 }),
  .out1({ S224 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_17_ (
  .in1({ CU_inst_11 }),
  .out1({ S225 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_18_ (
  .in1({ CU_rst }),
  .out1({ S226 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_19_ (
  .in1({ CU_inst_1 }),
  .out1({ S227 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_20_ (
  .in1({ CU_inst_3 }),
  .out1({ S228 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_21_ (
  .in1({ CU_enSKP }),
  .out1({ S229 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_49_ (
  .in1({ CU_pstate_1, CU_pstate_0 }),
  .out1({ CU_ldIR })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_50_ (
  .in1({ S219, CU_pstate_0 }),
  .out1({ S230 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_51_ (
  .in1({ CU_inst_15, S222 }),
  .out1({ S231 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_62_ (
  .in1({ S223, CU_inst_14 }),
  .out1({ S232 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_52_ (
  .in1({ S232, CU_inst_13 }),
  .out1({ S233 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_63_ (
  .in1({ S231, S221 }),
  .out1({ S234 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_64_ (
  .in1({ S233, S230 }),
  .out1({ S235 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_53_ (
  .in1({ S235, S220 }),
  .out1({ CU_selIN_MEM })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_54_ (
  .in1({ CU_inst_10, CU_inst_11 }),
  .out1({ S236 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_22_ (
  .in1({ S236 }),
  .out1({ S237 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_55_ (
  .in1({ CU_pstate_1, S218 }),
  .out1({ S238 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_65_ (
  .in1({ S219, CU_pstate_0 }),
  .out1({ S239 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_66_ (
  .in1({ CU_inst_15, CU_inst_14 }),
  .out1({ S240 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_23_ (
  .in1({ S240 }),
  .out1({ S241 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_56_ (
  .in1({ S221, S220 }),
  .out1({ S242 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_67_ (
  .in1({ CU_inst_13, CU_inst_12 }),
  .out1({ S243 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_57_ (
  .in1({ S243, S240 }),
  .out1({ S244 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_68_ (
  .in1({ S242, S241 }),
  .out1({ S245 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_58_ (
  .in1({ S245, S239 }),
  .out1({ S39 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_69_ (
  .in1({ S244, S238 }),
  .out1({ S40 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_59_ (
  .in1({ S40, S237 }),
  .out1({ S41 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_70_ (
  .in1({ S236, CU_inst_9 }),
  .out1({ S42 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_71_ (
  .in1({ S39, CU_inst_8 }),
  .out1({ S43 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_60_ (
  .in1({ S43, S42 }),
  .out1({ CU_SHF_0 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_72_ (
  .in1({ CU_inst_10, S225 }),
  .out1({ S44 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_24_ (
  .in1({ S44 }),
  .out1({ S45 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_61_ (
  .in1({ CU_inst_9, CU_inst_8 }),
  .out1({ S46 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_73_ (
  .in1({ S46, S45 }),
  .out1({ S47 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_62_ (
  .in1({ S47, S40 }),
  .out1({ CU_SHF_1 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_63_ (
  .in1({ S243, CU_inst_15 }),
  .out1({ S48 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_74_ (
  .in1({ S242, S223 }),
  .out1({ S49 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_64_ (
  .in1({ CU_inst_15, CU_inst_14 }),
  .out1({ S50 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_65_ (
  .in1({ S49, CU_inst_14 }),
  .out1({ S51 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_75_ (
  .in1({ S51, S238 }),
  .out1({ S52 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_66_ (
  .in1({ CU_inst_13, CU_inst_12 }),
  .out1({ S53 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_76_ (
  .in1({ S221, S220 }),
  .out1({ S54 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_67_ (
  .in1({ S54, S232 }),
  .out1({ S55 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_77_ (
  .in1({ S55, S230 }),
  .out1({ S56 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_78_ (
  .in1({ S56, S52 }),
  .out1({ CU_selAC_MEM })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_79_ (
  .in1({ S239, S226 }),
  .out1({ S57 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_68_ (
  .in1({ S57, S230 }),
  .out1({ S246 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_69_ (
  .in1({ S240, CU_inst_12 }),
  .out1({ S58 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_70_ (
  .in1({ S221, CU_inst_12 }),
  .out1({ S59 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_80_ (
  .in1({ CU_inst_13, S220 }),
  .out1({ S60 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_81_ (
  .in1({ S58, CU_inst_13 }),
  .out1({ S61 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_25_ (
  .in1({ S61 }),
  .out1({ S62 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_71_ (
  .in1({ S61, S239 }),
  .out1({ CU_selPC_MEM })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_72_ (
  .in1({ S60, CU_inst_14 }),
  .out1({ S63 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_82_ (
  .in1({ S59, S222 }),
  .out1({ S64 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_73_ (
  .in1({ S63, S233 }),
  .out1({ S65 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_83_ (
  .in1({ S64, S234 }),
  .out1({ S66 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_74_ (
  .in1({ S65, S239 }),
  .out1({ CU_ldIN })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_75_ (
  .in1({ S66, S62 }),
  .out1({ S67 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_84_ (
  .in1({ S65, S61 }),
  .out1({ S68 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_76_ (
  .in1({ S67, S239 }),
  .out1({ S247 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_85_ (
  .in1({ S63, S230 }),
  .out1({ S69 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_26_ (
  .in1({ S69 }),
  .out1({ S70 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_86_ (
  .in1({ S70, CU_inst_15 }),
  .out1({ S71 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_27_ (
  .in1({ S71 }),
  .out1({ S72 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_77_ (
  .in1({ S223, CU_inst_14 }),
  .out1({ S73 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_87_ (
  .in1({ CU_inst_15, S222 }),
  .out1({ S74 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_78_ (
  .in1({ S74, CU_inst_13 }),
  .out1({ S75 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_28_ (
  .in1({ S75 }),
  .out1({ S76 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_79_ (
  .in1({ S76, S239 }),
  .out1({ S77 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_88_ (
  .in1({ S75, S238 }),
  .out1({ S78 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_80_ (
  .in1({ S77, S72 }),
  .out1({ S79 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_81_ (
  .in1({ S44, CU_inst_8 }),
  .out1({ S80 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_89_ (
  .in1({ S80, CU_inst_9 }),
  .out1({ S81 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_82_ (
  .in1({ S81, S40 }),
  .out1({ CU_selSET_SR })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_90_ (
  .in1({ CU_selSET_SR, CU_inst_4 }),
  .out1({ S82 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_91_ (
  .in1({ S82, S79 }),
  .out1({ CU_ldSR_0 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_92_ (
  .in1({ CU_selSET_SR, CU_inst_5 }),
  .out1({ S83 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_93_ (
  .in1({ S83, S79 }),
  .out1({ CU_ldSR_1 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_83_ (
  .in1({ CU_inst_3, CU_inst_0 }),
  .out1({ S84 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_29_ (
  .in1({ S84 }),
  .out1({ S85 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_84_ (
  .in1({ CU_inst_2, CU_inst_3 }),
  .out1({ S86 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_85_ (
  .in1({ S85, CU_inst_2 }),
  .out1({ S87 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_94_ (
  .in1({ S46, S236 }),
  .out1({ S88 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_30_ (
  .in1({ S88 }),
  .out1({ S89 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_86_ (
  .in1({ CU_inst_5, CU_inst_4 }),
  .out1({ S90 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_87_ (
  .in1({ CU_inst_7, CU_inst_6 }),
  .out1({ S91 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_95_ (
  .in1({ S91, S90 }),
  .out1({ S92 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_31_ (
  .in1({ S92 }),
  .out1({ S93 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_88_ (
  .in1({ S92, S227 }),
  .out1({ S94 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_96_ (
  .in1({ S93, CU_inst_1 }),
  .out1({ S95 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_89_ (
  .in1({ S95, S88 }),
  .out1({ S96 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_97_ (
  .in1({ S94, S89 }),
  .out1({ S97 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_98_ (
  .in1({ S96, S87 }),
  .out1({ S98 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_90_ (
  .in1({ S98, S40 }),
  .out1({ CU_zeroAC })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_99_ (
  .in1({ S228, CU_inst_0 }),
  .out1({ S99 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_91_ (
  .in1({ S99, CU_inst_2 }),
  .out1({ S100 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_100_ (
  .in1({ S86, CU_inst_0 }),
  .out1({ S101 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_92_ (
  .in1({ S101, S97 }),
  .out1({ S102 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_101_ (
  .in1({ S102, S39 }),
  .out1({ S103 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_32_ (
  .in1({ S103 }),
  .out1({ CU_NOT })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_102_ (
  .in1({ S103, S71 }),
  .out1({ S104 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_93_ (
  .in1({ S104, CU_zeroAC }),
  .out1({ S105 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_103_ (
  .in1({ S231, CU_inst_13 }),
  .out1({ S106 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_33_ (
  .in1({ S106 }),
  .out1({ S107 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_94_ (
  .in1({ S106, S239 }),
  .out1({ CU_AND })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_34_ (
  .in1({ CU_AND }),
  .out1({ S108 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_104_ (
  .in1({ CU_selSET_SR, CU_inst_6 }),
  .out1({ S109 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_105_ (
  .in1({ S109, S78 }),
  .out1({ S110 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_95_ (
  .in1({ S110, CU_AND }),
  .out1({ S111 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_106_ (
  .in1({ S111, S105 }),
  .out1({ CU_ldSR_2 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_96_ (
  .in1({ S74, S59 }),
  .out1({ S112 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_107_ (
  .in1({ S112, S238 }),
  .out1({ S113 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_108_ (
  .in1({ S113, S108 }),
  .out1({ S114 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_109_ (
  .in1({ CU_selSET_SR, CU_inst_7 }),
  .out1({ S115 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_35_ (
  .in1({ S115 }),
  .out1({ S116 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_97_ (
  .in1({ S116, S114 }),
  .out1({ S117 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_110_ (
  .in1({ S117, S105 }),
  .out1({ CU_ldSR_3 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_111_ (
  .in1({ CU_pstate_1, CU_pstate_0 }),
  .out1({ S118 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_36_ (
  .in1({ S118 }),
  .out1({ S38 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_112_ (
  .in1({ S53, S50 }),
  .out1({ S119 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_37_ (
  .in1({ S119 }),
  .out1({ S120 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_113_ (
  .in1({ S119, S245 }),
  .out1({ S121 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_98_ (
  .in1({ S239, S220 }),
  .out1({ S122 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_114_ (
  .in1({ S238, CU_inst_12 }),
  .out1({ S123 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_99_ (
  .in1({ S60, S232 }),
  .out1({ S124 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_100_ (
  .in1({ S74, S54 }),
  .out1({ S125 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_101_ (
  .in1({ S125, S124 }),
  .out1({ S126 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_102_ (
  .in1({ S121, S239 }),
  .out1({ S127 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_115_ (
  .in1({ S127, S126 }),
  .out1({ S128 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_38_ (
  .in1({ S128 }),
  .out1({ S129 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_103_ (
  .in1({ S58, S51 }),
  .out1({ S130 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__1_ (
  .D({ S246 }),
  .E({ S38 }),
  .Q({ CU_nstate_0 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__2_ (
  .D({ S247 }),
  .E({ S38 }),
  .Q({ CU_nstate_1 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_1_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ CU_nstate_0 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_pstate_0 }),
  .Si({ S3365 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_2_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ CU_nstate_1 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_pstate_1 }),
  .Si({ S3366 }),
  .global_reset({ 1'b0 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_39_ (
  .in1({ DP_SR_V_out }),
  .out1({ S248 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_40_ (
  .in1({ DP_SR_C_out }),
  .out1({ S249 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_41_ (
  .in1({ DP_SR_N_out }),
  .out1({ S250 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_42_ (
  .in1({ DP_SR_Z_out }),
  .out1({ S251 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_104_ (
  .in1({ S250, CU_inst_2 }),
  .out1({ S252 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_116_ (
  .in1({ S250, CU_inst_2 }),
  .out1({ S253 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_117_ (
  .in1({ S253, CU_inst_6 }),
  .out1({ S254 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_105_ (
  .in1({ S254, S252 }),
  .out1({ S255 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_106_ (
  .in1({ S251, CU_inst_3 }),
  .out1({ S256 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_118_ (
  .in1({ S251, CU_inst_3 }),
  .out1({ S257 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_119_ (
  .in1({ S257, CU_inst_7 }),
  .out1({ S258 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_107_ (
  .in1({ S258, S256 }),
  .out1({ S259 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_108_ (
  .in1({ S259, S255 }),
  .out1({ S260 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_109_ (
  .in1({ S248, CU_inst_0 }),
  .out1({ S261 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_120_ (
  .in1({ S248, CU_inst_0 }),
  .out1({ S262 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_121_ (
  .in1({ S262, CU_inst_4 }),
  .out1({ S263 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_110_ (
  .in1({ S263, S261 }),
  .out1({ S264 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_111_ (
  .in1({ S249, CU_inst_1 }),
  .out1({ S265 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_122_ (
  .in1({ S249, CU_inst_1 }),
  .out1({ S266 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_123_ (
  .in1({ S266, CU_inst_5 }),
  .out1({ S267 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_112_ (
  .in1({ S267, S265 }),
  .out1({ S268 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_113_ (
  .in1({ S268, S264 }),
  .out1({ S269 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_124_ (
  .in1({ S269, S260 }),
  .out1({ CU_enSKP })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_43_ (
  .in1({ CU_ldAC }),
  .out1({ S287 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_114_ (
  .in1({ CU_ldAC, CU_zeroAC }),
  .out1({ S288 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_125_ (
  .in1({ S288, DP_AC_out_0 }),
  .out1({ S289 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_115_ (
  .in1({ S287, CU_zeroAC }),
  .out1({ S290 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_126_ (
  .in1({ S290, DP_AC_in_0 }),
  .out1({ S291 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_127_ (
  .in1({ S291, S289 }),
  .out1({ S270 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_128_ (
  .in1({ S288, DP_AC_out_1 }),
  .out1({ S292 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_129_ (
  .in1({ S290, DP_AC_in_1 }),
  .out1({ S293 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_130_ (
  .in1({ S293, S292 }),
  .out1({ S271 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_131_ (
  .in1({ S288, DP_AC_out_2 }),
  .out1({ S294 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_132_ (
  .in1({ S290, DP_AC_in_2 }),
  .out1({ S295 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_133_ (
  .in1({ S295, S294 }),
  .out1({ S272 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_134_ (
  .in1({ S288, DP_AC_out_3 }),
  .out1({ S296 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_135_ (
  .in1({ S290, DP_AC_in_3 }),
  .out1({ S297 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_136_ (
  .in1({ S297, S296 }),
  .out1({ S273 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_137_ (
  .in1({ S288, DP_AC_out_4 }),
  .out1({ S298 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_138_ (
  .in1({ S290, DP_AC_in_4 }),
  .out1({ S299 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_139_ (
  .in1({ S299, S298 }),
  .out1({ S274 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_140_ (
  .in1({ S288, DP_AC_out_5 }),
  .out1({ S300 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_141_ (
  .in1({ S290, DP_AC_in_5 }),
  .out1({ S301 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_142_ (
  .in1({ S301, S300 }),
  .out1({ S275 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_143_ (
  .in1({ S288, DP_AC_out_6 }),
  .out1({ S302 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_144_ (
  .in1({ S290, DP_AC_in_6 }),
  .out1({ S303 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_145_ (
  .in1({ S303, S302 }),
  .out1({ S276 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_146_ (
  .in1({ S288, DP_AC_out_7 }),
  .out1({ S304 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_147_ (
  .in1({ S290, DP_AC_in_7 }),
  .out1({ S305 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_148_ (
  .in1({ S305, S304 }),
  .out1({ S277 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_149_ (
  .in1({ S288, DP_AC_out_8 }),
  .out1({ S306 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_150_ (
  .in1({ S290, DP_AC_in_8 }),
  .out1({ S307 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_151_ (
  .in1({ S307, S306 }),
  .out1({ S278 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_152_ (
  .in1({ S288, DP_AC_out_9 }),
  .out1({ S308 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_153_ (
  .in1({ S290, DP_AC_in_9 }),
  .out1({ S309 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_154_ (
  .in1({ S309, S308 }),
  .out1({ S279 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_155_ (
  .in1({ S288, DP_AC_out_10 }),
  .out1({ S310 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_156_ (
  .in1({ S290, DP_AC_in_10 }),
  .out1({ S311 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_157_ (
  .in1({ S311, S310 }),
  .out1({ S280 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_158_ (
  .in1({ S288, DP_AC_out_11 }),
  .out1({ S312 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_159_ (
  .in1({ S290, DP_AC_in_11 }),
  .out1({ S313 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_160_ (
  .in1({ S313, S312 }),
  .out1({ S281 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_161_ (
  .in1({ S288, DP_AC_out_12 }),
  .out1({ S314 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_162_ (
  .in1({ S290, DP_AC_in_12 }),
  .out1({ S315 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_163_ (
  .in1({ S315, S314 }),
  .out1({ S282 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_164_ (
  .in1({ S288, DP_AC_out_13 }),
  .out1({ S316 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_165_ (
  .in1({ S290, DP_AC_in_13 }),
  .out1({ S317 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_166_ (
  .in1({ S317, S316 }),
  .out1({ S283 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_167_ (
  .in1({ S288, DP_AC_out_14 }),
  .out1({ S318 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_168_ (
  .in1({ S290, DP_AC_in_14 }),
  .out1({ S319 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_169_ (
  .in1({ S319, S318 }),
  .out1({ S284 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_170_ (
  .in1({ S288, DP_AC_out_15 }),
  .out1({ S320 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_171_ (
  .in1({ S290, DP_AC_in_15 }),
  .out1({ S286 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_172_ (
  .in1({ S286, S320 }),
  .out1({ S285 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_3_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S270 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_out_0 }),
  .Si({ S3307 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_4_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S271 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_out_1 }),
  .Si({ S3306 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_5_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S272 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_out_2 }),
  .Si({ S3305 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_6_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S273 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_out_3 }),
  .Si({ S3304 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_7_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S274 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_out_4 }),
  .Si({ S3303 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_8_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S275 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_out_5 }),
  .Si({ S3302 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_9_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S276 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_out_6 }),
  .Si({ S3301 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_10_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S277 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_out_7 }),
  .Si({ S3300 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_11_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S278 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_out_8 }),
  .Si({ S3299 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_12_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S279 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_out_9 }),
  .Si({ S3298 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_13_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S280 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_out_10 }),
  .Si({ S3297 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_14_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S281 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_out_11 }),
  .Si({ S3296 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_15_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S282 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_out_12 }),
  .Si({ S3295 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_16_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S283 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_out_13 }),
  .Si({ S3294 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_17_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S284 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_out_14 }),
  .Si({ S3293 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_18_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S285 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_out_15 }),
  .Si({ S3356 }),
  .global_reset({ 1'b0 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_44_ (
  .in1({ DP_AC_out_0 }),
  .out1({ S966 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_45_ (
  .in1({ DP_ARU1_in1_0 }),
  .out1({ S977 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_46_ (
  .in1({ CU_ADD }),
  .out1({ S988 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_47_ (
  .in1({ DP_AC_out_1 }),
  .out1({ S998 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_48_ (
  .in1({ DP_ARU1_in1_1 }),
  .out1({ S1009 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_49_ (
  .in1({ DP_AC_out_2 }),
  .out1({ S1020 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_50_ (
  .in1({ DP_ARU1_in1_2 }),
  .out1({ S1031 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_51_ (
  .in1({ DP_AC_out_3 }),
  .out1({ S1042 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_52_ (
  .in1({ DP_ARU1_in1_3 }),
  .out1({ S1053 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_53_ (
  .in1({ DP_AC_out_4 }),
  .out1({ S1064 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_54_ (
  .in1({ DP_ARU1_in1_4 }),
  .out1({ S1075 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_55_ (
  .in1({ DP_AC_out_5 }),
  .out1({ S1085 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_56_ (
  .in1({ DP_ARU1_in1_5 }),
  .out1({ S1096 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_57_ (
  .in1({ DP_AC_out_6 }),
  .out1({ S1107 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_58_ (
  .in1({ DP_ARU1_in1_6 }),
  .out1({ S1118 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_59_ (
  .in1({ DP_AC_out_7 }),
  .out1({ S1129 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_60_ (
  .in1({ DP_ARU1_in1_7 }),
  .out1({ S1140 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_61_ (
  .in1({ DP_AC_out_9 }),
  .out1({ S1150 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_62_ (
  .in1({ DP_ARU1_in1_9 }),
  .out1({ S1161 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_63_ (
  .in1({ DP_AC_out_11 }),
  .out1({ S1172 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_64_ (
  .in1({ DP_ARU1_in1_11 }),
  .out1({ S1183 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_65_ (
  .in1({ DP_AC_out_13 }),
  .out1({ S1194 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_66_ (
  .in1({ DP_ARU1_in1_13 }),
  .out1({ S1205 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_67_ (
  .in1({ DP_AC_out_14 }),
  .out1({ S1215 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_68_ (
  .in1({ DP_ARU1_in1_14 }),
  .out1({ S1226 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_116_ (
  .in1({ DP_ARU1_out_7, DP_ARU1_out_4 }),
  .out1({ S1237 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_117_ (
  .in1({ DP_ARU1_out_2, DP_ARU1_out_1 }),
  .out1({ S1248 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_173_ (
  .in1({ S1248, S1237 }),
  .out1({ S1258 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_118_ (
  .in1({ DP_ARU1_out_14, DP_ARU1_out_13 }),
  .out1({ S1269 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_119_ (
  .in1({ DP_ARU1_out_11, DP_ARU1_out_8 }),
  .out1({ S348 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_174_ (
  .in1({ S348, S1269 }),
  .out1({ S358 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_120_ (
  .in1({ S358, S1258 }),
  .out1({ S359 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_121_ (
  .in1({ DP_ARU1_out_6, DP_ARU1_out_5 }),
  .out1({ S360 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_122_ (
  .in1({ DP_ARU1_out_3, DP_ARU1_out_0 }),
  .out1({ S361 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_175_ (
  .in1({ S361, S360 }),
  .out1({ S362 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_123_ (
  .in1({ DP_ARU1_N, DP_ARU1_out_12 }),
  .out1({ S363 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_124_ (
  .in1({ DP_ARU1_out_10, DP_ARU1_out_9 }),
  .out1({ S364 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_176_ (
  .in1({ S364, S363 }),
  .out1({ S365 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_125_ (
  .in1({ S365, S362 }),
  .out1({ S366 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_177_ (
  .in1({ S366, S359 }),
  .out1({ S367 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_69_ (
  .in1({ S367 }),
  .out1({ DP_ARU1_Z })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_126_ (
  .in1({ DP_ARU1_in1_15, DP_AC_out_15 }),
  .out1({ S368 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_178_ (
  .in1({ S368, DP_ARU1_N }),
  .out1({ S369 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_179_ (
  .in1({ DP_ARU1_in1_15, DP_AC_out_15 }),
  .out1({ S370 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_70_ (
  .in1({ S370 }),
  .out1({ S371 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_127_ (
  .in1({ S370, DP_ARU1_N }),
  .out1({ S372 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_71_ (
  .in1({ S372 }),
  .out1({ S373 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_180_ (
  .in1({ S373, S369 }),
  .out1({ DP_ARU1_V })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_128_ (
  .in1({ DP_ARU1_in1_0, DP_AC_out_0 }),
  .out1({ S374 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_129_ (
  .in1({ S977, S966 }),
  .out1({ S375 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_181_ (
  .in1({ DP_ARU1_in1_0, DP_AC_out_0 }),
  .out1({ S376 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_130_ (
  .in1({ S376, S988 }),
  .out1({ S377 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_131_ (
  .in1({ S374, S988 }),
  .out1({ S378 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_132_ (
  .in1({ S378, S375 }),
  .out1({ S379 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_133_ (
  .in1({ S379, S377 }),
  .out1({ S321 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_134_ (
  .in1({ S1009, S998 }),
  .out1({ S380 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_182_ (
  .in1({ DP_ARU1_in1_1, DP_AC_out_1 }),
  .out1({ S381 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_135_ (
  .in1({ DP_ARU1_in1_1, DP_AC_out_1 }),
  .out1({ S382 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_136_ (
  .in1({ S382, S380 }),
  .out1({ S383 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_183_ (
  .in1({ S383, S375 }),
  .out1({ S384 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_137_ (
  .in1({ S383, S375 }),
  .out1({ S385 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_184_ (
  .in1({ DP_ARU1_in1_1, DP_AC_out_0 }),
  .out1({ S386 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_185_ (
  .in1({ DP_AC_out_1, DP_ARU1_in1_0 }),
  .out1({ S387 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_138_ (
  .in1({ S381, S376 }),
  .out1({ S388 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_186_ (
  .in1({ S387, S386 }),
  .out1({ S389 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_72_ (
  .in1({ S389 }),
  .out1({ S390 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_139_ (
  .in1({ S390, S388 }),
  .out1({ S391 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_187_ (
  .in1({ S391, S988 }),
  .out1({ S392 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_140_ (
  .in1({ S385, S988 }),
  .out1({ S393 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_188_ (
  .in1({ S393, S384 }),
  .out1({ S394 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_189_ (
  .in1({ S394, S392 }),
  .out1({ S328 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_190_ (
  .in1({ S384, S381 }),
  .out1({ S395 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_141_ (
  .in1({ DP_ARU1_in1_2, DP_AC_out_2 }),
  .out1({ S396 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_142_ (
  .in1({ S1031, S1020 }),
  .out1({ S397 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_191_ (
  .in1({ DP_ARU1_in1_2, DP_AC_out_2 }),
  .out1({ S398 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_143_ (
  .in1({ S397, S396 }),
  .out1({ S399 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_144_ (
  .in1({ S399, S395 }),
  .out1({ S400 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_192_ (
  .in1({ S399, S395 }),
  .out1({ S401 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_73_ (
  .in1({ S401 }),
  .out1({ S402 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_145_ (
  .in1({ S402, S400 }),
  .out1({ S403 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_193_ (
  .in1({ DP_ARU1_in1_2, DP_AC_out_0 }),
  .out1({ S404 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_194_ (
  .in1({ DP_AC_out_2, DP_ARU1_in1_0 }),
  .out1({ S405 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_195_ (
  .in1({ DP_AC_out_2, DP_ARU1_in1_1 }),
  .out1({ S406 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_74_ (
  .in1({ S406 }),
  .out1({ S407 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_146_ (
  .in1({ S405, S381 }),
  .out1({ S408 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_75_ (
  .in1({ S408 }),
  .out1({ S409 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_196_ (
  .in1({ S405, S381 }),
  .out1({ S410 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_197_ (
  .in1({ S410, S409 }),
  .out1({ S411 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_198_ (
  .in1({ S411, S404 }),
  .out1({ S412 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_76_ (
  .in1({ S412 }),
  .out1({ S413 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_147_ (
  .in1({ S411, S404 }),
  .out1({ S414 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_148_ (
  .in1({ S414, S413 }),
  .out1({ S415 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_199_ (
  .in1({ S415, S388 }),
  .out1({ S416 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_149_ (
  .in1({ S415, S388 }),
  .out1({ S417 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_150_ (
  .in1({ S417, CU_ADD }),
  .out1({ S418 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_200_ (
  .in1({ S418, S416 }),
  .out1({ S419 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_201_ (
  .in1({ S403, CU_ADD }),
  .out1({ S420 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_202_ (
  .in1({ S420, S419 }),
  .out1({ S329 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_203_ (
  .in1({ S401, S398 }),
  .out1({ S421 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_151_ (
  .in1({ DP_ARU1_in1_3, DP_AC_out_3 }),
  .out1({ S422 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_152_ (
  .in1({ S1053, S1042 }),
  .out1({ S423 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_204_ (
  .in1({ DP_ARU1_in1_3, DP_AC_out_3 }),
  .out1({ S424 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_153_ (
  .in1({ S423, S422 }),
  .out1({ S425 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_205_ (
  .in1({ S425, S421 }),
  .out1({ S426 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_77_ (
  .in1({ S426 }),
  .out1({ S427 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_154_ (
  .in1({ S425, S421 }),
  .out1({ S428 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_155_ (
  .in1({ S428, S427 }),
  .out1({ S429 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_206_ (
  .in1({ S429, CU_ADD }),
  .out1({ S430 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_207_ (
  .in1({ DP_ARU1_in1_3, DP_AC_out_0 }),
  .out1({ S431 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_78_ (
  .in1({ S431 }),
  .out1({ S432 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_156_ (
  .in1({ S414, S408 }),
  .out1({ S433 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_79_ (
  .in1({ S433 }),
  .out1({ S434 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_208_ (
  .in1({ DP_ARU1_in1_2, DP_AC_out_1 }),
  .out1({ S435 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_80_ (
  .in1({ S435 }),
  .out1({ S436 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_209_ (
  .in1({ DP_AC_out_3, DP_ARU1_in1_0 }),
  .out1({ S437 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_81_ (
  .in1({ S437 }),
  .out1({ S438 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_210_ (
  .in1({ DP_AC_out_3, DP_ARU1_in1_1 }),
  .out1({ S439 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_157_ (
  .in1({ S437, S406 }),
  .out1({ S440 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_211_ (
  .in1({ S438, S407 }),
  .out1({ S441 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_212_ (
  .in1({ S437, S406 }),
  .out1({ S442 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_82_ (
  .in1({ S442 }),
  .out1({ S443 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_158_ (
  .in1({ S443, S440 }),
  .out1({ S444 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_213_ (
  .in1({ S442, S441 }),
  .out1({ S445 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_214_ (
  .in1({ S445, S435 }),
  .out1({ S446 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_159_ (
  .in1({ S445, S435 }),
  .out1({ S447 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_215_ (
  .in1({ S444, S436 }),
  .out1({ S448 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_216_ (
  .in1({ S448, S446 }),
  .out1({ S449 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_83_ (
  .in1({ S449 }),
  .out1({ S450 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_217_ (
  .in1({ S450, S434 }),
  .out1({ S451 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_84_ (
  .in1({ S451 }),
  .out1({ S452 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_218_ (
  .in1({ S449, S433 }),
  .out1({ S453 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_219_ (
  .in1({ S453, S451 }),
  .out1({ S454 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_85_ (
  .in1({ S454 }),
  .out1({ S455 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_220_ (
  .in1({ S454, S431 }),
  .out1({ S456 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_160_ (
  .in1({ S454, S431 }),
  .out1({ S457 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_221_ (
  .in1({ S455, S432 }),
  .out1({ S458 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_222_ (
  .in1({ S458, S456 }),
  .out1({ S459 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_223_ (
  .in1({ S459, S416 }),
  .out1({ S460 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_161_ (
  .in1({ S459, S416 }),
  .out1({ S461 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_86_ (
  .in1({ S461 }),
  .out1({ S462 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_162_ (
  .in1({ S461, CU_ADD }),
  .out1({ S463 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_224_ (
  .in1({ S463, S460 }),
  .out1({ S464 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_225_ (
  .in1({ S464, S430 }),
  .out1({ S330 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_163_ (
  .in1({ DP_ARU1_in1_4, DP_AC_out_4 }),
  .out1({ S465 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_164_ (
  .in1({ S1075, S1064 }),
  .out1({ S466 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_226_ (
  .in1({ DP_ARU1_in1_4, DP_AC_out_4 }),
  .out1({ S467 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_165_ (
  .in1({ S466, S465 }),
  .out1({ S468 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_166_ (
  .in1({ S423, S421 }),
  .out1({ S469 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_167_ (
  .in1({ S469, S422 }),
  .out1({ S470 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_227_ (
  .in1({ S470, S468 }),
  .out1({ S471 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_87_ (
  .in1({ S471 }),
  .out1({ S472 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_168_ (
  .in1({ S470, S468 }),
  .out1({ S473 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_169_ (
  .in1({ S473, S472 }),
  .out1({ S474 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_170_ (
  .in1({ S474, S988 }),
  .out1({ S475 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_171_ (
  .in1({ S457, S452 }),
  .out1({ S476 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_228_ (
  .in1({ S458, S451 }),
  .out1({ S477 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_229_ (
  .in1({ DP_ARU1_in1_4, DP_AC_out_0 }),
  .out1({ S478 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_230_ (
  .in1({ DP_ARU1_in1_3, DP_AC_out_1 }),
  .out1({ S479 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_231_ (
  .in1({ S479, S478 }),
  .out1({ S480 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_88_ (
  .in1({ S480 }),
  .out1({ S481 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_232_ (
  .in1({ DP_ARU1_in1_4, DP_AC_out_1 }),
  .out1({ S482 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_89_ (
  .in1({ S482 }),
  .out1({ S483 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_172_ (
  .in1({ S482, S431 }),
  .out1({ S484 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_233_ (
  .in1({ S483, S432 }),
  .out1({ S485 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_173_ (
  .in1({ S484, S481 }),
  .out1({ S486 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_90_ (
  .in1({ S486 }),
  .out1({ S487 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_174_ (
  .in1({ S447, S440 }),
  .out1({ S488 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_234_ (
  .in1({ S448, S441 }),
  .out1({ S489 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_235_ (
  .in1({ DP_AC_out_4, DP_ARU1_in1_0 }),
  .out1({ S490 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_236_ (
  .in1({ DP_AC_out_4, DP_ARU1_in1_1 }),
  .out1({ S491 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_91_ (
  .in1({ S491 }),
  .out1({ S492 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_175_ (
  .in1({ S490, S439 }),
  .out1({ S493 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_237_ (
  .in1({ S492, S438 }),
  .out1({ S494 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_238_ (
  .in1({ S490, S439 }),
  .out1({ S495 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_92_ (
  .in1({ S495 }),
  .out1({ S496 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_176_ (
  .in1({ S496, S493 }),
  .out1({ S497 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_239_ (
  .in1({ S495, S494 }),
  .out1({ S498 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_177_ (
  .in1({ S497, S397 }),
  .out1({ S499 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_240_ (
  .in1({ S498, S398 }),
  .out1({ S500 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_178_ (
  .in1({ S498, S398 }),
  .out1({ S501 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_241_ (
  .in1({ S497, S397 }),
  .out1({ S502 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_179_ (
  .in1({ S501, S499 }),
  .out1({ S503 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_242_ (
  .in1({ S502, S500 }),
  .out1({ S504 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_180_ (
  .in1({ S504, S488 }),
  .out1({ S505 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_243_ (
  .in1({ S503, S489 }),
  .out1({ S506 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_181_ (
  .in1({ S503, S489 }),
  .out1({ S507 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_244_ (
  .in1({ S504, S488 }),
  .out1({ S508 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_182_ (
  .in1({ S507, S505 }),
  .out1({ S509 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_245_ (
  .in1({ S508, S506 }),
  .out1({ S510 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_183_ (
  .in1({ S509, S486 }),
  .out1({ S511 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_184_ (
  .in1({ S510, S487 }),
  .out1({ S512 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_246_ (
  .in1({ S509, S486 }),
  .out1({ S513 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_185_ (
  .in1({ S512, S511 }),
  .out1({ S514 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_93_ (
  .in1({ S514 }),
  .out1({ S515 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_186_ (
  .in1({ S515, S476 }),
  .out1({ S516 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_94_ (
  .in1({ S516 }),
  .out1({ S517 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_187_ (
  .in1({ S514, S477 }),
  .out1({ S518 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_188_ (
  .in1({ S518, S516 }),
  .out1({ S519 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_95_ (
  .in1({ S519 }),
  .out1({ S520 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_189_ (
  .in1({ S519, S461 }),
  .out1({ S521 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_190_ (
  .in1({ S520, S462 }),
  .out1({ S522 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_96_ (
  .in1({ S522 }),
  .out1({ S523 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_191_ (
  .in1({ S522, S521 }),
  .out1({ S524 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_192_ (
  .in1({ S524, CU_ADD }),
  .out1({ S525 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_193_ (
  .in1({ S525, S475 }),
  .out1({ S331 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_247_ (
  .in1({ S471, S467 }),
  .out1({ S526 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_194_ (
  .in1({ DP_ARU1_in1_5, DP_AC_out_5 }),
  .out1({ S527 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_195_ (
  .in1({ S1096, S1085 }),
  .out1({ S528 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_248_ (
  .in1({ DP_ARU1_in1_5, DP_AC_out_5 }),
  .out1({ S529 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_196_ (
  .in1({ S528, S527 }),
  .out1({ S530 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_197_ (
  .in1({ S530, S526 }),
  .out1({ S531 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_249_ (
  .in1({ S530, S526 }),
  .out1({ S532 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_97_ (
  .in1({ S532 }),
  .out1({ S533 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_198_ (
  .in1({ S533, S531 }),
  .out1({ S534 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_199_ (
  .in1({ S534, S988 }),
  .out1({ S535 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_200_ (
  .in1({ S512, S505 }),
  .out1({ S536 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_250_ (
  .in1({ S513, S506 }),
  .out1({ S537 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_251_ (
  .in1({ DP_ARU1_in1_5, DP_AC_out_0 }),
  .out1({ S538 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_252_ (
  .in1({ DP_ARU1_in1_3, DP_AC_out_2 }),
  .out1({ S539 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_253_ (
  .in1({ DP_ARU1_in1_4, DP_AC_out_2 }),
  .out1({ S540 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_201_ (
  .in1({ S539, S482 }),
  .out1({ S541 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_98_ (
  .in1({ S541 }),
  .out1({ S542 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_254_ (
  .in1({ S539, S482 }),
  .out1({ S543 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_255_ (
  .in1({ S543, S542 }),
  .out1({ S544 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_256_ (
  .in1({ S544, S538 }),
  .out1({ S545 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_99_ (
  .in1({ S545 }),
  .out1({ S546 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_202_ (
  .in1({ S544, S538 }),
  .out1({ S547 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_100_ (
  .in1({ S547 }),
  .out1({ S548 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_203_ (
  .in1({ S547, S546 }),
  .out1({ S549 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_257_ (
  .in1({ S548, S545 }),
  .out1({ S550 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_204_ (
  .in1({ S501, S493 }),
  .out1({ S551 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_258_ (
  .in1({ S502, S494 }),
  .out1({ S552 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_259_ (
  .in1({ DP_AC_out_3, DP_ARU1_in1_2 }),
  .out1({ S553 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_101_ (
  .in1({ S553 }),
  .out1({ S554 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_260_ (
  .in1({ DP_AC_out_5, DP_ARU1_in1_0 }),
  .out1({ S555 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_102_ (
  .in1({ S555 }),
  .out1({ S556 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_261_ (
  .in1({ DP_AC_out_5, DP_ARU1_in1_1 }),
  .out1({ S557 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_205_ (
  .in1({ S555, S491 }),
  .out1({ S558 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_262_ (
  .in1({ S556, S492 }),
  .out1({ S559 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_263_ (
  .in1({ S555, S491 }),
  .out1({ S560 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_103_ (
  .in1({ S560 }),
  .out1({ S561 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_206_ (
  .in1({ S561, S558 }),
  .out1({ S562 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_264_ (
  .in1({ S560, S559 }),
  .out1({ S563 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_207_ (
  .in1({ S562, S554 }),
  .out1({ S564 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_265_ (
  .in1({ S563, S553 }),
  .out1({ S565 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_208_ (
  .in1({ S563, S553 }),
  .out1({ S566 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_266_ (
  .in1({ S562, S554 }),
  .out1({ S567 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_209_ (
  .in1({ S566, S564 }),
  .out1({ S568 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_267_ (
  .in1({ S567, S565 }),
  .out1({ S569 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_210_ (
  .in1({ S569, S551 }),
  .out1({ S570 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_268_ (
  .in1({ S568, S552 }),
  .out1({ S571 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_211_ (
  .in1({ S568, S552 }),
  .out1({ S572 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_269_ (
  .in1({ S569, S551 }),
  .out1({ S573 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_212_ (
  .in1({ S572, S570 }),
  .out1({ S574 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_270_ (
  .in1({ S573, S571 }),
  .out1({ S575 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_213_ (
  .in1({ S574, S549 }),
  .out1({ S576 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_271_ (
  .in1({ S575, S550 }),
  .out1({ S577 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_214_ (
  .in1({ S575, S550 }),
  .out1({ S578 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_272_ (
  .in1({ S574, S549 }),
  .out1({ S579 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_215_ (
  .in1({ S578, S576 }),
  .out1({ S580 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_273_ (
  .in1({ S579, S577 }),
  .out1({ S581 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_216_ (
  .in1({ S581, S536 }),
  .out1({ S582 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_274_ (
  .in1({ S580, S537 }),
  .out1({ S583 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_217_ (
  .in1({ S580, S537 }),
  .out1({ S584 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_275_ (
  .in1({ S581, S536 }),
  .out1({ S585 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_218_ (
  .in1({ S584, S582 }),
  .out1({ S586 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_276_ (
  .in1({ S585, S583 }),
  .out1({ S587 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_219_ (
  .in1({ S587, S485 }),
  .out1({ S588 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_277_ (
  .in1({ S586, S484 }),
  .out1({ S589 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_220_ (
  .in1({ S586, S484 }),
  .out1({ S590 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_278_ (
  .in1({ S587, S485 }),
  .out1({ S591 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_221_ (
  .in1({ S590, S588 }),
  .out1({ S592 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_279_ (
  .in1({ S591, S589 }),
  .out1({ S593 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_222_ (
  .in1({ S593, S517 }),
  .out1({ S594 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_280_ (
  .in1({ S592, S516 }),
  .out1({ S595 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_223_ (
  .in1({ S592, S516 }),
  .out1({ S596 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_224_ (
  .in1({ S596, S594 }),
  .out1({ S597 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_104_ (
  .in1({ S597 }),
  .out1({ S598 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_225_ (
  .in1({ S597, S522 }),
  .out1({ S599 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_226_ (
  .in1({ S598, S523 }),
  .out1({ S600 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_281_ (
  .in1({ S597, S522 }),
  .out1({ S601 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_227_ (
  .in1({ S600, S599 }),
  .out1({ S602 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_228_ (
  .in1({ S602, CU_ADD }),
  .out1({ S603 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_229_ (
  .in1({ S603, S535 }),
  .out1({ S332 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_282_ (
  .in1({ S532, S529 }),
  .out1({ S604 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_230_ (
  .in1({ DP_ARU1_in1_6, DP_AC_out_6 }),
  .out1({ S605 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_231_ (
  .in1({ S1118, S1107 }),
  .out1({ S606 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_283_ (
  .in1({ DP_ARU1_in1_6, DP_AC_out_6 }),
  .out1({ S607 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_232_ (
  .in1({ S606, S605 }),
  .out1({ S608 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_233_ (
  .in1({ S608, S604 }),
  .out1({ S609 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_284_ (
  .in1({ S608, S604 }),
  .out1({ S610 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_234_ (
  .in1({ S588, S582 }),
  .out1({ S611 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_285_ (
  .in1({ S589, S583 }),
  .out1({ S612 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_286_ (
  .in1({ DP_ARU1_in1_6, DP_AC_out_0 }),
  .out1({ S613 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_105_ (
  .in1({ S613 }),
  .out1({ S614 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_235_ (
  .in1({ S547, S541 }),
  .out1({ S615 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_106_ (
  .in1({ S615 }),
  .out1({ S616 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_236_ (
  .in1({ S615, S613 }),
  .out1({ S617 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_287_ (
  .in1({ S616, S614 }),
  .out1({ S618 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_288_ (
  .in1({ S615, S613 }),
  .out1({ S619 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_107_ (
  .in1({ S619 }),
  .out1({ S620 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_237_ (
  .in1({ S620, S617 }),
  .out1({ S621 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_289_ (
  .in1({ S619, S618 }),
  .out1({ S622 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_238_ (
  .in1({ S578, S570 }),
  .out1({ S623 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_290_ (
  .in1({ S579, S571 }),
  .out1({ S624 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_291_ (
  .in1({ DP_ARU1_in1_5, DP_AC_out_1 }),
  .out1({ S625 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_292_ (
  .in1({ DP_ARU1_in1_4, DP_AC_out_3 }),
  .out1({ S626 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_239_ (
  .in1({ S540, S424 }),
  .out1({ S627 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_108_ (
  .in1({ S627 }),
  .out1({ S628 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_293_ (
  .in1({ S540, S424 }),
  .out1({ S629 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_294_ (
  .in1({ S629, S628 }),
  .out1({ S630 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_295_ (
  .in1({ S630, S625 }),
  .out1({ S631 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_109_ (
  .in1({ S631 }),
  .out1({ S632 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_240_ (
  .in1({ S630, S625 }),
  .out1({ S633 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_110_ (
  .in1({ S633 }),
  .out1({ S634 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_241_ (
  .in1({ S633, S632 }),
  .out1({ S635 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_296_ (
  .in1({ S634, S631 }),
  .out1({ S636 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_242_ (
  .in1({ S566, S558 }),
  .out1({ S637 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_297_ (
  .in1({ S567, S559 }),
  .out1({ S638 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_298_ (
  .in1({ DP_AC_out_4, DP_ARU1_in1_2 }),
  .out1({ S639 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_111_ (
  .in1({ S639 }),
  .out1({ S640 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_299_ (
  .in1({ DP_AC_out_6, DP_ARU1_in1_0 }),
  .out1({ S641 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_243_ (
  .in1({ S1107, S1009 }),
  .out1({ S642 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_300_ (
  .in1({ DP_AC_out_6, DP_ARU1_in1_1 }),
  .out1({ S643 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_244_ (
  .in1({ S643, S555 }),
  .out1({ S644 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_301_ (
  .in1({ S642, S556 }),
  .out1({ S645 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_302_ (
  .in1({ S641, S557 }),
  .out1({ S646 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_112_ (
  .in1({ S646 }),
  .out1({ S647 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_245_ (
  .in1({ S647, S644 }),
  .out1({ S648 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_303_ (
  .in1({ S646, S645 }),
  .out1({ S649 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_246_ (
  .in1({ S648, S640 }),
  .out1({ S650 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_304_ (
  .in1({ S649, S639 }),
  .out1({ S651 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_247_ (
  .in1({ S649, S639 }),
  .out1({ S652 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_305_ (
  .in1({ S648, S640 }),
  .out1({ S653 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_248_ (
  .in1({ S652, S650 }),
  .out1({ S654 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_306_ (
  .in1({ S653, S651 }),
  .out1({ S655 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_249_ (
  .in1({ S655, S637 }),
  .out1({ S656 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_307_ (
  .in1({ S654, S638 }),
  .out1({ S657 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_250_ (
  .in1({ S654, S638 }),
  .out1({ S658 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_308_ (
  .in1({ S655, S637 }),
  .out1({ S659 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_251_ (
  .in1({ S658, S656 }),
  .out1({ S660 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_309_ (
  .in1({ S659, S657 }),
  .out1({ S661 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_252_ (
  .in1({ S660, S635 }),
  .out1({ S662 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_310_ (
  .in1({ S661, S636 }),
  .out1({ S663 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_253_ (
  .in1({ S661, S636 }),
  .out1({ S664 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_311_ (
  .in1({ S660, S635 }),
  .out1({ S665 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_254_ (
  .in1({ S664, S662 }),
  .out1({ S666 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_312_ (
  .in1({ S665, S663 }),
  .out1({ S667 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_255_ (
  .in1({ S667, S623 }),
  .out1({ S668 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_313_ (
  .in1({ S666, S624 }),
  .out1({ S669 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_256_ (
  .in1({ S666, S624 }),
  .out1({ S670 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_314_ (
  .in1({ S667, S623 }),
  .out1({ S671 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_257_ (
  .in1({ S670, S668 }),
  .out1({ S672 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_315_ (
  .in1({ S671, S669 }),
  .out1({ S673 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_258_ (
  .in1({ S673, S622 }),
  .out1({ S674 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_316_ (
  .in1({ S672, S621 }),
  .out1({ S675 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_259_ (
  .in1({ S672, S621 }),
  .out1({ S676 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_317_ (
  .in1({ S673, S622 }),
  .out1({ S677 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_260_ (
  .in1({ S676, S674 }),
  .out1({ S678 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_318_ (
  .in1({ S677, S675 }),
  .out1({ S679 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_261_ (
  .in1({ S678, S612 }),
  .out1({ S680 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_319_ (
  .in1({ S679, S611 }),
  .out1({ S681 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_262_ (
  .in1({ S679, S611 }),
  .out1({ S682 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_320_ (
  .in1({ S678, S612 }),
  .out1({ S683 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_263_ (
  .in1({ S682, S680 }),
  .out1({ S684 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_321_ (
  .in1({ S683, S681 }),
  .out1({ S685 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_264_ (
  .in1({ S685, S595 }),
  .out1({ S686 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_322_ (
  .in1({ S684, S594 }),
  .out1({ S687 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_265_ (
  .in1({ S684, S594 }),
  .out1({ S688 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_323_ (
  .in1({ S685, S595 }),
  .out1({ S689 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_266_ (
  .in1({ S688, S686 }),
  .out1({ S690 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_324_ (
  .in1({ S689, S687 }),
  .out1({ S691 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_267_ (
  .in1({ S690, S600 }),
  .out1({ S692 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_268_ (
  .in1({ S691, S601 }),
  .out1({ S693 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_325_ (
  .in1({ S690, S600 }),
  .out1({ S694 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_269_ (
  .in1({ S693, S692 }),
  .out1({ S695 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_270_ (
  .in1({ S609, S988 }),
  .out1({ S696 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_326_ (
  .in1({ S696, S610 }),
  .out1({ S697 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_327_ (
  .in1({ S695, S988 }),
  .out1({ S698 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_328_ (
  .in1({ S698, S697 }),
  .out1({ S333 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_329_ (
  .in1({ S610, S607 }),
  .out1({ S699 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_271_ (
  .in1({ DP_ARU1_in1_7, DP_AC_out_7 }),
  .out1({ S700 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_272_ (
  .in1({ S1140, S1129 }),
  .out1({ S701 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_330_ (
  .in1({ DP_ARU1_in1_7, DP_AC_out_7 }),
  .out1({ S702 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_273_ (
  .in1({ S701, S700 }),
  .out1({ S703 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_331_ (
  .in1({ S703, S699 }),
  .out1({ S704 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_113_ (
  .in1({ S704 }),
  .out1({ S705 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_274_ (
  .in1({ S703, S699 }),
  .out1({ S706 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_275_ (
  .in1({ S706, S705 }),
  .out1({ S707 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_276_ (
  .in1({ S693, S686 }),
  .out1({ S708 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_332_ (
  .in1({ S694, S687 }),
  .out1({ S709 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_277_ (
  .in1({ S674, S668 }),
  .out1({ S710 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_333_ (
  .in1({ S675, S669 }),
  .out1({ S711 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_334_ (
  .in1({ DP_ARU1_in1_7, DP_AC_out_0 }),
  .out1({ S712 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_335_ (
  .in1({ DP_ARU1_in1_6, DP_AC_out_1 }),
  .out1({ S713 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_278_ (
  .in1({ S633, S627 }),
  .out1({ S714 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_279_ (
  .in1({ S714, S713 }),
  .out1({ S715 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_114_ (
  .in1({ S715 }),
  .out1({ S716 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_336_ (
  .in1({ S714, S713 }),
  .out1({ S717 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_337_ (
  .in1({ S717, S716 }),
  .out1({ S718 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_338_ (
  .in1({ S718, S712 }),
  .out1({ S719 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_115_ (
  .in1({ S719 }),
  .out1({ S720 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_280_ (
  .in1({ S718, S712 }),
  .out1({ S721 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_116_ (
  .in1({ S721 }),
  .out1({ S722 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_281_ (
  .in1({ S721, S720 }),
  .out1({ S723 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_339_ (
  .in1({ S722, S719 }),
  .out1({ S724 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_282_ (
  .in1({ S664, S656 }),
  .out1({ S725 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_340_ (
  .in1({ S665, S657 }),
  .out1({ S726 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_341_ (
  .in1({ DP_ARU1_in1_5, DP_AC_out_2 }),
  .out1({ S727 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_342_ (
  .in1({ DP_AC_out_4, DP_ARU1_in1_3 }),
  .out1({ S728 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_283_ (
  .in1({ S467, S424 }),
  .out1({ S729 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_117_ (
  .in1({ S729 }),
  .out1({ S730 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_343_ (
  .in1({ S728, S626 }),
  .out1({ S731 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_344_ (
  .in1({ S731, S730 }),
  .out1({ S732 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_345_ (
  .in1({ S732, S727 }),
  .out1({ S733 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_118_ (
  .in1({ S733 }),
  .out1({ S734 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_284_ (
  .in1({ S732, S727 }),
  .out1({ S735 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_119_ (
  .in1({ S735 }),
  .out1({ S736 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_285_ (
  .in1({ S735, S734 }),
  .out1({ S737 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_346_ (
  .in1({ S736, S733 }),
  .out1({ S738 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_286_ (
  .in1({ S652, S644 }),
  .out1({ S739 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_347_ (
  .in1({ S653, S645 }),
  .out1({ S740 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_348_ (
  .in1({ DP_AC_out_5, DP_ARU1_in1_2 }),
  .out1({ S741 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_120_ (
  .in1({ S741 }),
  .out1({ S742 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_349_ (
  .in1({ DP_AC_out_7, DP_ARU1_in1_0 }),
  .out1({ S743 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_350_ (
  .in1({ DP_AC_out_7, DP_ARU1_in1_1 }),
  .out1({ S744 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_287_ (
  .in1({ S744, S641 }),
  .out1({ S745 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_121_ (
  .in1({ S745 }),
  .out1({ S746 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_351_ (
  .in1({ S743, S643 }),
  .out1({ S747 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_122_ (
  .in1({ S747 }),
  .out1({ S748 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_288_ (
  .in1({ S748, S745 }),
  .out1({ S749 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_352_ (
  .in1({ S747, S746 }),
  .out1({ S750 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_289_ (
  .in1({ S749, S742 }),
  .out1({ S751 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_353_ (
  .in1({ S750, S741 }),
  .out1({ S752 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_290_ (
  .in1({ S750, S741 }),
  .out1({ S753 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_354_ (
  .in1({ S749, S742 }),
  .out1({ S754 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_291_ (
  .in1({ S753, S751 }),
  .out1({ S755 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_355_ (
  .in1({ S754, S752 }),
  .out1({ S756 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_292_ (
  .in1({ S756, S739 }),
  .out1({ S757 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_356_ (
  .in1({ S755, S740 }),
  .out1({ S758 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_293_ (
  .in1({ S755, S740 }),
  .out1({ S759 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_357_ (
  .in1({ S756, S739 }),
  .out1({ S760 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_294_ (
  .in1({ S759, S757 }),
  .out1({ S761 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_358_ (
  .in1({ S760, S758 }),
  .out1({ S762 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_295_ (
  .in1({ S761, S737 }),
  .out1({ S763 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_359_ (
  .in1({ S762, S738 }),
  .out1({ S764 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_296_ (
  .in1({ S762, S738 }),
  .out1({ S765 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_360_ (
  .in1({ S761, S737 }),
  .out1({ S766 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_297_ (
  .in1({ S765, S763 }),
  .out1({ S767 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_361_ (
  .in1({ S766, S764 }),
  .out1({ S768 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_298_ (
  .in1({ S768, S725 }),
  .out1({ S769 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_362_ (
  .in1({ S767, S726 }),
  .out1({ S770 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_299_ (
  .in1({ S767, S726 }),
  .out1({ S771 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_363_ (
  .in1({ S768, S725 }),
  .out1({ S772 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_300_ (
  .in1({ S771, S769 }),
  .out1({ S773 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_364_ (
  .in1({ S772, S770 }),
  .out1({ S774 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_301_ (
  .in1({ S773, S723 }),
  .out1({ S775 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_365_ (
  .in1({ S774, S724 }),
  .out1({ S776 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_302_ (
  .in1({ S774, S724 }),
  .out1({ S777 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_366_ (
  .in1({ S773, S723 }),
  .out1({ S778 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_303_ (
  .in1({ S777, S775 }),
  .out1({ S779 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_367_ (
  .in1({ S778, S776 }),
  .out1({ S780 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_304_ (
  .in1({ S780, S710 }),
  .out1({ S781 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_368_ (
  .in1({ S779, S711 }),
  .out1({ S782 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_305_ (
  .in1({ S779, S711 }),
  .out1({ S783 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_369_ (
  .in1({ S780, S710 }),
  .out1({ S784 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_306_ (
  .in1({ S783, S781 }),
  .out1({ S785 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_370_ (
  .in1({ S784, S782 }),
  .out1({ S786 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_307_ (
  .in1({ S785, S617 }),
  .out1({ S787 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_371_ (
  .in1({ S786, S618 }),
  .out1({ S788 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_308_ (
  .in1({ S786, S618 }),
  .out1({ S789 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_372_ (
  .in1({ S785, S617 }),
  .out1({ S790 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_309_ (
  .in1({ S789, S787 }),
  .out1({ S791 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_373_ (
  .in1({ S790, S788 }),
  .out1({ S792 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_310_ (
  .in1({ S792, S683 }),
  .out1({ S793 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_374_ (
  .in1({ S791, S682 }),
  .out1({ S794 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_311_ (
  .in1({ S791, S682 }),
  .out1({ S795 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_375_ (
  .in1({ S792, S683 }),
  .out1({ S796 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_312_ (
  .in1({ S795, S793 }),
  .out1({ S797 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_376_ (
  .in1({ S796, S794 }),
  .out1({ S798 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_313_ (
  .in1({ S798, S708 }),
  .out1({ S799 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_377_ (
  .in1({ S797, S709 }),
  .out1({ S800 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_314_ (
  .in1({ S797, S709 }),
  .out1({ S801 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_315_ (
  .in1({ S801, S799 }),
  .out1({ S802 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_316_ (
  .in1({ S802, CU_ADD }),
  .out1({ S803 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_317_ (
  .in1({ S707, S988 }),
  .out1({ S804 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_318_ (
  .in1({ S804, S803 }),
  .out1({ S334 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_319_ (
  .in1({ DP_ARU1_in1_8, DP_AC_out_8 }),
  .out1({ S805 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_378_ (
  .in1({ DP_ARU1_in1_8, DP_AC_out_8 }),
  .out1({ S806 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_123_ (
  .in1({ S806 }),
  .out1({ S807 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_320_ (
  .in1({ S807, S805 }),
  .out1({ S808 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_321_ (
  .in1({ S701, S699 }),
  .out1({ S809 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_322_ (
  .in1({ S809, S700 }),
  .out1({ S810 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_379_ (
  .in1({ S810, S808 }),
  .out1({ S811 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_323_ (
  .in1({ S810, S808 }),
  .out1({ S812 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_324_ (
  .in1({ S799, S793 }),
  .out1({ S813 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_380_ (
  .in1({ S800, S794 }),
  .out1({ S814 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_325_ (
  .in1({ S789, S781 }),
  .out1({ S815 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_381_ (
  .in1({ S790, S782 }),
  .out1({ S816 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_326_ (
  .in1({ S721, S715 }),
  .out1({ S817 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_327_ (
  .in1({ S777, S769 }),
  .out1({ S818 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_124_ (
  .in1({ S818 }),
  .out1({ S819 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_382_ (
  .in1({ DP_ARU1_in1_7, DP_AC_out_1 }),
  .out1({ S820 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_383_ (
  .in1({ DP_ARU1_in1_6, DP_AC_out_2 }),
  .out1({ S821 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_328_ (
  .in1({ S735, S729 }),
  .out1({ S822 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_329_ (
  .in1({ S822, S821 }),
  .out1({ S823 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_125_ (
  .in1({ S823 }),
  .out1({ S824 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_384_ (
  .in1({ S822, S821 }),
  .out1({ S825 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_385_ (
  .in1({ S825, S824 }),
  .out1({ S826 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_330_ (
  .in1({ S826, S820 }),
  .out1({ S827 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_126_ (
  .in1({ S827 }),
  .out1({ S828 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_386_ (
  .in1({ S826, S820 }),
  .out1({ S829 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_127_ (
  .in1({ S829 }),
  .out1({ S830 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_331_ (
  .in1({ S830, S827 }),
  .out1({ S831 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_387_ (
  .in1({ S829, S828 }),
  .out1({ S832 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_332_ (
  .in1({ S765, S757 }),
  .out1({ S833 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_388_ (
  .in1({ S766, S758 }),
  .out1({ S834 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_389_ (
  .in1({ DP_ARU1_in1_5, DP_AC_out_3 }),
  .out1({ S835 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_390_ (
  .in1({ DP_AC_out_5, DP_ARU1_in1_3 }),
  .out1({ S836 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_391_ (
  .in1({ DP_AC_out_5, DP_ARU1_in1_4 }),
  .out1({ S837 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_333_ (
  .in1({ S836, S467 }),
  .out1({ S838 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_128_ (
  .in1({ S838 }),
  .out1({ S839 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_392_ (
  .in1({ S836, S467 }),
  .out1({ S840 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_393_ (
  .in1({ S840, S839 }),
  .out1({ S841 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_394_ (
  .in1({ S841, S835 }),
  .out1({ S842 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_129_ (
  .in1({ S842 }),
  .out1({ S843 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_334_ (
  .in1({ S841, S835 }),
  .out1({ S844 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_130_ (
  .in1({ S844 }),
  .out1({ S845 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_335_ (
  .in1({ S844, S843 }),
  .out1({ S846 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_395_ (
  .in1({ S845, S842 }),
  .out1({ S847 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_336_ (
  .in1({ S753, S745 }),
  .out1({ S848 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_131_ (
  .in1({ S848 }),
  .out1({ S849 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_396_ (
  .in1({ DP_AC_out_6, DP_ARU1_in1_2 }),
  .out1({ S850 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_337_ (
  .in1({ S1129, S1031 }),
  .out1({ S851 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_397_ (
  .in1({ DP_AC_out_7, DP_ARU1_in1_2 }),
  .out1({ S852 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_338_ (
  .in1({ S852, S643 }),
  .out1({ S853 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_398_ (
  .in1({ S851, S642 }),
  .out1({ S854 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_399_ (
  .in1({ S850, S744 }),
  .out1({ S855 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_400_ (
  .in1({ S855, S854 }),
  .out1({ S856 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_132_ (
  .in1({ S856 }),
  .out1({ S857 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_339_ (
  .in1({ S856, S848 }),
  .out1({ S858 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_401_ (
  .in1({ S857, S849 }),
  .out1({ S859 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_402_ (
  .in1({ S856, S848 }),
  .out1({ S860 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_133_ (
  .in1({ S860 }),
  .out1({ S861 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_340_ (
  .in1({ S861, S858 }),
  .out1({ S862 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_403_ (
  .in1({ S860, S859 }),
  .out1({ S863 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_341_ (
  .in1({ S862, S846 }),
  .out1({ S864 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_404_ (
  .in1({ S863, S847 }),
  .out1({ S865 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_342_ (
  .in1({ S863, S847 }),
  .out1({ S866 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_405_ (
  .in1({ S862, S846 }),
  .out1({ S867 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_343_ (
  .in1({ S866, S864 }),
  .out1({ S868 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_406_ (
  .in1({ S867, S865 }),
  .out1({ S869 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_344_ (
  .in1({ S869, S833 }),
  .out1({ S870 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_407_ (
  .in1({ S868, S834 }),
  .out1({ S871 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_345_ (
  .in1({ S868, S834 }),
  .out1({ S872 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_408_ (
  .in1({ S869, S833 }),
  .out1({ S873 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_346_ (
  .in1({ S872, S870 }),
  .out1({ S874 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_409_ (
  .in1({ S873, S871 }),
  .out1({ S875 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_347_ (
  .in1({ S874, S831 }),
  .out1({ S876 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_410_ (
  .in1({ S875, S832 }),
  .out1({ S877 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_348_ (
  .in1({ S875, S832 }),
  .out1({ S878 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_411_ (
  .in1({ S874, S831 }),
  .out1({ S879 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_349_ (
  .in1({ S878, S876 }),
  .out1({ S880 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_412_ (
  .in1({ S879, S877 }),
  .out1({ S881 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_350_ (
  .in1({ S881, S818 }),
  .out1({ S882 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_413_ (
  .in1({ S880, S819 }),
  .out1({ S883 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_414_ (
  .in1({ S881, S818 }),
  .out1({ S884 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_415_ (
  .in1({ S884, S883 }),
  .out1({ S885 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_416_ (
  .in1({ S885, S817 }),
  .out1({ S886 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_134_ (
  .in1({ S886 }),
  .out1({ S887 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_351_ (
  .in1({ S885, S817 }),
  .out1({ S888 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_135_ (
  .in1({ S888 }),
  .out1({ S889 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_352_ (
  .in1({ S888, S887 }),
  .out1({ S890 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_417_ (
  .in1({ S889, S886 }),
  .out1({ S891 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_353_ (
  .in1({ S891, S815 }),
  .out1({ S892 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_418_ (
  .in1({ S890, S816 }),
  .out1({ S893 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_354_ (
  .in1({ S890, S816 }),
  .out1({ S894 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_419_ (
  .in1({ S891, S815 }),
  .out1({ S895 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_355_ (
  .in1({ S894, S892 }),
  .out1({ S896 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_420_ (
  .in1({ S895, S893 }),
  .out1({ S897 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_421_ (
  .in1({ S897, S813 }),
  .out1({ S898 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_356_ (
  .in1({ S897, S813 }),
  .out1({ S899 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_422_ (
  .in1({ S896, S814 }),
  .out1({ S900 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_423_ (
  .in1({ S900, S898 }),
  .out1({ S901 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_357_ (
  .in1({ S901, CU_ADD }),
  .out1({ S902 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_424_ (
  .in1({ S811, CU_ADD }),
  .out1({ S903 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_358_ (
  .in1({ S903, S812 }),
  .out1({ S904 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_359_ (
  .in1({ S904, S902 }),
  .out1({ S905 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_136_ (
  .in1({ S905 }),
  .out1({ S335 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_425_ (
  .in1({ S811, S806 }),
  .out1({ S906 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_426_ (
  .in1({ S1161, S1150 }),
  .out1({ S907 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_427_ (
  .in1({ DP_ARU1_in1_9, DP_AC_out_9 }),
  .out1({ S908 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_428_ (
  .in1({ S908, S907 }),
  .out1({ S909 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_429_ (
  .in1({ S909, S906 }),
  .out1({ S910 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_360_ (
  .in1({ S909, S906 }),
  .out1({ S911 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_137_ (
  .in1({ S911 }),
  .out1({ S912 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_430_ (
  .in1({ S912, S910 }),
  .out1({ S913 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_361_ (
  .in1({ S899, S892 }),
  .out1({ S914 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_431_ (
  .in1({ S900, S893 }),
  .out1({ S915 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_362_ (
  .in1({ S888, S882 }),
  .out1({ S916 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_138_ (
  .in1({ S916 }),
  .out1({ S917 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_363_ (
  .in1({ S827, S823 }),
  .out1({ S918 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_139_ (
  .in1({ S918 }),
  .out1({ S919 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_364_ (
  .in1({ S878, S870 }),
  .out1({ S920 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_432_ (
  .in1({ S879, S871 }),
  .out1({ S921 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_433_ (
  .in1({ DP_ARU1_in1_7, DP_AC_out_2 }),
  .out1({ S922 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_434_ (
  .in1({ DP_ARU1_in1_6, DP_AC_out_3 }),
  .out1({ S923 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_365_ (
  .in1({ S844, S838 }),
  .out1({ S924 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_366_ (
  .in1({ S924, S923 }),
  .out1({ S925 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_140_ (
  .in1({ S925 }),
  .out1({ S926 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_435_ (
  .in1({ S924, S923 }),
  .out1({ S927 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_436_ (
  .in1({ S927, S926 }),
  .out1({ S928 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_367_ (
  .in1({ S928, S922 }),
  .out1({ S929 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_141_ (
  .in1({ S929 }),
  .out1({ S930 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_437_ (
  .in1({ S928, S922 }),
  .out1({ S931 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_142_ (
  .in1({ S931 }),
  .out1({ S932 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_368_ (
  .in1({ S932, S929 }),
  .out1({ S933 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_438_ (
  .in1({ S931, S930 }),
  .out1({ S934 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_369_ (
  .in1({ S866, S858 }),
  .out1({ S935 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_439_ (
  .in1({ S867, S859 }),
  .out1({ S936 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_440_ (
  .in1({ DP_ARU1_in1_5, DP_AC_out_4 }),
  .out1({ S937 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_441_ (
  .in1({ DP_AC_out_6, DP_ARU1_in1_3 }),
  .out1({ S938 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_442_ (
  .in1({ DP_AC_out_6, DP_ARU1_in1_4 }),
  .out1({ S939 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_143_ (
  .in1({ S939 }),
  .out1({ S940 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_370_ (
  .in1({ S939, S836 }),
  .out1({ S941 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_144_ (
  .in1({ S941 }),
  .out1({ S942 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_443_ (
  .in1({ S938, S837 }),
  .out1({ S943 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_444_ (
  .in1({ S943, S942 }),
  .out1({ S944 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_445_ (
  .in1({ S944, S937 }),
  .out1({ S945 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_145_ (
  .in1({ S945 }),
  .out1({ S946 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_371_ (
  .in1({ S944, S937 }),
  .out1({ S947 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_146_ (
  .in1({ S947 }),
  .out1({ S948 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_372_ (
  .in1({ S947, S946 }),
  .out1({ S949 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_446_ (
  .in1({ S948, S945 }),
  .out1({ S950 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_373_ (
  .in1({ S852, S642 }),
  .out1({ S951 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_447_ (
  .in1({ S851, S643 }),
  .out1({ S952 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_374_ (
  .in1({ S951, S949 }),
  .out1({ S953 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_448_ (
  .in1({ S952, S950 }),
  .out1({ S954 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_375_ (
  .in1({ S952, S950 }),
  .out1({ S955 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_449_ (
  .in1({ S951, S949 }),
  .out1({ S956 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_376_ (
  .in1({ S955, S953 }),
  .out1({ S957 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_450_ (
  .in1({ S956, S954 }),
  .out1({ S958 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_377_ (
  .in1({ S958, S935 }),
  .out1({ S959 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_451_ (
  .in1({ S957, S936 }),
  .out1({ S960 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_378_ (
  .in1({ S957, S936 }),
  .out1({ S961 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_452_ (
  .in1({ S958, S935 }),
  .out1({ S962 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_379_ (
  .in1({ S961, S959 }),
  .out1({ S963 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_453_ (
  .in1({ S962, S960 }),
  .out1({ S964 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_380_ (
  .in1({ S963, S933 }),
  .out1({ S965 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_454_ (
  .in1({ S964, S934 }),
  .out1({ S967 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_381_ (
  .in1({ S964, S934 }),
  .out1({ S968 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_455_ (
  .in1({ S963, S933 }),
  .out1({ S969 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_382_ (
  .in1({ S968, S965 }),
  .out1({ S970 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_456_ (
  .in1({ S969, S967 }),
  .out1({ S971 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_457_ (
  .in1({ S970, S921 }),
  .out1({ S972 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_458_ (
  .in1({ S971, S920 }),
  .out1({ S973 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_459_ (
  .in1({ S973, S972 }),
  .out1({ S974 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_147_ (
  .in1({ S974 }),
  .out1({ S975 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_460_ (
  .in1({ S975, S919 }),
  .out1({ S976 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_461_ (
  .in1({ S974, S918 }),
  .out1({ S978 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_462_ (
  .in1({ S978, S976 }),
  .out1({ S979 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_148_ (
  .in1({ S979 }),
  .out1({ S980 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_463_ (
  .in1({ S979, S916 }),
  .out1({ S981 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_464_ (
  .in1({ S980, S917 }),
  .out1({ S982 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_149_ (
  .in1({ S982 }),
  .out1({ S983 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_465_ (
  .in1({ S982, S981 }),
  .out1({ S984 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_150_ (
  .in1({ S984 }),
  .out1({ S985 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_383_ (
  .in1({ S985, S915 }),
  .out1({ S986 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_384_ (
  .in1({ S984, S914 }),
  .out1({ S987 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_466_ (
  .in1({ S985, S915 }),
  .out1({ S989 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_385_ (
  .in1({ S987, S986 }),
  .out1({ S990 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_386_ (
  .in1({ S990, CU_ADD }),
  .out1({ S991 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_387_ (
  .in1({ S913, S988 }),
  .out1({ S992 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_388_ (
  .in1({ S992, S991 }),
  .out1({ S336 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_389_ (
  .in1({ DP_ARU1_in1_10, DP_AC_out_10 }),
  .out1({ S993 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_467_ (
  .in1({ DP_ARU1_in1_10, DP_AC_out_10 }),
  .out1({ S994 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_151_ (
  .in1({ S994 }),
  .out1({ S995 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_390_ (
  .in1({ S995, S993 }),
  .out1({ S996 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_152_ (
  .in1({ S996 }),
  .out1({ S997 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_468_ (
  .in1({ S907, S906 }),
  .out1({ S999 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_469_ (
  .in1({ S999, S908 }),
  .out1({ S1000 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_153_ (
  .in1({ S1000 }),
  .out1({ S1001 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_391_ (
  .in1({ S1000, S996 }),
  .out1({ S1002 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_392_ (
  .in1({ S1001, S997 }),
  .out1({ S1003 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_154_ (
  .in1({ S1003 }),
  .out1({ S1004 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_393_ (
  .in1({ S1003, S1002 }),
  .out1({ S1005 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_394_ (
  .in1({ S1005, S988 }),
  .out1({ S1006 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_395_ (
  .in1({ S987, S983 }),
  .out1({ S1007 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_470_ (
  .in1({ S989, S982 }),
  .out1({ S1008 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_471_ (
  .in1({ S976, S972 }),
  .out1({ S1010 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_155_ (
  .in1({ S1010 }),
  .out1({ S1011 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_396_ (
  .in1({ S929, S925 }),
  .out1({ S1012 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_397_ (
  .in1({ S968, S959 }),
  .out1({ S1013 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_472_ (
  .in1({ DP_ARU1_in1_7, DP_AC_out_3 }),
  .out1({ S1014 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_473_ (
  .in1({ DP_ARU1_in1_6, DP_AC_out_4 }),
  .out1({ S1015 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_398_ (
  .in1({ S947, S941 }),
  .out1({ S1016 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_399_ (
  .in1({ S1016, S1015 }),
  .out1({ S1017 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_156_ (
  .in1({ S1017 }),
  .out1({ S1018 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_474_ (
  .in1({ S1016, S1015 }),
  .out1({ S1019 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_475_ (
  .in1({ S1019, S1018 }),
  .out1({ S1021 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_400_ (
  .in1({ S1021, S1014 }),
  .out1({ S1022 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_157_ (
  .in1({ S1022 }),
  .out1({ S1023 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_476_ (
  .in1({ S1021, S1014 }),
  .out1({ S1024 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_158_ (
  .in1({ S1024 }),
  .out1({ S1025 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_401_ (
  .in1({ S1025, S1022 }),
  .out1({ S1026 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_477_ (
  .in1({ S1024, S1023 }),
  .out1({ S1027 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_402_ (
  .in1({ S955, S853 }),
  .out1({ S1028 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_478_ (
  .in1({ S956, S854 }),
  .out1({ S1029 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_479_ (
  .in1({ DP_AC_out_7, DP_ARU1_in1_3 }),
  .out1({ S1030 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_480_ (
  .in1({ S1030, S939 }),
  .out1({ S1032 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_159_ (
  .in1({ S1032 }),
  .out1({ S1033 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_481_ (
  .in1({ DP_AC_out_7, DP_ARU1_in1_4 }),
  .out1({ S1034 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_403_ (
  .in1({ S1034, S938 }),
  .out1({ S1035 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_160_ (
  .in1({ S1035 }),
  .out1({ S1036 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_404_ (
  .in1({ S1035, S1033 }),
  .out1({ S1037 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_482_ (
  .in1({ S1036, S1032 }),
  .out1({ S1038 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_405_ (
  .in1({ S1037, S528 }),
  .out1({ S1039 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_483_ (
  .in1({ S1038, S529 }),
  .out1({ S1040 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_406_ (
  .in1({ S1038, S529 }),
  .out1({ S1041 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_161_ (
  .in1({ S1041 }),
  .out1({ S1043 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_407_ (
  .in1({ S1041, S1039 }),
  .out1({ S1044 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_484_ (
  .in1({ S1043, S1040 }),
  .out1({ S1045 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_408_ (
  .in1({ S1045, S1028 }),
  .out1({ S1046 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_485_ (
  .in1({ S1044, S1029 }),
  .out1({ S1047 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_409_ (
  .in1({ S1044, S1029 }),
  .out1({ S1048 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_486_ (
  .in1({ S1045, S1028 }),
  .out1({ S1049 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_410_ (
  .in1({ S1048, S1046 }),
  .out1({ S1050 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_487_ (
  .in1({ S1049, S1047 }),
  .out1({ S1051 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_488_ (
  .in1({ S1051, S1027 }),
  .out1({ S1052 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_411_ (
  .in1({ S1051, S1027 }),
  .out1({ S1054 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_489_ (
  .in1({ S1050, S1026 }),
  .out1({ S1055 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_490_ (
  .in1({ S1055, S1052 }),
  .out1({ S1056 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_412_ (
  .in1({ S1056, S1013 }),
  .out1({ S1057 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_162_ (
  .in1({ S1057 }),
  .out1({ S1058 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_491_ (
  .in1({ S1056, S1013 }),
  .out1({ S1059 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_492_ (
  .in1({ S1059, S1058 }),
  .out1({ S1060 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_493_ (
  .in1({ S1060, S1012 }),
  .out1({ S1061 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_163_ (
  .in1({ S1061 }),
  .out1({ S1062 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_413_ (
  .in1({ S1060, S1012 }),
  .out1({ S1063 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_414_ (
  .in1({ S1063, S1062 }),
  .out1({ S1065 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_164_ (
  .in1({ S1065 }),
  .out1({ S1066 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_415_ (
  .in1({ S1066, S1011 }),
  .out1({ S1067 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_165_ (
  .in1({ S1067 }),
  .out1({ S1068 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_416_ (
  .in1({ S1065, S1010 }),
  .out1({ S1069 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_417_ (
  .in1({ S1069, S1067 }),
  .out1({ S1070 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_166_ (
  .in1({ S1070 }),
  .out1({ S1071 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_418_ (
  .in1({ S1070, S1008 }),
  .out1({ S1072 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_419_ (
  .in1({ S1071, S1007 }),
  .out1({ S1073 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_494_ (
  .in1({ S1070, S1008 }),
  .out1({ S1074 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_420_ (
  .in1({ S1073, S1072 }),
  .out1({ S1076 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_421_ (
  .in1({ S1076, CU_ADD }),
  .out1({ S1077 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_422_ (
  .in1({ S1077, S1006 }),
  .out1({ S322 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_495_ (
  .in1({ S1004, S994 }),
  .out1({ S1078 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_496_ (
  .in1({ S1183, S1172 }),
  .out1({ S1079 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_497_ (
  .in1({ DP_ARU1_in1_11, DP_AC_out_11 }),
  .out1({ S1080 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_498_ (
  .in1({ S1080, S1079 }),
  .out1({ S1081 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_499_ (
  .in1({ S1081, S1078 }),
  .out1({ S1082 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_423_ (
  .in1({ S1081, S1078 }),
  .out1({ S1083 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_167_ (
  .in1({ S1083 }),
  .out1({ S1084 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_500_ (
  .in1({ S1084, S1082 }),
  .out1({ S1086 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_424_ (
  .in1({ S1073, S1067 }),
  .out1({ S1087 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_501_ (
  .in1({ S1074, S1068 }),
  .out1({ S1088 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_425_ (
  .in1({ S1063, S1057 }),
  .out1({ S1089 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_168_ (
  .in1({ S1089 }),
  .out1({ S1090 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_426_ (
  .in1({ S1022, S1017 }),
  .out1({ S1091 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_169_ (
  .in1({ S1091 }),
  .out1({ S1092 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_427_ (
  .in1({ S1054, S1046 }),
  .out1({ S1093 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_502_ (
  .in1({ S1055, S1047 }),
  .out1({ S1094 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_503_ (
  .in1({ DP_ARU1_in1_7, DP_AC_out_4 }),
  .out1({ S1095 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_504_ (
  .in1({ DP_ARU1_in1_6, DP_AC_out_5 }),
  .out1({ S1097 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_428_ (
  .in1({ S1041, S1035 }),
  .out1({ S1098 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_429_ (
  .in1({ S1098, S1097 }),
  .out1({ S1099 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_170_ (
  .in1({ S1099 }),
  .out1({ S1100 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_505_ (
  .in1({ S1098, S1097 }),
  .out1({ S1101 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_506_ (
  .in1({ S1101, S1100 }),
  .out1({ S1102 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_430_ (
  .in1({ S1102, S1095 }),
  .out1({ S1103 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_171_ (
  .in1({ S1103 }),
  .out1({ S1104 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_507_ (
  .in1({ S1102, S1095 }),
  .out1({ S1105 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_172_ (
  .in1({ S1105 }),
  .out1({ S1106 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_431_ (
  .in1({ S1106, S1103 }),
  .out1({ S1108 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_508_ (
  .in1({ S1105, S1104 }),
  .out1({ S1109 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_509_ (
  .in1({ DP_AC_out_6, DP_ARU1_in1_5 }),
  .out1({ S1110 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_510_ (
  .in1({ S1110, S1034 }),
  .out1({ S1111 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_173_ (
  .in1({ S1111 }),
  .out1({ S1112 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_432_ (
  .in1({ S1129, S1096 }),
  .out1({ S1113 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_511_ (
  .in1({ DP_AC_out_7, DP_ARU1_in1_5 }),
  .out1({ S1114 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_433_ (
  .in1({ S1114, S939 }),
  .out1({ S1115 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_512_ (
  .in1({ S1113, S940 }),
  .out1({ S1116 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_434_ (
  .in1({ S1115, S1112 }),
  .out1({ S1117 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_513_ (
  .in1({ S1116, S1111 }),
  .out1({ S1119 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_514_ (
  .in1({ S1119, S1109 }),
  .out1({ S1120 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_435_ (
  .in1({ S1119, S1109 }),
  .out1({ S1121 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_515_ (
  .in1({ S1117, S1108 }),
  .out1({ S1122 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_516_ (
  .in1({ S1122, S1120 }),
  .out1({ S1123 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_174_ (
  .in1({ S1123 }),
  .out1({ S1124 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_517_ (
  .in1({ S1124, S1094 }),
  .out1({ S1125 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_518_ (
  .in1({ S1123, S1093 }),
  .out1({ S1126 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_519_ (
  .in1({ S1126, S1125 }),
  .out1({ S1127 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_175_ (
  .in1({ S1127 }),
  .out1({ S1128 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_520_ (
  .in1({ S1127, S1091 }),
  .out1({ S1130 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_521_ (
  .in1({ S1128, S1092 }),
  .out1({ S1131 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_522_ (
  .in1({ S1131, S1130 }),
  .out1({ S1132 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_176_ (
  .in1({ S1132 }),
  .out1({ S1133 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_523_ (
  .in1({ S1133, S1090 }),
  .out1({ S1134 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_177_ (
  .in1({ S1134 }),
  .out1({ S1135 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_524_ (
  .in1({ S1132, S1089 }),
  .out1({ S1136 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_525_ (
  .in1({ S1136, S1134 }),
  .out1({ S1137 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_178_ (
  .in1({ S1137 }),
  .out1({ S1138 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_436_ (
  .in1({ S1138, S1088 }),
  .out1({ S1139 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_437_ (
  .in1({ S1137, S1087 }),
  .out1({ S1141 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_526_ (
  .in1({ S1138, S1088 }),
  .out1({ S1142 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_438_ (
  .in1({ S1141, S1139 }),
  .out1({ S1143 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_439_ (
  .in1({ S1143, CU_ADD }),
  .out1({ S1144 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_440_ (
  .in1({ S1086, S988 }),
  .out1({ S1145 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_441_ (
  .in1({ S1145, S1144 }),
  .out1({ S323 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_442_ (
  .in1({ DP_ARU1_in1_12, DP_AC_out_12 }),
  .out1({ S1146 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_527_ (
  .in1({ DP_ARU1_in1_12, DP_AC_out_12 }),
  .out1({ S1147 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_179_ (
  .in1({ S1147 }),
  .out1({ S1148 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_443_ (
  .in1({ S1148, S1146 }),
  .out1({ S1149 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_528_ (
  .in1({ S1079, S1078 }),
  .out1({ S1151 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_529_ (
  .in1({ S1151, S1080 }),
  .out1({ S1152 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_530_ (
  .in1({ S1152, S1149 }),
  .out1({ S1153 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_444_ (
  .in1({ S1152, S1149 }),
  .out1({ S1154 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_445_ (
  .in1({ S1141, S1135 }),
  .out1({ S1155 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_531_ (
  .in1({ S1142, S1134 }),
  .out1({ S1156 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_532_ (
  .in1({ S1131, S1125 }),
  .out1({ S1157 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_180_ (
  .in1({ S1157 }),
  .out1({ S1158 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_446_ (
  .in1({ S1103, S1099 }),
  .out1({ S1159 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_533_ (
  .in1({ DP_ARU1_in1_7, DP_AC_out_5 }),
  .out1({ S1160 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_181_ (
  .in1({ S1160 }),
  .out1({ S1162 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_534_ (
  .in1({ S1115, DP_ARU1_in1_6 }),
  .out1({ S1163 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_182_ (
  .in1({ S1163 }),
  .out1({ S1164 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_535_ (
  .in1({ S1116, S607 }),
  .out1({ S1165 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_536_ (
  .in1({ S1165, S1163 }),
  .out1({ S1166 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_183_ (
  .in1({ S1166 }),
  .out1({ S1167 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_447_ (
  .in1({ S1166, S1160 }),
  .out1({ S1168 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_537_ (
  .in1({ S1167, S1162 }),
  .out1({ S1169 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_538_ (
  .in1({ S1166, S1160 }),
  .out1({ S1170 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_184_ (
  .in1({ S1170 }),
  .out1({ S1171 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_448_ (
  .in1({ S1171, S1168 }),
  .out1({ S1173 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_539_ (
  .in1({ S1170, S1169 }),
  .out1({ S1174 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_540_ (
  .in1({ S1174, S1114 }),
  .out1({ S1175 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_449_ (
  .in1({ S1174, S1114 }),
  .out1({ S1176 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_541_ (
  .in1({ S1173, S1113 }),
  .out1({ S1177 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_542_ (
  .in1({ S1177, S1175 }),
  .out1({ S1178 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_185_ (
  .in1({ S1178 }),
  .out1({ S1179 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_543_ (
  .in1({ S1179, S1121 }),
  .out1({ S1180 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_186_ (
  .in1({ S1180 }),
  .out1({ S1181 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_544_ (
  .in1({ S1178, S1122 }),
  .out1({ S1182 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_545_ (
  .in1({ S1182, S1180 }),
  .out1({ S1184 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_450_ (
  .in1({ S1184, S1159 }),
  .out1({ S1185 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_187_ (
  .in1({ S1185 }),
  .out1({ S1186 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_546_ (
  .in1({ S1184, S1159 }),
  .out1({ S1187 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_188_ (
  .in1({ S1187 }),
  .out1({ S1188 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_451_ (
  .in1({ S1188, S1185 }),
  .out1({ S1189 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_189_ (
  .in1({ S1189 }),
  .out1({ S1190 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_452_ (
  .in1({ S1190, S1158 }),
  .out1({ S1191 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_190_ (
  .in1({ S1191 }),
  .out1({ S1192 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_453_ (
  .in1({ S1189, S1157 }),
  .out1({ S1193 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_454_ (
  .in1({ S1193, S1191 }),
  .out1({ S1195 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_191_ (
  .in1({ S1195 }),
  .out1({ S1196 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_547_ (
  .in1({ S1196, S1155 }),
  .out1({ S1197 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_192_ (
  .in1({ S1197 }),
  .out1({ S1198 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_455_ (
  .in1({ S1196, S1155 }),
  .out1({ S1199 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_548_ (
  .in1({ S1195, S1156 }),
  .out1({ S1200 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_456_ (
  .in1({ S1199, S1198 }),
  .out1({ S1201 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_457_ (
  .in1({ S1154, S988 }),
  .out1({ S1202 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_549_ (
  .in1({ S1202, S1153 }),
  .out1({ S1203 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_550_ (
  .in1({ S1201, S988 }),
  .out1({ S1204 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_551_ (
  .in1({ S1204, S1203 }),
  .out1({ S324 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_552_ (
  .in1({ S1153, S1147 }),
  .out1({ S1206 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_553_ (
  .in1({ S1205, S1194 }),
  .out1({ S1207 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_554_ (
  .in1({ DP_ARU1_in1_13, DP_AC_out_13 }),
  .out1({ S1208 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_555_ (
  .in1({ S1208, S1207 }),
  .out1({ S1209 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_556_ (
  .in1({ S1209, S1206 }),
  .out1({ S1210 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_458_ (
  .in1({ S1209, S1206 }),
  .out1({ S1211 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_459_ (
  .in1({ S1199, S1191 }),
  .out1({ S1212 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_557_ (
  .in1({ S1200, S1192 }),
  .out1({ S1213 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_460_ (
  .in1({ S1185, S1181 }),
  .out1({ S1214 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_558_ (
  .in1({ S1186, S1180 }),
  .out1({ S1216 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_461_ (
  .in1({ S1168, S1164 }),
  .out1({ S1217 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_559_ (
  .in1({ S1169, S1163 }),
  .out1({ S1218 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_560_ (
  .in1({ DP_ARU1_in1_7, DP_AC_out_6 }),
  .out1({ S1219 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_561_ (
  .in1({ DP_AC_out_7, DP_ARU1_in1_6 }),
  .out1({ S1220 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_562_ (
  .in1({ S1220, S1219 }),
  .out1({ S1221 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_193_ (
  .in1({ S1221 }),
  .out1({ S1222 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_462_ (
  .in1({ S702, S607 }),
  .out1({ S1223 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_563_ (
  .in1({ S701, S606 }),
  .out1({ S1224 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_463_ (
  .in1({ S1223, S1222 }),
  .out1({ S1225 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_564_ (
  .in1({ S1224, S1221 }),
  .out1({ S1227 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_464_ (
  .in1({ S1227, S1177 }),
  .out1({ S1228 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_565_ (
  .in1({ S1225, S1176 }),
  .out1({ S1229 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_465_ (
  .in1({ S1225, S1176 }),
  .out1({ S1230 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_566_ (
  .in1({ S1227, S1177 }),
  .out1({ S1231 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_466_ (
  .in1({ S1230, S1228 }),
  .out1({ S1232 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_567_ (
  .in1({ S1231, S1229 }),
  .out1({ S1233 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_467_ (
  .in1({ S1233, S1217 }),
  .out1({ S1234 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_568_ (
  .in1({ S1232, S1218 }),
  .out1({ S1235 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_468_ (
  .in1({ S1232, S1218 }),
  .out1({ S1236 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_569_ (
  .in1({ S1233, S1217 }),
  .out1({ S1238 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_469_ (
  .in1({ S1236, S1234 }),
  .out1({ S1239 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_570_ (
  .in1({ S1238, S1235 }),
  .out1({ S1240 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_470_ (
  .in1({ S1240, S1214 }),
  .out1({ S1241 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_471_ (
  .in1({ S1239, S1216 }),
  .out1({ S1242 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_472_ (
  .in1({ S1242, S1241 }),
  .out1({ S1243 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_473_ (
  .in1({ S1243, S1212 }),
  .out1({ S1244 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_571_ (
  .in1({ S1243, S1212 }),
  .out1({ S1245 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_572_ (
  .in1({ S1210, CU_ADD }),
  .out1({ S1246 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_474_ (
  .in1({ S1246, S1211 }),
  .out1({ S1247 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_573_ (
  .in1({ S1245, S988 }),
  .out1({ S1249 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_475_ (
  .in1({ S1249, S1244 }),
  .out1({ S1250 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_476_ (
  .in1({ S1250, S1247 }),
  .out1({ S325 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_477_ (
  .in1({ S1234, S1228 }),
  .out1({ S1251 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_574_ (
  .in1({ S1235, S1229 }),
  .out1({ S1252 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_478_ (
  .in1({ S702, S606 }),
  .out1({ S1253 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_575_ (
  .in1({ S701, S607 }),
  .out1({ S1254 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_576_ (
  .in1({ S1253, S1252 }),
  .out1({ S1255 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_577_ (
  .in1({ S1254, S1251 }),
  .out1({ S1256 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_578_ (
  .in1({ S1256, S1255 }),
  .out1({ S1257 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_194_ (
  .in1({ S1257 }),
  .out1({ S1259 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_479_ (
  .in1({ S1242, S1212 }),
  .out1({ S1260 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_480_ (
  .in1({ S1241, S1213 }),
  .out1({ S1261 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_481_ (
  .in1({ S1260, S1241 }),
  .out1({ S1262 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_482_ (
  .in1({ S1261, S1242 }),
  .out1({ S1263 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_579_ (
  .in1({ S1262, S1257 }),
  .out1({ S1264 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_483_ (
  .in1({ S1262, S1257 }),
  .out1({ S1265 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_580_ (
  .in1({ S1263, S1259 }),
  .out1({ S1266 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_484_ (
  .in1({ S1265, CU_ADD }),
  .out1({ S1267 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_581_ (
  .in1({ S1266, S988 }),
  .out1({ S1268 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_582_ (
  .in1({ S1267, S1264 }),
  .out1({ S338 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_485_ (
  .in1({ DP_ARU1_in1_14, DP_AC_out_14 }),
  .out1({ S339 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_486_ (
  .in1({ S1226, S1215 }),
  .out1({ S340 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_487_ (
  .in1({ S340, S339 }),
  .out1({ S341 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_583_ (
  .in1({ S1207, S1206 }),
  .out1({ S342 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_584_ (
  .in1({ S342, S1208 }),
  .out1({ S343 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_488_ (
  .in1({ S343, S341 }),
  .out1({ S344 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_585_ (
  .in1({ S343, S341 }),
  .out1({ S345 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_195_ (
  .in1({ S345 }),
  .out1({ S346 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_489_ (
  .in1({ S344, S988 }),
  .out1({ S347 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_586_ (
  .in1({ S347, S345 }),
  .out1({ S349 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_587_ (
  .in1({ S349, S338 }),
  .out1({ S326 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_588_ (
  .in1({ S1255, S1224 }),
  .out1({ S350 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_490_ (
  .in1({ S350, S1268 }),
  .out1({ S351 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_491_ (
  .in1({ S346, S340 }),
  .out1({ S352 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_492_ (
  .in1({ S371, S368 }),
  .out1({ S353 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_493_ (
  .in1({ S353, S352 }),
  .out1({ S354 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_589_ (
  .in1({ S353, S352 }),
  .out1({ S355 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_590_ (
  .in1({ S355, CU_ADD }),
  .out1({ S356 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_494_ (
  .in1({ S356, S354 }),
  .out1({ S357 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_495_ (
  .in1({ S357, S351 }),
  .out1({ S327 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_496_ (
  .in1({ CU_MUL, CU_ADD }),
  .out1({ S337 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_591_ (
  .in1({ S355, S370 }),
  .out1({ S1270 })
);
$_DLATCH_P_ #() 
$_DLATCH_P__1_ (
  .D({ S1270 }),
  .E({ CU_ADD }),
  .Q({ DP_ARU1_C })
);
$_DLATCH_N_ #() 
$_DLATCH_N__3_ (
  .D({ S321 }),
  .E({ S337 }),
  .Q({ DP_ARU1_out_0 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__4_ (
  .D({ S328 }),
  .E({ S337 }),
  .Q({ DP_ARU1_out_1 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__5_ (
  .D({ S329 }),
  .E({ S337 }),
  .Q({ DP_ARU1_out_2 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__6_ (
  .D({ S330 }),
  .E({ S337 }),
  .Q({ DP_ARU1_out_3 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__7_ (
  .D({ S331 }),
  .E({ S337 }),
  .Q({ DP_ARU1_out_4 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__8_ (
  .D({ S332 }),
  .E({ S337 }),
  .Q({ DP_ARU1_out_5 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__9_ (
  .D({ S333 }),
  .E({ S337 }),
  .Q({ DP_ARU1_out_6 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__10_ (
  .D({ S334 }),
  .E({ S337 }),
  .Q({ DP_ARU1_out_7 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__11_ (
  .D({ S335 }),
  .E({ S337 }),
  .Q({ DP_ARU1_out_8 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__12_ (
  .D({ S336 }),
  .E({ S337 }),
  .Q({ DP_ARU1_out_9 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__13_ (
  .D({ S322 }),
  .E({ S337 }),
  .Q({ DP_ARU1_out_10 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__14_ (
  .D({ S323 }),
  .E({ S337 }),
  .Q({ DP_ARU1_out_11 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__15_ (
  .D({ S324 }),
  .E({ S337 }),
  .Q({ DP_ARU1_out_12 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__16_ (
  .D({ S325 }),
  .E({ S337 }),
  .Q({ DP_ARU1_out_13 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__17_ (
  .D({ S326 }),
  .E({ S337 }),
  .Q({ DP_ARU1_out_14 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__18_ (
  .D({ S327 }),
  .E({ S337 }),
  .Q({ DP_ARU1_N })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_196_ (
  .in1({ CU_inst_0 }),
  .out1({ S1290 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_197_ (
  .in1({ CU_LSB0E }),
  .out1({ S1291 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_198_ (
  .in1({ CU_conOF }),
  .out1({ S1292 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_199_ (
  .in1({ CU_inst_1 }),
  .out1({ S1293 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_200_ (
  .in1({ CU_inst_2 }),
  .out1({ S1294 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_201_ (
  .in1({ CU_inst_3 }),
  .out1({ S1295 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_202_ (
  .in1({ CU_inst_4 }),
  .out1({ S1296 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_203_ (
  .in1({ CU_SE12bits }),
  .out1({ S1297 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_497_ (
  .in1({ CU_conOF, S1291 }),
  .out1({ S1298 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_498_ (
  .in1({ S1298, S1290 }),
  .out1({ S1271 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_499_ (
  .in1({ S1298, S1293 }),
  .out1({ S1278 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_500_ (
  .in1({ S1298, S1294 }),
  .out1({ S1279 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_501_ (
  .in1({ S1298, S1295 }),
  .out1({ S1280 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_592_ (
  .in1({ S1292, S1291 }),
  .out1({ S1299 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_593_ (
  .in1({ CU_SE12bits, CU_inst_3 }),
  .out1({ S1300 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_594_ (
  .in1({ CU_SE12bits, S1292 }),
  .out1({ S1301 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_502_ (
  .in1({ S1300, S1299 }),
  .out1({ S1302 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_204_ (
  .in1({ S1302 }),
  .out1({ S1303 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_503_ (
  .in1({ S1298, S1296 }),
  .out1({ S1304 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_595_ (
  .in1({ S1304, S1301 }),
  .out1({ S1305 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_596_ (
  .in1({ S1305, S1303 }),
  .out1({ S1281 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_504_ (
  .in1({ S1299, CU_SE12bits }),
  .out1({ S1306 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_205_ (
  .in1({ S1306 }),
  .out1({ S1307 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_597_ (
  .in1({ S1306, CU_inst_5 }),
  .out1({ S1308 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_598_ (
  .in1({ CU_inst_5, CU_conOF }),
  .out1({ S1309 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_206_ (
  .in1({ S1309 }),
  .out1({ S1310 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_505_ (
  .in1({ S1310, S1302 }),
  .out1({ S1311 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_599_ (
  .in1({ S1311, S1308 }),
  .out1({ S1282 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_600_ (
  .in1({ S1306, CU_inst_6 }),
  .out1({ S1312 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_601_ (
  .in1({ CU_inst_6, CU_conOF }),
  .out1({ S1313 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_207_ (
  .in1({ S1313 }),
  .out1({ S1314 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_506_ (
  .in1({ S1314, S1302 }),
  .out1({ S1315 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_602_ (
  .in1({ S1315, S1312 }),
  .out1({ S1283 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_603_ (
  .in1({ S1306, CU_inst_7 }),
  .out1({ S1316 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_604_ (
  .in1({ CU_inst_7, CU_conOF }),
  .out1({ S1317 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_208_ (
  .in1({ S1317 }),
  .out1({ S1318 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_507_ (
  .in1({ S1318, S1302 }),
  .out1({ S1319 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_605_ (
  .in1({ S1319, S1316 }),
  .out1({ S1284 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_606_ (
  .in1({ S1306, CU_inst_8 }),
  .out1({ S1320 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_607_ (
  .in1({ CU_inst_8, CU_conOF }),
  .out1({ S1321 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_209_ (
  .in1({ S1321 }),
  .out1({ S1322 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_508_ (
  .in1({ S1322, S1302 }),
  .out1({ S1323 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_608_ (
  .in1({ S1323, S1320 }),
  .out1({ S1285 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_609_ (
  .in1({ S1306, CU_inst_9 }),
  .out1({ S1324 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_610_ (
  .in1({ CU_inst_9, CU_conOF }),
  .out1({ S1325 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_210_ (
  .in1({ S1325 }),
  .out1({ S1326 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_509_ (
  .in1({ S1326, S1302 }),
  .out1({ S1327 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_611_ (
  .in1({ S1327, S1324 }),
  .out1({ S1286 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_612_ (
  .in1({ S1306, CU_inst_10 }),
  .out1({ S1328 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_613_ (
  .in1({ CU_inst_10, CU_conOF }),
  .out1({ S1329 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_211_ (
  .in1({ S1329 }),
  .out1({ S1330 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_510_ (
  .in1({ S1330, S1302 }),
  .out1({ S1331 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_614_ (
  .in1({ S1331, S1328 }),
  .out1({ S1272 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_615_ (
  .in1({ CU_inst_11, CU_conOF }),
  .out1({ S1332 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_616_ (
  .in1({ CU_inst_11, S1297 }),
  .out1({ S1333 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_511_ (
  .in1({ S1333, S1299 }),
  .out1({ S1334 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_512_ (
  .in1({ S1334, S1302 }),
  .out1({ S1335 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_617_ (
  .in1({ S1335, S1332 }),
  .out1({ S1273 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_618_ (
  .in1({ S1299, DP_IMM1_in1_0 }),
  .out1({ S1336 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_619_ (
  .in1({ S1336, S1335 }),
  .out1({ S1274 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_620_ (
  .in1({ S1299, DP_IMM1_in1_1 }),
  .out1({ S1337 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_621_ (
  .in1({ S1337, S1335 }),
  .out1({ S1275 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_622_ (
  .in1({ S1299, DP_IMM1_in1_2 }),
  .out1({ S1288 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_623_ (
  .in1({ S1288, S1335 }),
  .out1({ S1276 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_624_ (
  .in1({ S1299, DP_IMM1_in1_3 }),
  .out1({ S1289 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_625_ (
  .in1({ S1289, S1335 }),
  .out1({ S1277 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_513_ (
  .in1({ S1307, CU_SE4bits }),
  .out1({ S1287 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__19_ (
  .D({ S1271 }),
  .E({ S1287 }),
  .Q({ DP_IMM1_out_0 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__20_ (
  .D({ S1278 }),
  .E({ S1287 }),
  .Q({ DP_IMM1_out_1 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__21_ (
  .D({ S1279 }),
  .E({ S1287 }),
  .Q({ DP_IMM1_out_2 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__22_ (
  .D({ S1280 }),
  .E({ S1287 }),
  .Q({ DP_IMM1_out_3 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__23_ (
  .D({ S1281 }),
  .E({ S1287 }),
  .Q({ DP_IMM1_out_4 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__24_ (
  .D({ S1282 }),
  .E({ S1287 }),
  .Q({ DP_IMM1_out_5 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__25_ (
  .D({ S1283 }),
  .E({ S1287 }),
  .Q({ DP_IMM1_out_6 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__26_ (
  .D({ S1284 }),
  .E({ S1287 }),
  .Q({ DP_IMM1_out_7 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__27_ (
  .D({ S1285 }),
  .E({ S1287 }),
  .Q({ DP_IMM1_out_8 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__28_ (
  .D({ S1286 }),
  .E({ S1287 }),
  .Q({ DP_IMM1_out_9 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__29_ (
  .D({ S1272 }),
  .E({ S1287 }),
  .Q({ DP_IMM1_out_10 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__30_ (
  .D({ S1273 }),
  .E({ S1287 }),
  .Q({ DP_IMM1_out_11 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__31_ (
  .D({ S1274 }),
  .E({ S1287 }),
  .Q({ DP_IMM1_out_12 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__32_ (
  .D({ S1275 }),
  .E({ S1287 }),
  .Q({ DP_IMM1_out_13 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__33_ (
  .D({ S1276 }),
  .E({ S1287 }),
  .Q({ DP_IMM1_out_14 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__34_ (
  .D({ S1277 }),
  .E({ S1287 }),
  .Q({ DP_IMM1_out_15 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_212_ (
  .in1({ CU_ldIN }),
  .out1({ S1355 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_514_ (
  .in1({ CU_ldIN, S6 }),
  .out1({ S1356 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_626_ (
  .in1({ S1356, DP_IN_out_0 }),
  .out1({ S1357 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_515_ (
  .in1({ S1355, S7 }),
  .out1({ S1358 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_627_ (
  .in1({ S1358, DP_IN_in_0 }),
  .out1({ S1359 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_628_ (
  .in1({ S1359, S1357 }),
  .out1({ S1338 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_629_ (
  .in1({ S1356, DP_IN_out_1 }),
  .out1({ S1360 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_630_ (
  .in1({ S1358, DP_IN_in_1 }),
  .out1({ S1361 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_631_ (
  .in1({ S1361, S1360 }),
  .out1({ S1339 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_632_ (
  .in1({ S1356, DP_IN_out_2 }),
  .out1({ S1362 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_633_ (
  .in1({ S1358, DP_IN_in_2 }),
  .out1({ S1363 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_634_ (
  .in1({ S1363, S1362 }),
  .out1({ S1340 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_635_ (
  .in1({ S1356, DP_IN_out_3 }),
  .out1({ S1364 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_636_ (
  .in1({ S1358, DP_IN_in_3 }),
  .out1({ S1365 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_637_ (
  .in1({ S1365, S1364 }),
  .out1({ S1341 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_638_ (
  .in1({ S1356, DP_IN_out_4 }),
  .out1({ S1366 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_639_ (
  .in1({ S1358, DP_IN_in_4 }),
  .out1({ S1367 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_640_ (
  .in1({ S1367, S1366 }),
  .out1({ S1342 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_641_ (
  .in1({ S1356, DP_IN_out_5 }),
  .out1({ S1368 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_642_ (
  .in1({ S1358, DP_IN_in_5 }),
  .out1({ S1369 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_643_ (
  .in1({ S1369, S1368 }),
  .out1({ S1343 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_644_ (
  .in1({ S1356, DP_IN_out_6 }),
  .out1({ S1370 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_645_ (
  .in1({ S1358, DP_IN_in_6 }),
  .out1({ S1371 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_646_ (
  .in1({ S1371, S1370 }),
  .out1({ S1344 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_647_ (
  .in1({ S1356, DP_IN_out_7 }),
  .out1({ S1372 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_648_ (
  .in1({ S1358, DP_IN_in_7 }),
  .out1({ S1373 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_649_ (
  .in1({ S1373, S1372 }),
  .out1({ S1345 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_650_ (
  .in1({ S1356, DP_IN_out_8 }),
  .out1({ S1374 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_651_ (
  .in1({ S1358, DP_IN_in_8 }),
  .out1({ S1375 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_652_ (
  .in1({ S1375, S1374 }),
  .out1({ S1346 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_653_ (
  .in1({ S1356, DP_IN_out_9 }),
  .out1({ S1376 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_654_ (
  .in1({ S1358, DP_IN_in_9 }),
  .out1({ S1377 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_655_ (
  .in1({ S1377, S1376 }),
  .out1({ S1347 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_656_ (
  .in1({ S1356, DP_IN_out_10 }),
  .out1({ S1378 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_657_ (
  .in1({ S1358, DP_IN_in_10 }),
  .out1({ S1379 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_658_ (
  .in1({ S1379, S1378 }),
  .out1({ S1348 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_659_ (
  .in1({ S1356, DP_IN_out_11 }),
  .out1({ S1380 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_660_ (
  .in1({ S1358, DP_IN_in_11 }),
  .out1({ S1381 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_661_ (
  .in1({ S1381, S1380 }),
  .out1({ S1349 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_662_ (
  .in1({ S1356, DP_IN_out_12 }),
  .out1({ S1382 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_663_ (
  .in1({ S1358, DP_IN_in_12 }),
  .out1({ S1383 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_664_ (
  .in1({ S1383, S1382 }),
  .out1({ S1350 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_665_ (
  .in1({ S1356, DP_IN_out_13 }),
  .out1({ S1384 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_666_ (
  .in1({ S1358, DP_IN_in_13 }),
  .out1({ S1385 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_667_ (
  .in1({ S1385, S1384 }),
  .out1({ S1351 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_668_ (
  .in1({ S1356, DP_IN_out_14 }),
  .out1({ S1386 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_669_ (
  .in1({ S1358, DP_IN_in_14 }),
  .out1({ S1387 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_670_ (
  .in1({ S1387, S1386 }),
  .out1({ S1352 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_671_ (
  .in1({ S1356, DP_IN_out_15 }),
  .out1({ S1388 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_672_ (
  .in1({ S1358, DP_IN_in_15 }),
  .out1({ S1354 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_673_ (
  .in1({ S1354, S1388 }),
  .out1({ S1353 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_19_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1338 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_out_0 }),
  .Si({ S3322 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_20_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1339 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_out_1 }),
  .Si({ S3321 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_21_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1340 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_out_2 }),
  .Si({ S3320 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_22_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1341 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_out_3 }),
  .Si({ S3319 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_23_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1342 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_out_4 }),
  .Si({ S3318 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_24_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1343 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_out_5 }),
  .Si({ S3317 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_25_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1344 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_out_6 }),
  .Si({ S3316 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_26_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1345 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_out_7 }),
  .Si({ S3315 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_27_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1346 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_out_8 }),
  .Si({ S3314 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_28_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1347 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_out_9 }),
  .Si({ S3313 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_29_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1348 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_out_10 }),
  .Si({ S3312 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_30_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1349 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_out_11 }),
  .Si({ S3311 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_31_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1350 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_out_12 }),
  .Si({ S3310 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_32_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1351 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_out_13 }),
  .Si({ S3309 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_33_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1352 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_out_14 }),
  .Si({ S3308 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_34_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1353 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_out_15 }),
  .Si({ S3357 }),
  .global_reset({ 1'b0 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_213_ (
  .in1({ DP_INC_1_in_0 }),
  .out1({ S1406 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_214_ (
  .in1({ DP_INC_1_inc_val_0 }),
  .out1({ S1407 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_215_ (
  .in1({ DP_INC_1_in_1 }),
  .out1({ S1408 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_216_ (
  .in1({ DP_INC_1_inc_val_1 }),
  .out1({ S1409 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_217_ (
  .in1({ DP_INC_1_in_2 }),
  .out1({ S1410 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_218_ (
  .in1({ DP_INC_1_in_3 }),
  .out1({ S1411 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_219_ (
  .in1({ DP_INC_1_in_4 }),
  .out1({ S1412 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_220_ (
  .in1({ DP_INC_1_in_5 }),
  .out1({ S1413 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_221_ (
  .in1({ DP_INC_1_in_6 }),
  .out1({ S1414 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_222_ (
  .in1({ DP_INC_1_in_7 }),
  .out1({ S1415 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_223_ (
  .in1({ DP_INC_1_in_8 }),
  .out1({ S1416 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_224_ (
  .in1({ DP_INC_1_in_9 }),
  .out1({ S1417 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_225_ (
  .in1({ DP_INC_1_in_10 }),
  .out1({ S1418 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_226_ (
  .in1({ DP_INC_1_in_11 }),
  .out1({ S1419 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_227_ (
  .in1({ DP_INC_1_in_12 }),
  .out1({ S1420 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_228_ (
  .in1({ DP_INC_1_in_13 }),
  .out1({ S1421 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_229_ (
  .in1({ DP_INC_1_in_14 }),
  .out1({ S1422 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_230_ (
  .in1({ DP_INC_1_in_15 }),
  .out1({ S1423 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_516_ (
  .in1({ S1407, S1406 }),
  .out1({ S1424 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_674_ (
  .in1({ DP_INC_1_inc_val_0, DP_INC_1_in_0 }),
  .out1({ S1425 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_517_ (
  .in1({ DP_INC_1_inc_val_0, DP_INC_1_in_0 }),
  .out1({ S1426 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_518_ (
  .in1({ S1426, S1424 }),
  .out1({ DP_INC_1_out_0 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_519_ (
  .in1({ S1409, S1408 }),
  .out1({ S1427 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_675_ (
  .in1({ DP_INC_1_inc_val_1, DP_INC_1_in_1 }),
  .out1({ S1428 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_520_ (
  .in1({ DP_INC_1_inc_val_1, DP_INC_1_in_1 }),
  .out1({ S1429 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_231_ (
  .in1({ S1429 }),
  .out1({ S1430 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_521_ (
  .in1({ S1429, S1427 }),
  .out1({ S1431 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_676_ (
  .in1({ S1430, S1428 }),
  .out1({ S1432 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_522_ (
  .in1({ S1432, S1425 }),
  .out1({ S1433 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_677_ (
  .in1({ S1431, S1424 }),
  .out1({ S1434 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_523_ (
  .in1({ S1431, S1424 }),
  .out1({ S1435 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_524_ (
  .in1({ S1435, S1433 }),
  .out1({ DP_INC_1_out_1 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_525_ (
  .in1({ S1433, S1427 }),
  .out1({ S1436 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_678_ (
  .in1({ S1434, S1428 }),
  .out1({ S1437 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_526_ (
  .in1({ S1436, S1410 }),
  .out1({ S1438 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_679_ (
  .in1({ S1437, DP_INC_1_in_2 }),
  .out1({ S1439 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_527_ (
  .in1({ S1437, DP_INC_1_in_2 }),
  .out1({ S1440 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_528_ (
  .in1({ S1440, S1438 }),
  .out1({ DP_INC_1_out_2 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_529_ (
  .in1({ S1439, S1411 }),
  .out1({ S1441 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_680_ (
  .in1({ S1438, DP_INC_1_in_3 }),
  .out1({ S1442 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_530_ (
  .in1({ S1438, DP_INC_1_in_3 }),
  .out1({ S1443 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_531_ (
  .in1({ S1443, S1441 }),
  .out1({ DP_INC_1_out_3 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_532_ (
  .in1({ S1442, S1412 }),
  .out1({ S1444 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_681_ (
  .in1({ S1441, DP_INC_1_in_4 }),
  .out1({ S1445 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_533_ (
  .in1({ S1441, DP_INC_1_in_4 }),
  .out1({ S1446 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_534_ (
  .in1({ S1446, S1444 }),
  .out1({ DP_INC_1_out_4 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_535_ (
  .in1({ S1445, S1413 }),
  .out1({ S1447 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_682_ (
  .in1({ S1444, DP_INC_1_in_5 }),
  .out1({ S1448 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_536_ (
  .in1({ S1444, DP_INC_1_in_5 }),
  .out1({ S1449 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_537_ (
  .in1({ S1449, S1447 }),
  .out1({ DP_INC_1_out_5 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_538_ (
  .in1({ S1448, S1414 }),
  .out1({ S1450 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_683_ (
  .in1({ S1447, DP_INC_1_in_6 }),
  .out1({ S1451 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_539_ (
  .in1({ S1447, DP_INC_1_in_6 }),
  .out1({ S1452 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_540_ (
  .in1({ S1452, S1450 }),
  .out1({ DP_INC_1_out_6 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_541_ (
  .in1({ S1451, S1415 }),
  .out1({ S1453 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_684_ (
  .in1({ S1450, DP_INC_1_in_7 }),
  .out1({ S1454 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_542_ (
  .in1({ S1450, DP_INC_1_in_7 }),
  .out1({ S1455 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_543_ (
  .in1({ S1455, S1453 }),
  .out1({ DP_INC_1_out_7 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_544_ (
  .in1({ S1454, S1416 }),
  .out1({ S1456 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_685_ (
  .in1({ S1453, DP_INC_1_in_8 }),
  .out1({ S1457 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_545_ (
  .in1({ S1453, DP_INC_1_in_8 }),
  .out1({ S1458 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_546_ (
  .in1({ S1458, S1456 }),
  .out1({ DP_INC_1_out_8 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_547_ (
  .in1({ S1457, S1417 }),
  .out1({ S1459 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_686_ (
  .in1({ S1456, DP_INC_1_in_9 }),
  .out1({ S1460 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_548_ (
  .in1({ S1456, DP_INC_1_in_9 }),
  .out1({ S1461 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_549_ (
  .in1({ S1461, S1459 }),
  .out1({ DP_INC_1_out_9 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_550_ (
  .in1({ S1460, S1418 }),
  .out1({ S1389 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_687_ (
  .in1({ S1459, DP_INC_1_in_10 }),
  .out1({ S1390 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_551_ (
  .in1({ S1459, DP_INC_1_in_10 }),
  .out1({ S1391 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_552_ (
  .in1({ S1391, S1389 }),
  .out1({ DP_INC_1_out_10 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_553_ (
  .in1({ S1390, S1419 }),
  .out1({ S1392 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_688_ (
  .in1({ S1389, DP_INC_1_in_11 }),
  .out1({ S1393 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_554_ (
  .in1({ S1389, DP_INC_1_in_11 }),
  .out1({ S1394 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_555_ (
  .in1({ S1394, S1392 }),
  .out1({ DP_INC_1_out_11 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_556_ (
  .in1({ S1393, S1420 }),
  .out1({ S1395 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_689_ (
  .in1({ S1392, DP_INC_1_in_12 }),
  .out1({ S1396 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_557_ (
  .in1({ S1392, DP_INC_1_in_12 }),
  .out1({ S1397 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_558_ (
  .in1({ S1397, S1395 }),
  .out1({ DP_INC_1_out_12 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_559_ (
  .in1({ S1396, S1421 }),
  .out1({ S1398 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_690_ (
  .in1({ S1395, DP_INC_1_in_13 }),
  .out1({ S1399 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_560_ (
  .in1({ S1395, DP_INC_1_in_13 }),
  .out1({ S1400 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_561_ (
  .in1({ S1400, S1398 }),
  .out1({ DP_INC_1_out_13 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_562_ (
  .in1({ S1399, S1422 }),
  .out1({ S1401 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_691_ (
  .in1({ S1398, DP_INC_1_in_14 }),
  .out1({ S1402 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_563_ (
  .in1({ S1398, DP_INC_1_in_14 }),
  .out1({ S1403 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_564_ (
  .in1({ S1403, S1401 }),
  .out1({ DP_INC_1_out_14 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_565_ (
  .in1({ S1401, DP_INC_1_in_15 }),
  .out1({ S1404 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_566_ (
  .in1({ S1402, S1423 }),
  .out1({ S1405 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_567_ (
  .in1({ S1405, S1404 }),
  .out1({ DP_INC_1_out_15 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_232_ (
  .in1({ dataBus[0] }),
  .out1({ S1479 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_233_ (
  .in1({ S0 }),
  .out1({ S1480 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_234_ (
  .in1({ dataBus[1] }),
  .out1({ S1481 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_235_ (
  .in1({ S8 }),
  .out1({ S1482 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_236_ (
  .in1({ dataBus[2] }),
  .out1({ S1483 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_237_ (
  .in1({ dataBus[3] }),
  .out1({ S1484 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_238_ (
  .in1({ dataBus[4] }),
  .out1({ S1485 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_239_ (
  .in1({ dataBus[5] }),
  .out1({ S1486 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_240_ (
  .in1({ dataBus[6] }),
  .out1({ S1487 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_241_ (
  .in1({ dataBus[7] }),
  .out1({ S1488 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_242_ (
  .in1({ dataBus[8] }),
  .out1({ S1489 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_243_ (
  .in1({ dataBus[9] }),
  .out1({ S1490 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_244_ (
  .in1({ dataBus[10] }),
  .out1({ S1491 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_245_ (
  .in1({ dataBus[11] }),
  .out1({ S1492 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_246_ (
  .in1({ dataBus[12] }),
  .out1({ S1493 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_247_ (
  .in1({ dataBus[13] }),
  .out1({ S1494 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_248_ (
  .in1({ dataBus[14] }),
  .out1({ S1495 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_249_ (
  .in1({ dataBus[15] }),
  .out1({ S1496 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_568_ (
  .in1({ S1480, S1479 }),
  .out1({ S1497 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_692_ (
  .in1({ S1, dataBus[0] }),
  .out1({ S1498 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_569_ (
  .in1({ S2, dataBus[0] }),
  .out1({ S1499 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_570_ (
  .in1({ S1499, S1497 }),
  .out1({ DP_INC2_out_0 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_571_ (
  .in1({ S1482, S1481 }),
  .out1({ S1500 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_693_ (
  .in1({ S9, dataBus[1] }),
  .out1({ S1501 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_572_ (
  .in1({ S10, dataBus[1] }),
  .out1({ S1502 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_250_ (
  .in1({ S1502 }),
  .out1({ S1503 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_573_ (
  .in1({ S1502, S1500 }),
  .out1({ S1504 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_694_ (
  .in1({ S1503, S1501 }),
  .out1({ S1505 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_574_ (
  .in1({ S1505, S1498 }),
  .out1({ S1506 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_695_ (
  .in1({ S1504, S1497 }),
  .out1({ S1507 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_575_ (
  .in1({ S1504, S1497 }),
  .out1({ S1508 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_576_ (
  .in1({ S1508, S1506 }),
  .out1({ DP_INC2_out_1 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_577_ (
  .in1({ S1506, S1500 }),
  .out1({ S1509 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_696_ (
  .in1({ S1507, S1501 }),
  .out1({ S1510 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_578_ (
  .in1({ S1509, S1483 }),
  .out1({ S1511 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_697_ (
  .in1({ S1510, dataBus[2] }),
  .out1({ S1512 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_579_ (
  .in1({ S1510, dataBus[2] }),
  .out1({ S1513 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_580_ (
  .in1({ S1513, S1511 }),
  .out1({ DP_INC2_out_2 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_581_ (
  .in1({ S1512, S1484 }),
  .out1({ S1514 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_698_ (
  .in1({ S1511, dataBus[3] }),
  .out1({ S1515 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_582_ (
  .in1({ S1511, dataBus[3] }),
  .out1({ S1516 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_583_ (
  .in1({ S1516, S1514 }),
  .out1({ DP_INC2_out_3 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_584_ (
  .in1({ S1515, S1485 }),
  .out1({ S1517 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_699_ (
  .in1({ S1514, dataBus[4] }),
  .out1({ S1518 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_585_ (
  .in1({ S1514, dataBus[4] }),
  .out1({ S1519 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_586_ (
  .in1({ S1519, S1517 }),
  .out1({ DP_INC2_out_4 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_587_ (
  .in1({ S1518, S1486 }),
  .out1({ S1520 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_700_ (
  .in1({ S1517, dataBus[5] }),
  .out1({ S1521 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_588_ (
  .in1({ S1517, dataBus[5] }),
  .out1({ S1522 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_589_ (
  .in1({ S1522, S1520 }),
  .out1({ DP_INC2_out_5 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_590_ (
  .in1({ S1521, S1487 }),
  .out1({ S1523 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_701_ (
  .in1({ S1520, dataBus[6] }),
  .out1({ S1524 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_591_ (
  .in1({ S1520, dataBus[6] }),
  .out1({ S1525 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_592_ (
  .in1({ S1525, S1523 }),
  .out1({ DP_INC2_out_6 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_593_ (
  .in1({ S1524, S1488 }),
  .out1({ S1526 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_702_ (
  .in1({ S1523, dataBus[7] }),
  .out1({ S1527 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_594_ (
  .in1({ S1523, dataBus[7] }),
  .out1({ S1528 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_595_ (
  .in1({ S1528, S1526 }),
  .out1({ DP_INC2_out_7 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_596_ (
  .in1({ S1527, S1489 }),
  .out1({ S1529 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_703_ (
  .in1({ S1526, dataBus[8] }),
  .out1({ S1530 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_597_ (
  .in1({ S1526, dataBus[8] }),
  .out1({ S1531 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_598_ (
  .in1({ S1531, S1529 }),
  .out1({ DP_INC2_out_8 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_599_ (
  .in1({ S1530, S1490 }),
  .out1({ S1532 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_704_ (
  .in1({ S1529, dataBus[9] }),
  .out1({ S1533 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_600_ (
  .in1({ S1529, dataBus[9] }),
  .out1({ S1534 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_601_ (
  .in1({ S1534, S1532 }),
  .out1({ DP_INC2_out_9 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_602_ (
  .in1({ S1533, S1491 }),
  .out1({ S1462 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_705_ (
  .in1({ S1532, dataBus[10] }),
  .out1({ S1463 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_603_ (
  .in1({ S1532, dataBus[10] }),
  .out1({ S1464 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_604_ (
  .in1({ S1464, S1462 }),
  .out1({ DP_INC2_out_10 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_605_ (
  .in1({ S1463, S1492 }),
  .out1({ S1465 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_706_ (
  .in1({ S1462, dataBus[11] }),
  .out1({ S1466 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_606_ (
  .in1({ S1462, dataBus[11] }),
  .out1({ S1467 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_607_ (
  .in1({ S1467, S1465 }),
  .out1({ DP_INC2_out_11 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_608_ (
  .in1({ S1466, S1493 }),
  .out1({ S1468 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_707_ (
  .in1({ S1465, dataBus[12] }),
  .out1({ S1469 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_609_ (
  .in1({ S1465, dataBus[12] }),
  .out1({ S1470 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_610_ (
  .in1({ S1470, S1468 }),
  .out1({ DP_INC2_out_12 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_611_ (
  .in1({ S1469, S1494 }),
  .out1({ S1471 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_708_ (
  .in1({ S1468, dataBus[13] }),
  .out1({ S1472 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_612_ (
  .in1({ S1468, dataBus[13] }),
  .out1({ S1473 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_613_ (
  .in1({ S1473, S1471 }),
  .out1({ DP_INC2_out_13 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_614_ (
  .in1({ S1472, S1495 }),
  .out1({ S1474 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_709_ (
  .in1({ S1471, dataBus[14] }),
  .out1({ S1475 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_615_ (
  .in1({ S1471, dataBus[14] }),
  .out1({ S1476 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_616_ (
  .in1({ S1476, S1474 }),
  .out1({ DP_INC2_out_14 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_617_ (
  .in1({ S1474, dataBus[15] }),
  .out1({ S1477 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_618_ (
  .in1({ S1475, S1496 }),
  .out1({ S1478 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_619_ (
  .in1({ S1478, S1477 }),
  .out1({ DP_INC2_out_15 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_251_ (
  .in1({ CU_ldIR }),
  .out1({ S1552 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_620_ (
  .in1({ CU_ldIR, S11 }),
  .out1({ S1553 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_710_ (
  .in1({ S1553, CU_inst_0 }),
  .out1({ S1554 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_621_ (
  .in1({ S1552, S12 }),
  .out1({ S1555 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_711_ (
  .in1({ S1555, dataBus[0] }),
  .out1({ S1556 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_712_ (
  .in1({ S1556, S1554 }),
  .out1({ S1535 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_713_ (
  .in1({ S1553, CU_inst_1 }),
  .out1({ S1557 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_714_ (
  .in1({ S1555, dataBus[1] }),
  .out1({ S1558 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_715_ (
  .in1({ S1558, S1557 }),
  .out1({ S1536 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_716_ (
  .in1({ S1553, CU_inst_2 }),
  .out1({ S1559 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_717_ (
  .in1({ S1555, dataBus[2] }),
  .out1({ S1560 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_718_ (
  .in1({ S1560, S1559 }),
  .out1({ S1537 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_719_ (
  .in1({ S1553, CU_inst_3 }),
  .out1({ S1561 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_720_ (
  .in1({ S1555, dataBus[3] }),
  .out1({ S1562 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_721_ (
  .in1({ S1562, S1561 }),
  .out1({ S1538 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_722_ (
  .in1({ S1553, CU_inst_4 }),
  .out1({ S1563 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_723_ (
  .in1({ S1555, dataBus[4] }),
  .out1({ S1564 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_724_ (
  .in1({ S1564, S1563 }),
  .out1({ S1539 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_725_ (
  .in1({ S1553, CU_inst_5 }),
  .out1({ S1565 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_726_ (
  .in1({ S1555, dataBus[5] }),
  .out1({ S1566 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_727_ (
  .in1({ S1566, S1565 }),
  .out1({ S1540 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_728_ (
  .in1({ S1553, CU_inst_6 }),
  .out1({ S1567 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_729_ (
  .in1({ S1555, dataBus[6] }),
  .out1({ S1568 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_730_ (
  .in1({ S1568, S1567 }),
  .out1({ S1541 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_731_ (
  .in1({ S1553, CU_inst_7 }),
  .out1({ S1569 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_732_ (
  .in1({ S1555, dataBus[7] }),
  .out1({ S1570 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_733_ (
  .in1({ S1570, S1569 }),
  .out1({ S1542 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_734_ (
  .in1({ S1553, CU_inst_8 }),
  .out1({ S1571 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_735_ (
  .in1({ S1555, dataBus[8] }),
  .out1({ S1572 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_736_ (
  .in1({ S1572, S1571 }),
  .out1({ S1543 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_737_ (
  .in1({ S1553, CU_inst_9 }),
  .out1({ S1573 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_738_ (
  .in1({ S1555, dataBus[9] }),
  .out1({ S1574 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_739_ (
  .in1({ S1574, S1573 }),
  .out1({ S1544 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_740_ (
  .in1({ S1553, CU_inst_10 }),
  .out1({ S1575 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_741_ (
  .in1({ S1555, dataBus[10] }),
  .out1({ S1576 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_742_ (
  .in1({ S1576, S1575 }),
  .out1({ S1545 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_743_ (
  .in1({ S1553, CU_inst_11 }),
  .out1({ S1577 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_744_ (
  .in1({ S1555, dataBus[11] }),
  .out1({ S1578 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_745_ (
  .in1({ S1578, S1577 }),
  .out1({ S1546 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_746_ (
  .in1({ S1553, CU_inst_12 }),
  .out1({ S1579 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_747_ (
  .in1({ S1555, dataBus[12] }),
  .out1({ S1580 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_748_ (
  .in1({ S1580, S1579 }),
  .out1({ S1547 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_749_ (
  .in1({ S1553, CU_inst_13 }),
  .out1({ S1581 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_750_ (
  .in1({ S1555, dataBus[13] }),
  .out1({ S1582 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_751_ (
  .in1({ S1582, S1581 }),
  .out1({ S1548 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_752_ (
  .in1({ S1553, CU_inst_14 }),
  .out1({ S1583 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_753_ (
  .in1({ S1555, dataBus[14] }),
  .out1({ S1584 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_754_ (
  .in1({ S1584, S1583 }),
  .out1({ S1549 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_755_ (
  .in1({ S1553, CU_inst_15 }),
  .out1({ S1585 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_756_ (
  .in1({ S1555, dataBus[15] }),
  .out1({ S1551 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_757_ (
  .in1({ S1551, S1585 }),
  .out1({ S1550 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_35_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1535 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_0 }),
  .Si({ S3337 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_36_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1536 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_1 }),
  .Si({ S3336 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_37_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1537 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_2 }),
  .Si({ S3335 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_38_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1538 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_3 }),
  .Si({ S3334 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_39_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1539 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_4 }),
  .Si({ S3333 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_40_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1540 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_5 }),
  .Si({ S3332 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_41_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1541 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_6 }),
  .Si({ S3331 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_42_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1542 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_7 }),
  .Si({ S3330 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_43_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1543 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_8 }),
  .Si({ S3329 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_44_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1544 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_9 }),
  .Si({ S3328 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_45_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1545 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_10 }),
  .Si({ S3327 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_46_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1546 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_11 }),
  .Si({ S3326 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_47_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1547 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_12 }),
  .Si({ S3325 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_48_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1548 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_13 }),
  .Si({ S3324 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_49_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1549 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_14 }),
  .Si({ S3323 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_50_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1550 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_15 }),
  .Si({ S3358 }),
  .global_reset({ 1'b0 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_252_ (
  .in1({ DP_AC_out_15 }),
  .out1({ S1652 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_253_ (
  .in1({ DP_LGU1_in1_0 }),
  .out1({ S1653 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_254_ (
  .in1({ DP_LGU1_in1_1 }),
  .out1({ S1654 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_255_ (
  .in1({ DP_AC_out_4 }),
  .out1({ S1655 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_256_ (
  .in1({ DP_AC_out_5 }),
  .out1({ S1656 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_257_ (
  .in1({ DP_LGU1_in1_2 }),
  .out1({ S1657 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_258_ (
  .in1({ DP_LGU1_in1_3 }),
  .out1({ S1658 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_259_ (
  .in1({ DP_LGU1_in1_4 }),
  .out1({ S1659 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_260_ (
  .in1({ CU_SHF_0 }),
  .out1({ S1660 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_261_ (
  .in1({ CU_SHF_1 }),
  .out1({ S1661 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_262_ (
  .in1({ CU_NOT }),
  .out1({ S1662 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_622_ (
  .in1({ DP_LGU1_out_7, DP_LGU1_out_4 }),
  .out1({ S1663 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_623_ (
  .in1({ DP_LGU1_out_2, DP_LGU1_out_1 }),
  .out1({ S1664 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_758_ (
  .in1({ S1664, S1663 }),
  .out1({ S1665 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_624_ (
  .in1({ DP_LGU1_out_14, DP_LGU1_out_13 }),
  .out1({ S1666 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_625_ (
  .in1({ DP_LGU1_out_11, DP_LGU1_out_8 }),
  .out1({ S1667 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_759_ (
  .in1({ S1667, S1666 }),
  .out1({ S1668 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_626_ (
  .in1({ S1668, S1665 }),
  .out1({ S1669 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_627_ (
  .in1({ DP_LGU1_out_6, DP_LGU1_out_5 }),
  .out1({ S1670 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_628_ (
  .in1({ DP_LGU1_out_3, DP_LGU1_out_0 }),
  .out1({ S1671 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_760_ (
  .in1({ S1671, S1670 }),
  .out1({ S1672 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_629_ (
  .in1({ DP_LGU1_N, DP_LGU1_out_12 }),
  .out1({ S1673 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_630_ (
  .in1({ DP_LGU1_out_10, DP_LGU1_out_9 }),
  .out1({ S1674 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_761_ (
  .in1({ S1674, S1673 }),
  .out1({ S1675 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_631_ (
  .in1({ S1675, S1672 }),
  .out1({ S1676 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_762_ (
  .in1({ S1676, S1669 }),
  .out1({ S1677 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_263_ (
  .in1({ S1677 }),
  .out1({ DP_LGU1_Z })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_632_ (
  .in1({ DP_LGU1_in1_15, DP_LGU1_in1_14 }),
  .out1({ S1678 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_264_ (
  .in1({ S1678 }),
  .out1({ S1679 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_633_ (
  .in1({ S1679, DP_LGU1_in1_13 }),
  .out1({ S1680 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_634_ (
  .in1({ DP_LGU1_in1_9, DP_LGU1_in1_10 }),
  .out1({ S1681 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_635_ (
  .in1({ DP_LGU1_in1_11, DP_LGU1_in1_12 }),
  .out1({ S1682 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_763_ (
  .in1({ S1682, S1681 }),
  .out1({ S1683 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_636_ (
  .in1({ DP_LGU1_in1_5, DP_LGU1_in1_6 }),
  .out1({ S1684 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_637_ (
  .in1({ DP_LGU1_in1_7, DP_LGU1_in1_8 }),
  .out1({ S1685 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_764_ (
  .in1({ S1685, S1684 }),
  .out1({ S1686 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_265_ (
  .in1({ S1686 }),
  .out1({ S1687 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_638_ (
  .in1({ S1686, S1683 }),
  .out1({ S1688 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_765_ (
  .in1({ S1687, S1680 }),
  .out1({ S1689 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_639_ (
  .in1({ S1689, S1683 }),
  .out1({ S1690 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_766_ (
  .in1({ S1688, S1680 }),
  .out1({ S1691 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_640_ (
  .in1({ S1691, S1655 }),
  .out1({ S1692 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_767_ (
  .in1({ S1690, DP_AC_out_4 }),
  .out1({ S1693 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_641_ (
  .in1({ S1693, DP_LGU1_in1_0 }),
  .out1({ S1694 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_768_ (
  .in1({ S1692, S1653 }),
  .out1({ S1695 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_642_ (
  .in1({ S1691, S1656 }),
  .out1({ S1696 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_769_ (
  .in1({ S1690, DP_AC_out_5 }),
  .out1({ S1697 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_643_ (
  .in1({ S1697, S1653 }),
  .out1({ S1698 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_770_ (
  .in1({ S1696, DP_LGU1_in1_0 }),
  .out1({ S1699 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_771_ (
  .in1({ S1699, S1695 }),
  .out1({ S1700 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_644_ (
  .in1({ S1700, DP_LGU1_in1_1 }),
  .out1({ S1701 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_266_ (
  .in1({ S1701 }),
  .out1({ S1702 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_772_ (
  .in1({ S1690, DP_AC_out_6 }),
  .out1({ S1703 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_645_ (
  .in1({ S1703, DP_LGU1_in1_0 }),
  .out1({ S1704 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_773_ (
  .in1({ S1690, DP_AC_out_7 }),
  .out1({ S1705 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_774_ (
  .in1({ S1703, S1653 }),
  .out1({ S1706 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_775_ (
  .in1({ S1705, DP_LGU1_in1_0 }),
  .out1({ S1707 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_776_ (
  .in1({ S1707, S1706 }),
  .out1({ S1708 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_267_ (
  .in1({ S1708 }),
  .out1({ S1709 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_777_ (
  .in1({ S1708, DP_LGU1_in1_1 }),
  .out1({ S1710 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_268_ (
  .in1({ S1710 }),
  .out1({ S1711 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_646_ (
  .in1({ S1711, S1701 }),
  .out1({ S1712 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_778_ (
  .in1({ S1710, S1702 }),
  .out1({ S1713 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_779_ (
  .in1({ S1712, DP_LGU1_in1_2 }),
  .out1({ S1714 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_780_ (
  .in1({ S1690, DP_AC_out_2 }),
  .out1({ S1715 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_647_ (
  .in1({ S1715, DP_LGU1_in1_0 }),
  .out1({ S1716 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_781_ (
  .in1({ S1690, DP_AC_out_3 }),
  .out1({ S1717 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_648_ (
  .in1({ S1717, S1653 }),
  .out1({ S1718 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_649_ (
  .in1({ S1718, S1716 }),
  .out1({ S1719 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_269_ (
  .in1({ S1719 }),
  .out1({ S1720 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_650_ (
  .in1({ S1719, S1654 }),
  .out1({ S1721 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_782_ (
  .in1({ S1690, DP_AC_out_1 }),
  .out1({ S1722 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_270_ (
  .in1({ S1722 }),
  .out1({ S1723 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_651_ (
  .in1({ S1722, S1653 }),
  .out1({ S1724 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_783_ (
  .in1({ S1723, DP_LGU1_in1_0 }),
  .out1({ S1725 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_652_ (
  .in1({ S1725, DP_LGU1_in1_1 }),
  .out1({ S1726 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_653_ (
  .in1({ S1726, S1721 }),
  .out1({ S1727 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_654_ (
  .in1({ S1727, DP_LGU1_in1_2 }),
  .out1({ S1728 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_784_ (
  .in1({ S1690, DP_AC_out_0 }),
  .out1({ S1729 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_655_ (
  .in1({ S1729, DP_LGU1_in1_0 }),
  .out1({ S1730 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_785_ (
  .in1({ S1730, S1654 }),
  .out1({ S1731 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_656_ (
  .in1({ S1731, DP_LGU1_in1_2 }),
  .out1({ S1732 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_657_ (
  .in1({ S1732, DP_LGU1_in1_3 }),
  .out1({ S1733 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_271_ (
  .in1({ S1733 }),
  .out1({ S1734 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_658_ (
  .in1({ S1734, S1728 }),
  .out1({ S1735 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_786_ (
  .in1({ S1733, S1714 }),
  .out1({ S1736 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_659_ (
  .in1({ S1736, S1728 }),
  .out1({ S1737 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_787_ (
  .in1({ S1735, S1714 }),
  .out1({ S1738 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_788_ (
  .in1({ S1690, DP_AC_out_8 }),
  .out1({ S1739 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_789_ (
  .in1({ S1739, S1653 }),
  .out1({ S1740 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_790_ (
  .in1({ S1690, DP_AC_out_9 }),
  .out1({ S1741 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_791_ (
  .in1({ S1741, DP_LGU1_in1_0 }),
  .out1({ S1742 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_792_ (
  .in1({ S1742, S1740 }),
  .out1({ S1743 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_793_ (
  .in1({ S1743, S1654 }),
  .out1({ S1744 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_794_ (
  .in1({ S1690, DP_AC_out_10 }),
  .out1({ S1745 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_795_ (
  .in1({ S1745, S1653 }),
  .out1({ S1746 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_796_ (
  .in1({ S1690, DP_AC_out_11 }),
  .out1({ S1747 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_797_ (
  .in1({ S1747, DP_LGU1_in1_0 }),
  .out1({ S1748 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_798_ (
  .in1({ S1748, S1746 }),
  .out1({ S1749 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_272_ (
  .in1({ S1749 }),
  .out1({ S1750 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_799_ (
  .in1({ S1749, DP_LGU1_in1_1 }),
  .out1({ S1751 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_800_ (
  .in1({ S1751, S1744 }),
  .out1({ S1752 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_801_ (
  .in1({ S1752, S1657 }),
  .out1({ S1753 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_802_ (
  .in1({ S1690, DP_AC_out_12 }),
  .out1({ S1754 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_803_ (
  .in1({ S1754, S1653 }),
  .out1({ S1755 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_804_ (
  .in1({ S1690, DP_AC_out_13 }),
  .out1({ S1756 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_805_ (
  .in1({ S1756, DP_LGU1_in1_0 }),
  .out1({ S1757 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_806_ (
  .in1({ S1757, S1755 }),
  .out1({ S1758 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_807_ (
  .in1({ S1758, S1654 }),
  .out1({ S1759 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_808_ (
  .in1({ S1690, DP_AC_out_14 }),
  .out1({ S1760 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_809_ (
  .in1({ S1760, S1653 }),
  .out1({ S1761 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_810_ (
  .in1({ S1690, DP_AC_out_15 }),
  .out1({ S1762 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_811_ (
  .in1({ S1762, DP_LGU1_in1_0 }),
  .out1({ S1763 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_812_ (
  .in1({ S1763, S1761 }),
  .out1({ S1764 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_813_ (
  .in1({ S1764, DP_LGU1_in1_1 }),
  .out1({ S1765 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_814_ (
  .in1({ S1765, S1759 }),
  .out1({ S1766 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_815_ (
  .in1({ S1766, DP_LGU1_in1_2 }),
  .out1({ S1767 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_816_ (
  .in1({ S1767, S1753 }),
  .out1({ S1768 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_817_ (
  .in1({ S1768, DP_LGU1_in1_3 }),
  .out1({ S1769 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_818_ (
  .in1({ S1769, S1738 }),
  .out1({ S1603 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_660_ (
  .in1({ CU_SHF_1, S1660 }),
  .out1({ S1604 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_819_ (
  .in1({ S1732, S1658 }),
  .out1({ S1605 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_820_ (
  .in1({ DP_AC_out_0, CU_AND }),
  .out1({ S1770 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_273_ (
  .in1({ S1770 }),
  .out1({ S1771 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_821_ (
  .in1({ S1771, DP_LGU1_in1_0 }),
  .out1({ S1772 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_661_ (
  .in1({ CU_NOT, CU_AND }),
  .out1({ S1773 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_822_ (
  .in1({ CU_NOT, DP_AC_out_0 }),
  .out1({ S1774 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_274_ (
  .in1({ S1774 }),
  .out1({ S1775 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_662_ (
  .in1({ S1775, CU_AND }),
  .out1({ S1776 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_663_ (
  .in1({ CU_SHF_1, CU_SHF_0 }),
  .out1({ S1777 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_823_ (
  .in1({ S1661, S1660 }),
  .out1({ S1778 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_824_ (
  .in1({ DP_LGU1_in1_0, S1652 }),
  .out1({ S1779 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_825_ (
  .in1({ S1779, S1761 }),
  .out1({ S1780 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_826_ (
  .in1({ S1780, DP_LGU1_in1_1 }),
  .out1({ S1781 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_827_ (
  .in1({ S1781, S1759 }),
  .out1({ S1782 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_828_ (
  .in1({ S1782, DP_LGU1_in1_2 }),
  .out1({ S1783 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_829_ (
  .in1({ S1783, S1753 }),
  .out1({ S1784 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_830_ (
  .in1({ S1784, DP_LGU1_in1_3 }),
  .out1({ S1785 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_664_ (
  .in1({ S1737, DP_LGU1_in1_4 }),
  .out1({ S1786 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_831_ (
  .in1({ S1786, S1785 }),
  .out1({ S1787 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_665_ (
  .in1({ S1659, S1652 }),
  .out1({ S1788 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_832_ (
  .in1({ DP_LGU1_in1_4, DP_AC_out_15 }),
  .out1({ S1789 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_666_ (
  .in1({ S1690, S1652 }),
  .out1({ S1790 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_833_ (
  .in1({ S1691, DP_AC_out_15 }),
  .out1({ S1791 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_667_ (
  .in1({ S1790, S1788 }),
  .out1({ S1792 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_834_ (
  .in1({ S1792, S1787 }),
  .out1({ S1793 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_835_ (
  .in1({ S1793, S1777 }),
  .out1({ S1794 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_836_ (
  .in1({ S1778, S1659 }),
  .out1({ S1795 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_668_ (
  .in1({ S1795, S1636 }),
  .out1({ S1796 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_669_ (
  .in1({ S1796, CU_NOT }),
  .out1({ S1797 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_837_ (
  .in1({ S1797, S1794 }),
  .out1({ S1798 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_838_ (
  .in1({ S1798, S1776 }),
  .out1({ S1799 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_839_ (
  .in1({ S1799, S1772 }),
  .out1({ S1586 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_840_ (
  .in1({ S1722, S1653 }),
  .out1({ S1800 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_841_ (
  .in1({ S1715, DP_LGU1_in1_0 }),
  .out1({ S1801 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_842_ (
  .in1({ S1801, S1800 }),
  .out1({ S1802 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_843_ (
  .in1({ S1802, S1654 }),
  .out1({ S1803 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_844_ (
  .in1({ S1717, S1653 }),
  .out1({ S1804 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_845_ (
  .in1({ S1693, DP_LGU1_in1_0 }),
  .out1({ S1805 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_846_ (
  .in1({ S1805, S1804 }),
  .out1({ S1806 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_847_ (
  .in1({ S1806, DP_LGU1_in1_1 }),
  .out1({ S1807 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_848_ (
  .in1({ S1807, S1803 }),
  .out1({ S1808 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_849_ (
  .in1({ S1808, S1657 }),
  .out1({ S1809 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_850_ (
  .in1({ S1697, S1653 }),
  .out1({ S1810 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_851_ (
  .in1({ S1703, DP_LGU1_in1_0 }),
  .out1({ S1811 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_852_ (
  .in1({ S1811, S1810 }),
  .out1({ S1812 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_853_ (
  .in1({ S1812, S1654 }),
  .out1({ S1813 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_854_ (
  .in1({ S1705, S1653 }),
  .out1({ S1814 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_855_ (
  .in1({ S1739, DP_LGU1_in1_0 }),
  .out1({ S1815 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_856_ (
  .in1({ S1815, S1814 }),
  .out1({ S1816 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_857_ (
  .in1({ S1816, DP_LGU1_in1_1 }),
  .out1({ S1817 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_858_ (
  .in1({ S1817, S1813 }),
  .out1({ S1818 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_859_ (
  .in1({ S1818, DP_LGU1_in1_2 }),
  .out1({ S1819 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_860_ (
  .in1({ S1819, S1809 }),
  .out1({ S1820 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_861_ (
  .in1({ S1820, S1658 }),
  .out1({ S1821 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_670_ (
  .in1({ S1745, S1653 }),
  .out1({ S1822 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_862_ (
  .in1({ S1741, S1653 }),
  .out1({ S1823 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_863_ (
  .in1({ S1745, DP_LGU1_in1_0 }),
  .out1({ S1824 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_864_ (
  .in1({ S1824, S1823 }),
  .out1({ S1825 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_275_ (
  .in1({ S1825 }),
  .out1({ S1826 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_671_ (
  .in1({ S1826, DP_LGU1_in1_1 }),
  .out1({ S1827 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_865_ (
  .in1({ S1825, S1654 }),
  .out1({ S1828 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_672_ (
  .in1({ S1754, S1653 }),
  .out1({ S1829 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_673_ (
  .in1({ S1747, DP_LGU1_in1_0 }),
  .out1({ S1830 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_674_ (
  .in1({ S1830, S1829 }),
  .out1({ S1831 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_866_ (
  .in1({ S1831, DP_LGU1_in1_1 }),
  .out1({ S1832 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_276_ (
  .in1({ S1832 }),
  .out1({ S1833 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_675_ (
  .in1({ S1833, S1827 }),
  .out1({ S1834 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_867_ (
  .in1({ S1832, S1828 }),
  .out1({ S1835 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_676_ (
  .in1({ S1834, DP_LGU1_in1_2 }),
  .out1({ S1836 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_868_ (
  .in1({ S1835, S1657 }),
  .out1({ S1837 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_677_ (
  .in1({ S1760, S1653 }),
  .out1({ S1838 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_678_ (
  .in1({ S1756, DP_LGU1_in1_0 }),
  .out1({ S1839 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_679_ (
  .in1({ S1839, S1838 }),
  .out1({ S1840 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_680_ (
  .in1({ S1840, DP_LGU1_in1_1 }),
  .out1({ S1841 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_681_ (
  .in1({ S1762, DP_LGU1_in1_0 }),
  .out1({ S1842 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_869_ (
  .in1({ S1842, DP_LGU1_in1_1 }),
  .out1({ S1843 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_277_ (
  .in1({ S1843 }),
  .out1({ S1844 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_682_ (
  .in1({ S1844, S1841 }),
  .out1({ S1845 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_870_ (
  .in1({ S1845, DP_LGU1_in1_2 }),
  .out1({ S1846 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_871_ (
  .in1({ S1846, S1837 }),
  .out1({ S1847 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_872_ (
  .in1({ S1847, DP_LGU1_in1_3 }),
  .out1({ S1848 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_873_ (
  .in1({ S1848, S1821 }),
  .out1({ S1606 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_874_ (
  .in1({ S1729, DP_LGU1_in1_0 }),
  .out1({ S1849 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_875_ (
  .in1({ S1849, S1800 }),
  .out1({ S1850 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_278_ (
  .in1({ S1850 }),
  .out1({ S1851 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_876_ (
  .in1({ S1851, S1654 }),
  .out1({ S1852 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_683_ (
  .in1({ S1852, DP_LGU1_in1_2 }),
  .out1({ S1853 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_279_ (
  .in1({ S1853 }),
  .out1({ S1854 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_877_ (
  .in1({ S1853, S1658 }),
  .out1({ S1607 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_878_ (
  .in1({ DP_AC_out_1, CU_AND }),
  .out1({ S1855 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_280_ (
  .in1({ S1855 }),
  .out1({ S1856 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_879_ (
  .in1({ S1856, DP_LGU1_in1_1 }),
  .out1({ S1857 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_684_ (
  .in1({ S1637, DP_LGU1_in1_4 }),
  .out1({ S1858 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_685_ (
  .in1({ S1858, S1777 }),
  .out1({ S1859 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_281_ (
  .in1({ S1859 }),
  .out1({ S1860 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_686_ (
  .in1({ S1788, S1778 }),
  .out1({ S1861 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_880_ (
  .in1({ S1789, S1777 }),
  .out1({ S1862 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_687_ (
  .in1({ S1821, S1790 }),
  .out1({ S1863 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_688_ (
  .in1({ S1837, S1790 }),
  .out1({ S1864 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_881_ (
  .in1({ S1836, S1791 }),
  .out1({ S1865 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_689_ (
  .in1({ S1691, DP_LGU1_in1_1 }),
  .out1({ S1866 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_690_ (
  .in1({ S1866, S1652 }),
  .out1({ S1867 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_691_ (
  .in1({ S1867, S1841 }),
  .out1({ S1868 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_882_ (
  .in1({ S1868, DP_LGU1_in1_2 }),
  .out1({ S1869 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_282_ (
  .in1({ S1869 }),
  .out1({ S1870 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_692_ (
  .in1({ S1870, S1864 }),
  .out1({ S1871 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_883_ (
  .in1({ S1869, S1865 }),
  .out1({ S1872 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_693_ (
  .in1({ S1871, S1658 }),
  .out1({ S1873 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_694_ (
  .in1({ S1873, S1863 }),
  .out1({ S1874 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_884_ (
  .in1({ S1874, S1659 }),
  .out1({ S1875 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_885_ (
  .in1({ S1875, S1861 }),
  .out1({ S1876 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_886_ (
  .in1({ S1876, S1860 }),
  .out1({ S1877 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_887_ (
  .in1({ S1877, S1662 }),
  .out1({ S1878 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_888_ (
  .in1({ CU_NOT, DP_AC_out_1 }),
  .out1({ S1879 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_283_ (
  .in1({ S1879 }),
  .out1({ S1880 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_695_ (
  .in1({ S1880, CU_AND }),
  .out1({ S1881 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_889_ (
  .in1({ S1881, S1878 }),
  .out1({ S1882 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_890_ (
  .in1({ S1882, S1857 }),
  .out1({ S1593 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_696_ (
  .in1({ S1700, S1654 }),
  .out1({ S1883 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_697_ (
  .in1({ S1720, DP_LGU1_in1_1 }),
  .out1({ S1884 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_698_ (
  .in1({ S1884, S1883 }),
  .out1({ S1885 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_699_ (
  .in1({ S1885, DP_LGU1_in1_2 }),
  .out1({ S1886 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_700_ (
  .in1({ S1709, DP_LGU1_in1_1 }),
  .out1({ S1887 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_891_ (
  .in1({ S1708, S1654 }),
  .out1({ S1888 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_892_ (
  .in1({ S1743, DP_LGU1_in1_1 }),
  .out1({ S1889 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_284_ (
  .in1({ S1889 }),
  .out1({ S1890 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_701_ (
  .in1({ S1890, S1887 }),
  .out1({ S1891 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_893_ (
  .in1({ S1889, S1888 }),
  .out1({ S1892 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_702_ (
  .in1({ S1891, S1657 }),
  .out1({ S1893 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_703_ (
  .in1({ S1893, S1886 }),
  .out1({ S1894 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_894_ (
  .in1({ S1891, DP_LGU1_in1_2 }),
  .out1({ S1895 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_704_ (
  .in1({ S1884, DP_LGU1_in1_2 }),
  .out1({ S1896 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_285_ (
  .in1({ S1896 }),
  .out1({ S1897 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_705_ (
  .in1({ S1897, S1883 }),
  .out1({ S1898 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_706_ (
  .in1({ S1898, DP_LGU1_in1_3 }),
  .out1({ S1899 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_707_ (
  .in1({ S1894, DP_LGU1_in1_3 }),
  .out1({ S1900 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_895_ (
  .in1({ S1899, S1895 }),
  .out1({ S1901 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_708_ (
  .in1({ S1750, DP_LGU1_in1_1 }),
  .out1({ S1902 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_896_ (
  .in1({ S1749, S1654 }),
  .out1({ S1903 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_897_ (
  .in1({ S1758, DP_LGU1_in1_1 }),
  .out1({ S1904 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_286_ (
  .in1({ S1904 }),
  .out1({ S1905 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_709_ (
  .in1({ S1905, S1902 }),
  .out1({ S1906 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_898_ (
  .in1({ S1904, S1903 }),
  .out1({ S1907 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_710_ (
  .in1({ S1906, DP_LGU1_in1_2 }),
  .out1({ S1908 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_899_ (
  .in1({ S1907, S1657 }),
  .out1({ S1909 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_711_ (
  .in1({ S1764, DP_LGU1_in1_1 }),
  .out1({ S1910 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_287_ (
  .in1({ S1910 }),
  .out1({ S1911 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_712_ (
  .in1({ S1910, S1657 }),
  .out1({ S1912 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_713_ (
  .in1({ S1912, S1908 }),
  .out1({ S1913 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_288_ (
  .in1({ S1913 }),
  .out1({ S1914 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_900_ (
  .in1({ S1914, DP_LGU1_in1_3 }),
  .out1({ S1915 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_901_ (
  .in1({ S1915, S1901 }),
  .out1({ S1608 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_714_ (
  .in1({ S1724, S1716 }),
  .out1({ S1916 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_715_ (
  .in1({ S1916, DP_LGU1_in1_1 }),
  .out1({ S1917 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_902_ (
  .in1({ S1730, DP_LGU1_in1_1 }),
  .out1({ S1918 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_289_ (
  .in1({ S1918 }),
  .out1({ S1919 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_716_ (
  .in1({ S1919, S1917 }),
  .out1({ S1920 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_717_ (
  .in1({ S1920, DP_LGU1_in1_2 }),
  .out1({ S1921 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_290_ (
  .in1({ S1921 }),
  .out1({ S1922 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_903_ (
  .in1({ S1921, S1658 }),
  .out1({ S1609 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_904_ (
  .in1({ DP_AC_out_2, CU_AND }),
  .out1({ S1923 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_291_ (
  .in1({ S1923 }),
  .out1({ S1924 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_905_ (
  .in1({ S1924, DP_LGU1_in1_2 }),
  .out1({ S1925 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_718_ (
  .in1({ S1638, DP_LGU1_in1_4 }),
  .out1({ S1926 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_719_ (
  .in1({ S1926, S1777 }),
  .out1({ S1927 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_292_ (
  .in1({ S1927 }),
  .out1({ S1928 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_906_ (
  .in1({ S1900, S1791 }),
  .out1({ S1929 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_720_ (
  .in1({ S1909, S1790 }),
  .out1({ S1930 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_907_ (
  .in1({ S1908, S1791 }),
  .out1({ S1931 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_721_ (
  .in1({ S1780, DP_LGU1_in1_1 }),
  .out1({ S1932 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_722_ (
  .in1({ S1932, S1867 }),
  .out1({ S1933 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_908_ (
  .in1({ S1933, DP_LGU1_in1_2 }),
  .out1({ S1934 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_293_ (
  .in1({ S1934 }),
  .out1({ S1935 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_723_ (
  .in1({ S1935, S1930 }),
  .out1({ S1936 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_909_ (
  .in1({ S1934, S1931 }),
  .out1({ S1937 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_724_ (
  .in1({ S1936, S1658 }),
  .out1({ S1938 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_725_ (
  .in1({ S1938, DP_LGU1_in1_4 }),
  .out1({ S1939 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_910_ (
  .in1({ S1939, S1929 }),
  .out1({ S1940 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_911_ (
  .in1({ S1940, S1861 }),
  .out1({ S1941 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_912_ (
  .in1({ S1941, S1928 }),
  .out1({ S1942 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_913_ (
  .in1({ S1942, S1662 }),
  .out1({ S1943 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_914_ (
  .in1({ CU_NOT, DP_AC_out_2 }),
  .out1({ S1944 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_294_ (
  .in1({ S1944 }),
  .out1({ S1945 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_726_ (
  .in1({ S1945, CU_AND }),
  .out1({ S1946 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_915_ (
  .in1({ S1946, S1943 }),
  .out1({ S1947 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_916_ (
  .in1({ S1947, S1925 }),
  .out1({ S1594 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_917_ (
  .in1({ S1806, S1654 }),
  .out1({ S1948 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_918_ (
  .in1({ S1812, DP_LGU1_in1_1 }),
  .out1({ S1949 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_919_ (
  .in1({ S1949, S1948 }),
  .out1({ S1950 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_920_ (
  .in1({ S1950, S1657 }),
  .out1({ S1951 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_921_ (
  .in1({ S1816, S1654 }),
  .out1({ S1952 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_922_ (
  .in1({ S1825, DP_LGU1_in1_1 }),
  .out1({ S1953 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_923_ (
  .in1({ S1953, S1952 }),
  .out1({ S1954 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_924_ (
  .in1({ S1954, DP_LGU1_in1_2 }),
  .out1({ S1955 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_925_ (
  .in1({ S1955, S1951 }),
  .out1({ S1956 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_926_ (
  .in1({ S1956, S1658 }),
  .out1({ S1957 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_927_ (
  .in1({ S1842, S1654 }),
  .out1({ S1958 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_727_ (
  .in1({ S1958, S1657 }),
  .out1({ S1959 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_928_ (
  .in1({ S1831, S1654 }),
  .out1({ S1960 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_929_ (
  .in1({ S1840, DP_LGU1_in1_1 }),
  .out1({ S1961 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_930_ (
  .in1({ S1961, S1960 }),
  .out1({ S1962 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_728_ (
  .in1({ S1962, DP_LGU1_in1_2 }),
  .out1({ S1963 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_729_ (
  .in1({ S1963, S1959 }),
  .out1({ S1964 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_931_ (
  .in1({ S1964, DP_LGU1_in1_3 }),
  .out1({ S1965 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_932_ (
  .in1({ S1965, S1957 }),
  .out1({ S1610 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_933_ (
  .in1({ S1804, S1801 }),
  .out1({ S1966 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_934_ (
  .in1({ S1966, S1654 }),
  .out1({ S1967 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_935_ (
  .in1({ S1850, DP_LGU1_in1_1 }),
  .out1({ S1968 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_936_ (
  .in1({ S1968, S1967 }),
  .out1({ S1969 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_730_ (
  .in1({ S1969, DP_LGU1_in1_2 }),
  .out1({ S1970 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_295_ (
  .in1({ S1970 }),
  .out1({ S1971 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_937_ (
  .in1({ S1970, S1658 }),
  .out1({ S1611 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_938_ (
  .in1({ DP_AC_out_3, CU_AND }),
  .out1({ S1972 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_296_ (
  .in1({ S1972 }),
  .out1({ S1973 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_939_ (
  .in1({ S1973, DP_LGU1_in1_3 }),
  .out1({ S1974 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_731_ (
  .in1({ S1639, DP_LGU1_in1_4 }),
  .out1({ S1975 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_732_ (
  .in1({ S1975, S1777 }),
  .out1({ S1976 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_733_ (
  .in1({ S1957, S1790 }),
  .out1({ S1977 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_940_ (
  .in1({ DP_LGU1_in1_2, DP_AC_out_15 }),
  .out1({ S1978 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_297_ (
  .in1({ S1978 }),
  .out1({ S1979 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_941_ (
  .in1({ S1978, S1791 }),
  .out1({ S1980 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_734_ (
  .in1({ S1980, S1963 }),
  .out1({ S1981 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_942_ (
  .in1({ S1981, DP_LGU1_in1_3 }),
  .out1({ S1982 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_943_ (
  .in1({ S1982, S1659 }),
  .out1({ S1983 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_735_ (
  .in1({ S1983, S1977 }),
  .out1({ S1984 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_736_ (
  .in1({ S1984, S1862 }),
  .out1({ S1985 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_737_ (
  .in1({ S1985, S1976 }),
  .out1({ S1986 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_738_ (
  .in1({ S1986, CU_NOT }),
  .out1({ S1987 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_298_ (
  .in1({ S1987 }),
  .out1({ S1988 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_944_ (
  .in1({ CU_NOT, DP_AC_out_3 }),
  .out1({ S1989 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_299_ (
  .in1({ S1989 }),
  .out1({ S1990 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_739_ (
  .in1({ S1990, CU_AND }),
  .out1({ S1991 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_945_ (
  .in1({ S1991, S1988 }),
  .out1({ S1992 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_946_ (
  .in1({ S1992, S1974 }),
  .out1({ S1595 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_947_ (
  .in1({ S1713, S1657 }),
  .out1({ S1993 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_948_ (
  .in1({ S1752, DP_LGU1_in1_2 }),
  .out1({ S1994 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_949_ (
  .in1({ S1994, S1993 }),
  .out1({ S1995 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_950_ (
  .in1({ S1995, S1658 }),
  .out1({ S1996 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_740_ (
  .in1({ S1766, DP_LGU1_in1_2 }),
  .out1({ S1997 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_300_ (
  .in1({ S1997 }),
  .out1({ S1998 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_951_ (
  .in1({ S1998, DP_LGU1_in1_3 }),
  .out1({ S1999 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_952_ (
  .in1({ S1999, S1996 }),
  .out1({ S1612 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_741_ (
  .in1({ S1718, S1694 }),
  .out1({ S2000 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_953_ (
  .in1({ S2000, S1654 }),
  .out1({ S2001 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_954_ (
  .in1({ S1916, DP_LGU1_in1_1 }),
  .out1({ S2002 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_955_ (
  .in1({ S2002, S2001 }),
  .out1({ S2003 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_956_ (
  .in1({ S2003, S1657 }),
  .out1({ S2004 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_957_ (
  .in1({ S1731, DP_LGU1_in1_2 }),
  .out1({ S2005 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_958_ (
  .in1({ S2005, S2004 }),
  .out1({ S2006 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_742_ (
  .in1({ S2006, DP_LGU1_in1_3 }),
  .out1({ S2007 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_301_ (
  .in1({ S2007 }),
  .out1({ S1613 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_743_ (
  .in1({ S1659, S1655 }),
  .out1({ S2008 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_959_ (
  .in1({ S2008, CU_AND }),
  .out1({ S2009 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_744_ (
  .in1({ S1640, DP_LGU1_in1_4 }),
  .out1({ S2010 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_745_ (
  .in1({ S2010, S1777 }),
  .out1({ S2011 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_746_ (
  .in1({ S1996, S1790 }),
  .out1({ S2012 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_747_ (
  .in1({ S1782, DP_LGU1_in1_2 }),
  .out1({ S2013 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_748_ (
  .in1({ S2013, S1980 }),
  .out1({ S2014 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_960_ (
  .in1({ S2014, DP_LGU1_in1_3 }),
  .out1({ S2015 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_961_ (
  .in1({ S2015, S1659 }),
  .out1({ S2016 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_749_ (
  .in1({ S2016, S2012 }),
  .out1({ S2017 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_750_ (
  .in1({ S2017, S1862 }),
  .out1({ S2018 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_751_ (
  .in1({ S2018, S2011 }),
  .out1({ S2019 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_752_ (
  .in1({ S2019, CU_NOT }),
  .out1({ S2020 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_302_ (
  .in1({ S2020 }),
  .out1({ S2021 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_962_ (
  .in1({ CU_NOT, DP_AC_out_4 }),
  .out1({ S2022 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_303_ (
  .in1({ S2022 }),
  .out1({ S2023 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_753_ (
  .in1({ S2023, CU_AND }),
  .out1({ S2024 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_963_ (
  .in1({ S2024, S2021 }),
  .out1({ S2025 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_964_ (
  .in1({ S2025, S2009 }),
  .out1({ S1596 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_754_ (
  .in1({ S1818, DP_LGU1_in1_2 }),
  .out1({ S2026 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_755_ (
  .in1({ S2026, DP_LGU1_in1_3 }),
  .out1({ S2027 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_965_ (
  .in1({ S1834, DP_LGU1_in1_2 }),
  .out1({ S2028 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_966_ (
  .in1({ S2028, S2027 }),
  .out1({ S2029 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_756_ (
  .in1({ S1845, DP_LGU1_in1_2 }),
  .out1({ S2030 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_304_ (
  .in1({ S2030 }),
  .out1({ S2031 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_967_ (
  .in1({ S2031, DP_LGU1_in1_3 }),
  .out1({ S2032 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_968_ (
  .in1({ S2032, S2029 }),
  .out1({ S1614 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_969_ (
  .in1({ S1810, S1805 }),
  .out1({ S2033 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_970_ (
  .in1({ S2033, S1654 }),
  .out1({ S2034 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_971_ (
  .in1({ S1966, DP_LGU1_in1_1 }),
  .out1({ S2035 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_972_ (
  .in1({ S2035, S2034 }),
  .out1({ S2036 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_973_ (
  .in1({ S2036, S1657 }),
  .out1({ S2037 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_974_ (
  .in1({ S1852, DP_LGU1_in1_2 }),
  .out1({ S2038 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_975_ (
  .in1({ S2038, S2037 }),
  .out1({ S2039 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_757_ (
  .in1({ S2039, DP_LGU1_in1_3 }),
  .out1({ S2040 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_305_ (
  .in1({ S2040 }),
  .out1({ S1615 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_976_ (
  .in1({ DP_LGU1_in1_5, CU_AND }),
  .out1({ S2041 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_306_ (
  .in1({ S2041 }),
  .out1({ S2042 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_977_ (
  .in1({ S2042, DP_AC_out_5 }),
  .out1({ S2043 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_758_ (
  .in1({ S1641, DP_LGU1_in1_4 }),
  .out1({ S2044 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_759_ (
  .in1({ S2044, S1777 }),
  .out1({ S2045 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_307_ (
  .in1({ S2045 }),
  .out1({ S2046 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_760_ (
  .in1({ S2029, S1790 }),
  .out1({ S2047 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_761_ (
  .in1({ S1868, DP_LGU1_in1_2 }),
  .out1({ S2048 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_308_ (
  .in1({ S2048 }),
  .out1({ S2049 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_762_ (
  .in1({ S2048, S1979 }),
  .out1({ S2050 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_978_ (
  .in1({ S2049, S1978 }),
  .out1({ S2051 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_763_ (
  .in1({ S2051, S1658 }),
  .out1({ S2052 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_764_ (
  .in1({ S2052, S2047 }),
  .out1({ S2053 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_979_ (
  .in1({ S2053, S1659 }),
  .out1({ S2054 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_980_ (
  .in1({ S2054, S1861 }),
  .out1({ S2055 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_981_ (
  .in1({ S2055, S2046 }),
  .out1({ S2056 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_982_ (
  .in1({ S2056, S1662 }),
  .out1({ S2057 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_983_ (
  .in1({ CU_NOT, DP_AC_out_5 }),
  .out1({ S2058 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_309_ (
  .in1({ S2058 }),
  .out1({ S2059 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_765_ (
  .in1({ S2059, CU_AND }),
  .out1({ S2060 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_984_ (
  .in1({ S2060, S2057 }),
  .out1({ S2061 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_985_ (
  .in1({ S2061, S2043 }),
  .out1({ S1597 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_766_ (
  .in1({ S1892, DP_LGU1_in1_2 }),
  .out1({ S2062 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_767_ (
  .in1({ S2062, DP_LGU1_in1_3 }),
  .out1({ S2063 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_986_ (
  .in1({ S1906, DP_LGU1_in1_2 }),
  .out1({ S2064 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_987_ (
  .in1({ S2064, S2063 }),
  .out1({ S2065 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_768_ (
  .in1({ S1911, DP_LGU1_in1_2 }),
  .out1({ S2066 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_988_ (
  .in1({ S1910, S1657 }),
  .out1({ S2067 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_989_ (
  .in1({ S2067, DP_LGU1_in1_3 }),
  .out1({ S2068 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_990_ (
  .in1({ S2068, S2065 }),
  .out1({ S1616 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_769_ (
  .in1({ S1704, S1698 }),
  .out1({ S2069 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_991_ (
  .in1({ S2069, S1654 }),
  .out1({ S2070 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_992_ (
  .in1({ S2000, DP_LGU1_in1_1 }),
  .out1({ S2071 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_993_ (
  .in1({ S2071, S2070 }),
  .out1({ S2072 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_994_ (
  .in1({ S2072, S1657 }),
  .out1({ S2073 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_995_ (
  .in1({ S1920, DP_LGU1_in1_2 }),
  .out1({ S2074 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_996_ (
  .in1({ S2074, S2073 }),
  .out1({ S2075 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_770_ (
  .in1({ S2075, DP_LGU1_in1_3 }),
  .out1({ S2076 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_310_ (
  .in1({ S2076 }),
  .out1({ S1617 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_997_ (
  .in1({ DP_LGU1_in1_6, CU_AND }),
  .out1({ S2077 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_311_ (
  .in1({ S2077 }),
  .out1({ S2078 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_998_ (
  .in1({ S2078, DP_AC_out_6 }),
  .out1({ S2079 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_771_ (
  .in1({ S1642, DP_LGU1_in1_4 }),
  .out1({ S2080 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_772_ (
  .in1({ S2080, S1777 }),
  .out1({ S2081 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_312_ (
  .in1({ S2081 }),
  .out1({ S2082 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_773_ (
  .in1({ S2065, S1790 }),
  .out1({ S2083 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_774_ (
  .in1({ S1933, DP_LGU1_in1_2 }),
  .out1({ S2084 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_313_ (
  .in1({ S2084 }),
  .out1({ S2085 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_775_ (
  .in1({ S2084, S1979 }),
  .out1({ S2086 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_999_ (
  .in1({ S2085, S1978 }),
  .out1({ S2087 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_776_ (
  .in1({ S2087, S1658 }),
  .out1({ S2088 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_777_ (
  .in1({ S2088, S2083 }),
  .out1({ S2089 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1000_ (
  .in1({ S2089, S1659 }),
  .out1({ S2090 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1001_ (
  .in1({ S2090, S1861 }),
  .out1({ S2091 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1002_ (
  .in1({ S2091, S2082 }),
  .out1({ S2092 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1003_ (
  .in1({ S2092, S1662 }),
  .out1({ S2093 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1004_ (
  .in1({ CU_NOT, DP_AC_out_6 }),
  .out1({ S2094 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_314_ (
  .in1({ S2094 }),
  .out1({ S2095 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_778_ (
  .in1({ S2095, CU_AND }),
  .out1({ S2096 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1005_ (
  .in1({ S2096, S2093 }),
  .out1({ S2097 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1006_ (
  .in1({ S2097, S2079 }),
  .out1({ S1598 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_779_ (
  .in1({ S1962, S1657 }),
  .out1({ S2098 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_780_ (
  .in1({ S1954, DP_LGU1_in1_2 }),
  .out1({ S2099 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_781_ (
  .in1({ S2099, S2098 }),
  .out1({ S2100 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_782_ (
  .in1({ S2100, DP_LGU1_in1_3 }),
  .out1({ S2101 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_315_ (
  .in1({ S2101 }),
  .out1({ S2102 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_783_ (
  .in1({ S1958, DP_LGU1_in1_2 }),
  .out1({ S2103 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1007_ (
  .in1({ S2103, DP_LGU1_in1_3 }),
  .out1({ S2104 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_316_ (
  .in1({ S2104 }),
  .out1({ S2105 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_784_ (
  .in1({ S2105, S2101 }),
  .out1({ S1618 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1008_ (
  .in1({ S1814, S1811 }),
  .out1({ S2106 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1009_ (
  .in1({ S2106, S1654 }),
  .out1({ S2107 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1010_ (
  .in1({ S2033, DP_LGU1_in1_1 }),
  .out1({ S2108 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1011_ (
  .in1({ S2108, S2107 }),
  .out1({ S2109 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1012_ (
  .in1({ S2109, S1657 }),
  .out1({ S2110 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1013_ (
  .in1({ S1969, DP_LGU1_in1_2 }),
  .out1({ S2111 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1014_ (
  .in1({ S2111, S2110 }),
  .out1({ S2112 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_785_ (
  .in1({ S2112, DP_LGU1_in1_3 }),
  .out1({ S2113 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_317_ (
  .in1({ S2113 }),
  .out1({ S1619 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_786_ (
  .in1({ S1643, DP_LGU1_in1_4 }),
  .out1({ S2114 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_787_ (
  .in1({ S2114, S1777 }),
  .out1({ S2115 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_788_ (
  .in1({ DP_LGU1_in1_4, DP_LGU1_in1_3 }),
  .out1({ S2116 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_318_ (
  .in1({ S2116 }),
  .out1({ S2117 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_789_ (
  .in1({ S2116, S1652 }),
  .out1({ S2118 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_790_ (
  .in1({ S2118, S1778 }),
  .out1({ S2119 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1015_ (
  .in1({ S2119, S1791 }),
  .out1({ S2120 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_791_ (
  .in1({ S2102, DP_LGU1_in1_4 }),
  .out1({ S2121 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_792_ (
  .in1({ S2121, S2120 }),
  .out1({ S2122 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_793_ (
  .in1({ S2122, S2115 }),
  .out1({ S2123 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_794_ (
  .in1({ S2123, CU_NOT }),
  .out1({ S2124 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_319_ (
  .in1({ S2124 }),
  .out1({ S2125 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1016_ (
  .in1({ CU_NOT, DP_AC_out_7 }),
  .out1({ S2126 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_320_ (
  .in1({ S2126 }),
  .out1({ S2127 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_795_ (
  .in1({ S2127, CU_AND }),
  .out1({ S2128 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1017_ (
  .in1({ S2128, S2125 }),
  .out1({ S2129 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1018_ (
  .in1({ DP_LGU1_in1_7, CU_AND }),
  .out1({ S2130 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_321_ (
  .in1({ S2130 }),
  .out1({ S2131 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1019_ (
  .in1({ S2131, DP_AC_out_7 }),
  .out1({ S2132 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1020_ (
  .in1({ S2132, S2129 }),
  .out1({ S1599 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_796_ (
  .in1({ S1768, DP_LGU1_in1_3 }),
  .out1({ S2133 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_322_ (
  .in1({ S2133 }),
  .out1({ S1620 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_797_ (
  .in1({ S2003, S1657 }),
  .out1({ S2134 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1021_ (
  .in1({ S1740, S1707 }),
  .out1({ S2135 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1022_ (
  .in1({ S2135, S1654 }),
  .out1({ S2136 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1023_ (
  .in1({ S2069, DP_LGU1_in1_1 }),
  .out1({ S2137 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1024_ (
  .in1({ S2137, S2136 }),
  .out1({ S2138 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_798_ (
  .in1({ S2138, DP_LGU1_in1_2 }),
  .out1({ S2139 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_799_ (
  .in1({ S2139, S2134 }),
  .out1({ S2140 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_800_ (
  .in1({ S2140, DP_LGU1_in1_3 }),
  .out1({ S2141 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1025_ (
  .in1({ S1732, DP_LGU1_in1_3 }),
  .out1({ S2142 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_323_ (
  .in1({ S2142 }),
  .out1({ S2143 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_801_ (
  .in1({ S2143, S2141 }),
  .out1({ S1621 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_802_ (
  .in1({ S1644, DP_LGU1_in1_4 }),
  .out1({ S2144 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_803_ (
  .in1({ S2144, S1777 }),
  .out1({ S2145 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_804_ (
  .in1({ S2117, S1784 }),
  .out1({ S2146 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_805_ (
  .in1({ S2146, S2120 }),
  .out1({ S2147 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_806_ (
  .in1({ S2147, S2145 }),
  .out1({ S2148 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_807_ (
  .in1({ S2148, CU_NOT }),
  .out1({ S2149 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_324_ (
  .in1({ S2149 }),
  .out1({ S2150 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1026_ (
  .in1({ CU_NOT, DP_AC_out_8 }),
  .out1({ S2151 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_325_ (
  .in1({ S2151 }),
  .out1({ S2152 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_808_ (
  .in1({ S2152, CU_AND }),
  .out1({ S2153 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1027_ (
  .in1({ S2153, S2150 }),
  .out1({ S2154 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1028_ (
  .in1({ DP_LGU1_in1_8, CU_AND }),
  .out1({ S2155 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_326_ (
  .in1({ S2155 }),
  .out1({ S2156 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1029_ (
  .in1({ S2156, DP_AC_out_8 }),
  .out1({ S2157 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1030_ (
  .in1({ S2157, S2154 }),
  .out1({ S1600 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_809_ (
  .in1({ S1847, DP_LGU1_in1_3 }),
  .out1({ S2158 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_327_ (
  .in1({ S2158 }),
  .out1({ S1622 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1031_ (
  .in1({ S1823, S1815 }),
  .out1({ S2159 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1032_ (
  .in1({ S2159, S1654 }),
  .out1({ S2160 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1033_ (
  .in1({ S2106, DP_LGU1_in1_1 }),
  .out1({ S2161 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1034_ (
  .in1({ S2161, S2160 }),
  .out1({ S2162 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1035_ (
  .in1({ S2162, S1657 }),
  .out1({ S2163 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1036_ (
  .in1({ S2036, DP_LGU1_in1_2 }),
  .out1({ S2164 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1037_ (
  .in1({ S2164, S2163 }),
  .out1({ S2165 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1038_ (
  .in1({ S2165, S1658 }),
  .out1({ S2166 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1039_ (
  .in1({ S1854, DP_LGU1_in1_3 }),
  .out1({ S2167 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1040_ (
  .in1({ S2167, S2166 }),
  .out1({ S1623 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1041_ (
  .in1({ CU_NOT, DP_AC_out_9 }),
  .out1({ S2168 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_328_ (
  .in1({ S2168 }),
  .out1({ S2169 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_810_ (
  .in1({ S2169, CU_AND }),
  .out1({ S2170 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1042_ (
  .in1({ S2116, S1872 }),
  .out1({ S2171 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1043_ (
  .in1({ S1777, DP_AC_out_15 }),
  .out1({ S2172 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_811_ (
  .in1({ S2116, DP_AC_out_15 }),
  .out1({ S2173 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_812_ (
  .in1({ S2173, S1778 }),
  .out1({ S2174 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1044_ (
  .in1({ S2174, S2171 }),
  .out1({ S2175 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_813_ (
  .in1({ S1795, S1645 }),
  .out1({ S2176 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_814_ (
  .in1({ S2176, CU_NOT }),
  .out1({ S2177 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1045_ (
  .in1({ S2177, S2175 }),
  .out1({ S2178 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1046_ (
  .in1({ S2178, S2170 }),
  .out1({ S2179 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1047_ (
  .in1({ DP_LGU1_in1_9, CU_AND }),
  .out1({ S2180 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_329_ (
  .in1({ S2180 }),
  .out1({ S2181 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1048_ (
  .in1({ S2181, DP_AC_out_9 }),
  .out1({ S2182 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1049_ (
  .in1({ S2182, S2179 }),
  .out1({ S1601 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1050_ (
  .in1({ S1913, S1658 }),
  .out1({ S1624 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1051_ (
  .in1({ S1746, S1742 }),
  .out1({ S2183 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1052_ (
  .in1({ S2183, S1654 }),
  .out1({ S2184 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1053_ (
  .in1({ S2135, DP_LGU1_in1_1 }),
  .out1({ S2185 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1054_ (
  .in1({ S2185, S2184 }),
  .out1({ S2186 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1055_ (
  .in1({ S2186, S1657 }),
  .out1({ S2187 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1056_ (
  .in1({ S2072, DP_LGU1_in1_2 }),
  .out1({ S2188 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1057_ (
  .in1({ S2188, S2187 }),
  .out1({ S2189 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1058_ (
  .in1({ S2189, S1658 }),
  .out1({ S2190 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1059_ (
  .in1({ S1922, DP_LGU1_in1_3 }),
  .out1({ S2191 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1060_ (
  .in1({ S2191, S2190 }),
  .out1({ S1625 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1061_ (
  .in1({ CU_NOT, DP_AC_out_10 }),
  .out1({ S2192 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_330_ (
  .in1({ S2192 }),
  .out1({ S2193 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_815_ (
  .in1({ S2193, CU_AND }),
  .out1({ S2194 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1062_ (
  .in1({ S2116, S1937 }),
  .out1({ S2195 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1063_ (
  .in1({ S2195, S2174 }),
  .out1({ S2196 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_816_ (
  .in1({ S1795, S1646 }),
  .out1({ S2197 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_817_ (
  .in1({ S2197, CU_NOT }),
  .out1({ S2198 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1064_ (
  .in1({ S2198, S2196 }),
  .out1({ S2199 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1065_ (
  .in1({ S2199, S2194 }),
  .out1({ S2200 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1066_ (
  .in1({ DP_LGU1_in1_10, CU_AND }),
  .out1({ S2201 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_331_ (
  .in1({ S2201 }),
  .out1({ S2202 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1067_ (
  .in1({ S2202, DP_AC_out_10 }),
  .out1({ S2203 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1068_ (
  .in1({ S2203, S2200 }),
  .out1({ S1587 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_818_ (
  .in1({ S1964, DP_LGU1_in1_3 }),
  .out1({ S2204 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_332_ (
  .in1({ S2204 }),
  .out1({ S1626 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_819_ (
  .in1({ S1830, S1822 }),
  .out1({ S2205 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1069_ (
  .in1({ S2205, S1654 }),
  .out1({ S2206 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1070_ (
  .in1({ S2159, DP_LGU1_in1_1 }),
  .out1({ S2207 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1071_ (
  .in1({ S2207, S2206 }),
  .out1({ S2208 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1072_ (
  .in1({ S2208, S1657 }),
  .out1({ S2209 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1073_ (
  .in1({ S2109, DP_LGU1_in1_2 }),
  .out1({ S2210 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1074_ (
  .in1({ S2210, S2209 }),
  .out1({ S2211 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1075_ (
  .in1({ S2211, S1658 }),
  .out1({ S2212 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1076_ (
  .in1({ S1971, DP_LGU1_in1_3 }),
  .out1({ S2213 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1077_ (
  .in1({ S2213, S2212 }),
  .out1({ S1627 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1078_ (
  .in1({ CU_NOT, DP_AC_out_11 }),
  .out1({ S2214 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_333_ (
  .in1({ S2214 }),
  .out1({ S2215 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_820_ (
  .in1({ S2215, CU_AND }),
  .out1({ S2216 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1079_ (
  .in1({ S2116, S1981 }),
  .out1({ S2217 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1080_ (
  .in1({ S2217, S2174 }),
  .out1({ S2218 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_821_ (
  .in1({ S1795, S1647 }),
  .out1({ S2219 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_822_ (
  .in1({ S2219, CU_NOT }),
  .out1({ S2220 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1081_ (
  .in1({ S2220, S2218 }),
  .out1({ S2221 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1082_ (
  .in1({ S2221, S2216 }),
  .out1({ S2222 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1083_ (
  .in1({ DP_LGU1_in1_11, CU_AND }),
  .out1({ S2223 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_334_ (
  .in1({ S2223 }),
  .out1({ S2224 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1084_ (
  .in1({ S2224, DP_AC_out_11 }),
  .out1({ S2225 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1085_ (
  .in1({ S2225, S2222 }),
  .out1({ S1588 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1086_ (
  .in1({ S1997, S1658 }),
  .out1({ S1628 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1087_ (
  .in1({ S1755, S1748 }),
  .out1({ S2226 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1088_ (
  .in1({ S2226, S1654 }),
  .out1({ S2227 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1089_ (
  .in1({ S2183, DP_LGU1_in1_1 }),
  .out1({ S2228 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1090_ (
  .in1({ S2228, S2227 }),
  .out1({ S2229 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1091_ (
  .in1({ S2229, S1657 }),
  .out1({ S2230 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1092_ (
  .in1({ S2138, DP_LGU1_in1_2 }),
  .out1({ S2231 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1093_ (
  .in1({ S2231, S2230 }),
  .out1({ S2232 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1094_ (
  .in1({ S2232, S1658 }),
  .out1({ S2233 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1095_ (
  .in1({ S2006, DP_LGU1_in1_3 }),
  .out1({ S2234 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1096_ (
  .in1({ S2234, S2233 }),
  .out1({ S1629 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1097_ (
  .in1({ CU_NOT, DP_AC_out_12 }),
  .out1({ S2235 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_335_ (
  .in1({ S2235 }),
  .out1({ S2236 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_823_ (
  .in1({ S2236, CU_AND }),
  .out1({ S2237 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1098_ (
  .in1({ S2116, S2014 }),
  .out1({ S2238 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1099_ (
  .in1({ S2238, S2174 }),
  .out1({ S2239 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_824_ (
  .in1({ S1795, S1648 }),
  .out1({ S2240 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_825_ (
  .in1({ S2240, CU_NOT }),
  .out1({ S2241 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1100_ (
  .in1({ S2241, S2239 }),
  .out1({ S2242 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1101_ (
  .in1({ S2242, S2237 }),
  .out1({ S2243 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1102_ (
  .in1({ DP_LGU1_in1_12, CU_AND }),
  .out1({ S2244 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_336_ (
  .in1({ S2244 }),
  .out1({ S2245 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1103_ (
  .in1({ S2245, DP_AC_out_12 }),
  .out1({ S2246 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1104_ (
  .in1({ S2246, S2243 }),
  .out1({ S1589 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1105_ (
  .in1({ S2030, S1658 }),
  .out1({ S1630 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_826_ (
  .in1({ S1839, S1829 }),
  .out1({ S2247 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1106_ (
  .in1({ S2247, S1654 }),
  .out1({ S2248 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1107_ (
  .in1({ S2205, DP_LGU1_in1_1 }),
  .out1({ S2249 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1108_ (
  .in1({ S2249, S2248 }),
  .out1({ S2250 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1109_ (
  .in1({ S2250, S1657 }),
  .out1({ S2251 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1110_ (
  .in1({ S2162, DP_LGU1_in1_2 }),
  .out1({ S2252 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1111_ (
  .in1({ S2252, S2251 }),
  .out1({ S2253 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1112_ (
  .in1({ S2253, S1658 }),
  .out1({ S2254 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1113_ (
  .in1({ S2039, DP_LGU1_in1_3 }),
  .out1({ S2255 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1114_ (
  .in1({ S2255, S2254 }),
  .out1({ S1631 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1115_ (
  .in1({ CU_NOT, DP_AC_out_13 }),
  .out1({ S2256 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_337_ (
  .in1({ S2256 }),
  .out1({ S2257 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_827_ (
  .in1({ S2257, CU_AND }),
  .out1({ S2258 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1116_ (
  .in1({ S2116, S2050 }),
  .out1({ S2259 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1117_ (
  .in1({ S2259, S2174 }),
  .out1({ S2260 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_828_ (
  .in1({ S1795, S1649 }),
  .out1({ S2261 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_829_ (
  .in1({ S2261, CU_NOT }),
  .out1({ S2262 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1118_ (
  .in1({ S2262, S2260 }),
  .out1({ S2263 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1119_ (
  .in1({ S2263, S2258 }),
  .out1({ S2264 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1120_ (
  .in1({ DP_LGU1_in1_13, CU_AND }),
  .out1({ S2265 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_338_ (
  .in1({ S2265 }),
  .out1({ S2266 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1121_ (
  .in1({ S2266, DP_AC_out_13 }),
  .out1({ S2267 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1122_ (
  .in1({ S2267, S2264 }),
  .out1({ S1590 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1123_ (
  .in1({ S2066, S1658 }),
  .out1({ S1632 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1124_ (
  .in1({ S1761, S1757 }),
  .out1({ S2268 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1125_ (
  .in1({ S2268, S1654 }),
  .out1({ S2269 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1126_ (
  .in1({ S2226, DP_LGU1_in1_1 }),
  .out1({ S2270 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1127_ (
  .in1({ S2270, S2269 }),
  .out1({ S2271 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1128_ (
  .in1({ S2271, S1657 }),
  .out1({ S2272 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1129_ (
  .in1({ S2186, DP_LGU1_in1_2 }),
  .out1({ S2273 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1130_ (
  .in1({ S2273, S2272 }),
  .out1({ S2274 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1131_ (
  .in1({ S2274, S1658 }),
  .out1({ S2275 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1132_ (
  .in1({ S2075, DP_LGU1_in1_3 }),
  .out1({ S2276 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1133_ (
  .in1({ S2276, S2275 }),
  .out1({ S1633 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1134_ (
  .in1({ CU_NOT, DP_AC_out_14 }),
  .out1({ S2277 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_339_ (
  .in1({ S2277 }),
  .out1({ S2278 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_830_ (
  .in1({ S2278, CU_AND }),
  .out1({ S2279 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1135_ (
  .in1({ S2116, S2086 }),
  .out1({ S2280 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1136_ (
  .in1({ S2280, S2174 }),
  .out1({ S2281 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_831_ (
  .in1({ S1795, S1650 }),
  .out1({ S2282 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_832_ (
  .in1({ S2282, CU_NOT }),
  .out1({ S2283 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1137_ (
  .in1({ S2283, S2281 }),
  .out1({ S2284 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1138_ (
  .in1({ S2284, S2279 }),
  .out1({ S2285 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1139_ (
  .in1({ DP_LGU1_in1_14, CU_AND }),
  .out1({ S2286 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_340_ (
  .in1({ S2286 }),
  .out1({ S2287 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1140_ (
  .in1({ S2287, DP_AC_out_14 }),
  .out1({ S2288 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1141_ (
  .in1({ S2288, S2285 }),
  .out1({ S1591 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1142_ (
  .in1({ S2103, S1658 }),
  .out1({ S1634 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_833_ (
  .in1({ S2112, S1658 }),
  .out1({ S2289 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_834_ (
  .in1({ S2247, S1654 }),
  .out1({ S2290 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1143_ (
  .in1({ S1838, S1654 }),
  .out1({ S2291 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1144_ (
  .in1({ S2291, S1958 }),
  .out1({ S2292 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_835_ (
  .in1({ S2292, S2290 }),
  .out1({ S2293 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_836_ (
  .in1({ S2293, DP_LGU1_in1_2 }),
  .out1({ S2294 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_837_ (
  .in1({ S2208, S1657 }),
  .out1({ S2295 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_838_ (
  .in1({ S2295, S2294 }),
  .out1({ S2296 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_839_ (
  .in1({ S2296, DP_LGU1_in1_3 }),
  .out1({ S2297 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_840_ (
  .in1({ S2297, S2289 }),
  .out1({ S1635 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1145_ (
  .in1({ DP_AC_out_15, DP_LGU1_in1_15 }),
  .out1({ S2298 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1146_ (
  .in1({ S2298, CU_AND }),
  .out1({ S2299 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_341_ (
  .in1({ S2299 }),
  .out1({ S2300 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_841_ (
  .in1({ S1795, S1651 }),
  .out1({ S2301 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1147_ (
  .in1({ S2172, S1662 }),
  .out1({ S2302 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_842_ (
  .in1({ S2302, S2301 }),
  .out1({ S2303 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1148_ (
  .in1({ CU_NOT, DP_AC_out_15 }),
  .out1({ S2304 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_342_ (
  .in1({ S2304 }),
  .out1({ S2305 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_843_ (
  .in1({ S2305, S2303 }),
  .out1({ S2306 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_844_ (
  .in1({ S2306, CU_AND }),
  .out1({ S2307 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_845_ (
  .in1({ S2307, S2300 }),
  .out1({ S1592 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1149_ (
  .in1({ S1773, CU_SHF_0 }),
  .out1({ S2308 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_846_ (
  .in1({ S2308, S1661 }),
  .out1({ S1602 })
);
$mux #( 
  .WIDTH(32'b00000000000000000000000000000001)) 
$mux_1_ (
  .A({ S1605 }),
  .B({ S1603 }),
  .S({ S1604 }),
  .Y({ S1636 })
);
$mux #( 
  .WIDTH(32'b00000000000000000000000000000001)) 
$mux_2_ (
  .A({ S1607 }),
  .B({ S1606 }),
  .S({ S1604 }),
  .Y({ S1637 })
);
$mux #( 
  .WIDTH(32'b00000000000000000000000000000001)) 
$mux_3_ (
  .A({ S1609 }),
  .B({ S1608 }),
  .S({ S1604 }),
  .Y({ S1638 })
);
$mux #( 
  .WIDTH(32'b00000000000000000000000000000001)) 
$mux_4_ (
  .A({ S1611 }),
  .B({ S1610 }),
  .S({ S1604 }),
  .Y({ S1639 })
);
$mux #( 
  .WIDTH(32'b00000000000000000000000000000001)) 
$mux_5_ (
  .A({ S1613 }),
  .B({ S1612 }),
  .S({ S1604 }),
  .Y({ S1640 })
);
$mux #( 
  .WIDTH(32'b00000000000000000000000000000001)) 
$mux_6_ (
  .A({ S1615 }),
  .B({ S1614 }),
  .S({ S1604 }),
  .Y({ S1641 })
);
$mux #( 
  .WIDTH(32'b00000000000000000000000000000001)) 
$mux_7_ (
  .A({ S1617 }),
  .B({ S1616 }),
  .S({ S1604 }),
  .Y({ S1642 })
);
$mux #( 
  .WIDTH(32'b00000000000000000000000000000001)) 
$mux_8_ (
  .A({ S1619 }),
  .B({ S1618 }),
  .S({ S1604 }),
  .Y({ S1643 })
);
$mux #( 
  .WIDTH(32'b00000000000000000000000000000001)) 
$mux_9_ (
  .A({ S1621 }),
  .B({ S1620 }),
  .S({ S1604 }),
  .Y({ S1644 })
);
$mux #( 
  .WIDTH(32'b00000000000000000000000000000001)) 
$mux_10_ (
  .A({ S1623 }),
  .B({ S1622 }),
  .S({ S1604 }),
  .Y({ S1645 })
);
$mux #( 
  .WIDTH(32'b00000000000000000000000000000001)) 
$mux_11_ (
  .A({ S1625 }),
  .B({ S1624 }),
  .S({ S1604 }),
  .Y({ S1646 })
);
$mux #( 
  .WIDTH(32'b00000000000000000000000000000001)) 
$mux_12_ (
  .A({ S1627 }),
  .B({ S1626 }),
  .S({ S1604 }),
  .Y({ S1647 })
);
$mux #( 
  .WIDTH(32'b00000000000000000000000000000001)) 
$mux_13_ (
  .A({ S1629 }),
  .B({ S1628 }),
  .S({ S1604 }),
  .Y({ S1648 })
);
$mux #( 
  .WIDTH(32'b00000000000000000000000000000001)) 
$mux_14_ (
  .A({ S1631 }),
  .B({ S1630 }),
  .S({ S1604 }),
  .Y({ S1649 })
);
$mux #( 
  .WIDTH(32'b00000000000000000000000000000001)) 
$mux_15_ (
  .A({ S1633 }),
  .B({ S1632 }),
  .S({ S1604 }),
  .Y({ S1650 })
);
$mux #( 
  .WIDTH(32'b00000000000000000000000000000001)) 
$mux_16_ (
  .A({ S1635 }),
  .B({ S1634 }),
  .S({ S1604 }),
  .Y({ S1651 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__35_ (
  .D({ S1586 }),
  .E({ S1602 }),
  .Q({ DP_LGU1_out_0 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__36_ (
  .D({ S1593 }),
  .E({ S1602 }),
  .Q({ DP_LGU1_out_1 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__37_ (
  .D({ S1594 }),
  .E({ S1602 }),
  .Q({ DP_LGU1_out_2 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__38_ (
  .D({ S1595 }),
  .E({ S1602 }),
  .Q({ DP_LGU1_out_3 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__39_ (
  .D({ S1596 }),
  .E({ S1602 }),
  .Q({ DP_LGU1_out_4 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__40_ (
  .D({ S1597 }),
  .E({ S1602 }),
  .Q({ DP_LGU1_out_5 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__41_ (
  .D({ S1598 }),
  .E({ S1602 }),
  .Q({ DP_LGU1_out_6 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__42_ (
  .D({ S1599 }),
  .E({ S1602 }),
  .Q({ DP_LGU1_out_7 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__43_ (
  .D({ S1600 }),
  .E({ S1602 }),
  .Q({ DP_LGU1_out_8 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__44_ (
  .D({ S1601 }),
  .E({ S1602 }),
  .Q({ DP_LGU1_out_9 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__45_ (
  .D({ S1587 }),
  .E({ S1602 }),
  .Q({ DP_LGU1_out_10 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__46_ (
  .D({ S1588 }),
  .E({ S1602 }),
  .Q({ DP_LGU1_out_11 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__47_ (
  .D({ S1589 }),
  .E({ S1602 }),
  .Q({ DP_LGU1_out_12 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__48_ (
  .D({ S1590 }),
  .E({ S1602 }),
  .Q({ DP_LGU1_out_13 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__49_ (
  .D({ S1591 }),
  .E({ S1602 }),
  .Q({ DP_LGU1_out_14 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__50_ (
  .D({ S1592 }),
  .E({ S1602 }),
  .Q({ DP_LGU1_N })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_343_ (
  .in1({ CU_ldOF }),
  .out1({ S2313 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_847_ (
  .in1({ CU_ldOF, S13 }),
  .out1({ S2314 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1150_ (
  .in1({ S2314, DP_IMM1_in1_0 }),
  .out1({ S2315 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_848_ (
  .in1({ S2313, S14 }),
  .out1({ S2316 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1151_ (
  .in1({ S2316, DP_OF_in_0 }),
  .out1({ S2317 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1152_ (
  .in1({ S2317, S2315 }),
  .out1({ S2309 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1153_ (
  .in1({ S2314, DP_IMM1_in1_1 }),
  .out1({ S2318 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1154_ (
  .in1({ S2316, DP_OF_in_1 }),
  .out1({ S2319 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1155_ (
  .in1({ S2319, S2318 }),
  .out1({ S2310 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1156_ (
  .in1({ S2314, DP_IMM1_in1_2 }),
  .out1({ S2320 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1157_ (
  .in1({ S2316, DP_OF_in_2 }),
  .out1({ S2321 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1158_ (
  .in1({ S2321, S2320 }),
  .out1({ S2311 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1159_ (
  .in1({ S2314, DP_IMM1_in1_3 }),
  .out1({ S2322 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1160_ (
  .in1({ S2316, DP_OF_in_3 }),
  .out1({ S2323 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1161_ (
  .in1({ S2323, S2322 }),
  .out1({ S2312 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_51_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2309 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IMM1_in1_0 }),
  .Si({ S3340 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_52_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2310 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IMM1_in1_1 }),
  .Si({ S3339 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_53_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2311 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IMM1_in1_2 }),
  .Si({ S3338 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_54_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2312 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IMM1_in1_3 }),
  .Si({ S3359 }),
  .global_reset({ 1'b0 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_344_ (
  .in1({ CU_ldPC }),
  .out1({ S2341 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_849_ (
  .in1({ CU_ldPC, S15 }),
  .out1({ S2342 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1162_ (
  .in1({ S2342, DP_INC_1_in_0 }),
  .out1({ S2343 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_850_ (
  .in1({ S2341, S16 }),
  .out1({ S2344 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1163_ (
  .in1({ S2344, DP_PC_in_0 }),
  .out1({ S2345 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1164_ (
  .in1({ S2345, S2343 }),
  .out1({ S2324 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1165_ (
  .in1({ S2342, DP_INC_1_in_1 }),
  .out1({ S2346 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1166_ (
  .in1({ S2344, DP_PC_in_1 }),
  .out1({ S2347 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1167_ (
  .in1({ S2347, S2346 }),
  .out1({ S2325 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1168_ (
  .in1({ S2342, DP_INC_1_in_2 }),
  .out1({ S2348 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1169_ (
  .in1({ S2344, DP_PC_in_2 }),
  .out1({ S2349 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1170_ (
  .in1({ S2349, S2348 }),
  .out1({ S2326 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1171_ (
  .in1({ S2342, DP_INC_1_in_3 }),
  .out1({ S2350 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1172_ (
  .in1({ S2344, DP_PC_in_3 }),
  .out1({ S2351 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1173_ (
  .in1({ S2351, S2350 }),
  .out1({ S2327 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1174_ (
  .in1({ S2342, DP_INC_1_in_4 }),
  .out1({ S2352 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1175_ (
  .in1({ S2344, DP_PC_in_4 }),
  .out1({ S2353 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1176_ (
  .in1({ S2353, S2352 }),
  .out1({ S2328 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1177_ (
  .in1({ S2342, DP_INC_1_in_5 }),
  .out1({ S2354 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1178_ (
  .in1({ S2344, DP_PC_in_5 }),
  .out1({ S2355 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1179_ (
  .in1({ S2355, S2354 }),
  .out1({ S2329 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1180_ (
  .in1({ S2342, DP_INC_1_in_6 }),
  .out1({ S2356 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1181_ (
  .in1({ S2344, DP_PC_in_6 }),
  .out1({ S2357 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1182_ (
  .in1({ S2357, S2356 }),
  .out1({ S2330 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1183_ (
  .in1({ S2342, DP_INC_1_in_7 }),
  .out1({ S2358 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1184_ (
  .in1({ S2344, DP_PC_in_7 }),
  .out1({ S2359 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1185_ (
  .in1({ S2359, S2358 }),
  .out1({ S2331 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1186_ (
  .in1({ S2342, DP_INC_1_in_8 }),
  .out1({ S2360 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1187_ (
  .in1({ S2344, DP_PC_in_8 }),
  .out1({ S2361 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1188_ (
  .in1({ S2361, S2360 }),
  .out1({ S2332 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1189_ (
  .in1({ S2342, DP_INC_1_in_9 }),
  .out1({ S2362 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1190_ (
  .in1({ S2344, DP_PC_in_9 }),
  .out1({ S2363 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1191_ (
  .in1({ S2363, S2362 }),
  .out1({ S2333 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1192_ (
  .in1({ S2342, DP_INC_1_in_10 }),
  .out1({ S2364 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1193_ (
  .in1({ S2344, DP_PC_in_10 }),
  .out1({ S2365 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1194_ (
  .in1({ S2365, S2364 }),
  .out1({ S2334 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1195_ (
  .in1({ S2342, DP_INC_1_in_11 }),
  .out1({ S2366 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1196_ (
  .in1({ S2344, DP_PC_in_11 }),
  .out1({ S2367 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1197_ (
  .in1({ S2367, S2366 }),
  .out1({ S2335 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1198_ (
  .in1({ S2342, DP_INC_1_in_12 }),
  .out1({ S2368 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1199_ (
  .in1({ S2344, DP_PC_in_12 }),
  .out1({ S2369 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1200_ (
  .in1({ S2369, S2368 }),
  .out1({ S2336 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1201_ (
  .in1({ S2342, DP_INC_1_in_13 }),
  .out1({ S2370 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1202_ (
  .in1({ S2344, DP_PC_in_13 }),
  .out1({ S2371 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1203_ (
  .in1({ S2371, S2370 }),
  .out1({ S2337 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1204_ (
  .in1({ S2342, DP_INC_1_in_14 }),
  .out1({ S2372 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1205_ (
  .in1({ S2344, DP_PC_in_14 }),
  .out1({ S2373 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1206_ (
  .in1({ S2373, S2372 }),
  .out1({ S2338 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1207_ (
  .in1({ S2342, DP_INC_1_in_15 }),
  .out1({ S2374 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1208_ (
  .in1({ S2344, DP_PC_in_15 }),
  .out1({ S2340 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1209_ (
  .in1({ S2340, S2374 }),
  .out1({ S2339 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_55_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2324 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_0 }),
  .Si({ S3355 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_56_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2325 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_1 }),
  .Si({ S3354 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_57_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2326 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_2 }),
  .Si({ S3353 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_58_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2327 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_3 }),
  .Si({ S3352 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_59_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2328 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_4 }),
  .Si({ S3351 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_60_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2329 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_5 }),
  .Si({ S3350 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_61_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2330 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_6 }),
  .Si({ S3349 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_62_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2331 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_7 }),
  .Si({ S3348 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_63_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2332 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_8 }),
  .Si({ S3347 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_64_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2333 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_9 }),
  .Si({ S3346 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_65_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2334 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_10 }),
  .Si({ S3345 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_66_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2335 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_11 }),
  .Si({ S3344 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_67_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2336 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_12 }),
  .Si({ S3343 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_68_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2337 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_13 }),
  .Si({ S3342 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_69_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2338 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_14 }),
  .Si({ S3341 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_70_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2339 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_15 }),
  .Si({ S3360 }),
  .global_reset({ 1'b0 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_345_ (
  .in1({ DP_SR_C_out }),
  .out1({ S2377 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1210_ (
  .in1({ DP_SR_C_in, CU_ldSR_1 }),
  .out1({ S2378 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_346_ (
  .in1({ S2378 }),
  .out1({ S2379 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_851_ (
  .in1({ S2377, CU_ldSR_1 }),
  .out1({ S2380 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_852_ (
  .in1({ S2380, S2379 }),
  .out1({ S2376 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_853_ (
  .in1({ S2376, S17 }),
  .out1({ S2375 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_71_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2375 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_SR_C_out }),
  .Si({ S3361 }),
  .global_reset({ 1'b0 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_347_ (
  .in1({ DP_SR_N_out }),
  .out1({ S2383 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1211_ (
  .in1({ DP_SR_N_in, CU_ldSR_2 }),
  .out1({ S2384 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_348_ (
  .in1({ S2384 }),
  .out1({ S2385 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_854_ (
  .in1({ S2383, CU_ldSR_2 }),
  .out1({ S2386 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_855_ (
  .in1({ S2386, S2385 }),
  .out1({ S2382 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_856_ (
  .in1({ S2382, S18 }),
  .out1({ S2381 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_72_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2381 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_SR_N_out }),
  .Si({ S3362 }),
  .global_reset({ 1'b0 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_349_ (
  .in1({ DP_SR_V_out }),
  .out1({ S2389 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1212_ (
  .in1({ DP_SR_V_in, CU_ldSR_0 }),
  .out1({ S2390 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_350_ (
  .in1({ S2390 }),
  .out1({ S2391 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_857_ (
  .in1({ S2389, CU_ldSR_0 }),
  .out1({ S2392 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_858_ (
  .in1({ S2392, S2391 }),
  .out1({ S2388 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_859_ (
  .in1({ S2388, S19 }),
  .out1({ S2387 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_73_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2387 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_SR_V_out }),
  .Si({ S3363 }),
  .global_reset({ 1'b0 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_351_ (
  .in1({ DP_SR_Z_out }),
  .out1({ S2395 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1213_ (
  .in1({ DP_SR_Z_in, CU_ldSR_3 }),
  .out1({ S2396 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_352_ (
  .in1({ S2396 }),
  .out1({ S2397 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_860_ (
  .in1({ S2395, CU_ldSR_3 }),
  .out1({ S2398 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_861_ (
  .in1({ S2398, S2397 }),
  .out1({ S2394 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_862_ (
  .in1({ S2394, S20 }),
  .out1({ S2393 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_74_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2393 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_SR_Z_out }),
  .Si({ S3364 }),
  .global_reset({ 1'b0 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_353_ (
  .in1({ CU_sel1_ARU }),
  .out1({ S2416 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1214_ (
  .in1({ CU_sel1_ARU, S3 }),
  .out1({ S2417 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1215_ (
  .in1({ S2416, DP_LGU1_in1_0 }),
  .out1({ S2418 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1216_ (
  .in1({ S2418, S2417 }),
  .out1({ S2399 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1217_ (
  .in1({ S21, CU_sel1_ARU }),
  .out1({ S2419 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1218_ (
  .in1({ DP_LGU1_in1_1, S2416 }),
  .out1({ S2420 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1219_ (
  .in1({ S2420, S2419 }),
  .out1({ S2406 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1220_ (
  .in1({ S22, CU_sel1_ARU }),
  .out1({ S2421 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1221_ (
  .in1({ DP_LGU1_in1_2, S2416 }),
  .out1({ S2422 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1222_ (
  .in1({ S2422, S2421 }),
  .out1({ S2407 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1223_ (
  .in1({ S23, CU_sel1_ARU }),
  .out1({ S2423 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1224_ (
  .in1({ DP_LGU1_in1_3, S2416 }),
  .out1({ S2424 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1225_ (
  .in1({ S2424, S2423 }),
  .out1({ S2408 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1226_ (
  .in1({ S24, CU_sel1_ARU }),
  .out1({ S2425 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1227_ (
  .in1({ DP_LGU1_in1_4, S2416 }),
  .out1({ S2426 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1228_ (
  .in1({ S2426, S2425 }),
  .out1({ S2409 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1229_ (
  .in1({ S25, CU_sel1_ARU }),
  .out1({ S2427 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1230_ (
  .in1({ DP_LGU1_in1_5, S2416 }),
  .out1({ S2428 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1231_ (
  .in1({ S2428, S2427 }),
  .out1({ S2410 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1232_ (
  .in1({ S26, CU_sel1_ARU }),
  .out1({ S2429 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1233_ (
  .in1({ DP_LGU1_in1_6, S2416 }),
  .out1({ S2430 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1234_ (
  .in1({ S2430, S2429 }),
  .out1({ S2411 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1235_ (
  .in1({ S27, CU_sel1_ARU }),
  .out1({ S2431 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1236_ (
  .in1({ DP_LGU1_in1_7, S2416 }),
  .out1({ S2432 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1237_ (
  .in1({ S2432, S2431 }),
  .out1({ S2412 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1238_ (
  .in1({ S28, CU_sel1_ARU }),
  .out1({ S2433 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1239_ (
  .in1({ DP_LGU1_in1_8, S2416 }),
  .out1({ S2434 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1240_ (
  .in1({ S2434, S2433 }),
  .out1({ S2413 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1241_ (
  .in1({ S29, CU_sel1_ARU }),
  .out1({ S2435 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1242_ (
  .in1({ DP_LGU1_in1_9, S2416 }),
  .out1({ S2436 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1243_ (
  .in1({ S2436, S2435 }),
  .out1({ S2414 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1244_ (
  .in1({ S30, CU_sel1_ARU }),
  .out1({ S2437 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1245_ (
  .in1({ DP_LGU1_in1_10, S2416 }),
  .out1({ S2438 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1246_ (
  .in1({ S2438, S2437 }),
  .out1({ S2400 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1247_ (
  .in1({ S31, CU_sel1_ARU }),
  .out1({ S2439 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1248_ (
  .in1({ DP_LGU1_in1_11, S2416 }),
  .out1({ S2440 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1249_ (
  .in1({ S2440, S2439 }),
  .out1({ S2401 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1250_ (
  .in1({ S32, CU_sel1_ARU }),
  .out1({ S2441 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1251_ (
  .in1({ DP_LGU1_in1_12, S2416 }),
  .out1({ S2442 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1252_ (
  .in1({ S2442, S2441 }),
  .out1({ S2402 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1253_ (
  .in1({ S33, CU_sel1_ARU }),
  .out1({ S2443 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1254_ (
  .in1({ DP_LGU1_in1_13, S2416 }),
  .out1({ S2444 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1255_ (
  .in1({ S2444, S2443 }),
  .out1({ S2403 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1256_ (
  .in1({ S34, CU_sel1_ARU }),
  .out1({ S2445 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1257_ (
  .in1({ DP_LGU1_in1_14, S2416 }),
  .out1({ S2446 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1258_ (
  .in1({ S2446, S2445 }),
  .out1({ S2404 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1259_ (
  .in1({ S35, CU_sel1_ARU }),
  .out1({ S2447 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1260_ (
  .in1({ DP_LGU1_in1_15, S2416 }),
  .out1({ S2448 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1261_ (
  .in1({ S2448, S2447 }),
  .out1({ S2405 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_863_ (
  .in1({ CU_selARU_SR, CU_sel1_ARU }),
  .out1({ S2415 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__51_ (
  .D({ S2399 }),
  .E({ S2415 }),
  .Q({ DP_ARU1_in1_0 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__52_ (
  .D({ S2406 }),
  .E({ S2415 }),
  .Q({ DP_ARU1_in1_1 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__53_ (
  .D({ S2407 }),
  .E({ S2415 }),
  .Q({ DP_ARU1_in1_2 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__54_ (
  .D({ S2408 }),
  .E({ S2415 }),
  .Q({ DP_ARU1_in1_3 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__55_ (
  .D({ S2409 }),
  .E({ S2415 }),
  .Q({ DP_ARU1_in1_4 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__56_ (
  .D({ S2410 }),
  .E({ S2415 }),
  .Q({ DP_ARU1_in1_5 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__57_ (
  .D({ S2411 }),
  .E({ S2415 }),
  .Q({ DP_ARU1_in1_6 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__58_ (
  .D({ S2412 }),
  .E({ S2415 }),
  .Q({ DP_ARU1_in1_7 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__59_ (
  .D({ S2413 }),
  .E({ S2415 }),
  .Q({ DP_ARU1_in1_8 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__60_ (
  .D({ S2414 }),
  .E({ S2415 }),
  .Q({ DP_ARU1_in1_9 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__61_ (
  .D({ S2400 }),
  .E({ S2415 }),
  .Q({ DP_ARU1_in1_10 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__62_ (
  .D({ S2401 }),
  .E({ S2415 }),
  .Q({ DP_ARU1_in1_11 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__63_ (
  .D({ S2402 }),
  .E({ S2415 }),
  .Q({ DP_ARU1_in1_12 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__64_ (
  .D({ S2403 }),
  .E({ S2415 }),
  .Q({ DP_ARU1_in1_13 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__65_ (
  .D({ S2404 }),
  .E({ S2415 }),
  .Q({ DP_ARU1_in1_14 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__66_ (
  .D({ S2405 }),
  .E({ S2415 }),
  .Q({ DP_ARU1_in1_15 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_354_ (
  .in1({ 1'bz }),
  .out1({ S2454 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_355_ (
  .in1({ 1'bz }),
  .out1({ S2455 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_356_ (
  .in1({ CU_selLGU_SR }),
  .out1({ S2456 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_357_ (
  .in1({ CU_inst_0 }),
  .out1({ S2457 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_358_ (
  .in1({ 1'bz }),
  .out1({ S2458 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_359_ (
  .in1({ 1'bz }),
  .out1({ S2459 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_360_ (
  .in1({ CU_inst_1 }),
  .out1({ S2460 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_361_ (
  .in1({ 1'bz }),
  .out1({ S2461 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_362_ (
  .in1({ DP_LGU1_N }),
  .out1({ S2462 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_363_ (
  .in1({ CU_inst_2 }),
  .out1({ S2463 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_364_ (
  .in1({ 1'bz }),
  .out1({ S2464 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_365_ (
  .in1({ DP_LGU1_Z }),
  .out1({ S2465 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_366_ (
  .in1({ CU_inst_3 }),
  .out1({ S2466 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_367_ (
  .in1({ 1'bz }),
  .out1({ S2467 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_864_ (
  .in1({ CU_selSET_SR, CU_selLGU_SR }),
  .out1({ S2468 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_865_ (
  .in1({ CU_selARU_SR, S2454 }),
  .out1({ S2469 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1262_ (
  .in1({ CU_selARU_SR, DP_ARU1_V }),
  .out1({ S2470 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1263_ (
  .in1({ S2470, S2468 }),
  .out1({ S2471 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_866_ (
  .in1({ S2471, S2469 }),
  .out1({ S2472 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1264_ (
  .in1({ CU_selSET_SR, S2457 }),
  .out1({ S2473 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_867_ (
  .in1({ CU_selSET_SR, S2456 }),
  .out1({ S2474 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1265_ (
  .in1({ S2474, S2455 }),
  .out1({ S2475 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1266_ (
  .in1({ S2475, S2473 }),
  .out1({ S2476 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_868_ (
  .in1({ S2476, S2472 }),
  .out1({ S2449 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_869_ (
  .in1({ S2458, CU_selARU_SR }),
  .out1({ S2477 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1267_ (
  .in1({ DP_ARU1_C, CU_selARU_SR }),
  .out1({ S2478 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1268_ (
  .in1({ S2478, S2468 }),
  .out1({ S2479 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_870_ (
  .in1({ S2479, S2477 }),
  .out1({ S2480 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1269_ (
  .in1({ S2460, CU_selSET_SR }),
  .out1({ S2481 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1270_ (
  .in1({ S2474, S2459 }),
  .out1({ S2482 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1271_ (
  .in1({ S2482, S2481 }),
  .out1({ S2483 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_871_ (
  .in1({ S2483, S2480 }),
  .out1({ S2450 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_872_ (
  .in1({ S2461, CU_selARU_SR }),
  .out1({ S2484 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1272_ (
  .in1({ DP_ARU1_N, CU_selARU_SR }),
  .out1({ S2485 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1273_ (
  .in1({ S2485, S2468 }),
  .out1({ S2486 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_873_ (
  .in1({ S2486, S2484 }),
  .out1({ S2487 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1274_ (
  .in1({ S2463, CU_selSET_SR }),
  .out1({ S2488 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1275_ (
  .in1({ S2474, S2462 }),
  .out1({ S2489 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1276_ (
  .in1({ S2489, S2488 }),
  .out1({ S2490 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_874_ (
  .in1({ S2490, S2487 }),
  .out1({ S2451 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_875_ (
  .in1({ S2464, CU_selARU_SR }),
  .out1({ S2491 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1277_ (
  .in1({ DP_ARU1_Z, CU_selARU_SR }),
  .out1({ S2492 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1278_ (
  .in1({ S2492, S2468 }),
  .out1({ S2493 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_876_ (
  .in1({ S2493, S2491 }),
  .out1({ S2494 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1279_ (
  .in1({ S2466, CU_selSET_SR }),
  .out1({ S2495 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1280_ (
  .in1({ S2474, S2465 }),
  .out1({ S2496 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1281_ (
  .in1({ S2496, S2495 }),
  .out1({ S2497 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_877_ (
  .in1({ S2497, S2494 }),
  .out1({ S2452 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1282_ (
  .in1({ S2468, S2467 }),
  .out1({ S2498 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_878_ (
  .in1({ S2498, CU_selARU_SR }),
  .out1({ S2453 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__67_ (
  .D({ S2449 }),
  .E({ S2453 }),
  .Q({ DP_SR_V_in })
);
$_DLATCH_N_ #() 
$_DLATCH_N__68_ (
  .D({ S2450 }),
  .E({ S2453 }),
  .Q({ DP_SR_C_in })
);
$_DLATCH_N_ #() 
$_DLATCH_N__69_ (
  .D({ S2451 }),
  .E({ S2453 }),
  .Q({ DP_SR_N_in })
);
$_DLATCH_N_ #() 
$_DLATCH_N__70_ (
  .D({ S2452 }),
  .E({ S2453 }),
  .Q({ DP_SR_Z_in })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_368_ (
  .in1({ CU_selIMM_LGU }),
  .out1({ S2516 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1283_ (
  .in1({ CU_selIMM_LGU, DP_IMM1_out_0 }),
  .out1({ S2517 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1284_ (
  .in1({ S2516, dataBus[0] }),
  .out1({ S2518 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1285_ (
  .in1({ S2518, S2517 }),
  .out1({ S2499 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1286_ (
  .in1({ DP_IMM1_out_1, CU_selIMM_LGU }),
  .out1({ S2519 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1287_ (
  .in1({ dataBus[1], S2516 }),
  .out1({ S2520 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1288_ (
  .in1({ S2520, S2519 }),
  .out1({ S2506 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1289_ (
  .in1({ DP_IMM1_out_2, CU_selIMM_LGU }),
  .out1({ S2521 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1290_ (
  .in1({ dataBus[2], S2516 }),
  .out1({ S2522 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1291_ (
  .in1({ S2522, S2521 }),
  .out1({ S2507 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1292_ (
  .in1({ DP_IMM1_out_3, CU_selIMM_LGU }),
  .out1({ S2523 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1293_ (
  .in1({ dataBus[3], S2516 }),
  .out1({ S2524 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1294_ (
  .in1({ S2524, S2523 }),
  .out1({ S2508 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1295_ (
  .in1({ DP_IMM1_out_4, CU_selIMM_LGU }),
  .out1({ S2525 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1296_ (
  .in1({ dataBus[4], S2516 }),
  .out1({ S2526 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1297_ (
  .in1({ S2526, S2525 }),
  .out1({ S2509 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1298_ (
  .in1({ DP_IMM1_out_5, CU_selIMM_LGU }),
  .out1({ S2527 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1299_ (
  .in1({ dataBus[5], S2516 }),
  .out1({ S2528 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1300_ (
  .in1({ S2528, S2527 }),
  .out1({ S2510 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1301_ (
  .in1({ DP_IMM1_out_6, CU_selIMM_LGU }),
  .out1({ S2529 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1302_ (
  .in1({ dataBus[6], S2516 }),
  .out1({ S2530 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1303_ (
  .in1({ S2530, S2529 }),
  .out1({ S2511 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1304_ (
  .in1({ DP_IMM1_out_7, CU_selIMM_LGU }),
  .out1({ S2531 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1305_ (
  .in1({ dataBus[7], S2516 }),
  .out1({ S2532 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1306_ (
  .in1({ S2532, S2531 }),
  .out1({ S2512 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1307_ (
  .in1({ DP_IMM1_out_8, CU_selIMM_LGU }),
  .out1({ S2533 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1308_ (
  .in1({ dataBus[8], S2516 }),
  .out1({ S2534 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1309_ (
  .in1({ S2534, S2533 }),
  .out1({ S2513 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1310_ (
  .in1({ DP_IMM1_out_9, CU_selIMM_LGU }),
  .out1({ S2535 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1311_ (
  .in1({ dataBus[9], S2516 }),
  .out1({ S2536 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1312_ (
  .in1({ S2536, S2535 }),
  .out1({ S2514 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1313_ (
  .in1({ DP_IMM1_out_10, CU_selIMM_LGU }),
  .out1({ S2537 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1314_ (
  .in1({ dataBus[10], S2516 }),
  .out1({ S2538 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1315_ (
  .in1({ S2538, S2537 }),
  .out1({ S2500 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1316_ (
  .in1({ DP_IMM1_out_11, CU_selIMM_LGU }),
  .out1({ S2539 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1317_ (
  .in1({ dataBus[11], S2516 }),
  .out1({ S2540 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1318_ (
  .in1({ S2540, S2539 }),
  .out1({ S2501 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1319_ (
  .in1({ DP_IMM1_out_12, CU_selIMM_LGU }),
  .out1({ S2541 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1320_ (
  .in1({ dataBus[12], S2516 }),
  .out1({ S2542 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1321_ (
  .in1({ S2542, S2541 }),
  .out1({ S2502 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1322_ (
  .in1({ DP_IMM1_out_13, CU_selIMM_LGU }),
  .out1({ S2543 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1323_ (
  .in1({ dataBus[13], S2516 }),
  .out1({ S2544 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1324_ (
  .in1({ S2544, S2543 }),
  .out1({ S2503 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1325_ (
  .in1({ DP_IMM1_out_14, CU_selIMM_LGU }),
  .out1({ S2545 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1326_ (
  .in1({ dataBus[14], S2516 }),
  .out1({ S2546 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1327_ (
  .in1({ S2546, S2545 }),
  .out1({ S2504 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1328_ (
  .in1({ DP_IMM1_out_15, CU_selIMM_LGU }),
  .out1({ S2547 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1329_ (
  .in1({ dataBus[15], S2516 }),
  .out1({ S2548 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1330_ (
  .in1({ S2548, S2547 }),
  .out1({ S2505 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_879_ (
  .in1({ CU_selMEM_LGU, CU_selIMM_LGU }),
  .out1({ S2515 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__71_ (
  .D({ S2499 }),
  .E({ S2515 }),
  .Q({ DP_LGU1_in1_0 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__72_ (
  .D({ S2506 }),
  .E({ S2515 }),
  .Q({ DP_LGU1_in1_1 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__73_ (
  .D({ S2507 }),
  .E({ S2515 }),
  .Q({ DP_LGU1_in1_2 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__74_ (
  .D({ S2508 }),
  .E({ S2515 }),
  .Q({ DP_LGU1_in1_3 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__75_ (
  .D({ S2509 }),
  .E({ S2515 }),
  .Q({ DP_LGU1_in1_4 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__76_ (
  .D({ S2510 }),
  .E({ S2515 }),
  .Q({ DP_LGU1_in1_5 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__77_ (
  .D({ S2511 }),
  .E({ S2515 }),
  .Q({ DP_LGU1_in1_6 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__78_ (
  .D({ S2512 }),
  .E({ S2515 }),
  .Q({ DP_LGU1_in1_7 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__79_ (
  .D({ S2513 }),
  .E({ S2515 }),
  .Q({ DP_LGU1_in1_8 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__80_ (
  .D({ S2514 }),
  .E({ S2515 }),
  .Q({ DP_LGU1_in1_9 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__81_ (
  .D({ S2500 }),
  .E({ S2515 }),
  .Q({ DP_LGU1_in1_10 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__82_ (
  .D({ S2501 }),
  .E({ S2515 }),
  .Q({ DP_LGU1_in1_11 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__83_ (
  .D({ S2502 }),
  .E({ S2515 }),
  .Q({ DP_LGU1_in1_12 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__84_ (
  .D({ S2503 }),
  .E({ S2515 }),
  .Q({ DP_LGU1_in1_13 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__85_ (
  .D({ S2504 }),
  .E({ S2515 }),
  .Q({ DP_LGU1_in1_14 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__86_ (
  .D({ S2505 }),
  .E({ S2515 }),
  .Q({ DP_LGU1_in1_15 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_369_ (
  .in1({ CU_selARU_AC }),
  .out1({ S2703 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_370_ (
  .in1({ dataBus[0] }),
  .out1({ S2704 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_371_ (
  .in1({ CU_selMEM_AC }),
  .out1({ S2705 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_372_ (
  .in1({ DP_IMM1_out_0 }),
  .out1({ S2706 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_373_ (
  .in1({ CU_selIMM_AC }),
  .out1({ S2707 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_374_ (
  .in1({ dataBus[1] }),
  .out1({ S2708 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_375_ (
  .in1({ DP_IMM1_out_1 }),
  .out1({ S2709 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_376_ (
  .in1({ dataBus[2] }),
  .out1({ S2710 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_377_ (
  .in1({ DP_IMM1_out_2 }),
  .out1({ S2711 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_378_ (
  .in1({ dataBus[3] }),
  .out1({ S2712 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_379_ (
  .in1({ DP_IMM1_out_3 }),
  .out1({ S2713 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_380_ (
  .in1({ dataBus[4] }),
  .out1({ S2714 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_381_ (
  .in1({ DP_IMM1_out_4 }),
  .out1({ S2715 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_382_ (
  .in1({ dataBus[5] }),
  .out1({ S2716 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_383_ (
  .in1({ DP_IMM1_out_5 }),
  .out1({ S2566 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_384_ (
  .in1({ dataBus[6] }),
  .out1({ S2567 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_385_ (
  .in1({ DP_IMM1_out_6 }),
  .out1({ S2568 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_386_ (
  .in1({ dataBus[7] }),
  .out1({ S2569 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_387_ (
  .in1({ DP_IMM1_out_7 }),
  .out1({ S2570 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_388_ (
  .in1({ dataBus[8] }),
  .out1({ S2571 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_389_ (
  .in1({ DP_IMM1_out_8 }),
  .out1({ S2572 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_390_ (
  .in1({ dataBus[9] }),
  .out1({ S2573 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_391_ (
  .in1({ DP_IMM1_out_9 }),
  .out1({ S2574 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_392_ (
  .in1({ dataBus[10] }),
  .out1({ S2575 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_393_ (
  .in1({ DP_IMM1_out_10 }),
  .out1({ S2576 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_394_ (
  .in1({ dataBus[11] }),
  .out1({ S2577 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_395_ (
  .in1({ DP_IMM1_out_11 }),
  .out1({ S2578 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_396_ (
  .in1({ dataBus[12] }),
  .out1({ S2579 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_397_ (
  .in1({ DP_IMM1_out_12 }),
  .out1({ S2580 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_398_ (
  .in1({ dataBus[13] }),
  .out1({ S2581 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_399_ (
  .in1({ DP_IMM1_out_13 }),
  .out1({ S2582 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_400_ (
  .in1({ dataBus[14] }),
  .out1({ S2583 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_401_ (
  .in1({ DP_IMM1_out_14 }),
  .out1({ S2584 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_402_ (
  .in1({ dataBus[15] }),
  .out1({ S2585 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_403_ (
  .in1({ DP_IMM1_out_15 }),
  .out1({ S2586 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_404_ (
  .in1({ CU_selLGU_AC }),
  .out1({ S2587 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1331_ (
  .in1({ S2707, S2705 }),
  .out1({ S2588 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1332_ (
  .in1({ CU_selARU_AC, DP_ARU1_out_0 }),
  .out1({ S2589 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1333_ (
  .in1({ S2703, DP_LGU1_out_0 }),
  .out1({ S2590 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1334_ (
  .in1({ S2590, S2589 }),
  .out1({ S2591 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_880_ (
  .in1({ S2591, S2588 }),
  .out1({ S2592 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1335_ (
  .in1({ CU_selIMM_AC, S2706 }),
  .out1({ S2593 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_881_ (
  .in1({ CU_selIMM_AC, S2705 }),
  .out1({ S2594 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1336_ (
  .in1({ S2594, S2704 }),
  .out1({ S2595 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1337_ (
  .in1({ S2595, S2593 }),
  .out1({ S2596 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_882_ (
  .in1({ S2596, S2592 }),
  .out1({ S2549 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1338_ (
  .in1({ DP_LGU1_out_1, S2703 }),
  .out1({ S2597 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1339_ (
  .in1({ DP_ARU1_out_1, CU_selARU_AC }),
  .out1({ S2598 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1340_ (
  .in1({ S2598, S2597 }),
  .out1({ S2599 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_883_ (
  .in1({ S2599, S2588 }),
  .out1({ S2600 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1341_ (
  .in1({ S2709, CU_selIMM_AC }),
  .out1({ S2601 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1342_ (
  .in1({ S2594, S2708 }),
  .out1({ S2602 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1343_ (
  .in1({ S2602, S2601 }),
  .out1({ S2603 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_884_ (
  .in1({ S2603, S2600 }),
  .out1({ S2556 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1344_ (
  .in1({ DP_LGU1_out_2, S2703 }),
  .out1({ S2604 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1345_ (
  .in1({ DP_ARU1_out_2, CU_selARU_AC }),
  .out1({ S2605 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1346_ (
  .in1({ S2605, S2604 }),
  .out1({ S2606 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_885_ (
  .in1({ S2606, S2588 }),
  .out1({ S2607 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1347_ (
  .in1({ S2711, CU_selIMM_AC }),
  .out1({ S2608 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1348_ (
  .in1({ S2594, S2710 }),
  .out1({ S2609 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1349_ (
  .in1({ S2609, S2608 }),
  .out1({ S2610 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_886_ (
  .in1({ S2610, S2607 }),
  .out1({ S2557 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1350_ (
  .in1({ DP_LGU1_out_3, S2703 }),
  .out1({ S2611 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1351_ (
  .in1({ DP_ARU1_out_3, CU_selARU_AC }),
  .out1({ S2612 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1352_ (
  .in1({ S2612, S2611 }),
  .out1({ S2613 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_887_ (
  .in1({ S2613, S2588 }),
  .out1({ S2614 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1353_ (
  .in1({ S2713, CU_selIMM_AC }),
  .out1({ S2615 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1354_ (
  .in1({ S2594, S2712 }),
  .out1({ S2616 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1355_ (
  .in1({ S2616, S2615 }),
  .out1({ S2617 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_888_ (
  .in1({ S2617, S2614 }),
  .out1({ S2558 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1356_ (
  .in1({ DP_LGU1_out_4, S2703 }),
  .out1({ S2618 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1357_ (
  .in1({ DP_ARU1_out_4, CU_selARU_AC }),
  .out1({ S2619 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1358_ (
  .in1({ S2619, S2618 }),
  .out1({ S2620 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_889_ (
  .in1({ S2620, S2588 }),
  .out1({ S2621 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1359_ (
  .in1({ S2715, CU_selIMM_AC }),
  .out1({ S2622 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1360_ (
  .in1({ S2594, S2714 }),
  .out1({ S2623 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1361_ (
  .in1({ S2623, S2622 }),
  .out1({ S2624 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_890_ (
  .in1({ S2624, S2621 }),
  .out1({ S2559 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1362_ (
  .in1({ DP_LGU1_out_5, S2703 }),
  .out1({ S2625 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1363_ (
  .in1({ DP_ARU1_out_5, CU_selARU_AC }),
  .out1({ S2626 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1364_ (
  .in1({ S2626, S2625 }),
  .out1({ S2627 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_891_ (
  .in1({ S2627, S2588 }),
  .out1({ S2628 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1365_ (
  .in1({ S2566, CU_selIMM_AC }),
  .out1({ S2629 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1366_ (
  .in1({ S2594, S2716 }),
  .out1({ S2630 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1367_ (
  .in1({ S2630, S2629 }),
  .out1({ S2631 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_892_ (
  .in1({ S2631, S2628 }),
  .out1({ S2560 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1368_ (
  .in1({ DP_LGU1_out_6, S2703 }),
  .out1({ S2632 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1369_ (
  .in1({ DP_ARU1_out_6, CU_selARU_AC }),
  .out1({ S2633 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1370_ (
  .in1({ S2633, S2632 }),
  .out1({ S2634 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_893_ (
  .in1({ S2634, S2588 }),
  .out1({ S2635 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1371_ (
  .in1({ S2568, CU_selIMM_AC }),
  .out1({ S2636 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1372_ (
  .in1({ S2594, S2567 }),
  .out1({ S2637 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1373_ (
  .in1({ S2637, S2636 }),
  .out1({ S2638 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_894_ (
  .in1({ S2638, S2635 }),
  .out1({ S2561 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1374_ (
  .in1({ DP_LGU1_out_7, S2703 }),
  .out1({ S2639 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1375_ (
  .in1({ DP_ARU1_out_7, CU_selARU_AC }),
  .out1({ S2640 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1376_ (
  .in1({ S2640, S2639 }),
  .out1({ S2641 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_895_ (
  .in1({ S2641, S2588 }),
  .out1({ S2642 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1377_ (
  .in1({ S2570, CU_selIMM_AC }),
  .out1({ S2643 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1378_ (
  .in1({ S2594, S2569 }),
  .out1({ S2644 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1379_ (
  .in1({ S2644, S2643 }),
  .out1({ S2645 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_896_ (
  .in1({ S2645, S2642 }),
  .out1({ S2562 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1380_ (
  .in1({ DP_ARU1_out_8, CU_selARU_AC }),
  .out1({ S2646 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1381_ (
  .in1({ DP_LGU1_out_8, S2703 }),
  .out1({ S2647 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1382_ (
  .in1({ S2647, S2646 }),
  .out1({ S2648 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_897_ (
  .in1({ S2648, S2588 }),
  .out1({ S2649 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1383_ (
  .in1({ S2572, CU_selIMM_AC }),
  .out1({ S2650 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1384_ (
  .in1({ S2594, S2571 }),
  .out1({ S2651 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1385_ (
  .in1({ S2651, S2650 }),
  .out1({ S2652 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_898_ (
  .in1({ S2652, S2649 }),
  .out1({ S2563 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1386_ (
  .in1({ DP_LGU1_out_9, S2703 }),
  .out1({ S2653 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1387_ (
  .in1({ DP_ARU1_out_9, CU_selARU_AC }),
  .out1({ S2654 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1388_ (
  .in1({ S2654, S2653 }),
  .out1({ S2655 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_899_ (
  .in1({ S2655, S2588 }),
  .out1({ S2656 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1389_ (
  .in1({ S2574, CU_selIMM_AC }),
  .out1({ S2657 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1390_ (
  .in1({ S2594, S2573 }),
  .out1({ S2658 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1391_ (
  .in1({ S2658, S2657 }),
  .out1({ S2659 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_900_ (
  .in1({ S2659, S2656 }),
  .out1({ S2564 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1392_ (
  .in1({ DP_ARU1_out_10, CU_selARU_AC }),
  .out1({ S2660 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1393_ (
  .in1({ DP_LGU1_out_10, S2703 }),
  .out1({ S2661 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1394_ (
  .in1({ S2661, S2660 }),
  .out1({ S2662 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_901_ (
  .in1({ S2662, S2588 }),
  .out1({ S2663 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1395_ (
  .in1({ S2576, CU_selIMM_AC }),
  .out1({ S2664 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1396_ (
  .in1({ S2594, S2575 }),
  .out1({ S2665 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1397_ (
  .in1({ S2665, S2664 }),
  .out1({ S2666 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_902_ (
  .in1({ S2666, S2663 }),
  .out1({ S2550 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1398_ (
  .in1({ DP_LGU1_out_11, S2703 }),
  .out1({ S2667 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1399_ (
  .in1({ DP_ARU1_out_11, CU_selARU_AC }),
  .out1({ S2668 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1400_ (
  .in1({ S2668, S2667 }),
  .out1({ S2669 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_903_ (
  .in1({ S2669, S2588 }),
  .out1({ S2670 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1401_ (
  .in1({ S2578, CU_selIMM_AC }),
  .out1({ S2671 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1402_ (
  .in1({ S2594, S2577 }),
  .out1({ S2672 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1403_ (
  .in1({ S2672, S2671 }),
  .out1({ S2673 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_904_ (
  .in1({ S2673, S2670 }),
  .out1({ S2551 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1404_ (
  .in1({ DP_ARU1_out_12, CU_selARU_AC }),
  .out1({ S2674 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1405_ (
  .in1({ DP_LGU1_out_12, S2703 }),
  .out1({ S2675 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1406_ (
  .in1({ S2675, S2674 }),
  .out1({ S2676 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_905_ (
  .in1({ S2676, S2588 }),
  .out1({ S2677 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1407_ (
  .in1({ S2580, CU_selIMM_AC }),
  .out1({ S2678 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1408_ (
  .in1({ S2594, S2579 }),
  .out1({ S2679 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1409_ (
  .in1({ S2679, S2678 }),
  .out1({ S2680 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_906_ (
  .in1({ S2680, S2677 }),
  .out1({ S2552 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1410_ (
  .in1({ DP_LGU1_out_13, S2703 }),
  .out1({ S2681 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1411_ (
  .in1({ DP_ARU1_out_13, CU_selARU_AC }),
  .out1({ S2682 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1412_ (
  .in1({ S2682, S2681 }),
  .out1({ S2683 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_907_ (
  .in1({ S2683, S2588 }),
  .out1({ S2684 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1413_ (
  .in1({ S2582, CU_selIMM_AC }),
  .out1({ S2685 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1414_ (
  .in1({ S2594, S2581 }),
  .out1({ S2686 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1415_ (
  .in1({ S2686, S2685 }),
  .out1({ S2687 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_908_ (
  .in1({ S2687, S2684 }),
  .out1({ S2553 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1416_ (
  .in1({ DP_ARU1_out_14, CU_selARU_AC }),
  .out1({ S2688 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1417_ (
  .in1({ DP_LGU1_out_14, S2703 }),
  .out1({ S2689 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1418_ (
  .in1({ S2689, S2688 }),
  .out1({ S2690 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_909_ (
  .in1({ S2690, S2588 }),
  .out1({ S2691 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1419_ (
  .in1({ S2584, CU_selIMM_AC }),
  .out1({ S2692 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1420_ (
  .in1({ S2594, S2583 }),
  .out1({ S2693 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1421_ (
  .in1({ S2693, S2692 }),
  .out1({ S2694 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_910_ (
  .in1({ S2694, S2691 }),
  .out1({ S2554 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1422_ (
  .in1({ DP_LGU1_N, S2703 }),
  .out1({ S2695 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1423_ (
  .in1({ DP_ARU1_N, CU_selARU_AC }),
  .out1({ S2696 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1424_ (
  .in1({ S2696, S2695 }),
  .out1({ S2697 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_911_ (
  .in1({ S2697, S2588 }),
  .out1({ S2698 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1425_ (
  .in1({ S2586, CU_selIMM_AC }),
  .out1({ S2699 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1426_ (
  .in1({ S2594, S2585 }),
  .out1({ S2700 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1427_ (
  .in1({ S2700, S2699 }),
  .out1({ S2701 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_912_ (
  .in1({ S2701, S2698 }),
  .out1({ S2555 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1428_ (
  .in1({ S2587, S2703 }),
  .out1({ S2702 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_913_ (
  .in1({ S2702, S2588 }),
  .out1({ S2565 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__87_ (
  .D({ S2549 }),
  .E({ S2565 }),
  .Q({ DP_AC_in_0 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__88_ (
  .D({ S2556 }),
  .E({ S2565 }),
  .Q({ DP_AC_in_1 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__89_ (
  .D({ S2557 }),
  .E({ S2565 }),
  .Q({ DP_AC_in_2 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__90_ (
  .D({ S2558 }),
  .E({ S2565 }),
  .Q({ DP_AC_in_3 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__91_ (
  .D({ S2559 }),
  .E({ S2565 }),
  .Q({ DP_AC_in_4 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__92_ (
  .D({ S2560 }),
  .E({ S2565 }),
  .Q({ DP_AC_in_5 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__93_ (
  .D({ S2561 }),
  .E({ S2565 }),
  .Q({ DP_AC_in_6 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__94_ (
  .D({ S2562 }),
  .E({ S2565 }),
  .Q({ DP_AC_in_7 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__95_ (
  .D({ S2563 }),
  .E({ S2565 }),
  .Q({ DP_AC_in_8 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__96_ (
  .D({ S2564 }),
  .E({ S2565 }),
  .Q({ DP_AC_in_9 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__97_ (
  .D({ S2550 }),
  .E({ S2565 }),
  .Q({ DP_AC_in_10 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__98_ (
  .D({ S2551 }),
  .E({ S2565 }),
  .Q({ DP_AC_in_11 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__99_ (
  .D({ S2552 }),
  .E({ S2565 }),
  .Q({ DP_AC_in_12 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__100_ (
  .D({ S2553 }),
  .E({ S2565 }),
  .Q({ DP_AC_in_13 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__101_ (
  .D({ S2554 }),
  .E({ S2565 }),
  .Q({ DP_AC_in_14 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__102_ (
  .D({ S2555 }),
  .E({ S2565 }),
  .Q({ DP_AC_in_15 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_405_ (
  .in1({ CU_selPC_OF }),
  .out1({ S2722 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1429_ (
  .in1({ CU_selPC_OF, DP_INC_1_in_12 }),
  .out1({ S2723 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1430_ (
  .in1({ S2722, DP_IMM1_out_0 }),
  .out1({ S2724 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1431_ (
  .in1({ S2724, S2723 }),
  .out1({ S2717 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1432_ (
  .in1({ DP_INC_1_in_13, CU_selPC_OF }),
  .out1({ S2725 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1433_ (
  .in1({ DP_IMM1_out_1, S2722 }),
  .out1({ S2726 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1434_ (
  .in1({ S2726, S2725 }),
  .out1({ S2718 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1435_ (
  .in1({ DP_INC_1_in_14, CU_selPC_OF }),
  .out1({ S2727 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1436_ (
  .in1({ DP_IMM1_out_2, S2722 }),
  .out1({ S2728 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1437_ (
  .in1({ S2728, S2727 }),
  .out1({ S2719 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1438_ (
  .in1({ DP_INC_1_in_15, CU_selPC_OF }),
  .out1({ S2729 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1439_ (
  .in1({ DP_IMM1_out_3, S2722 }),
  .out1({ S2730 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1440_ (
  .in1({ S2730, S2729 }),
  .out1({ S2720 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_914_ (
  .in1({ CU_selIMM_OF, CU_selPC_OF }),
  .out1({ S2721 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__103_ (
  .D({ S2717 }),
  .E({ S2721 }),
  .Q({ DP_OF_in_0 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__104_ (
  .D({ S2718 }),
  .E({ S2721 }),
  .Q({ DP_OF_in_1 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__105_ (
  .D({ S2719 }),
  .E({ S2721 }),
  .Q({ DP_OF_in_2 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__106_ (
  .D({ S2720 }),
  .E({ S2721 }),
  .Q({ DP_OF_in_3 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_406_ (
  .in1({ CU_selIMM_PC }),
  .out1({ S2885 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_407_ (
  .in1({ dataBus[0] }),
  .out1({ S2886 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_408_ (
  .in1({ CU_selMEM_PC }),
  .out1({ S2887 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_409_ (
  .in1({ DP_INC_1_out_0 }),
  .out1({ S2888 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_410_ (
  .in1({ CU_selINC_PC }),
  .out1({ S2889 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_411_ (
  .in1({ dataBus[1] }),
  .out1({ S2890 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_412_ (
  .in1({ DP_INC_1_out_1 }),
  .out1({ S2891 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_413_ (
  .in1({ dataBus[2] }),
  .out1({ S2892 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_414_ (
  .in1({ DP_INC_1_out_2 }),
  .out1({ S2893 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_415_ (
  .in1({ dataBus[3] }),
  .out1({ S2894 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_416_ (
  .in1({ DP_INC_1_out_3 }),
  .out1({ S2895 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_417_ (
  .in1({ dataBus[4] }),
  .out1({ S2896 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_418_ (
  .in1({ DP_INC_1_out_4 }),
  .out1({ S2897 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_419_ (
  .in1({ dataBus[5] }),
  .out1({ S2898 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_420_ (
  .in1({ DP_INC_1_out_5 }),
  .out1({ S2748 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_421_ (
  .in1({ dataBus[6] }),
  .out1({ S2749 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_422_ (
  .in1({ DP_INC_1_out_6 }),
  .out1({ S2750 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_423_ (
  .in1({ dataBus[7] }),
  .out1({ S2751 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_424_ (
  .in1({ DP_INC_1_out_7 }),
  .out1({ S2752 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_425_ (
  .in1({ dataBus[8] }),
  .out1({ S2753 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_426_ (
  .in1({ DP_INC_1_out_8 }),
  .out1({ S2754 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_427_ (
  .in1({ dataBus[9] }),
  .out1({ S2755 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_428_ (
  .in1({ DP_INC_1_out_9 }),
  .out1({ S2756 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_429_ (
  .in1({ dataBus[10] }),
  .out1({ S2757 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_430_ (
  .in1({ DP_INC_1_out_10 }),
  .out1({ S2758 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_431_ (
  .in1({ dataBus[11] }),
  .out1({ S2759 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_432_ (
  .in1({ DP_INC_1_out_11 }),
  .out1({ S2760 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_433_ (
  .in1({ dataBus[12] }),
  .out1({ S2761 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_434_ (
  .in1({ DP_INC_1_out_12 }),
  .out1({ S2762 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_435_ (
  .in1({ dataBus[13] }),
  .out1({ S2763 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_436_ (
  .in1({ DP_INC_1_out_13 }),
  .out1({ S2764 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_437_ (
  .in1({ dataBus[14] }),
  .out1({ S2765 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_438_ (
  .in1({ DP_INC_1_out_14 }),
  .out1({ S2766 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_439_ (
  .in1({ dataBus[15] }),
  .out1({ S2767 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_440_ (
  .in1({ DP_INC_1_out_15 }),
  .out1({ S2768 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_441_ (
  .in1({ 1'bz }),
  .out1({ S2769 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1441_ (
  .in1({ S2889, S2887 }),
  .out1({ S2770 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1442_ (
  .in1({ CU_selIMM_PC, DP_IMM1_out_0 }),
  .out1({ S2771 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1443_ (
  .in1({ S2885, 1'bz }),
  .out1({ S2772 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1444_ (
  .in1({ S2772, S2771 }),
  .out1({ S2773 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_915_ (
  .in1({ S2773, S2770 }),
  .out1({ S2774 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1445_ (
  .in1({ CU_selINC_PC, S2888 }),
  .out1({ S2775 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_916_ (
  .in1({ CU_selINC_PC, S2887 }),
  .out1({ S2776 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1446_ (
  .in1({ S2776, S2886 }),
  .out1({ S2777 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1447_ (
  .in1({ S2777, S2775 }),
  .out1({ S2778 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_917_ (
  .in1({ S2778, S2774 }),
  .out1({ S2731 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1448_ (
  .in1({ 1'bz, S2885 }),
  .out1({ S2779 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1449_ (
  .in1({ DP_IMM1_out_1, CU_selIMM_PC }),
  .out1({ S2780 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1450_ (
  .in1({ S2780, S2779 }),
  .out1({ S2781 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_918_ (
  .in1({ S2781, S2770 }),
  .out1({ S2782 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1451_ (
  .in1({ S2891, CU_selINC_PC }),
  .out1({ S2783 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1452_ (
  .in1({ S2776, S2890 }),
  .out1({ S2784 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1453_ (
  .in1({ S2784, S2783 }),
  .out1({ S2785 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_919_ (
  .in1({ S2785, S2782 }),
  .out1({ S2738 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1454_ (
  .in1({ 1'bz, S2885 }),
  .out1({ S2786 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1455_ (
  .in1({ DP_IMM1_out_2, CU_selIMM_PC }),
  .out1({ S2787 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1456_ (
  .in1({ S2787, S2786 }),
  .out1({ S2788 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_920_ (
  .in1({ S2788, S2770 }),
  .out1({ S2789 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1457_ (
  .in1({ S2893, CU_selINC_PC }),
  .out1({ S2790 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1458_ (
  .in1({ S2776, S2892 }),
  .out1({ S2791 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1459_ (
  .in1({ S2791, S2790 }),
  .out1({ S2792 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_921_ (
  .in1({ S2792, S2789 }),
  .out1({ S2739 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1460_ (
  .in1({ 1'bz, S2885 }),
  .out1({ S2793 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1461_ (
  .in1({ DP_IMM1_out_3, CU_selIMM_PC }),
  .out1({ S2794 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1462_ (
  .in1({ S2794, S2793 }),
  .out1({ S2795 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_922_ (
  .in1({ S2795, S2770 }),
  .out1({ S2796 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1463_ (
  .in1({ S2895, CU_selINC_PC }),
  .out1({ S2797 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1464_ (
  .in1({ S2776, S2894 }),
  .out1({ S2798 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1465_ (
  .in1({ S2798, S2797 }),
  .out1({ S2799 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_923_ (
  .in1({ S2799, S2796 }),
  .out1({ S2740 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1466_ (
  .in1({ 1'bz, S2885 }),
  .out1({ S2800 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1467_ (
  .in1({ DP_IMM1_out_4, CU_selIMM_PC }),
  .out1({ S2801 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1468_ (
  .in1({ S2801, S2800 }),
  .out1({ S2802 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_924_ (
  .in1({ S2802, S2770 }),
  .out1({ S2803 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1469_ (
  .in1({ S2897, CU_selINC_PC }),
  .out1({ S2804 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1470_ (
  .in1({ S2776, S2896 }),
  .out1({ S2805 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1471_ (
  .in1({ S2805, S2804 }),
  .out1({ S2806 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_925_ (
  .in1({ S2806, S2803 }),
  .out1({ S2741 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1472_ (
  .in1({ 1'bz, S2885 }),
  .out1({ S2807 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1473_ (
  .in1({ DP_IMM1_out_5, CU_selIMM_PC }),
  .out1({ S2808 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1474_ (
  .in1({ S2808, S2807 }),
  .out1({ S2809 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_926_ (
  .in1({ S2809, S2770 }),
  .out1({ S2810 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1475_ (
  .in1({ S2748, CU_selINC_PC }),
  .out1({ S2811 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1476_ (
  .in1({ S2776, S2898 }),
  .out1({ S2812 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1477_ (
  .in1({ S2812, S2811 }),
  .out1({ S2813 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_927_ (
  .in1({ S2813, S2810 }),
  .out1({ S2742 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1478_ (
  .in1({ 1'bz, S2885 }),
  .out1({ S2814 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1479_ (
  .in1({ DP_IMM1_out_6, CU_selIMM_PC }),
  .out1({ S2815 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1480_ (
  .in1({ S2815, S2814 }),
  .out1({ S2816 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_928_ (
  .in1({ S2816, S2770 }),
  .out1({ S2817 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1481_ (
  .in1({ S2750, CU_selINC_PC }),
  .out1({ S2818 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1482_ (
  .in1({ S2776, S2749 }),
  .out1({ S2819 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1483_ (
  .in1({ S2819, S2818 }),
  .out1({ S2820 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_929_ (
  .in1({ S2820, S2817 }),
  .out1({ S2743 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1484_ (
  .in1({ 1'bz, S2885 }),
  .out1({ S2821 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1485_ (
  .in1({ DP_IMM1_out_7, CU_selIMM_PC }),
  .out1({ S2822 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1486_ (
  .in1({ S2822, S2821 }),
  .out1({ S2823 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_930_ (
  .in1({ S2823, S2770 }),
  .out1({ S2824 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1487_ (
  .in1({ S2752, CU_selINC_PC }),
  .out1({ S2825 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1488_ (
  .in1({ S2776, S2751 }),
  .out1({ S2826 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1489_ (
  .in1({ S2826, S2825 }),
  .out1({ S2827 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_931_ (
  .in1({ S2827, S2824 }),
  .out1({ S2744 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1490_ (
  .in1({ DP_IMM1_out_8, CU_selIMM_PC }),
  .out1({ S2828 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1491_ (
  .in1({ 1'bz, S2885 }),
  .out1({ S2829 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1492_ (
  .in1({ S2829, S2828 }),
  .out1({ S2830 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_932_ (
  .in1({ S2830, S2770 }),
  .out1({ S2831 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1493_ (
  .in1({ S2754, CU_selINC_PC }),
  .out1({ S2832 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1494_ (
  .in1({ S2776, S2753 }),
  .out1({ S2833 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1495_ (
  .in1({ S2833, S2832 }),
  .out1({ S2834 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_933_ (
  .in1({ S2834, S2831 }),
  .out1({ S2745 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1496_ (
  .in1({ 1'bz, S2885 }),
  .out1({ S2835 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1497_ (
  .in1({ DP_IMM1_out_9, CU_selIMM_PC }),
  .out1({ S2836 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1498_ (
  .in1({ S2836, S2835 }),
  .out1({ S2837 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_934_ (
  .in1({ S2837, S2770 }),
  .out1({ S2838 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1499_ (
  .in1({ S2756, CU_selINC_PC }),
  .out1({ S2839 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1500_ (
  .in1({ S2776, S2755 }),
  .out1({ S2840 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1501_ (
  .in1({ S2840, S2839 }),
  .out1({ S2841 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_935_ (
  .in1({ S2841, S2838 }),
  .out1({ S2746 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1502_ (
  .in1({ DP_IMM1_out_10, CU_selIMM_PC }),
  .out1({ S2842 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1503_ (
  .in1({ 1'bz, S2885 }),
  .out1({ S2843 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1504_ (
  .in1({ S2843, S2842 }),
  .out1({ S2844 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_936_ (
  .in1({ S2844, S2770 }),
  .out1({ S2845 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1505_ (
  .in1({ S2758, CU_selINC_PC }),
  .out1({ S2846 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1506_ (
  .in1({ S2776, S2757 }),
  .out1({ S2847 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1507_ (
  .in1({ S2847, S2846 }),
  .out1({ S2848 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_937_ (
  .in1({ S2848, S2845 }),
  .out1({ S2732 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1508_ (
  .in1({ 1'bz, S2885 }),
  .out1({ S2849 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1509_ (
  .in1({ DP_IMM1_out_11, CU_selIMM_PC }),
  .out1({ S2850 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1510_ (
  .in1({ S2850, S2849 }),
  .out1({ S2851 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_938_ (
  .in1({ S2851, S2770 }),
  .out1({ S2852 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1511_ (
  .in1({ S2760, CU_selINC_PC }),
  .out1({ S2853 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1512_ (
  .in1({ S2776, S2759 }),
  .out1({ S2854 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1513_ (
  .in1({ S2854, S2853 }),
  .out1({ S2855 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_939_ (
  .in1({ S2855, S2852 }),
  .out1({ S2733 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1514_ (
  .in1({ DP_IMM1_out_12, CU_selIMM_PC }),
  .out1({ S2856 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1515_ (
  .in1({ 1'bz, S2885 }),
  .out1({ S2857 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1516_ (
  .in1({ S2857, S2856 }),
  .out1({ S2858 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_940_ (
  .in1({ S2858, S2770 }),
  .out1({ S2859 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1517_ (
  .in1({ S2762, CU_selINC_PC }),
  .out1({ S2860 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1518_ (
  .in1({ S2776, S2761 }),
  .out1({ S2861 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1519_ (
  .in1({ S2861, S2860 }),
  .out1({ S2862 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_941_ (
  .in1({ S2862, S2859 }),
  .out1({ S2734 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1520_ (
  .in1({ 1'bz, S2885 }),
  .out1({ S2863 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1521_ (
  .in1({ DP_IMM1_out_13, CU_selIMM_PC }),
  .out1({ S2864 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1522_ (
  .in1({ S2864, S2863 }),
  .out1({ S2865 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_942_ (
  .in1({ S2865, S2770 }),
  .out1({ S2866 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1523_ (
  .in1({ S2764, CU_selINC_PC }),
  .out1({ S2867 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1524_ (
  .in1({ S2776, S2763 }),
  .out1({ S2868 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1525_ (
  .in1({ S2868, S2867 }),
  .out1({ S2869 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_943_ (
  .in1({ S2869, S2866 }),
  .out1({ S2735 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1526_ (
  .in1({ DP_IMM1_out_14, CU_selIMM_PC }),
  .out1({ S2870 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1527_ (
  .in1({ 1'bz, S2885 }),
  .out1({ S2871 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1528_ (
  .in1({ S2871, S2870 }),
  .out1({ S2872 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_944_ (
  .in1({ S2872, S2770 }),
  .out1({ S2873 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1529_ (
  .in1({ S2766, CU_selINC_PC }),
  .out1({ S2874 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1530_ (
  .in1({ S2776, S2765 }),
  .out1({ S2875 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1531_ (
  .in1({ S2875, S2874 }),
  .out1({ S2876 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_945_ (
  .in1({ S2876, S2873 }),
  .out1({ S2736 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1532_ (
  .in1({ 1'bz, S2885 }),
  .out1({ S2877 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1533_ (
  .in1({ DP_IMM1_out_15, CU_selIMM_PC }),
  .out1({ S2878 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1534_ (
  .in1({ S2878, S2877 }),
  .out1({ S2879 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_946_ (
  .in1({ S2879, S2770 }),
  .out1({ S2880 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1535_ (
  .in1({ S2768, CU_selINC_PC }),
  .out1({ S2881 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1536_ (
  .in1({ S2776, S2767 }),
  .out1({ S2882 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1537_ (
  .in1({ S2882, S2881 }),
  .out1({ S2883 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_947_ (
  .in1({ S2883, S2880 }),
  .out1({ S2737 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1538_ (
  .in1({ S2769, S2885 }),
  .out1({ S2884 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_948_ (
  .in1({ S2884, S2770 }),
  .out1({ S2747 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__107_ (
  .D({ S2731 }),
  .E({ S2747 }),
  .Q({ DP_PC_in_0 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__108_ (
  .D({ S2738 }),
  .E({ S2747 }),
  .Q({ DP_PC_in_1 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__109_ (
  .D({ S2739 }),
  .E({ S2747 }),
  .Q({ DP_PC_in_2 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__110_ (
  .D({ S2740 }),
  .E({ S2747 }),
  .Q({ DP_PC_in_3 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__111_ (
  .D({ S2741 }),
  .E({ S2747 }),
  .Q({ DP_PC_in_4 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__112_ (
  .D({ S2742 }),
  .E({ S2747 }),
  .Q({ DP_PC_in_5 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__113_ (
  .D({ S2743 }),
  .E({ S2747 }),
  .Q({ DP_PC_in_6 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__114_ (
  .D({ S2744 }),
  .E({ S2747 }),
  .Q({ DP_PC_in_7 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__115_ (
  .D({ S2745 }),
  .E({ S2747 }),
  .Q({ DP_PC_in_8 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__116_ (
  .D({ S2746 }),
  .E({ S2747 }),
  .Q({ DP_PC_in_9 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__117_ (
  .D({ S2732 }),
  .E({ S2747 }),
  .Q({ DP_PC_in_10 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__118_ (
  .D({ S2733 }),
  .E({ S2747 }),
  .Q({ DP_PC_in_11 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__119_ (
  .D({ S2734 }),
  .E({ S2747 }),
  .Q({ DP_PC_in_12 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__120_ (
  .D({ S2735 }),
  .E({ S2747 }),
  .Q({ DP_PC_in_13 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__121_ (
  .D({ S2736 }),
  .E({ S2747 }),
  .Q({ DP_PC_in_14 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__122_ (
  .D({ S2737 }),
  .E({ S2747 }),
  .Q({ DP_PC_in_15 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_442_ (
  .in1({ CU_selINC_IN }),
  .out1({ S2916 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1539_ (
  .in1({ CU_selINC_IN, DP_INC2_out_0 }),
  .out1({ S2917 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1540_ (
  .in1({ S2916, dataBus[0] }),
  .out1({ S2918 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1541_ (
  .in1({ S2918, S2917 }),
  .out1({ S2899 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1542_ (
  .in1({ DP_INC2_out_1, CU_selINC_IN }),
  .out1({ S2919 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1543_ (
  .in1({ dataBus[1], S2916 }),
  .out1({ S2920 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1544_ (
  .in1({ S2920, S2919 }),
  .out1({ S2906 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1545_ (
  .in1({ DP_INC2_out_2, CU_selINC_IN }),
  .out1({ S2921 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1546_ (
  .in1({ dataBus[2], S2916 }),
  .out1({ S2922 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1547_ (
  .in1({ S2922, S2921 }),
  .out1({ S2907 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1548_ (
  .in1({ DP_INC2_out_3, CU_selINC_IN }),
  .out1({ S2923 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1549_ (
  .in1({ dataBus[3], S2916 }),
  .out1({ S2924 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1550_ (
  .in1({ S2924, S2923 }),
  .out1({ S2908 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1551_ (
  .in1({ DP_INC2_out_4, CU_selINC_IN }),
  .out1({ S2925 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1552_ (
  .in1({ dataBus[4], S2916 }),
  .out1({ S2926 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1553_ (
  .in1({ S2926, S2925 }),
  .out1({ S2909 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1554_ (
  .in1({ DP_INC2_out_5, CU_selINC_IN }),
  .out1({ S2927 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1555_ (
  .in1({ dataBus[5], S2916 }),
  .out1({ S2928 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1556_ (
  .in1({ S2928, S2927 }),
  .out1({ S2910 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1557_ (
  .in1({ DP_INC2_out_6, CU_selINC_IN }),
  .out1({ S2929 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1558_ (
  .in1({ dataBus[6], S2916 }),
  .out1({ S2930 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1559_ (
  .in1({ S2930, S2929 }),
  .out1({ S2911 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1560_ (
  .in1({ DP_INC2_out_7, CU_selINC_IN }),
  .out1({ S2931 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1561_ (
  .in1({ dataBus[7], S2916 }),
  .out1({ S2932 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1562_ (
  .in1({ S2932, S2931 }),
  .out1({ S2912 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1563_ (
  .in1({ DP_INC2_out_8, CU_selINC_IN }),
  .out1({ S2933 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1564_ (
  .in1({ dataBus[8], S2916 }),
  .out1({ S2934 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1565_ (
  .in1({ S2934, S2933 }),
  .out1({ S2913 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1566_ (
  .in1({ DP_INC2_out_9, CU_selINC_IN }),
  .out1({ S2935 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1567_ (
  .in1({ dataBus[9], S2916 }),
  .out1({ S2936 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1568_ (
  .in1({ S2936, S2935 }),
  .out1({ S2914 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1569_ (
  .in1({ DP_INC2_out_10, CU_selINC_IN }),
  .out1({ S2937 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1570_ (
  .in1({ dataBus[10], S2916 }),
  .out1({ S2938 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1571_ (
  .in1({ S2938, S2937 }),
  .out1({ S2900 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1572_ (
  .in1({ DP_INC2_out_11, CU_selINC_IN }),
  .out1({ S2939 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1573_ (
  .in1({ dataBus[11], S2916 }),
  .out1({ S2940 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1574_ (
  .in1({ S2940, S2939 }),
  .out1({ S2901 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1575_ (
  .in1({ DP_INC2_out_12, CU_selINC_IN }),
  .out1({ S2941 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1576_ (
  .in1({ dataBus[12], S2916 }),
  .out1({ S2942 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1577_ (
  .in1({ S2942, S2941 }),
  .out1({ S2902 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1578_ (
  .in1({ DP_INC2_out_13, CU_selINC_IN }),
  .out1({ S2943 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1579_ (
  .in1({ dataBus[13], S2916 }),
  .out1({ S2944 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1580_ (
  .in1({ S2944, S2943 }),
  .out1({ S2903 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1581_ (
  .in1({ DP_INC2_out_14, CU_selINC_IN }),
  .out1({ S2945 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1582_ (
  .in1({ dataBus[14], S2916 }),
  .out1({ S2946 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1583_ (
  .in1({ S2946, S2945 }),
  .out1({ S2904 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1584_ (
  .in1({ DP_INC2_out_15, CU_selINC_IN }),
  .out1({ S2947 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1585_ (
  .in1({ dataBus[15], S2916 }),
  .out1({ S2948 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1586_ (
  .in1({ S2948, S2947 }),
  .out1({ S2905 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_949_ (
  .in1({ CU_selMEM_IN, CU_selINC_IN }),
  .out1({ S2915 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__123_ (
  .D({ S2899 }),
  .E({ S2915 }),
  .Q({ DP_IN_in_0 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__124_ (
  .D({ S2906 }),
  .E({ S2915 }),
  .Q({ DP_IN_in_1 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__125_ (
  .D({ S2907 }),
  .E({ S2915 }),
  .Q({ DP_IN_in_2 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__126_ (
  .D({ S2908 }),
  .E({ S2915 }),
  .Q({ DP_IN_in_3 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__127_ (
  .D({ S2909 }),
  .E({ S2915 }),
  .Q({ DP_IN_in_4 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__128_ (
  .D({ S2910 }),
  .E({ S2915 }),
  .Q({ DP_IN_in_5 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__129_ (
  .D({ S2911 }),
  .E({ S2915 }),
  .Q({ DP_IN_in_6 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__130_ (
  .D({ S2912 }),
  .E({ S2915 }),
  .Q({ DP_IN_in_7 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__131_ (
  .D({ S2913 }),
  .E({ S2915 }),
  .Q({ DP_IN_in_8 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__132_ (
  .D({ S2914 }),
  .E({ S2915 }),
  .Q({ DP_IN_in_9 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__133_ (
  .D({ S2900 }),
  .E({ S2915 }),
  .Q({ DP_IN_in_10 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__134_ (
  .D({ S2901 }),
  .E({ S2915 }),
  .Q({ DP_IN_in_11 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__135_ (
  .D({ S2902 }),
  .E({ S2915 }),
  .Q({ DP_IN_in_12 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__136_ (
  .D({ S2903 }),
  .E({ S2915 }),
  .Q({ DP_IN_in_13 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__137_ (
  .D({ S2904 }),
  .E({ S2915 }),
  .Q({ DP_IN_in_14 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__138_ (
  .D({ S2905 }),
  .E({ S2915 }),
  .Q({ DP_IN_in_15 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_443_ (
  .in1({ CU_selAC_MEM }),
  .out1({ S3103 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_444_ (
  .in1({ DP_INC_1_out_0 }),
  .out1({ S3104 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_445_ (
  .in1({ CU_selPC_MEM }),
  .out1({ S3105 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_446_ (
  .in1({ DP_IN_out_0 }),
  .out1({ S3106 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_447_ (
  .in1({ CU_selIN_MEM }),
  .out1({ S3107 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_448_ (
  .in1({ DP_INC_1_out_1 }),
  .out1({ S3108 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_449_ (
  .in1({ DP_IN_out_1 }),
  .out1({ S3109 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_450_ (
  .in1({ DP_INC_1_out_2 }),
  .out1({ S3110 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_451_ (
  .in1({ DP_IN_out_2 }),
  .out1({ S3111 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_452_ (
  .in1({ DP_INC_1_out_3 }),
  .out1({ S3112 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_453_ (
  .in1({ DP_IN_out_3 }),
  .out1({ S3113 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_454_ (
  .in1({ DP_INC_1_out_4 }),
  .out1({ S3114 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_455_ (
  .in1({ DP_IN_out_4 }),
  .out1({ S3115 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_456_ (
  .in1({ DP_INC_1_out_5 }),
  .out1({ S3116 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_457_ (
  .in1({ DP_IN_out_5 }),
  .out1({ S2966 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_458_ (
  .in1({ DP_INC_1_out_6 }),
  .out1({ S2967 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_459_ (
  .in1({ DP_IN_out_6 }),
  .out1({ S2968 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_460_ (
  .in1({ DP_INC_1_out_7 }),
  .out1({ S2969 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_461_ (
  .in1({ DP_IN_out_7 }),
  .out1({ S2970 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_462_ (
  .in1({ DP_INC_1_out_8 }),
  .out1({ S2971 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_463_ (
  .in1({ DP_IN_out_8 }),
  .out1({ S2972 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_464_ (
  .in1({ DP_INC_1_out_9 }),
  .out1({ S2973 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_465_ (
  .in1({ DP_IN_out_9 }),
  .out1({ S2974 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_466_ (
  .in1({ DP_INC_1_out_10 }),
  .out1({ S2975 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_467_ (
  .in1({ DP_IN_out_10 }),
  .out1({ S2976 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_468_ (
  .in1({ DP_INC_1_out_11 }),
  .out1({ S2977 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_469_ (
  .in1({ DP_IN_out_11 }),
  .out1({ S2978 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_470_ (
  .in1({ DP_INC_1_out_12 }),
  .out1({ S2979 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_471_ (
  .in1({ DP_IN_out_12 }),
  .out1({ S2980 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_472_ (
  .in1({ DP_INC_1_out_13 }),
  .out1({ S2981 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_473_ (
  .in1({ DP_IN_out_13 }),
  .out1({ S2982 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_474_ (
  .in1({ DP_INC_1_out_14 }),
  .out1({ S2983 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_475_ (
  .in1({ DP_IN_out_14 }),
  .out1({ S2984 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_476_ (
  .in1({ DP_INC_1_out_15 }),
  .out1({ S2985 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_477_ (
  .in1({ DP_IN_out_15 }),
  .out1({ S2986 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_478_ (
  .in1({ 1'bz }),
  .out1({ S2987 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1587_ (
  .in1({ S3107, S3105 }),
  .out1({ S2988 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1588_ (
  .in1({ CU_selAC_MEM, DP_AC_out_0 }),
  .out1({ S2989 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1589_ (
  .in1({ S3103, 1'bz }),
  .out1({ S2990 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1590_ (
  .in1({ S2990, S2989 }),
  .out1({ S2991 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_950_ (
  .in1({ S2991, S2988 }),
  .out1({ S2992 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1591_ (
  .in1({ CU_selIN_MEM, S3106 }),
  .out1({ S2993 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_951_ (
  .in1({ CU_selIN_MEM, S3105 }),
  .out1({ S2994 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1592_ (
  .in1({ S2994, S3104 }),
  .out1({ S2995 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1593_ (
  .in1({ S2995, S2993 }),
  .out1({ S2996 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_952_ (
  .in1({ S2996, S2992 }),
  .out1({ S2949 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1594_ (
  .in1({ 1'bz, S3103 }),
  .out1({ S2997 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1595_ (
  .in1({ DP_AC_out_1, CU_selAC_MEM }),
  .out1({ S2998 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1596_ (
  .in1({ S2998, S2997 }),
  .out1({ S2999 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_953_ (
  .in1({ S2999, S2988 }),
  .out1({ S3000 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1597_ (
  .in1({ S3109, CU_selIN_MEM }),
  .out1({ S3001 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1598_ (
  .in1({ S2994, S3108 }),
  .out1({ S3002 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1599_ (
  .in1({ S3002, S3001 }),
  .out1({ S3003 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_954_ (
  .in1({ S3003, S3000 }),
  .out1({ S2956 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1600_ (
  .in1({ 1'bz, S3103 }),
  .out1({ S3004 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1601_ (
  .in1({ DP_AC_out_2, CU_selAC_MEM }),
  .out1({ S3005 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1602_ (
  .in1({ S3005, S3004 }),
  .out1({ S3006 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_955_ (
  .in1({ S3006, S2988 }),
  .out1({ S3007 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1603_ (
  .in1({ S3111, CU_selIN_MEM }),
  .out1({ S3008 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1604_ (
  .in1({ S2994, S3110 }),
  .out1({ S3009 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1605_ (
  .in1({ S3009, S3008 }),
  .out1({ S3010 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_956_ (
  .in1({ S3010, S3007 }),
  .out1({ S2957 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1606_ (
  .in1({ 1'bz, S3103 }),
  .out1({ S3011 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1607_ (
  .in1({ DP_AC_out_3, CU_selAC_MEM }),
  .out1({ S3012 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1608_ (
  .in1({ S3012, S3011 }),
  .out1({ S3013 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_957_ (
  .in1({ S3013, S2988 }),
  .out1({ S3014 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1609_ (
  .in1({ S3113, CU_selIN_MEM }),
  .out1({ S3015 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1610_ (
  .in1({ S2994, S3112 }),
  .out1({ S3016 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1611_ (
  .in1({ S3016, S3015 }),
  .out1({ S3017 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_958_ (
  .in1({ S3017, S3014 }),
  .out1({ S2958 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1612_ (
  .in1({ 1'bz, S3103 }),
  .out1({ S3018 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1613_ (
  .in1({ DP_AC_out_4, CU_selAC_MEM }),
  .out1({ S3019 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1614_ (
  .in1({ S3019, S3018 }),
  .out1({ S3020 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_959_ (
  .in1({ S3020, S2988 }),
  .out1({ S3021 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1615_ (
  .in1({ S3115, CU_selIN_MEM }),
  .out1({ S3022 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1616_ (
  .in1({ S2994, S3114 }),
  .out1({ S3023 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1617_ (
  .in1({ S3023, S3022 }),
  .out1({ S3024 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_960_ (
  .in1({ S3024, S3021 }),
  .out1({ S2959 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1618_ (
  .in1({ 1'bz, S3103 }),
  .out1({ S3025 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1619_ (
  .in1({ DP_AC_out_5, CU_selAC_MEM }),
  .out1({ S3026 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1620_ (
  .in1({ S3026, S3025 }),
  .out1({ S3027 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_961_ (
  .in1({ S3027, S2988 }),
  .out1({ S3028 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1621_ (
  .in1({ S2966, CU_selIN_MEM }),
  .out1({ S3029 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1622_ (
  .in1({ S2994, S3116 }),
  .out1({ S3030 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1623_ (
  .in1({ S3030, S3029 }),
  .out1({ S3031 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_962_ (
  .in1({ S3031, S3028 }),
  .out1({ S2960 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1624_ (
  .in1({ 1'bz, S3103 }),
  .out1({ S3032 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1625_ (
  .in1({ DP_AC_out_6, CU_selAC_MEM }),
  .out1({ S3033 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1626_ (
  .in1({ S3033, S3032 }),
  .out1({ S3034 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_963_ (
  .in1({ S3034, S2988 }),
  .out1({ S3035 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1627_ (
  .in1({ S2968, CU_selIN_MEM }),
  .out1({ S3036 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1628_ (
  .in1({ S2994, S2967 }),
  .out1({ S3037 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1629_ (
  .in1({ S3037, S3036 }),
  .out1({ S3038 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_964_ (
  .in1({ S3038, S3035 }),
  .out1({ S2961 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1630_ (
  .in1({ 1'bz, S3103 }),
  .out1({ S3039 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1631_ (
  .in1({ DP_AC_out_7, CU_selAC_MEM }),
  .out1({ S3040 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1632_ (
  .in1({ S3040, S3039 }),
  .out1({ S3041 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_965_ (
  .in1({ S3041, S2988 }),
  .out1({ S3042 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1633_ (
  .in1({ S2970, CU_selIN_MEM }),
  .out1({ S3043 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1634_ (
  .in1({ S2994, S2969 }),
  .out1({ S3044 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1635_ (
  .in1({ S3044, S3043 }),
  .out1({ S3045 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_966_ (
  .in1({ S3045, S3042 }),
  .out1({ S2962 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1636_ (
  .in1({ DP_AC_out_8, CU_selAC_MEM }),
  .out1({ S3046 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1637_ (
  .in1({ 1'bz, S3103 }),
  .out1({ S3047 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1638_ (
  .in1({ S3047, S3046 }),
  .out1({ S3048 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_967_ (
  .in1({ S3048, S2988 }),
  .out1({ S3049 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1639_ (
  .in1({ S2972, CU_selIN_MEM }),
  .out1({ S3050 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1640_ (
  .in1({ S2994, S2971 }),
  .out1({ S3051 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1641_ (
  .in1({ S3051, S3050 }),
  .out1({ S3052 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_968_ (
  .in1({ S3052, S3049 }),
  .out1({ S2963 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1642_ (
  .in1({ 1'bz, S3103 }),
  .out1({ S3053 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1643_ (
  .in1({ DP_AC_out_9, CU_selAC_MEM }),
  .out1({ S3054 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1644_ (
  .in1({ S3054, S3053 }),
  .out1({ S3055 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_969_ (
  .in1({ S3055, S2988 }),
  .out1({ S3056 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1645_ (
  .in1({ S2974, CU_selIN_MEM }),
  .out1({ S3057 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1646_ (
  .in1({ S2994, S2973 }),
  .out1({ S3058 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1647_ (
  .in1({ S3058, S3057 }),
  .out1({ S3059 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_970_ (
  .in1({ S3059, S3056 }),
  .out1({ S2964 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1648_ (
  .in1({ DP_AC_out_10, CU_selAC_MEM }),
  .out1({ S3060 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1649_ (
  .in1({ 1'bz, S3103 }),
  .out1({ S3061 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1650_ (
  .in1({ S3061, S3060 }),
  .out1({ S3062 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_971_ (
  .in1({ S3062, S2988 }),
  .out1({ S3063 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1651_ (
  .in1({ S2976, CU_selIN_MEM }),
  .out1({ S3064 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1652_ (
  .in1({ S2994, S2975 }),
  .out1({ S3065 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1653_ (
  .in1({ S3065, S3064 }),
  .out1({ S3066 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_972_ (
  .in1({ S3066, S3063 }),
  .out1({ S2950 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1654_ (
  .in1({ 1'bz, S3103 }),
  .out1({ S3067 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1655_ (
  .in1({ DP_AC_out_11, CU_selAC_MEM }),
  .out1({ S3068 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1656_ (
  .in1({ S3068, S3067 }),
  .out1({ S3069 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_973_ (
  .in1({ S3069, S2988 }),
  .out1({ S3070 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1657_ (
  .in1({ S2978, CU_selIN_MEM }),
  .out1({ S3071 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1658_ (
  .in1({ S2994, S2977 }),
  .out1({ S3072 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1659_ (
  .in1({ S3072, S3071 }),
  .out1({ S3073 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_974_ (
  .in1({ S3073, S3070 }),
  .out1({ S2951 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1660_ (
  .in1({ DP_AC_out_12, CU_selAC_MEM }),
  .out1({ S3074 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1661_ (
  .in1({ 1'bz, S3103 }),
  .out1({ S3075 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1662_ (
  .in1({ S3075, S3074 }),
  .out1({ S3076 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_975_ (
  .in1({ S3076, S2988 }),
  .out1({ S3077 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1663_ (
  .in1({ S2980, CU_selIN_MEM }),
  .out1({ S3078 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1664_ (
  .in1({ S2994, S2979 }),
  .out1({ S3079 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1665_ (
  .in1({ S3079, S3078 }),
  .out1({ S3080 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_976_ (
  .in1({ S3080, S3077 }),
  .out1({ S2952 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1666_ (
  .in1({ 1'bz, S3103 }),
  .out1({ S3081 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1667_ (
  .in1({ DP_AC_out_13, CU_selAC_MEM }),
  .out1({ S3082 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1668_ (
  .in1({ S3082, S3081 }),
  .out1({ S3083 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_977_ (
  .in1({ S3083, S2988 }),
  .out1({ S3084 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1669_ (
  .in1({ S2982, CU_selIN_MEM }),
  .out1({ S3085 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1670_ (
  .in1({ S2994, S2981 }),
  .out1({ S3086 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1671_ (
  .in1({ S3086, S3085 }),
  .out1({ S3087 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_978_ (
  .in1({ S3087, S3084 }),
  .out1({ S2953 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1672_ (
  .in1({ DP_AC_out_14, CU_selAC_MEM }),
  .out1({ S3088 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1673_ (
  .in1({ 1'bz, S3103 }),
  .out1({ S3089 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1674_ (
  .in1({ S3089, S3088 }),
  .out1({ S3090 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_979_ (
  .in1({ S3090, S2988 }),
  .out1({ S3091 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1675_ (
  .in1({ S2984, CU_selIN_MEM }),
  .out1({ S3092 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1676_ (
  .in1({ S2994, S2983 }),
  .out1({ S3093 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1677_ (
  .in1({ S3093, S3092 }),
  .out1({ S3094 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_980_ (
  .in1({ S3094, S3091 }),
  .out1({ S2954 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1678_ (
  .in1({ 1'bz, S3103 }),
  .out1({ S3095 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1679_ (
  .in1({ DP_AC_out_15, CU_selAC_MEM }),
  .out1({ S3096 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1680_ (
  .in1({ S3096, S3095 }),
  .out1({ S3097 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_981_ (
  .in1({ S3097, S2988 }),
  .out1({ S3098 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1681_ (
  .in1({ S2986, CU_selIN_MEM }),
  .out1({ S3099 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1682_ (
  .in1({ S2994, S2985 }),
  .out1({ S3100 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1683_ (
  .in1({ S3100, S3099 }),
  .out1({ S3101 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_982_ (
  .in1({ S3101, S3098 }),
  .out1({ S2955 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1684_ (
  .in1({ S2987, S3103 }),
  .out1({ S3102 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_983_ (
  .in1({ S3102, S2988 }),
  .out1({ S2965 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__139_ (
  .D({ S2949 }),
  .E({ S2965 }),
  .Q({ dataBus[0] })
);
$_DLATCH_N_ #() 
$_DLATCH_N__140_ (
  .D({ S2956 }),
  .E({ S2965 }),
  .Q({ dataBus[1] })
);
$_DLATCH_N_ #() 
$_DLATCH_N__141_ (
  .D({ S2957 }),
  .E({ S2965 }),
  .Q({ dataBus[2] })
);
$_DLATCH_N_ #() 
$_DLATCH_N__142_ (
  .D({ S2958 }),
  .E({ S2965 }),
  .Q({ dataBus[3] })
);
$_DLATCH_N_ #() 
$_DLATCH_N__143_ (
  .D({ S2959 }),
  .E({ S2965 }),
  .Q({ dataBus[4] })
);
$_DLATCH_N_ #() 
$_DLATCH_N__144_ (
  .D({ S2960 }),
  .E({ S2965 }),
  .Q({ dataBus[5] })
);
$_DLATCH_N_ #() 
$_DLATCH_N__145_ (
  .D({ S2961 }),
  .E({ S2965 }),
  .Q({ dataBus[6] })
);
$_DLATCH_N_ #() 
$_DLATCH_N__146_ (
  .D({ S2962 }),
  .E({ S2965 }),
  .Q({ dataBus[7] })
);
$_DLATCH_N_ #() 
$_DLATCH_N__147_ (
  .D({ S2963 }),
  .E({ S2965 }),
  .Q({ dataBus[8] })
);
$_DLATCH_N_ #() 
$_DLATCH_N__148_ (
  .D({ S2964 }),
  .E({ S2965 }),
  .Q({ dataBus[9] })
);
$_DLATCH_N_ #() 
$_DLATCH_N__149_ (
  .D({ S2950 }),
  .E({ S2965 }),
  .Q({ dataBus[10] })
);
$_DLATCH_N_ #() 
$_DLATCH_N__150_ (
  .D({ S2951 }),
  .E({ S2965 }),
  .Q({ dataBus[11] })
);
$_DLATCH_N_ #() 
$_DLATCH_N__151_ (
  .D({ S2952 }),
  .E({ S2965 }),
  .Q({ dataBus[12] })
);
$_DLATCH_N_ #() 
$_DLATCH_N__152_ (
  .D({ S2953 }),
  .E({ S2965 }),
  .Q({ dataBus[13] })
);
$_DLATCH_N_ #() 
$_DLATCH_N__153_ (
  .D({ S2954 }),
  .E({ S2965 }),
  .Q({ dataBus[14] })
);
$_DLATCH_N_ #() 
$_DLATCH_N__154_ (
  .D({ S2955 }),
  .E({ S2965 }),
  .Q({ dataBus[15] })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_479_ (
  .in1({ CU_ldIR }),
  .out1({ S3271 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_480_ (
  .in1({ DP_IMM1_out_0 }),
  .out1({ S3272 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_481_ (
  .in1({ CU_selIR_ADR }),
  .out1({ S3273 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_482_ (
  .in1({ DP_IN_out_0 }),
  .out1({ S3274 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_483_ (
  .in1({ CU_selIN_ADR }),
  .out1({ S3275 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_484_ (
  .in1({ DP_IMM1_out_1 }),
  .out1({ S3276 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_485_ (
  .in1({ DP_IN_out_1 }),
  .out1({ S3277 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_486_ (
  .in1({ DP_IMM1_out_2 }),
  .out1({ S3278 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_487_ (
  .in1({ DP_IN_out_2 }),
  .out1({ S3279 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_488_ (
  .in1({ DP_IMM1_out_3 }),
  .out1({ S3280 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_489_ (
  .in1({ DP_IN_out_3 }),
  .out1({ S3281 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_490_ (
  .in1({ DP_IMM1_out_4 }),
  .out1({ S3282 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_491_ (
  .in1({ DP_IN_out_4 }),
  .out1({ S3283 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_492_ (
  .in1({ DP_IMM1_out_5 }),
  .out1({ S3284 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_493_ (
  .in1({ DP_IN_out_5 }),
  .out1({ S3134 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_494_ (
  .in1({ DP_IMM1_out_6 }),
  .out1({ S3135 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_495_ (
  .in1({ DP_IN_out_6 }),
  .out1({ S3136 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_496_ (
  .in1({ DP_IMM1_out_7 }),
  .out1({ S3137 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_497_ (
  .in1({ DP_IN_out_7 }),
  .out1({ S3138 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_498_ (
  .in1({ DP_IMM1_out_8 }),
  .out1({ S3139 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_499_ (
  .in1({ DP_IN_out_8 }),
  .out1({ S3140 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_500_ (
  .in1({ DP_IMM1_out_9 }),
  .out1({ S3141 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_501_ (
  .in1({ DP_IN_out_9 }),
  .out1({ S3142 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_502_ (
  .in1({ DP_IMM1_out_10 }),
  .out1({ S3143 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_503_ (
  .in1({ DP_IN_out_10 }),
  .out1({ S3144 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_504_ (
  .in1({ DP_IMM1_out_11 }),
  .out1({ S3145 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_505_ (
  .in1({ DP_IN_out_11 }),
  .out1({ S3146 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_506_ (
  .in1({ DP_IMM1_out_12 }),
  .out1({ S3147 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_507_ (
  .in1({ DP_IN_out_12 }),
  .out1({ S3148 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_508_ (
  .in1({ DP_IMM1_out_13 }),
  .out1({ S3149 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_509_ (
  .in1({ DP_IN_out_13 }),
  .out1({ S3150 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_510_ (
  .in1({ DP_IMM1_out_14 }),
  .out1({ S3151 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_511_ (
  .in1({ DP_IN_out_14 }),
  .out1({ S3152 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_512_ (
  .in1({ DP_IMM1_out_15 }),
  .out1({ S3153 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_513_ (
  .in1({ DP_IN_out_15 }),
  .out1({ S3154 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_514_ (
  .in1({ 1'bz }),
  .out1({ S3155 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1685_ (
  .in1({ S3275, S3273 }),
  .out1({ S3156 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1686_ (
  .in1({ CU_ldIR, DP_INC_1_in_0 }),
  .out1({ S3157 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1687_ (
  .in1({ S3271, 1'bz }),
  .out1({ S3158 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1688_ (
  .in1({ S3158, S3157 }),
  .out1({ S3159 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_984_ (
  .in1({ S3159, S3156 }),
  .out1({ S3160 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1689_ (
  .in1({ CU_selIN_ADR, S3274 }),
  .out1({ S3161 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_985_ (
  .in1({ CU_selIN_ADR, S3273 }),
  .out1({ S3162 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1690_ (
  .in1({ S3162, S3272 }),
  .out1({ S3163 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1691_ (
  .in1({ S3163, S3161 }),
  .out1({ S3164 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_986_ (
  .in1({ S3164, S3160 }),
  .out1({ S3117 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1692_ (
  .in1({ 1'bz, S3271 }),
  .out1({ S3165 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1693_ (
  .in1({ DP_INC_1_in_1, CU_ldIR }),
  .out1({ S3166 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1694_ (
  .in1({ S3166, S3165 }),
  .out1({ S3167 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_987_ (
  .in1({ S3167, S3156 }),
  .out1({ S3168 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1695_ (
  .in1({ S3277, CU_selIN_ADR }),
  .out1({ S3169 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1696_ (
  .in1({ S3162, S3276 }),
  .out1({ S3170 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1697_ (
  .in1({ S3170, S3169 }),
  .out1({ S3171 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_988_ (
  .in1({ S3171, S3168 }),
  .out1({ S3124 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1698_ (
  .in1({ 1'bz, S3271 }),
  .out1({ S3172 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1699_ (
  .in1({ DP_INC_1_in_2, CU_ldIR }),
  .out1({ S3173 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1700_ (
  .in1({ S3173, S3172 }),
  .out1({ S3174 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_989_ (
  .in1({ S3174, S3156 }),
  .out1({ S3175 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1701_ (
  .in1({ S3279, CU_selIN_ADR }),
  .out1({ S3176 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1702_ (
  .in1({ S3162, S3278 }),
  .out1({ S3177 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1703_ (
  .in1({ S3177, S3176 }),
  .out1({ S3178 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_990_ (
  .in1({ S3178, S3175 }),
  .out1({ S3125 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1704_ (
  .in1({ 1'bz, S3271 }),
  .out1({ S3179 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1705_ (
  .in1({ DP_INC_1_in_3, CU_ldIR }),
  .out1({ S3180 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1706_ (
  .in1({ S3180, S3179 }),
  .out1({ S3181 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_991_ (
  .in1({ S3181, S3156 }),
  .out1({ S3182 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1707_ (
  .in1({ S3281, CU_selIN_ADR }),
  .out1({ S3183 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1708_ (
  .in1({ S3162, S3280 }),
  .out1({ S3184 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1709_ (
  .in1({ S3184, S3183 }),
  .out1({ S3185 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_992_ (
  .in1({ S3185, S3182 }),
  .out1({ S3126 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1710_ (
  .in1({ 1'bz, S3271 }),
  .out1({ S3186 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1711_ (
  .in1({ DP_INC_1_in_4, CU_ldIR }),
  .out1({ S3187 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1712_ (
  .in1({ S3187, S3186 }),
  .out1({ S3188 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_993_ (
  .in1({ S3188, S3156 }),
  .out1({ S3189 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1713_ (
  .in1({ S3283, CU_selIN_ADR }),
  .out1({ S3190 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1714_ (
  .in1({ S3162, S3282 }),
  .out1({ S3191 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1715_ (
  .in1({ S3191, S3190 }),
  .out1({ S3192 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_994_ (
  .in1({ S3192, S3189 }),
  .out1({ S3127 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1716_ (
  .in1({ 1'bz, S3271 }),
  .out1({ S3193 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1717_ (
  .in1({ DP_INC_1_in_5, CU_ldIR }),
  .out1({ S3194 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1718_ (
  .in1({ S3194, S3193 }),
  .out1({ S3195 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_995_ (
  .in1({ S3195, S3156 }),
  .out1({ S3196 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1719_ (
  .in1({ S3134, CU_selIN_ADR }),
  .out1({ S3197 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1720_ (
  .in1({ S3162, S3284 }),
  .out1({ S3198 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1721_ (
  .in1({ S3198, S3197 }),
  .out1({ S3199 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_996_ (
  .in1({ S3199, S3196 }),
  .out1({ S3128 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1722_ (
  .in1({ 1'bz, S3271 }),
  .out1({ S3200 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1723_ (
  .in1({ DP_INC_1_in_6, CU_ldIR }),
  .out1({ S3201 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1724_ (
  .in1({ S3201, S3200 }),
  .out1({ S3202 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_997_ (
  .in1({ S3202, S3156 }),
  .out1({ S3203 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1725_ (
  .in1({ S3136, CU_selIN_ADR }),
  .out1({ S3204 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1726_ (
  .in1({ S3162, S3135 }),
  .out1({ S3205 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1727_ (
  .in1({ S3205, S3204 }),
  .out1({ S3206 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_998_ (
  .in1({ S3206, S3203 }),
  .out1({ S3129 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1728_ (
  .in1({ 1'bz, S3271 }),
  .out1({ S3207 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1729_ (
  .in1({ DP_INC_1_in_7, CU_ldIR }),
  .out1({ S3208 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1730_ (
  .in1({ S3208, S3207 }),
  .out1({ S3209 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_999_ (
  .in1({ S3209, S3156 }),
  .out1({ S3210 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1731_ (
  .in1({ S3138, CU_selIN_ADR }),
  .out1({ S3211 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1732_ (
  .in1({ S3162, S3137 }),
  .out1({ S3212 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1733_ (
  .in1({ S3212, S3211 }),
  .out1({ S3213 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1000_ (
  .in1({ S3213, S3210 }),
  .out1({ S3130 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1734_ (
  .in1({ DP_INC_1_in_8, CU_ldIR }),
  .out1({ S3214 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1735_ (
  .in1({ 1'bz, S3271 }),
  .out1({ S3215 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1736_ (
  .in1({ S3215, S3214 }),
  .out1({ S3216 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1001_ (
  .in1({ S3216, S3156 }),
  .out1({ S3217 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1737_ (
  .in1({ S3140, CU_selIN_ADR }),
  .out1({ S3218 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1738_ (
  .in1({ S3162, S3139 }),
  .out1({ S3219 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1739_ (
  .in1({ S3219, S3218 }),
  .out1({ S3220 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1002_ (
  .in1({ S3220, S3217 }),
  .out1({ S3131 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1740_ (
  .in1({ 1'bz, S3271 }),
  .out1({ S3221 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1741_ (
  .in1({ DP_INC_1_in_9, CU_ldIR }),
  .out1({ S3222 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1742_ (
  .in1({ S3222, S3221 }),
  .out1({ S3223 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1003_ (
  .in1({ S3223, S3156 }),
  .out1({ S3224 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1743_ (
  .in1({ S3142, CU_selIN_ADR }),
  .out1({ S3225 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1744_ (
  .in1({ S3162, S3141 }),
  .out1({ S3226 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1745_ (
  .in1({ S3226, S3225 }),
  .out1({ S3227 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1004_ (
  .in1({ S3227, S3224 }),
  .out1({ S3132 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1746_ (
  .in1({ DP_INC_1_in_10, CU_ldIR }),
  .out1({ S3228 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1747_ (
  .in1({ 1'bz, S3271 }),
  .out1({ S3229 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1748_ (
  .in1({ S3229, S3228 }),
  .out1({ S3230 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1005_ (
  .in1({ S3230, S3156 }),
  .out1({ S3231 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1749_ (
  .in1({ S3144, CU_selIN_ADR }),
  .out1({ S3232 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1750_ (
  .in1({ S3162, S3143 }),
  .out1({ S3233 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1751_ (
  .in1({ S3233, S3232 }),
  .out1({ S3234 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1006_ (
  .in1({ S3234, S3231 }),
  .out1({ S3118 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1752_ (
  .in1({ 1'bz, S3271 }),
  .out1({ S3235 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1753_ (
  .in1({ DP_INC_1_in_11, CU_ldIR }),
  .out1({ S3236 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1754_ (
  .in1({ S3236, S3235 }),
  .out1({ S3237 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1007_ (
  .in1({ S3237, S3156 }),
  .out1({ S3238 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1755_ (
  .in1({ S3146, CU_selIN_ADR }),
  .out1({ S3239 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1756_ (
  .in1({ S3162, S3145 }),
  .out1({ S3240 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1757_ (
  .in1({ S3240, S3239 }),
  .out1({ S3241 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1008_ (
  .in1({ S3241, S3238 }),
  .out1({ S3119 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1758_ (
  .in1({ DP_INC_1_in_12, CU_ldIR }),
  .out1({ S3242 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1759_ (
  .in1({ 1'bz, S3271 }),
  .out1({ S3243 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1760_ (
  .in1({ S3243, S3242 }),
  .out1({ S3244 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1009_ (
  .in1({ S3244, S3156 }),
  .out1({ S3245 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1761_ (
  .in1({ S3148, CU_selIN_ADR }),
  .out1({ S3246 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1762_ (
  .in1({ S3162, S3147 }),
  .out1({ S3247 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1763_ (
  .in1({ S3247, S3246 }),
  .out1({ S3248 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1010_ (
  .in1({ S3248, S3245 }),
  .out1({ S3120 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1764_ (
  .in1({ 1'bz, S3271 }),
  .out1({ S3249 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1765_ (
  .in1({ DP_INC_1_in_13, CU_ldIR }),
  .out1({ S3250 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1766_ (
  .in1({ S3250, S3249 }),
  .out1({ S3251 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1011_ (
  .in1({ S3251, S3156 }),
  .out1({ S3252 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1767_ (
  .in1({ S3150, CU_selIN_ADR }),
  .out1({ S3253 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1768_ (
  .in1({ S3162, S3149 }),
  .out1({ S3254 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1769_ (
  .in1({ S3254, S3253 }),
  .out1({ S3255 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1012_ (
  .in1({ S3255, S3252 }),
  .out1({ S3121 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1770_ (
  .in1({ DP_INC_1_in_14, CU_ldIR }),
  .out1({ S3256 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1771_ (
  .in1({ 1'bz, S3271 }),
  .out1({ S3257 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1772_ (
  .in1({ S3257, S3256 }),
  .out1({ S3258 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1013_ (
  .in1({ S3258, S3156 }),
  .out1({ S3259 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1773_ (
  .in1({ S3152, CU_selIN_ADR }),
  .out1({ S3260 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1774_ (
  .in1({ S3162, S3151 }),
  .out1({ S3261 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1775_ (
  .in1({ S3261, S3260 }),
  .out1({ S3262 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1014_ (
  .in1({ S3262, S3259 }),
  .out1({ S3122 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1776_ (
  .in1({ 1'bz, S3271 }),
  .out1({ S3263 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1777_ (
  .in1({ DP_INC_1_in_15, CU_ldIR }),
  .out1({ S3264 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1778_ (
  .in1({ S3264, S3263 }),
  .out1({ S3265 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1015_ (
  .in1({ S3265, S3156 }),
  .out1({ S3266 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1779_ (
  .in1({ S3154, CU_selIN_ADR }),
  .out1({ S3267 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1780_ (
  .in1({ S3162, S3153 }),
  .out1({ S3268 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1781_ (
  .in1({ S3268, S3267 }),
  .out1({ S3269 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1016_ (
  .in1({ S3269, S3266 }),
  .out1({ S3123 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1782_ (
  .in1({ S3155, S3271 }),
  .out1({ S3270 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1017_ (
  .in1({ S3270, S3156 }),
  .out1({ S3133 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__155_ (
  .D({ S3117 }),
  .E({ S3133 }),
  .Q({ DP_addrBus_0 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__156_ (
  .D({ S3124 }),
  .E({ S3133 }),
  .Q({ DP_addrBus_1 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__157_ (
  .D({ S3125 }),
  .E({ S3133 }),
  .Q({ DP_addrBus_2 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__158_ (
  .D({ S3126 }),
  .E({ S3133 }),
  .Q({ DP_addrBus_3 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__159_ (
  .D({ S3127 }),
  .E({ S3133 }),
  .Q({ DP_addrBus_4 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__160_ (
  .D({ S3128 }),
  .E({ S3133 }),
  .Q({ DP_addrBus_5 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__161_ (
  .D({ S3129 }),
  .E({ S3133 }),
  .Q({ DP_addrBus_6 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__162_ (
  .D({ S3130 }),
  .E({ S3133 }),
  .Q({ DP_addrBus_7 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__163_ (
  .D({ S3131 }),
  .E({ S3133 }),
  .Q({ DP_addrBus_8 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__164_ (
  .D({ S3132 }),
  .E({ S3133 }),
  .Q({ DP_addrBus_9 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__165_ (
  .D({ S3118 }),
  .E({ S3133 }),
  .Q({ DP_addrBus_10 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__166_ (
  .D({ S3119 }),
  .E({ S3133 }),
  .Q({ DP_addrBus_11 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__167_ (
  .D({ S3120 }),
  .E({ S3133 }),
  .Q({ DP_addrBus_12 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__168_ (
  .D({ S3121 }),
  .E({ S3133 }),
  .Q({ DP_addrBus_13 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__169_ (
  .D({ S3122 }),
  .E({ S3133 }),
  .Q({ DP_addrBus_14 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__170_ (
  .D({ S3123 }),
  .E({ S3133 }),
  .Q({ DP_addrBus_15 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_515_ (
  .in1({ CU_INC2 }),
  .out1({ S3288 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1783_ (
  .in1({ CU_INC2, S36 }),
  .out1({ S3289 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1784_ (
  .in1({ S3288, S4 }),
  .out1({ S3290 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1785_ (
  .in1({ S3290, S3289 }),
  .out1({ S3285 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1786_ (
  .in1({ S5, CU_INC2 }),
  .out1({ S3291 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1787_ (
  .in1({ S37, S3288 }),
  .out1({ S3292 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1788_ (
  .in1({ S3292, S3291 }),
  .out1({ S3286 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1018_ (
  .in1({ CU_INC1, CU_INC2 }),
  .out1({ S3287 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__171_ (
  .D({ S3285 }),
  .E({ S3287 }),
  .Q({ DP_INC_1_inc_val_0 })
);
$_DLATCH_N_ #() 
$_DLATCH_N__172_ (
  .D({ S3286 }),
  .E({ S3287 }),
  .Q({ DP_INC_1_inc_val_1 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_39_ (
  .in1({ DP_addrBus_0 }),
  .out1({ addrBus[0] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_40_ (
  .in1({ DP_addrBus_1 }),
  .out1({ addrBus[1] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_41_ (
  .in1({ DP_addrBus_10 }),
  .out1({ addrBus[10] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_42_ (
  .in1({ DP_addrBus_11 }),
  .out1({ addrBus[11] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_43_ (
  .in1({ DP_addrBus_12 }),
  .out1({ addrBus[12] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_44_ (
  .in1({ DP_addrBus_13 }),
  .out1({ addrBus[13] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_45_ (
  .in1({ DP_addrBus_14 }),
  .out1({ addrBus[14] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_46_ (
  .in1({ DP_addrBus_15 }),
  .out1({ addrBus[15] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_47_ (
  .in1({ DP_addrBus_2 }),
  .out1({ addrBus[2] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_48_ (
  .in1({ DP_addrBus_3 }),
  .out1({ addrBus[3] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_49_ (
  .in1({ DP_addrBus_4 }),
  .out1({ addrBus[4] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_50_ (
  .in1({ DP_addrBus_5 }),
  .out1({ addrBus[5] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_51_ (
  .in1({ DP_addrBus_6 }),
  .out1({ addrBus[6] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_52_ (
  .in1({ DP_addrBus_7 }),
  .out1({ addrBus[7] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_53_ (
  .in1({ DP_addrBus_8 }),
  .out1({ addrBus[8] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_54_ (
  .in1({ DP_addrBus_9 }),
  .out1({ addrBus[9] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_55_ (
  .in1({ clk }),
  .out1({ CU_clk })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_56_ (
  .in1({ CU_readMEM }),
  .out1({ readMEM })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_57_ (
  .in1({ rst }),
  .out1({ CU_rst })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_58_ (
  .in1({ CU_seldataBus }),
  .out1({ writeMEM })
);

endmodule