module fulladder(i0, i1, ci, s, co);

wire S0;
wire S1;
wire S2;
wire S3;
wire S4;
wire S5;
wire S6;
wire S7;
wire S8;
wire S9;
wire S10;
wire S11;
wire S12;
wire S13;
wire S14;
wire S15;
wire S16;
input i0;
input i1;
input ci;
output s;
output co;

nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_0_ (
  .in({ S12, S15 }),
  .out({ S11 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1_ (
  .in({ S10, S8 }),
  .out({ S0 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2_ (
  .in({ S12, S15 }),
  .out({ S1 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3_ (
  .in({ S1 }),
  .out({ S2 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4_ (
  .in({ S2, S11 }),
  .out({ S3 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5_ (
  .in({ S1, S0 }),
  .out({ S4 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6_ (
  .in({ S4, S14 }),
  .out({ S5 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_7_ (
  .in({ S3, S9 }),
  .out({ S6 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_8_ (
  .in({ S6, S5 }),
  .out({ S16 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_9_ (
  .in({ S0, S14 }),
  .out({ S7 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_10_ (
  .in({ S7, S1 }),
  .out({ S13 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_11_ (
  .in({ S15 }),
  .out({ S8 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_12_ (
  .in({ S14 }),
  .out({ S9 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_13_ (
  .in({ S12 }),
  .out({ S10 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_14_ (
  .in({ ci }),
  .out({ S12 })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_15_ (
  .in({ S13 }),
  .out({ co })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_16_ (
  .in({ i0 }),
  .out({ S14 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_17_ (
  .in({ i1 }),
  .out({ S15 })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_18_ (
  .in({ S16 }),
  .out({ s })
);

endmodule