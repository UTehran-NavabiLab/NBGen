module c432 (N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, N421, N430, N431, N432);

input N1;
input N4;
input N8;
input N11;
input N14;
input N17;
input N21;
input N24;
input N27;
input N30;
input N34;
input N37;
input N40;
input N43;
input N47;
input N50;
input N53;
input N56;
input N60;
input N63;
input N66;
input N69;
input N73;
input N76;
input N79;
input N82;
input N86;
input N89;
input N92;
input N95;
input N99;
input N102;
input N105;
input N108;
input N112;
input N115;
output N223;
output N329;
output N370;
output N421;
output N430;
output N431;
output N432;

INV_X1 INV_X1_1 ( .A(N56), .ZN(_69_) );
NOR2_X1 NOR2_X1_1 ( .A1(_69_), .A2(N60), .ZN(_70_) );
INV_X1 INV_X1_2 ( .A(N50), .ZN(_71_) );
INV_X1 INV_X1_3 ( .A(N89), .ZN(_72_) );
AOI22_X1 AOI22_X1_1 ( .A1(N56), .A2(_71_), .B1(_72_), .B2(N95), .ZN(_73_) );
INV_X1 INV_X1_4 ( .A(N1), .ZN(_74_) );
INV_X1 INV_X1_5 ( .A(N37), .ZN(_75_) );
AOI22_X1 AOI22_X1_2 ( .A1(_74_), .A2(N4), .B1(_75_), .B2(N43), .ZN(_76_) );
INV_X1 INV_X1_6 ( .A(N11), .ZN(_77_) );
INV_X1 INV_X1_7 ( .A(N24), .ZN(_78_) );
AOI22_X1 AOI22_X1_3 ( .A1(N17), .A2(_77_), .B1(_78_), .B2(N30), .ZN(_79_) );
INV_X1 INV_X1_8 ( .A(N63), .ZN(_80_) );
INV_X1 INV_X1_9 ( .A(N76), .ZN(_81_) );
AOI22_X1 AOI22_X1_4 ( .A1(N69), .A2(_80_), .B1(_81_), .B2(N82), .ZN(_82_) );
NAND4_X1 NAND4_X1_1 ( .A1(_73_), .A2(_76_), .A3(_79_), .A4(_82_), .ZN(_83_) );
INV_X1 INV_X1_10 ( .A(N102), .ZN(_84_) );
AND2_X1 AND2_X1_1 ( .A1(_84_), .A2(N108), .ZN(_85_) );
OAI21_X1 OAI21_X1_1 ( .A(N50), .B1(_83_), .B2(_85_), .ZN(_86_) );
NAND2_X1 NAND2_X1_1 ( .A1(_86_), .A2(_70_), .ZN(_87_) );
INV_X1 INV_X1_11 ( .A(_87_), .ZN(_88_) );
NOR2_X1 NOR2_X1_2 ( .A1(_83_), .A2(_85_), .ZN(_89_) );
OAI21_X1 OAI21_X1_2 ( .A(N108), .B1(_89_), .B2(_84_), .ZN(_90_) );
NOR2_X1 NOR2_X1_3 ( .A1(_90_), .A2(N112), .ZN(_91_) );
INV_X1 INV_X1_12 ( .A(N43), .ZN(_92_) );
NOR2_X1 NOR2_X1_4 ( .A1(_92_), .A2(N47), .ZN(_93_) );
OAI21_X1 OAI21_X1_3 ( .A(N37), .B1(_83_), .B2(_85_), .ZN(_94_) );
INV_X1 INV_X1_13 ( .A(N82), .ZN(_95_) );
NOR2_X1 NOR2_X1_5 ( .A1(_95_), .A2(N86), .ZN(_96_) );
OAI21_X1 OAI21_X1_4 ( .A(N76), .B1(_83_), .B2(_85_), .ZN(_97_) );
AOI22_X1 AOI22_X1_5 ( .A1(_93_), .A2(_94_), .B1(_97_), .B2(_96_), .ZN(_98_) );
INV_X1 INV_X1_14 ( .A(N69), .ZN(_99_) );
NOR2_X1 NOR2_X1_6 ( .A1(_99_), .A2(N73), .ZN(_100_) );
OAI21_X1 OAI21_X1_5 ( .A(N63), .B1(_83_), .B2(_85_), .ZN(_101_) );
AOI22_X1 AOI22_X1_6 ( .A1(_100_), .A2(_101_), .B1(_86_), .B2(_70_), .ZN(_102_) );
INV_X1 INV_X1_15 ( .A(N4), .ZN(_103_) );
NOR2_X1 NOR2_X1_7 ( .A1(_103_), .A2(N8), .ZN(_104_) );
OAI21_X1 OAI21_X1_6 ( .A(N1), .B1(_83_), .B2(_85_), .ZN(_105_) );
INV_X1 INV_X1_16 ( .A(N17), .ZN(_106_) );
NOR2_X1 NOR2_X1_8 ( .A1(_106_), .A2(N21), .ZN(_107_) );
OAI21_X1 OAI21_X1_7 ( .A(N11), .B1(_83_), .B2(_85_), .ZN(_108_) );
AOI22_X1 AOI22_X1_7 ( .A1(_104_), .A2(_105_), .B1(_108_), .B2(_107_), .ZN(_109_) );
INV_X1 INV_X1_17 ( .A(N95), .ZN(_110_) );
NOR2_X1 NOR2_X1_9 ( .A1(_110_), .A2(N99), .ZN(_111_) );
OAI21_X1 OAI21_X1_8 ( .A(N89), .B1(_83_), .B2(_85_), .ZN(_112_) );
INV_X1 INV_X1_18 ( .A(N30), .ZN(_113_) );
NOR2_X1 NOR2_X1_10 ( .A1(_113_), .A2(N34), .ZN(_114_) );
OAI21_X1 OAI21_X1_9 ( .A(N24), .B1(_83_), .B2(_85_), .ZN(_115_) );
AOI22_X1 AOI22_X1_8 ( .A1(_111_), .A2(_112_), .B1(_115_), .B2(_114_), .ZN(_116_) );
NAND4_X1 NAND4_X1_2 ( .A1(_98_), .A2(_102_), .A3(_109_), .A4(_116_), .ZN(_117_) );
NOR2_X1 NOR2_X1_11 ( .A1(_117_), .A2(_91_), .ZN(_118_) );
NAND2_X1 NAND2_X1_2 ( .A1(_86_), .A2(N56), .ZN(_119_) );
NOR2_X1 NOR2_X1_12 ( .A1(_119_), .A2(N66), .ZN(_120_) );
OAI21_X1 OAI21_X1_10 ( .A(_120_), .B1(_118_), .B2(_88_), .ZN(_121_) );
INV_X1 INV_X1_19 ( .A(N115), .ZN(_122_) );
AOI21_X1 AOI21_X1_1 ( .A(_90_), .B1(_117_), .B2(N112), .ZN(_123_) );
NAND2_X1 NAND2_X1_3 ( .A1(_123_), .A2(_122_), .ZN(_124_) );
NAND2_X1 NAND2_X1_4 ( .A1(_108_), .A2(_107_), .ZN(_0_) );
INV_X1 INV_X1_20 ( .A(_0_), .ZN(_1_) );
NAND2_X1 NAND2_X1_5 ( .A1(_108_), .A2(N17), .ZN(_2_) );
NOR2_X1 NOR2_X1_13 ( .A1(_2_), .A2(N27), .ZN(_3_) );
OAI21_X1 OAI21_X1_11 ( .A(_3_), .B1(_118_), .B2(_1_), .ZN(_4_) );
NAND2_X1 NAND2_X1_6 ( .A1(_105_), .A2(_104_), .ZN(_5_) );
INV_X1 INV_X1_21 ( .A(_5_), .ZN(_6_) );
NAND2_X1 NAND2_X1_7 ( .A1(_105_), .A2(N4), .ZN(_7_) );
NOR2_X1 NOR2_X1_14 ( .A1(_7_), .A2(N14), .ZN(_8_) );
OAI21_X1 OAI21_X1_12 ( .A(_8_), .B1(_118_), .B2(_6_), .ZN(_9_) );
NAND4_X1 NAND4_X1_3 ( .A1(_121_), .A2(_4_), .A3(_9_), .A4(_124_), .ZN(_10_) );
NAND2_X1 NAND2_X1_8 ( .A1(_97_), .A2(_96_), .ZN(_11_) );
INV_X1 INV_X1_22 ( .A(_11_), .ZN(_12_) );
NAND2_X1 NAND2_X1_9 ( .A1(_97_), .A2(N82), .ZN(_13_) );
NOR2_X1 NOR2_X1_15 ( .A1(_13_), .A2(N92), .ZN(_14_) );
OAI21_X1 OAI21_X1_13 ( .A(_14_), .B1(_118_), .B2(_12_), .ZN(_15_) );
NAND2_X1 NAND2_X1_10 ( .A1(_101_), .A2(_100_), .ZN(_16_) );
OAI21_X1 OAI21_X1_14 ( .A(_16_), .B1(_117_), .B2(_91_), .ZN(_17_) );
NAND2_X1 NAND2_X1_11 ( .A1(_101_), .A2(N69), .ZN(_18_) );
NOR2_X1 NOR2_X1_16 ( .A1(_18_), .A2(N79), .ZN(_19_) );
NAND2_X1 NAND2_X1_12 ( .A1(_112_), .A2(_111_), .ZN(_20_) );
OAI21_X1 OAI21_X1_15 ( .A(_20_), .B1(_117_), .B2(_91_), .ZN(_21_) );
NAND2_X1 NAND2_X1_13 ( .A1(_112_), .A2(N95), .ZN(_22_) );
NOR2_X1 NOR2_X1_17 ( .A1(_22_), .A2(N105), .ZN(_23_) );
AOI22_X1 AOI22_X1_9 ( .A1(_17_), .A2(_19_), .B1(_21_), .B2(_23_), .ZN(_24_) );
NAND2_X1 NAND2_X1_14 ( .A1(_94_), .A2(_93_), .ZN(_25_) );
OAI21_X1 OAI21_X1_16 ( .A(_25_), .B1(_117_), .B2(_91_), .ZN(_26_) );
NAND2_X1 NAND2_X1_15 ( .A1(_94_), .A2(N43), .ZN(_27_) );
NOR2_X1 NOR2_X1_18 ( .A1(_27_), .A2(N53), .ZN(_28_) );
NAND2_X1 NAND2_X1_16 ( .A1(_115_), .A2(_114_), .ZN(_29_) );
OAI21_X1 OAI21_X1_17 ( .A(_29_), .B1(_117_), .B2(_91_), .ZN(_30_) );
NAND2_X1 NAND2_X1_17 ( .A1(_115_), .A2(N30), .ZN(_31_) );
NOR2_X1 NOR2_X1_19 ( .A1(_31_), .A2(N40), .ZN(_32_) );
AOI22_X1 AOI22_X1_10 ( .A1(_26_), .A2(_28_), .B1(_30_), .B2(_32_), .ZN(_33_) );
NAND3_X1 NAND3_X1_1 ( .A1(_24_), .A2(_33_), .A3(_15_), .ZN(_34_) );
OAI21_X1 OAI21_X1_18 ( .A(N40), .B1(_34_), .B2(_10_), .ZN(_35_) );
INV_X1 INV_X1_23 ( .A(_118_), .ZN(_126_) );
AOI21_X1 AOI21_X1_2 ( .A(_31_), .B1(_126_), .B2(N34), .ZN(_36_) );
NAND2_X1 NAND2_X1_18 ( .A1(_35_), .A2(_36_), .ZN(_37_) );
OAI21_X1 OAI21_X1_19 ( .A(N27), .B1(_34_), .B2(_10_), .ZN(_38_) );
AOI21_X1 AOI21_X1_3 ( .A(_2_), .B1(_126_), .B2(N21), .ZN(_39_) );
NAND2_X1 NAND2_X1_19 ( .A1(_38_), .A2(_39_), .ZN(_40_) );
OAI21_X1 OAI21_X1_20 ( .A(N66), .B1(_34_), .B2(_10_), .ZN(_41_) );
AOI21_X1 AOI21_X1_4 ( .A(_119_), .B1(_126_), .B2(N60), .ZN(_42_) );
NAND2_X1 NAND2_X1_20 ( .A1(_41_), .A2(_42_), .ZN(_43_) );
OAI21_X1 OAI21_X1_21 ( .A(N53), .B1(_34_), .B2(_10_), .ZN(_44_) );
AOI21_X1 AOI21_X1_5 ( .A(_27_), .B1(_126_), .B2(N47), .ZN(_45_) );
NAND2_X1 NAND2_X1_21 ( .A1(_44_), .A2(_45_), .ZN(_46_) );
AND4_X1 AND4_X1_1 ( .A1(_37_), .A2(_40_), .A3(_43_), .A4(_46_), .ZN(_47_) );
OAI21_X1 OAI21_X1_22 ( .A(N115), .B1(_34_), .B2(_10_), .ZN(_48_) );
NAND2_X1 NAND2_X1_22 ( .A1(_48_), .A2(_123_), .ZN(_49_) );
AOI21_X1 AOI21_X1_6 ( .A(_22_), .B1(_126_), .B2(N99), .ZN(_50_) );
OAI21_X1 OAI21_X1_23 ( .A(N105), .B1(_34_), .B2(_10_), .ZN(_51_) );
NAND2_X1 NAND2_X1_23 ( .A1(_51_), .A2(_50_), .ZN(_52_) );
OAI21_X1 OAI21_X1_24 ( .A(N92), .B1(_34_), .B2(_10_), .ZN(_53_) );
AOI21_X1 AOI21_X1_7 ( .A(_13_), .B1(_126_), .B2(N86), .ZN(_54_) );
NAND2_X1 NAND2_X1_24 ( .A1(_53_), .A2(_54_), .ZN(_55_) );
AOI21_X1 AOI21_X1_8 ( .A(_18_), .B1(_126_), .B2(N73), .ZN(_56_) );
OAI21_X1 OAI21_X1_25 ( .A(N79), .B1(_34_), .B2(_10_), .ZN(_57_) );
NAND2_X1 NAND2_X1_25 ( .A1(_57_), .A2(_56_), .ZN(_58_) );
AND4_X1 AND4_X1_2 ( .A1(_49_), .A2(_52_), .A3(_55_), .A4(_58_), .ZN(_59_) );
OR2_X1 OR2_X1_1 ( .A1(_34_), .A2(_10_), .ZN(_127_) );
AND2_X1 AND2_X1_2 ( .A1(_126_), .A2(N8), .ZN(_60_) );
AOI211_X1 AOI211_X1_1 ( .A(_7_), .B(_60_), .C1(_127_), .C2(N14), .ZN(_61_) );
AOI21_X1 AOI21_X1_9 ( .A(_61_), .B1(_47_), .B2(_59_), .ZN(_128_) );
INV_X1 INV_X1_24 ( .A(_47_), .ZN(_129_) );
AND2_X1 AND2_X1_3 ( .A1(_37_), .A2(_40_), .ZN(_62_) );
NAND2_X1 NAND2_X1_26 ( .A1(_43_), .A2(_46_), .ZN(_63_) );
INV_X1 INV_X1_25 ( .A(_58_), .ZN(_64_) );
NAND4_X1 NAND4_X1_4 ( .A1(_64_), .A2(_37_), .A3(_43_), .A4(_46_), .ZN(_65_) );
OAI211_X1 OAI211_X1_1 ( .A(_65_), .B(_62_), .C1(_63_), .C2(_55_), .ZN(_130_) );
NAND3_X1 NAND3_X1_2 ( .A1(_37_), .A2(_46_), .A3(_55_), .ZN(_66_) );
AND2_X1 AND2_X1_4 ( .A1(_44_), .A2(_45_), .ZN(_67_) );
AOI22_X1 AOI22_X1_11 ( .A1(_67_), .A2(_37_), .B1(_38_), .B2(_39_), .ZN(_68_) );
OAI211_X1 OAI211_X1_2 ( .A(_65_), .B(_68_), .C1(_52_), .C2(_66_), .ZN(_131_) );
INV_X1 INV_X1_26 ( .A(_89_), .ZN(_125_) );
BUF_X1 BUF_X1_1 ( .A(_125_), .Z(N223) );
BUF_X1 BUF_X1_2 ( .A(_126_), .Z(N329) );
BUF_X1 BUF_X1_3 ( .A(_127_), .Z(N370) );
BUF_X1 BUF_X1_4 ( .A(_128_), .Z(N421) );
BUF_X1 BUF_X1_5 ( .A(_129_), .Z(N430) );
BUF_X1 BUF_X1_6 ( .A(_130_), .Z(N431) );
BUF_X1 BUF_X1_7 ( .A(_131_), .Z(N432) );
endmodule
