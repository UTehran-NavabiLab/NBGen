LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

ENTITY AES IS
    PORT (
        enable : IN STD_LOGIC;
        in : IN STD_LOGIC_VECTOR (127 DOWNTO 0);
        key128 : IN STD_LOGIC_VECTOR (127 DOWNTO 0);
        expected128 : IN STD_LOGIC_VECTOR (127 DOWNTO 0);
        decrypted128 : OUT STD_LOGIC_VECTOR (127 DOWNTO 0);
        encrypted128 : OUT STD_LOGIC_VECTOR (127 DOWNTO 0);
        e128 : OUT STD_LOGIC;
        d128 : OUT STD_LOGIC);
END ENTITY AES;

ARCHITECTURE arch OF AES IS
    SIGNAL S0 : STD_LOGIC;
    SIGNAL S1 : STD_LOGIC;
    SIGNAL S2 : STD_LOGIC;
    SIGNAL S3 : STD_LOGIC;
    SIGNAL S4 : STD_LOGIC;
    SIGNAL S5 : STD_LOGIC;
    SIGNAL S6 : STD_LOGIC;
    SIGNAL S7 : STD_LOGIC;
    SIGNAL S8 : STD_LOGIC;
    SIGNAL S9 : STD_LOGIC;
    SIGNAL S10 : STD_LOGIC;
    SIGNAL S11 : STD_LOGIC;
    SIGNAL S12 : STD_LOGIC;
    SIGNAL S13 : STD_LOGIC;
    SIGNAL S14 : STD_LOGIC;
    SIGNAL S15 : STD_LOGIC;
    SIGNAL S16 : STD_LOGIC;
    SIGNAL S17 : STD_LOGIC;
    SIGNAL S18 : STD_LOGIC;
    SIGNAL S19 : STD_LOGIC;
    SIGNAL S20 : STD_LOGIC;
    SIGNAL S21 : STD_LOGIC;
    SIGNAL S22 : STD_LOGIC;
    SIGNAL S23 : STD_LOGIC;
    SIGNAL S24 : STD_LOGIC;
    SIGNAL S25 : STD_LOGIC;
    SIGNAL S26 : STD_LOGIC;
    SIGNAL S27 : STD_LOGIC;
    SIGNAL S28 : STD_LOGIC;
    SIGNAL S29 : STD_LOGIC;
    SIGNAL S30 : STD_LOGIC;
    SIGNAL S31 : STD_LOGIC;
    SIGNAL S32 : STD_LOGIC;
    SIGNAL S33 : STD_LOGIC;
    SIGNAL S34 : STD_LOGIC;
    SIGNAL S35 : STD_LOGIC;
    SIGNAL S36 : STD_LOGIC;
    SIGNAL S37 : STD_LOGIC;
    SIGNAL S38 : STD_LOGIC;
    SIGNAL S39 : STD_LOGIC;
    SIGNAL S40 : STD_LOGIC;
    SIGNAL S41 : STD_LOGIC;
    SIGNAL S42 : STD_LOGIC;
    SIGNAL S43 : STD_LOGIC;
    SIGNAL S44 : STD_LOGIC;
    SIGNAL S45 : STD_LOGIC;
    SIGNAL S46 : STD_LOGIC;
    SIGNAL S47 : STD_LOGIC;
    SIGNAL S48 : STD_LOGIC;
    SIGNAL S49 : STD_LOGIC;
    SIGNAL S50 : STD_LOGIC;
    SIGNAL S51 : STD_LOGIC;
    SIGNAL S52 : STD_LOGIC;
    SIGNAL S53 : STD_LOGIC;
    SIGNAL S54 : STD_LOGIC;
    SIGNAL S55 : STD_LOGIC;
    SIGNAL S56 : STD_LOGIC;
    SIGNAL S57 : STD_LOGIC;
    SIGNAL S58 : STD_LOGIC;
    SIGNAL S59 : STD_LOGIC;
    SIGNAL S60 : STD_LOGIC;
    SIGNAL S61 : STD_LOGIC;
    SIGNAL S62 : STD_LOGIC;
    SIGNAL S63 : STD_LOGIC;
    SIGNAL S64 : STD_LOGIC;
    SIGNAL S65 : STD_LOGIC;
    SIGNAL S66 : STD_LOGIC;
    SIGNAL S67 : STD_LOGIC;
    SIGNAL S68 : STD_LOGIC;
    SIGNAL S69 : STD_LOGIC;
    SIGNAL S70 : STD_LOGIC;
    SIGNAL S71 : STD_LOGIC;
    SIGNAL S72 : STD_LOGIC;
    SIGNAL S73 : STD_LOGIC;
    SIGNAL S74 : STD_LOGIC;
    SIGNAL S75 : STD_LOGIC;
    SIGNAL S76 : STD_LOGIC;
    SIGNAL S77 : STD_LOGIC;
    SIGNAL S78 : STD_LOGIC;
    SIGNAL S79 : STD_LOGIC;
    SIGNAL S80 : STD_LOGIC;
    SIGNAL S81 : STD_LOGIC;
    SIGNAL S82 : STD_LOGIC;
    SIGNAL S83 : STD_LOGIC;
    SIGNAL S84 : STD_LOGIC;
    SIGNAL S85 : STD_LOGIC;
    SIGNAL S86 : STD_LOGIC;
    SIGNAL S87 : STD_LOGIC;
    SIGNAL S88 : STD_LOGIC;
    SIGNAL S89 : STD_LOGIC;
    SIGNAL S90 : STD_LOGIC;
    SIGNAL S91 : STD_LOGIC;
    SIGNAL S92 : STD_LOGIC;
    SIGNAL S93 : STD_LOGIC;
    SIGNAL S94 : STD_LOGIC;
    SIGNAL S95 : STD_LOGIC;
    SIGNAL S96 : STD_LOGIC;
    SIGNAL S97 : STD_LOGIC;
    SIGNAL S98 : STD_LOGIC;
    SIGNAL S99 : STD_LOGIC;
    SIGNAL S100 : STD_LOGIC;
    SIGNAL S101 : STD_LOGIC;
    SIGNAL S102 : STD_LOGIC;
    SIGNAL S103 : STD_LOGIC;
    SIGNAL S104 : STD_LOGIC;
    SIGNAL S105 : STD_LOGIC;
    SIGNAL S106 : STD_LOGIC;
    SIGNAL S107 : STD_LOGIC;
    SIGNAL S108 : STD_LOGIC;
    SIGNAL S109 : STD_LOGIC;
    SIGNAL S110 : STD_LOGIC;
    SIGNAL S111 : STD_LOGIC;
    SIGNAL S112 : STD_LOGIC;
    SIGNAL S113 : STD_LOGIC;
    SIGNAL S114 : STD_LOGIC;
    SIGNAL S115 : STD_LOGIC;
    SIGNAL S116 : STD_LOGIC;
    SIGNAL S117 : STD_LOGIC;
    SIGNAL S118 : STD_LOGIC;
    SIGNAL S119 : STD_LOGIC;
    SIGNAL S120 : STD_LOGIC;
    SIGNAL S121 : STD_LOGIC;
    SIGNAL S122 : STD_LOGIC;
    SIGNAL S123 : STD_LOGIC;
    SIGNAL S124 : STD_LOGIC;
    SIGNAL S125 : STD_LOGIC;
    SIGNAL S126 : STD_LOGIC;
    SIGNAL S127 : STD_LOGIC;
    SIGNAL S128 : STD_LOGIC;
    SIGNAL S129 : STD_LOGIC;
    SIGNAL S130 : STD_LOGIC;
    SIGNAL S131 : STD_LOGIC;
    SIGNAL S132 : STD_LOGIC;
    SIGNAL S133 : STD_LOGIC;
    SIGNAL S134 : STD_LOGIC;
    SIGNAL S135 : STD_LOGIC;
    SIGNAL S136 : STD_LOGIC;
    SIGNAL S137 : STD_LOGIC;
    SIGNAL S138 : STD_LOGIC;
    SIGNAL S139 : STD_LOGIC;
    SIGNAL S140 : STD_LOGIC;
    SIGNAL S141 : STD_LOGIC;
    SIGNAL S142 : STD_LOGIC;
    SIGNAL S143 : STD_LOGIC;
    SIGNAL S144 : STD_LOGIC;
    SIGNAL S145 : STD_LOGIC;
    SIGNAL S146 : STD_LOGIC;
    SIGNAL S147 : STD_LOGIC;
    SIGNAL S148 : STD_LOGIC;
    SIGNAL S149 : STD_LOGIC;
    SIGNAL S150 : STD_LOGIC;
    SIGNAL S151 : STD_LOGIC;
    SIGNAL S152 : STD_LOGIC;
    SIGNAL S153 : STD_LOGIC;
    SIGNAL S154 : STD_LOGIC;
    SIGNAL S155 : STD_LOGIC;
    SIGNAL S156 : STD_LOGIC;
    SIGNAL S157 : STD_LOGIC;
    SIGNAL S158 : STD_LOGIC;
    SIGNAL S159 : STD_LOGIC;
    SIGNAL S160 : STD_LOGIC;
    SIGNAL S161 : STD_LOGIC;
    SIGNAL S162 : STD_LOGIC;
    SIGNAL S163 : STD_LOGIC;
    SIGNAL S164 : STD_LOGIC;
    SIGNAL S165 : STD_LOGIC;
    SIGNAL S166 : STD_LOGIC;
    SIGNAL S167 : STD_LOGIC;
    SIGNAL S168 : STD_LOGIC;
    SIGNAL S169 : STD_LOGIC;
    SIGNAL S170 : STD_LOGIC;
    SIGNAL S171 : STD_LOGIC;
    SIGNAL S172 : STD_LOGIC;
    SIGNAL S173 : STD_LOGIC;
    SIGNAL S174 : STD_LOGIC;
    SIGNAL S175 : STD_LOGIC;
    SIGNAL S176 : STD_LOGIC;
    SIGNAL S177 : STD_LOGIC;
    SIGNAL S178 : STD_LOGIC;
    SIGNAL S179 : STD_LOGIC;
    SIGNAL S180 : STD_LOGIC;
    SIGNAL S181 : STD_LOGIC;
    SIGNAL S182 : STD_LOGIC;
    SIGNAL S183 : STD_LOGIC;
    SIGNAL S184 : STD_LOGIC;
    SIGNAL S185 : STD_LOGIC;
    SIGNAL S186 : STD_LOGIC;
    SIGNAL S187 : STD_LOGIC;
    SIGNAL S188 : STD_LOGIC;
    SIGNAL S189 : STD_LOGIC;
    SIGNAL S190 : STD_LOGIC;
    SIGNAL S191 : STD_LOGIC;
    SIGNAL S192 : STD_LOGIC;
    SIGNAL S193 : STD_LOGIC;
    SIGNAL S194 : STD_LOGIC;
    SIGNAL S195 : STD_LOGIC;
    SIGNAL S196 : STD_LOGIC;
    SIGNAL S197 : STD_LOGIC;
    SIGNAL S198 : STD_LOGIC;
    SIGNAL S199 : STD_LOGIC;
    SIGNAL S200 : STD_LOGIC;
    SIGNAL S201 : STD_LOGIC;
    SIGNAL S202 : STD_LOGIC;
    SIGNAL S203 : STD_LOGIC;
    SIGNAL S204 : STD_LOGIC;
    SIGNAL S205 : STD_LOGIC;
    SIGNAL S206 : STD_LOGIC;
    SIGNAL S207 : STD_LOGIC;
    SIGNAL S208 : STD_LOGIC;
    SIGNAL S209 : STD_LOGIC;
    SIGNAL S210 : STD_LOGIC;
    SIGNAL S211 : STD_LOGIC;
    SIGNAL S212 : STD_LOGIC;
    SIGNAL S213 : STD_LOGIC;
    SIGNAL S214 : STD_LOGIC;
    SIGNAL S215 : STD_LOGIC;
    SIGNAL S216 : STD_LOGIC;
    SIGNAL S217 : STD_LOGIC;
    SIGNAL S218 : STD_LOGIC;
    SIGNAL S219 : STD_LOGIC;
    SIGNAL S220 : STD_LOGIC;
    SIGNAL S221 : STD_LOGIC;
    SIGNAL S222 : STD_LOGIC;
    SIGNAL S223 : STD_LOGIC;
    SIGNAL S224 : STD_LOGIC;
    SIGNAL S225 : STD_LOGIC;
    SIGNAL S226 : STD_LOGIC;
    SIGNAL S227 : STD_LOGIC;
    SIGNAL S228 : STD_LOGIC;
    SIGNAL S229 : STD_LOGIC;
    SIGNAL S230 : STD_LOGIC;
    SIGNAL S231 : STD_LOGIC;
    SIGNAL S232 : STD_LOGIC;
    SIGNAL S233 : STD_LOGIC;
    SIGNAL S234 : STD_LOGIC;
    SIGNAL S235 : STD_LOGIC;
    SIGNAL S236 : STD_LOGIC;
    SIGNAL S237 : STD_LOGIC;
    SIGNAL S238 : STD_LOGIC;
    SIGNAL S239 : STD_LOGIC;
    SIGNAL S240 : STD_LOGIC;
    SIGNAL S241 : STD_LOGIC;
    SIGNAL S242 : STD_LOGIC;
    SIGNAL S243 : STD_LOGIC;
    SIGNAL S244 : STD_LOGIC;
    SIGNAL S245 : STD_LOGIC;
    SIGNAL S246 : STD_LOGIC;
    SIGNAL S247 : STD_LOGIC;
    SIGNAL S248 : STD_LOGIC;
    SIGNAL S249 : STD_LOGIC;
    SIGNAL S250 : STD_LOGIC;
    SIGNAL S251 : STD_LOGIC;
    SIGNAL S252 : STD_LOGIC;
    SIGNAL S253 : STD_LOGIC;
    SIGNAL S254 : STD_LOGIC;
    SIGNAL S255 : STD_LOGIC;
    SIGNAL S256 : STD_LOGIC;
    SIGNAL S257 : STD_LOGIC;
    SIGNAL S258 : STD_LOGIC;
    SIGNAL S259 : STD_LOGIC;
    SIGNAL S260 : STD_LOGIC;
    SIGNAL S261 : STD_LOGIC;
    SIGNAL S262 : STD_LOGIC;
    SIGNAL S263 : STD_LOGIC;
    SIGNAL S264 : STD_LOGIC;
    SIGNAL S265 : STD_LOGIC;
    SIGNAL S266 : STD_LOGIC;
    SIGNAL S267 : STD_LOGIC;
    SIGNAL S268 : STD_LOGIC;
    SIGNAL S269 : STD_LOGIC;
    SIGNAL S270 : STD_LOGIC;
    SIGNAL S271 : STD_LOGIC;
    SIGNAL S272 : STD_LOGIC;
    SIGNAL S273 : STD_LOGIC;
    SIGNAL S274 : STD_LOGIC;
    SIGNAL S275 : STD_LOGIC;
    SIGNAL S276 : STD_LOGIC;
    SIGNAL S277 : STD_LOGIC;
    SIGNAL S278 : STD_LOGIC;
    SIGNAL S279 : STD_LOGIC;
    SIGNAL S280 : STD_LOGIC;
    SIGNAL S281 : STD_LOGIC;
    SIGNAL S282 : STD_LOGIC;
    SIGNAL S283 : STD_LOGIC;
    SIGNAL S284 : STD_LOGIC;
    SIGNAL S285 : STD_LOGIC;
    SIGNAL S286 : STD_LOGIC;
    SIGNAL S287 : STD_LOGIC;
    SIGNAL S288 : STD_LOGIC;
    SIGNAL S289 : STD_LOGIC;
    SIGNAL S290 : STD_LOGIC;
    SIGNAL S291 : STD_LOGIC;
    SIGNAL S292 : STD_LOGIC;
    SIGNAL S293 : STD_LOGIC;
    SIGNAL S294 : STD_LOGIC;
    SIGNAL S295 : STD_LOGIC;
    SIGNAL S296 : STD_LOGIC;
    SIGNAL S297 : STD_LOGIC;
    SIGNAL S298 : STD_LOGIC;
    SIGNAL S299 : STD_LOGIC;
    SIGNAL S300 : STD_LOGIC;
    SIGNAL S301 : STD_LOGIC;
    SIGNAL S302 : STD_LOGIC;
    SIGNAL S303 : STD_LOGIC;
    SIGNAL S304 : STD_LOGIC;
    SIGNAL S305 : STD_LOGIC;
    SIGNAL S306 : STD_LOGIC;
    SIGNAL S307 : STD_LOGIC;
    SIGNAL S308 : STD_LOGIC;
    SIGNAL S309 : STD_LOGIC;
    SIGNAL S310 : STD_LOGIC;
    SIGNAL S311 : STD_LOGIC;
    SIGNAL S312 : STD_LOGIC;
    SIGNAL S313 : STD_LOGIC;
    SIGNAL S314 : STD_LOGIC;
    SIGNAL S315 : STD_LOGIC;
    SIGNAL S316 : STD_LOGIC;
    SIGNAL S317 : STD_LOGIC;
    SIGNAL S318 : STD_LOGIC;
    SIGNAL S319 : STD_LOGIC;
    SIGNAL S320 : STD_LOGIC;
    SIGNAL S321 : STD_LOGIC;
    SIGNAL S322 : STD_LOGIC;
    SIGNAL S323 : STD_LOGIC;
    SIGNAL S324 : STD_LOGIC;
    SIGNAL S325 : STD_LOGIC;
    SIGNAL S326 : STD_LOGIC;
    SIGNAL S327 : STD_LOGIC;
    SIGNAL S328 : STD_LOGIC;
    SIGNAL S329 : STD_LOGIC;
    SIGNAL S330 : STD_LOGIC;
    SIGNAL S331 : STD_LOGIC;
    SIGNAL S332 : STD_LOGIC;
    SIGNAL S333 : STD_LOGIC;
    SIGNAL S334 : STD_LOGIC;
    SIGNAL S335 : STD_LOGIC;
    SIGNAL S336 : STD_LOGIC;
    SIGNAL S337 : STD_LOGIC;
    SIGNAL S338 : STD_LOGIC;
    SIGNAL S339 : STD_LOGIC;
    SIGNAL S340 : STD_LOGIC;
    SIGNAL S341 : STD_LOGIC;
    SIGNAL S342 : STD_LOGIC;
    SIGNAL S343 : STD_LOGIC;
    SIGNAL S344 : STD_LOGIC;
    SIGNAL S345 : STD_LOGIC;
    SIGNAL S346 : STD_LOGIC;
    SIGNAL S347 : STD_LOGIC;
    SIGNAL S348 : STD_LOGIC;
    SIGNAL S349 : STD_LOGIC;
    SIGNAL S350 : STD_LOGIC;
    SIGNAL S351 : STD_LOGIC;
    SIGNAL S352 : STD_LOGIC;
    SIGNAL S353 : STD_LOGIC;
    SIGNAL S354 : STD_LOGIC;
    SIGNAL S355 : STD_LOGIC;
    SIGNAL S356 : STD_LOGIC;
    SIGNAL S357 : STD_LOGIC;
    SIGNAL S358 : STD_LOGIC;
    SIGNAL S359 : STD_LOGIC;
    SIGNAL S360 : STD_LOGIC;
    SIGNAL S361 : STD_LOGIC;
    SIGNAL S362 : STD_LOGIC;
    SIGNAL S363 : STD_LOGIC;
    SIGNAL S364 : STD_LOGIC;
    SIGNAL S365 : STD_LOGIC;
    SIGNAL S366 : STD_LOGIC;
    SIGNAL S367 : STD_LOGIC;
    SIGNAL S368 : STD_LOGIC;
    SIGNAL S369 : STD_LOGIC;
    SIGNAL S370 : STD_LOGIC;
    SIGNAL S371 : STD_LOGIC;
    SIGNAL S372 : STD_LOGIC;
    SIGNAL S373 : STD_LOGIC;
    SIGNAL S374 : STD_LOGIC;
    SIGNAL S375 : STD_LOGIC;
    SIGNAL S376 : STD_LOGIC;
    SIGNAL S377 : STD_LOGIC;
    SIGNAL S378 : STD_LOGIC;
    SIGNAL S379 : STD_LOGIC;
    SIGNAL S380 : STD_LOGIC;
    SIGNAL S381 : STD_LOGIC;
    SIGNAL S382 : STD_LOGIC;
    SIGNAL S383 : STD_LOGIC;
    SIGNAL S384 : STD_LOGIC;
    SIGNAL S385 : STD_LOGIC;
    SIGNAL S386 : STD_LOGIC;
    SIGNAL S387 : STD_LOGIC;
    SIGNAL S388 : STD_LOGIC;
    SIGNAL S389 : STD_LOGIC;
    SIGNAL S390 : STD_LOGIC;
    SIGNAL S391 : STD_LOGIC;
    SIGNAL S392 : STD_LOGIC;
    SIGNAL S393 : STD_LOGIC;
    SIGNAL S394 : STD_LOGIC;
    SIGNAL S395 : STD_LOGIC;
    SIGNAL S396 : STD_LOGIC;
    SIGNAL S397 : STD_LOGIC;
    SIGNAL S398 : STD_LOGIC;
    SIGNAL S399 : STD_LOGIC;
    SIGNAL S400 : STD_LOGIC;
    SIGNAL S401 : STD_LOGIC;
    SIGNAL S402 : STD_LOGIC;
    SIGNAL S403 : STD_LOGIC;
    SIGNAL S404 : STD_LOGIC;
    SIGNAL S405 : STD_LOGIC;
    SIGNAL S406 : STD_LOGIC;
    SIGNAL S407 : STD_LOGIC;
    SIGNAL S408 : STD_LOGIC;
    SIGNAL S409 : STD_LOGIC;
    SIGNAL S410 : STD_LOGIC;
    SIGNAL S411 : STD_LOGIC;
    SIGNAL S412 : STD_LOGIC;
    SIGNAL S413 : STD_LOGIC;
    SIGNAL S414 : STD_LOGIC;
    SIGNAL S415 : STD_LOGIC;
    SIGNAL S416 : STD_LOGIC;
    SIGNAL S417 : STD_LOGIC;
    SIGNAL S418 : STD_LOGIC;
    SIGNAL S419 : STD_LOGIC;
    SIGNAL S420 : STD_LOGIC;
    SIGNAL S421 : STD_LOGIC;
    SIGNAL S422 : STD_LOGIC;
    SIGNAL S423 : STD_LOGIC;
    SIGNAL S424 : STD_LOGIC;
    SIGNAL S425 : STD_LOGIC;
    SIGNAL S426 : STD_LOGIC;
    SIGNAL S427 : STD_LOGIC;
    SIGNAL S428 : STD_LOGIC;
    SIGNAL S429 : STD_LOGIC;
    SIGNAL S430 : STD_LOGIC;
    SIGNAL S431 : STD_LOGIC;
    SIGNAL S432 : STD_LOGIC;
    SIGNAL S433 : STD_LOGIC;
    SIGNAL S434 : STD_LOGIC;
    SIGNAL S435 : STD_LOGIC;
    SIGNAL S436 : STD_LOGIC;
    SIGNAL S437 : STD_LOGIC;
    SIGNAL S438 : STD_LOGIC;
    SIGNAL S439 : STD_LOGIC;
    SIGNAL S440 : STD_LOGIC;
    SIGNAL S441 : STD_LOGIC;
    SIGNAL S442 : STD_LOGIC;
    SIGNAL S443 : STD_LOGIC;
    SIGNAL S444 : STD_LOGIC;
    SIGNAL S445 : STD_LOGIC;
    SIGNAL S446 : STD_LOGIC;
    SIGNAL S447 : STD_LOGIC;
    SIGNAL S448 : STD_LOGIC;
    SIGNAL S449 : STD_LOGIC;
    SIGNAL S450 : STD_LOGIC;
    SIGNAL S451 : STD_LOGIC;
    SIGNAL S452 : STD_LOGIC;
    SIGNAL S453 : STD_LOGIC;
    SIGNAL S454 : STD_LOGIC;
    SIGNAL S455 : STD_LOGIC;
    SIGNAL S456 : STD_LOGIC;
    SIGNAL S457 : STD_LOGIC;
    SIGNAL S458 : STD_LOGIC;
    SIGNAL S459 : STD_LOGIC;
    SIGNAL S460 : STD_LOGIC;
    SIGNAL S461 : STD_LOGIC;
    SIGNAL S462 : STD_LOGIC;
    SIGNAL S463 : STD_LOGIC;
    SIGNAL S464 : STD_LOGIC;
    SIGNAL S465 : STD_LOGIC;
    SIGNAL S466 : STD_LOGIC;
    SIGNAL S467 : STD_LOGIC;
    SIGNAL S468 : STD_LOGIC;
    SIGNAL S469 : STD_LOGIC;
    SIGNAL S470 : STD_LOGIC;
    SIGNAL S471 : STD_LOGIC;
    SIGNAL S472 : STD_LOGIC;
    SIGNAL S473 : STD_LOGIC;
    SIGNAL S474 : STD_LOGIC;
    SIGNAL S475 : STD_LOGIC;
    SIGNAL S476 : STD_LOGIC;
    SIGNAL S477 : STD_LOGIC;
    SIGNAL S478 : STD_LOGIC;
    SIGNAL S479 : STD_LOGIC;
    SIGNAL S480 : STD_LOGIC;
    SIGNAL S481 : STD_LOGIC;
    SIGNAL S482 : STD_LOGIC;
    SIGNAL S483 : STD_LOGIC;
    SIGNAL S484 : STD_LOGIC;
    SIGNAL S485 : STD_LOGIC;
    SIGNAL S486 : STD_LOGIC;
    SIGNAL S487 : STD_LOGIC;
    SIGNAL S488 : STD_LOGIC;
    SIGNAL S489 : STD_LOGIC;
    SIGNAL S490 : STD_LOGIC;
    SIGNAL S491 : STD_LOGIC;
    SIGNAL S492 : STD_LOGIC;
    SIGNAL S493 : STD_LOGIC;
    SIGNAL S494 : STD_LOGIC;
    SIGNAL S495 : STD_LOGIC;
    SIGNAL S496 : STD_LOGIC;
    SIGNAL S497 : STD_LOGIC;
    SIGNAL S498 : STD_LOGIC;
    SIGNAL S499 : STD_LOGIC;
    SIGNAL S500 : STD_LOGIC;
    SIGNAL S501 : STD_LOGIC;
    SIGNAL S502 : STD_LOGIC;
    SIGNAL S503 : STD_LOGIC;
    SIGNAL S504 : STD_LOGIC;
    SIGNAL S505 : STD_LOGIC;
    SIGNAL S506 : STD_LOGIC;
    SIGNAL S507 : STD_LOGIC;
    SIGNAL S508 : STD_LOGIC;
    SIGNAL S509 : STD_LOGIC;
    SIGNAL S510 : STD_LOGIC;
    SIGNAL S511 : STD_LOGIC;
    SIGNAL S512 : STD_LOGIC;
    SIGNAL S513 : STD_LOGIC;
    SIGNAL S514 : STD_LOGIC;
    SIGNAL S515 : STD_LOGIC;
    SIGNAL S516 : STD_LOGIC;
    SIGNAL S517 : STD_LOGIC;
    SIGNAL S518 : STD_LOGIC;
    SIGNAL S519 : STD_LOGIC;
    SIGNAL S520 : STD_LOGIC;
    SIGNAL S521 : STD_LOGIC;
    SIGNAL S522 : STD_LOGIC;
    SIGNAL S523 : STD_LOGIC;
    SIGNAL S524 : STD_LOGIC;
    SIGNAL S525 : STD_LOGIC;
    SIGNAL S526 : STD_LOGIC;
    SIGNAL S527 : STD_LOGIC;
    SIGNAL S528 : STD_LOGIC;
    SIGNAL S529 : STD_LOGIC;
    SIGNAL S530 : STD_LOGIC;
    SIGNAL S531 : STD_LOGIC;
    SIGNAL S532 : STD_LOGIC;
    SIGNAL S533 : STD_LOGIC;
    SIGNAL S534 : STD_LOGIC;
    SIGNAL S535 : STD_LOGIC;
    SIGNAL S536 : STD_LOGIC;
    SIGNAL S537 : STD_LOGIC;
    SIGNAL S538 : STD_LOGIC;
    SIGNAL S539 : STD_LOGIC;
    SIGNAL S540 : STD_LOGIC;
    SIGNAL S541 : STD_LOGIC;
    SIGNAL S542 : STD_LOGIC;
    SIGNAL S543 : STD_LOGIC;
    SIGNAL S544 : STD_LOGIC;
    SIGNAL S545 : STD_LOGIC;
    SIGNAL S546 : STD_LOGIC;
    SIGNAL S547 : STD_LOGIC;
    SIGNAL S548 : STD_LOGIC;
    SIGNAL S549 : STD_LOGIC;
    SIGNAL S550 : STD_LOGIC;
    SIGNAL S551 : STD_LOGIC;
    SIGNAL S552 : STD_LOGIC;
    SIGNAL S553 : STD_LOGIC;
    SIGNAL S554 : STD_LOGIC;
    SIGNAL S555 : STD_LOGIC;
    SIGNAL S556 : STD_LOGIC;
    SIGNAL S557 : STD_LOGIC;
    SIGNAL S558 : STD_LOGIC;
    SIGNAL S559 : STD_LOGIC;
    SIGNAL S560 : STD_LOGIC;
    SIGNAL S561 : STD_LOGIC;
    SIGNAL S562 : STD_LOGIC;
    SIGNAL S563 : STD_LOGIC;
    SIGNAL S564 : STD_LOGIC;
    SIGNAL S565 : STD_LOGIC;
    SIGNAL S566 : STD_LOGIC;
    SIGNAL S567 : STD_LOGIC;
    SIGNAL S568 : STD_LOGIC;
    SIGNAL S569 : STD_LOGIC;
    SIGNAL S570 : STD_LOGIC;
    SIGNAL S571 : STD_LOGIC;
    SIGNAL S572 : STD_LOGIC;
    SIGNAL S573 : STD_LOGIC;
    SIGNAL S574 : STD_LOGIC;
    SIGNAL S575 : STD_LOGIC;
    SIGNAL S576 : STD_LOGIC;
    SIGNAL S577 : STD_LOGIC;
    SIGNAL S578 : STD_LOGIC;
    SIGNAL S579 : STD_LOGIC;
    SIGNAL S580 : STD_LOGIC;
    SIGNAL S581 : STD_LOGIC;
    SIGNAL S582 : STD_LOGIC;
    SIGNAL S583 : STD_LOGIC;
    SIGNAL S584 : STD_LOGIC;
    SIGNAL S585 : STD_LOGIC;
    SIGNAL S586 : STD_LOGIC;
    SIGNAL S587 : STD_LOGIC;
    SIGNAL S588 : STD_LOGIC;
    SIGNAL S589 : STD_LOGIC;
    SIGNAL S590 : STD_LOGIC;
    SIGNAL S591 : STD_LOGIC;
    SIGNAL S592 : STD_LOGIC;
    SIGNAL S593 : STD_LOGIC;
    SIGNAL S594 : STD_LOGIC;
    SIGNAL S595 : STD_LOGIC;
    SIGNAL S596 : STD_LOGIC;
    SIGNAL S597 : STD_LOGIC;
    SIGNAL S598 : STD_LOGIC;
    SIGNAL S599 : STD_LOGIC;
    SIGNAL S600 : STD_LOGIC;
    SIGNAL S601 : STD_LOGIC;
    SIGNAL S602 : STD_LOGIC;
    SIGNAL S603 : STD_LOGIC;
    SIGNAL S604 : STD_LOGIC;
    SIGNAL S605 : STD_LOGIC;
    SIGNAL S606 : STD_LOGIC;
    SIGNAL S607 : STD_LOGIC;
    SIGNAL S608 : STD_LOGIC;
    SIGNAL S609 : STD_LOGIC;
    SIGNAL S610 : STD_LOGIC;
    SIGNAL S611 : STD_LOGIC;
    SIGNAL S612 : STD_LOGIC;
    SIGNAL S613 : STD_LOGIC;
    SIGNAL S614 : STD_LOGIC;
    SIGNAL S615 : STD_LOGIC;
    SIGNAL S616 : STD_LOGIC;
    SIGNAL S617 : STD_LOGIC;
    SIGNAL S618 : STD_LOGIC;
    SIGNAL S619 : STD_LOGIC;
    SIGNAL S620 : STD_LOGIC;
    SIGNAL S621 : STD_LOGIC;
    SIGNAL S622 : STD_LOGIC;
    SIGNAL S623 : STD_LOGIC;
    SIGNAL S624 : STD_LOGIC;
    SIGNAL S625 : STD_LOGIC;
    SIGNAL S626 : STD_LOGIC;
    SIGNAL S627 : STD_LOGIC;
    SIGNAL S628 : STD_LOGIC;
    SIGNAL S629 : STD_LOGIC;
    SIGNAL S630 : STD_LOGIC;
    SIGNAL S631 : STD_LOGIC;
    SIGNAL S632 : STD_LOGIC;
    SIGNAL S633 : STD_LOGIC;
    SIGNAL S634 : STD_LOGIC;
    SIGNAL S635 : STD_LOGIC;
    SIGNAL S636 : STD_LOGIC;
    SIGNAL S637 : STD_LOGIC;
    SIGNAL S638 : STD_LOGIC;
    SIGNAL S639 : STD_LOGIC;
    SIGNAL S640 : STD_LOGIC;
    SIGNAL S641 : STD_LOGIC;
    SIGNAL S642 : STD_LOGIC;
    SIGNAL S643 : STD_LOGIC;
    SIGNAL S644 : STD_LOGIC;
    SIGNAL S645 : STD_LOGIC;
    SIGNAL S646 : STD_LOGIC;
    SIGNAL S647 : STD_LOGIC;
    SIGNAL S648 : STD_LOGIC;
    SIGNAL S649 : STD_LOGIC;
    SIGNAL S650 : STD_LOGIC;
    SIGNAL S651 : STD_LOGIC;
    SIGNAL S652 : STD_LOGIC;
    SIGNAL S653 : STD_LOGIC;
    SIGNAL S654 : STD_LOGIC;
    SIGNAL S655 : STD_LOGIC;
    SIGNAL S656 : STD_LOGIC;
    SIGNAL S657 : STD_LOGIC;
    SIGNAL S658 : STD_LOGIC;
    SIGNAL S659 : STD_LOGIC;
    SIGNAL S660 : STD_LOGIC;
    SIGNAL S661 : STD_LOGIC;
    SIGNAL S662 : STD_LOGIC;
    SIGNAL S663 : STD_LOGIC;
    SIGNAL S664 : STD_LOGIC;
    SIGNAL S665 : STD_LOGIC;
    SIGNAL S666 : STD_LOGIC;
    SIGNAL S667 : STD_LOGIC;
    SIGNAL S668 : STD_LOGIC;
    SIGNAL S669 : STD_LOGIC;
    SIGNAL S670 : STD_LOGIC;
    SIGNAL S671 : STD_LOGIC;
    SIGNAL S672 : STD_LOGIC;
    SIGNAL S673 : STD_LOGIC;
    SIGNAL S674 : STD_LOGIC;
    SIGNAL S675 : STD_LOGIC;
    SIGNAL S676 : STD_LOGIC;
    SIGNAL S677 : STD_LOGIC;
    SIGNAL S678 : STD_LOGIC;
    SIGNAL S679 : STD_LOGIC;
    SIGNAL S680 : STD_LOGIC;
    SIGNAL S681 : STD_LOGIC;
    SIGNAL S682 : STD_LOGIC;
    SIGNAL S683 : STD_LOGIC;
    SIGNAL S684 : STD_LOGIC;
    SIGNAL S685 : STD_LOGIC;
    SIGNAL S686 : STD_LOGIC;
    SIGNAL S687 : STD_LOGIC;
    SIGNAL S688 : STD_LOGIC;
    SIGNAL S689 : STD_LOGIC;
    SIGNAL S690 : STD_LOGIC;
    SIGNAL S691 : STD_LOGIC;
    SIGNAL S692 : STD_LOGIC;
    SIGNAL S693 : STD_LOGIC;
    SIGNAL S694 : STD_LOGIC;
    SIGNAL S695 : STD_LOGIC;
    SIGNAL S696 : STD_LOGIC;
    SIGNAL S697 : STD_LOGIC;
    SIGNAL S698 : STD_LOGIC;
    SIGNAL S699 : STD_LOGIC;
    SIGNAL S700 : STD_LOGIC;
    SIGNAL S701 : STD_LOGIC;
    SIGNAL S702 : STD_LOGIC;
    SIGNAL S703 : STD_LOGIC;
    SIGNAL S704 : STD_LOGIC;
    SIGNAL S705 : STD_LOGIC;
    SIGNAL S706 : STD_LOGIC;
    SIGNAL S707 : STD_LOGIC;
    SIGNAL S708 : STD_LOGIC;
    SIGNAL S709 : STD_LOGIC;
    SIGNAL S710 : STD_LOGIC;
    SIGNAL S711 : STD_LOGIC;
    SIGNAL S712 : STD_LOGIC;
    SIGNAL S713 : STD_LOGIC;
    SIGNAL S714 : STD_LOGIC;
    SIGNAL S715 : STD_LOGIC;
    SIGNAL S716 : STD_LOGIC;
    SIGNAL S717 : STD_LOGIC;
    SIGNAL S718 : STD_LOGIC;
    SIGNAL S719 : STD_LOGIC;
    SIGNAL S720 : STD_LOGIC;
    SIGNAL S721 : STD_LOGIC;
    SIGNAL S722 : STD_LOGIC;
    SIGNAL S723 : STD_LOGIC;
    SIGNAL S724 : STD_LOGIC;
    SIGNAL S725 : STD_LOGIC;
    SIGNAL S726 : STD_LOGIC;
    SIGNAL S727 : STD_LOGIC;
    SIGNAL S728 : STD_LOGIC;
    SIGNAL S729 : STD_LOGIC;
    SIGNAL S730 : STD_LOGIC;
    SIGNAL S731 : STD_LOGIC;
    SIGNAL S732 : STD_LOGIC;
    SIGNAL S733 : STD_LOGIC;
    SIGNAL S734 : STD_LOGIC;
    SIGNAL S735 : STD_LOGIC;
    SIGNAL S736 : STD_LOGIC;
    SIGNAL S737 : STD_LOGIC;
    SIGNAL S738 : STD_LOGIC;
    SIGNAL S739 : STD_LOGIC;
    SIGNAL S740 : STD_LOGIC;
    SIGNAL S741 : STD_LOGIC;
    SIGNAL S742 : STD_LOGIC;
    SIGNAL S743 : STD_LOGIC;
    SIGNAL S744 : STD_LOGIC;
    SIGNAL S745 : STD_LOGIC;
    SIGNAL S746 : STD_LOGIC;
    SIGNAL S747 : STD_LOGIC;
    SIGNAL S748 : STD_LOGIC;
    SIGNAL S749 : STD_LOGIC;
    SIGNAL S750 : STD_LOGIC;
    SIGNAL S751 : STD_LOGIC;
    SIGNAL S752 : STD_LOGIC;
    SIGNAL S753 : STD_LOGIC;
    SIGNAL S754 : STD_LOGIC;
    SIGNAL S755 : STD_LOGIC;
    SIGNAL S756 : STD_LOGIC;
    SIGNAL S757 : STD_LOGIC;
    SIGNAL S758 : STD_LOGIC;
    SIGNAL S759 : STD_LOGIC;
    SIGNAL S760 : STD_LOGIC;
    SIGNAL S761 : STD_LOGIC;
    SIGNAL S762 : STD_LOGIC;
    SIGNAL S763 : STD_LOGIC;
    SIGNAL S764 : STD_LOGIC;
    SIGNAL S765 : STD_LOGIC;
    SIGNAL S766 : STD_LOGIC;
    SIGNAL S767 : STD_LOGIC;
    SIGNAL S768 : STD_LOGIC;
    SIGNAL S769 : STD_LOGIC;
    SIGNAL S770 : STD_LOGIC;
    SIGNAL S771 : STD_LOGIC;
    SIGNAL S772 : STD_LOGIC;
    SIGNAL S773 : STD_LOGIC;
    SIGNAL S774 : STD_LOGIC;
    SIGNAL S775 : STD_LOGIC;
    SIGNAL S776 : STD_LOGIC;
    SIGNAL S777 : STD_LOGIC;
    SIGNAL S778 : STD_LOGIC;
    SIGNAL S779 : STD_LOGIC;
    SIGNAL S780 : STD_LOGIC;
    SIGNAL S781 : STD_LOGIC;
    SIGNAL S782 : STD_LOGIC;
    SIGNAL S783 : STD_LOGIC;
    SIGNAL S784 : STD_LOGIC;
    SIGNAL S785 : STD_LOGIC;
    SIGNAL S786 : STD_LOGIC;
    SIGNAL S787 : STD_LOGIC;
    SIGNAL S788 : STD_LOGIC;
    SIGNAL S789 : STD_LOGIC;
    SIGNAL S790 : STD_LOGIC;
    SIGNAL S791 : STD_LOGIC;
    SIGNAL S792 : STD_LOGIC;
    SIGNAL S793 : STD_LOGIC;

BEGIN
XNOR2_X1_1: ENTITY WORK.XNOR2_X1
    PORT MAP (
        A => S791(72),
        B => S790(72),
        ZN => S303
    );
XNOR2_X1_2: ENTITY WORK.XNOR2_X1
    PORT MAP (
        A => S791(98),
        B => S790(98),
        ZN => S304
    );
XNOR2_X1_3: ENTITY WORK.XNOR2_X1
    PORT MAP (
        A => S791(100),
        B => S790(100),
        ZN => S305
    );
NAND3_X1_1: ENTITY WORK.NAND3_X1
    PORT MAP (
        A1 => S303,
        A2 => S304,
        A3 => S305,
        ZN => S306
    );
XNOR2_X1_4: ENTITY WORK.XNOR2_X1
    PORT MAP (
        A => S791(96),
        B => S790(96),
        ZN => S307
    );
INV_X1_1: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(34),
        ZN => S308
    );
INV_X1_2: ENTITY WORK.INV_X1
    PORT MAP (
        A => S789,
        ZN => S309
    );
AOI21_X1_1: ENTITY WORK.AOI21_X1
    PORT MAP (
        A => S309,
        B1 => S308,
        B2 => S791(34),
        ZN => S310
    );
XNOR2_X1_5: ENTITY WORK.XNOR2_X1
    PORT MAP (
        A => S791(26),
        B => S790(26),
        ZN => S311
    );
XNOR2_X1_6: ENTITY WORK.XNOR2_X1
    PORT MAP (
        A => S791(28),
        B => S790(28),
        ZN => S312
    );
NAND4_X1_1: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S311,
        A2 => S312,
        A3 => S307,
        A4 => S310,
        ZN => S313
    );
INV_X1_3: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(56),
        ZN => S314
    );
INV_X1_4: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(66),
        ZN => S315
    );
AOI22_X1_1: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S314,
        A2 => S790(56),
        B1 => S315,
        B2 => S791(66),
        ZN => S316
    );
XNOR2_X1_7: ENTITY WORK.XNOR2_X1
    PORT MAP (
        A => S791(36),
        B => S790(36),
        ZN => S317
    );
INV_X1_5: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(34),
        ZN => S318
    );
INV_X1_6: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(54),
        ZN => S319
    );
AOI22_X1_2: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S318,
        A2 => S790(34),
        B1 => S319,
        B2 => S791(54),
        ZN => S320
    );
INV_X1_7: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(54),
        ZN => S321
    );
INV_X1_8: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(56),
        ZN => S322
    );
AOI22_X1_3: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S321,
        A2 => S790(54),
        B1 => S322,
        B2 => S791(56),
        ZN => S323
    );
NAND4_X1_2: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S323,
        A2 => S320,
        A3 => S317,
        A4 => S316,
        ZN => S324
    );
NOR3_X1_1: ENTITY WORK.NOR3_X1
    PORT MAP (
        A1 => S324,
        A2 => S313,
        A3 => S306,
        ZN => S325
    );
INV_X1_9: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(60),
        ZN => S326
    );
INV_X1_10: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(64),
        ZN => S327
    );
AOI22_X1_4: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S327,
        A2 => S790(64),
        B1 => S326,
        B2 => S791(60),
        ZN => S328
    );
INV_X1_11: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(58),
        ZN => S329
    );
INV_X1_12: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(60),
        ZN => S330
    );
AOI22_X1_5: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S330,
        A2 => S790(60),
        B1 => S329,
        B2 => S791(58),
        ZN => S331
    );
INV_X1_13: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(74),
        ZN => S332
    );
INV_X1_14: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(76),
        ZN => S333
    );
AOI22_X1_6: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S333,
        A2 => S790(76),
        B1 => S332,
        B2 => S791(74),
        ZN => S334
    );
INV_X1_15: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(64),
        ZN => S335
    );
INV_X1_16: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(74),
        ZN => S336
    );
AOI22_X1_7: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S336,
        A2 => S790(74),
        B1 => S335,
        B2 => S791(64),
        ZN => S337
    );
AND4_X1_1: ENTITY WORK.AND4_X1
    PORT MAP (
        A1 => S328,
        A2 => S334,
        A3 => S337,
        A4 => S331,
        ZN => S338
    );
INV_X1_17: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(82),
        ZN => S339
    );
NAND2_X1_1: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S339,
        A2 => S790(82),
        ZN => S340
    );
INV_X1_18: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(8),
        ZN => S341
    );
NAND2_X1_2: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S341,
        A2 => S791(8),
        ZN => S342
    );
INV_X1_19: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(8),
        ZN => S343
    );
NAND2_X1_3: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S343,
        A2 => S790(8),
        ZN => S344
    );
INV_X1_20: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(12),
        ZN => S345
    );
NAND2_X1_4: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S345,
        A2 => S791(12),
        ZN => S346
    );
NAND4_X1_3: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S344,
        A2 => S346,
        A3 => S340,
        A4 => S342,
        ZN => S347
    );
INV_X1_21: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(58),
        ZN => S348
    );
NAND2_X1_5: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S348,
        A2 => S790(58),
        ZN => S349
    );
INV_X1_22: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(62),
        ZN => S350
    );
NAND2_X1_6: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S350,
        A2 => S791(62),
        ZN => S351
    );
INV_X1_23: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(62),
        ZN => S352
    );
NAND2_X1_7: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S352,
        A2 => S790(62),
        ZN => S353
    );
INV_X1_24: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(82),
        ZN => S354
    );
NAND2_X1_8: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S354,
        A2 => S791(82),
        ZN => S355
    );
NAND4_X1_4: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S353,
        A2 => S355,
        A3 => S349,
        A4 => S351,
        ZN => S356
    );
NOR2_X1_1: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S347,
        A2 => S356,
        ZN => S357
    );
INV_X1_25: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(32),
        ZN => S358
    );
NAND2_X1_9: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S358,
        A2 => S790(32),
        ZN => S359
    );
INV_X1_26: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(22),
        ZN => S360
    );
NAND2_X1_10: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S360,
        A2 => S791(22),
        ZN => S361
    );
INV_X1_27: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(22),
        ZN => S362
    );
NAND2_X1_11: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S362,
        A2 => S790(22),
        ZN => S363
    );
INV_X1_28: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(80),
        ZN => S364
    );
NAND2_X1_12: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S364,
        A2 => S791(80),
        ZN => S365
    );
NAND4_X1_5: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S363,
        A2 => S365,
        A3 => S359,
        A4 => S361,
        ZN => S366
    );
INV_X1_29: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(32),
        ZN => S367
    );
NAND2_X1_13: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S367,
        A2 => S791(32),
        ZN => S368
    );
INV_X1_30: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(66),
        ZN => S369
    );
NAND2_X1_14: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S369,
        A2 => S790(66),
        ZN => S370
    );
AND2_X1_1: ENTITY WORK.AND2_X1
    PORT MAP (
        A1 => S790(68),
        A2 => S791(68),
        ZN => S371
    );
NOR2_X1_2: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S791(68),
        A2 => S790(68),
        ZN => S372
    );
OAI211_X1_1: ENTITY WORK.OAI211_X1
    PORT MAP (
        A => S370,
        B => S368,
        C1 => S371,
        C2 => S372,
        ZN => S373
    );
NOR2_X1_3: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S366,
        A2 => S373,
        ZN => S374
    );
INV_X1_31: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(70),
        ZN => S375
    );
NAND2_X1_15: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S375,
        A2 => S790(70),
        ZN => S376
    );
INV_X1_32: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(84),
        ZN => S377
    );
NAND2_X1_16: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S377,
        A2 => S791(84),
        ZN => S378
    );
INV_X1_33: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(84),
        ZN => S379
    );
NAND2_X1_17: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S379,
        A2 => S790(84),
        ZN => S380
    );
INV_X1_34: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(76),
        ZN => S381
    );
NAND2_X1_18: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S381,
        A2 => S791(76),
        ZN => S382
    );
NAND4_X1_6: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S380,
        A2 => S382,
        A3 => S376,
        A4 => S378,
        ZN => S383
    );
INV_X1_35: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(80),
        ZN => S384
    );
NAND2_X1_19: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S384,
        A2 => S790(80),
        ZN => S385
    );
INV_X1_36: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(78),
        ZN => S386
    );
NAND2_X1_20: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S386,
        A2 => S791(78),
        ZN => S387
    );
INV_X1_37: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(78),
        ZN => S388
    );
NAND2_X1_21: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S388,
        A2 => S790(78),
        ZN => S389
    );
INV_X1_38: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(70),
        ZN => S390
    );
NAND2_X1_22: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S390,
        A2 => S791(70),
        ZN => S391
    );
NAND4_X1_7: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S389,
        A2 => S391,
        A3 => S385,
        A4 => S387,
        ZN => S392
    );
NOR2_X1_4: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S383,
        A2 => S392,
        ZN => S393
    );
AND4_X1_2: ENTITY WORK.AND4_X1
    PORT MAP (
        A1 => S338,
        A2 => S393,
        A3 => S357,
        A4 => S374,
        ZN => S394
    );
INV_X1_39: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(59),
        ZN => S395
    );
INV_X1_40: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(75),
        ZN => S396
    );
OAI22_X1_1: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S395,
        A2 => S791(59),
        B1 => S396,
        B2 => S790(75),
        ZN => S397
    );
INV_X1_41: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(63),
        ZN => S398
    );
AND2_X1_2: ENTITY WORK.AND2_X1
    PORT MAP (
        A1 => S398,
        A2 => S790(63),
        ZN => S399
    );
NOR2_X1_5: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S398,
        A2 => S790(63),
        ZN => S400
    );
NOR3_X1_2: ENTITY WORK.NOR3_X1
    PORT MAP (
        A1 => S397,
        A2 => S399,
        A3 => S400,
        ZN => S401
    );
INV_X1_42: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(73),
        ZN => S402
    );
INV_X1_43: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(83),
        ZN => S403
    );
AOI22_X1_8: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S402,
        A2 => S790(73),
        B1 => S403,
        B2 => S791(83),
        ZN => S404
    );
INV_X1_44: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(69),
        ZN => S405
    );
AOI22_X1_9: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S790(69),
        A2 => S405,
        B1 => S396,
        B2 => S790(75),
        ZN => S406
    );
AND2_X1_3: ENTITY WORK.AND2_X1
    PORT MAP (
        A1 => S406,
        A2 => S404,
        ZN => S407
    );
INV_X1_45: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(57),
        ZN => S408
    );
INV_X1_46: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(65),
        ZN => S409
    );
OAI22_X1_2: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S408,
        A2 => S791(57),
        B1 => S409,
        B2 => S790(65),
        ZN => S410
    );
INV_X1_47: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(61),
        ZN => S411
    );
OAI22_X1_3: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S411,
        A2 => S790(61),
        B1 => S403,
        B2 => S791(83),
        ZN => S412
    );
NOR2_X1_6: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S410,
        A2 => S412,
        ZN => S413
    );
INV_X1_48: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(71),
        ZN => S414
    );
INV_X1_49: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(77),
        ZN => S415
    );
AOI22_X1_10: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S791(77),
        A2 => S415,
        B1 => S414,
        B2 => S791(71),
        ZN => S416
    );
INV_X1_50: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(31),
        ZN => S417
    );
AOI22_X1_11: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S790(31),
        A2 => S417,
        B1 => S411,
        B2 => S790(61),
        ZN => S418
    );
AND2_X1_4: ENTITY WORK.AND2_X1
    PORT MAP (
        A1 => S418,
        A2 => S416,
        ZN => S419
    );
NAND4_X1_8: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S419,
        A2 => S407,
        A3 => S401,
        A4 => S413,
        ZN => S420
    );
INV_X1_51: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(42),
        ZN => S421
    );
INV_X1_52: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(46),
        ZN => S422
    );
OAI22_X1_4: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S421,
        A2 => S790(42),
        B1 => S422,
        B2 => S791(46),
        ZN => S423
    );
INV_X1_53: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(40),
        ZN => S424
    );
INV_X1_54: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(42),
        ZN => S425
    );
OAI22_X1_5: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S424,
        A2 => S790(40),
        B1 => S425,
        B2 => S791(42),
        ZN => S426
    );
NOR2_X1_7: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S423,
        A2 => S426,
        ZN => S427
    );
INV_X1_55: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(10),
        ZN => S428
    );
OAI22_X1_6: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S428,
        A2 => S790(10),
        B1 => S345,
        B2 => S791(12),
        ZN => S429
    );
INV_X1_56: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(10),
        ZN => S430
    );
INV_X1_57: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(46),
        ZN => S431
    );
OAI22_X1_7: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S430,
        A2 => S791(10),
        B1 => S431,
        B2 => S790(46),
        ZN => S432
    );
NOR2_X1_8: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S429,
        A2 => S432,
        ZN => S433
    );
INV_X1_58: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(6),
        ZN => S434
    );
AOI22_X1_12: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S434,
        A2 => S790(6),
        B1 => S395,
        B2 => S791(59),
        ZN => S435
    );
INV_X1_59: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(41),
        ZN => S436
    );
INV_X1_60: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(81),
        ZN => S437
    );
AOI22_X1_13: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S437,
        A2 => S790(81),
        B1 => S436,
        B2 => S791(41),
        ZN => S438
    );
AND2_X1_5: ENTITY WORK.AND2_X1
    PORT MAP (
        A1 => S438,
        A2 => S435,
        ZN => S439
    );
INV_X1_61: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(40),
        ZN => S440
    );
INV_X1_62: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(44),
        ZN => S441
    );
OAI22_X1_8: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S440,
        A2 => S791(40),
        B1 => S441,
        B2 => S790(44),
        ZN => S442
    );
INV_X1_63: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(44),
        ZN => S443
    );
OAI22_X1_9: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S434,
        A2 => S790(6),
        B1 => S443,
        B2 => S791(44),
        ZN => S444
    );
NOR2_X1_9: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S442,
        A2 => S444,
        ZN => S445
    );
NAND4_X1_9: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S439,
        A2 => S445,
        A3 => S427,
        A4 => S433,
        ZN => S446
    );
NOR2_X1_10: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S420,
        A2 => S446,
        ZN => S447
    );
NAND3_X1_2: ENTITY WORK.NAND3_X1
    PORT MAP (
        A1 => S447,
        A2 => S394,
        A3 => S325,
        ZN => S448
    );
INV_X1_64: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(127),
        ZN => S449
    );
INV_X1_65: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(125),
        ZN => S450
    );
AOI22_X1_14: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S450,
        A2 => S790(125),
        B1 => S449,
        B2 => S791(127),
        ZN => S451
    );
OAI21_X1_1: ENTITY WORK.OAI21_X1
    PORT MAP (
        A => S451,
        B1 => S791(127),
        B2 => S449,
        ZN => S452
    );
INV_X1_66: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(122),
        ZN => S453
    );
INV_X1_67: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(126),
        ZN => S454
    );
NAND2_X1_23: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S454,
        A2 => S790(126),
        ZN => S455
    );
INV_X1_68: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(123),
        ZN => S456
    );
AOI22_X1_15: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S790(122),
        A2 => S453,
        B1 => S456,
        B2 => S790(123),
        ZN => S457
    );
OAI211_X1_2: ENTITY WORK.OAI211_X1
    PORT MAP (
        A => S457,
        B => S455,
        C1 => S790(122),
        C2 => S453,
        ZN => S458
    );
INV_X1_69: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(117),
        ZN => S459
    );
INV_X1_70: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(109),
        ZN => S460
    );
AOI22_X1_16: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S459,
        A2 => S790(117),
        B1 => S460,
        B2 => S791(109),
        ZN => S461
    );
OAI221_X1_1: ENTITY WORK.OAI221_X1
    PORT MAP (
        A => S461,
        B1 => S454,
        B2 => S790(126),
        C1 => S790(117),
        C2 => S459,
        ZN => S462
    );
NOR3_X1_3: ENTITY WORK.NOR3_X1
    PORT MAP (
        A1 => S462,
        A2 => S458,
        A3 => S452,
        ZN => S463
    );
INV_X1_71: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(16),
        ZN => S464
    );
INV_X1_72: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(18),
        ZN => S465
    );
OAI22_X1_10: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S464,
        A2 => S790(16),
        B1 => S465,
        B2 => S791(18),
        ZN => S466
    );
INV_X1_73: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(14),
        ZN => S467
    );
INV_X1_74: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(16),
        ZN => S468
    );
OAI22_X1_11: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S467,
        A2 => S790(14),
        B1 => S468,
        B2 => S791(16),
        ZN => S469
    );
INV_X1_75: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(106),
        ZN => S470
    );
INV_X1_76: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(124),
        ZN => S471
    );
AOI22_X1_17: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S471,
        A2 => S790(124),
        B1 => S470,
        B2 => S791(106),
        ZN => S472
    );
INV_X1_77: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(106),
        ZN => S473
    );
AOI22_X1_18: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S473,
        A2 => S790(106),
        B1 => S465,
        B2 => S791(18),
        ZN => S474
    );
NAND2_X1_24: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S472,
        A2 => S474,
        ZN => S475
    );
INV_X1_78: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(115),
        ZN => S476
    );
INV_X1_79: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(121),
        ZN => S477
    );
AOI22_X1_19: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S476,
        A2 => S790(115),
        B1 => S477,
        B2 => S791(121),
        ZN => S478
    );
INV_X1_80: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(105),
        ZN => S479
    );
INV_X1_81: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(113),
        ZN => S480
    );
AOI22_X1_20: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S790(105),
        A2 => S479,
        B1 => S480,
        B2 => S790(113),
        ZN => S481
    );
INV_X1_82: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(4),
        ZN => S482
    );
AOI22_X1_21: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S467,
        A2 => S790(14),
        B1 => S482,
        B2 => S791(4),
        ZN => S483
    );
INV_X1_83: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(4),
        ZN => S484
    );
INV_X1_84: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(115),
        ZN => S485
    );
AOI22_X1_22: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S484,
        A2 => S790(4),
        B1 => S485,
        B2 => S791(115),
        ZN => S486
    );
NAND4_X1_10: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S483,
        A2 => S486,
        A3 => S478,
        A4 => S481,
        ZN => S487
    );
NOR4_X1_1: ENTITY WORK.NOR4_X1
    PORT MAP (
        A1 => S487,
        A2 => S475,
        A3 => S469,
        A4 => S466,
        ZN => S488
    );
INV_X1_85: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(37),
        ZN => S489
    );
INV_X1_86: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(77),
        ZN => S490
    );
AOI22_X1_23: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S490,
        A2 => S790(77),
        B1 => S489,
        B2 => S791(37),
        ZN => S491
    );
INV_X1_87: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(53),
        ZN => S492
    );
INV_X1_88: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(81),
        ZN => S493
    );
AOI22_X1_24: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S492,
        A2 => S790(53),
        B1 => S493,
        B2 => S791(81),
        ZN => S494
    );
INV_X1_89: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(91),
        ZN => S495
    );
INV_X1_90: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(93),
        ZN => S496
    );
AOI22_X1_25: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S495,
        A2 => S790(91),
        B1 => S496,
        B2 => S791(93),
        ZN => S497
    );
INV_X1_91: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(33),
        ZN => S498
    );
INV_X1_92: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(87),
        ZN => S499
    );
AOI22_X1_26: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S790(33),
        A2 => S498,
        B1 => S499,
        B2 => S790(87),
        ZN => S500
    );
NAND4_X1_11: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S497,
        A2 => S500,
        A3 => S491,
        A4 => S494,
        ZN => S501
    );
INV_X1_93: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(110),
        ZN => S502
    );
INV_X1_94: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(116),
        ZN => S503
    );
OAI22_X1_12: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S502,
        A2 => S790(110),
        B1 => S503,
        B2 => S791(116),
        ZN => S504
    );
INV_X1_95: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(110),
        ZN => S505
    );
OAI22_X1_13: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S505,
        A2 => S791(110),
        B1 => S471,
        B2 => S790(124),
        ZN => S506
    );
INV_X1_96: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(55),
        ZN => S507
    );
AOI22_X1_27: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S507,
        A2 => S790(55),
        B1 => S408,
        B2 => S791(57),
        ZN => S508
    );
INV_X1_97: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(67),
        ZN => S509
    );
AOI22_X1_28: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S791(116),
        A2 => S503,
        B1 => S509,
        B2 => S791(67),
        ZN => S510
    );
NAND2_X1_25: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S508,
        A2 => S510,
        ZN => S511
    );
NOR4_X1_2: ENTITY WORK.NOR4_X1
    PORT MAP (
        A1 => S501,
        A2 => S511,
        A3 => S506,
        A4 => S504,
        ZN => S512
    );
NAND3_X1_3: ENTITY WORK.NAND3_X1
    PORT MAP (
        A1 => S488,
        A2 => S512,
        A3 => S463,
        ZN => S513
    );
INV_X1_98: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(94),
        ZN => S514
    );
NAND2_X1_26: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S514,
        A2 => S791(94),
        ZN => S515
    );
INV_X1_99: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(24),
        ZN => S516
    );
NAND2_X1_27: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S516,
        A2 => S790(24),
        ZN => S517
    );
INV_X1_100: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(24),
        ZN => S518
    );
NAND2_X1_28: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S518,
        A2 => S791(24),
        ZN => S519
    );
INV_X1_101: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(33),
        ZN => S520
    );
NAND2_X1_29: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S520,
        A2 => S791(33),
        ZN => S521
    );
NAND4_X1_12: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S519,
        A2 => S521,
        A3 => S515,
        A4 => S517,
        ZN => S522
    );
INV_X1_102: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(90),
        ZN => S523
    );
NAND2_X1_30: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S523,
        A2 => S790(90),
        ZN => S524
    );
INV_X1_103: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(94),
        ZN => S525
    );
NAND2_X1_31: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S525,
        A2 => S790(94),
        ZN => S526
    );
INV_X1_104: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(88),
        ZN => S527
    );
NAND2_X1_32: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S527,
        A2 => S791(88),
        ZN => S528
    );
INV_X1_105: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(92),
        ZN => S529
    );
NAND2_X1_33: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S529,
        A2 => S790(92),
        ZN => S530
    );
NAND4_X1_13: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S528,
        A2 => S530,
        A3 => S524,
        A4 => S526,
        ZN => S531
    );
NOR2_X1_11: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S522,
        A2 => S531,
        ZN => S532
    );
INV_X1_106: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(27),
        ZN => S533
    );
INV_X1_107: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(29),
        ZN => S534
    );
AOI22_X1_29: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S533,
        A2 => S790(27),
        B1 => S534,
        B2 => S791(29),
        ZN => S535
    );
INV_X1_108: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(51),
        ZN => S536
    );
INV_X1_109: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(95),
        ZN => S537
    );
AOI22_X1_30: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S790(51),
        A2 => S536,
        B1 => S537,
        B2 => S790(95),
        ZN => S538
    );
INV_X1_110: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(21),
        ZN => S539
    );
INV_X1_111: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(25),
        ZN => S540
    );
AOI22_X1_31: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S790(21),
        A2 => S539,
        B1 => S540,
        B2 => S790(25),
        ZN => S541
    );
INV_X1_112: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(23),
        ZN => S542
    );
INV_X1_113: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(27),
        ZN => S543
    );
AOI22_X1_32: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S791(27),
        A2 => S543,
        B1 => S542,
        B2 => S791(23),
        ZN => S544
    );
AND4_X1_3: ENTITY WORK.AND4_X1
    PORT MAP (
        A1 => S535,
        A2 => S541,
        A3 => S544,
        A4 => S538,
        ZN => S545
    );
INV_X1_114: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(92),
        ZN => S546
    );
NAND2_X1_34: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S546,
        A2 => S791(92),
        ZN => S547
    );
INV_X1_115: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(52),
        ZN => S548
    );
NAND2_X1_35: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S548,
        A2 => S790(52),
        ZN => S549
    );
INV_X1_116: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(50),
        ZN => S550
    );
NAND2_X1_36: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S550,
        A2 => S791(50),
        ZN => S551
    );
INV_X1_117: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(48),
        ZN => S552
    );
NAND2_X1_37: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S552,
        A2 => S791(48),
        ZN => S553
    );
NAND4_X1_14: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S551,
        A2 => S553,
        A3 => S547,
        A4 => S549,
        ZN => S554
    );
INV_X1_118: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(120),
        ZN => S555
    );
NAND2_X1_38: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S555,
        A2 => S790(120),
        ZN => S556
    );
INV_X1_119: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(118),
        ZN => S557
    );
NAND2_X1_39: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S557,
        A2 => S791(118),
        ZN => S558
    );
INV_X1_120: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(118),
        ZN => S559
    );
NAND2_X1_40: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S559,
        A2 => S790(118),
        ZN => S560
    );
INV_X1_121: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(88),
        ZN => S561
    );
NAND2_X1_41: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S561,
        A2 => S790(88),
        ZN => S562
    );
NAND4_X1_15: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S560,
        A2 => S562,
        A3 => S556,
        A4 => S558,
        ZN => S563
    );
NOR2_X1_12: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S554,
        A2 => S563,
        ZN => S564
    );
AND2_X1_6: ENTITY WORK.AND2_X1
    PORT MAP (
        A1 => S790(86),
        A2 => S791(86),
        ZN => S565
    );
NOR2_X1_13: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S791(86),
        A2 => S790(86),
        ZN => S566
    );
INV_X1_122: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(30),
        ZN => S567
    );
NAND2_X1_42: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S567,
        A2 => S791(30),
        ZN => S568
    );
INV_X1_123: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(90),
        ZN => S569
    );
NAND2_X1_43: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S569,
        A2 => S791(90),
        ZN => S570
    );
OAI211_X1_3: ENTITY WORK.OAI211_X1
    PORT MAP (
        A => S570,
        B => S568,
        C1 => S565,
        C2 => S566,
        ZN => S571
    );
INV_X1_124: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(48),
        ZN => S572
    );
NAND2_X1_44: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S572,
        A2 => S790(48),
        ZN => S573
    );
INV_X1_125: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(30),
        ZN => S574
    );
NAND2_X1_45: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S574,
        A2 => S790(30),
        ZN => S575
    );
INV_X1_126: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(52),
        ZN => S576
    );
NAND2_X1_46: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S576,
        A2 => S791(52),
        ZN => S577
    );
INV_X1_127: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(50),
        ZN => S578
    );
NAND2_X1_47: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S578,
        A2 => S790(50),
        ZN => S579
    );
NAND4_X1_16: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S577,
        A2 => S579,
        A3 => S573,
        A4 => S575,
        ZN => S580
    );
NOR2_X1_14: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S580,
        A2 => S571,
        ZN => S581
    );
AND4_X1_4: ENTITY WORK.AND4_X1
    PORT MAP (
        A1 => S545,
        A2 => S532,
        A3 => S564,
        A4 => S581,
        ZN => S582
    );
INV_X1_128: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(15),
        ZN => S583
    );
INV_X1_129: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(19),
        ZN => S584
    );
AOI22_X1_33: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S584,
        A2 => S790(19),
        B1 => S583,
        B2 => S791(15),
        ZN => S585
    );
INV_X1_130: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(7),
        ZN => S586
    );
INV_X1_131: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(49),
        ZN => S587
    );
AOI22_X1_34: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S790(7),
        A2 => S586,
        B1 => S587,
        B2 => S790(49),
        ZN => S588
    );
AND2_X1_7: ENTITY WORK.AND2_X1
    PORT MAP (
        A1 => S588,
        A2 => S585,
        ZN => S589
    );
XOR2_X1_1: ENTITY WORK.XOR2_X1
    PORT MAP (
        A => S791(1),
        B => S790(1),
        Z => S590
    );
INV_X1_132: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(111),
        ZN => S591
    );
OAI22_X1_14: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S591,
        A2 => S791(111),
        B1 => S480,
        B2 => S790(113),
        ZN => S592
    );
NOR2_X1_15: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S590,
        A2 => S592,
        ZN => S593
    );
INV_X1_133: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(87),
        ZN => S594
    );
INV_X1_134: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(97),
        ZN => S595
    );
AOI22_X1_35: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S791(97),
        A2 => S595,
        B1 => S594,
        B2 => S791(87),
        ZN => S596
    );
INV_X1_135: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(89),
        ZN => S597
    );
INV_X1_136: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(101),
        ZN => S598
    );
AOI22_X1_36: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S597,
        A2 => S790(89),
        B1 => S598,
        B2 => S791(101),
        ZN => S599
    );
AND2_X1_8: ENTITY WORK.AND2_X1
    PORT MAP (
        A1 => S599,
        A2 => S596,
        ZN => S600
    );
INV_X1_137: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(11),
        ZN => S601
    );
INV_X1_138: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(45),
        ZN => S602
    );
OAI22_X1_15: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S791(11),
        A2 => S601,
        B1 => S602,
        B2 => S791(45),
        ZN => S603
    );
OAI22_X1_16: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S492,
        A2 => S790(53),
        B1 => S595,
        B2 => S791(97),
        ZN => S604
    );
NOR2_X1_16: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S603,
        A2 => S604,
        ZN => S605
    );
NAND4_X1_17: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S593,
        A2 => S589,
        A3 => S600,
        A4 => S605,
        ZN => S606
    );
INV_X1_139: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(9),
        ZN => S607
    );
NAND2_X1_48: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S607,
        A2 => S790(9),
        ZN => S608
    );
OR2_X1_1: ENTITY WORK.OR2_X1
    PORT MAP (
        A1 => S607,
        A2 => S790(9),
        ZN => S609
    );
INV_X1_140: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(13),
        ZN => S610
    );
INV_X1_141: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(17),
        ZN => S611
    );
AOI22_X1_37: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S610,
        A2 => S790(13),
        B1 => S611,
        B2 => S791(17),
        ZN => S612
    );
AND3_X1_1: ENTITY WORK.AND3_X1
    PORT MAP (
        A1 => S612,
        A2 => S609,
        A3 => S608,
        ZN => S613
    );
INV_X1_142: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(11),
        ZN => S614
    );
OAI22_X1_17: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S790(7),
        A2 => S586,
        B1 => S614,
        B2 => S790(11),
        ZN => S615
    );
OAI22_X1_18: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S790(13),
        A2 => S610,
        B1 => S536,
        B2 => S790(51),
        ZN => S616
    );
NOR2_X1_17: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S615,
        A2 => S616,
        ZN => S617
    );
OAI22_X1_19: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S542,
        A2 => S791(23),
        B1 => S417,
        B2 => S790(31),
        ZN => S618
    );
INV_X1_143: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(3),
        ZN => S619
    );
INV_X1_144: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(5),
        ZN => S620
    );
OAI22_X1_20: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S790(3),
        A2 => S619,
        B1 => S620,
        B2 => S790(5),
        ZN => S621
    );
NOR2_X1_18: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S618,
        A2 => S621,
        ZN => S622
    );
INV_X1_145: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(45),
        ZN => S623
    );
OAI22_X1_21: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S436,
        A2 => S791(41),
        B1 => S623,
        B2 => S790(45),
        ZN => S624
    );
INV_X1_146: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(47),
        ZN => S625
    );
OAI22_X1_22: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S540,
        A2 => S790(25),
        B1 => S625,
        B2 => S791(47),
        ZN => S626
    );
NOR2_X1_19: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S624,
        A2 => S626,
        ZN => S627
    );
NAND4_X1_18: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S613,
        A2 => S617,
        A3 => S622,
        A4 => S627,
        ZN => S628
    );
NOR2_X1_20: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S606,
        A2 => S628,
        ZN => S629
    );
INV_X1_147: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(99),
        ZN => S630
    );
OAI22_X1_23: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S790(95),
        A2 => S537,
        B1 => S630,
        B2 => S790(99),
        ZN => S631
    );
INV_X1_148: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(85),
        ZN => S632
    );
INV_X1_149: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(99),
        ZN => S633
    );
OAI22_X1_24: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S791(85),
        A2 => S632,
        B1 => S633,
        B2 => S791(99),
        ZN => S634
    );
NOR2_X1_21: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S631,
        A2 => S634,
        ZN => S635
    );
INV_X1_150: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(103),
        ZN => S636
    );
OAI22_X1_25: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S636,
        A2 => S791(103),
        B1 => S479,
        B2 => S790(105),
        ZN => S637
    );
OAI22_X1_26: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S611,
        A2 => S791(17),
        B1 => S539,
        B2 => S790(21),
        ZN => S638
    );
NOR2_X1_22: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S637,
        A2 => S638,
        ZN => S639
    );
INV_X1_151: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(79),
        ZN => S640
    );
OAI22_X1_27: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S790(55),
        A2 => S507,
        B1 => S640,
        B2 => S790(79),
        ZN => S641
    );
INV_X1_152: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(79),
        ZN => S642
    );
OAI22_X1_28: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S791(71),
        A2 => S414,
        B1 => S642,
        B2 => S791(79),
        ZN => S643
    );
NOR2_X1_23: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S641,
        A2 => S643,
        ZN => S644
    );
OAI22_X1_29: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S509,
        A2 => S791(67),
        B1 => S495,
        B2 => S790(91),
        ZN => S645
    );
OAI22_X1_30: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S597,
        A2 => S790(89),
        B1 => S496,
        B2 => S791(93),
        ZN => S646
    );
NOR2_X1_24: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S645,
        A2 => S646,
        ZN => S647
    );
NAND4_X1_19: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S644,
        A2 => S647,
        A3 => S635,
        A4 => S639,
        ZN => S648
    );
INV_X1_153: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(43),
        ZN => S649
    );
OAI22_X1_31: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S790(43),
        A2 => S649,
        B1 => S587,
        B2 => S790(49),
        ZN => S650
    );
INV_X1_154: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(43),
        ZN => S651
    );
OAI22_X1_32: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S791(37),
        A2 => S489,
        B1 => S651,
        B2 => S791(43),
        ZN => S652
    );
NOR2_X1_25: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S650,
        A2 => S652,
        ZN => S653
    );
NAND2_X1_49: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S632,
        A2 => S791(85),
        ZN => S654
    );
NAND2_X1_50: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S625,
        A2 => S791(47),
        ZN => S655
    );
INV_X1_155: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(39),
        ZN => S656
    );
NAND2_X1_51: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S656,
        A2 => S790(39),
        ZN => S657
    );
NAND2_X1_52: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S620,
        A2 => S790(5),
        ZN => S658
    );
AND4_X1_5: ENTITY WORK.AND4_X1
    PORT MAP (
        A1 => S654,
        A2 => S657,
        A3 => S658,
        A4 => S655,
        ZN => S659
    );
INV_X1_156: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(3),
        ZN => S660
    );
OAI22_X1_33: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S660,
        A2 => S791(3),
        B1 => S584,
        B2 => S790(19),
        ZN => S661
    );
INV_X1_157: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(0),
        ZN => S662
    );
AND2_X1_9: ENTITY WORK.AND2_X1
    PORT MAP (
        A1 => S662,
        A2 => S791(0),
        ZN => S663
    );
NOR2_X1_26: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S662,
        A2 => S791(0),
        ZN => S664
    );
NOR3_X1_4: ENTITY WORK.NOR3_X1
    PORT MAP (
        A1 => S661,
        A2 => S663,
        A3 => S664,
        ZN => S665
    );
OAI22_X1_34: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S583,
        A2 => S791(15),
        B1 => S656,
        B2 => S790(39),
        ZN => S666
    );
INV_X1_158: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(35),
        ZN => S667
    );
OAI22_X1_35: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S534,
        A2 => S791(29),
        B1 => S667,
        B2 => S790(35),
        ZN => S668
    );
NOR2_X1_27: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S666,
        A2 => S668,
        ZN => S669
    );
NAND4_X1_20: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S665,
        A2 => S669,
        A3 => S659,
        A4 => S653,
        ZN => S670
    );
NOR2_X1_28: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S648,
        A2 => S670,
        ZN => S671
    );
INV_X1_159: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(103),
        ZN => S672
    );
OAI22_X1_36: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S598,
        A2 => S791(101),
        B1 => S672,
        B2 => S790(103),
        ZN => S673
    );
INV_X1_160: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(111),
        ZN => S674
    );
OAI22_X1_37: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S460,
        A2 => S791(109),
        B1 => S674,
        B2 => S790(111),
        ZN => S675
    );
NOR2_X1_29: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S673,
        A2 => S675,
        ZN => S676
    );
NAND2_X1_53: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S791(112),
        A2 => S790(112),
        ZN => S677
    );
OR2_X1_2: ENTITY WORK.OR2_X1
    PORT MAP (
        A1 => S791(112),
        A2 => S790(112),
        ZN => S678
    );
NAND2_X1_54: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S791(2),
        A2 => S790(2),
        ZN => S679
    );
OR2_X1_3: ENTITY WORK.OR2_X1
    PORT MAP (
        A1 => S791(2),
        A2 => S790(2),
        ZN => S680
    );
AOI22_X1_38: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S679,
        A2 => S680,
        B1 => S678,
        B2 => S677,
        ZN => S681
    );
OAI22_X1_38: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S477,
        A2 => S791(121),
        B1 => S456,
        B2 => S790(123),
        ZN => S682
    );
OAI22_X1_39: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S790(120),
        A2 => S555,
        B1 => S450,
        B2 => S790(125),
        ZN => S683
    );
NOR2_X1_30: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S682,
        A2 => S683,
        ZN => S684
    );
INV_X1_161: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(107),
        ZN => S685
    );
NAND2_X1_55: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S685,
        A2 => S791(107),
        ZN => S686
    );
INV_X1_162: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(107),
        ZN => S687
    );
NAND2_X1_56: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S687,
        A2 => S790(107),
        ZN => S688
    );
INV_X1_163: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(119),
        ZN => S689
    );
NAND2_X1_57: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S689,
        A2 => S791(119),
        ZN => S690
    );
INV_X1_164: ENTITY WORK.INV_X1
    PORT MAP (
        A => S791(119),
        ZN => S691
    );
NAND2_X1_58: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S691,
        A2 => S790(119),
        ZN => S692
    );
AND4_X1_6: ENTITY WORK.AND4_X1
    PORT MAP (
        A1 => S686,
        A2 => S690,
        A3 => S692,
        A4 => S688,
        ZN => S693
    );
NAND4_X1_21: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S684,
        A2 => S693,
        A3 => S676,
        A4 => S681,
        ZN => S694
    );
NAND2_X1_59: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S791(114),
        A2 => S790(114),
        ZN => S695
    );
OR2_X1_4: ENTITY WORK.OR2_X1
    PORT MAP (
        A1 => S791(114),
        A2 => S790(114),
        ZN => S696
    );
NAND2_X1_60: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S791(104),
        A2 => S790(104),
        ZN => S697
    );
OR2_X1_5: ENTITY WORK.OR2_X1
    PORT MAP (
        A1 => S791(104),
        A2 => S790(104),
        ZN => S698
    );
AOI22_X1_39: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S697,
        A2 => S698,
        B1 => S696,
        B2 => S695,
        ZN => S699
    );
INV_X1_165: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(35),
        ZN => S700
    );
OAI22_X1_40: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S700,
        A2 => S791(35),
        B1 => S402,
        B2 => S790(73),
        ZN => S701
    );
INV_X1_166: ENTITY WORK.INV_X1
    PORT MAP (
        A => S790(65),
        ZN => S702
    );
OAI22_X1_41: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S702,
        A2 => S791(65),
        B1 => S405,
        B2 => S790(69),
        ZN => S703
    );
NOR2_X1_31: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S701,
        A2 => S703,
        ZN => S704
    );
NAND2_X1_61: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S791(38),
        A2 => S790(38),
        ZN => S705
    );
OR2_X1_6: ENTITY WORK.OR2_X1
    PORT MAP (
        A1 => S791(38),
        A2 => S790(38),
        ZN => S706
    );
NAND2_X1_62: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S791(20),
        A2 => S790(20),
        ZN => S707
    );
OR2_X1_7: ENTITY WORK.OR2_X1
    PORT MAP (
        A1 => S791(20),
        A2 => S790(20),
        ZN => S708
    );
AOI22_X1_40: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S707,
        A2 => S708,
        B1 => S706,
        B2 => S705,
        ZN => S709
    );
NAND2_X1_63: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S791(108),
        A2 => S790(108),
        ZN => S710
    );
OR2_X1_8: ENTITY WORK.OR2_X1
    PORT MAP (
        A1 => S791(108),
        A2 => S790(108),
        ZN => S711
    );
NAND2_X1_64: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S791(102),
        A2 => S790(102),
        ZN => S712
    );
OR2_X1_9: ENTITY WORK.OR2_X1
    PORT MAP (
        A1 => S791(102),
        A2 => S790(102),
        ZN => S713
    );
AOI22_X1_41: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S712,
        A2 => S713,
        B1 => S711,
        B2 => S710,
        ZN => S714
    );
NAND4_X1_22: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S704,
        A2 => S699,
        A3 => S709,
        A4 => S714,
        ZN => S715
    );
NOR2_X1_32: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S694,
        A2 => S715,
        ZN => S716
    );
NAND4_X1_23: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S629,
        A2 => S671,
        A3 => S582,
        A4 => S716,
        ZN => S717
    );
NOR3_X1_5: ENTITY WORK.NOR3_X1
    PORT MAP (
        A1 => S717,
        A2 => S448,
        A3 => S513,
        ZN => S788
    );
XNOR2_X1_8: ENTITY WORK.XNOR2_X1
    PORT MAP (
        A => S792(72),
        B => S787(72),
        ZN => S718
    );
XNOR2_X1_9: ENTITY WORK.XNOR2_X1
    PORT MAP (
        A => S792(18),
        B => S787(18),
        ZN => S719
    );
XNOR2_X1_10: ENTITY WORK.XNOR2_X1
    PORT MAP (
        A => S792(20),
        B => S787(20),
        ZN => S720
    );
NAND3_X1_4: ENTITY WORK.NAND3_X1
    PORT MAP (
        A1 => S718,
        A2 => S719,
        A3 => S720,
        ZN => S721
    );
XNOR2_X1_11: ENTITY WORK.XNOR2_X1
    PORT MAP (
        A => S792(70),
        B => S787(70),
        ZN => S722
    );
XNOR2_X1_12: ENTITY WORK.XNOR2_X1
    PORT MAP (
        A => S792(16),
        B => S787(16),
        ZN => S723
    );
XNOR2_X1_13: ENTITY WORK.XNOR2_X1
    PORT MAP (
        A => S792(30),
        B => S787(30),
        ZN => S724
    );
XNOR2_X1_14: ENTITY WORK.XNOR2_X1
    PORT MAP (
        A => S792(36),
        B => S787(36),
        ZN => S725
    );
NAND4_X1_24: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S724,
        A2 => S725,
        A3 => S722,
        A4 => S723,
        ZN => S726
    );
INV_X1_167: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(56),
        ZN => S727
    );
INV_X1_168: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(60),
        ZN => S728
    );
AOI22_X1_42: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S727,
        A2 => S787(56),
        B1 => S728,
        B2 => S792(60),
        ZN => S729
    );
INV_X1_169: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(60),
        ZN => S730
    );
INV_X1_170: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(66),
        ZN => S731
    );
AOI22_X1_43: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S730,
        A2 => S787(60),
        B1 => S731,
        B2 => S792(66),
        ZN => S732
    );
INV_X1_171: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(76),
        ZN => S733
    );
AOI21_X1_2: ENTITY WORK.AOI21_X1
    PORT MAP (
        A => S309,
        B1 => S792(76),
        B2 => S733,
        ZN => S734
    );
INV_X1_172: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(56),
        ZN => S735
    );
INV_X1_173: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(76),
        ZN => S736
    );
AOI22_X1_44: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S736,
        A2 => S787(76),
        B1 => S735,
        B2 => S792(56),
        ZN => S737
    );
NAND4_X1_25: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S737,
        A2 => S732,
        A3 => S729,
        A4 => S734,
        ZN => S738
    );
NOR3_X1_6: ENTITY WORK.NOR3_X1
    PORT MAP (
        A1 => S726,
        A2 => S738,
        A3 => S721,
        ZN => S739
    );
INV_X1_174: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(88),
        ZN => S740
    );
INV_X1_175: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(92),
        ZN => S741
    );
AOI22_X1_45: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S740,
        A2 => S787(88),
        B1 => S741,
        B2 => S792(92),
        ZN => S742
    );
INV_X1_176: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(22),
        ZN => S743
    );
INV_X1_177: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(40),
        ZN => S744
    );
AOI22_X1_46: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S743,
        A2 => S787(22),
        B1 => S744,
        B2 => S792(40),
        ZN => S745
    );
INV_X1_178: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(86),
        ZN => S746
    );
INV_X1_179: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(98),
        ZN => S747
    );
AOI22_X1_47: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S746,
        A2 => S787(86),
        B1 => S747,
        B2 => S792(98),
        ZN => S748
    );
INV_X1_180: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(88),
        ZN => S749
    );
INV_X1_181: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(98),
        ZN => S750
    );
AOI22_X1_48: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S750,
        A2 => S787(98),
        B1 => S749,
        B2 => S792(88),
        ZN => S751
    );
AND4_X1_7: ENTITY WORK.AND4_X1
    PORT MAP (
        A1 => S742,
        A2 => S748,
        A3 => S751,
        A4 => S745,
        ZN => S752
    );
INV_X1_182: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(94),
        ZN => S753
    );
INV_X1_183: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(100),
        ZN => S754
    );
AOI22_X1_49: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S753,
        A2 => S787(94),
        B1 => S754,
        B2 => S792(100),
        ZN => S755
    );
INV_X1_184: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(92),
        ZN => S756
    );
INV_X1_185: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(100),
        ZN => S757
    );
AOI22_X1_50: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S787(92),
        A2 => S756,
        B1 => S757,
        B2 => S787(100),
        ZN => S758
    );
INV_X1_186: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(40),
        ZN => S759
    );
INV_X1_187: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(96),
        ZN => S760
    );
AOI22_X1_51: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S759,
        A2 => S787(40),
        B1 => S760,
        B2 => S792(96),
        ZN => S761
    );
INV_X1_188: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(94),
        ZN => S762
    );
INV_X1_189: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(96),
        ZN => S763
    );
AOI22_X1_52: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S763,
        A2 => S787(96),
        B1 => S762,
        B2 => S792(94),
        ZN => S764
    );
AND4_X1_8: ENTITY WORK.AND4_X1
    PORT MAP (
        A1 => S755,
        A2 => S761,
        A3 => S764,
        A4 => S758,
        ZN => S765
    );
AND2_X1_10: ENTITY WORK.AND2_X1
    PORT MAP (
        A1 => S787(68),
        A2 => S792(68),
        ZN => S766
    );
NOR2_X1_33: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S792(68),
        A2 => S787(68),
        ZN => S767
    );
INV_X1_190: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(74),
        ZN => S768
    );
NAND2_X1_65: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S768,
        A2 => S787(74),
        ZN => S769
    );
INV_X1_191: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(34),
        ZN => S770
    );
NAND2_X1_66: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S770,
        A2 => S792(34),
        ZN => S771
    );
OAI211_X1_4: ENTITY WORK.OAI211_X1
    PORT MAP (
        A => S771,
        B => S769,
        C1 => S766,
        C2 => S767,
        ZN => S772
    );
AND2_X1_11: ENTITY WORK.AND2_X1
    PORT MAP (
        A1 => S787(80),
        A2 => S792(80),
        ZN => S773
    );
NOR2_X1_34: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S792(80),
        A2 => S787(80),
        ZN => S774
    );
INV_X1_192: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(74),
        ZN => S775
    );
NAND2_X1_67: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S775,
        A2 => S792(74),
        ZN => S776
    );
INV_X1_193: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(66),
        ZN => S777
    );
NAND2_X1_68: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S777,
        A2 => S787(66),
        ZN => S778
    );
OAI211_X1_5: ENTITY WORK.OAI211_X1
    PORT MAP (
        A => S778,
        B => S776,
        C1 => S773,
        C2 => S774,
        ZN => S779
    );
NOR2_X1_35: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S772,
        A2 => S779,
        ZN => S780
    );
INV_X1_194: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(82),
        ZN => S781
    );
INV_X1_195: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(84),
        ZN => S782
    );
AOI22_X1_53: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S782,
        A2 => S787(84),
        B1 => S781,
        B2 => S792(82),
        ZN => S783
    );
INV_X1_196: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(82),
        ZN => S784
    );
INV_X1_197: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(86),
        ZN => S785
    );
AOI22_X1_54: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S784,
        A2 => S787(82),
        B1 => S785,
        B2 => S792(86),
        ZN => S0
    );
INV_X1_198: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(34),
        ZN => S1
    );
INV_X1_199: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(58),
        ZN => S2
    );
AOI22_X1_55: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S1,
        A2 => S787(34),
        B1 => S2,
        B2 => S792(58),
        ZN => S3
    );
INV_X1_200: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(58),
        ZN => S4
    );
INV_X1_201: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(84),
        ZN => S5
    );
AOI22_X1_56: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S4,
        A2 => S787(58),
        B1 => S5,
        B2 => S792(84),
        ZN => S6
    );
AND4_X1_9: ENTITY WORK.AND4_X1
    PORT MAP (
        A1 => S783,
        A2 => S3,
        A3 => S6,
        A4 => S0,
        ZN => S7
    );
AND4_X1_10: ENTITY WORK.AND4_X1
    PORT MAP (
        A1 => S752,
        A2 => S7,
        A3 => S765,
        A4 => S780,
        ZN => S8
    );
INV_X1_202: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(57),
        ZN => S9
    );
NAND2_X1_69: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S9,
        A2 => S792(57),
        ZN => S10
    );
INV_X1_203: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(73),
        ZN => S11
    );
NAND2_X1_70: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S11,
        A2 => S792(73),
        ZN => S12
    );
INV_X1_204: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(79),
        ZN => S13
    );
NAND2_X1_71: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S13,
        A2 => S787(79),
        ZN => S14
    );
INV_X1_205: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(71),
        ZN => S15
    );
NAND2_X1_72: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S15,
        A2 => S787(71),
        ZN => S16
    );
NAND4_X1_26: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S14,
        A2 => S16,
        A3 => S10,
        A4 => S12,
        ZN => S17
    );
INV_X1_206: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(63),
        ZN => S18
    );
NAND2_X1_73: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S18,
        A2 => S792(63),
        ZN => S19
    );
INV_X1_207: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(63),
        ZN => S20
    );
NAND2_X1_74: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S20,
        A2 => S787(63),
        ZN => S21
    );
INV_X1_208: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(61),
        ZN => S22
    );
NAND2_X1_75: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S22,
        A2 => S787(61),
        ZN => S23
    );
INV_X1_209: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(65),
        ZN => S24
    );
NAND2_X1_76: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S24,
        A2 => S792(65),
        ZN => S25
    );
NAND4_X1_27: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S23,
        A2 => S25,
        A3 => S19,
        A4 => S21,
        ZN => S26
    );
NOR2_X1_36: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S17,
        A2 => S26,
        ZN => S27
    );
INV_X1_210: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(1),
        ZN => S28
    );
INV_X1_211: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(15),
        ZN => S29
    );
AOI22_X1_57: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S792(15),
        A2 => S29,
        B1 => S28,
        B2 => S792(1),
        ZN => S30
    );
XNOR2_X1_15: ENTITY WORK.XNOR2_X1
    PORT MAP (
        A => S792(0),
        B => S787(0),
        ZN => S31
    );
INV_X1_212: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(69),
        ZN => S32
    );
INV_X1_213: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(81),
        ZN => S33
    );
AOI22_X1_58: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S32,
        A2 => S787(69),
        B1 => S33,
        B2 => S792(81),
        ZN => S34
    );
INV_X1_214: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(13),
        ZN => S35
    );
INV_X1_215: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(21),
        ZN => S36
    );
AOI22_X1_59: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S35,
        A2 => S787(13),
        B1 => S36,
        B2 => S792(21),
        ZN => S37
    );
AND4_X1_11: ENTITY WORK.AND4_X1
    PORT MAP (
        A1 => S30,
        A2 => S37,
        A3 => S31,
        A4 => S34,
        ZN => S38
    );
INV_X1_216: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(2),
        ZN => S39
    );
NAND2_X1_77: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S39,
        A2 => S787(2),
        ZN => S40
    );
INV_X1_217: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(42),
        ZN => S41
    );
NAND2_X1_78: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S41,
        A2 => S787(42),
        ZN => S42
    );
AND2_X1_12: ENTITY WORK.AND2_X1
    PORT MAP (
        A1 => S787(4),
        A2 => S792(4),
        ZN => S43
    );
NOR2_X1_37: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S792(4),
        A2 => S787(4),
        ZN => S44
    );
OAI211_X1_6: ENTITY WORK.OAI211_X1
    PORT MAP (
        A => S42,
        B => S40,
        C1 => S43,
        C2 => S44,
        ZN => S45
    );
AND2_X1_13: ENTITY WORK.AND2_X1
    PORT MAP (
        A1 => S787(90),
        A2 => S792(90),
        ZN => S46
    );
NOR2_X1_38: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S792(90),
        A2 => S787(90),
        ZN => S47
    );
INV_X1_218: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(42),
        ZN => S48
    );
NAND2_X1_79: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S48,
        A2 => S792(42),
        ZN => S49
    );
INV_X1_219: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(2),
        ZN => S50
    );
NAND2_X1_80: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S50,
        A2 => S792(2),
        ZN => S51
    );
OAI211_X1_7: ENTITY WORK.OAI211_X1
    PORT MAP (
        A => S51,
        B => S49,
        C1 => S46,
        C2 => S47,
        ZN => S52
    );
NOR2_X1_39: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S45,
        A2 => S52,
        ZN => S53
    );
AND2_X1_14: ENTITY WORK.AND2_X1
    PORT MAP (
        A1 => S787(44),
        A2 => S792(44),
        ZN => S54
    );
NOR2_X1_40: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S792(44),
        A2 => S787(44),
        ZN => S55
    );
INV_X1_220: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(22),
        ZN => S56
    );
NAND2_X1_81: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S56,
        A2 => S792(22),
        ZN => S57
    );
INV_X1_221: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(55),
        ZN => S58
    );
NAND2_X1_82: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S58,
        A2 => S787(55),
        ZN => S59
    );
OAI211_X1_8: ENTITY WORK.OAI211_X1
    PORT MAP (
        A => S59,
        B => S57,
        C1 => S54,
        C2 => S55,
        ZN => S60
    );
INV_X1_222: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(32),
        ZN => S61
    );
NAND2_X1_83: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S61,
        A2 => S792(32),
        ZN => S62
    );
INV_X1_223: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(32),
        ZN => S63
    );
NAND2_X1_84: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S63,
        A2 => S787(32),
        ZN => S64
    );
AND2_X1_15: ENTITY WORK.AND2_X1
    PORT MAP (
        A1 => S787(46),
        A2 => S792(46),
        ZN => S65
    );
NOR2_X1_41: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S792(46),
        A2 => S787(46),
        ZN => S66
    );
OAI211_X1_9: ENTITY WORK.OAI211_X1
    PORT MAP (
        A => S64,
        B => S62,
        C1 => S65,
        C2 => S66,
        ZN => S67
    );
NOR2_X1_42: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S60,
        A2 => S67,
        ZN => S68
    );
AND4_X1_12: ENTITY WORK.AND4_X1
    PORT MAP (
        A1 => S38,
        A2 => S27,
        A3 => S53,
        A4 => S68,
        ZN => S69
    );
NAND3_X1_5: ENTITY WORK.NAND3_X1
    PORT MAP (
        A1 => S8,
        A2 => S739,
        A3 => S69,
        ZN => S70
    );
INV_X1_224: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(39),
        ZN => S71
    );
INV_X1_225: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(5),
        ZN => S72
    );
NAND2_X1_85: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S72,
        A2 => S792(5),
        ZN => S73
    );
OAI221_X1_2: ENTITY WORK.OAI221_X1
    PORT MAP (
        A => S73,
        B1 => S792(39),
        B2 => S71,
        C1 => S29,
        C2 => S792(15),
        ZN => S74
    );
INV_X1_226: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(122),
        ZN => S75
    );
NAND2_X1_86: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S75,
        A2 => S787(122),
        ZN => S76
    );
INV_X1_227: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(35),
        ZN => S77
    );
INV_X1_228: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(41),
        ZN => S78
    );
AOI22_X1_60: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S792(41),
        A2 => S78,
        B1 => S77,
        B2 => S792(35),
        ZN => S79
    );
OAI211_X1_10: ENTITY WORK.OAI211_X1
    PORT MAP (
        A => S79,
        B => S76,
        C1 => S787(71),
        C2 => S15,
        ZN => S80
    );
INV_X1_229: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(124),
        ZN => S81
    );
INV_X1_230: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(125),
        ZN => S82
    );
AOI22_X1_61: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S792(125),
        A2 => S82,
        B1 => S81,
        B2 => S792(124),
        ZN => S83
    );
OAI221_X1_3: ENTITY WORK.OAI221_X1
    PORT MAP (
        A => S83,
        B1 => S792(124),
        B2 => S81,
        C1 => S787(122),
        C2 => S75,
        ZN => S84
    );
NOR3_X1_7: ENTITY WORK.NOR3_X1
    PORT MAP (
        A1 => S84,
        A2 => S80,
        A3 => S74,
        ZN => S85
    );
XNOR2_X1_16: ENTITY WORK.XNOR2_X1
    PORT MAP (
        A => S792(48),
        B => S787(48),
        ZN => S86
    );
INV_X1_231: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(113),
        ZN => S87
    );
INV_X1_232: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(117),
        ZN => S88
    );
AOI22_X1_62: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S87,
        A2 => S787(113),
        B1 => S88,
        B2 => S792(117),
        ZN => S89
    );
XNOR2_X1_17: ENTITY WORK.XNOR2_X1
    PORT MAP (
        A => S792(24),
        B => S787(24),
        ZN => S90
    );
XNOR2_X1_18: ENTITY WORK.XNOR2_X1
    PORT MAP (
        A => S792(50),
        B => S787(50),
        ZN => S91
    );
NAND4_X1_28: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S90,
        A2 => S91,
        A3 => S86,
        A4 => S89,
        ZN => S92
    );
XNOR2_X1_19: ENTITY WORK.XNOR2_X1
    PORT MAP (
        A => S792(107),
        B => S787(107),
        ZN => S93
    );
INV_X1_233: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(119),
        ZN => S94
    );
INV_X1_234: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(123),
        ZN => S95
    );
AOI22_X1_63: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S95,
        A2 => S787(123),
        B1 => S94,
        B2 => S792(119),
        ZN => S96
    );
XNOR2_X1_20: ENTITY WORK.XNOR2_X1
    PORT MAP (
        A => S792(115),
        B => S787(115),
        ZN => S97
    );
INV_X1_235: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(125),
        ZN => S98
    );
INV_X1_236: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(127),
        ZN => S99
    );
AOI22_X1_64: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S787(125),
        A2 => S98,
        B1 => S99,
        B2 => S787(127),
        ZN => S100
    );
NAND4_X1_29: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S97,
        A2 => S100,
        A3 => S93,
        A4 => S96,
        ZN => S101
    );
NOR2_X1_43: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S92,
        A2 => S101,
        ZN => S102
    );
INV_X1_237: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(93),
        ZN => S103
    );
INV_X1_238: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(97),
        ZN => S104
    );
AOI22_X1_65: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S104,
        A2 => S787(97),
        B1 => S103,
        B2 => S792(93),
        ZN => S105
    );
XNOR2_X1_21: ENTITY WORK.XNOR2_X1
    PORT MAP (
        A => S792(116),
        B => S787(116),
        ZN => S106
    );
XNOR2_X1_22: ENTITY WORK.XNOR2_X1
    PORT MAP (
        A => S792(89),
        B => S787(89),
        ZN => S107
    );
INV_X1_239: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(59),
        ZN => S108
    );
INV_X1_240: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(61),
        ZN => S109
    );
AOI22_X1_66: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S108,
        A2 => S787(59),
        B1 => S109,
        B2 => S792(61),
        ZN => S110
    );
NAND4_X1_30: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S110,
        A2 => S107,
        A3 => S106,
        A4 => S105,
        ZN => S111
    );
XNOR2_X1_23: ENTITY WORK.XNOR2_X1
    PORT MAP (
        A => S792(106),
        B => S787(106),
        ZN => S112
    );
XNOR2_X1_24: ENTITY WORK.XNOR2_X1
    PORT MAP (
        A => S792(52),
        B => S787(52),
        ZN => S113
    );
XNOR2_X1_25: ENTITY WORK.XNOR2_X1
    PORT MAP (
        A => S792(110),
        B => S787(110),
        ZN => S114
    );
XNOR2_X1_26: ENTITY WORK.XNOR2_X1
    PORT MAP (
        A => S792(126),
        B => S787(126),
        ZN => S115
    );
NAND4_X1_31: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S114,
        A2 => S115,
        A3 => S112,
        A4 => S113,
        ZN => S116
    );
NOR2_X1_44: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S116,
        A2 => S111,
        ZN => S117
    );
NAND3_X1_6: ENTITY WORK.NAND3_X1
    PORT MAP (
        A1 => S85,
        A2 => S102,
        A3 => S117,
        ZN => S118
    );
NAND2_X1_87: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S792(78),
        A2 => S787(78),
        ZN => S119
    );
OR2_X1_10: ENTITY WORK.OR2_X1
    PORT MAP (
        A1 => S792(78),
        A2 => S787(78),
        ZN => S120
    );
NAND2_X1_88: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S792(6),
        A2 => S787(6),
        ZN => S121
    );
OR2_X1_11: ENTITY WORK.OR2_X1
    PORT MAP (
        A1 => S792(6),
        A2 => S787(6),
        ZN => S122
    );
AOI22_X1_67: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S121,
        A2 => S122,
        B1 => S120,
        B2 => S119,
        ZN => S123
    );
NAND2_X1_89: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S792(54),
        A2 => S787(54),
        ZN => S124
    );
OR2_X1_12: ENTITY WORK.OR2_X1
    PORT MAP (
        A1 => S792(54),
        A2 => S787(54),
        ZN => S125
    );
NAND2_X1_90: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S792(10),
        A2 => S787(10),
        ZN => S126
    );
OR2_X1_13: ENTITY WORK.OR2_X1
    PORT MAP (
        A1 => S792(10),
        A2 => S787(10),
        ZN => S127
    );
AOI22_X1_68: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S126,
        A2 => S127,
        B1 => S125,
        B2 => S124,
        ZN => S128
    );
INV_X1_241: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(64),
        ZN => S129
    );
NOR2_X1_45: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S129,
        A2 => S792(64),
        ZN => S130
    );
AND2_X1_16: ENTITY WORK.AND2_X1
    PORT MAP (
        A1 => S129,
        A2 => S792(64),
        ZN => S131
    );
INV_X1_242: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(31),
        ZN => S132
    );
INV_X1_243: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(51),
        ZN => S133
    );
OAI22_X1_42: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S792(31),
        A2 => S132,
        B1 => S133,
        B2 => S792(51),
        ZN => S134
    );
NOR3_X1_8: ENTITY WORK.NOR3_X1
    PORT MAP (
        A1 => S134,
        A2 => S131,
        A3 => S130,
        ZN => S135
    );
INV_X1_244: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(12),
        ZN => S136
    );
INV_X1_245: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(14),
        ZN => S137
    );
OAI22_X1_43: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S136,
        A2 => S787(12),
        B1 => S137,
        B2 => S792(14),
        ZN => S138
    );
INV_X1_246: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(8),
        ZN => S139
    );
INV_X1_247: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(14),
        ZN => S140
    );
OAI22_X1_44: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S139,
        A2 => S792(8),
        B1 => S140,
        B2 => S787(14),
        ZN => S141
    );
NOR2_X1_46: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S138,
        A2 => S141,
        ZN => S142
    );
NAND4_X1_32: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S135,
        A2 => S142,
        A3 => S123,
        A4 => S128,
        ZN => S143
    );
OAI22_X1_45: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S88,
        A2 => S792(117),
        B1 => S99,
        B2 => S787(127),
        ZN => S144
    );
INV_X1_248: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(121),
        ZN => S145
    );
OAI22_X1_46: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S145,
        A2 => S792(121),
        B1 => S95,
        B2 => S787(123),
        ZN => S146
    );
NOR2_X1_47: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S144,
        A2 => S146,
        ZN => S147
    );
INV_X1_249: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(119),
        ZN => S148
    );
AOI22_X1_69: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S148,
        A2 => S787(119),
        B1 => S145,
        B2 => S792(121),
        ZN => S149
    );
INV_X1_250: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(101),
        ZN => S150
    );
INV_X1_251: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(111),
        ZN => S151
    );
AOI22_X1_70: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S150,
        A2 => S787(101),
        B1 => S151,
        B2 => S792(111),
        ZN => S152
    );
AND2_X1_17: ENTITY WORK.AND2_X1
    PORT MAP (
        A1 => S152,
        A2 => S149,
        ZN => S153
    );
INV_X1_252: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(8),
        ZN => S154
    );
INV_X1_253: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(12),
        ZN => S155
    );
OAI22_X1_47: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S154,
        A2 => S787(8),
        B1 => S155,
        B2 => S792(12),
        ZN => S156
    );
AND2_X1_18: ENTITY WORK.AND2_X1
    PORT MAP (
        A1 => S787(62),
        A2 => S792(62),
        ZN => S157
    );
NOR2_X1_48: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S792(62),
        A2 => S787(62),
        ZN => S158
    );
NOR2_X1_49: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S157,
        A2 => S158,
        ZN => S159
    );
NOR2_X1_50: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S159,
        A2 => S156,
        ZN => S160
    );
NAND2_X1_91: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S792(120),
        A2 => S787(120),
        ZN => S161
    );
OR2_X1_14: ENTITY WORK.OR2_X1
    PORT MAP (
        A1 => S792(120),
        A2 => S787(120),
        ZN => S162
    );
NAND2_X1_92: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S792(118),
        A2 => S787(118),
        ZN => S163
    );
OR2_X1_15: ENTITY WORK.OR2_X1
    PORT MAP (
        A1 => S792(118),
        A2 => S787(118),
        ZN => S164
    );
AOI22_X1_71: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S163,
        A2 => S164,
        B1 => S162,
        B2 => S161,
        ZN => S165
    );
NAND4_X1_33: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S153,
        A2 => S147,
        A3 => S160,
        A4 => S165,
        ZN => S166
    );
NOR2_X1_51: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S166,
        A2 => S143,
        ZN => S167
    );
INV_X1_254: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(29),
        ZN => S168
    );
INV_X1_255: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(31),
        ZN => S169
    );
OAI22_X1_48: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S168,
        A2 => S792(29),
        B1 => S169,
        B2 => S787(31),
        ZN => S170
    );
OAI22_X1_49: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S787(13),
        A2 => S35,
        B1 => S104,
        B2 => S787(97),
        ZN => S171
    );
NOR2_X1_52: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S170,
        A2 => S171,
        ZN => S172
    );
INV_X1_256: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(37),
        ZN => S173
    );
AOI22_X1_72: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S173,
        A2 => S787(37),
        B1 => S71,
        B2 => S792(39),
        ZN => S174
    );
INV_X1_257: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(43),
        ZN => S175
    );
INV_X1_258: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(45),
        ZN => S176
    );
AOI22_X1_73: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S175,
        A2 => S787(43),
        B1 => S176,
        B2 => S792(45),
        ZN => S177
    );
AND2_X1_19: ENTITY WORK.AND2_X1
    PORT MAP (
        A1 => S177,
        A2 => S174,
        ZN => S178
    );
XNOR2_X1_27: ENTITY WORK.XNOR2_X1
    PORT MAP (
        A => S792(11),
        B => S787(11),
        ZN => S179
    );
INV_X1_259: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(87),
        ZN => S180
    );
INV_X1_260: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(99),
        ZN => S181
    );
AOI22_X1_74: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S180,
        A2 => S787(87),
        B1 => S181,
        B2 => S792(99),
        ZN => S182
    );
AND2_X1_20: ENTITY WORK.AND2_X1
    PORT MAP (
        A1 => S179,
        A2 => S182,
        ZN => S183
    );
INV_X1_261: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(9),
        ZN => S184
    );
INV_X1_262: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(93),
        ZN => S185
    );
AOI22_X1_75: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S787(9),
        A2 => S184,
        B1 => S185,
        B2 => S787(93),
        ZN => S186
    );
INV_X1_263: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(17),
        ZN => S187
    );
INV_X1_264: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(19),
        ZN => S188
    );
AOI22_X1_76: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S187,
        A2 => S787(17),
        B1 => S188,
        B2 => S792(19),
        ZN => S189
    );
AND2_X1_21: ENTITY WORK.AND2_X1
    PORT MAP (
        A1 => S189,
        A2 => S186,
        ZN => S190
    );
NAND4_X1_34: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S190,
        A2 => S183,
        A3 => S178,
        A4 => S172,
        ZN => S191
    );
INV_X1_265: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(77),
        ZN => S192
    );
AND2_X1_22: ENTITY WORK.AND2_X1
    PORT MAP (
        A1 => S192,
        A2 => S792(77),
        ZN => S193
    );
NOR2_X1_53: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S192,
        A2 => S792(77),
        ZN => S194
    );
OAI22_X1_50: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S77,
        A2 => S792(35),
        B1 => S173,
        B2 => S787(37),
        ZN => S195
    );
NOR3_X1_9: ENTITY WORK.NOR3_X1
    PORT MAP (
        A1 => S195,
        A2 => S193,
        A3 => S194,
        ZN => S196
    );
INV_X1_266: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(3),
        ZN => S197
    );
OAI22_X1_51: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S792(1),
        A2 => S28,
        B1 => S197,
        B2 => S792(3),
        ZN => S198
    );
OAI22_X1_52: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S9,
        A2 => S792(57),
        B1 => S108,
        B2 => S787(59),
        ZN => S199
    );
NOR2_X1_54: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S198,
        A2 => S199,
        ZN => S200
    );
INV_X1_267: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(47),
        ZN => S201
    );
OAI22_X1_53: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S787(17),
        A2 => S187,
        B1 => S201,
        B2 => S787(47),
        ZN => S202
    );
OAI22_X1_54: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S151,
        A2 => S792(111),
        B1 => S87,
        B2 => S787(113),
        ZN => S203
    );
NOR2_X1_55: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S202,
        A2 => S203,
        ZN => S204
    );
INV_X1_268: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(85),
        ZN => S205
    );
OAI22_X1_55: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S33,
        A2 => S792(81),
        B1 => S205,
        B2 => S787(85),
        ZN => S206
    );
INV_X1_269: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(23),
        ZN => S207
    );
INV_X1_270: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(27),
        ZN => S208
    );
OAI22_X1_56: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S787(23),
        A2 => S207,
        B1 => S208,
        B2 => S787(27),
        ZN => S209
    );
NOR2_X1_56: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S206,
        A2 => S209,
        ZN => S210
    );
NAND4_X1_35: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S196,
        A2 => S200,
        A3 => S204,
        A4 => S210,
        ZN => S211
    );
NOR2_X1_57: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S191,
        A2 => S211,
        ZN => S212
    );
INV_X1_271: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(103),
        ZN => S213
    );
INV_X1_272: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(105),
        ZN => S214
    );
OAI22_X1_57: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S213,
        A2 => S792(103),
        B1 => S214,
        B2 => S787(105),
        ZN => S215
    );
OAI22_X1_58: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S78,
        A2 => S792(41),
        B1 => S175,
        B2 => S787(43),
        ZN => S216
    );
NOR2_X1_58: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S215,
        A2 => S216,
        ZN => S217
    );
INV_X1_273: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(53),
        ZN => S218
    );
OAI22_X1_59: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S218,
        A2 => S792(53),
        B1 => S58,
        B2 => S787(55),
        ZN => S219
    );
INV_X1_274: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(83),
        ZN => S220
    );
AND2_X1_23: ENTITY WORK.AND2_X1
    PORT MAP (
        A1 => S220,
        A2 => S792(83),
        ZN => S221
    );
NOR2_X1_59: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S220,
        A2 => S792(83),
        ZN => S222
    );
NOR3_X1_10: ENTITY WORK.NOR3_X1
    PORT MAP (
        A1 => S219,
        A2 => S221,
        A3 => S222,
        ZN => S223
    );
OAI22_X1_60: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S72,
        A2 => S792(5),
        B1 => S184,
        B2 => S787(9),
        ZN => S224
    );
XOR2_X1_2: ENTITY WORK.XOR2_X1
    PORT MAP (
        A => S792(7),
        B => S787(7),
        Z => S225
    );
NOR2_X1_60: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S225,
        A2 => S224,
        ZN => S226
    );
INV_X1_275: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(49),
        ZN => S227
    );
NAND2_X1_93: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S227,
        A2 => S792(49),
        ZN => S228
    );
NAND2_X1_94: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S201,
        A2 => S787(47),
        ZN => S229
    );
INV_X1_276: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(25),
        ZN => S230
    );
NAND2_X1_95: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S230,
        A2 => S792(25),
        ZN => S231
    );
NAND2_X1_96: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S207,
        A2 => S787(23),
        ZN => S232
    );
AND4_X1_13: ENTITY WORK.AND4_X1
    PORT MAP (
        A1 => S228,
        A2 => S231,
        A3 => S232,
        A4 => S229,
        ZN => S233
    );
NAND4_X1_36: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S226,
        A2 => S223,
        A3 => S217,
        A4 => S233,
        ZN => S234
    );
INV_X1_277: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(29),
        ZN => S235
    );
OAI22_X1_61: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S235,
        A2 => S787(29),
        B1 => S176,
        B2 => S792(45),
        ZN => S236
    );
OAI22_X1_62: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S792(21),
        A2 => S36,
        B1 => S227,
        B2 => S792(49),
        ZN => S237
    );
NOR2_X1_61: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S236,
        A2 => S237,
        ZN => S238
    );
INV_X1_278: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(3),
        ZN => S239
    );
OAI22_X1_63: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S239,
        A2 => S787(3),
        B1 => S188,
        B2 => S792(19),
        ZN => S240
    );
INV_X1_279: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(27),
        ZN => S241
    );
INV_X1_280: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(33),
        ZN => S242
    );
OAI22_X1_64: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S792(27),
        A2 => S241,
        B1 => S242,
        B2 => S792(33),
        ZN => S243
    );
NOR2_X1_62: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S240,
        A2 => S243,
        ZN => S244
    );
OAI22_X1_65: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S11,
        A2 => S792(73),
        B1 => S13,
        B2 => S787(79),
        ZN => S245
    );
INV_X1_281: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(75),
        ZN => S246
    );
AND2_X1_24: ENTITY WORK.AND2_X1
    PORT MAP (
        A1 => S246,
        A2 => S792(75),
        ZN => S247
    );
NOR2_X1_63: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S246,
        A2 => S792(75),
        ZN => S248
    );
NOR3_X1_11: ENTITY WORK.NOR3_X1
    PORT MAP (
        A1 => S245,
        A2 => S247,
        A3 => S248,
        ZN => S249
    );
INV_X1_282: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(33),
        ZN => S250
    );
OAI22_X1_66: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S230,
        A2 => S792(25),
        B1 => S250,
        B2 => S787(33),
        ZN => S251
    );
INV_X1_283: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(51),
        ZN => S252
    );
INV_X1_284: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(53),
        ZN => S253
    );
OAI22_X1_67: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S787(51),
        A2 => S252,
        B1 => S253,
        B2 => S787(53),
        ZN => S254
    );
NOR2_X1_64: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S251,
        A2 => S254,
        ZN => S255
    );
NAND4_X1_37: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S249,
        A2 => S255,
        A3 => S238,
        A4 => S244,
        ZN => S256
    );
NOR2_X1_65: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S234,
        A2 => S256,
        ZN => S257
    );
NAND2_X1_97: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S792(28),
        A2 => S787(28),
        ZN => S258
    );
OR2_X1_16: ENTITY WORK.OR2_X1
    PORT MAP (
        A1 => S792(28),
        A2 => S787(28),
        ZN => S259
    );
NAND2_X1_98: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S792(26),
        A2 => S787(26),
        ZN => S260
    );
OR2_X1_17: ENTITY WORK.OR2_X1
    PORT MAP (
        A1 => S792(26),
        A2 => S787(26),
        ZN => S261
    );
AOI22_X1_77: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S260,
        A2 => S261,
        B1 => S259,
        B2 => S258,
        ZN => S262
    );
NAND2_X1_99: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S792(108),
        A2 => S787(108),
        ZN => S263
    );
OR2_X1_18: ENTITY WORK.OR2_X1
    PORT MAP (
        A1 => S792(108),
        A2 => S787(108),
        ZN => S264
    );
NAND2_X1_100: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S792(102),
        A2 => S787(102),
        ZN => S265
    );
OR2_X1_19: ENTITY WORK.OR2_X1
    PORT MAP (
        A1 => S792(102),
        A2 => S787(102),
        ZN => S266
    );
AOI22_X1_78: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S265,
        A2 => S266,
        B1 => S264,
        B2 => S263,
        ZN => S267
    );
INV_X1_285: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(103),
        ZN => S268
    );
INV_X1_286: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(109),
        ZN => S269
    );
OAI22_X1_68: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S787(103),
        A2 => S268,
        B1 => S269,
        B2 => S787(109),
        ZN => S270
    );
INV_X1_287: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(105),
        ZN => S271
    );
INV_X1_288: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(109),
        ZN => S272
    );
OAI22_X1_69: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S792(105),
        A2 => S271,
        B1 => S272,
        B2 => S792(109),
        ZN => S273
    );
NOR2_X1_66: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S270,
        A2 => S273,
        ZN => S274
    );
NAND2_X1_101: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S792(112),
        A2 => S787(112),
        ZN => S275
    );
OR2_X1_20: ENTITY WORK.OR2_X1
    PORT MAP (
        A1 => S792(112),
        A2 => S787(112),
        ZN => S276
    );
NAND2_X1_102: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S792(38),
        A2 => S787(38),
        ZN => S277
    );
OR2_X1_21: ENTITY WORK.OR2_X1
    PORT MAP (
        A1 => S792(38),
        A2 => S787(38),
        ZN => S278
    );
AOI22_X1_79: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S277,
        A2 => S278,
        B1 => S276,
        B2 => S275,
        ZN => S279
    );
NAND4_X1_38: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S274,
        A2 => S279,
        A3 => S262,
        A4 => S267,
        ZN => S280
    );
INV_X1_289: ENTITY WORK.INV_X1
    PORT MAP (
        A => S792(67),
        ZN => S281
    );
OAI22_X1_70: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S24,
        A2 => S792(65),
        B1 => S281,
        B2 => S787(67),
        ZN => S282
    );
INV_X1_290: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(67),
        ZN => S283
    );
OAI22_X1_71: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S283,
        A2 => S792(67),
        B1 => S32,
        B2 => S787(69),
        ZN => S284
    );
NOR2_X1_67: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S282,
        A2 => S284,
        ZN => S285
    );
OAI22_X1_72: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S181,
        A2 => S792(99),
        B1 => S150,
        B2 => S787(101),
        ZN => S286
    );
INV_X1_291: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(95),
        ZN => S287
    );
AND2_X1_25: ENTITY WORK.AND2_X1
    PORT MAP (
        A1 => S287,
        A2 => S792(95),
        ZN => S288
    );
NOR2_X1_68: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S287,
        A2 => S792(95),
        ZN => S289
    );
NOR3_X1_12: ENTITY WORK.NOR3_X1
    PORT MAP (
        A1 => S286,
        A2 => S288,
        A3 => S289,
        ZN => S290
    );
NAND2_X1_103: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S792(114),
        A2 => S787(114),
        ZN => S291
    );
OR2_X1_22: ENTITY WORK.OR2_X1
    PORT MAP (
        A1 => S792(114),
        A2 => S787(114),
        ZN => S292
    );
NAND2_X1_104: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => S792(104),
        A2 => S787(104),
        ZN => S293
    );
OR2_X1_23: ENTITY WORK.OR2_X1
    PORT MAP (
        A1 => S792(104),
        A2 => S787(104),
        ZN => S294
    );
AOI22_X1_80: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => S293,
        A2 => S294,
        B1 => S292,
        B2 => S291,
        ZN => S295
    );
INV_X1_292: ENTITY WORK.INV_X1
    PORT MAP (
        A => S787(85),
        ZN => S296
    );
OAI22_X1_73: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => S296,
        A2 => S792(85),
        B1 => S180,
        B2 => S787(87),
        ZN => S297
    );
XOR2_X1_3: ENTITY WORK.XOR2_X1
    PORT MAP (
        A => S792(91),
        B => S787(91),
        Z => S298
    );
NOR2_X1_69: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S298,
        A2 => S297,
        ZN => S299
    );
NAND4_X1_39: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S299,
        A2 => S290,
        A3 => S295,
        A4 => S285,
        ZN => S300
    );
NOR2_X1_70: ENTITY WORK.NOR2_X1
    PORT MAP (
        A1 => S300,
        A2 => S280,
        ZN => S301
    );
NAND4_X1_40: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => S212,
        A2 => S257,
        A3 => S167,
        A4 => S301,
        ZN => S302
    );
NOR3_X1_13: ENTITY WORK.NOR3_X1
    PORT MAP (
        A1 => S302,
        A2 => S70,
        A3 => S118,
        ZN => S786
    );
BUF_X1_1: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S786,
        Z => d128
    );
BUF_X1_2: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(0),
        Z => decrypted128(0)
    );
BUF_X1_3: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(1),
        Z => decrypted128(1)
    );
BUF_X1_4: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(10),
        Z => decrypted128(10)
    );
BUF_X1_5: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(100),
        Z => decrypted128(100)
    );
BUF_X1_6: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(101),
        Z => decrypted128(101)
    );
BUF_X1_7: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(102),
        Z => decrypted128(102)
    );
BUF_X1_8: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(103),
        Z => decrypted128(103)
    );
BUF_X1_9: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(104),
        Z => decrypted128(104)
    );
BUF_X1_10: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(105),
        Z => decrypted128(105)
    );
BUF_X1_11: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(106),
        Z => decrypted128(106)
    );
BUF_X1_12: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(107),
        Z => decrypted128(107)
    );
BUF_X1_13: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(108),
        Z => decrypted128(108)
    );
BUF_X1_14: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(109),
        Z => decrypted128(109)
    );
BUF_X1_15: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(11),
        Z => decrypted128(11)
    );
BUF_X1_16: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(110),
        Z => decrypted128(110)
    );
BUF_X1_17: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(111),
        Z => decrypted128(111)
    );
BUF_X1_18: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(112),
        Z => decrypted128(112)
    );
BUF_X1_19: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(113),
        Z => decrypted128(113)
    );
BUF_X1_20: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(114),
        Z => decrypted128(114)
    );
BUF_X1_21: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(115),
        Z => decrypted128(115)
    );
BUF_X1_22: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(116),
        Z => decrypted128(116)
    );
BUF_X1_23: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(117),
        Z => decrypted128(117)
    );
BUF_X1_24: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(118),
        Z => decrypted128(118)
    );
BUF_X1_25: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(119),
        Z => decrypted128(119)
    );
BUF_X1_26: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(12),
        Z => decrypted128(12)
    );
BUF_X1_27: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(120),
        Z => decrypted128(120)
    );
BUF_X1_28: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(121),
        Z => decrypted128(121)
    );
BUF_X1_29: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(122),
        Z => decrypted128(122)
    );
BUF_X1_30: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(123),
        Z => decrypted128(123)
    );
BUF_X1_31: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(124),
        Z => decrypted128(124)
    );
BUF_X1_32: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(125),
        Z => decrypted128(125)
    );
BUF_X1_33: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(126),
        Z => decrypted128(126)
    );
BUF_X1_34: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(127),
        Z => decrypted128(127)
    );
BUF_X1_35: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(13),
        Z => decrypted128(13)
    );
BUF_X1_36: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(14),
        Z => decrypted128(14)
    );
BUF_X1_37: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(15),
        Z => decrypted128(15)
    );
BUF_X1_38: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(16),
        Z => decrypted128(16)
    );
BUF_X1_39: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(17),
        Z => decrypted128(17)
    );
BUF_X1_40: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(18),
        Z => decrypted128(18)
    );
BUF_X1_41: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(19),
        Z => decrypted128(19)
    );
BUF_X1_42: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(2),
        Z => decrypted128(2)
    );
BUF_X1_43: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(20),
        Z => decrypted128(20)
    );
BUF_X1_44: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(21),
        Z => decrypted128(21)
    );
BUF_X1_45: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(22),
        Z => decrypted128(22)
    );
BUF_X1_46: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(23),
        Z => decrypted128(23)
    );
BUF_X1_47: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(24),
        Z => decrypted128(24)
    );
BUF_X1_48: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(25),
        Z => decrypted128(25)
    );
BUF_X1_49: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(26),
        Z => decrypted128(26)
    );
BUF_X1_50: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(27),
        Z => decrypted128(27)
    );
BUF_X1_51: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(28),
        Z => decrypted128(28)
    );
BUF_X1_52: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(29),
        Z => decrypted128(29)
    );
BUF_X1_53: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(3),
        Z => decrypted128(3)
    );
BUF_X1_54: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(30),
        Z => decrypted128(30)
    );
BUF_X1_55: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(31),
        Z => decrypted128(31)
    );
BUF_X1_56: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(32),
        Z => decrypted128(32)
    );
BUF_X1_57: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(33),
        Z => decrypted128(33)
    );
BUF_X1_58: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(34),
        Z => decrypted128(34)
    );
BUF_X1_59: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(35),
        Z => decrypted128(35)
    );
BUF_X1_60: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(36),
        Z => decrypted128(36)
    );
BUF_X1_61: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(37),
        Z => decrypted128(37)
    );
BUF_X1_62: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(38),
        Z => decrypted128(38)
    );
BUF_X1_63: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(39),
        Z => decrypted128(39)
    );
BUF_X1_64: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(4),
        Z => decrypted128(4)
    );
BUF_X1_65: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(40),
        Z => decrypted128(40)
    );
BUF_X1_66: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(41),
        Z => decrypted128(41)
    );
BUF_X1_67: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(42),
        Z => decrypted128(42)
    );
BUF_X1_68: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(43),
        Z => decrypted128(43)
    );
BUF_X1_69: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(44),
        Z => decrypted128(44)
    );
BUF_X1_70: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(45),
        Z => decrypted128(45)
    );
BUF_X1_71: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(46),
        Z => decrypted128(46)
    );
BUF_X1_72: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(47),
        Z => decrypted128(47)
    );
BUF_X1_73: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(48),
        Z => decrypted128(48)
    );
BUF_X1_74: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(49),
        Z => decrypted128(49)
    );
BUF_X1_75: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(5),
        Z => decrypted128(5)
    );
BUF_X1_76: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(50),
        Z => decrypted128(50)
    );
BUF_X1_77: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(51),
        Z => decrypted128(51)
    );
BUF_X1_78: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(52),
        Z => decrypted128(52)
    );
BUF_X1_79: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(53),
        Z => decrypted128(53)
    );
BUF_X1_80: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(54),
        Z => decrypted128(54)
    );
BUF_X1_81: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(55),
        Z => decrypted128(55)
    );
BUF_X1_82: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(56),
        Z => decrypted128(56)
    );
BUF_X1_83: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(57),
        Z => decrypted128(57)
    );
BUF_X1_84: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(58),
        Z => decrypted128(58)
    );
BUF_X1_85: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(59),
        Z => decrypted128(59)
    );
BUF_X1_86: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(6),
        Z => decrypted128(6)
    );
BUF_X1_87: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(60),
        Z => decrypted128(60)
    );
BUF_X1_88: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(61),
        Z => decrypted128(61)
    );
BUF_X1_89: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(62),
        Z => decrypted128(62)
    );
BUF_X1_90: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(63),
        Z => decrypted128(63)
    );
BUF_X1_91: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(64),
        Z => decrypted128(64)
    );
BUF_X1_92: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(65),
        Z => decrypted128(65)
    );
BUF_X1_93: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(66),
        Z => decrypted128(66)
    );
BUF_X1_94: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(67),
        Z => decrypted128(67)
    );
BUF_X1_95: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(68),
        Z => decrypted128(68)
    );
BUF_X1_96: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(69),
        Z => decrypted128(69)
    );
BUF_X1_97: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(7),
        Z => decrypted128(7)
    );
BUF_X1_98: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(70),
        Z => decrypted128(70)
    );
BUF_X1_99: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(71),
        Z => decrypted128(71)
    );
BUF_X1_100: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(72),
        Z => decrypted128(72)
    );
BUF_X1_101: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(73),
        Z => decrypted128(73)
    );
BUF_X1_102: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(74),
        Z => decrypted128(74)
    );
BUF_X1_103: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(75),
        Z => decrypted128(75)
    );
BUF_X1_104: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(76),
        Z => decrypted128(76)
    );
BUF_X1_105: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(77),
        Z => decrypted128(77)
    );
BUF_X1_106: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(78),
        Z => decrypted128(78)
    );
BUF_X1_107: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(79),
        Z => decrypted128(79)
    );
BUF_X1_108: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(8),
        Z => decrypted128(8)
    );
BUF_X1_109: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(80),
        Z => decrypted128(80)
    );
BUF_X1_110: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(81),
        Z => decrypted128(81)
    );
BUF_X1_111: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(82),
        Z => decrypted128(82)
    );
BUF_X1_112: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(83),
        Z => decrypted128(83)
    );
BUF_X1_113: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(84),
        Z => decrypted128(84)
    );
BUF_X1_114: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(85),
        Z => decrypted128(85)
    );
BUF_X1_115: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(86),
        Z => decrypted128(86)
    );
BUF_X1_116: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(87),
        Z => decrypted128(87)
    );
BUF_X1_117: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(88),
        Z => decrypted128(88)
    );
BUF_X1_118: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(89),
        Z => decrypted128(89)
    );
BUF_X1_119: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(9),
        Z => decrypted128(9)
    );
BUF_X1_120: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(90),
        Z => decrypted128(90)
    );
BUF_X1_121: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(91),
        Z => decrypted128(91)
    );
BUF_X1_122: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(92),
        Z => decrypted128(92)
    );
BUF_X1_123: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(93),
        Z => decrypted128(93)
    );
BUF_X1_124: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(94),
        Z => decrypted128(94)
    );
BUF_X1_125: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(95),
        Z => decrypted128(95)
    );
BUF_X1_126: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(96),
        Z => decrypted128(96)
    );
BUF_X1_127: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(97),
        Z => decrypted128(97)
    );
BUF_X1_128: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(98),
        Z => decrypted128(98)
    );
BUF_X1_129: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S787(99),
        Z => decrypted128(99)
    );
BUF_X1_130: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S788,
        Z => e128
    );
BUF_X1_131: ENTITY WORK.BUF_X1
    PORT MAP (
        A => enable,
        Z => S789
    );
BUF_X1_132: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(0),
        Z => encrypted128(0)
    );
BUF_X1_133: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(1),
        Z => encrypted128(1)
    );
BUF_X1_134: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(10),
        Z => encrypted128(10)
    );
BUF_X1_135: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(100),
        Z => encrypted128(100)
    );
BUF_X1_136: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(101),
        Z => encrypted128(101)
    );
BUF_X1_137: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(102),
        Z => encrypted128(102)
    );
BUF_X1_138: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(103),
        Z => encrypted128(103)
    );
BUF_X1_139: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(104),
        Z => encrypted128(104)
    );
BUF_X1_140: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(105),
        Z => encrypted128(105)
    );
BUF_X1_141: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(106),
        Z => encrypted128(106)
    );
BUF_X1_142: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(107),
        Z => encrypted128(107)
    );
BUF_X1_143: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(108),
        Z => encrypted128(108)
    );
BUF_X1_144: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(109),
        Z => encrypted128(109)
    );
BUF_X1_145: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(11),
        Z => encrypted128(11)
    );
BUF_X1_146: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(110),
        Z => encrypted128(110)
    );
BUF_X1_147: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(111),
        Z => encrypted128(111)
    );
BUF_X1_148: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(112),
        Z => encrypted128(112)
    );
BUF_X1_149: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(113),
        Z => encrypted128(113)
    );
BUF_X1_150: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(114),
        Z => encrypted128(114)
    );
BUF_X1_151: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(115),
        Z => encrypted128(115)
    );
BUF_X1_152: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(116),
        Z => encrypted128(116)
    );
BUF_X1_153: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(117),
        Z => encrypted128(117)
    );
BUF_X1_154: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(118),
        Z => encrypted128(118)
    );
BUF_X1_155: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(119),
        Z => encrypted128(119)
    );
BUF_X1_156: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(12),
        Z => encrypted128(12)
    );
BUF_X1_157: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(120),
        Z => encrypted128(120)
    );
BUF_X1_158: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(121),
        Z => encrypted128(121)
    );
BUF_X1_159: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(122),
        Z => encrypted128(122)
    );
BUF_X1_160: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(123),
        Z => encrypted128(123)
    );
BUF_X1_161: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(124),
        Z => encrypted128(124)
    );
BUF_X1_162: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(125),
        Z => encrypted128(125)
    );
BUF_X1_163: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(126),
        Z => encrypted128(126)
    );
BUF_X1_164: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(127),
        Z => encrypted128(127)
    );
BUF_X1_165: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(13),
        Z => encrypted128(13)
    );
BUF_X1_166: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(14),
        Z => encrypted128(14)
    );
BUF_X1_167: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(15),
        Z => encrypted128(15)
    );
BUF_X1_168: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(16),
        Z => encrypted128(16)
    );
BUF_X1_169: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(17),
        Z => encrypted128(17)
    );
BUF_X1_170: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(18),
        Z => encrypted128(18)
    );
BUF_X1_171: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(19),
        Z => encrypted128(19)
    );
BUF_X1_172: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(2),
        Z => encrypted128(2)
    );
BUF_X1_173: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(20),
        Z => encrypted128(20)
    );
BUF_X1_174: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(21),
        Z => encrypted128(21)
    );
BUF_X1_175: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(22),
        Z => encrypted128(22)
    );
BUF_X1_176: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(23),
        Z => encrypted128(23)
    );
BUF_X1_177: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(24),
        Z => encrypted128(24)
    );
BUF_X1_178: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(25),
        Z => encrypted128(25)
    );
BUF_X1_179: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(26),
        Z => encrypted128(26)
    );
BUF_X1_180: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(27),
        Z => encrypted128(27)
    );
BUF_X1_181: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(28),
        Z => encrypted128(28)
    );
BUF_X1_182: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(29),
        Z => encrypted128(29)
    );
BUF_X1_183: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(3),
        Z => encrypted128(3)
    );
BUF_X1_184: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(30),
        Z => encrypted128(30)
    );
BUF_X1_185: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(31),
        Z => encrypted128(31)
    );
BUF_X1_186: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(32),
        Z => encrypted128(32)
    );
BUF_X1_187: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(33),
        Z => encrypted128(33)
    );
BUF_X1_188: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(34),
        Z => encrypted128(34)
    );
BUF_X1_189: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(35),
        Z => encrypted128(35)
    );
BUF_X1_190: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(36),
        Z => encrypted128(36)
    );
BUF_X1_191: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(37),
        Z => encrypted128(37)
    );
BUF_X1_192: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(38),
        Z => encrypted128(38)
    );
BUF_X1_193: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(39),
        Z => encrypted128(39)
    );
BUF_X1_194: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(4),
        Z => encrypted128(4)
    );
BUF_X1_195: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(40),
        Z => encrypted128(40)
    );
BUF_X1_196: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(41),
        Z => encrypted128(41)
    );
BUF_X1_197: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(42),
        Z => encrypted128(42)
    );
BUF_X1_198: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(43),
        Z => encrypted128(43)
    );
BUF_X1_199: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(44),
        Z => encrypted128(44)
    );
BUF_X1_200: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(45),
        Z => encrypted128(45)
    );
BUF_X1_201: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(46),
        Z => encrypted128(46)
    );
BUF_X1_202: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(47),
        Z => encrypted128(47)
    );
BUF_X1_203: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(48),
        Z => encrypted128(48)
    );
BUF_X1_204: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(49),
        Z => encrypted128(49)
    );
BUF_X1_205: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(5),
        Z => encrypted128(5)
    );
BUF_X1_206: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(50),
        Z => encrypted128(50)
    );
BUF_X1_207: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(51),
        Z => encrypted128(51)
    );
BUF_X1_208: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(52),
        Z => encrypted128(52)
    );
BUF_X1_209: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(53),
        Z => encrypted128(53)
    );
BUF_X1_210: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(54),
        Z => encrypted128(54)
    );
BUF_X1_211: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(55),
        Z => encrypted128(55)
    );
BUF_X1_212: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(56),
        Z => encrypted128(56)
    );
BUF_X1_213: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(57),
        Z => encrypted128(57)
    );
BUF_X1_214: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(58),
        Z => encrypted128(58)
    );
BUF_X1_215: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(59),
        Z => encrypted128(59)
    );
BUF_X1_216: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(6),
        Z => encrypted128(6)
    );
BUF_X1_217: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(60),
        Z => encrypted128(60)
    );
BUF_X1_218: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(61),
        Z => encrypted128(61)
    );
BUF_X1_219: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(62),
        Z => encrypted128(62)
    );
BUF_X1_220: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(63),
        Z => encrypted128(63)
    );
BUF_X1_221: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(64),
        Z => encrypted128(64)
    );
BUF_X1_222: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(65),
        Z => encrypted128(65)
    );
BUF_X1_223: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(66),
        Z => encrypted128(66)
    );
BUF_X1_224: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(67),
        Z => encrypted128(67)
    );
BUF_X1_225: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(68),
        Z => encrypted128(68)
    );
BUF_X1_226: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(69),
        Z => encrypted128(69)
    );
BUF_X1_227: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(7),
        Z => encrypted128(7)
    );
BUF_X1_228: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(70),
        Z => encrypted128(70)
    );
BUF_X1_229: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(71),
        Z => encrypted128(71)
    );
BUF_X1_230: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(72),
        Z => encrypted128(72)
    );
BUF_X1_231: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(73),
        Z => encrypted128(73)
    );
BUF_X1_232: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(74),
        Z => encrypted128(74)
    );
BUF_X1_233: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(75),
        Z => encrypted128(75)
    );
BUF_X1_234: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(76),
        Z => encrypted128(76)
    );
BUF_X1_235: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(77),
        Z => encrypted128(77)
    );
BUF_X1_236: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(78),
        Z => encrypted128(78)
    );
BUF_X1_237: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(79),
        Z => encrypted128(79)
    );
BUF_X1_238: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(8),
        Z => encrypted128(8)
    );
BUF_X1_239: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(80),
        Z => encrypted128(80)
    );
BUF_X1_240: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(81),
        Z => encrypted128(81)
    );
BUF_X1_241: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(82),
        Z => encrypted128(82)
    );
BUF_X1_242: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(83),
        Z => encrypted128(83)
    );
BUF_X1_243: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(84),
        Z => encrypted128(84)
    );
BUF_X1_244: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(85),
        Z => encrypted128(85)
    );
BUF_X1_245: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(86),
        Z => encrypted128(86)
    );
BUF_X1_246: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(87),
        Z => encrypted128(87)
    );
BUF_X1_247: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(88),
        Z => encrypted128(88)
    );
BUF_X1_248: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(89),
        Z => encrypted128(89)
    );
BUF_X1_249: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(9),
        Z => encrypted128(9)
    );
BUF_X1_250: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(90),
        Z => encrypted128(90)
    );
BUF_X1_251: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(91),
        Z => encrypted128(91)
    );
BUF_X1_252: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(92),
        Z => encrypted128(92)
    );
BUF_X1_253: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(93),
        Z => encrypted128(93)
    );
BUF_X1_254: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(94),
        Z => encrypted128(94)
    );
BUF_X1_255: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(95),
        Z => encrypted128(95)
    );
BUF_X1_256: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(96),
        Z => encrypted128(96)
    );
BUF_X1_257: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(97),
        Z => encrypted128(97)
    );
BUF_X1_258: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(98),
        Z => encrypted128(98)
    );
BUF_X1_259: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S790(99),
        Z => encrypted128(99)
    );
BUF_X1_260: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(0),
        Z => S791(0)
    );
BUF_X1_261: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(1),
        Z => S791(1)
    );
BUF_X1_262: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(10),
        Z => S791(10)
    );
BUF_X1_263: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(100),
        Z => S791(100)
    );
BUF_X1_264: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(101),
        Z => S791(101)
    );
BUF_X1_265: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(102),
        Z => S791(102)
    );
BUF_X1_266: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(103),
        Z => S791(103)
    );
BUF_X1_267: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(104),
        Z => S791(104)
    );
BUF_X1_268: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(105),
        Z => S791(105)
    );
BUF_X1_269: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(106),
        Z => S791(106)
    );
BUF_X1_270: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(107),
        Z => S791(107)
    );
BUF_X1_271: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(108),
        Z => S791(108)
    );
BUF_X1_272: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(109),
        Z => S791(109)
    );
BUF_X1_273: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(11),
        Z => S791(11)
    );
BUF_X1_274: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(110),
        Z => S791(110)
    );
BUF_X1_275: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(111),
        Z => S791(111)
    );
BUF_X1_276: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(112),
        Z => S791(112)
    );
BUF_X1_277: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(113),
        Z => S791(113)
    );
BUF_X1_278: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(114),
        Z => S791(114)
    );
BUF_X1_279: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(115),
        Z => S791(115)
    );
BUF_X1_280: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(116),
        Z => S791(116)
    );
BUF_X1_281: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(117),
        Z => S791(117)
    );
BUF_X1_282: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(118),
        Z => S791(118)
    );
BUF_X1_283: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(119),
        Z => S791(119)
    );
BUF_X1_284: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(12),
        Z => S791(12)
    );
BUF_X1_285: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(120),
        Z => S791(120)
    );
BUF_X1_286: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(121),
        Z => S791(121)
    );
BUF_X1_287: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(122),
        Z => S791(122)
    );
BUF_X1_288: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(123),
        Z => S791(123)
    );
BUF_X1_289: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(124),
        Z => S791(124)
    );
BUF_X1_290: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(125),
        Z => S791(125)
    );
BUF_X1_291: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(126),
        Z => S791(126)
    );
BUF_X1_292: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(127),
        Z => S791(127)
    );
BUF_X1_293: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(13),
        Z => S791(13)
    );
BUF_X1_294: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(14),
        Z => S791(14)
    );
BUF_X1_295: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(15),
        Z => S791(15)
    );
BUF_X1_296: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(16),
        Z => S791(16)
    );
BUF_X1_297: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(17),
        Z => S791(17)
    );
BUF_X1_298: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(18),
        Z => S791(18)
    );
BUF_X1_299: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(19),
        Z => S791(19)
    );
BUF_X1_300: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(2),
        Z => S791(2)
    );
BUF_X1_301: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(20),
        Z => S791(20)
    );
BUF_X1_302: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(21),
        Z => S791(21)
    );
BUF_X1_303: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(22),
        Z => S791(22)
    );
BUF_X1_304: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(23),
        Z => S791(23)
    );
BUF_X1_305: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(24),
        Z => S791(24)
    );
BUF_X1_306: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(25),
        Z => S791(25)
    );
BUF_X1_307: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(26),
        Z => S791(26)
    );
BUF_X1_308: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(27),
        Z => S791(27)
    );
BUF_X1_309: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(28),
        Z => S791(28)
    );
BUF_X1_310: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(29),
        Z => S791(29)
    );
BUF_X1_311: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(3),
        Z => S791(3)
    );
BUF_X1_312: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(30),
        Z => S791(30)
    );
BUF_X1_313: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(31),
        Z => S791(31)
    );
BUF_X1_314: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(32),
        Z => S791(32)
    );
BUF_X1_315: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(33),
        Z => S791(33)
    );
BUF_X1_316: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(34),
        Z => S791(34)
    );
BUF_X1_317: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(35),
        Z => S791(35)
    );
BUF_X1_318: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(36),
        Z => S791(36)
    );
BUF_X1_319: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(37),
        Z => S791(37)
    );
BUF_X1_320: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(38),
        Z => S791(38)
    );
BUF_X1_321: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(39),
        Z => S791(39)
    );
BUF_X1_322: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(4),
        Z => S791(4)
    );
BUF_X1_323: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(40),
        Z => S791(40)
    );
BUF_X1_324: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(41),
        Z => S791(41)
    );
BUF_X1_325: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(42),
        Z => S791(42)
    );
BUF_X1_326: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(43),
        Z => S791(43)
    );
BUF_X1_327: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(44),
        Z => S791(44)
    );
BUF_X1_328: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(45),
        Z => S791(45)
    );
BUF_X1_329: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(46),
        Z => S791(46)
    );
BUF_X1_330: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(47),
        Z => S791(47)
    );
BUF_X1_331: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(48),
        Z => S791(48)
    );
BUF_X1_332: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(49),
        Z => S791(49)
    );
BUF_X1_333: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(5),
        Z => S791(5)
    );
BUF_X1_334: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(50),
        Z => S791(50)
    );
BUF_X1_335: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(51),
        Z => S791(51)
    );
BUF_X1_336: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(52),
        Z => S791(52)
    );
BUF_X1_337: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(53),
        Z => S791(53)
    );
BUF_X1_338: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(54),
        Z => S791(54)
    );
BUF_X1_339: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(55),
        Z => S791(55)
    );
BUF_X1_340: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(56),
        Z => S791(56)
    );
BUF_X1_341: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(57),
        Z => S791(57)
    );
BUF_X1_342: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(58),
        Z => S791(58)
    );
BUF_X1_343: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(59),
        Z => S791(59)
    );
BUF_X1_344: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(6),
        Z => S791(6)
    );
BUF_X1_345: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(60),
        Z => S791(60)
    );
BUF_X1_346: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(61),
        Z => S791(61)
    );
BUF_X1_347: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(62),
        Z => S791(62)
    );
BUF_X1_348: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(63),
        Z => S791(63)
    );
BUF_X1_349: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(64),
        Z => S791(64)
    );
BUF_X1_350: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(65),
        Z => S791(65)
    );
BUF_X1_351: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(66),
        Z => S791(66)
    );
BUF_X1_352: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(67),
        Z => S791(67)
    );
BUF_X1_353: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(68),
        Z => S791(68)
    );
BUF_X1_354: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(69),
        Z => S791(69)
    );
BUF_X1_355: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(7),
        Z => S791(7)
    );
BUF_X1_356: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(70),
        Z => S791(70)
    );
BUF_X1_357: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(71),
        Z => S791(71)
    );
BUF_X1_358: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(72),
        Z => S791(72)
    );
BUF_X1_359: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(73),
        Z => S791(73)
    );
BUF_X1_360: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(74),
        Z => S791(74)
    );
BUF_X1_361: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(75),
        Z => S791(75)
    );
BUF_X1_362: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(76),
        Z => S791(76)
    );
BUF_X1_363: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(77),
        Z => S791(77)
    );
BUF_X1_364: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(78),
        Z => S791(78)
    );
BUF_X1_365: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(79),
        Z => S791(79)
    );
BUF_X1_366: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(8),
        Z => S791(8)
    );
BUF_X1_367: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(80),
        Z => S791(80)
    );
BUF_X1_368: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(81),
        Z => S791(81)
    );
BUF_X1_369: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(82),
        Z => S791(82)
    );
BUF_X1_370: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(83),
        Z => S791(83)
    );
BUF_X1_371: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(84),
        Z => S791(84)
    );
BUF_X1_372: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(85),
        Z => S791(85)
    );
BUF_X1_373: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(86),
        Z => S791(86)
    );
BUF_X1_374: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(87),
        Z => S791(87)
    );
BUF_X1_375: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(88),
        Z => S791(88)
    );
BUF_X1_376: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(89),
        Z => S791(89)
    );
BUF_X1_377: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(9),
        Z => S791(9)
    );
BUF_X1_378: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(90),
        Z => S791(90)
    );
BUF_X1_379: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(91),
        Z => S791(91)
    );
BUF_X1_380: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(92),
        Z => S791(92)
    );
BUF_X1_381: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(93),
        Z => S791(93)
    );
BUF_X1_382: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(94),
        Z => S791(94)
    );
BUF_X1_383: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(95),
        Z => S791(95)
    );
BUF_X1_384: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(96),
        Z => S791(96)
    );
BUF_X1_385: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(97),
        Z => S791(97)
    );
BUF_X1_386: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(98),
        Z => S791(98)
    );
BUF_X1_387: ENTITY WORK.BUF_X1
    PORT MAP (
        A => expected128(99),
        Z => S791(99)
    );
BUF_X1_388: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(0),
        Z => S792(0)
    );
BUF_X1_389: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(1),
        Z => S792(1)
    );
BUF_X1_390: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(10),
        Z => S792(10)
    );
BUF_X1_391: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(100),
        Z => S792(100)
    );
BUF_X1_392: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(101),
        Z => S792(101)
    );
BUF_X1_393: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(102),
        Z => S792(102)
    );
BUF_X1_394: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(103),
        Z => S792(103)
    );
BUF_X1_395: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(104),
        Z => S792(104)
    );
BUF_X1_396: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(105),
        Z => S792(105)
    );
BUF_X1_397: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(106),
        Z => S792(106)
    );
BUF_X1_398: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(107),
        Z => S792(107)
    );
BUF_X1_399: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(108),
        Z => S792(108)
    );
BUF_X1_400: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(109),
        Z => S792(109)
    );
BUF_X1_401: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(11),
        Z => S792(11)
    );
BUF_X1_402: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(110),
        Z => S792(110)
    );
BUF_X1_403: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(111),
        Z => S792(111)
    );
BUF_X1_404: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(112),
        Z => S792(112)
    );
BUF_X1_405: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(113),
        Z => S792(113)
    );
BUF_X1_406: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(114),
        Z => S792(114)
    );
BUF_X1_407: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(115),
        Z => S792(115)
    );
BUF_X1_408: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(116),
        Z => S792(116)
    );
BUF_X1_409: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(117),
        Z => S792(117)
    );
BUF_X1_410: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(118),
        Z => S792(118)
    );
BUF_X1_411: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(119),
        Z => S792(119)
    );
BUF_X1_412: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(12),
        Z => S792(12)
    );
BUF_X1_413: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(120),
        Z => S792(120)
    );
BUF_X1_414: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(121),
        Z => S792(121)
    );
BUF_X1_415: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(122),
        Z => S792(122)
    );
BUF_X1_416: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(123),
        Z => S792(123)
    );
BUF_X1_417: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(124),
        Z => S792(124)
    );
BUF_X1_418: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(125),
        Z => S792(125)
    );
BUF_X1_419: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(126),
        Z => S792(126)
    );
BUF_X1_420: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(127),
        Z => S792(127)
    );
BUF_X1_421: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(13),
        Z => S792(13)
    );
BUF_X1_422: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(14),
        Z => S792(14)
    );
BUF_X1_423: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(15),
        Z => S792(15)
    );
BUF_X1_424: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(16),
        Z => S792(16)
    );
BUF_X1_425: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(17),
        Z => S792(17)
    );
BUF_X1_426: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(18),
        Z => S792(18)
    );
BUF_X1_427: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(19),
        Z => S792(19)
    );
BUF_X1_428: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(2),
        Z => S792(2)
    );
BUF_X1_429: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(20),
        Z => S792(20)
    );
BUF_X1_430: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(21),
        Z => S792(21)
    );
BUF_X1_431: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(22),
        Z => S792(22)
    );
BUF_X1_432: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(23),
        Z => S792(23)
    );
BUF_X1_433: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(24),
        Z => S792(24)
    );
BUF_X1_434: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(25),
        Z => S792(25)
    );
BUF_X1_435: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(26),
        Z => S792(26)
    );
BUF_X1_436: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(27),
        Z => S792(27)
    );
BUF_X1_437: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(28),
        Z => S792(28)
    );
BUF_X1_438: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(29),
        Z => S792(29)
    );
BUF_X1_439: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(3),
        Z => S792(3)
    );
BUF_X1_440: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(30),
        Z => S792(30)
    );
BUF_X1_441: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(31),
        Z => S792(31)
    );
BUF_X1_442: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(32),
        Z => S792(32)
    );
BUF_X1_443: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(33),
        Z => S792(33)
    );
BUF_X1_444: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(34),
        Z => S792(34)
    );
BUF_X1_445: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(35),
        Z => S792(35)
    );
BUF_X1_446: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(36),
        Z => S792(36)
    );
BUF_X1_447: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(37),
        Z => S792(37)
    );
BUF_X1_448: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(38),
        Z => S792(38)
    );
BUF_X1_449: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(39),
        Z => S792(39)
    );
BUF_X1_450: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(4),
        Z => S792(4)
    );
BUF_X1_451: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(40),
        Z => S792(40)
    );
BUF_X1_452: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(41),
        Z => S792(41)
    );
BUF_X1_453: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(42),
        Z => S792(42)
    );
BUF_X1_454: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(43),
        Z => S792(43)
    );
BUF_X1_455: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(44),
        Z => S792(44)
    );
BUF_X1_456: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(45),
        Z => S792(45)
    );
BUF_X1_457: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(46),
        Z => S792(46)
    );
BUF_X1_458: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(47),
        Z => S792(47)
    );
BUF_X1_459: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(48),
        Z => S792(48)
    );
BUF_X1_460: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(49),
        Z => S792(49)
    );
BUF_X1_461: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(5),
        Z => S792(5)
    );
BUF_X1_462: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(50),
        Z => S792(50)
    );
BUF_X1_463: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(51),
        Z => S792(51)
    );
BUF_X1_464: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(52),
        Z => S792(52)
    );
BUF_X1_465: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(53),
        Z => S792(53)
    );
BUF_X1_466: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(54),
        Z => S792(54)
    );
BUF_X1_467: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(55),
        Z => S792(55)
    );
BUF_X1_468: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(56),
        Z => S792(56)
    );
BUF_X1_469: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(57),
        Z => S792(57)
    );
BUF_X1_470: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(58),
        Z => S792(58)
    );
BUF_X1_471: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(59),
        Z => S792(59)
    );
BUF_X1_472: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(6),
        Z => S792(6)
    );
BUF_X1_473: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(60),
        Z => S792(60)
    );
BUF_X1_474: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(61),
        Z => S792(61)
    );
BUF_X1_475: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(62),
        Z => S792(62)
    );
BUF_X1_476: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(63),
        Z => S792(63)
    );
BUF_X1_477: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(64),
        Z => S792(64)
    );
BUF_X1_478: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(65),
        Z => S792(65)
    );
BUF_X1_479: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(66),
        Z => S792(66)
    );
BUF_X1_480: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(67),
        Z => S792(67)
    );
BUF_X1_481: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(68),
        Z => S792(68)
    );
BUF_X1_482: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(69),
        Z => S792(69)
    );
BUF_X1_483: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(7),
        Z => S792(7)
    );
BUF_X1_484: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(70),
        Z => S792(70)
    );
BUF_X1_485: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(71),
        Z => S792(71)
    );
BUF_X1_486: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(72),
        Z => S792(72)
    );
BUF_X1_487: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(73),
        Z => S792(73)
    );
BUF_X1_488: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(74),
        Z => S792(74)
    );
BUF_X1_489: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(75),
        Z => S792(75)
    );
BUF_X1_490: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(76),
        Z => S792(76)
    );
BUF_X1_491: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(77),
        Z => S792(77)
    );
BUF_X1_492: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(78),
        Z => S792(78)
    );
BUF_X1_493: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(79),
        Z => S792(79)
    );
BUF_X1_494: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(8),
        Z => S792(8)
    );
BUF_X1_495: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(80),
        Z => S792(80)
    );
BUF_X1_496: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(81),
        Z => S792(81)
    );
BUF_X1_497: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(82),
        Z => S792(82)
    );
BUF_X1_498: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(83),
        Z => S792(83)
    );
BUF_X1_499: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(84),
        Z => S792(84)
    );
BUF_X1_500: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(85),
        Z => S792(85)
    );
BUF_X1_501: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(86),
        Z => S792(86)
    );
BUF_X1_502: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(87),
        Z => S792(87)
    );
BUF_X1_503: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(88),
        Z => S792(88)
    );
BUF_X1_504: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(89),
        Z => S792(89)
    );
BUF_X1_505: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(9),
        Z => S792(9)
    );
BUF_X1_506: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(90),
        Z => S792(90)
    );
BUF_X1_507: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(91),
        Z => S792(91)
    );
BUF_X1_508: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(92),
        Z => S792(92)
    );
BUF_X1_509: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(93),
        Z => S792(93)
    );
BUF_X1_510: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(94),
        Z => S792(94)
    );
BUF_X1_511: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(95),
        Z => S792(95)
    );
BUF_X1_512: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(96),
        Z => S792(96)
    );
BUF_X1_513: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(97),
        Z => S792(97)
    );
BUF_X1_514: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(98),
        Z => S792(98)
    );
BUF_X1_515: ENTITY WORK.BUF_X1
    PORT MAP (
        A => in(99),
        Z => S792(99)
    );
BUF_X1_516: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(0),
        Z => S793(0)
    );
BUF_X1_517: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(1),
        Z => S793(1)
    );
BUF_X1_518: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(10),
        Z => S793(10)
    );
BUF_X1_519: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(100),
        Z => S793(100)
    );
BUF_X1_520: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(101),
        Z => S793(101)
    );
BUF_X1_521: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(102),
        Z => S793(102)
    );
BUF_X1_522: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(103),
        Z => S793(103)
    );
BUF_X1_523: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(104),
        Z => S793(104)
    );
BUF_X1_524: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(105),
        Z => S793(105)
    );
BUF_X1_525: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(106),
        Z => S793(106)
    );
BUF_X1_526: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(107),
        Z => S793(107)
    );
BUF_X1_527: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(108),
        Z => S793(108)
    );
BUF_X1_528: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(109),
        Z => S793(109)
    );
BUF_X1_529: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(11),
        Z => S793(11)
    );
BUF_X1_530: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(110),
        Z => S793(110)
    );
BUF_X1_531: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(111),
        Z => S793(111)
    );
BUF_X1_532: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(112),
        Z => S793(112)
    );
BUF_X1_533: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(113),
        Z => S793(113)
    );
BUF_X1_534: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(114),
        Z => S793(114)
    );
BUF_X1_535: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(115),
        Z => S793(115)
    );
BUF_X1_536: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(116),
        Z => S793(116)
    );
BUF_X1_537: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(117),
        Z => S793(117)
    );
BUF_X1_538: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(118),
        Z => S793(118)
    );
BUF_X1_539: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(119),
        Z => S793(119)
    );
BUF_X1_540: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(12),
        Z => S793(12)
    );
BUF_X1_541: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(120),
        Z => S793(120)
    );
BUF_X1_542: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(121),
        Z => S793(121)
    );
BUF_X1_543: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(122),
        Z => S793(122)
    );
BUF_X1_544: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(123),
        Z => S793(123)
    );
BUF_X1_545: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(124),
        Z => S793(124)
    );
BUF_X1_546: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(125),
        Z => S793(125)
    );
BUF_X1_547: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(126),
        Z => S793(126)
    );
BUF_X1_548: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(127),
        Z => S793(127)
    );
BUF_X1_549: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(13),
        Z => S793(13)
    );
BUF_X1_550: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(14),
        Z => S793(14)
    );
BUF_X1_551: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(15),
        Z => S793(15)
    );
BUF_X1_552: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(16),
        Z => S793(16)
    );
BUF_X1_553: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(17),
        Z => S793(17)
    );
BUF_X1_554: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(18),
        Z => S793(18)
    );
BUF_X1_555: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(19),
        Z => S793(19)
    );
BUF_X1_556: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(2),
        Z => S793(2)
    );
BUF_X1_557: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(20),
        Z => S793(20)
    );
BUF_X1_558: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(21),
        Z => S793(21)
    );
BUF_X1_559: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(22),
        Z => S793(22)
    );
BUF_X1_560: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(23),
        Z => S793(23)
    );
BUF_X1_561: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(24),
        Z => S793(24)
    );
BUF_X1_562: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(25),
        Z => S793(25)
    );
BUF_X1_563: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(26),
        Z => S793(26)
    );
BUF_X1_564: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(27),
        Z => S793(27)
    );
BUF_X1_565: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(28),
        Z => S793(28)
    );
BUF_X1_566: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(29),
        Z => S793(29)
    );
BUF_X1_567: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(3),
        Z => S793(3)
    );
BUF_X1_568: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(30),
        Z => S793(30)
    );
BUF_X1_569: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(31),
        Z => S793(31)
    );
BUF_X1_570: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(32),
        Z => S793(32)
    );
BUF_X1_571: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(33),
        Z => S793(33)
    );
BUF_X1_572: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(34),
        Z => S793(34)
    );
BUF_X1_573: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(35),
        Z => S793(35)
    );
BUF_X1_574: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(36),
        Z => S793(36)
    );
BUF_X1_575: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(37),
        Z => S793(37)
    );
BUF_X1_576: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(38),
        Z => S793(38)
    );
BUF_X1_577: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(39),
        Z => S793(39)
    );
BUF_X1_578: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(4),
        Z => S793(4)
    );
BUF_X1_579: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(40),
        Z => S793(40)
    );
BUF_X1_580: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(41),
        Z => S793(41)
    );
BUF_X1_581: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(42),
        Z => S793(42)
    );
BUF_X1_582: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(43),
        Z => S793(43)
    );
BUF_X1_583: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(44),
        Z => S793(44)
    );
BUF_X1_584: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(45),
        Z => S793(45)
    );
BUF_X1_585: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(46),
        Z => S793(46)
    );
BUF_X1_586: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(47),
        Z => S793(47)
    );
BUF_X1_587: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(48),
        Z => S793(48)
    );
BUF_X1_588: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(49),
        Z => S793(49)
    );
BUF_X1_589: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(5),
        Z => S793(5)
    );
BUF_X1_590: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(50),
        Z => S793(50)
    );
BUF_X1_591: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(51),
        Z => S793(51)
    );
BUF_X1_592: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(52),
        Z => S793(52)
    );
BUF_X1_593: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(53),
        Z => S793(53)
    );
BUF_X1_594: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(54),
        Z => S793(54)
    );
BUF_X1_595: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(55),
        Z => S793(55)
    );
BUF_X1_596: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(56),
        Z => S793(56)
    );
BUF_X1_597: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(57),
        Z => S793(57)
    );
BUF_X1_598: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(58),
        Z => S793(58)
    );
BUF_X1_599: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(59),
        Z => S793(59)
    );
BUF_X1_600: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(6),
        Z => S793(6)
    );
BUF_X1_601: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(60),
        Z => S793(60)
    );
BUF_X1_602: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(61),
        Z => S793(61)
    );
BUF_X1_603: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(62),
        Z => S793(62)
    );
BUF_X1_604: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(63),
        Z => S793(63)
    );
BUF_X1_605: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(64),
        Z => S793(64)
    );
BUF_X1_606: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(65),
        Z => S793(65)
    );
BUF_X1_607: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(66),
        Z => S793(66)
    );
BUF_X1_608: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(67),
        Z => S793(67)
    );
BUF_X1_609: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(68),
        Z => S793(68)
    );
BUF_X1_610: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(69),
        Z => S793(69)
    );
BUF_X1_611: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(7),
        Z => S793(7)
    );
BUF_X1_612: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(70),
        Z => S793(70)
    );
BUF_X1_613: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(71),
        Z => S793(71)
    );
BUF_X1_614: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(72),
        Z => S793(72)
    );
BUF_X1_615: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(73),
        Z => S793(73)
    );
BUF_X1_616: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(74),
        Z => S793(74)
    );
BUF_X1_617: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(75),
        Z => S793(75)
    );
BUF_X1_618: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(76),
        Z => S793(76)
    );
BUF_X1_619: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(77),
        Z => S793(77)
    );
BUF_X1_620: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(78),
        Z => S793(78)
    );
BUF_X1_621: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(79),
        Z => S793(79)
    );
BUF_X1_622: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(8),
        Z => S793(8)
    );
BUF_X1_623: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(80),
        Z => S793(80)
    );
BUF_X1_624: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(81),
        Z => S793(81)
    );
BUF_X1_625: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(82),
        Z => S793(82)
    );
BUF_X1_626: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(83),
        Z => S793(83)
    );
BUF_X1_627: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(84),
        Z => S793(84)
    );
BUF_X1_628: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(85),
        Z => S793(85)
    );
BUF_X1_629: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(86),
        Z => S793(86)
    );
BUF_X1_630: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(87),
        Z => S793(87)
    );
BUF_X1_631: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(88),
        Z => S793(88)
    );
BUF_X1_632: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(89),
        Z => S793(89)
    );
BUF_X1_633: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(9),
        Z => S793(9)
    );
BUF_X1_634: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(90),
        Z => S793(90)
    );
BUF_X1_635: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(91),
        Z => S793(91)
    );
BUF_X1_636: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(92),
        Z => S793(92)
    );
BUF_X1_637: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(93),
        Z => S793(93)
    );
BUF_X1_638: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(94),
        Z => S793(94)
    );
BUF_X1_639: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(95),
        Z => S793(95)
    );
BUF_X1_640: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(96),
        Z => S793(96)
    );
BUF_X1_641: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(97),
        Z => S793(97)
    );
BUF_X1_642: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(98),
        Z => S793(98)
    );
BUF_X1_643: ENTITY WORK.BUF_X1
    PORT MAP (
        A => key128(99),
        Z => S793(99)
    );
AES_Encrypt_1: ENTITY WORK.AES_Encrypt
    PORT MAP (
        in(0) => S792(0),
        in(1) => S792(1),
        in(2) => S792(2),
        in(3) => S792(3),
        in(4) => S792(4),
        in(5) => S792(5),
        in(6) => S792(6),
        in(7) => S792(7),
        in(8) => S792(8),
        in(9) => S792(9),
        in(10) => S792(10),
        in(11) => S792(11),
        in(12) => S792(12),
        in(13) => S792(13),
        in(14) => S792(14),
        in(15) => S792(15),
        in(16) => S792(16),
        in(17) => S792(17),
        in(18) => S792(18),
        in(19) => S792(19),
        in(20) => S792(20),
        in(21) => S792(21),
        in(22) => S792(22),
        in(23) => S792(23),
        in(24) => S792(24),
        in(25) => S792(25),
        in(26) => S792(26),
        in(27) => S792(27),
        in(28) => S792(28),
        in(29) => S792(29),
        in(30) => S792(30),
        in(31) => S792(31),
        in(32) => S792(32),
        in(33) => S792(33),
        in(34) => S792(34),
        in(35) => S792(35),
        in(36) => S792(36),
        in(37) => S792(37),
        in(38) => S792(38),
        in(39) => S792(39),
        in(40) => S792(40),
        in(41) => S792(41),
        in(42) => S792(42),
        in(43) => S792(43),
        in(44) => S792(44),
        in(45) => S792(45),
        in(46) => S792(46),
        in(47) => S792(47),
        in(48) => S792(48),
        in(49) => S792(49),
        in(50) => S792(50),
        in(51) => S792(51),
        in(52) => S792(52),
        in(53) => S792(53),
        in(54) => S792(54),
        in(55) => S792(55),
        in(56) => S792(56),
        in(57) => S792(57),
        in(58) => S792(58),
        in(59) => S792(59),
        in(60) => S792(60),
        in(61) => S792(61),
        in(62) => S792(62),
        in(63) => S792(63),
        in(64) => S792(64),
        in(65) => S792(65),
        in(66) => S792(66),
        in(67) => S792(67),
        in(68) => S792(68),
        in(69) => S792(69),
        in(70) => S792(70),
        in(71) => S792(71),
        in(72) => S792(72),
        in(73) => S792(73),
        in(74) => S792(74),
        in(75) => S792(75),
        in(76) => S792(76),
        in(77) => S792(77),
        in(78) => S792(78),
        in(79) => S792(79),
        in(80) => S792(80),
        in(81) => S792(81),
        in(82) => S792(82),
        in(83) => S792(83),
        in(84) => S792(84),
        in(85) => S792(85),
        in(86) => S792(86),
        in(87) => S792(87),
        in(88) => S792(88),
        in(89) => S792(89),
        in(90) => S792(90),
        in(91) => S792(91),
        in(92) => S792(92),
        in(93) => S792(93),
        in(94) => S792(94),
        in(95) => S792(95),
        in(96) => S792(96),
        in(97) => S792(97),
        in(98) => S792(98),
        in(99) => S792(99),
        in(100) => S792(100),
        in(101) => S792(101),
        in(102) => S792(102),
        in(103) => S792(103),
        in(104) => S792(104),
        in(105) => S792(105),
        in(106) => S792(106),
        in(107) => S792(107),
        in(108) => S792(108),
        in(109) => S792(109),
        in(110) => S792(110),
        in(111) => S792(111),
        in(112) => S792(112),
        in(113) => S792(113),
        in(114) => S792(114),
        in(115) => S792(115),
        in(116) => S792(116),
        in(117) => S792(117),
        in(118) => S792(118),
        in(119) => S792(119),
        in(120) => S792(120),
        in(121) => S792(121),
        in(122) => S792(122),
        in(123) => S792(123),
        in(124) => S792(124),
        in(125) => S792(125),
        in(126) => S792(126),
        in(127) => S792(127),
        key(0) => S793(0),
        key(1) => S793(1),
        key(2) => S793(2),
        key(3) => S793(3),
        key(4) => S793(4),
        key(5) => S793(5),
        key(6) => S793(6),
        key(7) => S793(7),
        key(8) => S793(8),
        key(9) => S793(9),
        key(10) => S793(10),
        key(11) => S793(11),
        key(12) => S793(12),
        key(13) => S793(13),
        key(14) => S793(14),
        key(15) => S793(15),
        key(16) => S793(16),
        key(17) => S793(17),
        key(18) => S793(18),
        key(19) => S793(19),
        key(20) => S793(20),
        key(21) => S793(21),
        key(22) => S793(22),
        key(23) => S793(23),
        key(24) => S793(24),
        key(25) => S793(25),
        key(26) => S793(26),
        key(27) => S793(27),
        key(28) => S793(28),
        key(29) => S793(29),
        key(30) => S793(30),
        key(31) => S793(31),
        key(32) => S793(32),
        key(33) => S793(33),
        key(34) => S793(34),
        key(35) => S793(35),
        key(36) => S793(36),
        key(37) => S793(37),
        key(38) => S793(38),
        key(39) => S793(39),
        key(40) => S793(40),
        key(41) => S793(41),
        key(42) => S793(42),
        key(43) => S793(43),
        key(44) => S793(44),
        key(45) => S793(45),
        key(46) => S793(46),
        key(47) => S793(47),
        key(48) => S793(48),
        key(49) => S793(49),
        key(50) => S793(50),
        key(51) => S793(51),
        key(52) => S793(52),
        key(53) => S793(53),
        key(54) => S793(54),
        key(55) => S793(55),
        key(56) => S793(56),
        key(57) => S793(57),
        key(58) => S793(58),
        key(59) => S793(59),
        key(60) => S793(60),
        key(61) => S793(61),
        key(62) => S793(62),
        key(63) => S793(63),
        key(64) => S793(64),
        key(65) => S793(65),
        key(66) => S793(66),
        key(67) => S793(67),
        key(68) => S793(68),
        key(69) => S793(69),
        key(70) => S793(70),
        key(71) => S793(71),
        key(72) => S793(72),
        key(73) => S793(73),
        key(74) => S793(74),
        key(75) => S793(75),
        key(76) => S793(76),
        key(77) => S793(77),
        key(78) => S793(78),
        key(79) => S793(79),
        key(80) => S793(80),
        key(81) => S793(81),
        key(82) => S793(82),
        key(83) => S793(83),
        key(84) => S793(84),
        key(85) => S793(85),
        key(86) => S793(86),
        key(87) => S793(87),
        key(88) => S793(88),
        key(89) => S793(89),
        key(90) => S793(90),
        key(91) => S793(91),
        key(92) => S793(92),
        key(93) => S793(93),
        key(94) => S793(94),
        key(95) => S793(95),
        key(96) => S793(96),
        key(97) => S793(97),
        key(98) => S793(98),
        key(99) => S793(99),
        key(100) => S793(100),
        key(101) => S793(101),
        key(102) => S793(102),
        key(103) => S793(103),
        key(104) => S793(104),
        key(105) => S793(105),
        key(106) => S793(106),
        key(107) => S793(107),
        key(108) => S793(108),
        key(109) => S793(109),
        key(110) => S793(110),
        key(111) => S793(111),
        key(112) => S793(112),
        key(113) => S793(113),
        key(114) => S793(114),
        key(115) => S793(115),
        key(116) => S793(116),
        key(117) => S793(117),
        key(118) => S793(118),
        key(119) => S793(119),
        key(120) => S793(120),
        key(121) => S793(121),
        key(122) => S793(122),
        key(123) => S793(123),
        key(124) => S793(124),
        key(125) => S793(125),
        key(126) => S793(126),
        key(127) => S793(127),
        out(0) => S790(0),
        out(1) => S790(1),
        out(2) => S790(2),
        out(3) => S790(3),
        out(4) => S790(4),
        out(5) => S790(5),
        out(6) => S790(6),
        out(7) => S790(7),
        out(8) => S790(8),
        out(9) => S790(9),
        out(10) => S790(10),
        out(11) => S790(11),
        out(12) => S790(12),
        out(13) => S790(13),
        out(14) => S790(14),
        out(15) => S790(15),
        out(16) => S790(16),
        out(17) => S790(17),
        out(18) => S790(18),
        out(19) => S790(19),
        out(20) => S790(20),
        out(21) => S790(21),
        out(22) => S790(22),
        out(23) => S790(23),
        out(24) => S790(24),
        out(25) => S790(25),
        out(26) => S790(26),
        out(27) => S790(27),
        out(28) => S790(28),
        out(29) => S790(29),
        out(30) => S790(30),
        out(31) => S790(31),
        out(32) => S790(32),
        out(33) => S790(33),
        out(34) => S790(34),
        out(35) => S790(35),
        out(36) => S790(36),
        out(37) => S790(37),
        out(38) => S790(38),
        out(39) => S790(39),
        out(40) => S790(40),
        out(41) => S790(41),
        out(42) => S790(42),
        out(43) => S790(43),
        out(44) => S790(44),
        out(45) => S790(45),
        out(46) => S790(46),
        out(47) => S790(47),
        out(48) => S790(48),
        out(49) => S790(49),
        out(50) => S790(50),
        out(51) => S790(51),
        out(52) => S790(52),
        out(53) => S790(53),
        out(54) => S790(54),
        out(55) => S790(55),
        out(56) => S790(56),
        out(57) => S790(57),
        out(58) => S790(58),
        out(59) => S790(59),
        out(60) => S790(60),
        out(61) => S790(61),
        out(62) => S790(62),
        out(63) => S790(63),
        out(64) => S790(64),
        out(65) => S790(65),
        out(66) => S790(66),
        out(67) => S790(67),
        out(68) => S790(68),
        out(69) => S790(69),
        out(70) => S790(70),
        out(71) => S790(71),
        out(72) => S790(72),
        out(73) => S790(73),
        out(74) => S790(74),
        out(75) => S790(75),
        out(76) => S790(76),
        out(77) => S790(77),
        out(78) => S790(78),
        out(79) => S790(79),
        out(80) => S790(80),
        out(81) => S790(81),
        out(82) => S790(82),
        out(83) => S790(83),
        out(84) => S790(84),
        out(85) => S790(85),
        out(86) => S790(86),
        out(87) => S790(87),
        out(88) => S790(88),
        out(89) => S790(89),
        out(90) => S790(90),
        out(91) => S790(91),
        out(92) => S790(92),
        out(93) => S790(93),
        out(94) => S790(94),
        out(95) => S790(95),
        out(96) => S790(96),
        out(97) => S790(97),
        out(98) => S790(98),
        out(99) => S790(99),
        out(100) => S790(100),
        out(101) => S790(101),
        out(102) => S790(102),
        out(103) => S790(103),
        out(104) => S790(104),
        out(105) => S790(105),
        out(106) => S790(106),
        out(107) => S790(107),
        out(108) => S790(108),
        out(109) => S790(109),
        out(110) => S790(110),
        out(111) => S790(111),
        out(112) => S790(112),
        out(113) => S790(113),
        out(114) => S790(114),
        out(115) => S790(115),
        out(116) => S790(116),
        out(117) => S790(117),
        out(118) => S790(118),
        out(119) => S790(119),
        out(120) => S790(120),
        out(121) => S790(121),
        out(122) => S790(122),
        out(123) => S790(123),
        out(124) => S790(124),
        out(125) => S790(125),
        out(126) => S790(126),
        out(127) => S790(127)
    );
AES_Decrypt_1: ENTITY WORK.AES_Decrypt
    PORT MAP (
        in(0) => S790(0),
        in(1) => S790(1),
        in(2) => S790(2),
        in(3) => S790(3),
        in(4) => S790(4),
        in(5) => S790(5),
        in(6) => S790(6),
        in(7) => S790(7),
        in(8) => S790(8),
        in(9) => S790(9),
        in(10) => S790(10),
        in(11) => S790(11),
        in(12) => S790(12),
        in(13) => S790(13),
        in(14) => S790(14),
        in(15) => S790(15),
        in(16) => S790(16),
        in(17) => S790(17),
        in(18) => S790(18),
        in(19) => S790(19),
        in(20) => S790(20),
        in(21) => S790(21),
        in(22) => S790(22),
        in(23) => S790(23),
        in(24) => S790(24),
        in(25) => S790(25),
        in(26) => S790(26),
        in(27) => S790(27),
        in(28) => S790(28),
        in(29) => S790(29),
        in(30) => S790(30),
        in(31) => S790(31),
        in(32) => S790(32),
        in(33) => S790(33),
        in(34) => S790(34),
        in(35) => S790(35),
        in(36) => S790(36),
        in(37) => S790(37),
        in(38) => S790(38),
        in(39) => S790(39),
        in(40) => S790(40),
        in(41) => S790(41),
        in(42) => S790(42),
        in(43) => S790(43),
        in(44) => S790(44),
        in(45) => S790(45),
        in(46) => S790(46),
        in(47) => S790(47),
        in(48) => S790(48),
        in(49) => S790(49),
        in(50) => S790(50),
        in(51) => S790(51),
        in(52) => S790(52),
        in(53) => S790(53),
        in(54) => S790(54),
        in(55) => S790(55),
        in(56) => S790(56),
        in(57) => S790(57),
        in(58) => S790(58),
        in(59) => S790(59),
        in(60) => S790(60),
        in(61) => S790(61),
        in(62) => S790(62),
        in(63) => S790(63),
        in(64) => S790(64),
        in(65) => S790(65),
        in(66) => S790(66),
        in(67) => S790(67),
        in(68) => S790(68),
        in(69) => S790(69),
        in(70) => S790(70),
        in(71) => S790(71),
        in(72) => S790(72),
        in(73) => S790(73),
        in(74) => S790(74),
        in(75) => S790(75),
        in(76) => S790(76),
        in(77) => S790(77),
        in(78) => S790(78),
        in(79) => S790(79),
        in(80) => S790(80),
        in(81) => S790(81),
        in(82) => S790(82),
        in(83) => S790(83),
        in(84) => S790(84),
        in(85) => S790(85),
        in(86) => S790(86),
        in(87) => S790(87),
        in(88) => S790(88),
        in(89) => S790(89),
        in(90) => S790(90),
        in(91) => S790(91),
        in(92) => S790(92),
        in(93) => S790(93),
        in(94) => S790(94),
        in(95) => S790(95),
        in(96) => S790(96),
        in(97) => S790(97),
        in(98) => S790(98),
        in(99) => S790(99),
        in(100) => S790(100),
        in(101) => S790(101),
        in(102) => S790(102),
        in(103) => S790(103),
        in(104) => S790(104),
        in(105) => S790(105),
        in(106) => S790(106),
        in(107) => S790(107),
        in(108) => S790(108),
        in(109) => S790(109),
        in(110) => S790(110),
        in(111) => S790(111),
        in(112) => S790(112),
        in(113) => S790(113),
        in(114) => S790(114),
        in(115) => S790(115),
        in(116) => S790(116),
        in(117) => S790(117),
        in(118) => S790(118),
        in(119) => S790(119),
        in(120) => S790(120),
        in(121) => S790(121),
        in(122) => S790(122),
        in(123) => S790(123),
        in(124) => S790(124),
        in(125) => S790(125),
        in(126) => S790(126),
        in(127) => S790(127),
        key(0) => S793(0),
        key(1) => S793(1),
        key(2) => S793(2),
        key(3) => S793(3),
        key(4) => S793(4),
        key(5) => S793(5),
        key(6) => S793(6),
        key(7) => S793(7),
        key(8) => S793(8),
        key(9) => S793(9),
        key(10) => S793(10),
        key(11) => S793(11),
        key(12) => S793(12),
        key(13) => S793(13),
        key(14) => S793(14),
        key(15) => S793(15),
        key(16) => S793(16),
        key(17) => S793(17),
        key(18) => S793(18),
        key(19) => S793(19),
        key(20) => S793(20),
        key(21) => S793(21),
        key(22) => S793(22),
        key(23) => S793(23),
        key(24) => S793(24),
        key(25) => S793(25),
        key(26) => S793(26),
        key(27) => S793(27),
        key(28) => S793(28),
        key(29) => S793(29),
        key(30) => S793(30),
        key(31) => S793(31),
        key(32) => S793(32),
        key(33) => S793(33),
        key(34) => S793(34),
        key(35) => S793(35),
        key(36) => S793(36),
        key(37) => S793(37),
        key(38) => S793(38),
        key(39) => S793(39),
        key(40) => S793(40),
        key(41) => S793(41),
        key(42) => S793(42),
        key(43) => S793(43),
        key(44) => S793(44),
        key(45) => S793(45),
        key(46) => S793(46),
        key(47) => S793(47),
        key(48) => S793(48),
        key(49) => S793(49),
        key(50) => S793(50),
        key(51) => S793(51),
        key(52) => S793(52),
        key(53) => S793(53),
        key(54) => S793(54),
        key(55) => S793(55),
        key(56) => S793(56),
        key(57) => S793(57),
        key(58) => S793(58),
        key(59) => S793(59),
        key(60) => S793(60),
        key(61) => S793(61),
        key(62) => S793(62),
        key(63) => S793(63),
        key(64) => S793(64),
        key(65) => S793(65),
        key(66) => S793(66),
        key(67) => S793(67),
        key(68) => S793(68),
        key(69) => S793(69),
        key(70) => S793(70),
        key(71) => S793(71),
        key(72) => S793(72),
        key(73) => S793(73),
        key(74) => S793(74),
        key(75) => S793(75),
        key(76) => S793(76),
        key(77) => S793(77),
        key(78) => S793(78),
        key(79) => S793(79),
        key(80) => S793(80),
        key(81) => S793(81),
        key(82) => S793(82),
        key(83) => S793(83),
        key(84) => S793(84),
        key(85) => S793(85),
        key(86) => S793(86),
        key(87) => S793(87),
        key(88) => S793(88),
        key(89) => S793(89),
        key(90) => S793(90),
        key(91) => S793(91),
        key(92) => S793(92),
        key(93) => S793(93),
        key(94) => S793(94),
        key(95) => S793(95),
        key(96) => S793(96),
        key(97) => S793(97),
        key(98) => S793(98),
        key(99) => S793(99),
        key(100) => S793(100),
        key(101) => S793(101),
        key(102) => S793(102),
        key(103) => S793(103),
        key(104) => S793(104),
        key(105) => S793(105),
        key(106) => S793(106),
        key(107) => S793(107),
        key(108) => S793(108),
        key(109) => S793(109),
        key(110) => S793(110),
        key(111) => S793(111),
        key(112) => S793(112),
        key(113) => S793(113),
        key(114) => S793(114),
        key(115) => S793(115),
        key(116) => S793(116),
        key(117) => S793(117),
        key(118) => S793(118),
        key(119) => S793(119),
        key(120) => S793(120),
        key(121) => S793(121),
        key(122) => S793(122),
        key(123) => S793(123),
        key(124) => S793(124),
        key(125) => S793(125),
        key(126) => S793(126),
        key(127) => S793(127),
        out(0) => S787(0),
        out(1) => S787(1),
        out(2) => S787(2),
        out(3) => S787(3),
        out(4) => S787(4),
        out(5) => S787(5),
        out(6) => S787(6),
        out(7) => S787(7),
        out(8) => S787(8),
        out(9) => S787(9),
        out(10) => S787(10),
        out(11) => S787(11),
        out(12) => S787(12),
        out(13) => S787(13),
        out(14) => S787(14),
        out(15) => S787(15),
        out(16) => S787(16),
        out(17) => S787(17),
        out(18) => S787(18),
        out(19) => S787(19),
        out(20) => S787(20),
        out(21) => S787(21),
        out(22) => S787(22),
        out(23) => S787(23),
        out(24) => S787(24),
        out(25) => S787(25),
        out(26) => S787(26),
        out(27) => S787(27),
        out(28) => S787(28),
        out(29) => S787(29),
        out(30) => S787(30),
        out(31) => S787(31),
        out(32) => S787(32),
        out(33) => S787(33),
        out(34) => S787(34),
        out(35) => S787(35),
        out(36) => S787(36),
        out(37) => S787(37),
        out(38) => S787(38),
        out(39) => S787(39),
        out(40) => S787(40),
        out(41) => S787(41),
        out(42) => S787(42),
        out(43) => S787(43),
        out(44) => S787(44),
        out(45) => S787(45),
        out(46) => S787(46),
        out(47) => S787(47),
        out(48) => S787(48),
        out(49) => S787(49),
        out(50) => S787(50),
        out(51) => S787(51),
        out(52) => S787(52),
        out(53) => S787(53),
        out(54) => S787(54),
        out(55) => S787(55),
        out(56) => S787(56),
        out(57) => S787(57),
        out(58) => S787(58),
        out(59) => S787(59),
        out(60) => S787(60),
        out(61) => S787(61),
        out(62) => S787(62),
        out(63) => S787(63),
        out(64) => S787(64),
        out(65) => S787(65),
        out(66) => S787(66),
        out(67) => S787(67),
        out(68) => S787(68),
        out(69) => S787(69),
        out(70) => S787(70),
        out(71) => S787(71),
        out(72) => S787(72),
        out(73) => S787(73),
        out(74) => S787(74),
        out(75) => S787(75),
        out(76) => S787(76),
        out(77) => S787(77),
        out(78) => S787(78),
        out(79) => S787(79),
        out(80) => S787(80),
        out(81) => S787(81),
        out(82) => S787(82),
        out(83) => S787(83),
        out(84) => S787(84),
        out(85) => S787(85),
        out(86) => S787(86),
        out(87) => S787(87),
        out(88) => S787(88),
        out(89) => S787(89),
        out(90) => S787(90),
        out(91) => S787(91),
        out(92) => S787(92),
        out(93) => S787(93),
        out(94) => S787(94),
        out(95) => S787(95),
        out(96) => S787(96),
        out(97) => S787(97),
        out(98) => S787(98),
        out(99) => S787(99),
        out(100) => S787(100),
        out(101) => S787(101),
        out(102) => S787(102),
        out(103) => S787(103),
        out(104) => S787(104),
        out(105) => S787(105),
        out(106) => S787(106),
        out(107) => S787(107),
        out(108) => S787(108),
        out(109) => S787(109),
        out(110) => S787(110),
        out(111) => S787(111),
        out(112) => S787(112),
        out(113) => S787(113),
        out(114) => S787(114),
        out(115) => S787(115),
        out(116) => S787(116),
        out(117) => S787(117),
        out(118) => S787(118),
        out(119) => S787(119),
        out(120) => S787(120),
        out(121) => S787(121),
        out(122) => S787(122),
        out(123) => S787(123),
        out(124) => S787(124),
        out(125) => S787(125),
        out(126) => S787(126),
        out(127) => S787(127)
    );

END ARCHITECTURE arch;
