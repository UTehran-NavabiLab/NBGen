`timescale 1ns/1ps

module C432_tb;
 
	reg [35:0]IN_Vector=36'd0;
	wire out223, out329, out370, out421, out430, out431, out432;

    initial begin
		#10  IN_Vector=35'b 111111111011111111011111111011111111;
		#10  IN_Vector=35'b 111111111101111111101111111101111111;
		#10  IN_Vector=35'b 111111111110111111110111111110111111;
		#10  IN_Vector=35'b 111111111111011111111011111111011111;
		#10  IN_Vector=35'b 111111111111101111111101111111101111;
		#10  IN_Vector=35'b 111111111111110111111110111111110111;
		#10  IN_Vector=35'b 111111111111111011111111011111111011;
		#10  IN_Vector=35'b 111111111111111101111111101111111101;
		#10  IN_Vector=35'b 111111111111111110111111110111111110;
		#10  IN_Vector=35'b 111111111111111111010011111101111111;
		#10  IN_Vector=35'b 111111111111111111101111111010000000;
		#10  IN_Vector=35'b 111111111111111111110110101111111111;
		#10  IN_Vector=35'b 111111111111111111111010111111111111;
		#10  IN_Vector=35'b 111111111111111111111100111111111111;
		#10  IN_Vector=35'b 111111111111111111111110111111111111;
		#10  IN_Vector=35'b 111111111111111111111111011111111111;
		#10  IN_Vector=35'b 111111111111111111111111101111111111;
		#10  IN_Vector=35'b 111111111111111111111111110111111111;
		#10  IN_Vector=35'b 111111111111111111111111111011111111;
		#10  IN_Vector=35'b 111111111111111111111111111101111111;
		#10  IN_Vector=35'b 111111111111111111111111111110111111;
		#10  IN_Vector=35'b 111111111111111111111111111111011111;
		#10  IN_Vector=35'b 111111111111111111111111111111101111;
		#10  IN_Vector=35'b 111111111111111111111111111111110111;
		#10  IN_Vector=35'b 111111111111111111111111111111111011;
		#10  IN_Vector=35'b 100000010100000010100000010100000000;
		#10  IN_Vector=35'b 011111101011111101011111101011111100;
		#10  IN_Vector=35'b 111111111111011011000100100000100100;
		#10  IN_Vector=35'b 111111111111101001111111111111111111;
		#10  IN_Vector=35'b 111111111011111111100000000100000000;
		#10  IN_Vector=35'b 111111111001111111111111111001111111;
		#10  IN_Vector=35'b 000000000000000000000000000000000000;
	end
    Circuit432  UUT( IN_Vector[35], IN_Vector[34], IN_Vector[33],
	IN_Vector[32], IN_Vector[31], IN_Vector[30], IN_Vector[29], IN_Vector[28], IN_Vector[27],
	IN_Vector[26], IN_Vector[25], IN_Vector[24], IN_Vector[23], IN_Vector[22], IN_Vector[21],
	IN_Vector[20], IN_Vector[19], IN_Vector[18], IN_Vector[17], IN_Vector[16], IN_Vector[15],
	IN_Vector[14], IN_Vector[13], IN_Vector[12], IN_Vector[11], IN_Vector[10], IN_Vector[9],
	IN_Vector[8], IN_Vector[7], IN_Vector[6], IN_Vector[5], IN_Vector[4], IN_Vector[3], IN_Vector[2],
	IN_Vector[1], IN_Vector[0], out223, out329, out370, out421, out430, out431, out432);

endmodule