module counter(clk, rst, en, co, counter);

wire S0;
wire S1;
wire S2;
wire S3;
wire S4;
wire S5;
wire S6;
wire S7;
wire S8;
wire S9;
wire S10;
wire S11;
wire S12;
wire S13;
wire S14;
wire S15;
wire S16;
wire S17;
wire S18;
wire S19;
wire S20;
wire S21;
wire S22;
wire S23;
wire S24;
wire S25;
wire new_counter_reg_0;
wire new_counter_reg_1;
wire new_counter_reg_2;
wire new_counter_reg_3;
input clk;
input rst;
input en;
output co;
output [3:0] counter;
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_0_ (
  .in({ new_counter_reg_0 }),
  .out({ S4 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1_ (
  .in({ new_counter_reg_3 }),
  .out({ S5 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2_ (
  .in({ S20 }),
  .out({ S6 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3_ (
  .in({ new_counter_reg_1, new_counter_reg_0 }),
  .out({ S7 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4_ (
  .in({ new_counter_reg_2, new_counter_reg_3 }),
  .out({ S8 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5_ (
  .in({ S8, S7 }),
  .out({ S19 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6_ (
  .in({ S6, S4 }),
  .out({ S9 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_7_ (
  .in({ S20, new_counter_reg_0 }),
  .out({ S10 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_8_ (
  .in({ S10, S9 }),
  .out({ S0 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_9_ (
  .in({ S7, S6 }),
  .out({ S11 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_10_ (
  .in({ S9, new_counter_reg_1 }),
  .out({ S12 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_11_ (
  .in({ S12, S11 }),
  .out({ S1 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_12_ (
  .in({ S11, new_counter_reg_2 }),
  .out({ S13 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_13_ (
  .in({ S13 }),
  .out({ S14 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_14_ (
  .in({ S11, new_counter_reg_2 }),
  .out({ S15 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_15_ (
  .in({ S15, S14 }),
  .out({ S2 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_16_ (
  .in({ S14, new_counter_reg_3 }),
  .out({ S16 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_17_ (
  .in({ S13, S5 }),
  .out({ S17 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_18_ (
  .in({ S17, S16 }),
  .out({ S3 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_19_ (
  .C({ S18 }),
  .CE({ 1'b1 }),
  .CLR({ S21 }),
  .D({ S0 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_counter_reg_0 }),
  .Si({ S22 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_20_ (
  .C({ S18 }),
  .CE({ 1'b1 }),
  .CLR({ S21 }),
  .D({ S1 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_counter_reg_1 }),
  .Si({ S23 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_21_ (
  .C({ S18 }),
  .CE({ 1'b1 }),
  .CLR({ S21 }),
  .D({ S2 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_counter_reg_2 }),
  .Si({ S24 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_22_ (
  .C({ S18 }),
  .CE({ 1'b1 }),
  .CLR({ S21 }),
  .D({ S3 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_counter_reg_3 }),
  .Si({ S25 }),
  .global_reset({ 1'b0 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_23_ (
  .in({ clk }),
  .out({ S18 })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_24_ (
  .in({ S19 }),
  .out({ co })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_25_ (
  .in({ new_counter_reg_0 }),
  .out({ counter[0] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_26_ (
  .in({ new_counter_reg_1 }),
  .out({ counter[1] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_27_ (
  .in({ new_counter_reg_2 }),
  .out({ counter[2] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_28_ (
  .in({ new_counter_reg_3 }),
  .out({ counter[3] })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_29_ (
  .in({ en }),
  .out({ S20 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_30_ (
  .in({ rst }),
  .out({ S21 })
);

endmodule