module PUNEH_Top_Module(clk, rst, writeMEM, readMEM, dataBus_in, dataBus_out, addrBus);

wire S0;
wire S1;
wire S2;
wire S3;
wire S4;
wire S5;
wire S6;
wire S7;
wire S8;
wire S9;
wire S10;
wire S11;
wire S12;
wire S13;
wire S14;
wire S15;
wire S16;
wire S17;
wire S18;
wire S19;
wire S20;
wire S21;
wire S22;
wire S23;
wire S24;
wire S25;
wire S26;
wire S27;
wire S28;
wire S29;
wire S30;
wire S31;
wire S32;
wire S33;
wire S34;
wire S35;
wire S36;
wire S37;
wire S38;
wire S39;
wire S40;
wire S41;
wire S42;
wire S43;
wire S44;
wire S45;
wire S46;
wire S47;
wire S48;
wire S49;
wire S50;
wire S51;
wire S52;
wire S53;
wire S54;
wire S55;
wire S56;
wire S57;
wire S58;
wire S59;
wire S60;
wire S61;
wire S62;
wire S63;
wire S64;
wire S65;
wire S66;
wire S67;
wire S68;
wire S69;
wire S70;
wire S71;
wire S72;
wire S73;
wire S74;
wire S75;
wire S76;
wire S77;
wire S78;
wire S79;
wire S80;
wire S81;
wire S82;
wire S83;
wire S84;
wire S85;
wire S86;
wire S87;
wire S88;
wire S89;
wire S90;
wire S91;
wire S92;
wire S93;
wire S94;
wire S95;
wire S96;
wire S97;
wire S98;
wire S99;
wire S100;
wire S101;
wire S102;
wire S103;
wire S104;
wire S105;
wire S106;
wire S107;
wire S108;
wire S109;
wire S110;
wire S111;
wire S112;
wire S113;
wire S114;
wire S115;
wire S116;
wire S117;
wire S118;
wire S119;
wire S120;
wire S121;
wire S122;
wire S123;
wire S124;
wire S125;
wire S126;
wire S127;
wire S128;
wire S129;
wire S130;
wire S131;
wire S132;
wire S133;
wire S134;
wire S135;
wire S136;
wire S137;
wire S138;
wire S139;
wire S140;
wire S141;
wire S142;
wire S143;
wire S144;
wire S145;
wire S146;
wire S147;
wire S148;
wire S149;
wire S150;
wire S151;
wire S152;
wire S153;
wire S154;
wire S155;
wire S156;
wire S157;
wire S158;
wire S159;
wire S160;
wire S161;
wire S162;
wire S163;
wire S164;
wire S165;
wire S166;
wire S167;
wire S168;
wire S169;
wire S170;
wire S171;
wire S172;
wire S173;
wire S174;
wire S175;
wire S176;
wire S177;
wire S178;
wire S179;
wire S180;
wire S181;
wire S182;
wire S183;
wire S184;
wire S185;
wire S186;
wire S187;
wire S188;
wire S189;
wire S190;
wire S191;
wire S192;
wire S193;
wire S194;
wire S195;
wire S196;
wire S197;
wire S198;
wire S199;
wire S200;
wire S201;
wire S202;
wire S203;
wire S204;
wire S205;
wire S206;
wire S207;
wire S208;
wire S209;
wire S210;
wire S211;
wire S212;
wire S213;
wire S214;
wire S215;
wire S216;
wire S217;
wire S218;
wire S219;
wire S220;
wire S221;
wire S222;
wire S223;
wire S224;
wire S225;
wire S226;
wire S227;
wire S228;
wire S229;
wire S230;
wire S231;
wire S232;
wire S233;
wire S234;
wire S235;
wire S236;
wire S237;
wire S238;
wire S239;
wire S240;
wire S241;
wire S242;
wire S243;
wire S244;
wire S245;
wire S246;
wire S247;
wire S248;
wire S249;
wire S250;
wire S251;
wire S252;
wire S253;
wire S254;
wire S255;
wire S256;
wire S257;
wire S258;
wire S259;
wire S260;
wire S261;
wire S262;
wire S263;
wire S264;
wire S265;
wire S266;
wire S267;
wire S268;
wire S269;
wire S270;
wire S271;
wire S272;
wire S273;
wire S274;
wire S275;
wire S276;
wire S277;
wire S278;
wire S279;
wire S280;
wire S281;
wire S282;
wire S283;
wire S284;
wire S285;
wire S286;
wire S287;
wire S288;
wire S289;
wire S290;
wire S291;
wire S292;
wire S293;
wire S294;
wire S295;
wire S296;
wire S297;
wire S298;
wire S299;
wire S300;
wire S301;
wire S302;
wire S303;
wire S304;
wire S305;
wire S306;
wire S307;
wire S308;
wire S309;
wire S310;
wire S311;
wire S312;
wire S313;
wire S314;
wire S315;
wire S316;
wire S317;
wire S318;
wire S319;
wire S320;
wire S321;
wire S322;
wire S323;
wire S324;
wire S325;
wire S326;
wire S327;
wire S328;
wire S329;
wire S330;
wire S331;
wire S332;
wire S333;
wire S334;
wire S335;
wire S336;
wire S337;
wire S338;
wire S339;
wire S340;
wire S341;
wire S342;
wire S343;
wire S344;
wire S345;
wire S346;
wire S347;
wire S348;
wire S349;
wire S350;
wire S351;
wire S352;
wire S353;
wire S354;
wire S355;
wire S356;
wire S357;
wire S358;
wire S359;
wire S360;
wire S361;
wire S362;
wire S363;
wire S364;
wire S365;
wire S366;
wire S367;
wire S368;
wire S369;
wire S370;
wire S371;
wire S372;
wire S373;
wire S374;
wire S375;
wire S376;
wire S377;
wire S378;
wire S379;
wire S380;
wire S381;
wire S382;
wire S383;
wire S384;
wire S385;
wire S386;
wire S387;
wire S388;
wire S389;
wire S390;
wire S391;
wire S392;
wire S393;
wire S394;
wire S395;
wire S396;
wire S397;
wire S398;
wire S399;
wire S400;
wire S401;
wire S402;
wire S403;
wire S404;
wire S405;
wire S406;
wire S407;
wire S408;
wire S409;
wire S410;
wire S411;
wire S412;
wire S413;
wire S414;
wire S415;
wire S416;
wire S417;
wire S418;
wire S419;
wire S420;
wire S421;
wire S422;
wire S423;
wire S424;
wire S425;
wire S426;
wire S427;
wire S428;
wire S429;
wire S430;
wire S431;
wire S432;
wire S433;
wire S434;
wire S435;
wire S436;
wire S437;
wire S438;
wire S439;
wire S440;
wire S441;
wire S442;
wire S443;
wire S444;
wire S445;
wire S446;
wire S447;
wire S448;
wire S449;
wire S450;
wire S451;
wire S452;
wire S453;
wire S454;
wire S455;
wire S456;
wire S457;
wire S458;
wire S459;
wire S460;
wire S461;
wire S462;
wire S463;
wire S464;
wire S465;
wire S466;
wire S467;
wire S468;
wire S469;
wire S470;
wire S471;
wire S472;
wire S473;
wire S474;
wire S475;
wire S476;
wire S477;
wire S478;
wire S479;
wire S480;
wire S481;
wire S482;
wire S483;
wire S484;
wire S485;
wire S486;
wire S487;
wire S488;
wire S489;
wire S490;
wire S491;
wire S492;
wire S493;
wire S494;
wire S495;
wire S496;
wire S497;
wire S498;
wire S499;
wire S500;
wire S501;
wire S502;
wire S503;
wire S504;
wire S505;
wire S506;
wire S507;
wire S508;
wire S509;
wire S510;
wire S511;
wire S512;
wire S513;
wire S514;
wire S515;
wire S516;
wire S517;
wire S518;
wire S519;
wire S520;
wire S521;
wire S522;
wire S523;
wire S524;
wire S525;
wire S526;
wire S527;
wire S528;
wire S529;
wire S530;
wire S531;
wire S532;
wire S533;
wire S534;
wire S535;
wire S536;
wire S537;
wire S538;
wire S539;
wire S540;
wire S541;
wire S542;
wire S543;
wire S544;
wire S545;
wire S546;
wire S547;
wire S548;
wire S549;
wire S550;
wire S551;
wire S552;
wire S553;
wire S554;
wire S555;
wire S556;
wire S557;
wire S558;
wire S559;
wire S560;
wire S561;
wire S562;
wire S563;
wire S564;
wire S565;
wire S566;
wire S567;
wire S568;
wire S569;
wire S570;
wire S571;
wire S572;
wire S573;
wire S574;
wire S575;
wire S576;
wire S577;
wire S578;
wire S579;
wire S580;
wire S581;
wire S582;
wire S583;
wire S584;
wire S585;
wire S586;
wire S587;
wire S588;
wire S589;
wire S590;
wire S591;
wire S592;
wire S593;
wire S594;
wire S595;
wire S596;
wire S597;
wire S598;
wire S599;
wire S600;
wire S601;
wire S602;
wire S603;
wire S604;
wire S605;
wire S606;
wire S607;
wire S608;
wire S609;
wire S610;
wire S611;
wire S612;
wire S613;
wire S614;
wire S615;
wire S616;
wire S617;
wire S618;
wire S619;
wire S620;
wire S621;
wire S622;
wire S623;
wire S624;
wire S625;
wire S626;
wire S627;
wire S628;
wire S629;
wire S630;
wire S631;
wire S632;
wire S633;
wire S634;
wire S635;
wire S636;
wire S637;
wire S638;
wire S639;
wire S640;
wire S641;
wire S642;
wire S643;
wire S644;
wire S645;
wire S646;
wire S647;
wire S648;
wire S649;
wire S650;
wire S651;
wire S652;
wire S653;
wire S654;
wire S655;
wire S656;
wire S657;
wire S658;
wire S659;
wire S660;
wire S661;
wire S662;
wire S663;
wire S664;
wire S665;
wire S666;
wire S667;
wire S668;
wire S669;
wire S670;
wire S671;
wire S672;
wire S673;
wire S674;
wire S675;
wire S676;
wire S677;
wire S678;
wire S679;
wire S680;
wire S681;
wire S682;
wire S683;
wire S684;
wire S685;
wire S686;
wire S687;
wire S688;
wire S689;
wire S690;
wire S691;
wire S692;
wire S693;
wire S694;
wire S695;
wire S696;
wire S697;
wire S698;
wire S699;
wire S700;
wire S701;
wire S702;
wire S703;
wire S704;
wire S705;
wire S706;
wire S707;
wire S708;
wire S709;
wire S710;
wire S711;
wire S712;
wire S713;
wire S714;
wire S715;
wire S716;
wire S717;
wire S718;
wire S719;
wire S720;
wire S721;
wire S722;
wire S723;
wire S724;
wire S725;
wire S726;
wire S727;
wire S728;
wire S729;
wire S730;
wire S731;
wire S732;
wire S733;
wire S734;
wire S735;
wire S736;
wire S737;
wire S738;
wire S739;
wire S740;
wire S741;
wire S742;
wire S743;
wire S744;
wire S745;
wire S746;
wire S747;
wire S748;
wire S749;
wire S750;
wire S751;
wire S752;
wire S753;
wire S754;
wire S755;
wire S756;
wire S757;
wire S758;
wire S759;
wire S760;
wire S761;
wire S762;
wire S763;
wire S764;
wire S765;
wire S766;
wire S767;
wire S768;
wire S769;
wire S770;
wire S771;
wire S772;
wire S773;
wire S774;
wire S775;
wire S776;
wire S777;
wire S778;
wire S779;
wire S780;
wire S781;
wire S782;
wire S783;
wire S784;
wire S785;
wire S786;
wire S787;
wire S788;
wire S789;
wire S790;
wire S791;
wire S792;
wire S793;
wire S794;
wire S795;
wire S796;
wire S797;
wire S798;
wire S799;
wire S800;
wire S801;
wire S802;
wire S803;
wire S804;
wire S805;
wire S806;
wire S807;
wire S808;
wire S809;
wire S810;
wire S811;
wire S812;
wire S813;
wire S814;
wire S815;
wire S816;
wire S817;
wire S818;
wire S819;
wire S820;
wire S821;
wire S822;
wire S823;
wire S824;
wire S825;
wire S826;
wire S827;
wire S828;
wire S829;
wire S830;
wire S831;
wire S832;
wire S833;
wire S834;
wire S835;
wire S836;
wire S837;
wire S838;
wire S839;
wire S840;
wire S841;
wire S842;
wire S843;
wire S844;
wire S845;
wire S846;
wire S847;
wire S848;
wire S849;
wire S850;
wire S851;
wire S852;
wire S853;
wire S854;
wire S855;
wire S856;
wire S857;
wire S858;
wire S859;
wire S860;
wire S861;
wire S862;
wire S863;
wire S864;
wire S865;
wire S866;
wire S867;
wire S868;
wire S869;
wire S870;
wire S871;
wire S872;
wire S873;
wire S874;
wire S875;
wire S876;
wire S877;
wire S878;
wire S879;
wire S880;
wire S881;
wire S882;
wire S883;
wire S884;
wire S885;
wire S886;
wire S887;
wire S888;
wire S889;
wire S890;
wire S891;
wire S892;
wire S893;
wire S894;
wire S895;
wire S896;
wire S897;
wire S898;
wire S899;
wire S900;
wire S901;
wire S902;
wire S903;
wire S904;
wire S905;
wire S906;
wire S907;
wire S908;
wire S909;
wire S910;
wire S911;
wire S912;
wire S913;
wire S914;
wire S915;
wire S916;
wire S917;
wire S918;
wire S919;
wire S920;
wire S921;
wire S922;
wire S923;
wire S924;
wire S925;
wire S926;
wire S927;
wire S928;
wire S929;
wire S930;
wire S931;
wire S932;
wire S933;
wire S934;
wire S935;
wire S936;
wire S937;
wire S938;
wire S939;
wire S940;
wire S941;
wire S942;
wire S943;
wire S944;
wire S945;
wire S946;
wire S947;
wire S948;
wire S949;
wire S950;
wire S951;
wire S952;
wire S953;
wire S954;
wire S955;
wire S956;
wire S957;
wire S958;
wire S959;
wire S960;
wire S961;
wire S962;
wire S963;
wire S964;
wire S965;
wire S966;
wire S967;
wire S968;
wire S969;
wire S970;
wire S971;
wire S972;
wire S973;
wire S974;
wire S975;
wire S976;
wire S977;
wire S978;
wire S979;
wire S980;
wire S981;
wire S982;
wire S983;
wire S984;
wire S985;
wire S986;
wire S987;
wire S988;
wire S989;
wire S990;
wire S991;
wire S992;
wire S993;
wire S994;
wire S995;
wire S996;
wire S997;
wire S998;
wire S999;
wire S1000;
wire S1001;
wire S1002;
wire S1003;
wire S1004;
wire S1005;
wire S1006;
wire S1007;
wire S1008;
wire S1009;
wire S1010;
wire S1011;
wire S1012;
wire S1013;
wire S1014;
wire S1015;
wire S1016;
wire S1017;
wire S1018;
wire S1019;
wire S1020;
wire S1021;
wire S1022;
wire S1023;
wire S1024;
wire S1025;
wire S1026;
wire S1027;
wire S1028;
wire S1029;
wire S1030;
wire S1031;
wire S1032;
wire S1033;
wire S1034;
wire S1035;
wire S1036;
wire S1037;
wire S1038;
wire S1039;
wire S1040;
wire S1041;
wire S1042;
wire S1043;
wire S1044;
wire S1045;
wire S1046;
wire S1047;
wire S1048;
wire S1049;
wire S1050;
wire S1051;
wire S1052;
wire S1053;
wire S1054;
wire S1055;
wire S1056;
wire S1057;
wire S1058;
wire S1059;
wire S1060;
wire S1061;
wire S1062;
wire S1063;
wire S1064;
wire S1065;
wire S1066;
wire S1067;
wire S1068;
wire S1069;
wire S1070;
wire S1071;
wire S1072;
wire S1073;
wire S1074;
wire S1075;
wire S1076;
wire S1077;
wire S1078;
wire S1079;
wire S1080;
wire S1081;
wire S1082;
wire S1083;
wire S1084;
wire S1085;
wire S1086;
wire S1087;
wire S1088;
wire S1089;
wire S1090;
wire S1091;
wire S1092;
wire S1093;
wire S1094;
wire S1095;
wire S1096;
wire S1097;
wire S1098;
wire S1099;
wire S1100;
wire S1101;
wire S1102;
wire S1103;
wire S1104;
wire S1105;
wire S1106;
wire S1107;
wire S1108;
wire S1109;
wire S1110;
wire S1111;
wire S1112;
wire S1113;
wire S1114;
wire S1115;
wire S1116;
wire S1117;
wire S1118;
wire S1119;
wire S1120;
wire S1121;
wire S1122;
wire S1123;
wire S1124;
wire S1125;
wire S1126;
wire S1127;
wire S1128;
wire S1129;
wire S1130;
wire S1131;
wire S1132;
wire S1133;
wire S1134;
wire S1135;
wire S1136;
wire S1137;
wire S1138;
wire S1139;
wire S1140;
wire S1141;
wire S1142;
wire S1143;
wire S1144;
wire S1145;
wire S1146;
wire S1147;
wire S1148;
wire S1149;
wire S1150;
wire S1151;
wire S1152;
wire S1153;
wire S1154;
wire S1155;
wire S1156;
wire S1157;
wire S1158;
wire S1159;
wire S1160;
wire S1161;
wire S1162;
wire S1163;
wire S1164;
wire S1165;
wire S1166;
wire S1167;
wire S1168;
wire S1169;
wire S1170;
wire S1171;
wire S1172;
wire S1173;
wire S1174;
wire S1175;
wire S1176;
wire S1177;
wire S1178;
wire S1179;
wire S1180;
wire S1181;
wire S1182;
wire S1183;
wire S1184;
wire S1185;
wire S1186;
wire S1187;
wire S1188;
wire S1189;
wire S1190;
wire S1191;
wire S1192;
wire S1193;
wire S1194;
wire S1195;
wire S1196;
wire S1197;
wire S1198;
wire S1199;
wire S1200;
wire S1201;
wire S1202;
wire S1203;
wire S1204;
wire S1205;
wire S1206;
wire S1207;
wire S1208;
wire S1209;
wire S1210;
wire S1211;
wire S1212;
wire S1213;
wire S1214;
wire S1215;
wire S1216;
wire S1217;
wire S1218;
wire S1219;
wire S1220;
wire S1221;
wire S1222;
wire S1223;
wire S1224;
wire S1225;
wire S1226;
wire S1227;
wire S1228;
wire S1229;
wire S1230;
wire S1231;
wire S1232;
wire S1233;
wire S1234;
wire S1235;
wire S1236;
wire S1237;
wire S1238;
wire S1239;
wire S1240;
wire S1241;
wire S1242;
wire S1243;
wire S1244;
wire S1245;
wire S1246;
wire S1247;
wire S1248;
wire S1249;
wire S1250;
wire S1251;
wire S1252;
wire S1253;
wire S1254;
wire S1255;
wire S1256;
wire S1257;
wire S1258;
wire S1259;
wire S1260;
wire S1261;
wire S1262;
wire S1263;
wire S1264;
wire S1265;
wire S1266;
wire S1267;
wire S1268;
wire S1269;
wire S1270;
wire S1271;
wire S1272;
wire S1273;
wire S1274;
wire S1275;
wire S1276;
wire S1277;
wire S1278;
wire S1279;
wire S1280;
wire S1281;
wire S1282;
wire S1283;
wire S1284;
wire S1285;
wire S1286;
wire S1287;
wire S1288;
wire S1289;
wire S1290;
wire S1291;
wire S1292;
wire S1293;
wire S1294;
wire S1295;
wire S1296;
wire S1297;
wire S1298;
wire S1299;
wire S1300;
wire S1301;
wire S1302;
wire S1303;
wire S1304;
wire S1305;
wire S1306;
wire S1307;
wire S1308;
wire S1309;
wire S1310;
wire S1311;
wire S1312;
wire S1313;
wire S1314;
wire S1315;
wire S1316;
wire S1317;
wire S1318;
wire S1319;
wire S1320;
wire S1321;
wire S1322;
wire S1323;
wire S1324;
wire S1325;
wire S1326;
wire S1327;
wire S1328;
wire S1329;
wire S1330;
wire S1331;
wire S1332;
wire S1333;
wire S1334;
wire S1335;
wire S1336;
wire S1337;
wire S1338;
wire S1339;
wire S1340;
wire S1341;
wire S1342;
wire S1343;
wire S1344;
wire S1345;
wire S1346;
wire S1347;
wire S1348;
wire S1349;
wire S1350;
wire S1351;
wire S1352;
wire S1353;
wire S1354;
wire S1355;
wire S1356;
wire S1357;
wire S1358;
wire S1359;
wire S1360;
wire S1361;
wire S1362;
wire S1363;
wire S1364;
wire S1365;
wire S1366;
wire S1367;
wire S1368;
wire S1369;
wire S1370;
wire S1371;
wire S1372;
wire S1373;
wire S1374;
wire S1375;
wire S1376;
wire S1377;
wire S1378;
wire S1379;
wire S1380;
wire S1381;
wire S1382;
wire S1383;
wire S1384;
wire S1385;
wire S1386;
wire S1387;
wire S1388;
wire S1389;
wire S1390;
wire S1391;
wire S1392;
wire S1393;
wire S1394;
wire S1395;
wire S1396;
wire S1397;
wire S1398;
wire S1399;
wire S1400;
wire S1401;
wire S1402;
wire S1403;
wire S1404;
wire S1405;
wire S1406;
wire S1407;
wire S1408;
wire S1409;
wire S1410;
wire S1411;
wire S1412;
wire S1413;
wire S1414;
wire S1415;
wire S1416;
wire S1417;
wire S1418;
wire S1419;
wire S1420;
wire S1421;
wire S1422;
wire S1423;
wire S1424;
wire S1425;
wire S1426;
wire S1427;
wire S1428;
wire S1429;
wire S1430;
wire S1431;
wire S1432;
wire S1433;
wire S1434;
wire S1435;
wire S1436;
wire S1437;
wire S1438;
wire S1439;
wire S1440;
wire S1441;
wire S1442;
wire S1443;
wire S1444;
wire S1445;
wire S1446;
wire S1447;
wire S1448;
wire S1449;
wire S1450;
wire S1451;
wire S1452;
wire S1453;
wire S1454;
wire S1455;
wire S1456;
wire S1457;
wire S1458;
wire S1459;
wire S1460;
wire S1461;
wire S1462;
wire S1463;
wire S1464;
wire S1465;
wire S1466;
wire S1467;
wire S1468;
wire S1469;
wire S1470;
wire S1471;
wire S1472;
wire S1473;
wire S1474;
wire S1475;
wire S1476;
wire S1477;
wire S1478;
wire S1479;
wire S1480;
wire S1481;
wire S1482;
wire S1483;
wire S1484;
wire S1485;
wire S1486;
wire S1487;
wire S1488;
wire S1489;
wire S1490;
wire S1491;
wire S1492;
wire S1493;
wire S1494;
wire S1495;
wire S1496;
wire S1497;
wire S1498;
wire S1499;
wire S1500;
wire S1501;
wire S1502;
wire S1503;
wire S1504;
wire S1505;
wire S1506;
wire S1507;
wire S1508;
wire S1509;
wire S1510;
wire S1511;
wire S1512;
wire S1513;
wire S1514;
wire S1515;
wire S1516;
wire S1517;
wire S1518;
wire S1519;
wire S1520;
wire S1521;
wire S1522;
wire S1523;
wire S1524;
wire S1525;
wire S1526;
wire S1527;
wire S1528;
wire S1529;
wire S1530;
wire S1531;
wire S1532;
wire S1533;
wire S1534;
wire S1535;
wire S1536;
wire S1537;
wire S1538;
wire S1539;
wire S1540;
wire S1541;
wire S1542;
wire S1543;
wire S1544;
wire S1545;
wire S1546;
wire S1547;
wire S1548;
wire S1549;
wire S1550;
wire S1551;
wire S1552;
wire S1553;
wire S1554;
wire S1555;
wire S1556;
wire S1557;
wire S1558;
wire S1559;
wire S1560;
wire S1561;
wire S1562;
wire S1563;
wire S1564;
wire S1565;
wire S1566;
wire S1567;
wire S1568;
wire S1569;
wire S1570;
wire S1571;
wire S1572;
wire S1573;
wire S1574;
wire S1575;
wire S1576;
wire S1577;
wire S1578;
wire S1579;
wire S1580;
wire S1581;
wire S1582;
wire S1583;
wire S1584;
wire S1585;
wire S1586;
wire S1587;
wire S1588;
wire S1589;
wire S1590;
wire S1591;
wire S1592;
wire S1593;
wire S1594;
wire S1595;
wire S1596;
wire S1597;
wire S1598;
wire S1599;
wire S1600;
wire S1601;
wire S1602;
wire S1603;
wire S1604;
wire S1605;
wire S1606;
wire S1607;
wire S1608;
wire S1609;
wire S1610;
wire S1611;
wire S1612;
wire S1613;
wire S1614;
wire S1615;
wire S1616;
wire S1617;
wire S1618;
wire S1619;
wire S1620;
wire S1621;
wire S1622;
wire S1623;
wire S1624;
wire S1625;
wire S1626;
wire S1627;
wire S1628;
wire S1629;
wire S1630;
wire S1631;
wire S1632;
wire S1633;
wire S1634;
wire S1635;
wire S1636;
wire S1637;
wire S1638;
wire S1639;
wire S1640;
wire S1641;
wire S1642;
wire S1643;
wire S1644;
wire S1645;
wire S1646;
wire S1647;
wire S1648;
wire S1649;
wire S1650;
wire S1651;
wire S1652;
wire S1653;
wire S1654;
wire S1655;
wire S1656;
wire S1657;
wire S1658;
wire S1659;
wire S1660;
wire S1661;
wire S1662;
wire S1663;
wire S1664;
wire S1665;
wire S1666;
wire S1667;
wire S1668;
wire S1669;
wire S1670;
wire S1671;
wire S1672;
wire S1673;
wire S1674;
wire S1675;
wire S1676;
wire S1677;
wire S1678;
wire S1679;
wire S1680;
wire S1681;
wire S1682;
wire S1683;
wire S1684;
wire S1685;
wire S1686;
wire S1687;
wire S1688;
wire S1689;
wire S1690;
wire S1691;
wire S1692;
wire S1693;
wire S1694;
wire S1695;
wire S1696;
wire S1697;
wire S1698;
wire S1699;
wire S1700;
wire S1701;
wire S1702;
wire S1703;
wire S1704;
wire S1705;
wire S1706;
wire S1707;
wire S1708;
wire S1709;
wire S1710;
wire S1711;
wire S1712;
wire S1713;
wire S1714;
wire S1715;
wire S1716;
wire S1717;
wire S1718;
wire S1719;
wire S1720;
wire S1721;
wire S1722;
wire S1723;
wire S1724;
wire S1725;
wire S1726;
wire S1727;
wire S1728;
wire S1729;
wire S1730;
wire S1731;
wire S1732;
wire S1733;
wire S1734;
wire S1735;
wire S1736;
wire S1737;
wire S1738;
wire S1739;
wire S1740;
wire S1741;
wire S1742;
wire S1743;
wire S1744;
wire S1745;
wire S1746;
wire S1747;
wire S1748;
wire S1749;
wire S1750;
wire S1751;
wire S1752;
wire S1753;
wire S1754;
wire S1755;
wire S1756;
wire S1757;
wire S1758;
wire S1759;
wire S1760;
wire S1761;
wire S1762;
wire S1763;
wire S1764;
wire S1765;
wire S1766;
wire S1767;
wire S1768;
wire S1769;
wire S1770;
wire S1771;
wire S1772;
wire S1773;
wire S1774;
wire S1775;
wire S1776;
wire S1777;
wire S1778;
wire S1779;
wire S1780;
wire S1781;
wire S1782;
wire S1783;
wire S1784;
wire S1785;
wire S1786;
wire S1787;
wire S1788;
wire S1789;
wire S1790;
wire S1791;
wire S1792;
wire S1793;
wire S1794;
wire S1795;
wire S1796;
wire S1797;
wire S1798;
wire S1799;
wire S1800;
wire S1801;
wire S1802;
wire S1803;
wire S1804;
wire S1805;
wire S1806;
wire S1807;
wire S1808;
wire S1809;
wire S1810;
wire S1811;
wire S1812;
wire S1813;
wire S1814;
wire S1815;
wire S1816;
wire S1817;
wire S1818;
wire S1819;
wire S1820;
wire S1821;
wire S1822;
wire S1823;
wire S1824;
wire S1825;
wire S1826;
wire S1827;
wire S1828;
wire S1829;
wire S1830;
wire S1831;
wire S1832;
wire S1833;
wire S1834;
wire S1835;
wire S1836;
wire S1837;
wire S1838;
wire S1839;
wire S1840;
wire S1841;
wire S1842;
wire S1843;
wire S1844;
wire S1845;
wire S1846;
wire S1847;
wire S1848;
wire S1849;
wire S1850;
wire S1851;
wire S1852;
wire S1853;
wire S1854;
wire S1855;
wire S1856;
wire S1857;
wire S1858;
wire S1859;
wire S1860;
wire S1861;
wire S1862;
wire S1863;
wire S1864;
wire S1865;
wire S1866;
wire S1867;
wire S1868;
wire S1869;
wire S1870;
wire S1871;
wire S1872;
wire S1873;
wire S1874;
wire S1875;
wire S1876;
wire S1877;
wire S1878;
wire S1879;
wire S1880;
wire S1881;
wire S1882;
wire S1883;
wire S1884;
wire S1885;
wire S1886;
wire S1887;
wire S1888;
wire S1889;
wire S1890;
wire S1891;
wire S1892;
wire S1893;
wire S1894;
wire S1895;
wire S1896;
wire S1897;
wire S1898;
wire S1899;
wire S1900;
wire S1901;
wire S1902;
wire S1903;
wire S1904;
wire S1905;
wire S1906;
wire S1907;
wire S1908;
wire S1909;
wire S1910;
wire S1911;
wire S1912;
wire S1913;
wire S1914;
wire S1915;
wire S1916;
wire S1917;
wire S1918;
wire S1919;
wire S1920;
wire S1921;
wire S1922;
wire S1923;
wire S1924;
wire S1925;
wire S1926;
wire S1927;
wire S1928;
wire S1929;
wire S1930;
wire S1931;
wire S1932;
wire S1933;
wire S1934;
wire S1935;
wire S1936;
wire S1937;
wire S1938;
wire S1939;
wire S1940;
wire S1941;
wire S1942;
wire S1943;
wire S1944;
wire S1945;
wire S1946;
wire S1947;
wire S1948;
wire S1949;
wire S1950;
wire S1951;
wire S1952;
wire S1953;
wire S1954;
wire S1955;
wire S1956;
wire S1957;
wire S1958;
wire S1959;
wire S1960;
wire S1961;
wire S1962;
wire S1963;
wire S1964;
wire S1965;
wire S1966;
wire S1967;
wire S1968;
wire S1969;
wire S1970;
wire S1971;
wire S1972;
wire S1973;
wire S1974;
wire S1975;
wire S1976;
wire S1977;
wire S1978;
wire S1979;
wire S1980;
wire S1981;
wire S1982;
wire S1983;
wire S1984;
wire S1985;
wire S1986;
wire S1987;
wire S1988;
wire S1989;
wire S1990;
wire S1991;
wire S1992;
wire S1993;
wire S1994;
wire S1995;
wire S1996;
wire S1997;
wire S1998;
wire S1999;
wire S2000;
wire S2001;
wire S2002;
wire S2003;
wire S2004;
wire S2005;
wire S2006;
wire S2007;
wire S2008;
wire S2009;
wire S2010;
wire S2011;
wire S2012;
wire S2013;
wire S2014;
wire S2015;
wire S2016;
wire S2017;
wire S2018;
wire S2019;
wire S2020;
wire S2021;
wire S2022;
wire S2023;
wire S2024;
wire S2025;
wire S2026;
wire S2027;
wire S2028;
wire S2029;
wire S2030;
wire S2031;
wire S2032;
wire S2033;
wire S2034;
wire S2035;
wire S2036;
wire S2037;
wire S2038;
wire S2039;
wire S2040;
wire S2041;
wire S2042;
wire S2043;
wire S2044;
wire S2045;
wire S2046;
wire S2047;
wire S2048;
wire S2049;
wire S2050;
wire S2051;
wire S2052;
wire S2053;
wire S2054;
wire S2055;
wire S2056;
wire S2057;
wire S2058;
wire S2059;
wire S2060;
wire S2061;
wire S2062;
wire S2063;
wire S2064;
wire S2065;
wire S2066;
wire S2067;
wire S2068;
wire S2069;
wire S2070;
wire S2071;
wire S2072;
wire S2073;
wire S2074;
wire S2075;
wire S2076;
wire S2077;
wire S2078;
wire S2079;
wire S2080;
wire S2081;
wire S2082;
wire S2083;
wire S2084;
wire S2085;
wire S2086;
wire S2087;
wire S2088;
wire S2089;
wire S2090;
wire S2091;
wire S2092;
wire S2093;
wire S2094;
wire S2095;
wire S2096;
wire S2097;
wire S2098;
wire S2099;
wire S2100;
wire S2101;
wire S2102;
wire S2103;
wire S2104;
wire S2105;
wire S2106;
wire S2107;
wire S2108;
wire S2109;
wire S2110;
wire S2111;
wire S2112;
wire S2113;
wire S2114;
wire S2115;
wire S2116;
wire S2117;
wire S2118;
wire S2119;
wire S2120;
wire S2121;
wire S2122;
wire S2123;
wire S2124;
wire S2125;
wire S2126;
wire S2127;
wire S2128;
wire S2129;
wire S2130;
wire S2131;
wire S2132;
wire S2133;
wire S2134;
wire S2135;
wire S2136;
wire S2137;
wire S2138;
wire S2139;
wire S2140;
wire S2141;
wire S2142;
wire S2143;
wire S2144;
wire S2145;
wire S2146;
wire S2147;
wire S2148;
wire S2149;
wire S2150;
wire S2151;
wire S2152;
wire S2153;
wire S2154;
wire S2155;
wire S2156;
wire S2157;
wire S2158;
wire S2159;
wire S2160;
wire S2161;
wire S2162;
wire S2163;
wire S2164;
wire S2165;
wire S2166;
wire S2167;
wire S2168;
wire S2169;
wire S2170;
wire S2171;
wire S2172;
wire S2173;
wire S2174;
wire S2175;
wire S2176;
wire S2177;
wire S2178;
wire S2179;
wire S2180;
wire S2181;
wire S2182;
wire S2183;
wire S2184;
wire S2185;
wire S2186;
wire S2187;
wire S2188;
wire S2189;
wire S2190;
wire S2191;
wire S2192;
wire S2193;
wire S2194;
wire S2195;
wire S2196;
wire S2197;
wire S2198;
wire S2199;
wire S2200;
wire S2201;
wire S2202;
wire S2203;
wire S2204;
wire S2205;
wire S2206;
wire S2207;
wire S2208;
wire S2209;
wire S2210;
wire S2211;
wire S2212;
wire S2213;
wire S2214;
wire S2215;
wire S2216;
wire S2217;
wire S2218;
wire S2219;
wire S2220;
wire S2221;
wire S2222;
wire S2223;
wire S2224;
wire S2225;
wire S2226;
wire S2227;
wire S2228;
wire S2229;
wire S2230;
wire S2231;
wire S2232;
wire S2233;
wire S2234;
wire S2235;
wire S2236;
wire S2237;
wire S2238;
wire S2239;
wire S2240;
wire S2241;
wire S2242;
wire S2243;
wire S2244;
wire S2245;
wire S2246;
wire S2247;
wire S2248;
wire S2249;
wire S2250;
wire S2251;
wire S2252;
wire S2253;
wire S2254;
wire S2255;
wire S2256;
wire S2257;
wire S2258;
wire S2259;
wire S2260;
wire S2261;
wire S2262;
wire S2263;
wire S2264;
wire S2265;
wire S2266;
wire S2267;
wire S2268;
wire S2269;
wire S2270;
wire S2271;
wire S2272;
wire S2273;
wire S2274;
wire S2275;
wire S2276;
wire S2277;
wire S2278;
wire S2279;
wire S2280;
wire S2281;
wire S2282;
wire S2283;
wire S2284;
wire S2285;
wire S2286;
wire S2287;
wire S2288;
wire S2289;
wire S2290;
wire S2291;
wire S2292;
wire S2293;
wire S2294;
wire S2295;
wire S2296;
wire S2297;
wire S2298;
wire S2299;
wire S2300;
wire S2301;
wire S2302;
wire S2303;
wire S2304;
wire S2305;
wire S2306;
wire S2307;
wire S2308;
wire S2309;
wire S2310;
wire S2311;
wire S2312;
wire S2313;
wire S2314;
wire S2315;
wire S2316;
wire S2317;
wire S2318;
wire S2319;
wire S2320;
wire S2321;
wire S2322;
wire S2323;
wire S2324;
wire S2325;
wire S2326;
wire S2327;
wire S2328;
wire S2329;
wire S2330;
wire S2331;
wire S2332;
wire S2333;
wire S2334;
wire S2335;
wire S2336;
wire S2337;
wire S2338;
wire S2339;
wire S2340;
wire S2341;
wire S2342;
wire S2343;
wire S2344;
wire S2345;
wire S2346;
wire S2347;
wire S2348;
wire S2349;
wire S2350;
wire S2351;
wire S2352;
wire S2353;
wire S2354;
wire S2355;
wire S2356;
wire S2357;
wire S2358;
wire S2359;
wire S2360;
wire S2361;
wire S2362;
wire S2363;
wire S2364;
wire S2365;
wire S2366;
wire S2367;
wire S2368;
wire S2369;
wire S2370;
wire S2371;
wire S2372;
wire S2373;
wire S2374;
wire S2375;
wire S2376;
wire S2377;
wire S2378;
wire S2379;
wire S2380;
wire S2381;
wire S2382;
wire S2383;
wire S2384;
wire S2385;
wire S2386;
wire S2387;
wire S2388;
wire S2389;
wire S2390;
wire S2391;
wire S2392;
wire S2393;
wire S2394;
wire S2395;
wire S2396;
wire S2397;
wire S2398;
wire S2399;
wire S2400;
wire S2401;
wire S2402;
wire S2403;
wire S2404;
wire S2405;
wire S2406;
wire S2407;
wire S2408;
wire S2409;
wire S2410;
wire S2411;
wire S2412;
wire S2413;
wire S2414;
wire S2415;
wire S2416;
wire S2417;
wire S2418;
wire S2419;
wire S2420;
wire S2421;
wire S2422;
wire S2423;
wire S2424;
wire S2425;
wire S2426;
wire S2427;
wire S2428;
wire S2429;
wire S2430;
wire S2431;
wire S2432;
wire S2433;
wire S2434;
wire S2435;
wire S2436;
wire S2437;
wire S2438;
wire S2439;
wire S2440;
wire S2441;
wire S2442;
wire S2443;
wire S2444;
wire S2445;
wire S2446;
wire S2447;
wire S2448;
wire S2449;
wire S2450;
wire S2451;
wire S2452;
wire S2453;
wire S2454;
wire S2455;
wire S2456;
wire S2457;
wire S2458;
wire S2459;
wire S2460;
wire S2461;
wire S2462;
wire S2463;
wire S2464;
wire S2465;
wire S2466;
wire S2467;
wire S2468;
wire S2469;
wire S2470;
wire S2471;
wire S2472;
wire S2473;
wire S2474;
wire S2475;
wire S2476;
wire S2477;
wire S2478;
wire S2479;
wire S2480;
wire S2481;
wire S2482;
wire S2483;
wire S2484;
wire S2485;
wire S2486;
wire S2487;
wire S2488;
wire S2489;
wire S2490;
wire S2491;
wire S2492;
wire S2493;
wire S2494;
wire S2495;
wire S2496;
wire S2497;
wire S2498;
wire S2499;
wire S2500;
wire S2501;
wire S2502;
wire S2503;
wire S2504;
wire S2505;
wire S2506;
wire S2507;
wire S2508;
wire S2509;
wire S2510;
wire S2511;
wire S2512;
wire S2513;
wire S2514;
wire S2515;
wire S2516;
wire S2517;
wire S2518;
wire S2519;
wire S2520;
wire S2521;
wire S2522;
wire S2523;
wire S2524;
wire S2525;
wire S2526;
wire S2527;
wire S2528;
wire S2529;
wire S2530;
wire S2531;
wire S2532;
wire S2533;
wire S2534;
wire S2535;
wire S2536;
wire S2537;
wire S2538;
wire S2539;
wire S2540;
wire S2541;
wire S2542;
wire S2543;
wire S2544;
wire S2545;
wire S2546;
wire S2547;
wire S2548;
wire S2549;
wire S2550;
wire S2551;
wire S2552;
wire S2553;
wire S2554;
wire S2555;
wire S2556;
wire S2557;
wire S2558;
wire S2559;
wire S2560;
wire S2561;
wire S2562;
wire S2563;
wire S2564;
wire S2565;
wire S2566;
wire S2567;
wire S2568;
wire S2569;
wire S2570;
wire S2571;
wire S2572;
wire S2573;
wire S2574;
wire S2575;
wire S2576;
wire S2577;
wire S2578;
wire S2579;
wire S2580;
wire S2581;
wire S2582;
wire S2583;
wire S2584;
wire S2585;
wire S2586;
wire S2587;
wire S2588;
wire S2589;
wire S2590;
wire S2591;
wire S2592;
wire S2593;
wire S2594;
wire S2595;
wire S2596;
wire S2597;
wire S2598;
wire S2599;
wire S2600;
wire S2601;
wire S2602;
wire S2603;
wire S2604;
wire S2605;
wire S2606;
wire S2607;
wire S2608;
wire S2609;
wire S2610;
wire S2611;
wire S2612;
wire S2613;
wire S2614;
wire S2615;
wire S2616;
wire S2617;
wire S2618;
wire S2619;
wire S2620;
wire S2621;
wire S2622;
wire S2623;
wire S2624;
wire S2625;
wire S2626;
wire S2627;
wire S2628;
wire S2629;
wire S2630;
wire S2631;
wire S2632;
wire S2633;
wire S2634;
wire S2635;
wire S2636;
wire S2637;
wire S2638;
wire S2639;
wire S2640;
wire S2641;
wire S2642;
wire S2643;
wire S2644;
wire S2645;
wire S2646;
wire S2647;
wire S2648;
wire S2649;
wire S2650;
wire S2651;
wire S2652;
wire S2653;
wire S2654;
wire S2655;
wire S2656;
wire S2657;
wire S2658;
wire S2659;
wire S2660;
wire S2661;
wire S2662;
wire S2663;
wire S2664;
wire S2665;
wire S2666;
wire S2667;
wire S2668;
wire S2669;
wire S2670;
wire S2671;
wire S2672;
wire S2673;
wire S2674;
wire S2675;
wire S2676;
wire S2677;
wire S2678;
wire S2679;
wire S2680;
wire S2681;
wire S2682;
wire S2683;
wire S2684;
wire S2685;
wire S2686;
wire S2687;
wire S2688;
wire S2689;
wire S2690;
wire S2691;
wire S2692;
wire S2693;
wire S2694;
wire S2695;
wire S2696;
wire S2697;
wire S2698;
wire S2699;
wire S2700;
wire S2701;
wire S2702;
wire S2703;
wire S2704;
wire S2705;
wire S2706;
wire S2707;
wire S2708;
wire S2709;
wire S2710;
wire S2711;
wire S2712;
wire S2713;
wire S2714;
wire S2715;
wire S2716;
wire S2717;
wire S2718;
wire S2719;
wire S2720;
wire S2721;
wire S2722;
wire S2723;
wire S2724;
wire S2725;
wire S2726;
wire S2727;
wire S2728;
wire S2729;
wire S2730;
wire S2731;
wire S2732;
wire S2733;
wire S2734;
wire S2735;
wire S2736;
wire S2737;
wire S2738;
wire S2739;
wire S2740;
wire S2741;
wire S2742;
wire S2743;
wire S2744;
wire S2745;
wire S2746;
wire S2747;
wire S2748;
wire S2749;
wire S2750;
wire S2751;
wire S2752;
wire S2753;
wire S2754;
wire S2755;
wire S2756;
wire S2757;
wire S2758;
wire S2759;
wire S2760;
wire S2761;
wire S2762;
wire S2763;
wire S2764;
wire S2765;
wire S2766;
wire S2767;
wire S2768;
wire S2769;
wire S2770;
wire S2771;
wire S2772;
wire S2773;
wire S2774;
wire S2775;
wire S2776;
wire S2777;
wire S2778;
wire S2779;
wire S2780;
wire S2781;
wire S2782;
wire S2783;
wire S2784;
wire S2785;
wire S2786;
wire S2787;
wire S2788;
wire S2789;
wire S2790;
wire S2791;
wire S2792;
wire S2793;
wire S2794;
wire S2795;
wire S2796;
wire S2797;
wire S2798;
wire S2799;
wire S2800;
wire S2801;
wire S2802;
wire S2803;
wire S2804;
wire S2805;
wire S2806;
wire S2807;
wire S2808;
wire S2809;
wire S2810;
wire S2811;
wire S2812;
wire S2813;
wire S2814;
wire S2815;
wire S2816;
wire S2817;
wire S2818;
wire S2819;
wire S2820;
wire S2821;
wire S2822;
wire S2823;
wire S2824;
wire S2825;
wire S2826;
wire S2827;
wire S2828;
wire S2829;
wire S2830;
wire S2831;
wire S2832;
wire S2833;
wire S2834;
wire S2835;
wire S2836;
wire S2837;
wire S2838;
wire S2839;
wire S2840;
wire S2841;
wire S2842;
wire S2843;
wire S2844;
wire S2845;
wire S2846;
wire S2847;
wire S2848;
wire S2849;
wire S2850;
wire S2851;
wire S2852;
wire S2853;
wire S2854;
wire S2855;
wire S2856;
wire S2857;
wire S2858;
wire S2859;
wire S2860;
wire S2861;
wire S2862;
wire S2863;
wire S2864;
wire S2865;
wire S2866;
wire S2867;
wire S2868;
wire S2869;
wire S2870;
wire S2871;
wire S2872;
wire S2873;
wire S2874;
wire S2875;
wire S2876;
wire S2877;
wire S2878;
wire S2879;
wire S2880;
wire S2881;
wire S2882;
wire S2883;
wire S2884;
wire S2885;
wire S2886;
wire S2887;
wire S2888;
wire S2889;
wire S2890;
wire S2891;
wire S2892;
wire S2893;
wire S2894;
wire S2895;
wire S2896;
wire S2897;
wire S2898;
wire S2899;
wire S2900;
wire S2901;
wire S2902;
wire S2903;
wire S2904;
wire S2905;
wire S2906;
wire S2907;
wire S2908;
wire S2909;
wire S2910;
wire S2911;
wire S2912;
wire S2913;
wire S2914;
wire S2915;
wire S2916;
wire S2917;
wire S2918;
wire S2919;
wire S2920;
wire S2921;
wire S2922;
wire S2923;
wire S2924;
wire S2925;
wire S2926;
wire S2927;
wire S2928;
wire S2929;
wire S2930;
wire S2931;
wire S2932;
wire S2933;
wire S2934;
wire S2935;
wire S2936;
wire S2937;
wire S2938;
wire S2939;
wire S2940;
wire S2941;
wire S2942;
wire S2943;
wire S2944;
wire S2945;
wire S2946;
wire S2947;
wire S2948;
wire S2949;
wire S2950;
wire S2951;
wire S2952;
wire S2953;
wire S2954;
wire S2955;
wire S2956;
wire S2957;
wire S2958;
wire S2959;
wire S2960;
wire S2961;
wire S2962;
wire S2963;
wire S2964;
wire S2965;
wire S2966;
wire S2967;
wire S2968;
wire S2969;
wire S2970;
wire S2971;
wire S2972;
wire S2973;
wire S2974;
wire S2975;
wire S2976;
wire S2977;
wire S2978;
wire S2979;
wire S2980;
wire S2981;
wire S2982;
wire S2983;
wire S2984;
wire S2985;
wire S2986;
wire S2987;
wire S2988;
wire S2989;
wire S2990;
wire S2991;
wire S2992;
wire S2993;
wire S2994;
wire S2995;
wire S2996;
wire S2997;
wire S2998;
wire S2999;
wire S3000;
wire S3001;
wire S3002;
wire S3003;
wire S3004;
wire S3005;
wire S3006;
wire S3007;
wire S3008;
wire S3009;
wire S3010;
wire S3011;
wire S3012;
wire S3013;
wire S3014;
wire S3015;
wire S3016;
wire S3017;
wire S3018;
wire S3019;
wire S3020;
wire S3021;
wire S3022;
wire S3023;
wire S3024;
wire S3025;
wire S3026;
wire S3027;
wire S3028;
wire S3029;
wire S3030;
wire S3031;
wire S3032;
wire S3033;
wire S3034;
wire S3035;
wire S3036;
wire S3037;
wire S3038;
wire S3039;
wire S3040;
wire S3041;
wire S3042;
wire S3043;
wire S3044;
wire S3045;
wire S3046;
wire S3047;
wire S3048;
wire S3049;
wire S3050;
wire S3051;
wire S3052;
wire S3053;
wire S3054;
wire S3055;
wire S3056;
wire S3057;
wire S3058;
wire S3059;
wire S3060;
wire S3061;
wire S3062;
wire S3063;
wire S3064;
wire S3065;
wire S3066;
wire S3067;
wire S3068;
wire S3069;
wire S3070;
wire S3071;
wire S3072;
wire S3073;
wire S3074;
wire S3075;
wire S3076;
wire S3077;
wire S3078;
wire S3079;
wire S3080;
wire S3081;
wire S3082;
wire S3083;
wire S3084;
wire S3085;
wire S3086;
wire S3087;
wire S3088;
wire S3089;
wire S3090;
wire S3091;
wire S3092;
wire S3093;
wire S3094;
wire S3095;
wire S3096;
wire S3097;
wire S3098;
wire S3099;
wire S3100;
wire S3101;
wire S3102;
wire S3103;
wire S3104;
wire S3105;
wire S3106;
wire S3107;
wire S3108;
wire S3109;
wire S3110;
wire S3111;
wire S3112;
wire S3113;
wire S3114;
wire S3115;
wire S3116;
wire S3117;
wire S3118;
wire S3119;
wire S3120;
wire S3121;
wire S3122;
wire S3123;
wire S3124;
wire S3125;
wire S3126;
wire S3127;
wire S3128;
wire S3129;
wire S3130;
wire S3131;
wire S3132;
wire S3133;
wire S3134;
wire S3135;
wire S3136;
wire S3137;
wire S3138;
wire S3139;
wire S3140;
wire S3141;
wire S3142;
wire S3143;
wire S3144;
wire S3145;
wire S3146;
wire S3147;
wire S3148;
wire S3149;
wire S3150;
wire S3151;
wire S3152;
wire S3153;
wire S3154;
wire S3155;
wire S3156;
wire S3157;
wire S3158;
wire S3159;
wire S3160;
wire S3161;
wire S3162;
wire S3163;
wire S3164;
wire S3165;
wire S3166;
wire S3167;
wire S3168;
wire S3169;
wire S3170;
wire S3171;
wire S3172;
wire S3173;
wire S3174;
wire S3175;
wire S3176;
wire S3177;
wire S3178;
wire S3179;
wire S3180;
wire S3181;
wire S3182;
wire S3183;
wire S3184;
wire S3185;
wire S3186;
wire S3187;
wire S3188;
wire S3189;
wire S3190;
wire S3191;
wire S3192;
wire S3193;
wire S3194;
wire S3195;
wire S3196;
wire S3197;
wire S3198;
wire S3199;
wire S3200;
wire S3201;
wire S3202;
wire S3203;
wire S3204;
wire S3205;
wire S3206;
wire S3207;
wire S3208;
wire S3209;
wire S3210;
wire S3211;
wire S3212;
wire S3213;
wire S3214;
wire S3215;
wire S3216;
wire S3217;
wire S3218;
wire S3219;
wire S3220;
wire S3221;
wire S3222;
wire S3223;
wire S3224;
wire S3225;
wire S3226;
wire S3227;
wire S3228;
wire S3229;
wire S3230;
wire S3231;
wire S3232;
wire S3233;
wire S3234;
wire S3235;
wire S3236;
wire S3237;
wire S3238;
wire S3239;
wire S3240;
wire S3241;
wire S3242;
wire S3243;
wire S3244;
wire S3245;
wire S3246;
wire S3247;
wire S3248;
wire S3249;
wire S3250;
wire S3251;
wire S3252;
wire S3253;
wire S3254;
wire S3255;
wire S3256;
wire S3257;
wire S3258;
wire S3259;
wire S3260;
wire S3261;
wire S3262;
wire S3263;
wire S3264;
wire S3265;
wire S3266;
wire S3267;
wire S3268;
wire S3269;
wire S3270;
wire S3271;
wire S3272;
wire S3273;
wire S3274;
wire S3275;
wire S3276;
wire S3277;
wire S3278;
wire S3279;
wire S3280;
wire S3281;
wire S3282;
wire S3283;
wire S3284;
wire S3285;
wire S3286;
wire S3287;
wire S3288;
wire S3289;
wire S3290;
wire S3291;
wire S3292;
wire S3293;
wire S3294;
wire S3295;
wire S3296;
wire S3297;
wire S3298;
wire S3299;
wire S3300;
wire S3301;
wire S3302;
wire S3303;
wire S3304;
wire S3305;
wire S3306;
wire S3307;
wire S3308;
wire S3309;
wire S3310;
wire S3311;
wire S3312;
wire S3313;
wire S3314;
wire S3315;
wire S3316;
wire S3317;
wire S3318;
wire S3319;
wire S3320;
wire S3321;
wire S3322;
wire S3323;
wire S3324;
wire S3325;
wire S3326;
wire S3327;
wire S3328;
wire S3329;
wire S3330;
wire S3331;
wire S3332;
wire S3333;
wire S3334;
wire S3335;
wire S3336;
wire S3337;
wire S3338;
wire S3339;
wire S3340;
wire S3341;
wire S3342;
wire S3343;
wire S3344;
wire S3345;
wire S3346;
wire S3347;
wire S3348;
wire S3349;
wire S3350;
wire S3351;
wire S3352;
wire S3353;
wire S3354;
wire S3355;
wire S3356;
wire S3357;
wire S3358;
wire S3359;
wire S3360;
wire S3361;
wire S3362;
wire S3363;
wire S3364;
wire S3365;
wire S3366;
wire S3367;
wire S3368;
wire S3369;
wire S3370;
wire S3371;
wire S3372;
wire S3373;
wire S3374;
wire S3375;
wire S3376;
wire S3377;
wire S3378;
wire S3379;
wire S3380;
wire S3381;
wire S3382;
wire S3383;
wire S3384;
wire S3385;
wire S3386;
wire S3387;
wire S3388;
wire S3389;
wire S3390;
wire S3391;
wire S3392;
wire S3393;
wire S3394;
wire S3395;
wire S3396;
wire S3397;
wire S3398;
wire S3399;
wire S3400;
wire S3401;
wire S3402;
wire S3403;
wire S3404;
wire S3405;
wire S3406;
wire S3407;
wire S3408;
wire S3409;
wire S3410;
wire S3411;
wire S3412;
wire S3413;
wire S3414;
wire S3415;
wire S3416;
wire S3417;
wire S3418;
wire S3419;
wire S3420;
wire S3421;
wire S3422;
wire S3423;
wire S3424;
wire S3425;
wire S3426;
wire S3427;
wire S3428;
wire S3429;
wire S3430;
wire S3431;
wire S3432;
wire CU_clk;
wire CU_enSKP;
wire CU_inst_0;
wire CU_inst_10;
wire CU_inst_11;
wire CU_inst_12;
wire CU_inst_13;
wire CU_inst_14;
wire CU_inst_15;
wire CU_inst_1;
wire CU_inst_2;
wire CU_inst_3;
wire CU_inst_4;
wire CU_inst_5;
wire CU_inst_6;
wire CU_inst_7;
wire CU_inst_8;
wire CU_inst_9;
wire CU_rst;
wire DP_AC_din_0;
wire DP_AC_din_10;
wire DP_AC_din_11;
wire DP_AC_din_12;
wire DP_AC_din_13;
wire DP_AC_din_14;
wire DP_AC_din_15;
wire DP_AC_din_1;
wire DP_AC_din_2;
wire DP_AC_din_3;
wire DP_AC_din_4;
wire DP_AC_din_5;
wire DP_AC_din_6;
wire DP_AC_din_7;
wire DP_AC_din_8;
wire DP_AC_din_9;
wire DP_AC_dout_0;
wire DP_AC_dout_10;
wire DP_AC_dout_11;
wire DP_AC_dout_12;
wire DP_AC_dout_13;
wire DP_AC_dout_14;
wire DP_AC_dout_15;
wire DP_AC_dout_1;
wire DP_AC_dout_2;
wire DP_AC_dout_3;
wire DP_AC_dout_4;
wire DP_AC_dout_5;
wire DP_AC_dout_6;
wire DP_AC_dout_7;
wire DP_AC_dout_8;
wire DP_AC_dout_9;
wire DP_ARU1_C;
wire DP_ARU1_N;
wire DP_ARU1_V;
wire DP_ARU1_Z;
wire DP_ARU1_in1_0;
wire DP_ARU1_in1_10;
wire DP_ARU1_in1_11;
wire DP_ARU1_in1_12;
wire DP_ARU1_in1_13;
wire DP_ARU1_in1_14;
wire DP_ARU1_in1_15;
wire DP_ARU1_in1_1;
wire DP_ARU1_in1_2;
wire DP_ARU1_in1_3;
wire DP_ARU1_in1_4;
wire DP_ARU1_in1_5;
wire DP_ARU1_in1_6;
wire DP_ARU1_in1_7;
wire DP_ARU1_in1_8;
wire DP_ARU1_in1_9;
wire DP_ARU1_out_0;
wire DP_ARU1_out_10;
wire DP_ARU1_out_11;
wire DP_ARU1_out_12;
wire DP_ARU1_out_13;
wire DP_ARU1_out_14;
wire DP_ARU1_out_1;
wire DP_ARU1_out_2;
wire DP_ARU1_out_3;
wire DP_ARU1_out_4;
wire DP_ARU1_out_5;
wire DP_ARU1_out_6;
wire DP_ARU1_out_7;
wire DP_ARU1_out_8;
wire DP_ARU1_out_9;
wire DP_IMM1_in1_0;
wire DP_IMM1_in1_1;
wire DP_IMM1_in1_2;
wire DP_IMM1_in1_3;
wire DP_IMM1_out_0;
wire DP_IMM1_out_10;
wire DP_IMM1_out_11;
wire DP_IMM1_out_12;
wire DP_IMM1_out_13;
wire DP_IMM1_out_14;
wire DP_IMM1_out_15;
wire DP_IMM1_out_1;
wire DP_IMM1_out_2;
wire DP_IMM1_out_3;
wire DP_IMM1_out_4;
wire DP_IMM1_out_5;
wire DP_IMM1_out_6;
wire DP_IMM1_out_7;
wire DP_IMM1_out_8;
wire DP_IMM1_out_9;
wire DP_IN_din_0;
wire DP_IN_din_10;
wire DP_IN_din_11;
wire DP_IN_din_12;
wire DP_IN_din_13;
wire DP_IN_din_14;
wire DP_IN_din_15;
wire DP_IN_din_1;
wire DP_IN_din_2;
wire DP_IN_din_3;
wire DP_IN_din_4;
wire DP_IN_din_5;
wire DP_IN_din_6;
wire DP_IN_din_7;
wire DP_IN_din_8;
wire DP_IN_din_9;
wire DP_IN_dout_0;
wire DP_IN_dout_10;
wire DP_IN_dout_11;
wire DP_IN_dout_12;
wire DP_IN_dout_13;
wire DP_IN_dout_14;
wire DP_IN_dout_15;
wire DP_IN_dout_1;
wire DP_IN_dout_2;
wire DP_IN_dout_3;
wire DP_IN_dout_4;
wire DP_IN_dout_5;
wire DP_IN_dout_6;
wire DP_IN_dout_7;
wire DP_IN_dout_8;
wire DP_IN_dout_9;
wire DP_INC2_out_0;
wire DP_INC2_out_10;
wire DP_INC2_out_11;
wire DP_INC2_out_12;
wire DP_INC2_out_13;
wire DP_INC2_out_14;
wire DP_INC2_out_15;
wire DP_INC2_out_1;
wire DP_INC2_out_2;
wire DP_INC2_out_3;
wire DP_INC2_out_4;
wire DP_INC2_out_5;
wire DP_INC2_out_6;
wire DP_INC2_out_7;
wire DP_INC2_out_8;
wire DP_INC2_out_9;
wire DP_INC_1_in_0;
wire DP_INC_1_in_10;
wire DP_INC_1_in_11;
wire DP_INC_1_in_12;
wire DP_INC_1_in_13;
wire DP_INC_1_in_14;
wire DP_INC_1_in_15;
wire DP_INC_1_in_1;
wire DP_INC_1_in_2;
wire DP_INC_1_in_3;
wire DP_INC_1_in_4;
wire DP_INC_1_in_5;
wire DP_INC_1_in_6;
wire DP_INC_1_in_7;
wire DP_INC_1_in_8;
wire DP_INC_1_in_9;
wire DP_INC_1_inc_value_0;
wire DP_INC_1_inc_value_1;
wire DP_INC_1_out_0;
wire DP_INC_1_out_10;
wire DP_INC_1_out_11;
wire DP_INC_1_out_12;
wire DP_INC_1_out_13;
wire DP_INC_1_out_14;
wire DP_INC_1_out_15;
wire DP_INC_1_out_1;
wire DP_INC_1_out_2;
wire DP_INC_1_out_3;
wire DP_INC_1_out_4;
wire DP_INC_1_out_5;
wire DP_INC_1_out_6;
wire DP_INC_1_out_7;
wire DP_INC_1_out_8;
wire DP_INC_1_out_9;
wire DP_INC_2_in_0;
wire DP_INC_2_in_10;
wire DP_INC_2_in_11;
wire DP_INC_2_in_12;
wire DP_INC_2_in_13;
wire DP_INC_2_in_14;
wire DP_INC_2_in_15;
wire DP_INC_2_in_1;
wire DP_INC_2_in_2;
wire DP_INC_2_in_3;
wire DP_INC_2_in_4;
wire DP_INC_2_in_5;
wire DP_INC_2_in_6;
wire DP_INC_2_in_7;
wire DP_INC_2_in_8;
wire DP_INC_2_in_9;
wire DP_LGU1_N;
wire DP_LGU1_Z;
wire DP_LGU1_in1_0;
wire DP_LGU1_in1_10;
wire DP_LGU1_in1_11;
wire DP_LGU1_in1_12;
wire DP_LGU1_in1_13;
wire DP_LGU1_in1_14;
wire DP_LGU1_in1_15;
wire DP_LGU1_in1_1;
wire DP_LGU1_in1_2;
wire DP_LGU1_in1_3;
wire DP_LGU1_in1_4;
wire DP_LGU1_in1_5;
wire DP_LGU1_in1_6;
wire DP_LGU1_in1_7;
wire DP_LGU1_in1_8;
wire DP_LGU1_in1_9;
wire DP_LGU1_out_0;
wire DP_LGU1_out_10;
wire DP_LGU1_out_11;
wire DP_LGU1_out_12;
wire DP_LGU1_out_13;
wire DP_LGU1_out_14;
wire DP_LGU1_out_1;
wire DP_LGU1_out_2;
wire DP_LGU1_out_3;
wire DP_LGU1_out_4;
wire DP_LGU1_out_5;
wire DP_LGU1_out_6;
wire DP_LGU1_out_7;
wire DP_LGU1_out_8;
wire DP_LGU1_out_9;
wire DP_OF_din_0;
wire DP_OF_din_1;
wire DP_OF_din_2;
wire DP_OF_din_3;
wire DP_PC_din_0;
wire DP_PC_din_10;
wire DP_PC_din_11;
wire DP_PC_din_12;
wire DP_PC_din_13;
wire DP_PC_din_14;
wire DP_PC_din_15;
wire DP_PC_din_1;
wire DP_PC_din_2;
wire DP_PC_din_3;
wire DP_PC_din_4;
wire DP_PC_din_5;
wire DP_PC_din_6;
wire DP_PC_din_7;
wire DP_PC_din_8;
wire DP_PC_din_9;
wire DP_SR_C_din;
wire DP_SR_C_dout;
wire DP_SR_N_din;
wire DP_SR_N_dout;
wire DP_SR_V_din;
wire DP_SR_V_dout;
wire DP_SR_Z_din;
wire DP_SR_Z_dout;
wire DP_TriBuff_in_0;
wire DP_TriBuff_in_10;
wire DP_TriBuff_in_11;
wire DP_TriBuff_in_12;
wire DP_TriBuff_in_13;
wire DP_TriBuff_in_14;
wire DP_TriBuff_in_15;
wire DP_TriBuff_in_1;
wire DP_TriBuff_in_2;
wire DP_TriBuff_in_3;
wire DP_TriBuff_in_4;
wire DP_TriBuff_in_5;
wire DP_TriBuff_in_6;
wire DP_TriBuff_in_7;
wire DP_TriBuff_in_8;
wire DP_TriBuff_in_9;
wire DP_TriBuff_out_0;
wire DP_TriBuff_out_10;
wire DP_TriBuff_out_11;
wire DP_TriBuff_out_12;
wire DP_TriBuff_out_13;
wire DP_TriBuff_out_14;
wire DP_TriBuff_out_15;
wire DP_TriBuff_out_1;
wire DP_TriBuff_out_2;
wire DP_TriBuff_out_3;
wire DP_TriBuff_out_4;
wire DP_TriBuff_out_5;
wire DP_TriBuff_out_6;
wire DP_TriBuff_out_7;
wire DP_TriBuff_out_8;
wire DP_TriBuff_out_9;
wire DP_addrBus_0;
wire DP_addrBus_10;
wire DP_addrBus_11;
wire DP_addrBus_12;
wire DP_addrBus_13;
wire DP_addrBus_14;
wire DP_addrBus_15;
wire DP_addrBus_1;
wire DP_addrBus_2;
wire DP_addrBus_3;
wire DP_addrBus_4;
wire DP_addrBus_5;
wire DP_addrBus_6;
wire DP_addrBus_7;
wire DP_addrBus_8;
wire DP_addrBus_9;
input clk;
input rst;
output writeMEM;
output readMEM;
input [15:0] dataBus_in;output [15:0] dataBus_out;output [15:0] addrBus;
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_1_ (
  .in1({ 1'b1 }),
  .out1({ S0 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_2_ (
  .in1({ 1'b1 }),
  .out1({ S1 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_3_ (
  .in1({ 1'b1 }),
  .out1({ S2 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_4_ (
  .in1({ 1'b1 }),
  .out1({ S3 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_5_ (
  .in1({ 1'b1 }),
  .out1({ S4 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_6_ (
  .in1({ 1'b1 }),
  .out1({ S5 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_7_ (
  .in1({ 1'b1 }),
  .out1({ S6 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_8_ (
  .in1({ 1'b1 }),
  .out1({ S7 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_9_ (
  .in1({ 1'b1 }),
  .out1({ S8 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_10_ (
  .in1({ 1'b1 }),
  .out1({ S9 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_11_ (
  .in1({ 1'b1 }),
  .out1({ S10 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_12_ (
  .in1({ 1'b1 }),
  .out1({ S11 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_13_ (
  .in1({ 1'b1 }),
  .out1({ S12 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_14_ (
  .in1({ 1'b1 }),
  .out1({ S13 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_15_ (
  .in1({ 1'b1 }),
  .out1({ S14 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_16_ (
  .in1({ 1'b1 }),
  .out1({ S15 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_17_ (
  .in1({ 1'b1 }),
  .out1({ S16 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_18_ (
  .in1({ 1'b1 }),
  .out1({ S17 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_19_ (
  .in1({ 1'b1 }),
  .out1({ S18 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_20_ (
  .in1({ 1'b1 }),
  .out1({ S19 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_21_ (
  .in1({ 1'b1 }),
  .out1({ S20 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_22_ (
  .in1({ 1'b1 }),
  .out1({ S21 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_23_ (
  .in1({ 1'b1 }),
  .out1({ S22 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_24_ (
  .in1({ 1'b1 }),
  .out1({ S23 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_25_ (
  .in1({ 1'b1 }),
  .out1({ S24 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_26_ (
  .in1({ 1'b1 }),
  .out1({ S25 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_27_ (
  .in1({ 1'b1 }),
  .out1({ S26 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_28_ (
  .in1({ 1'b1 }),
  .out1({ S27 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_29_ (
  .in1({ 1'b1 }),
  .out1({ S28 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_30_ (
  .in1({ 1'b1 }),
  .out1({ S29 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_31_ (
  .in1({ 1'b1 }),
  .out1({ S30 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_32_ (
  .in1({ 1'b1 }),
  .out1({ S31 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_33_ (
  .in1({ 1'b1 }),
  .out1({ S32 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_34_ (
  .in1({ 1'b1 }),
  .out1({ S33 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_35_ (
  .in1({ 1'b1 }),
  .out1({ S34 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_36_ (
  .in1({ 1'b1 }),
  .out1({ S35 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_37_ (
  .in1({ 1'b1 }),
  .out1({ S36 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_38_ (
  .in1({ 1'b1 }),
  .out1({ S37 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_39_ (
  .in1({ 1'b1 }),
  .out1({ S38 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_40_ (
  .in1({ 1'b1 }),
  .out1({ S39 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_41_ (
  .in1({ 1'b1 }),
  .out1({ S40 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_42_ (
  .in1({ 1'b1 }),
  .out1({ S41 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_43_ (
  .in1({ 1'b0 }),
  .out1({ S42 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_44_ (
  .in1({ 1'b0 }),
  .out1({ S43 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_45_ (
  .in1({ 1'b0 }),
  .out1({ S44 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_46_ (
  .in1({ 1'b0 }),
  .out1({ S45 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_47_ (
  .in1({ 1'b0 }),
  .out1({ S46 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_48_ (
  .in1({ 1'b0 }),
  .out1({ S47 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_49_ (
  .in1({ 1'b0 }),
  .out1({ S48 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_50_ (
  .in1({ 1'b0 }),
  .out1({ S49 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_51_ (
  .in1({ 1'b0 }),
  .out1({ S50 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_52_ (
  .in1({ 1'b0 }),
  .out1({ S51 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_53_ (
  .in1({ 1'b0 }),
  .out1({ S52 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_54_ (
  .in1({ 1'b0 }),
  .out1({ S53 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_55_ (
  .in1({ 1'b0 }),
  .out1({ S54 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_56_ (
  .in1({ 1'b0 }),
  .out1({ S55 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_57_ (
  .in1({ 1'b0 }),
  .out1({ S56 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_58_ (
  .in1({ 1'b0 }),
  .out1({ S57 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_59_ (
  .in1({ 1'b0 }),
  .out1({ S58 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_60_ (
  .in1({ 1'b0 }),
  .out1({ S59 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_61_ (
  .in1({ 1'b0 }),
  .out1({ S60 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_62_ (
  .in1({ 1'b0 }),
  .out1({ S61 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_63_ (
  .in1({ 1'b0 }),
  .out1({ S62 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_64_ (
  .in1({ 1'b0 }),
  .out1({ S63 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_65_ (
  .in1({ 1'b0 }),
  .out1({ S64 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_66_ (
  .in1({ 1'b0 }),
  .out1({ S65 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_67_ (
  .in1({ 1'b0 }),
  .out1({ S66 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_68_ (
  .in1({ 1'b0 }),
  .out1({ S67 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_69_ (
  .in1({ 1'b0 }),
  .out1({ S68 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_70_ (
  .in1({ 1'b0 }),
  .out1({ S69 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_71_ (
  .in1({ 1'b0 }),
  .out1({ S70 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_72_ (
  .in1({ 1'b0 }),
  .out1({ S71 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_73_ (
  .in1({ 1'b0 }),
  .out1({ S72 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_74_ (
  .in1({ 1'b0 }),
  .out1({ S73 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_75_ (
  .in1({ 1'b0 }),
  .out1({ S74 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_76_ (
  .in1({ 1'b0 }),
  .out1({ S75 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_77_ (
  .in1({ 1'b0 }),
  .out1({ S76 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_78_ (
  .in1({ 1'b0 }),
  .out1({ S77 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_79_ (
  .in1({ 1'b0 }),
  .out1({ S78 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_80_ (
  .in1({ 1'b0 }),
  .out1({ S79 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_81_ (
  .in1({ 1'b0 }),
  .out1({ S80 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_82_ (
  .in1({ 1'b0 }),
  .out1({ S81 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_83_ (
  .in1({ 1'b0 }),
  .out1({ S82 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_84_ (
  .in1({ 1'b0 }),
  .out1({ S83 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_85_ (
  .in1({ 1'b0 }),
  .out1({ S84 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_86_ (
  .in1({ 1'b0 }),
  .out1({ S85 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_87_ (
  .in1({ 1'b0 }),
  .out1({ S86 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_88_ (
  .in1({ 1'b0 }),
  .out1({ S87 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_89_ (
  .in1({ 1'b0 }),
  .out1({ S88 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_90_ (
  .in1({ 1'b0 }),
  .out1({ S89 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_91_ (
  .in1({ 1'b0 }),
  .out1({ S90 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_92_ (
  .in1({ 1'b0 }),
  .out1({ S91 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_93_ (
  .in1({ 1'b0 }),
  .out1({ S92 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_94_ (
  .in1({ 1'b0 }),
  .out1({ S93 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_95_ (
  .in1({ 1'b0 }),
  .out1({ S94 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_96_ (
  .in1({ 1'b0 }),
  .out1({ S95 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_97_ (
  .in1({ 1'b0 }),
  .out1({ S96 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_98_ (
  .in1({ 1'b0 }),
  .out1({ S97 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_99_ (
  .in1({ 1'b0 }),
  .out1({ S98 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_100_ (
  .in1({ 1'b0 }),
  .out1({ S99 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_101_ (
  .in1({ 1'b0 }),
  .out1({ S100 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_102_ (
  .in1({ 1'b0 }),
  .out1({ S101 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_103_ (
  .in1({ 1'b0 }),
  .out1({ S102 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_104_ (
  .in1({ 1'b0 }),
  .out1({ S103 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_105_ (
  .in1({ 1'b0 }),
  .out1({ S104 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_106_ (
  .in1({ 1'b0 }),
  .out1({ S105 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_107_ (
  .in1({ 1'b0 }),
  .out1({ S106 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_108_ (
  .in1({ 1'b0 }),
  .out1({ S107 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_109_ (
  .in1({ 1'b0 }),
  .out1({ S108 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_110_ (
  .in1({ 1'b0 }),
  .out1({ S109 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_111_ (
  .in1({ 1'b0 }),
  .out1({ S110 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_112_ (
  .in1({ 1'b0 }),
  .out1({ S111 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_113_ (
  .in1({ 1'b0 }),
  .out1({ S112 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_114_ (
  .in1({ 1'b0 }),
  .out1({ S113 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_115_ (
  .in1({ 1'b0 }),
  .out1({ S114 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_116_ (
  .in1({ 1'b0 }),
  .out1({ S115 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_117_ (
  .in1({ 1'b0 }),
  .out1({ S116 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_118_ (
  .in1({ 1'b0 }),
  .out1({ S117 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_119_ (
  .in1({ 1'b0 }),
  .out1({ S118 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_120_ (
  .in1({ 1'b0 }),
  .out1({ S119 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_121_ (
  .in1({ 1'b0 }),
  .out1({ S120 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_122_ (
  .in1({ 1'b0 }),
  .out1({ S121 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_123_ (
  .in1({ 1'b0 }),
  .out1({ S122 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_124_ (
  .in1({ 1'b0 }),
  .out1({ S123 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_125_ (
  .in1({ 1'b0 }),
  .out1({ S124 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_126_ (
  .in1({ 1'b0 }),
  .out1({ S125 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_127_ (
  .in1({ 1'b0 }),
  .out1({ S126 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_128_ (
  .in1({ 1'b0 }),
  .out1({ S127 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_129_ (
  .in1({ 1'b0 }),
  .out1({ S128 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_130_ (
  .in1({ 1'b0 }),
  .out1({ S129 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_131_ (
  .in1({ 1'b0 }),
  .out1({ S130 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_132_ (
  .in1({ 1'b0 }),
  .out1({ S131 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_133_ (
  .in1({ 1'b0 }),
  .out1({ S132 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_134_ (
  .in1({ 1'b0 }),
  .out1({ S133 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_135_ (
  .in1({ 1'b0 }),
  .out1({ S134 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_136_ (
  .in1({ 1'b0 }),
  .out1({ S135 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_137_ (
  .in1({ 1'b0 }),
  .out1({ S136 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_138_ (
  .in1({ 1'b0 }),
  .out1({ S137 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_139_ (
  .in1({ 1'b0 }),
  .out1({ S138 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_140_ (
  .in1({ 1'b0 }),
  .out1({ S139 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_141_ (
  .in1({ 1'b0 }),
  .out1({ S140 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_142_ (
  .in1({ 1'b0 }),
  .out1({ S141 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_143_ (
  .in1({ 1'b0 }),
  .out1({ S142 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_144_ (
  .in1({ 1'b0 }),
  .out1({ S143 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_145_ (
  .in1({ 1'b0 }),
  .out1({ S144 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_146_ (
  .in1({ 1'b0 }),
  .out1({ S145 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_147_ (
  .in1({ 1'b0 }),
  .out1({ S146 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_148_ (
  .in1({ 1'b0 }),
  .out1({ S147 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_149_ (
  .in1({ 1'b0 }),
  .out1({ S148 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_150_ (
  .in1({ 1'b0 }),
  .out1({ S149 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_151_ (
  .in1({ 1'b0 }),
  .out1({ S150 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_152_ (
  .in1({ 1'b0 }),
  .out1({ S151 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_153_ (
  .in1({ 1'b0 }),
  .out1({ S152 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_154_ (
  .in1({ 1'b0 }),
  .out1({ S153 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_155_ (
  .in1({ 1'b0 }),
  .out1({ S154 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_156_ (
  .in1({ 1'b0 }),
  .out1({ S155 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_157_ (
  .in1({ 1'b0 }),
  .out1({ S156 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_158_ (
  .in1({ 1'b0 }),
  .out1({ S157 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_159_ (
  .in1({ 1'b0 }),
  .out1({ S158 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_160_ (
  .in1({ 1'b0 }),
  .out1({ S159 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_161_ (
  .in1({ 1'b0 }),
  .out1({ S160 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_162_ (
  .in1({ 1'b0 }),
  .out1({ S161 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_163_ (
  .in1({ 1'b0 }),
  .out1({ S162 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_164_ (
  .in1({ 1'b0 }),
  .out1({ S163 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_165_ (
  .in1({ 1'b0 }),
  .out1({ S164 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_166_ (
  .in1({ 1'b0 }),
  .out1({ S165 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_167_ (
  .in1({ 1'b0 }),
  .out1({ S166 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_168_ (
  .in1({ 1'b0 }),
  .out1({ S167 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_169_ (
  .in1({ 1'b0 }),
  .out1({ S168 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_170_ (
  .in1({ 1'b0 }),
  .out1({ S169 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_171_ (
  .in1({ 1'b0 }),
  .out1({ S170 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_172_ (
  .in1({ 1'b0 }),
  .out1({ S171 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_173_ (
  .in1({ 1'b0 }),
  .out1({ S172 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_174_ (
  .in1({ 1'b0 }),
  .out1({ S173 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_175_ (
  .in1({ 1'b0 }),
  .out1({ S174 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_176_ (
  .in1({ 1'b0 }),
  .out1({ S175 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_177_ (
  .in1({ 1'b0 }),
  .out1({ S176 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_178_ (
  .in1({ 1'b0 }),
  .out1({ S177 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_179_ (
  .in1({ 1'b0 }),
  .out1({ S178 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_180_ (
  .in1({ 1'b0 }),
  .out1({ S179 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_181_ (
  .in1({ 1'b0 }),
  .out1({ S180 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_182_ (
  .in1({ 1'b0 }),
  .out1({ S181 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_183_ (
  .in1({ 1'b0 }),
  .out1({ S182 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_184_ (
  .in1({ 1'b0 }),
  .out1({ S183 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_185_ (
  .in1({ 1'b0 }),
  .out1({ S184 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_186_ (
  .in1({ 1'b0 }),
  .out1({ S185 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_187_ (
  .in1({ 1'b0 }),
  .out1({ S186 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_188_ (
  .in1({ 1'b0 }),
  .out1({ S187 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_189_ (
  .in1({ 1'b0 }),
  .out1({ S188 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_190_ (
  .in1({ 1'b0 }),
  .out1({ S189 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_191_ (
  .in1({ 1'b0 }),
  .out1({ S190 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_192_ (
  .in1({ 1'b0 }),
  .out1({ S191 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_193_ (
  .in1({ 1'b0 }),
  .out1({ S192 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_194_ (
  .in1({ 1'b0 }),
  .out1({ S193 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_195_ (
  .in1({ 1'b0 }),
  .out1({ S194 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_196_ (
  .in1({ 1'b0 }),
  .out1({ S195 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_197_ (
  .in1({ 1'b0 }),
  .out1({ S196 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_198_ (
  .in1({ 1'b0 }),
  .out1({ S197 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_199_ (
  .in1({ 1'b0 }),
  .out1({ S198 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_200_ (
  .in1({ 1'b0 }),
  .out1({ S199 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_201_ (
  .in1({ 1'b0 }),
  .out1({ S200 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_202_ (
  .in1({ 1'b0 }),
  .out1({ S201 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_203_ (
  .in1({ 1'b0 }),
  .out1({ S202 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_204_ (
  .in1({ 1'b0 }),
  .out1({ S203 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_205_ (
  .in1({ 1'b0 }),
  .out1({ S204 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_206_ (
  .in1({ 1'b0 }),
  .out1({ S205 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_207_ (
  .in1({ 1'b0 }),
  .out1({ S206 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_208_ (
  .in1({ 1'b0 }),
  .out1({ S207 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_209_ (
  .in1({ 1'b0 }),
  .out1({ S208 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_210_ (
  .in1({ 1'b0 }),
  .out1({ S209 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_211_ (
  .in1({ 1'b0 }),
  .out1({ S210 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_212_ (
  .in1({ 1'b0 }),
  .out1({ S211 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_213_ (
  .in1({ 1'b0 }),
  .out1({ S212 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_214_ (
  .in1({ 1'b0 }),
  .out1({ S213 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_215_ (
  .in1({ 1'b0 }),
  .out1({ S214 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_216_ (
  .in1({ 1'b0 }),
  .out1({ S215 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_217_ (
  .in1({ 1'b0 }),
  .out1({ S216 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_218_ (
  .in1({ 1'b0 }),
  .out1({ S217 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_219_ (
  .in1({ 1'b0 }),
  .out1({ S218 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_220_ (
  .in1({ 1'b0 }),
  .out1({ S219 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_221_ (
  .in1({ 1'b0 }),
  .out1({ S220 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_222_ (
  .in1({ 1'b0 }),
  .out1({ S221 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_223_ (
  .in1({ 1'b0 }),
  .out1({ S222 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_224_ (
  .in1({ 1'b0 }),
  .out1({ S223 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_225_ (
  .in1({ 1'b0 }),
  .out1({ S224 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_226_ (
  .in1({ 1'b0 }),
  .out1({ S225 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_227_ (
  .in1({ 1'b0 }),
  .out1({ S226 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_228_ (
  .in1({ 1'b0 }),
  .out1({ S227 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_229_ (
  .in1({ 1'b0 }),
  .out1({ S228 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_230_ (
  .in1({ 1'b0 }),
  .out1({ S229 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_231_ (
  .in1({ 1'b0 }),
  .out1({ S230 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_232_ (
  .in1({ 1'b0 }),
  .out1({ S231 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_233_ (
  .in1({ 1'b0 }),
  .out1({ S232 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_234_ (
  .in1({ 1'b0 }),
  .out1({ S233 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_235_ (
  .in1({ 1'b0 }),
  .out1({ S234 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_236_ (
  .in1({ 1'b0 }),
  .out1({ S235 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_237_ (
  .in1({ 1'b0 }),
  .out1({ S236 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_238_ (
  .in1({ 1'b0 }),
  .out1({ S237 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_239_ (
  .in1({ 1'b0 }),
  .out1({ S238 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_240_ (
  .in1({ 1'b0 }),
  .out1({ S239 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_241_ (
  .in1({ 1'b0 }),
  .out1({ S240 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_242_ (
  .in1({ 1'b0 }),
  .out1({ S241 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_243_ (
  .in1({ 1'b0 }),
  .out1({ S242 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_244_ (
  .in1({ 1'b0 }),
  .out1({ S243 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_245_ (
  .in1({ 1'b0 }),
  .out1({ S244 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_246_ (
  .in1({ 1'b0 }),
  .out1({ S245 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_247_ (
  .in1({ 1'b0 }),
  .out1({ S246 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_248_ (
  .in1({ 1'b0 }),
  .out1({ S247 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_249_ (
  .in1({ 1'b0 }),
  .out1({ S248 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_250_ (
  .in1({ 1'b0 }),
  .out1({ S249 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_251_ (
  .in1({ 1'b0 }),
  .out1({ S250 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_252_ (
  .in1({ 1'b0 }),
  .out1({ S251 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_253_ (
  .in1({ 1'b0 }),
  .out1({ S252 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_254_ (
  .in1({ 1'b0 }),
  .out1({ S253 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_255_ (
  .in1({ 1'b0 }),
  .out1({ S254 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_256_ (
  .in1({ 1'b0 }),
  .out1({ S255 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_257_ (
  .in1({ 1'b0 }),
  .out1({ S256 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_258_ (
  .in1({ 1'b0 }),
  .out1({ S257 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_259_ (
  .in1({ 1'b0 }),
  .out1({ S258 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_260_ (
  .in1({ 1'b0 }),
  .out1({ S259 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_261_ (
  .in1({ 1'b0 }),
  .out1({ S260 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_262_ (
  .in1({ 1'b0 }),
  .out1({ S261 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_263_ (
  .in1({ 1'b0 }),
  .out1({ S262 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_264_ (
  .in1({ 1'b0 }),
  .out1({ S263 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_265_ (
  .in1({ 1'b0 }),
  .out1({ S264 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_266_ (
  .in1({ 1'b0 }),
  .out1({ S265 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_267_ (
  .in1({ 1'b0 }),
  .out1({ S266 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_268_ (
  .in1({ 1'b0 }),
  .out1({ S267 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_269_ (
  .in1({ 1'b0 }),
  .out1({ S268 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_270_ (
  .in1({ 1'b0 }),
  .out1({ S269 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_271_ (
  .in1({ 1'b0 }),
  .out1({ S270 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_272_ (
  .in1({ 1'b0 }),
  .out1({ S271 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_273_ (
  .in1({ 1'b0 }),
  .out1({ S272 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_274_ (
  .in1({ 1'b0 }),
  .out1({ S273 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_275_ (
  .in1({ 1'b0 }),
  .out1({ S274 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_276_ (
  .in1({ 1'b0 }),
  .out1({ S275 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_277_ (
  .in1({ 1'b0 }),
  .out1({ S276 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_278_ (
  .in1({ 1'b0 }),
  .out1({ S277 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_279_ (
  .in1({ 1'b0 }),
  .out1({ S278 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_280_ (
  .in1({ 1'b0 }),
  .out1({ S279 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_281_ (
  .in1({ 1'b0 }),
  .out1({ S280 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_282_ (
  .in1({ 1'b0 }),
  .out1({ S281 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_283_ (
  .in1({ 1'b0 }),
  .out1({ S282 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_284_ (
  .in1({ 1'b0 }),
  .out1({ S283 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_285_ (
  .in1({ 1'b0 }),
  .out1({ S284 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_286_ (
  .in1({ 1'b0 }),
  .out1({ S285 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_287_ (
  .in1({ 1'b0 }),
  .out1({ S286 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_288_ (
  .in1({ 1'b0 }),
  .out1({ S287 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_289_ (
  .in1({ 1'b0 }),
  .out1({ S288 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_290_ (
  .in1({ 1'b0 }),
  .out1({ S289 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_291_ (
  .in1({ 1'b0 }),
  .out1({ S290 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_292_ (
  .in1({ 1'b0 }),
  .out1({ S291 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_293_ (
  .in1({ 1'b0 }),
  .out1({ S292 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_294_ (
  .in1({ 1'b0 }),
  .out1({ S293 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_295_ (
  .in1({ 1'b0 }),
  .out1({ S294 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_296_ (
  .in1({ 1'b0 }),
  .out1({ S295 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_297_ (
  .in1({ 1'b0 }),
  .out1({ S296 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_298_ (
  .in1({ 1'b0 }),
  .out1({ S297 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_299_ (
  .in1({ 1'b0 }),
  .out1({ S298 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_300_ (
  .in1({ 1'b0 }),
  .out1({ S299 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_301_ (
  .in1({ 1'b0 }),
  .out1({ S300 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_302_ (
  .in1({ 1'b0 }),
  .out1({ S301 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_303_ (
  .in1({ 1'b0 }),
  .out1({ S302 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_304_ (
  .in1({ 1'b0 }),
  .out1({ S303 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_305_ (
  .in1({ 1'b0 }),
  .out1({ S304 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_306_ (
  .in1({ 1'b0 }),
  .out1({ S305 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_307_ (
  .in1({ 1'b0 }),
  .out1({ S306 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_308_ (
  .in1({ 1'b0 }),
  .out1({ S307 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_309_ (
  .in1({ 1'b0 }),
  .out1({ S308 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_310_ (
  .in1({ 1'b0 }),
  .out1({ S309 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_311_ (
  .in1({ 1'b0 }),
  .out1({ S310 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_312_ (
  .in1({ 1'b0 }),
  .out1({ S311 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_313_ (
  .in1({ 1'b0 }),
  .out1({ S312 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_314_ (
  .in1({ 1'b0 }),
  .out1({ S313 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_315_ (
  .in1({ 1'b0 }),
  .out1({ S314 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_316_ (
  .in1({ 1'b0 }),
  .out1({ S315 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_317_ (
  .in1({ 1'b0 }),
  .out1({ S316 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_318_ (
  .in1({ 1'b0 }),
  .out1({ S317 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_319_ (
  .in1({ 1'b0 }),
  .out1({ S318 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_320_ (
  .in1({ 1'b0 }),
  .out1({ S319 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_321_ (
  .in1({ 1'b0 }),
  .out1({ S320 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_322_ (
  .in1({ 1'b0 }),
  .out1({ S321 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_323_ (
  .in1({ 1'b0 }),
  .out1({ S322 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_324_ (
  .in1({ 1'b0 }),
  .out1({ S323 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_325_ (
  .in1({ 1'b0 }),
  .out1({ S324 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_326_ (
  .in1({ 1'b0 }),
  .out1({ S325 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_327_ (
  .in1({ 1'b0 }),
  .out1({ S326 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_328_ (
  .in1({ 1'b0 }),
  .out1({ S327 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_329_ (
  .in1({ 1'b0 }),
  .out1({ S328 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_330_ (
  .in1({ 1'b0 }),
  .out1({ S329 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_331_ (
  .in1({ 1'b0 }),
  .out1({ S330 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_332_ (
  .in1({ 1'b0 }),
  .out1({ S331 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_333_ (
  .in1({ 1'b0 }),
  .out1({ S332 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_334_ (
  .in1({ 1'b0 }),
  .out1({ S333 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_335_ (
  .in1({ 1'b0 }),
  .out1({ S334 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_336_ (
  .in1({ 1'b0 }),
  .out1({ S335 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_337_ (
  .in1({ 1'b0 }),
  .out1({ S336 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_338_ (
  .in1({ 1'b0 }),
  .out1({ S337 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_339_ (
  .in1({ 1'b0 }),
  .out1({ S338 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_340_ (
  .in1({ 1'b0 }),
  .out1({ S339 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_341_ (
  .in1({ 1'b0 }),
  .out1({ S340 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_342_ (
  .in1({ 1'b0 }),
  .out1({ S341 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_343_ (
  .in1({ 1'b0 }),
  .out1({ S342 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_344_ (
  .in1({ 1'b0 }),
  .out1({ S343 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_345_ (
  .in1({ 1'b0 }),
  .out1({ S344 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_346_ (
  .in1({ 1'b0 }),
  .out1({ S345 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_347_ (
  .in1({ 1'b0 }),
  .out1({ S346 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_348_ (
  .in1({ 1'b0 }),
  .out1({ S347 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_349_ (
  .in1({ 1'b0 }),
  .out1({ S348 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_350_ (
  .in1({ 1'b0 }),
  .out1({ S349 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_351_ (
  .in1({ 1'b0 }),
  .out1({ S350 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_352_ (
  .in1({ 1'b0 }),
  .out1({ S351 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_353_ (
  .in1({ 1'b0 }),
  .out1({ S352 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_354_ (
  .in1({ 1'b0 }),
  .out1({ S353 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_355_ (
  .in1({ 1'b0 }),
  .out1({ S354 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_356_ (
  .in1({ 1'b0 }),
  .out1({ S355 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_357_ (
  .in1({ 1'b0 }),
  .out1({ S356 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_358_ (
  .in1({ 1'b0 }),
  .out1({ S357 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_359_ (
  .in1({ 1'b0 }),
  .out1({ S358 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_360_ (
  .in1({ 1'b0 }),
  .out1({ S359 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_361_ (
  .in1({ 1'b0 }),
  .out1({ S360 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_362_ (
  .in1({ 1'b0 }),
  .out1({ S361 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_363_ (
  .in1({ 1'b0 }),
  .out1({ S362 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_364_ (
  .in1({ 1'b0 }),
  .out1({ S363 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_365_ (
  .in1({ 1'b0 }),
  .out1({ S364 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_366_ (
  .in1({ 1'b0 }),
  .out1({ S365 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_367_ (
  .in1({ 1'b0 }),
  .out1({ S366 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_368_ (
  .in1({ 1'b0 }),
  .out1({ S367 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_369_ (
  .in1({ 1'b0 }),
  .out1({ S368 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_370_ (
  .in1({ 1'b0 }),
  .out1({ S369 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_371_ (
  .in1({ 1'b0 }),
  .out1({ S370 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_372_ (
  .in1({ 1'b0 }),
  .out1({ S371 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_373_ (
  .in1({ 1'b0 }),
  .out1({ S372 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_374_ (
  .in1({ 1'b0 }),
  .out1({ S373 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_375_ (
  .in1({ 1'b0 }),
  .out1({ S374 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_376_ (
  .in1({ 1'b0 }),
  .out1({ S375 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_377_ (
  .in1({ 1'b0 }),
  .out1({ S376 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_378_ (
  .in1({ 1'b0 }),
  .out1({ S377 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_379_ (
  .in1({ 1'b0 }),
  .out1({ S378 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_380_ (
  .in1({ 1'b0 }),
  .out1({ S379 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_381_ (
  .in1({ 1'b0 }),
  .out1({ S380 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_382_ (
  .in1({ 1'b0 }),
  .out1({ S381 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_383_ (
  .in1({ 1'b0 }),
  .out1({ S382 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_384_ (
  .in1({ 1'b0 }),
  .out1({ S383 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_385_ (
  .in1({ 1'b0 }),
  .out1({ S384 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_386_ (
  .in1({ 1'b0 }),
  .out1({ S385 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_387_ (
  .in1({ 1'b0 }),
  .out1({ S386 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_388_ (
  .in1({ 1'b0 }),
  .out1({ S387 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_389_ (
  .in1({ 1'b0 }),
  .out1({ S388 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_390_ (
  .in1({ 1'b0 }),
  .out1({ S389 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_391_ (
  .in1({ 1'b0 }),
  .out1({ S390 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_392_ (
  .in1({ 1'b0 }),
  .out1({ S391 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_393_ (
  .in1({ 1'b0 }),
  .out1({ S392 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_394_ (
  .in1({ 1'b0 }),
  .out1({ S393 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_395_ (
  .in1({ 1'b0 }),
  .out1({ S394 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_396_ (
  .in1({ 1'b0 }),
  .out1({ S395 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_397_ (
  .in1({ 1'b0 }),
  .out1({ S396 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_398_ (
  .in1({ 1'b0 }),
  .out1({ S397 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_399_ (
  .in1({ 1'b0 }),
  .out1({ S398 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_400_ (
  .in1({ 1'b0 }),
  .out1({ S399 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_401_ (
  .in1({ 1'b0 }),
  .out1({ S400 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_402_ (
  .in1({ 1'b0 }),
  .out1({ S401 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_403_ (
  .in1({ 1'b0 }),
  .out1({ S402 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_404_ (
  .in1({ 1'b0 }),
  .out1({ S403 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_405_ (
  .in1({ 1'b0 }),
  .out1({ S404 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_406_ (
  .in1({ 1'b0 }),
  .out1({ S405 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_407_ (
  .in1({ 1'b0 }),
  .out1({ S406 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_408_ (
  .in1({ 1'b0 }),
  .out1({ S407 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_409_ (
  .in1({ 1'b0 }),
  .out1({ S408 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_410_ (
  .in1({ 1'b0 }),
  .out1({ S409 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_411_ (
  .in1({ 1'b0 }),
  .out1({ S410 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_412_ (
  .in1({ 1'b0 }),
  .out1({ S411 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_413_ (
  .in1({ 1'b0 }),
  .out1({ S412 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_414_ (
  .in1({ 1'b0 }),
  .out1({ S413 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_415_ (
  .in1({ 1'b0 }),
  .out1({ S414 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_416_ (
  .in1({ 1'b0 }),
  .out1({ S415 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_417_ (
  .in1({ 1'b0 }),
  .out1({ S416 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_418_ (
  .in1({ 1'b0 }),
  .out1({ S417 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_419_ (
  .in1({ 1'b0 }),
  .out1({ S418 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_420_ (
  .in1({ 1'b0 }),
  .out1({ S419 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_421_ (
  .in1({ 1'b0 }),
  .out1({ S420 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_422_ (
  .in1({ 1'b0 }),
  .out1({ S421 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_423_ (
  .in1({ 1'b0 }),
  .out1({ S422 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_424_ (
  .in1({ 1'b0 }),
  .out1({ S423 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_425_ (
  .in1({ 1'b0 }),
  .out1({ S424 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_426_ (
  .in1({ 1'b0 }),
  .out1({ S425 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_427_ (
  .in1({ 1'b0 }),
  .out1({ S426 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_428_ (
  .in1({ 1'b0 }),
  .out1({ S427 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_429_ (
  .in1({ 1'b0 }),
  .out1({ S428 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_430_ (
  .in1({ 1'b0 }),
  .out1({ S429 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_431_ (
  .in1({ 1'b0 }),
  .out1({ S430 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_432_ (
  .in1({ 1'b0 }),
  .out1({ S431 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_433_ (
  .in1({ 1'b0 }),
  .out1({ S432 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_434_ (
  .in1({ 1'b0 }),
  .out1({ S433 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_435_ (
  .in1({ 1'b0 }),
  .out1({ S434 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_436_ (
  .in1({ 1'b0 }),
  .out1({ S435 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_437_ (
  .in1({ 1'b0 }),
  .out1({ S436 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_438_ (
  .in1({ 1'b0 }),
  .out1({ S437 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_439_ (
  .in1({ 1'b0 }),
  .out1({ S438 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_440_ (
  .in1({ 1'b0 }),
  .out1({ S439 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_441_ (
  .in1({ 1'b0 }),
  .out1({ S440 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_442_ (
  .in1({ 1'b0 }),
  .out1({ S441 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_443_ (
  .in1({ 1'b0 }),
  .out1({ S442 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_444_ (
  .in1({ 1'b0 }),
  .out1({ S443 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_445_ (
  .in1({ 1'b0 }),
  .out1({ S444 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_446_ (
  .in1({ 1'b0 }),
  .out1({ S445 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_447_ (
  .in1({ 1'b0 }),
  .out1({ S446 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_448_ (
  .in1({ 1'b0 }),
  .out1({ S447 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_449_ (
  .in1({ 1'b0 }),
  .out1({ S448 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_450_ (
  .in1({ 1'b0 }),
  .out1({ S449 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_451_ (
  .in1({ 1'b0 }),
  .out1({ S450 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_452_ (
  .in1({ 1'b0 }),
  .out1({ S451 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_453_ (
  .in1({ 1'b0 }),
  .out1({ S452 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_454_ (
  .in1({ 1'b0 }),
  .out1({ S453 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_455_ (
  .in1({ 1'b0 }),
  .out1({ S454 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_456_ (
  .in1({ 1'b0 }),
  .out1({ S455 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_457_ (
  .in1({ 1'b0 }),
  .out1({ S456 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_458_ (
  .in1({ 1'b0 }),
  .out1({ S457 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_459_ (
  .in1({ 1'b0 }),
  .out1({ S458 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_460_ (
  .in1({ 1'b0 }),
  .out1({ S459 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_461_ (
  .in1({ 1'b0 }),
  .out1({ S460 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_462_ (
  .in1({ 1'b0 }),
  .out1({ S461 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_463_ (
  .in1({ 1'b0 }),
  .out1({ S462 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_464_ (
  .in1({ 1'b0 }),
  .out1({ S463 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_465_ (
  .in1({ 1'b0 }),
  .out1({ S464 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_466_ (
  .in1({ 1'b0 }),
  .out1({ S465 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_467_ (
  .in1({ 1'b0 }),
  .out1({ S466 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_468_ (
  .in1({ 1'b0 }),
  .out1({ S467 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_469_ (
  .in1({ 1'b0 }),
  .out1({ S468 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_470_ (
  .in1({ 1'b0 }),
  .out1({ S469 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_471_ (
  .in1({ 1'b0 }),
  .out1({ S470 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_472_ (
  .in1({ 1'b0 }),
  .out1({ S471 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_473_ (
  .in1({ 1'b0 }),
  .out1({ S472 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_474_ (
  .in1({ 1'b0 }),
  .out1({ S473 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_475_ (
  .in1({ 1'b0 }),
  .out1({ S474 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_476_ (
  .in1({ 1'b0 }),
  .out1({ S475 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_477_ (
  .in1({ 1'b0 }),
  .out1({ S476 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_478_ (
  .in1({ 1'b0 }),
  .out1({ S477 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_479_ (
  .in1({ 1'b0 }),
  .out1({ S478 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_480_ (
  .in1({ 1'b0 }),
  .out1({ S479 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_481_ (
  .in1({ 1'b0 }),
  .out1({ S480 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_482_ (
  .in1({ 1'b0 }),
  .out1({ S481 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_483_ (
  .in1({ 1'b0 }),
  .out1({ S482 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_484_ (
  .in1({ 1'b0 }),
  .out1({ S483 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_485_ (
  .in1({ 1'b0 }),
  .out1({ S484 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_486_ (
  .in1({ 1'b0 }),
  .out1({ S485 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_487_ (
  .in1({ 1'b0 }),
  .out1({ S486 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_488_ (
  .in1({ 1'b0 }),
  .out1({ S487 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_489_ (
  .in1({ 1'b0 }),
  .out1({ S488 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_490_ (
  .in1({ 1'b0 }),
  .out1({ S489 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_491_ (
  .in1({ 1'b0 }),
  .out1({ S490 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_492_ (
  .in1({ 1'b0 }),
  .out1({ S491 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_493_ (
  .in1({ 1'b0 }),
  .out1({ S492 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_494_ (
  .in1({ 1'b0 }),
  .out1({ S493 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_495_ (
  .in1({ 1'b0 }),
  .out1({ S494 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_496_ (
  .in1({ 1'b0 }),
  .out1({ S495 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_497_ (
  .in1({ 1'b0 }),
  .out1({ S496 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_498_ (
  .in1({ 1'b0 }),
  .out1({ S497 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_499_ (
  .in1({ 1'b0 }),
  .out1({ S498 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_500_ (
  .in1({ 1'b0 }),
  .out1({ S499 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_501_ (
  .in1({ 1'b0 }),
  .out1({ S500 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_502_ (
  .in1({ 1'b0 }),
  .out1({ S501 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_503_ (
  .in1({ 1'b0 }),
  .out1({ S502 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_504_ (
  .in1({ 1'b0 }),
  .out1({ S503 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_505_ (
  .in1({ 1'b0 }),
  .out1({ S504 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_1_ (
  .in1({ DP_SR_V_dout }),
  .out1({ S505 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_2_ (
  .in1({ DP_SR_C_dout }),
  .out1({ S506 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_3_ (
  .in1({ DP_SR_N_dout }),
  .out1({ S507 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_4_ (
  .in1({ DP_SR_Z_dout }),
  .out1({ S508 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1_ (
  .in1({ S507, CU_inst_2 }),
  .out1({ S509 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1_ (
  .in1({ S507, CU_inst_2 }),
  .out1({ S510 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_2_ (
  .in1({ S510, CU_inst_6 }),
  .out1({ S511 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_2_ (
  .in1({ S511, S509 }),
  .out1({ S512 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_3_ (
  .in1({ S508, CU_inst_3 }),
  .out1({ S513 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_3_ (
  .in1({ S508, CU_inst_3 }),
  .out1({ S514 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_4_ (
  .in1({ S514, CU_inst_7 }),
  .out1({ S515 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_4_ (
  .in1({ S515, S513 }),
  .out1({ S516 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_5_ (
  .in1({ S516, S512 }),
  .out1({ S517 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_6_ (
  .in1({ S505, CU_inst_0 }),
  .out1({ S518 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_5_ (
  .in1({ S505, CU_inst_0 }),
  .out1({ S519 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_6_ (
  .in1({ S519, CU_inst_4 }),
  .out1({ S520 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_7_ (
  .in1({ S520, S518 }),
  .out1({ S521 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_8_ (
  .in1({ S506, CU_inst_1 }),
  .out1({ S522 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_7_ (
  .in1({ S506, CU_inst_1 }),
  .out1({ S523 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_8_ (
  .in1({ S523, CU_inst_5 }),
  .out1({ S524 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_9_ (
  .in1({ S524, S522 }),
  .out1({ S525 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_10_ (
  .in1({ S525, S521 }),
  .out1({ S526 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_9_ (
  .in1({ S526, S517 }),
  .out1({ CU_enSKP })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_5_ (
  .in1({ S42 }),
  .out1({ S544 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_11_ (
  .in1({ S44, S43 }),
  .out1({ S545 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_10_ (
  .in1({ S545, DP_AC_dout_0 }),
  .out1({ S546 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_12_ (
  .in1({ S544, S45 }),
  .out1({ S547 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_11_ (
  .in1({ S547, DP_AC_din_0 }),
  .out1({ S548 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_12_ (
  .in1({ S548, S546 }),
  .out1({ S527 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_13_ (
  .in1({ S545, DP_AC_dout_1 }),
  .out1({ S549 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_14_ (
  .in1({ S547, DP_AC_din_1 }),
  .out1({ S550 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_15_ (
  .in1({ S550, S549 }),
  .out1({ S528 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_16_ (
  .in1({ S545, DP_AC_dout_2 }),
  .out1({ S551 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_17_ (
  .in1({ S547, DP_AC_din_2 }),
  .out1({ S552 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_18_ (
  .in1({ S552, S551 }),
  .out1({ S529 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_19_ (
  .in1({ S545, DP_AC_dout_3 }),
  .out1({ S553 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_20_ (
  .in1({ S547, DP_AC_din_3 }),
  .out1({ S554 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_21_ (
  .in1({ S554, S553 }),
  .out1({ S530 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_22_ (
  .in1({ S545, DP_AC_dout_4 }),
  .out1({ S555 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_23_ (
  .in1({ S547, DP_AC_din_4 }),
  .out1({ S556 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_24_ (
  .in1({ S556, S555 }),
  .out1({ S531 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_25_ (
  .in1({ S545, DP_AC_dout_5 }),
  .out1({ S557 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_26_ (
  .in1({ S547, DP_AC_din_5 }),
  .out1({ S558 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_27_ (
  .in1({ S558, S557 }),
  .out1({ S532 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_28_ (
  .in1({ S545, DP_AC_dout_6 }),
  .out1({ S559 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_29_ (
  .in1({ S547, DP_AC_din_6 }),
  .out1({ S560 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_30_ (
  .in1({ S560, S559 }),
  .out1({ S533 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_31_ (
  .in1({ S545, DP_AC_dout_7 }),
  .out1({ S561 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_32_ (
  .in1({ S547, DP_AC_din_7 }),
  .out1({ S562 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_33_ (
  .in1({ S562, S561 }),
  .out1({ S534 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_34_ (
  .in1({ S545, DP_AC_dout_8 }),
  .out1({ S563 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_35_ (
  .in1({ S547, DP_AC_din_8 }),
  .out1({ S564 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_36_ (
  .in1({ S564, S563 }),
  .out1({ S535 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_37_ (
  .in1({ S545, DP_AC_dout_9 }),
  .out1({ S565 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_38_ (
  .in1({ S547, DP_AC_din_9 }),
  .out1({ S566 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_39_ (
  .in1({ S566, S565 }),
  .out1({ S536 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_40_ (
  .in1({ S545, DP_AC_dout_10 }),
  .out1({ S567 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_41_ (
  .in1({ S547, DP_AC_din_10 }),
  .out1({ S568 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_42_ (
  .in1({ S568, S567 }),
  .out1({ S537 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_43_ (
  .in1({ S545, DP_AC_dout_11 }),
  .out1({ S569 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_44_ (
  .in1({ S547, DP_AC_din_11 }),
  .out1({ S570 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_45_ (
  .in1({ S570, S569 }),
  .out1({ S538 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_46_ (
  .in1({ S545, DP_AC_dout_12 }),
  .out1({ S571 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_47_ (
  .in1({ S547, DP_AC_din_12 }),
  .out1({ S572 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_48_ (
  .in1({ S572, S571 }),
  .out1({ S539 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_49_ (
  .in1({ S545, DP_AC_dout_13 }),
  .out1({ S573 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_50_ (
  .in1({ S547, DP_AC_din_13 }),
  .out1({ S574 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_51_ (
  .in1({ S574, S573 }),
  .out1({ S540 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_52_ (
  .in1({ S545, DP_AC_dout_14 }),
  .out1({ S575 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_53_ (
  .in1({ S547, DP_AC_din_14 }),
  .out1({ S576 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_54_ (
  .in1({ S576, S575 }),
  .out1({ S541 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_55_ (
  .in1({ S545, DP_AC_dout_15 }),
  .out1({ S577 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_56_ (
  .in1({ S547, DP_AC_din_15 }),
  .out1({ S543 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_57_ (
  .in1({ S543, S577 }),
  .out1({ S542 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_1_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S527 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_dout_0 }),
  .Si({ S3375 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_2_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S528 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_dout_1 }),
  .Si({ S3374 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_3_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S529 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_dout_2 }),
  .Si({ S3373 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_4_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S530 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_dout_3 }),
  .Si({ S3372 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_5_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S531 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_dout_4 }),
  .Si({ S3371 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_6_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S532 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_dout_5 }),
  .Si({ S3370 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_7_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S533 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_dout_6 }),
  .Si({ S3369 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_8_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S534 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_dout_7 }),
  .Si({ S3368 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_9_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S535 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_dout_8 }),
  .Si({ S3367 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_10_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S536 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_dout_9 }),
  .Si({ S3366 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_11_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S537 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_dout_10 }),
  .Si({ S3365 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_12_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S538 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_dout_11 }),
  .Si({ S3364 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_13_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S539 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_dout_12 }),
  .Si({ S3363 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_14_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S540 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_dout_13 }),
  .Si({ S3362 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_15_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S541 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_dout_14 }),
  .Si({ S3361 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_16_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S542 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_AC_dout_15 }),
  .Si({ S3424 }),
  .global_reset({ 1'b0 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_6_ (
  .in1({ DP_AC_dout_0 }),
  .out1({ S1099 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_7_ (
  .in1({ DP_ARU1_in1_0 }),
  .out1({ S1109 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_8_ (
  .in1({ S46 }),
  .out1({ S1120 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_9_ (
  .in1({ S47 }),
  .out1({ S1131 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_10_ (
  .in1({ DP_ARU1_in1_1 }),
  .out1({ S1142 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_11_ (
  .in1({ DP_AC_dout_1 }),
  .out1({ S1153 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_12_ (
  .in1({ DP_ARU1_in1_2 }),
  .out1({ S1164 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_13_ (
  .in1({ DP_AC_dout_2 }),
  .out1({ S1175 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_14_ (
  .in1({ DP_AC_dout_3 }),
  .out1({ S1186 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_15_ (
  .in1({ DP_ARU1_in1_3 }),
  .out1({ S1197 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_16_ (
  .in1({ DP_ARU1_in1_4 }),
  .out1({ S1208 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_17_ (
  .in1({ DP_AC_dout_4 }),
  .out1({ S1218 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_18_ (
  .in1({ DP_ARU1_in1_5 }),
  .out1({ S1229 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_19_ (
  .in1({ DP_AC_dout_5 }),
  .out1({ S1240 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_20_ (
  .in1({ DP_ARU1_in1_6 }),
  .out1({ S1251 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_21_ (
  .in1({ DP_AC_dout_6 }),
  .out1({ S1262 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_22_ (
  .in1({ DP_ARU1_in1_7 }),
  .out1({ S1273 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_23_ (
  .in1({ DP_AC_dout_7 }),
  .out1({ S1284 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_24_ (
  .in1({ DP_AC_dout_11 }),
  .out1({ S1295 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_25_ (
  .in1({ DP_ARU1_in1_11 }),
  .out1({ S1306 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_26_ (
  .in1({ DP_AC_dout_15 }),
  .out1({ S1316 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_27_ (
  .in1({ DP_ARU1_in1_15 }),
  .out1({ S1327 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_13_ (
  .in1({ DP_ARU1_in1_0, DP_AC_dout_0 }),
  .out1({ S1338 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_28_ (
  .in1({ S1338 }),
  .out1({ S1349 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_14_ (
  .in1({ S1109, S1099 }),
  .out1({ S1360 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_58_ (
  .in1({ DP_ARU1_in1_0, DP_AC_dout_0 }),
  .out1({ S1371 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_59_ (
  .in1({ S1371, S48 }),
  .out1({ S1382 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_15_ (
  .in1({ S49, S1120 }),
  .out1({ S1393 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_60_ (
  .in1({ S1131, S50 }),
  .out1({ S1404 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_61_ (
  .in1({ S1393, S1360 }),
  .out1({ S1414 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_62_ (
  .in1({ S1414, S1382 }),
  .out1({ S1425 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_63_ (
  .in1({ S1425, S1349 }),
  .out1({ S1436 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_29_ (
  .in1({ S1436 }),
  .out1({ DP_ARU1_out_0 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_16_ (
  .in1({ S1153, S1142 }),
  .out1({ S1457 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_64_ (
  .in1({ DP_AC_dout_1, DP_ARU1_in1_1 }),
  .out1({ S1468 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_17_ (
  .in1({ DP_AC_dout_1, DP_ARU1_in1_1 }),
  .out1({ S1479 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_18_ (
  .in1({ S1479, S1457 }),
  .out1({ S1489 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_19_ (
  .in1({ S1489, S1360 }),
  .out1({ S1500 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_65_ (
  .in1({ S1489, S1360 }),
  .out1({ S1511 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_66_ (
  .in1({ S1511, S51 }),
  .out1({ S1522 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_20_ (
  .in1({ S1522, S1500 }),
  .out1({ S1533 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_67_ (
  .in1({ DP_AC_dout_1, DP_ARU1_in1_0 }),
  .out1({ S1544 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_30_ (
  .in1({ S1544 }),
  .out1({ S1555 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_68_ (
  .in1({ DP_ARU1_in1_1, DP_AC_dout_0 }),
  .out1({ S1565 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_31_ (
  .in1({ S1565 }),
  .out1({ S1576 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_69_ (
  .in1({ S1565, S1544 }),
  .out1({ S1587 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_21_ (
  .in1({ S1468, S1371 }),
  .out1({ S588 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_70_ (
  .in1({ S1587, S1393 }),
  .out1({ S598 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_22_ (
  .in1({ S598, S588 }),
  .out1({ S609 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_23_ (
  .in1({ S609, S1533 }),
  .out1({ S620 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_32_ (
  .in1({ S620 }),
  .out1({ DP_ARU1_out_1 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_71_ (
  .in1({ S1511, S1468 }),
  .out1({ S640 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_24_ (
  .in1({ S1175, S1164 }),
  .out1({ S650 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_72_ (
  .in1({ DP_AC_dout_2, DP_ARU1_in1_2 }),
  .out1({ S659 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_25_ (
  .in1({ DP_AC_dout_2, DP_ARU1_in1_2 }),
  .out1({ S662 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_26_ (
  .in1({ S662, S650 }),
  .out1({ S663 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_27_ (
  .in1({ S663, S640 }),
  .out1({ S664 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_73_ (
  .in1({ S663, S640 }),
  .out1({ S665 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_28_ (
  .in1({ S664, S1131 }),
  .out1({ S666 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_74_ (
  .in1({ S666, S665 }),
  .out1({ S667 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_75_ (
  .in1({ DP_AC_dout_2, DP_ARU1_in1_0 }),
  .out1({ S668 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_33_ (
  .in1({ S668 }),
  .out1({ S669 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_29_ (
  .in1({ S1164, S1099 }),
  .out1({ S670 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_76_ (
  .in1({ DP_ARU1_in1_2, DP_AC_dout_0 }),
  .out1({ S671 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_77_ (
  .in1({ S671, S1468 }),
  .out1({ S672 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_78_ (
  .in1({ DP_ARU1_in1_2, DP_AC_dout_1 }),
  .out1({ S673 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_30_ (
  .in1({ S671, S1468 }),
  .out1({ S674 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_79_ (
  .in1({ S670, S1457 }),
  .out1({ S675 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_80_ (
  .in1({ S675, S672 }),
  .out1({ S676 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_34_ (
  .in1({ S676 }),
  .out1({ S677 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_81_ (
  .in1({ S677, S669 }),
  .out1({ S678 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_82_ (
  .in1({ S676, S668 }),
  .out1({ S679 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_83_ (
  .in1({ S679, S678 }),
  .out1({ S680 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_35_ (
  .in1({ S680 }),
  .out1({ S681 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_31_ (
  .in1({ S681, S588 }),
  .out1({ S682 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_84_ (
  .in1({ S681, S588 }),
  .out1({ S683 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_36_ (
  .in1({ S683 }),
  .out1({ S684 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_32_ (
  .in1({ S684, S682 }),
  .out1({ S685 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_85_ (
  .in1({ S685, S1393 }),
  .out1({ S686 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_86_ (
  .in1({ S686, S667 }),
  .out1({ DP_ARU1_out_2 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_87_ (
  .in1({ DP_ARU1_in1_3, DP_AC_dout_0 }),
  .out1({ S687 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_88_ (
  .in1({ DP_AC_dout_3, DP_ARU1_in1_0 }),
  .out1({ S688 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_33_ (
  .in1({ S1197, S1186 }),
  .out1({ S689 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_89_ (
  .in1({ DP_ARU1_in1_3, DP_AC_dout_3 }),
  .out1({ S690 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_34_ (
  .in1({ S690, S1371 }),
  .out1({ S691 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_90_ (
  .in1({ S689, S1360 }),
  .out1({ S692 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_91_ (
  .in1({ S688, S687 }),
  .out1({ S693 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_92_ (
  .in1({ S693, S692 }),
  .out1({ S694 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_37_ (
  .in1({ S694 }),
  .out1({ S695 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_93_ (
  .in1({ DP_AC_dout_2, DP_ARU1_in1_1 }),
  .out1({ S696 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_38_ (
  .in1({ S696 }),
  .out1({ S697 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_35_ (
  .in1({ S659, S1468 }),
  .out1({ S698 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_94_ (
  .in1({ S650, S1457 }),
  .out1({ S699 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_95_ (
  .in1({ S696, S673 }),
  .out1({ S700 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_39_ (
  .in1({ S700 }),
  .out1({ S701 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_36_ (
  .in1({ S701, S698 }),
  .out1({ S702 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_96_ (
  .in1({ S700, S699 }),
  .out1({ S703 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_37_ (
  .in1({ S703, S675 }),
  .out1({ S704 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_97_ (
  .in1({ S702, S674 }),
  .out1({ S705 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_98_ (
  .in1({ S703, S675 }),
  .out1({ S706 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_99_ (
  .in1({ S706, S705 }),
  .out1({ S707 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_40_ (
  .in1({ S707 }),
  .out1({ S708 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_100_ (
  .in1({ S707, S694 }),
  .out1({ S709 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_101_ (
  .in1({ S708, S695 }),
  .out1({ S710 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_41_ (
  .in1({ S710 }),
  .out1({ S711 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_102_ (
  .in1({ S710, S709 }),
  .out1({ S712 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_38_ (
  .in1({ S712, S678 }),
  .out1({ S713 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_42_ (
  .in1({ S713 }),
  .out1({ S714 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_103_ (
  .in1({ S712, S678 }),
  .out1({ S715 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_104_ (
  .in1({ S715, S714 }),
  .out1({ S716 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_105_ (
  .in1({ S716, S683 }),
  .out1({ S717 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_39_ (
  .in1({ S716, S683 }),
  .out1({ S718 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_106_ (
  .in1({ S717, S1393 }),
  .out1({ S719 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_40_ (
  .in1({ S719, S718 }),
  .out1({ S720 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_107_ (
  .in1({ S665, S659 }),
  .out1({ S721 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_43_ (
  .in1({ S721 }),
  .out1({ S722 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_41_ (
  .in1({ DP_ARU1_in1_3, DP_AC_dout_3 }),
  .out1({ S723 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_42_ (
  .in1({ S723, S689 }),
  .out1({ S724 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_43_ (
  .in1({ S724, S721 }),
  .out1({ S725 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_108_ (
  .in1({ S724, S721 }),
  .out1({ S726 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_109_ (
  .in1({ S726, S52 }),
  .out1({ S727 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_44_ (
  .in1({ S727, S725 }),
  .out1({ S728 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_45_ (
  .in1({ S728, S720 }),
  .out1({ S729 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_44_ (
  .in1({ S729 }),
  .out1({ DP_ARU1_out_3 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_46_ (
  .in1({ S711, S704 }),
  .out1({ S730 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_110_ (
  .in1({ S710, S705 }),
  .out1({ S731 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_111_ (
  .in1({ DP_ARU1_in1_3, DP_AC_dout_1 }),
  .out1({ S732 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_112_ (
  .in1({ DP_AC_dout_4, DP_ARU1_in1_0 }),
  .out1({ S733 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_47_ (
  .in1({ S1218, S1197 }),
  .out1({ S734 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_113_ (
  .in1({ DP_AC_dout_4, DP_ARU1_in1_3 }),
  .out1({ S735 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_48_ (
  .in1({ S735, S1544 }),
  .out1({ S736 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_114_ (
  .in1({ S734, S1555 }),
  .out1({ S737 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_115_ (
  .in1({ S733, S732 }),
  .out1({ S738 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_45_ (
  .in1({ S738 }),
  .out1({ S739 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_49_ (
  .in1({ S739, S736 }),
  .out1({ S740 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_116_ (
  .in1({ S738, S737 }),
  .out1({ S741 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_117_ (
  .in1({ DP_AC_dout_3, DP_ARU1_in1_1 }),
  .out1({ S742 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_118_ (
  .in1({ DP_ARU1_in1_4, DP_AC_dout_0 }),
  .out1({ S743 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_119_ (
  .in1({ S743, S742 }),
  .out1({ S744 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_46_ (
  .in1({ S744 }),
  .out1({ S745 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_120_ (
  .in1({ DP_ARU1_in1_4, DP_AC_dout_3 }),
  .out1({ S746 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_47_ (
  .in1({ S746 }),
  .out1({ S747 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_50_ (
  .in1({ S746, S1565 }),
  .out1({ S748 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_121_ (
  .in1({ S747, S1576 }),
  .out1({ S749 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_51_ (
  .in1({ S748, S745 }),
  .out1({ S750 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_122_ (
  .in1({ S749, S744 }),
  .out1({ S751 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_52_ (
  .in1({ S659, S1457 }),
  .out1({ S752 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_123_ (
  .in1({ S650, S1468 }),
  .out1({ S753 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_53_ (
  .in1({ S752, S751 }),
  .out1({ S754 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_124_ (
  .in1({ S753, S750 }),
  .out1({ S755 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_54_ (
  .in1({ S753, S750 }),
  .out1({ S756 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_125_ (
  .in1({ S752, S751 }),
  .out1({ S757 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_55_ (
  .in1({ S756, S754 }),
  .out1({ S758 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_126_ (
  .in1({ S757, S755 }),
  .out1({ S759 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_127_ (
  .in1({ S758, S741 }),
  .out1({ S760 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_56_ (
  .in1({ S758, S741 }),
  .out1({ S761 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_128_ (
  .in1({ S759, S740 }),
  .out1({ S762 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_129_ (
  .in1({ S762, S760 }),
  .out1({ S763 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_48_ (
  .in1({ S763 }),
  .out1({ S764 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_130_ (
  .in1({ S764, S731 }),
  .out1({ S765 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_131_ (
  .in1({ S763, S730 }),
  .out1({ S766 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_132_ (
  .in1({ S766, S765 }),
  .out1({ S767 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_49_ (
  .in1({ S767 }),
  .out1({ S768 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_133_ (
  .in1({ S767, S692 }),
  .out1({ S769 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_134_ (
  .in1({ S768, S691 }),
  .out1({ S770 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_135_ (
  .in1({ S770, S769 }),
  .out1({ S771 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_57_ (
  .in1({ S718, S713 }),
  .out1({ S772 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_136_ (
  .in1({ S772, S771 }),
  .out1({ S773 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_58_ (
  .in1({ S772, S771 }),
  .out1({ S774 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_50_ (
  .in1({ S774 }),
  .out1({ S775 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_59_ (
  .in1({ S774, S1404 }),
  .out1({ S776 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_137_ (
  .in1({ S776, S773 }),
  .out1({ S777 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_60_ (
  .in1({ S1218, S1208 }),
  .out1({ S778 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_138_ (
  .in1({ DP_AC_dout_4, DP_ARU1_in1_4 }),
  .out1({ S779 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_61_ (
  .in1({ DP_AC_dout_4, DP_ARU1_in1_4 }),
  .out1({ S780 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_51_ (
  .in1({ S780 }),
  .out1({ S781 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_139_ (
  .in1({ S781, S779 }),
  .out1({ S782 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_62_ (
  .in1({ S723, S722 }),
  .out1({ S783 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_63_ (
  .in1({ S783, S689 }),
  .out1({ S784 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_140_ (
  .in1({ S784, S782 }),
  .out1({ S785 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_64_ (
  .in1({ S784, S782 }),
  .out1({ S786 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_52_ (
  .in1({ S786 }),
  .out1({ S787 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_65_ (
  .in1({ S786, S1131 }),
  .out1({ S788 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_141_ (
  .in1({ S788, S785 }),
  .out1({ S789 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_142_ (
  .in1({ S789, S777 }),
  .out1({ DP_ARU1_out_4 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_143_ (
  .in1({ S787, S779 }),
  .out1({ S790 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_66_ (
  .in1({ S1240, S1229 }),
  .out1({ S791 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_144_ (
  .in1({ DP_AC_dout_5, DP_ARU1_in1_5 }),
  .out1({ S792 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_67_ (
  .in1({ DP_AC_dout_5, DP_ARU1_in1_5 }),
  .out1({ S793 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_68_ (
  .in1({ S793, S791 }),
  .out1({ S794 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_69_ (
  .in1({ S794, S790 }),
  .out1({ S795 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_145_ (
  .in1({ S794, S790 }),
  .out1({ S796 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_146_ (
  .in1({ S796, S53 }),
  .out1({ S797 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_70_ (
  .in1({ S797, S795 }),
  .out1({ S798 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_147_ (
  .in1({ S770, S765 }),
  .out1({ S799 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_53_ (
  .in1({ S799 }),
  .out1({ S800 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_71_ (
  .in1({ S750, S699 }),
  .out1({ S801 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_148_ (
  .in1({ S751, S698 }),
  .out1({ S802 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_72_ (
  .in1({ S801, S761 }),
  .out1({ S803 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_149_ (
  .in1({ S802, S762 }),
  .out1({ S804 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_150_ (
  .in1({ DP_ARU1_in1_3, DP_AC_dout_2 }),
  .out1({ S805 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_151_ (
  .in1({ DP_AC_dout_5, DP_ARU1_in1_0 }),
  .out1({ S806 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_152_ (
  .in1({ DP_AC_dout_5, DP_ARU1_in1_3 }),
  .out1({ S807 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_54_ (
  .in1({ S807 }),
  .out1({ S808 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_73_ (
  .in1({ S807, S668 }),
  .out1({ S809 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_153_ (
  .in1({ S808, S669 }),
  .out1({ S810 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_154_ (
  .in1({ S806, S805 }),
  .out1({ S811 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_55_ (
  .in1({ S811 }),
  .out1({ S812 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_74_ (
  .in1({ S812, S809 }),
  .out1({ S813 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_155_ (
  .in1({ S811, S810 }),
  .out1({ S814 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_75_ (
  .in1({ S751, S659 }),
  .out1({ S815 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_156_ (
  .in1({ S750, S650 }),
  .out1({ S816 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_157_ (
  .in1({ DP_ARU1_in1_5, DP_AC_dout_0 }),
  .out1({ S817 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_158_ (
  .in1({ DP_AC_dout_3, DP_ARU1_in1_2 }),
  .out1({ S818 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_159_ (
  .in1({ S818, S817 }),
  .out1({ S819 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_56_ (
  .in1({ S819 }),
  .out1({ S820 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_160_ (
  .in1({ DP_ARU1_in1_5, DP_AC_dout_3 }),
  .out1({ S821 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_57_ (
  .in1({ S821 }),
  .out1({ S822 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_76_ (
  .in1({ S821, S671 }),
  .out1({ S823 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_161_ (
  .in1({ S822, S670 }),
  .out1({ S824 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_77_ (
  .in1({ S823, S820 }),
  .out1({ S825 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_162_ (
  .in1({ S824, S819 }),
  .out1({ S826 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_163_ (
  .in1({ DP_AC_dout_4, DP_ARU1_in1_1 }),
  .out1({ S827 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_164_ (
  .in1({ DP_ARU1_in1_4, DP_AC_dout_1 }),
  .out1({ S828 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_165_ (
  .in1({ S828, S827 }),
  .out1({ S829 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_58_ (
  .in1({ S829 }),
  .out1({ S830 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_78_ (
  .in1({ S779, S1468 }),
  .out1({ S831 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_166_ (
  .in1({ S778, S1457 }),
  .out1({ S832 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_79_ (
  .in1({ S831, S830 }),
  .out1({ S833 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_167_ (
  .in1({ S832, S829 }),
  .out1({ S834 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_80_ (
  .in1({ S834, S749 }),
  .out1({ S835 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_168_ (
  .in1({ S833, S748 }),
  .out1({ S836 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_81_ (
  .in1({ S833, S748 }),
  .out1({ S837 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_169_ (
  .in1({ S834, S749 }),
  .out1({ S838 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_82_ (
  .in1({ S837, S835 }),
  .out1({ S839 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_170_ (
  .in1({ S838, S836 }),
  .out1({ S840 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_83_ (
  .in1({ S839, S825 }),
  .out1({ S841 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_171_ (
  .in1({ S840, S826 }),
  .out1({ S842 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_84_ (
  .in1({ S840, S826 }),
  .out1({ S843 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_172_ (
  .in1({ S839, S825 }),
  .out1({ S844 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_85_ (
  .in1({ S843, S841 }),
  .out1({ S845 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_173_ (
  .in1({ S844, S842 }),
  .out1({ S846 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_86_ (
  .in1({ S846, S816 }),
  .out1({ S847 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_174_ (
  .in1({ S845, S815 }),
  .out1({ S848 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_87_ (
  .in1({ S845, S815 }),
  .out1({ S849 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_175_ (
  .in1({ S846, S816 }),
  .out1({ S850 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_88_ (
  .in1({ S849, S847 }),
  .out1({ S851 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_176_ (
  .in1({ S850, S848 }),
  .out1({ S852 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_89_ (
  .in1({ S851, S813 }),
  .out1({ S853 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_177_ (
  .in1({ S852, S814 }),
  .out1({ S854 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_90_ (
  .in1({ S852, S814 }),
  .out1({ S855 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_178_ (
  .in1({ S851, S813 }),
  .out1({ S856 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_91_ (
  .in1({ S855, S853 }),
  .out1({ S857 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_179_ (
  .in1({ S856, S854 }),
  .out1({ S858 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_92_ (
  .in1({ S858, S803 }),
  .out1({ S859 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_180_ (
  .in1({ S857, S804 }),
  .out1({ S860 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_93_ (
  .in1({ S857, S804 }),
  .out1({ S861 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_181_ (
  .in1({ S858, S803 }),
  .out1({ S862 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_94_ (
  .in1({ S861, S859 }),
  .out1({ S863 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_182_ (
  .in1({ S862, S860 }),
  .out1({ S864 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_95_ (
  .in1({ S863, S736 }),
  .out1({ S865 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_183_ (
  .in1({ S864, S737 }),
  .out1({ S866 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_96_ (
  .in1({ S864, S737 }),
  .out1({ S867 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_184_ (
  .in1({ S863, S736 }),
  .out1({ S868 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_97_ (
  .in1({ S867, S865 }),
  .out1({ S869 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_185_ (
  .in1({ S868, S866 }),
  .out1({ S870 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_98_ (
  .in1({ S870, S800 }),
  .out1({ S871 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_186_ (
  .in1({ S869, S799 }),
  .out1({ S872 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_99_ (
  .in1({ S869, S799 }),
  .out1({ S873 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_187_ (
  .in1({ S870, S800 }),
  .out1({ S874 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_100_ (
  .in1({ S873, S871 }),
  .out1({ S875 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_188_ (
  .in1({ S874, S872 }),
  .out1({ S876 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_101_ (
  .in1({ S875, S774 }),
  .out1({ S877 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_102_ (
  .in1({ S876, S775 }),
  .out1({ S878 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_189_ (
  .in1({ S875, S774 }),
  .out1({ S879 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_190_ (
  .in1({ S879, S1393 }),
  .out1({ S880 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_103_ (
  .in1({ S880, S877 }),
  .out1({ S881 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_104_ (
  .in1({ S881, S798 }),
  .out1({ S882 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_59_ (
  .in1({ S882 }),
  .out1({ DP_ARU1_out_5 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_191_ (
  .in1({ S796, S792 }),
  .out1({ S883 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_60_ (
  .in1({ S883 }),
  .out1({ S884 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_105_ (
  .in1({ S1262, S1251 }),
  .out1({ S885 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_192_ (
  .in1({ DP_AC_dout_6, DP_ARU1_in1_6 }),
  .out1({ S886 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_106_ (
  .in1({ DP_AC_dout_6, DP_ARU1_in1_6 }),
  .out1({ S887 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_107_ (
  .in1({ S887, S885 }),
  .out1({ S888 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_61_ (
  .in1({ S888 }),
  .out1({ S889 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_108_ (
  .in1({ S888, S883 }),
  .out1({ S890 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_109_ (
  .in1({ S889, S884 }),
  .out1({ S891 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_110_ (
  .in1({ S891, S890 }),
  .out1({ S892 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_193_ (
  .in1({ S892, S54 }),
  .out1({ S893 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_111_ (
  .in1({ S878, S871 }),
  .out1({ S894 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_194_ (
  .in1({ S879, S872 }),
  .out1({ S895 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_112_ (
  .in1({ S867, S859 }),
  .out1({ S896 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_62_ (
  .in1({ S896 }),
  .out1({ S897 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_113_ (
  .in1({ S855, S847 }),
  .out1({ S898 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_195_ (
  .in1({ S856, S848 }),
  .out1({ S899 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_196_ (
  .in1({ DP_AC_dout_6, DP_ARU1_in1_0 }),
  .out1({ S900 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_63_ (
  .in1({ S900 }),
  .out1({ S901 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_114_ (
  .in1({ S900, S824 }),
  .out1({ S902 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_197_ (
  .in1({ S901, S823 }),
  .out1({ S903 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_115_ (
  .in1({ S901, S823 }),
  .out1({ S904 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_198_ (
  .in1({ S900, S824 }),
  .out1({ S905 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_116_ (
  .in1({ S904, S902 }),
  .out1({ S906 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_199_ (
  .in1({ S905, S903 }),
  .out1({ S907 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_117_ (
  .in1({ S906, S689 }),
  .out1({ S908 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_200_ (
  .in1({ S907, S690 }),
  .out1({ S909 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_118_ (
  .in1({ S907, S690 }),
  .out1({ S910 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_201_ (
  .in1({ S906, S689 }),
  .out1({ S911 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_119_ (
  .in1({ S910, S908 }),
  .out1({ S912 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_202_ (
  .in1({ S911, S909 }),
  .out1({ S913 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_120_ (
  .in1({ S843, S835 }),
  .out1({ S914 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_203_ (
  .in1({ S844, S836 }),
  .out1({ S915 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_204_ (
  .in1({ DP_ARU1_in1_5, DP_AC_dout_1 }),
  .out1({ S916 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_205_ (
  .in1({ DP_AC_dout_4, DP_ARU1_in1_2 }),
  .out1({ S917 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_206_ (
  .in1({ DP_ARU1_in1_6, DP_AC_dout_0 }),
  .out1({ S918 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_207_ (
  .in1({ DP_ARU1_in1_6, DP_AC_dout_4 }),
  .out1({ S919 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_64_ (
  .in1({ S919 }),
  .out1({ S920 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_121_ (
  .in1({ S919, S671 }),
  .out1({ S921 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_65_ (
  .in1({ S921 }),
  .out1({ S922 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_208_ (
  .in1({ S918, S917 }),
  .out1({ S923 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_209_ (
  .in1({ S923, S922 }),
  .out1({ S924 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_210_ (
  .in1({ S924, S916 }),
  .out1({ S925 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_66_ (
  .in1({ S925 }),
  .out1({ S926 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_122_ (
  .in1({ S924, S916 }),
  .out1({ S927 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_67_ (
  .in1({ S927 }),
  .out1({ S928 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_123_ (
  .in1({ S927, S926 }),
  .out1({ S929 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_211_ (
  .in1({ S928, S925 }),
  .out1({ S930 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_212_ (
  .in1({ DP_AC_dout_5, DP_ARU1_in1_1 }),
  .out1({ S931 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_213_ (
  .in1({ DP_ARU1_in1_4, DP_AC_dout_2 }),
  .out1({ S932 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_214_ (
  .in1({ S932, S931 }),
  .out1({ S933 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_68_ (
  .in1({ S933 }),
  .out1({ S934 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_215_ (
  .in1({ DP_AC_dout_5, DP_ARU1_in1_4 }),
  .out1({ S935 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_69_ (
  .in1({ S935 }),
  .out1({ S936 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_124_ (
  .in1({ S935, S696 }),
  .out1({ S937 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_216_ (
  .in1({ S936, S697 }),
  .out1({ S938 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_125_ (
  .in1({ S937, S934 }),
  .out1({ S939 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_217_ (
  .in1({ S938, S933 }),
  .out1({ S940 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_126_ (
  .in1({ S940, S832 }),
  .out1({ S941 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_218_ (
  .in1({ S939, S831 }),
  .out1({ S942 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_127_ (
  .in1({ S939, S831 }),
  .out1({ S943 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_219_ (
  .in1({ S940, S832 }),
  .out1({ S944 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_128_ (
  .in1({ S943, S941 }),
  .out1({ S945 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_220_ (
  .in1({ S944, S942 }),
  .out1({ S946 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_129_ (
  .in1({ S945, S929 }),
  .out1({ S947 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_221_ (
  .in1({ S946, S930 }),
  .out1({ S948 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_130_ (
  .in1({ S946, S930 }),
  .out1({ S949 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_222_ (
  .in1({ S945, S929 }),
  .out1({ S950 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_131_ (
  .in1({ S949, S947 }),
  .out1({ S951 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_223_ (
  .in1({ S950, S948 }),
  .out1({ S952 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_132_ (
  .in1({ S952, S914 }),
  .out1({ S953 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_224_ (
  .in1({ S951, S915 }),
  .out1({ S954 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_133_ (
  .in1({ S951, S915 }),
  .out1({ S955 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_225_ (
  .in1({ S952, S914 }),
  .out1({ S956 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_134_ (
  .in1({ S955, S953 }),
  .out1({ S957 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_226_ (
  .in1({ S956, S954 }),
  .out1({ S958 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_135_ (
  .in1({ S957, S912 }),
  .out1({ S959 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_227_ (
  .in1({ S958, S913 }),
  .out1({ S960 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_136_ (
  .in1({ S958, S913 }),
  .out1({ S961 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_228_ (
  .in1({ S957, S912 }),
  .out1({ S962 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_137_ (
  .in1({ S961, S959 }),
  .out1({ S963 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_229_ (
  .in1({ S962, S960 }),
  .out1({ S964 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_138_ (
  .in1({ S964, S898 }),
  .out1({ S965 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_230_ (
  .in1({ S963, S899 }),
  .out1({ S966 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_139_ (
  .in1({ S963, S899 }),
  .out1({ S967 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_231_ (
  .in1({ S964, S898 }),
  .out1({ S968 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_140_ (
  .in1({ S967, S965 }),
  .out1({ S969 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_232_ (
  .in1({ S968, S966 }),
  .out1({ S970 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_141_ (
  .in1({ S969, S809 }),
  .out1({ S971 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_233_ (
  .in1({ S970, S810 }),
  .out1({ S972 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_142_ (
  .in1({ S970, S810 }),
  .out1({ S973 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_234_ (
  .in1({ S969, S809 }),
  .out1({ S974 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_143_ (
  .in1({ S973, S971 }),
  .out1({ S975 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_235_ (
  .in1({ S974, S972 }),
  .out1({ S976 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_236_ (
  .in1({ S976, S896 }),
  .out1({ S977 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_237_ (
  .in1({ S975, S897 }),
  .out1({ S978 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_70_ (
  .in1({ S978 }),
  .out1({ S979 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_238_ (
  .in1({ S978, S977 }),
  .out1({ S980 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_71_ (
  .in1({ S980 }),
  .out1({ S981 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_144_ (
  .in1({ S981, S895 }),
  .out1({ S982 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_72_ (
  .in1({ S982 }),
  .out1({ S983 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_145_ (
  .in1({ S980, S894 }),
  .out1({ S984 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_239_ (
  .in1({ S981, S895 }),
  .out1({ S985 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_146_ (
  .in1({ S984, S1404 }),
  .out1({ S986 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_240_ (
  .in1({ S986, S983 }),
  .out1({ S987 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_241_ (
  .in1({ S987, S893 }),
  .out1({ DP_ARU1_out_6 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_147_ (
  .in1({ S891, S885 }),
  .out1({ S988 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_148_ (
  .in1({ S1284, S1273 }),
  .out1({ S989 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_242_ (
  .in1({ DP_AC_dout_7, DP_ARU1_in1_7 }),
  .out1({ S990 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_149_ (
  .in1({ DP_AC_dout_7, DP_ARU1_in1_7 }),
  .out1({ S991 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_73_ (
  .in1({ S991 }),
  .out1({ S992 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_243_ (
  .in1({ S992, S990 }),
  .out1({ S993 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_150_ (
  .in1({ S993, S988 }),
  .out1({ S994 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_244_ (
  .in1({ S993, S988 }),
  .out1({ S995 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_245_ (
  .in1({ S995, S55 }),
  .out1({ S996 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_151_ (
  .in1({ S996, S994 }),
  .out1({ S997 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_152_ (
  .in1({ S984, S979 }),
  .out1({ S998 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_246_ (
  .in1({ S985, S978 }),
  .out1({ S999 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_153_ (
  .in1({ S973, S965 }),
  .out1({ S1000 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_74_ (
  .in1({ S1000 }),
  .out1({ S1001 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_154_ (
  .in1({ S910, S902 }),
  .out1({ S1002 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_247_ (
  .in1({ S911, S903 }),
  .out1({ S1003 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_155_ (
  .in1({ S961, S953 }),
  .out1({ S1004 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_248_ (
  .in1({ S962, S954 }),
  .out1({ S1005 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_249_ (
  .in1({ DP_AC_dout_7, DP_ARU1_in1_0 }),
  .out1({ S1006 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_75_ (
  .in1({ S1006 }),
  .out1({ S1007 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_156_ (
  .in1({ S927, S921 }),
  .out1({ S1008 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_76_ (
  .in1({ S1008 }),
  .out1({ S1009 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_157_ (
  .in1({ S1008, S1006 }),
  .out1({ S1010 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_250_ (
  .in1({ S1009, S1007 }),
  .out1({ S1011 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_251_ (
  .in1({ S1008, S1006 }),
  .out1({ S1012 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_77_ (
  .in1({ S1012 }),
  .out1({ S1013 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_158_ (
  .in1({ S1013, S1010 }),
  .out1({ S1014 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_252_ (
  .in1({ S1012, S1011 }),
  .out1({ S1015 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_159_ (
  .in1({ S1014, S734 }),
  .out1({ S1016 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_253_ (
  .in1({ S1015, S735 }),
  .out1({ S1017 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_160_ (
  .in1({ S1015, S735 }),
  .out1({ S1018 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_254_ (
  .in1({ S1014, S734 }),
  .out1({ S1019 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_161_ (
  .in1({ S1018, S1016 }),
  .out1({ S1020 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_255_ (
  .in1({ S1019, S1017 }),
  .out1({ S1021 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_162_ (
  .in1({ S949, S941 }),
  .out1({ S1022 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_256_ (
  .in1({ S950, S942 }),
  .out1({ S1023 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_257_ (
  .in1({ DP_ARU1_in1_5, DP_AC_dout_2 }),
  .out1({ S1024 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_258_ (
  .in1({ DP_AC_dout_5, DP_ARU1_in1_2 }),
  .out1({ S1025 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_259_ (
  .in1({ DP_ARU1_in1_6, DP_AC_dout_1 }),
  .out1({ S1026 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_260_ (
  .in1({ DP_ARU1_in1_6, DP_AC_dout_5 }),
  .out1({ S1027 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_163_ (
  .in1({ S1027, S673 }),
  .out1({ S1028 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_78_ (
  .in1({ S1028 }),
  .out1({ S1029 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_261_ (
  .in1({ S1026, S1025 }),
  .out1({ S1030 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_262_ (
  .in1({ S1030, S1029 }),
  .out1({ S1031 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_263_ (
  .in1({ S1031, S1024 }),
  .out1({ S1032 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_79_ (
  .in1({ S1032 }),
  .out1({ S1033 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_164_ (
  .in1({ S1031, S1024 }),
  .out1({ S1034 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_80_ (
  .in1({ S1034 }),
  .out1({ S1035 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_165_ (
  .in1({ S1034, S1033 }),
  .out1({ S1036 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_264_ (
  .in1({ S1035, S1032 }),
  .out1({ S1037 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_265_ (
  .in1({ DP_AC_dout_6, DP_ARU1_in1_1 }),
  .out1({ S1038 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_81_ (
  .in1({ S1038 }),
  .out1({ S1039 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_266_ (
  .in1({ DP_ARU1_in1_7, DP_AC_dout_0 }),
  .out1({ S1040 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_267_ (
  .in1({ DP_ARU1_in1_7, DP_AC_dout_3 }),
  .out1({ S1041 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_166_ (
  .in1({ S1041, S743 }),
  .out1({ S1042 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_82_ (
  .in1({ S1042 }),
  .out1({ S1043 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_268_ (
  .in1({ S1040, S746 }),
  .out1({ S1044 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_83_ (
  .in1({ S1044 }),
  .out1({ S1045 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_167_ (
  .in1({ S1045, S1042 }),
  .out1({ S1046 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_269_ (
  .in1({ S1044, S1043 }),
  .out1({ S1047 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_168_ (
  .in1({ S1046, S1039 }),
  .out1({ S1048 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_270_ (
  .in1({ S1047, S1038 }),
  .out1({ S1049 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_169_ (
  .in1({ S1047, S1038 }),
  .out1({ S1050 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_84_ (
  .in1({ S1050 }),
  .out1({ S1051 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_170_ (
  .in1({ S1050, S1048 }),
  .out1({ S1052 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_271_ (
  .in1({ S1051, S1049 }),
  .out1({ S1053 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_171_ (
  .in1({ S1053, S938 }),
  .out1({ S1054 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_272_ (
  .in1({ S1052, S937 }),
  .out1({ S1055 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_172_ (
  .in1({ S1052, S937 }),
  .out1({ S1056 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_273_ (
  .in1({ S1053, S938 }),
  .out1({ S1057 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_173_ (
  .in1({ S1056, S1054 }),
  .out1({ S1058 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_274_ (
  .in1({ S1057, S1055 }),
  .out1({ S1059 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_174_ (
  .in1({ S1058, S1036 }),
  .out1({ S1060 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_275_ (
  .in1({ S1059, S1037 }),
  .out1({ S1061 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_175_ (
  .in1({ S1059, S1037 }),
  .out1({ S1062 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_276_ (
  .in1({ S1058, S1036 }),
  .out1({ S1063 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_176_ (
  .in1({ S1062, S1060 }),
  .out1({ S1064 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_277_ (
  .in1({ S1063, S1061 }),
  .out1({ S1065 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_177_ (
  .in1({ S1065, S1022 }),
  .out1({ S1066 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_278_ (
  .in1({ S1064, S1023 }),
  .out1({ S1067 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_178_ (
  .in1({ S1064, S1023 }),
  .out1({ S1068 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_279_ (
  .in1({ S1065, S1022 }),
  .out1({ S1069 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_179_ (
  .in1({ S1068, S1066 }),
  .out1({ S1070 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_280_ (
  .in1({ S1069, S1067 }),
  .out1({ S1071 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_180_ (
  .in1({ S1070, S1020 }),
  .out1({ S1072 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_281_ (
  .in1({ S1071, S1021 }),
  .out1({ S1073 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_181_ (
  .in1({ S1071, S1021 }),
  .out1({ S1074 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_282_ (
  .in1({ S1070, S1020 }),
  .out1({ S1075 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_182_ (
  .in1({ S1074, S1072 }),
  .out1({ S1076 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_283_ (
  .in1({ S1075, S1073 }),
  .out1({ S1077 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_183_ (
  .in1({ S1077, S1004 }),
  .out1({ S1078 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_284_ (
  .in1({ S1076, S1005 }),
  .out1({ S1079 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_184_ (
  .in1({ S1076, S1005 }),
  .out1({ S1080 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_285_ (
  .in1({ S1077, S1004 }),
  .out1({ S1081 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_185_ (
  .in1({ S1080, S1078 }),
  .out1({ S1082 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_286_ (
  .in1({ S1081, S1079 }),
  .out1({ S1083 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_186_ (
  .in1({ S1082, S1003 }),
  .out1({ S1084 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_287_ (
  .in1({ S1083, S1002 }),
  .out1({ S1085 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_187_ (
  .in1({ S1083, S1002 }),
  .out1({ S1086 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_288_ (
  .in1({ S1082, S1003 }),
  .out1({ S1087 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_188_ (
  .in1({ S1086, S1084 }),
  .out1({ S1088 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_289_ (
  .in1({ S1087, S1085 }),
  .out1({ S1089 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_290_ (
  .in1({ S1088, S1001 }),
  .out1({ S1090 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_85_ (
  .in1({ S1090 }),
  .out1({ S1091 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_291_ (
  .in1({ S1089, S1000 }),
  .out1({ S1092 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_292_ (
  .in1({ S1092, S1090 }),
  .out1({ S1093 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_86_ (
  .in1({ S1093 }),
  .out1({ S1094 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_293_ (
  .in1({ S1093, S998 }),
  .out1({ S1095 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_189_ (
  .in1({ S1093, S998 }),
  .out1({ S1096 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_294_ (
  .in1({ S1094, S999 }),
  .out1({ S1097 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_190_ (
  .in1({ S1096, S1404 }),
  .out1({ S1098 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_295_ (
  .in1({ S1098, S1095 }),
  .out1({ S1100 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_87_ (
  .in1({ S1100 }),
  .out1({ S1101 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_191_ (
  .in1({ S1101, S997 }),
  .out1({ S1102 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_88_ (
  .in1({ S1102 }),
  .out1({ DP_ARU1_out_7 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_192_ (
  .in1({ S1096, S1091 }),
  .out1({ S1103 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_296_ (
  .in1({ S1097, S1090 }),
  .out1({ S1104 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_193_ (
  .in1({ S1086, S1078 }),
  .out1({ S1105 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_89_ (
  .in1({ S1105 }),
  .out1({ S1106 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_194_ (
  .in1({ S1018, S1010 }),
  .out1({ S1107 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_90_ (
  .in1({ S1107 }),
  .out1({ S1108 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_195_ (
  .in1({ S1074, S1066 }),
  .out1({ S1110 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_297_ (
  .in1({ S1075, S1067 }),
  .out1({ S1111 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_196_ (
  .in1({ S1034, S1028 }),
  .out1({ S1112 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_91_ (
  .in1({ S1112 }),
  .out1({ S1113 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_197_ (
  .in1({ S1112, S807 }),
  .out1({ S1114 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_298_ (
  .in1({ S1113, S808 }),
  .out1({ S1115 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_299_ (
  .in1({ S1112, S807 }),
  .out1({ S1116 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_92_ (
  .in1({ S1116 }),
  .out1({ S1117 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_198_ (
  .in1({ S1117, S1114 }),
  .out1({ S1118 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_300_ (
  .in1({ S1116, S1115 }),
  .out1({ S1119 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_199_ (
  .in1({ S1062, S1054 }),
  .out1({ S1121 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_301_ (
  .in1({ S1063, S1055 }),
  .out1({ S1122 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_302_ (
  .in1({ DP_AC_dout_6, DP_ARU1_in1_2 }),
  .out1({ S1123 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_303_ (
  .in1({ DP_ARU1_in1_6, DP_AC_dout_2 }),
  .out1({ S1124 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_200_ (
  .in1({ S886, S659 }),
  .out1({ S1125 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_304_ (
  .in1({ S885, S650 }),
  .out1({ S1126 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_305_ (
  .in1({ S1124, S1123 }),
  .out1({ S1127 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_306_ (
  .in1({ S1127, S1126 }),
  .out1({ S1128 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_307_ (
  .in1({ S1128, S821 }),
  .out1({ S1129 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_93_ (
  .in1({ S1129 }),
  .out1({ S1130 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_201_ (
  .in1({ S1128, S821 }),
  .out1({ S1132 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_94_ (
  .in1({ S1132 }),
  .out1({ S1133 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_202_ (
  .in1({ S1132, S1130 }),
  .out1({ S1134 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_308_ (
  .in1({ S1133, S1129 }),
  .out1({ S1135 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_203_ (
  .in1({ S1050, S1042 }),
  .out1({ S1136 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_95_ (
  .in1({ S1136 }),
  .out1({ S1137 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_309_ (
  .in1({ DP_AC_dout_7, DP_ARU1_in1_1 }),
  .out1({ S1138 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_310_ (
  .in1({ DP_ARU1_in1_7, DP_AC_dout_1 }),
  .out1({ S1139 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_311_ (
  .in1({ DP_ARU1_in1_7, DP_AC_dout_4 }),
  .out1({ S1140 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_204_ (
  .in1({ S1140, S828 }),
  .out1({ S1141 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_96_ (
  .in1({ S1141 }),
  .out1({ S1143 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_312_ (
  .in1({ S1139, S779 }),
  .out1({ S1144 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_313_ (
  .in1({ S1144, S1143 }),
  .out1({ S1145 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_314_ (
  .in1({ S1145, S1138 }),
  .out1({ S1146 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_205_ (
  .in1({ S1145, S1138 }),
  .out1({ S1147 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_97_ (
  .in1({ S1147 }),
  .out1({ S1148 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_315_ (
  .in1({ S1148, S1146 }),
  .out1({ S1149 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_98_ (
  .in1({ S1149 }),
  .out1({ S1150 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_206_ (
  .in1({ S1149, S1136 }),
  .out1({ S1151 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_316_ (
  .in1({ S1150, S1137 }),
  .out1({ S1152 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_317_ (
  .in1({ S1149, S1136 }),
  .out1({ S1154 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_99_ (
  .in1({ S1154 }),
  .out1({ S1155 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_207_ (
  .in1({ S1155, S1151 }),
  .out1({ S1156 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_318_ (
  .in1({ S1154, S1152 }),
  .out1({ S1157 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_208_ (
  .in1({ S1156, S1134 }),
  .out1({ S1158 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_319_ (
  .in1({ S1157, S1135 }),
  .out1({ S1159 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_209_ (
  .in1({ S1157, S1135 }),
  .out1({ S1160 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_320_ (
  .in1({ S1156, S1134 }),
  .out1({ S1161 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_210_ (
  .in1({ S1160, S1158 }),
  .out1({ S1162 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_321_ (
  .in1({ S1161, S1159 }),
  .out1({ S1163 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_211_ (
  .in1({ S1163, S1121 }),
  .out1({ S1165 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_322_ (
  .in1({ S1162, S1122 }),
  .out1({ S1166 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_212_ (
  .in1({ S1162, S1122 }),
  .out1({ S1167 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_323_ (
  .in1({ S1163, S1121 }),
  .out1({ S1168 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_213_ (
  .in1({ S1167, S1165 }),
  .out1({ S1169 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_324_ (
  .in1({ S1168, S1166 }),
  .out1({ S1170 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_214_ (
  .in1({ S1169, S1118 }),
  .out1({ S1171 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_325_ (
  .in1({ S1170, S1119 }),
  .out1({ S1172 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_215_ (
  .in1({ S1170, S1119 }),
  .out1({ S1173 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_326_ (
  .in1({ S1169, S1118 }),
  .out1({ S1174 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_216_ (
  .in1({ S1173, S1171 }),
  .out1({ S1176 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_327_ (
  .in1({ S1174, S1172 }),
  .out1({ S1177 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_217_ (
  .in1({ S1177, S1110 }),
  .out1({ S1178 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_328_ (
  .in1({ S1176, S1111 }),
  .out1({ S1179 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_218_ (
  .in1({ S1176, S1111 }),
  .out1({ S1180 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_329_ (
  .in1({ S1177, S1110 }),
  .out1({ S1181 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_219_ (
  .in1({ S1180, S1178 }),
  .out1({ S1182 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_330_ (
  .in1({ S1181, S1179 }),
  .out1({ S1183 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_331_ (
  .in1({ S1183, S1107 }),
  .out1({ S1184 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_220_ (
  .in1({ S1183, S1107 }),
  .out1({ S1185 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_332_ (
  .in1({ S1182, S1108 }),
  .out1({ S1187 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_333_ (
  .in1({ S1187, S1184 }),
  .out1({ S1188 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_100_ (
  .in1({ S1188 }),
  .out1({ S1189 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_334_ (
  .in1({ S1188, S1105 }),
  .out1({ S1190 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_335_ (
  .in1({ S1189, S1106 }),
  .out1({ S1191 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_101_ (
  .in1({ S1191 }),
  .out1({ S1192 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_336_ (
  .in1({ S1191, S1190 }),
  .out1({ S1193 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_102_ (
  .in1({ S1193 }),
  .out1({ S1194 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_221_ (
  .in1({ S1193, S1103 }),
  .out1({ S1195 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_337_ (
  .in1({ S1194, S1104 }),
  .out1({ S1196 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_222_ (
  .in1({ S1194, S1104 }),
  .out1({ S1198 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_223_ (
  .in1({ S1198, S1404 }),
  .out1({ S1199 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_338_ (
  .in1({ S1199, S1196 }),
  .out1({ S1200 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_339_ (
  .in1({ DP_ARU1_in1_8, DP_AC_dout_8 }),
  .out1({ S1201 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_103_ (
  .in1({ S1201 }),
  .out1({ S1202 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_224_ (
  .in1({ DP_ARU1_in1_8, DP_AC_dout_8 }),
  .out1({ S1203 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_225_ (
  .in1({ S1203, S1202 }),
  .out1({ S1204 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_226_ (
  .in1({ S991, S988 }),
  .out1({ S1205 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_104_ (
  .in1({ S1205 }),
  .out1({ S1206 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_340_ (
  .in1({ S1206, S990 }),
  .out1({ S1207 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_227_ (
  .in1({ S1207, S1204 }),
  .out1({ S1209 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_341_ (
  .in1({ S1207, S1204 }),
  .out1({ S1210 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_105_ (
  .in1({ S1210 }),
  .out1({ S1211 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_228_ (
  .in1({ S1211, S1209 }),
  .out1({ S1212 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_342_ (
  .in1({ S1212, S56 }),
  .out1({ S1213 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_343_ (
  .in1({ S1213, S1200 }),
  .out1({ DP_ARU1_out_8 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_344_ (
  .in1({ S1210, S1201 }),
  .out1({ S1214 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_345_ (
  .in1({ DP_ARU1_in1_9, DP_AC_dout_9 }),
  .out1({ S1215 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_106_ (
  .in1({ S1215 }),
  .out1({ S1216 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_229_ (
  .in1({ DP_ARU1_in1_9, DP_AC_dout_9 }),
  .out1({ S1217 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_230_ (
  .in1({ S1217, S1216 }),
  .out1({ S1219 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_231_ (
  .in1({ S1219, S1214 }),
  .out1({ S1220 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_346_ (
  .in1({ S1219, S1214 }),
  .out1({ S1221 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_347_ (
  .in1({ S1221, S57 }),
  .out1({ S1222 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_232_ (
  .in1({ S1222, S1220 }),
  .out1({ S1223 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_233_ (
  .in1({ S1195, S1192 }),
  .out1({ S1224 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_348_ (
  .in1({ S1196, S1191 }),
  .out1({ S1225 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_234_ (
  .in1({ S1185, S1178 }),
  .out1({ S1226 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_107_ (
  .in1({ S1226 }),
  .out1({ S1227 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_235_ (
  .in1({ S1173, S1165 }),
  .out1({ S1228 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_349_ (
  .in1({ DP_AC_dout_6, DP_ARU1_in1_3 }),
  .out1({ S1230 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_108_ (
  .in1({ S1230 }),
  .out1({ S1231 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_236_ (
  .in1({ S1132, S1125 }),
  .out1({ S1232 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_109_ (
  .in1({ S1232 }),
  .out1({ S1233 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_237_ (
  .in1({ S1232, S1230 }),
  .out1({ S1234 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_350_ (
  .in1({ S1233, S1231 }),
  .out1({ S1235 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_351_ (
  .in1({ S1232, S1230 }),
  .out1({ S1236 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_110_ (
  .in1({ S1236 }),
  .out1({ S1237 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_238_ (
  .in1({ S1237, S1234 }),
  .out1({ S1238 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_352_ (
  .in1({ S1236, S1235 }),
  .out1({ S1239 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_239_ (
  .in1({ S1160, S1151 }),
  .out1({ S1241 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_353_ (
  .in1({ S1161, S1152 }),
  .out1({ S1242 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_354_ (
  .in1({ DP_ARU1_in1_5, DP_AC_dout_4 }),
  .out1({ S1243 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_355_ (
  .in1({ DP_AC_dout_7, DP_ARU1_in1_2 }),
  .out1({ S1244 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_356_ (
  .in1({ DP_ARU1_in1_6, DP_AC_dout_3 }),
  .out1({ S1245 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_357_ (
  .in1({ DP_AC_dout_7, DP_ARU1_in1_6 }),
  .out1({ S1246 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_240_ (
  .in1({ S1246, S818 }),
  .out1({ S1247 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_111_ (
  .in1({ S1247 }),
  .out1({ S1248 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_358_ (
  .in1({ S1245, S1244 }),
  .out1({ S1249 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_359_ (
  .in1({ S1249, S1248 }),
  .out1({ S1250 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_360_ (
  .in1({ S1250, S1243 }),
  .out1({ S1252 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_112_ (
  .in1({ S1252 }),
  .out1({ S1253 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_241_ (
  .in1({ S1250, S1243 }),
  .out1({ S1254 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_113_ (
  .in1({ S1254 }),
  .out1({ S1255 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_242_ (
  .in1({ S1254, S1253 }),
  .out1({ S1256 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_361_ (
  .in1({ S1255, S1252 }),
  .out1({ S1257 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_243_ (
  .in1({ S1147, S1141 }),
  .out1({ S1258 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_114_ (
  .in1({ S1258 }),
  .out1({ S1259 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_244_ (
  .in1({ S1273, S1175 }),
  .out1({ S1260 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_362_ (
  .in1({ DP_ARU1_in1_7, DP_AC_dout_2 }),
  .out1({ S1261 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_363_ (
  .in1({ DP_ARU1_in1_7, DP_AC_dout_5 }),
  .out1({ S1263 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_245_ (
  .in1({ S1263, S932 }),
  .out1({ S1264 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_364_ (
  .in1({ S1260, S936 }),
  .out1({ S1265 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_365_ (
  .in1({ S1261, S935 }),
  .out1({ S1266 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_366_ (
  .in1({ S1266, S1265 }),
  .out1({ S1267 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_115_ (
  .in1({ S1267 }),
  .out1({ S1268 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_246_ (
  .in1({ S1267, S1258 }),
  .out1({ S1269 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_367_ (
  .in1({ S1268, S1259 }),
  .out1({ S1270 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_368_ (
  .in1({ S1267, S1258 }),
  .out1({ S1271 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_116_ (
  .in1({ S1271 }),
  .out1({ S1272 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_247_ (
  .in1({ S1272, S1269 }),
  .out1({ S1274 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_369_ (
  .in1({ S1271, S1270 }),
  .out1({ S1275 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_248_ (
  .in1({ S1274, S1256 }),
  .out1({ S1276 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_370_ (
  .in1({ S1275, S1257 }),
  .out1({ S1277 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_249_ (
  .in1({ S1275, S1257 }),
  .out1({ S1278 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_371_ (
  .in1({ S1274, S1256 }),
  .out1({ S1279 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_250_ (
  .in1({ S1278, S1276 }),
  .out1({ S1280 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_372_ (
  .in1({ S1279, S1277 }),
  .out1({ S1281 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_251_ (
  .in1({ S1281, S1241 }),
  .out1({ S1282 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_373_ (
  .in1({ S1280, S1242 }),
  .out1({ S1283 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_252_ (
  .in1({ S1280, S1242 }),
  .out1({ S1285 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_374_ (
  .in1({ S1281, S1241 }),
  .out1({ S1286 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_253_ (
  .in1({ S1285, S1282 }),
  .out1({ S1287 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_375_ (
  .in1({ S1286, S1283 }),
  .out1({ S1288 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_376_ (
  .in1({ S1288, S1239 }),
  .out1({ S1289 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_254_ (
  .in1({ S1288, S1239 }),
  .out1({ S1290 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_377_ (
  .in1({ S1287, S1238 }),
  .out1({ S1291 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_378_ (
  .in1({ S1291, S1289 }),
  .out1({ S1292 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_255_ (
  .in1({ S1292, S1228 }),
  .out1({ S1293 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_117_ (
  .in1({ S1293 }),
  .out1({ S1294 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_379_ (
  .in1({ S1292, S1228 }),
  .out1({ S1296 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_380_ (
  .in1({ S1296, S1294 }),
  .out1({ S1297 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_118_ (
  .in1({ S1297 }),
  .out1({ S1298 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_381_ (
  .in1({ S1297, S1115 }),
  .out1({ S1299 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_256_ (
  .in1({ S1297, S1115 }),
  .out1({ S1300 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_382_ (
  .in1({ S1298, S1114 }),
  .out1({ S1301 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_383_ (
  .in1({ S1301, S1299 }),
  .out1({ S1302 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_119_ (
  .in1({ S1302 }),
  .out1({ S1303 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_384_ (
  .in1({ S1303, S1227 }),
  .out1({ S1304 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_120_ (
  .in1({ S1304 }),
  .out1({ S1305 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_385_ (
  .in1({ S1302, S1226 }),
  .out1({ S1307 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_386_ (
  .in1({ S1307, S1304 }),
  .out1({ S1308 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_121_ (
  .in1({ S1308 }),
  .out1({ S1309 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_257_ (
  .in1({ S1308, S1224 }),
  .out1({ S1310 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_387_ (
  .in1({ S1309, S1225 }),
  .out1({ S1311 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_388_ (
  .in1({ S1308, S1224 }),
  .out1({ S1312 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_389_ (
  .in1({ S1312, S1393 }),
  .out1({ S1313 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_258_ (
  .in1({ S1313, S1310 }),
  .out1({ S1314 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_259_ (
  .in1({ S1314, S1223 }),
  .out1({ S1315 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_122_ (
  .in1({ S1315 }),
  .out1({ DP_ARU1_out_9 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_390_ (
  .in1({ DP_ARU1_in1_10, DP_AC_dout_10 }),
  .out1({ S1317 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_123_ (
  .in1({ S1317 }),
  .out1({ S1318 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_260_ (
  .in1({ DP_ARU1_in1_10, DP_AC_dout_10 }),
  .out1({ S1319 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_261_ (
  .in1({ S1319, S1318 }),
  .out1({ S1320 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_262_ (
  .in1({ S1216, S1214 }),
  .out1({ S1321 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_263_ (
  .in1({ S1321, S1217 }),
  .out1({ S1322 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_264_ (
  .in1({ S1322, S1320 }),
  .out1({ S1323 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_391_ (
  .in1({ S1322, S1320 }),
  .out1({ S1324 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_265_ (
  .in1({ S1323, S1131 }),
  .out1({ S1325 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_392_ (
  .in1({ S1325, S1324 }),
  .out1({ S1326 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_266_ (
  .in1({ S1310, S1305 }),
  .out1({ S1328 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_393_ (
  .in1({ S1311, S1304 }),
  .out1({ S1329 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_267_ (
  .in1({ S1300, S1293 }),
  .out1({ S1330 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_124_ (
  .in1({ S1330 }),
  .out1({ S1331 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_268_ (
  .in1({ S1290, S1282 }),
  .out1({ S1332 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_394_ (
  .in1({ DP_AC_dout_7, DP_ARU1_in1_3 }),
  .out1({ S1333 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_125_ (
  .in1({ S1333 }),
  .out1({ S1334 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_269_ (
  .in1({ S1254, S1247 }),
  .out1({ S1335 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_126_ (
  .in1({ S1335 }),
  .out1({ S1336 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_270_ (
  .in1({ S1335, S1333 }),
  .out1({ S1337 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_395_ (
  .in1({ S1336, S1334 }),
  .out1({ S1339 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_396_ (
  .in1({ S1335, S1333 }),
  .out1({ S1340 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_127_ (
  .in1({ S1340 }),
  .out1({ S1341 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_271_ (
  .in1({ S1341, S1337 }),
  .out1({ S1342 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_397_ (
  .in1({ S1340, S1339 }),
  .out1({ S1343 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_272_ (
  .in1({ S1278, S1269 }),
  .out1({ S1344 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_398_ (
  .in1({ S1279, S1270 }),
  .out1({ S1345 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_273_ (
  .in1({ S919, S792 }),
  .out1({ S1346 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_399_ (
  .in1({ S920, S791 }),
  .out1({ S1347 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_400_ (
  .in1({ S919, S792 }),
  .out1({ S1348 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_128_ (
  .in1({ S1348 }),
  .out1({ S1350 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_274_ (
  .in1({ S1350, S1346 }),
  .out1({ S1351 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_401_ (
  .in1({ S1348, S1347 }),
  .out1({ S1352 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_402_ (
  .in1({ DP_AC_dout_6, DP_ARU1_in1_4 }),
  .out1({ S1353 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_403_ (
  .in1({ DP_ARU1_in1_7, DP_AC_dout_6 }),
  .out1({ S1354 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_129_ (
  .in1({ S1354 }),
  .out1({ S1355 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_275_ (
  .in1({ S1354, S746 }),
  .out1({ S1356 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_404_ (
  .in1({ S1355, S747 }),
  .out1({ S1357 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_405_ (
  .in1({ S1353, S1041 }),
  .out1({ S1358 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_130_ (
  .in1({ S1358 }),
  .out1({ S1359 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_276_ (
  .in1({ S1359, S1356 }),
  .out1({ S1361 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_406_ (
  .in1({ S1358, S1357 }),
  .out1({ S1362 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_277_ (
  .in1({ S1362, S1265 }),
  .out1({ S1363 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_407_ (
  .in1({ S1361, S1264 }),
  .out1({ S1364 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_278_ (
  .in1({ S1361, S1264 }),
  .out1({ S1365 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_408_ (
  .in1({ S1362, S1265 }),
  .out1({ S1366 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_279_ (
  .in1({ S1365, S1363 }),
  .out1({ S1367 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_409_ (
  .in1({ S1366, S1364 }),
  .out1({ S1368 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_280_ (
  .in1({ S1367, S1351 }),
  .out1({ S1369 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_410_ (
  .in1({ S1368, S1352 }),
  .out1({ S1370 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_281_ (
  .in1({ S1368, S1352 }),
  .out1({ S1372 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_411_ (
  .in1({ S1367, S1351 }),
  .out1({ S1373 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_282_ (
  .in1({ S1372, S1369 }),
  .out1({ S1374 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_412_ (
  .in1({ S1373, S1370 }),
  .out1({ S1375 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_283_ (
  .in1({ S1375, S1344 }),
  .out1({ S1376 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_413_ (
  .in1({ S1374, S1345 }),
  .out1({ S1377 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_284_ (
  .in1({ S1374, S1345 }),
  .out1({ S1378 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_414_ (
  .in1({ S1375, S1344 }),
  .out1({ S1379 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_285_ (
  .in1({ S1378, S1376 }),
  .out1({ S1380 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_415_ (
  .in1({ S1379, S1377 }),
  .out1({ S1381 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_416_ (
  .in1({ S1381, S1343 }),
  .out1({ S1383 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_286_ (
  .in1({ S1381, S1343 }),
  .out1({ S1384 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_417_ (
  .in1({ S1380, S1342 }),
  .out1({ S1385 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_418_ (
  .in1({ S1385, S1383 }),
  .out1({ S1386 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_287_ (
  .in1({ S1386, S1332 }),
  .out1({ S1387 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_131_ (
  .in1({ S1387 }),
  .out1({ S1388 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_419_ (
  .in1({ S1386, S1332 }),
  .out1({ S1389 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_420_ (
  .in1({ S1389, S1388 }),
  .out1({ S1390 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_132_ (
  .in1({ S1390 }),
  .out1({ S1391 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_421_ (
  .in1({ S1390, S1235 }),
  .out1({ S1392 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_288_ (
  .in1({ S1390, S1235 }),
  .out1({ S1394 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_422_ (
  .in1({ S1391, S1234 }),
  .out1({ S1395 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_423_ (
  .in1({ S1395, S1392 }),
  .out1({ S1396 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_133_ (
  .in1({ S1396 }),
  .out1({ S1397 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_424_ (
  .in1({ S1396, S1330 }),
  .out1({ S1398 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_425_ (
  .in1({ S1397, S1331 }),
  .out1({ S1399 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_134_ (
  .in1({ S1399 }),
  .out1({ S1400 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_426_ (
  .in1({ S1399, S1398 }),
  .out1({ S1401 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_135_ (
  .in1({ S1401 }),
  .out1({ S1402 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_427_ (
  .in1({ S1401, S1328 }),
  .out1({ S1403 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_289_ (
  .in1({ S1401, S1328 }),
  .out1({ S1405 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_428_ (
  .in1({ S1402, S1329 }),
  .out1({ S1406 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_290_ (
  .in1({ S1405, S1404 }),
  .out1({ S1407 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_429_ (
  .in1({ S1407, S1403 }),
  .out1({ S1408 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_430_ (
  .in1({ S1408, S1326 }),
  .out1({ DP_ARU1_out_10 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_431_ (
  .in1({ S1324, S1317 }),
  .out1({ S1409 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_291_ (
  .in1({ S1306, S1295 }),
  .out1({ S1410 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_292_ (
  .in1({ DP_ARU1_in1_11, DP_AC_dout_11 }),
  .out1({ S1411 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_293_ (
  .in1({ S1411, S1410 }),
  .out1({ S1412 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_294_ (
  .in1({ S1412, S1409 }),
  .out1({ S1413 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_432_ (
  .in1({ S1412, S1409 }),
  .out1({ S1415 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_433_ (
  .in1({ S1415, S58 }),
  .out1({ S1416 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_295_ (
  .in1({ S1416, S1413 }),
  .out1({ S1417 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_296_ (
  .in1({ S1405, S1400 }),
  .out1({ S1418 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_434_ (
  .in1({ S1406, S1399 }),
  .out1({ S1419 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_297_ (
  .in1({ S1394, S1387 }),
  .out1({ S1420 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_136_ (
  .in1({ S1420 }),
  .out1({ S1421 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_298_ (
  .in1({ S1384, S1376 }),
  .out1({ S1422 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_299_ (
  .in1({ S1372, S1363 }),
  .out1({ S1423 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_435_ (
  .in1({ S1373, S1364 }),
  .out1({ S1424 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_436_ (
  .in1({ DP_AC_dout_6, DP_ARU1_in1_5 }),
  .out1({ S1426 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_300_ (
  .in1({ S886, S792 }),
  .out1({ S1427 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_437_ (
  .in1({ S885, S791 }),
  .out1({ S1428 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_438_ (
  .in1({ S1426, S1027 }),
  .out1({ S1429 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_137_ (
  .in1({ S1429 }),
  .out1({ S1430 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_301_ (
  .in1({ S1430, S1427 }),
  .out1({ S1431 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_439_ (
  .in1({ S1429, S1428 }),
  .out1({ S1432 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_440_ (
  .in1({ DP_AC_dout_7, DP_ARU1_in1_4 }),
  .out1({ S1433 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_302_ (
  .in1({ S990, S779 }),
  .out1({ S1434 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_441_ (
  .in1({ S989, S778 }),
  .out1({ S1435 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_442_ (
  .in1({ S1433, S1140 }),
  .out1({ S1437 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_138_ (
  .in1({ S1437 }),
  .out1({ S1438 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_303_ (
  .in1({ S1438, S1434 }),
  .out1({ S1439 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_443_ (
  .in1({ S1437, S1435 }),
  .out1({ S1440 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_304_ (
  .in1({ S1440, S1357 }),
  .out1({ S1441 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_444_ (
  .in1({ S1439, S1356 }),
  .out1({ S1442 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_305_ (
  .in1({ S1439, S1356 }),
  .out1({ S1443 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_445_ (
  .in1({ S1440, S1357 }),
  .out1({ S1444 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_306_ (
  .in1({ S1443, S1441 }),
  .out1({ S1445 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_446_ (
  .in1({ S1444, S1442 }),
  .out1({ S1446 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_307_ (
  .in1({ S1445, S1431 }),
  .out1({ S1447 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_447_ (
  .in1({ S1446, S1432 }),
  .out1({ S1448 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_308_ (
  .in1({ S1446, S1432 }),
  .out1({ S1449 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_448_ (
  .in1({ S1445, S1431 }),
  .out1({ S1450 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_309_ (
  .in1({ S1449, S1447 }),
  .out1({ S1451 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_449_ (
  .in1({ S1450, S1448 }),
  .out1({ S1452 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_310_ (
  .in1({ S1452, S1423 }),
  .out1({ S1453 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_450_ (
  .in1({ S1451, S1424 }),
  .out1({ S1454 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_311_ (
  .in1({ S1451, S1424 }),
  .out1({ S1455 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_451_ (
  .in1({ S1452, S1423 }),
  .out1({ S1456 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_312_ (
  .in1({ S1455, S1453 }),
  .out1({ S1458 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_452_ (
  .in1({ S1456, S1454 }),
  .out1({ S1459 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_453_ (
  .in1({ S1459, S1347 }),
  .out1({ S1460 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_313_ (
  .in1({ S1459, S1347 }),
  .out1({ S1461 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_454_ (
  .in1({ S1458, S1346 }),
  .out1({ S1462 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_455_ (
  .in1({ S1462, S1460 }),
  .out1({ S1463 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_314_ (
  .in1({ S1463, S1422 }),
  .out1({ S1464 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_139_ (
  .in1({ S1464 }),
  .out1({ S1465 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_456_ (
  .in1({ S1463, S1422 }),
  .out1({ S1466 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_457_ (
  .in1({ S1466, S1465 }),
  .out1({ S1467 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_140_ (
  .in1({ S1467 }),
  .out1({ S1469 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_458_ (
  .in1({ S1467, S1339 }),
  .out1({ S1470 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_315_ (
  .in1({ S1467, S1339 }),
  .out1({ S1471 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_459_ (
  .in1({ S1469, S1337 }),
  .out1({ S1472 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_460_ (
  .in1({ S1472, S1470 }),
  .out1({ S1473 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_141_ (
  .in1({ S1473 }),
  .out1({ S1474 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_461_ (
  .in1({ S1474, S1421 }),
  .out1({ S1475 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_142_ (
  .in1({ S1475 }),
  .out1({ S1476 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_462_ (
  .in1({ S1473, S1420 }),
  .out1({ S1477 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_463_ (
  .in1({ S1477, S1475 }),
  .out1({ S1478 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_143_ (
  .in1({ S1478 }),
  .out1({ S1480 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_464_ (
  .in1({ S1478, S1418 }),
  .out1({ S1481 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_316_ (
  .in1({ S1478, S1418 }),
  .out1({ S1482 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_465_ (
  .in1({ S1480, S1419 }),
  .out1({ S1483 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_466_ (
  .in1({ S1481, S1393 }),
  .out1({ S1484 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_317_ (
  .in1({ S1484, S1482 }),
  .out1({ S1485 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_318_ (
  .in1({ S1485, S1417 }),
  .out1({ S1486 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_144_ (
  .in1({ S1486 }),
  .out1({ DP_ARU1_out_11 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_319_ (
  .in1({ S1482, S1476 }),
  .out1({ S1487 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_467_ (
  .in1({ S1483, S1475 }),
  .out1({ S1488 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_320_ (
  .in1({ S1471, S1464 }),
  .out1({ S1490 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_145_ (
  .in1({ S1490 }),
  .out1({ S1491 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_321_ (
  .in1({ S1461, S1453 }),
  .out1({ S1492 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_468_ (
  .in1({ S1462, S1454 }),
  .out1({ S1493 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_322_ (
  .in1({ S1449, S1441 }),
  .out1({ S1494 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_469_ (
  .in1({ S1450, S1442 }),
  .out1({ S1495 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_470_ (
  .in1({ DP_AC_dout_7, DP_ARU1_in1_5 }),
  .out1({ S1496 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_146_ (
  .in1({ S1496 }),
  .out1({ S1497 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_471_ (
  .in1({ S1497, S885 }),
  .out1({ S1498 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_472_ (
  .in1({ S1496, S886 }),
  .out1({ S1499 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_473_ (
  .in1({ S1499, S1498 }),
  .out1({ S1501 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_147_ (
  .in1({ S1501 }),
  .out1({ S1502 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_474_ (
  .in1({ S1434, DP_AC_dout_5 }),
  .out1({ S1503 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_148_ (
  .in1({ S1503 }),
  .out1({ S1504 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_475_ (
  .in1({ S1435, S1263 }),
  .out1({ S1505 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_476_ (
  .in1({ S1505, S1503 }),
  .out1({ S1506 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_149_ (
  .in1({ S1506 }),
  .out1({ S1507 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_477_ (
  .in1({ S1506, S1501 }),
  .out1({ S1508 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_150_ (
  .in1({ S1508 }),
  .out1({ S1509 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_323_ (
  .in1({ S1506, S1501 }),
  .out1({ S1510 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_478_ (
  .in1({ S1507, S1502 }),
  .out1({ S1512 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_324_ (
  .in1({ S1510, S1509 }),
  .out1({ S1513 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_479_ (
  .in1({ S1512, S1508 }),
  .out1({ S1514 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_325_ (
  .in1({ S1513, S1495 }),
  .out1({ S1515 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_480_ (
  .in1({ S1514, S1494 }),
  .out1({ S1516 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_326_ (
  .in1({ S1514, S1494 }),
  .out1({ S1517 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_481_ (
  .in1({ S1513, S1495 }),
  .out1({ S1518 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_327_ (
  .in1({ S1517, S1515 }),
  .out1({ S1519 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_482_ (
  .in1({ S1518, S1516 }),
  .out1({ S1520 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_328_ (
  .in1({ S1520, S1428 }),
  .out1({ S1521 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_483_ (
  .in1({ S1519, S1427 }),
  .out1({ S1523 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_329_ (
  .in1({ S1519, S1427 }),
  .out1({ S1524 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_484_ (
  .in1({ S1520, S1428 }),
  .out1({ S1525 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_330_ (
  .in1({ S1524, S1521 }),
  .out1({ S1526 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_485_ (
  .in1({ S1525, S1523 }),
  .out1({ S1527 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_486_ (
  .in1({ S1527, S1492 }),
  .out1({ S1528 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_487_ (
  .in1({ S1526, S1493 }),
  .out1({ S1529 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_151_ (
  .in1({ S1529 }),
  .out1({ S1530 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_488_ (
  .in1({ S1529, S1528 }),
  .out1({ S1531 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_152_ (
  .in1({ S1531 }),
  .out1({ S1532 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_489_ (
  .in1({ S1531, S1490 }),
  .out1({ S1534 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_490_ (
  .in1({ S1532, S1491 }),
  .out1({ S1535 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_153_ (
  .in1({ S1535 }),
  .out1({ S1536 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_491_ (
  .in1({ S1535, S1534 }),
  .out1({ S1537 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_154_ (
  .in1({ S1537 }),
  .out1({ S1538 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_331_ (
  .in1({ S1538, S1488 }),
  .out1({ S1539 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_332_ (
  .in1({ S1537, S1487 }),
  .out1({ S1540 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_492_ (
  .in1({ S1538, S1488 }),
  .out1({ S1541 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_333_ (
  .in1({ S1540, S1539 }),
  .out1({ S1542 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_493_ (
  .in1({ S1542, S1393 }),
  .out1({ S1543 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_494_ (
  .in1({ DP_ARU1_in1_12, DP_AC_dout_12 }),
  .out1({ S1545 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_155_ (
  .in1({ S1545 }),
  .out1({ S1546 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_334_ (
  .in1({ DP_ARU1_in1_12, DP_AC_dout_12 }),
  .out1({ S1547 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_335_ (
  .in1({ S1547, S1546 }),
  .out1({ S1548 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_336_ (
  .in1({ S1410, S1409 }),
  .out1({ S1549 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_337_ (
  .in1({ S1549, S1411 }),
  .out1({ S1550 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_338_ (
  .in1({ S1550, S1548 }),
  .out1({ S1551 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_495_ (
  .in1({ S1550, S1548 }),
  .out1({ S1552 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_156_ (
  .in1({ S1552 }),
  .out1({ S1553 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_339_ (
  .in1({ S1553, S1551 }),
  .out1({ S1554 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_496_ (
  .in1({ S1554, S59 }),
  .out1({ S1556 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_497_ (
  .in1({ S1556, S1543 }),
  .out1({ DP_ARU1_out_12 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_498_ (
  .in1({ S1552, S1545 }),
  .out1({ S1557 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_499_ (
  .in1({ DP_ARU1_in1_13, DP_AC_dout_13 }),
  .out1({ S1558 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_157_ (
  .in1({ S1558 }),
  .out1({ S1559 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_340_ (
  .in1({ DP_ARU1_in1_13, DP_AC_dout_13 }),
  .out1({ S1560 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_341_ (
  .in1({ S1560, S1559 }),
  .out1({ S1561 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_342_ (
  .in1({ S1561, S1557 }),
  .out1({ S1562 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_500_ (
  .in1({ S1561, S1557 }),
  .out1({ S1563 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_501_ (
  .in1({ S1563, S60 }),
  .out1({ S1564 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_343_ (
  .in1({ S1564, S1562 }),
  .out1({ S1566 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_344_ (
  .in1({ S1540, S1536 }),
  .out1({ S1567 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_502_ (
  .in1({ S1541, S1535 }),
  .out1({ S1568 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_345_ (
  .in1({ S1521, S1517 }),
  .out1({ S1569 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_158_ (
  .in1({ S1569 }),
  .out1({ S1570 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_346_ (
  .in1({ S1510, S1504 }),
  .out1({ S1571 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_347_ (
  .in1({ S990, S886 }),
  .out1({ S1572 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_503_ (
  .in1({ S989, S885 }),
  .out1({ S1573 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_504_ (
  .in1({ S1354, S1246 }),
  .out1({ S1574 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_505_ (
  .in1({ S1574, S1573 }),
  .out1({ S1575 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_506_ (
  .in1({ S1575, S1571 }),
  .out1({ S1577 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_348_ (
  .in1({ S1575, S1571 }),
  .out1({ S1578 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_159_ (
  .in1({ S1578 }),
  .out1({ S1579 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_507_ (
  .in1({ S1579, S1577 }),
  .out1({ S1580 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_349_ (
  .in1({ S1580, S1498 }),
  .out1({ S1581 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_160_ (
  .in1({ S1581 }),
  .out1({ S1582 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_508_ (
  .in1({ S1580, S1498 }),
  .out1({ S1583 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_509_ (
  .in1({ S1583, S1582 }),
  .out1({ S1584 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_161_ (
  .in1({ S1584 }),
  .out1({ S1585 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_510_ (
  .in1({ S1584, S1569 }),
  .out1({ S1586 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_511_ (
  .in1({ S1585, S1570 }),
  .out1({ S578 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_162_ (
  .in1({ S578 }),
  .out1({ S579 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_512_ (
  .in1({ S578, S1586 }),
  .out1({ S580 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_163_ (
  .in1({ S580 }),
  .out1({ S581 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_513_ (
  .in1({ S581, S1530 }),
  .out1({ S582 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_164_ (
  .in1({ S582 }),
  .out1({ S583 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_514_ (
  .in1({ S580, S1529 }),
  .out1({ S584 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_515_ (
  .in1({ S584, S582 }),
  .out1({ S585 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_165_ (
  .in1({ S585 }),
  .out1({ S586 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_516_ (
  .in1({ S585, S1567 }),
  .out1({ S587 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_350_ (
  .in1({ S585, S1567 }),
  .out1({ S589 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_517_ (
  .in1({ S586, S1568 }),
  .out1({ S590 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_518_ (
  .in1({ S590, S587 }),
  .out1({ S591 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_351_ (
  .in1({ S591, S1404 }),
  .out1({ S592 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_352_ (
  .in1({ S592, S1566 }),
  .out1({ S593 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_166_ (
  .in1({ S593 }),
  .out1({ DP_ARU1_out_13 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_519_ (
  .in1({ DP_ARU1_in1_14, DP_AC_dout_14 }),
  .out1({ S594 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_167_ (
  .in1({ S594 }),
  .out1({ S595 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_353_ (
  .in1({ DP_ARU1_in1_14, DP_AC_dout_14 }),
  .out1({ S596 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_354_ (
  .in1({ S596, S595 }),
  .out1({ S597 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_355_ (
  .in1({ S1559, S1557 }),
  .out1({ S599 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_356_ (
  .in1({ S599, S1560 }),
  .out1({ S600 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_520_ (
  .in1({ S600, S597 }),
  .out1({ S601 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_357_ (
  .in1({ S600, S597 }),
  .out1({ S602 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_521_ (
  .in1({ S601, S61 }),
  .out1({ S603 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_358_ (
  .in1({ S603, S602 }),
  .out1({ S604 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_359_ (
  .in1({ S589, S583 }),
  .out1({ S605 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_522_ (
  .in1({ S590, S582 }),
  .out1({ S606 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_360_ (
  .in1({ S1581, S1578 }),
  .out1({ S607 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_523_ (
  .in1({ S989, S886 }),
  .out1({ S608 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_524_ (
  .in1({ S608, S607 }),
  .out1({ S610 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_168_ (
  .in1({ S610 }),
  .out1({ S611 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_361_ (
  .in1({ S608, S607 }),
  .out1({ S612 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_169_ (
  .in1({ S612 }),
  .out1({ S613 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_362_ (
  .in1({ S612, S611 }),
  .out1({ S614 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_525_ (
  .in1({ S613, S610 }),
  .out1({ S615 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_526_ (
  .in1({ S614, S579 }),
  .out1({ S616 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_527_ (
  .in1({ S615, S578 }),
  .out1({ S617 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_528_ (
  .in1({ S617, S616 }),
  .out1({ S618 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_170_ (
  .in1({ S618 }),
  .out1({ S619 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_529_ (
  .in1({ S618, S605 }),
  .out1({ S621 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_363_ (
  .in1({ S618, S605 }),
  .out1({ S622 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_530_ (
  .in1({ S619, S606 }),
  .out1({ S623 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_531_ (
  .in1({ S623, S621 }),
  .out1({ S624 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_364_ (
  .in1({ S624, S1404 }),
  .out1({ S625 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_365_ (
  .in1({ S625, S604 }),
  .out1({ S626 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_171_ (
  .in1({ S626 }),
  .out1({ DP_ARU1_out_14 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_366_ (
  .in1({ S612, S1572 }),
  .out1({ S627 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_532_ (
  .in1({ S627, S616 }),
  .out1({ S628 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_367_ (
  .in1({ S628, S622 }),
  .out1({ S629 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_368_ (
  .in1({ S629, S1404 }),
  .out1({ S630 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_533_ (
  .in1({ S601, S594 }),
  .out1({ S631 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_369_ (
  .in1({ S1327, S1316 }),
  .out1({ S632 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_370_ (
  .in1({ DP_ARU1_in1_15, DP_AC_dout_15 }),
  .out1({ S633 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_534_ (
  .in1({ S1327, S1316 }),
  .out1({ S634 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_371_ (
  .in1({ S633, S632 }),
  .out1({ S635 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_535_ (
  .in1({ S635, S631 }),
  .out1({ S636 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_372_ (
  .in1({ S635, S631 }),
  .out1({ S637 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_536_ (
  .in1({ S636, S62 }),
  .out1({ S638 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_373_ (
  .in1({ S638, S637 }),
  .out1({ S639 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_374_ (
  .in1({ S639, S630 }),
  .out1({ S641 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_172_ (
  .in1({ S641 }),
  .out1({ DP_ARU1_N })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_537_ (
  .in1({ S620, S1436 }),
  .out1({ S642 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_375_ (
  .in1({ S642, DP_ARU1_out_2 }),
  .out1({ S643 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_538_ (
  .in1({ S643, S729 }),
  .out1({ S644 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_376_ (
  .in1({ S644, DP_ARU1_out_4 }),
  .out1({ S645 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_539_ (
  .in1({ S645, S882 }),
  .out1({ S646 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_377_ (
  .in1({ S646, DP_ARU1_out_6 }),
  .out1({ S647 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_540_ (
  .in1({ S647, S1102 }),
  .out1({ S648 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_378_ (
  .in1({ S648, DP_ARU1_out_8 }),
  .out1({ S649 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_541_ (
  .in1({ S649, S1315 }),
  .out1({ S651 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_379_ (
  .in1({ S651, DP_ARU1_out_10 }),
  .out1({ S652 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_542_ (
  .in1({ S652, S1486 }),
  .out1({ S653 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_380_ (
  .in1({ S653, DP_ARU1_out_12 }),
  .out1({ S654 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_543_ (
  .in1({ S654, S593 }),
  .out1({ S655 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_544_ (
  .in1({ S641, S626 }),
  .out1({ S656 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_381_ (
  .in1({ S656, S655 }),
  .out1({ DP_ARU1_Z })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_545_ (
  .in1({ S641, S632 }),
  .out1({ S657 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_546_ (
  .in1({ DP_ARU1_N, S633 }),
  .out1({ S658 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_547_ (
  .in1({ S658, S657 }),
  .out1({ DP_ARU1_V })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_382_ (
  .in1({ S632, S631 }),
  .out1({ S660 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_548_ (
  .in1({ S634, S63 }),
  .out1({ S661 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_383_ (
  .in1({ S661, S660 }),
  .out1({ DP_ARU1_C })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_173_ (
  .in1({ CU_inst_0 }),
  .out1({ S1588 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_174_ (
  .in1({ S64 }),
  .out1({ S1589 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_175_ (
  .in1({ S65 }),
  .out1({ S1590 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_176_ (
  .in1({ CU_inst_1 }),
  .out1({ S1591 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_177_ (
  .in1({ CU_inst_2 }),
  .out1({ S1592 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_178_ (
  .in1({ CU_inst_3 }),
  .out1({ S1593 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_384_ (
  .in1({ S67, S66 }),
  .out1({ S1594 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_179_ (
  .in1({ S1594 }),
  .out1({ S1595 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_385_ (
  .in1({ S1595, S68 }),
  .out1({ S1596 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_386_ (
  .in1({ S1596, S1588 }),
  .out1({ DP_IMM1_out_0 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_387_ (
  .in1({ S1596, S1591 }),
  .out1({ DP_IMM1_out_1 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_388_ (
  .in1({ S1596, S1592 }),
  .out1({ DP_IMM1_out_2 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_389_ (
  .in1({ S1596, S1593 }),
  .out1({ DP_IMM1_out_3 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_549_ (
  .in1({ S1589, S69 }),
  .out1({ S1597 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_550_ (
  .in1({ S1597, S1590 }),
  .out1({ S1598 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_551_ (
  .in1({ S1598, CU_inst_4 }),
  .out1({ S1599 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_390_ (
  .in1({ S70, S1589 }),
  .out1({ S1600 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_552_ (
  .in1({ CU_inst_3, S71 }),
  .out1({ S1601 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_391_ (
  .in1({ S1601, S72 }),
  .out1({ S1602 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_553_ (
  .in1({ S1600, CU_inst_3 }),
  .out1({ S1603 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_554_ (
  .in1({ S1603, S1599 }),
  .out1({ DP_IMM1_out_4 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_555_ (
  .in1({ S1598, CU_inst_5 }),
  .out1({ S1604 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_556_ (
  .in1({ S1604, S1603 }),
  .out1({ DP_IMM1_out_5 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_557_ (
  .in1({ S1598, CU_inst_6 }),
  .out1({ S1605 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_558_ (
  .in1({ S1605, S1603 }),
  .out1({ DP_IMM1_out_6 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_559_ (
  .in1({ S1598, CU_inst_7 }),
  .out1({ S1606 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_560_ (
  .in1({ S1606, S1603 }),
  .out1({ DP_IMM1_out_7 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_561_ (
  .in1({ S1598, CU_inst_8 }),
  .out1({ S1607 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_562_ (
  .in1({ S1607, S1603 }),
  .out1({ DP_IMM1_out_8 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_563_ (
  .in1({ S1598, CU_inst_9 }),
  .out1({ S1608 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_564_ (
  .in1({ S1608, S1603 }),
  .out1({ DP_IMM1_out_9 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_565_ (
  .in1({ S1598, CU_inst_10 }),
  .out1({ S1609 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_566_ (
  .in1({ S1609, S1603 }),
  .out1({ DP_IMM1_out_10 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_567_ (
  .in1({ S1598, CU_inst_11 }),
  .out1({ S1610 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_568_ (
  .in1({ S1610, S1603 }),
  .out1({ DP_IMM1_out_11 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_569_ (
  .in1({ S1594, S73 }),
  .out1({ S1611 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_570_ (
  .in1({ S1611, S1590 }),
  .out1({ S1612 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_571_ (
  .in1({ S1612, DP_IMM1_in1_0 }),
  .out1({ S1613 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_572_ (
  .in1({ CU_inst_11, S1590 }),
  .out1({ S1614 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_392_ (
  .in1({ S1614, S1597 }),
  .out1({ S1615 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_393_ (
  .in1({ S1615, S1602 }),
  .out1({ S1616 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_573_ (
  .in1({ S1616, S1613 }),
  .out1({ DP_IMM1_out_12 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_574_ (
  .in1({ S1612, DP_IMM1_in1_1 }),
  .out1({ S1617 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_575_ (
  .in1({ S1617, S1616 }),
  .out1({ DP_IMM1_out_13 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_576_ (
  .in1({ S1612, DP_IMM1_in1_2 }),
  .out1({ S1618 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_577_ (
  .in1({ S1618, S1616 }),
  .out1({ DP_IMM1_out_14 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_578_ (
  .in1({ S1612, DP_IMM1_in1_3 }),
  .out1({ S1619 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_579_ (
  .in1({ S1619, S1616 }),
  .out1({ DP_IMM1_out_15 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_180_ (
  .in1({ S74 }),
  .out1({ S1637 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_394_ (
  .in1({ S76, S75 }),
  .out1({ S1638 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_580_ (
  .in1({ S1638, DP_IN_dout_0 }),
  .out1({ S1639 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_395_ (
  .in1({ S1637, S77 }),
  .out1({ S1640 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_581_ (
  .in1({ S1640, DP_IN_din_0 }),
  .out1({ S1641 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_582_ (
  .in1({ S1641, S1639 }),
  .out1({ S1620 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_583_ (
  .in1({ S1638, DP_IN_dout_1 }),
  .out1({ S1642 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_584_ (
  .in1({ S1640, DP_IN_din_1 }),
  .out1({ S1643 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_585_ (
  .in1({ S1643, S1642 }),
  .out1({ S1621 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_586_ (
  .in1({ S1638, DP_IN_dout_2 }),
  .out1({ S1644 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_587_ (
  .in1({ S1640, DP_IN_din_2 }),
  .out1({ S1645 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_588_ (
  .in1({ S1645, S1644 }),
  .out1({ S1622 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_589_ (
  .in1({ S1638, DP_IN_dout_3 }),
  .out1({ S1646 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_590_ (
  .in1({ S1640, DP_IN_din_3 }),
  .out1({ S1647 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_591_ (
  .in1({ S1647, S1646 }),
  .out1({ S1623 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_592_ (
  .in1({ S1638, DP_IN_dout_4 }),
  .out1({ S1648 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_593_ (
  .in1({ S1640, DP_IN_din_4 }),
  .out1({ S1649 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_594_ (
  .in1({ S1649, S1648 }),
  .out1({ S1624 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_595_ (
  .in1({ S1638, DP_IN_dout_5 }),
  .out1({ S1650 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_596_ (
  .in1({ S1640, DP_IN_din_5 }),
  .out1({ S1651 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_597_ (
  .in1({ S1651, S1650 }),
  .out1({ S1625 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_598_ (
  .in1({ S1638, DP_IN_dout_6 }),
  .out1({ S1652 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_599_ (
  .in1({ S1640, DP_IN_din_6 }),
  .out1({ S1653 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_600_ (
  .in1({ S1653, S1652 }),
  .out1({ S1626 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_601_ (
  .in1({ S1638, DP_IN_dout_7 }),
  .out1({ S1654 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_602_ (
  .in1({ S1640, DP_IN_din_7 }),
  .out1({ S1655 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_603_ (
  .in1({ S1655, S1654 }),
  .out1({ S1627 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_604_ (
  .in1({ S1638, DP_IN_dout_8 }),
  .out1({ S1656 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_605_ (
  .in1({ S1640, DP_IN_din_8 }),
  .out1({ S1657 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_606_ (
  .in1({ S1657, S1656 }),
  .out1({ S1628 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_607_ (
  .in1({ S1638, DP_IN_dout_9 }),
  .out1({ S1658 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_608_ (
  .in1({ S1640, DP_IN_din_9 }),
  .out1({ S1659 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_609_ (
  .in1({ S1659, S1658 }),
  .out1({ S1629 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_610_ (
  .in1({ S1638, DP_IN_dout_10 }),
  .out1({ S1660 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_611_ (
  .in1({ S1640, DP_IN_din_10 }),
  .out1({ S1661 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_612_ (
  .in1({ S1661, S1660 }),
  .out1({ S1630 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_613_ (
  .in1({ S1638, DP_IN_dout_11 }),
  .out1({ S1662 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_614_ (
  .in1({ S1640, DP_IN_din_11 }),
  .out1({ S1663 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_615_ (
  .in1({ S1663, S1662 }),
  .out1({ S1631 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_616_ (
  .in1({ S1638, DP_IN_dout_12 }),
  .out1({ S1664 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_617_ (
  .in1({ S1640, DP_IN_din_12 }),
  .out1({ S1665 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_618_ (
  .in1({ S1665, S1664 }),
  .out1({ S1632 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_619_ (
  .in1({ S1638, DP_IN_dout_13 }),
  .out1({ S1666 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_620_ (
  .in1({ S1640, DP_IN_din_13 }),
  .out1({ S1667 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_621_ (
  .in1({ S1667, S1666 }),
  .out1({ S1633 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_622_ (
  .in1({ S1638, DP_IN_dout_14 }),
  .out1({ S1668 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_623_ (
  .in1({ S1640, DP_IN_din_14 }),
  .out1({ S1669 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_624_ (
  .in1({ S1669, S1668 }),
  .out1({ S1634 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_625_ (
  .in1({ S1638, DP_IN_dout_15 }),
  .out1({ S1670 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_626_ (
  .in1({ S1640, DP_IN_din_15 }),
  .out1({ S1636 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_627_ (
  .in1({ S1636, S1670 }),
  .out1({ S1635 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_17_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1620 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_dout_0 }),
  .Si({ S3390 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_18_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1621 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_dout_1 }),
  .Si({ S3389 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_19_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1622 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_dout_2 }),
  .Si({ S3388 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_20_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1623 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_dout_3 }),
  .Si({ S3387 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_21_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1624 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_dout_4 }),
  .Si({ S3386 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_22_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1625 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_dout_5 }),
  .Si({ S3385 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_23_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1626 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_dout_6 }),
  .Si({ S3384 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_24_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1627 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_dout_7 }),
  .Si({ S3383 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_25_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1628 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_dout_8 }),
  .Si({ S3382 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_26_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1629 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_dout_9 }),
  .Si({ S3381 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_27_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1630 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_dout_10 }),
  .Si({ S3380 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_28_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1631 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_dout_11 }),
  .Si({ S3379 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_29_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1632 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_dout_12 }),
  .Si({ S3378 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_30_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1633 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_dout_13 }),
  .Si({ S3377 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_31_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1634 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_dout_14 }),
  .Si({ S3376 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_32_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1635 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IN_dout_15 }),
  .Si({ S3425 }),
  .global_reset({ 1'b0 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_181_ (
  .in1({ DP_INC_1_in_1 }),
  .out1({ S1688 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_182_ (
  .in1({ DP_INC_1_inc_value_1 }),
  .out1({ S1689 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_183_ (
  .in1({ DP_INC_1_in_0 }),
  .out1({ S1690 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_184_ (
  .in1({ DP_INC_1_inc_value_0 }),
  .out1({ S1691 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_185_ (
  .in1({ DP_INC_1_in_2 }),
  .out1({ S1692 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_186_ (
  .in1({ DP_INC_1_in_3 }),
  .out1({ S1693 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_187_ (
  .in1({ DP_INC_1_in_4 }),
  .out1({ S1694 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_188_ (
  .in1({ DP_INC_1_in_5 }),
  .out1({ S1695 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_189_ (
  .in1({ DP_INC_1_in_6 }),
  .out1({ S1696 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_190_ (
  .in1({ DP_INC_1_in_7 }),
  .out1({ S1697 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_191_ (
  .in1({ DP_INC_1_in_8 }),
  .out1({ S1698 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_192_ (
  .in1({ DP_INC_1_in_9 }),
  .out1({ S1699 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_193_ (
  .in1({ DP_INC_1_in_10 }),
  .out1({ S1700 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_194_ (
  .in1({ DP_INC_1_in_11 }),
  .out1({ S1701 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_195_ (
  .in1({ DP_INC_1_in_12 }),
  .out1({ S1702 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_196_ (
  .in1({ DP_INC_1_in_13 }),
  .out1({ S1703 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_197_ (
  .in1({ DP_INC_1_in_14 }),
  .out1({ S1704 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_198_ (
  .in1({ DP_INC_1_in_15 }),
  .out1({ S1705 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_396_ (
  .in1({ S1691, S1690 }),
  .out1({ S1706 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_628_ (
  .in1({ DP_INC_1_inc_value_0, DP_INC_1_in_0 }),
  .out1({ S1707 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_397_ (
  .in1({ S1689, S1688 }),
  .out1({ S1708 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_629_ (
  .in1({ DP_INC_1_inc_value_1, DP_INC_1_in_1 }),
  .out1({ S1709 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_398_ (
  .in1({ DP_INC_1_inc_value_1, DP_INC_1_in_1 }),
  .out1({ S1710 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_199_ (
  .in1({ S1710 }),
  .out1({ S1711 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_399_ (
  .in1({ S1710, S1708 }),
  .out1({ S1712 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_630_ (
  .in1({ S1711, S1709 }),
  .out1({ S1713 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_400_ (
  .in1({ S1713, S1707 }),
  .out1({ S1714 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_631_ (
  .in1({ S1712, S1706 }),
  .out1({ S1715 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_401_ (
  .in1({ S1712, S1706 }),
  .out1({ S1716 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_402_ (
  .in1({ S1716, S1714 }),
  .out1({ DP_INC_1_out_1 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_403_ (
  .in1({ S1714, S1708 }),
  .out1({ S1717 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_632_ (
  .in1({ S1715, S1709 }),
  .out1({ S1718 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_404_ (
  .in1({ S1717, S1692 }),
  .out1({ S1719 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_633_ (
  .in1({ S1718, DP_INC_1_in_2 }),
  .out1({ S1720 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_405_ (
  .in1({ S1718, DP_INC_1_in_2 }),
  .out1({ S1721 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_406_ (
  .in1({ S1721, S1719 }),
  .out1({ DP_INC_1_out_2 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_407_ (
  .in1({ S1720, S1693 }),
  .out1({ S1722 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_634_ (
  .in1({ S1719, DP_INC_1_in_3 }),
  .out1({ S1723 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_408_ (
  .in1({ S1719, DP_INC_1_in_3 }),
  .out1({ S1724 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_409_ (
  .in1({ S1724, S1722 }),
  .out1({ DP_INC_1_out_3 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_410_ (
  .in1({ S1723, S1694 }),
  .out1({ S1725 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_635_ (
  .in1({ S1722, DP_INC_1_in_4 }),
  .out1({ S1726 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_411_ (
  .in1({ S1722, DP_INC_1_in_4 }),
  .out1({ S1727 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_412_ (
  .in1({ S1727, S1725 }),
  .out1({ DP_INC_1_out_4 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_413_ (
  .in1({ S1726, S1695 }),
  .out1({ S1728 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_636_ (
  .in1({ S1725, DP_INC_1_in_5 }),
  .out1({ S1729 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_414_ (
  .in1({ S1725, DP_INC_1_in_5 }),
  .out1({ S1730 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_415_ (
  .in1({ S1730, S1728 }),
  .out1({ DP_INC_1_out_5 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_416_ (
  .in1({ S1729, S1696 }),
  .out1({ S1731 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_637_ (
  .in1({ S1728, DP_INC_1_in_6 }),
  .out1({ S1732 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_417_ (
  .in1({ S1728, DP_INC_1_in_6 }),
  .out1({ S1733 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_418_ (
  .in1({ S1733, S1731 }),
  .out1({ DP_INC_1_out_6 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_419_ (
  .in1({ S1732, S1697 }),
  .out1({ S1734 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_638_ (
  .in1({ S1731, DP_INC_1_in_7 }),
  .out1({ S1735 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_420_ (
  .in1({ S1731, DP_INC_1_in_7 }),
  .out1({ S1736 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_421_ (
  .in1({ S1736, S1734 }),
  .out1({ DP_INC_1_out_7 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_422_ (
  .in1({ S1735, S1698 }),
  .out1({ S1737 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_639_ (
  .in1({ S1734, DP_INC_1_in_8 }),
  .out1({ S1738 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_423_ (
  .in1({ S1734, DP_INC_1_in_8 }),
  .out1({ S1739 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_424_ (
  .in1({ S1739, S1737 }),
  .out1({ DP_INC_1_out_8 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_425_ (
  .in1({ S1738, S1699 }),
  .out1({ S1740 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_640_ (
  .in1({ S1737, DP_INC_1_in_9 }),
  .out1({ S1741 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_426_ (
  .in1({ S1737, DP_INC_1_in_9 }),
  .out1({ S1742 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_427_ (
  .in1({ S1742, S1740 }),
  .out1({ DP_INC_1_out_9 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_428_ (
  .in1({ S1741, S1700 }),
  .out1({ S1743 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_641_ (
  .in1({ S1740, DP_INC_1_in_10 }),
  .out1({ S1671 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_429_ (
  .in1({ S1740, DP_INC_1_in_10 }),
  .out1({ S1672 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_430_ (
  .in1({ S1672, S1743 }),
  .out1({ DP_INC_1_out_10 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_431_ (
  .in1({ S1671, S1701 }),
  .out1({ S1673 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_642_ (
  .in1({ S1743, DP_INC_1_in_11 }),
  .out1({ S1674 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_432_ (
  .in1({ S1743, DP_INC_1_in_11 }),
  .out1({ S1675 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_433_ (
  .in1({ S1675, S1673 }),
  .out1({ DP_INC_1_out_11 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_434_ (
  .in1({ S1674, S1702 }),
  .out1({ S1676 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_643_ (
  .in1({ S1673, DP_INC_1_in_12 }),
  .out1({ S1677 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_435_ (
  .in1({ S1673, DP_INC_1_in_12 }),
  .out1({ S1678 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_436_ (
  .in1({ S1678, S1676 }),
  .out1({ DP_INC_1_out_12 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_437_ (
  .in1({ S1677, S1703 }),
  .out1({ S1679 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_644_ (
  .in1({ S1676, DP_INC_1_in_13 }),
  .out1({ S1680 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_438_ (
  .in1({ S1676, DP_INC_1_in_13 }),
  .out1({ S1681 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_439_ (
  .in1({ S1681, S1679 }),
  .out1({ DP_INC_1_out_13 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_440_ (
  .in1({ S1680, S1704 }),
  .out1({ S1682 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_645_ (
  .in1({ S1679, DP_INC_1_in_14 }),
  .out1({ S1683 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_441_ (
  .in1({ S1679, DP_INC_1_in_14 }),
  .out1({ S1684 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_442_ (
  .in1({ S1684, S1682 }),
  .out1({ DP_INC_1_out_14 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_443_ (
  .in1({ S1682, DP_INC_1_in_15 }),
  .out1({ S1685 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_444_ (
  .in1({ S1683, S1705 }),
  .out1({ S1686 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_445_ (
  .in1({ S1686, S1685 }),
  .out1({ DP_INC_1_out_15 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_446_ (
  .in1({ DP_INC_1_inc_value_0, DP_INC_1_in_0 }),
  .out1({ S1687 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_447_ (
  .in1({ S1687, S1706 }),
  .out1({ DP_INC_1_out_0 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_200_ (
  .in1({ DP_INC_2_in_1 }),
  .out1({ S1761 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_201_ (
  .in1({ S78 }),
  .out1({ S1762 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_202_ (
  .in1({ DP_INC_2_in_0 }),
  .out1({ S1763 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_203_ (
  .in1({ S0 }),
  .out1({ S1764 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_204_ (
  .in1({ DP_INC_2_in_2 }),
  .out1({ S1765 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_205_ (
  .in1({ DP_INC_2_in_3 }),
  .out1({ S1766 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_206_ (
  .in1({ DP_INC_2_in_4 }),
  .out1({ S1767 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_207_ (
  .in1({ DP_INC_2_in_5 }),
  .out1({ S1768 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_208_ (
  .in1({ DP_INC_2_in_6 }),
  .out1({ S1769 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_209_ (
  .in1({ DP_INC_2_in_7 }),
  .out1({ S1770 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_210_ (
  .in1({ DP_INC_2_in_8 }),
  .out1({ S1771 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_211_ (
  .in1({ DP_INC_2_in_9 }),
  .out1({ S1772 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_212_ (
  .in1({ DP_INC_2_in_10 }),
  .out1({ S1773 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_213_ (
  .in1({ DP_INC_2_in_11 }),
  .out1({ S1774 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_214_ (
  .in1({ DP_INC_2_in_12 }),
  .out1({ S1775 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_215_ (
  .in1({ DP_INC_2_in_13 }),
  .out1({ S1776 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_216_ (
  .in1({ DP_INC_2_in_14 }),
  .out1({ S1777 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_217_ (
  .in1({ DP_INC_2_in_15 }),
  .out1({ S1778 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_448_ (
  .in1({ S1764, S1763 }),
  .out1({ S1779 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_646_ (
  .in1({ S1, DP_INC_2_in_0 }),
  .out1({ S1780 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_449_ (
  .in1({ S1762, S1761 }),
  .out1({ S1781 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_647_ (
  .in1({ S79, DP_INC_2_in_1 }),
  .out1({ S1782 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_450_ (
  .in1({ S80, DP_INC_2_in_1 }),
  .out1({ S1783 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_218_ (
  .in1({ S1783 }),
  .out1({ S1784 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_451_ (
  .in1({ S1783, S1781 }),
  .out1({ S1785 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_648_ (
  .in1({ S1784, S1782 }),
  .out1({ S1786 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_452_ (
  .in1({ S1786, S1780 }),
  .out1({ S1787 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_649_ (
  .in1({ S1785, S1779 }),
  .out1({ S1788 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_453_ (
  .in1({ S1785, S1779 }),
  .out1({ S1789 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_454_ (
  .in1({ S1789, S1787 }),
  .out1({ DP_INC2_out_1 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_455_ (
  .in1({ S1787, S1781 }),
  .out1({ S1790 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_650_ (
  .in1({ S1788, S1782 }),
  .out1({ S1791 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_456_ (
  .in1({ S1790, S1765 }),
  .out1({ S1792 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_651_ (
  .in1({ S1791, DP_INC_2_in_2 }),
  .out1({ S1793 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_457_ (
  .in1({ S1791, DP_INC_2_in_2 }),
  .out1({ S1794 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_458_ (
  .in1({ S1794, S1792 }),
  .out1({ DP_INC2_out_2 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_459_ (
  .in1({ S1793, S1766 }),
  .out1({ S1795 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_652_ (
  .in1({ S1792, DP_INC_2_in_3 }),
  .out1({ S1796 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_460_ (
  .in1({ S1792, DP_INC_2_in_3 }),
  .out1({ S1797 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_461_ (
  .in1({ S1797, S1795 }),
  .out1({ DP_INC2_out_3 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_462_ (
  .in1({ S1796, S1767 }),
  .out1({ S1798 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_653_ (
  .in1({ S1795, DP_INC_2_in_4 }),
  .out1({ S1799 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_463_ (
  .in1({ S1795, DP_INC_2_in_4 }),
  .out1({ S1800 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_464_ (
  .in1({ S1800, S1798 }),
  .out1({ DP_INC2_out_4 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_465_ (
  .in1({ S1799, S1768 }),
  .out1({ S1801 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_654_ (
  .in1({ S1798, DP_INC_2_in_5 }),
  .out1({ S1802 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_466_ (
  .in1({ S1798, DP_INC_2_in_5 }),
  .out1({ S1803 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_467_ (
  .in1({ S1803, S1801 }),
  .out1({ DP_INC2_out_5 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_468_ (
  .in1({ S1802, S1769 }),
  .out1({ S1804 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_655_ (
  .in1({ S1801, DP_INC_2_in_6 }),
  .out1({ S1805 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_469_ (
  .in1({ S1801, DP_INC_2_in_6 }),
  .out1({ S1806 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_470_ (
  .in1({ S1806, S1804 }),
  .out1({ DP_INC2_out_6 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_471_ (
  .in1({ S1805, S1770 }),
  .out1({ S1807 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_656_ (
  .in1({ S1804, DP_INC_2_in_7 }),
  .out1({ S1808 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_472_ (
  .in1({ S1804, DP_INC_2_in_7 }),
  .out1({ S1809 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_473_ (
  .in1({ S1809, S1807 }),
  .out1({ DP_INC2_out_7 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_474_ (
  .in1({ S1808, S1771 }),
  .out1({ S1810 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_657_ (
  .in1({ S1807, DP_INC_2_in_8 }),
  .out1({ S1811 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_475_ (
  .in1({ S1807, DP_INC_2_in_8 }),
  .out1({ S1812 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_476_ (
  .in1({ S1812, S1810 }),
  .out1({ DP_INC2_out_8 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_477_ (
  .in1({ S1811, S1772 }),
  .out1({ S1813 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_658_ (
  .in1({ S1810, DP_INC_2_in_9 }),
  .out1({ S1814 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_478_ (
  .in1({ S1810, DP_INC_2_in_9 }),
  .out1({ S1815 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_479_ (
  .in1({ S1815, S1813 }),
  .out1({ DP_INC2_out_9 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_480_ (
  .in1({ S1814, S1773 }),
  .out1({ S1816 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_659_ (
  .in1({ S1813, DP_INC_2_in_10 }),
  .out1({ S1744 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_481_ (
  .in1({ S1813, DP_INC_2_in_10 }),
  .out1({ S1745 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_482_ (
  .in1({ S1745, S1816 }),
  .out1({ DP_INC2_out_10 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_483_ (
  .in1({ S1744, S1774 }),
  .out1({ S1746 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_660_ (
  .in1({ S1816, DP_INC_2_in_11 }),
  .out1({ S1747 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_484_ (
  .in1({ S1816, DP_INC_2_in_11 }),
  .out1({ S1748 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_485_ (
  .in1({ S1748, S1746 }),
  .out1({ DP_INC2_out_11 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_486_ (
  .in1({ S1747, S1775 }),
  .out1({ S1749 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_661_ (
  .in1({ S1746, DP_INC_2_in_12 }),
  .out1({ S1750 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_487_ (
  .in1({ S1746, DP_INC_2_in_12 }),
  .out1({ S1751 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_488_ (
  .in1({ S1751, S1749 }),
  .out1({ DP_INC2_out_12 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_489_ (
  .in1({ S1750, S1776 }),
  .out1({ S1752 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_662_ (
  .in1({ S1749, DP_INC_2_in_13 }),
  .out1({ S1753 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_490_ (
  .in1({ S1749, DP_INC_2_in_13 }),
  .out1({ S1754 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_491_ (
  .in1({ S1754, S1752 }),
  .out1({ DP_INC2_out_13 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_492_ (
  .in1({ S1753, S1777 }),
  .out1({ S1755 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_663_ (
  .in1({ S1752, DP_INC_2_in_14 }),
  .out1({ S1756 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_493_ (
  .in1({ S1752, DP_INC_2_in_14 }),
  .out1({ S1757 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_494_ (
  .in1({ S1757, S1755 }),
  .out1({ DP_INC2_out_14 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_495_ (
  .in1({ S1755, DP_INC_2_in_15 }),
  .out1({ S1758 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_496_ (
  .in1({ S1756, S1778 }),
  .out1({ S1759 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_497_ (
  .in1({ S1759, S1758 }),
  .out1({ DP_INC2_out_15 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_498_ (
  .in1({ S2, DP_INC_2_in_0 }),
  .out1({ S1760 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_499_ (
  .in1({ S1760, S1779 }),
  .out1({ DP_INC2_out_0 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_219_ (
  .in1({ S3 }),
  .out1({ S1834 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_500_ (
  .in1({ S4, S81 }),
  .out1({ S1835 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_664_ (
  .in1({ S1835, CU_inst_0 }),
  .out1({ S1836 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_501_ (
  .in1({ S1834, S82 }),
  .out1({ S1837 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_665_ (
  .in1({ S1837, DP_INC_2_in_0 }),
  .out1({ S1838 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_666_ (
  .in1({ S1838, S1836 }),
  .out1({ S1817 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_667_ (
  .in1({ S1835, CU_inst_1 }),
  .out1({ S1839 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_668_ (
  .in1({ S1837, DP_INC_2_in_1 }),
  .out1({ S1840 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_669_ (
  .in1({ S1840, S1839 }),
  .out1({ S1818 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_670_ (
  .in1({ S1835, CU_inst_2 }),
  .out1({ S1841 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_671_ (
  .in1({ S1837, DP_INC_2_in_2 }),
  .out1({ S1842 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_672_ (
  .in1({ S1842, S1841 }),
  .out1({ S1819 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_673_ (
  .in1({ S1835, CU_inst_3 }),
  .out1({ S1843 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_674_ (
  .in1({ S1837, DP_INC_2_in_3 }),
  .out1({ S1844 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_675_ (
  .in1({ S1844, S1843 }),
  .out1({ S1820 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_676_ (
  .in1({ S1835, CU_inst_4 }),
  .out1({ S1845 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_677_ (
  .in1({ S1837, DP_INC_2_in_4 }),
  .out1({ S1846 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_678_ (
  .in1({ S1846, S1845 }),
  .out1({ S1821 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_679_ (
  .in1({ S1835, CU_inst_5 }),
  .out1({ S1847 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_680_ (
  .in1({ S1837, DP_INC_2_in_5 }),
  .out1({ S1848 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_681_ (
  .in1({ S1848, S1847 }),
  .out1({ S1822 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_682_ (
  .in1({ S1835, CU_inst_6 }),
  .out1({ S1849 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_683_ (
  .in1({ S1837, DP_INC_2_in_6 }),
  .out1({ S1850 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_684_ (
  .in1({ S1850, S1849 }),
  .out1({ S1823 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_685_ (
  .in1({ S1835, CU_inst_7 }),
  .out1({ S1851 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_686_ (
  .in1({ S1837, DP_INC_2_in_7 }),
  .out1({ S1852 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_687_ (
  .in1({ S1852, S1851 }),
  .out1({ S1824 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_688_ (
  .in1({ S1835, CU_inst_8 }),
  .out1({ S1853 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_689_ (
  .in1({ S1837, DP_INC_2_in_8 }),
  .out1({ S1854 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_690_ (
  .in1({ S1854, S1853 }),
  .out1({ S1825 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_691_ (
  .in1({ S1835, CU_inst_9 }),
  .out1({ S1855 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_692_ (
  .in1({ S1837, DP_INC_2_in_9 }),
  .out1({ S1856 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_693_ (
  .in1({ S1856, S1855 }),
  .out1({ S1826 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_694_ (
  .in1({ S1835, CU_inst_10 }),
  .out1({ S1857 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_695_ (
  .in1({ S1837, DP_INC_2_in_10 }),
  .out1({ S1858 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_696_ (
  .in1({ S1858, S1857 }),
  .out1({ S1827 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_697_ (
  .in1({ S1835, CU_inst_11 }),
  .out1({ S1859 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_698_ (
  .in1({ S1837, DP_INC_2_in_11 }),
  .out1({ S1860 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_699_ (
  .in1({ S1860, S1859 }),
  .out1({ S1828 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_700_ (
  .in1({ S1835, CU_inst_12 }),
  .out1({ S1861 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_701_ (
  .in1({ S1837, DP_INC_2_in_12 }),
  .out1({ S1862 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_702_ (
  .in1({ S1862, S1861 }),
  .out1({ S1829 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_703_ (
  .in1({ S1835, CU_inst_13 }),
  .out1({ S1863 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_704_ (
  .in1({ S1837, DP_INC_2_in_13 }),
  .out1({ S1864 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_705_ (
  .in1({ S1864, S1863 }),
  .out1({ S1830 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_706_ (
  .in1({ S1835, CU_inst_14 }),
  .out1({ S1865 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_707_ (
  .in1({ S1837, DP_INC_2_in_14 }),
  .out1({ S1866 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_708_ (
  .in1({ S1866, S1865 }),
  .out1({ S1831 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_709_ (
  .in1({ S1835, CU_inst_15 }),
  .out1({ S1867 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_710_ (
  .in1({ S1837, DP_INC_2_in_15 }),
  .out1({ S1833 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_711_ (
  .in1({ S1833, S1867 }),
  .out1({ S1832 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_33_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1817 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_0 }),
  .Si({ S3405 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_34_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1818 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_1 }),
  .Si({ S3404 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_35_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1819 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_2 }),
  .Si({ S3403 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_36_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1820 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_3 }),
  .Si({ S3402 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_37_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1821 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_4 }),
  .Si({ S3401 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_38_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1822 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_5 }),
  .Si({ S3400 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_39_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1823 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_6 }),
  .Si({ S3399 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_40_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1824 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_7 }),
  .Si({ S3398 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_41_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1825 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_8 }),
  .Si({ S3397 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_42_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1826 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_9 }),
  .Si({ S3396 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_43_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1827 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_10 }),
  .Si({ S3395 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_44_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1828 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_11 }),
  .Si({ S3394 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_45_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1829 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_12 }),
  .Si({ S3393 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_46_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1830 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_13 }),
  .Si({ S3392 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_47_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1831 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_14 }),
  .Si({ S3391 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_48_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S1832 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ CU_inst_15 }),
  .Si({ S3426 }),
  .global_reset({ 1'b0 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_220_ (
  .in1({ DP_AC_dout_0 }),
  .out1({ S2306 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_221_ (
  .in1({ DP_LGU1_in1_3 }),
  .out1({ S2317 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_222_ (
  .in1({ DP_LGU1_in1_1 }),
  .out1({ S2327 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_223_ (
  .in1({ DP_AC_dout_1 }),
  .out1({ S2338 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_224_ (
  .in1({ DP_LGU1_in1_0 }),
  .out1({ S2348 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_225_ (
  .in1({ DP_AC_dout_4 }),
  .out1({ S2359 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_226_ (
  .in1({ DP_AC_dout_5 }),
  .out1({ S2369 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_227_ (
  .in1({ DP_LGU1_in1_2 }),
  .out1({ S2380 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_228_ (
  .in1({ DP_AC_dout_11 }),
  .out1({ S2390 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_229_ (
  .in1({ DP_AC_dout_15 }),
  .out1({ S2401 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_230_ (
  .in1({ S83 }),
  .out1({ S2406 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_231_ (
  .in1({ S84 }),
  .out1({ S2407 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_232_ (
  .in1({ S85 }),
  .out1({ S2408 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_233_ (
  .in1({ S86 }),
  .out1({ S2409 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_234_ (
  .in1({ DP_LGU1_in1_9 }),
  .out1({ S2410 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_235_ (
  .in1({ DP_LGU1_in1_11 }),
  .out1({ S2411 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_502_ (
  .in1({ S2348, S2306 }),
  .out1({ S2412 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_712_ (
  .in1({ DP_LGU1_in1_0, DP_AC_dout_0 }),
  .out1({ S2413 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_713_ (
  .in1({ S2412, S87 }),
  .out1({ S2414 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_503_ (
  .in1({ S88, DP_LGU1_in1_3 }),
  .out1({ S2415 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_236_ (
  .in1({ S2415 }),
  .out1({ S2416 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_714_ (
  .in1({ DP_AC_dout_8, S2348 }),
  .out1({ S2417 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_715_ (
  .in1({ DP_AC_dout_9, DP_LGU1_in1_0 }),
  .out1({ S2418 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_716_ (
  .in1({ S2418, S2417 }),
  .out1({ S2419 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_717_ (
  .in1({ S2419, S2327 }),
  .out1({ S2420 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_718_ (
  .in1({ DP_AC_dout_10, S2348 }),
  .out1({ S2421 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_719_ (
  .in1({ DP_AC_dout_11, DP_LGU1_in1_0 }),
  .out1({ S2422 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_720_ (
  .in1({ S2422, S2421 }),
  .out1({ S2423 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_721_ (
  .in1({ S2423, DP_LGU1_in1_1 }),
  .out1({ S2424 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_722_ (
  .in1({ S2424, S2420 }),
  .out1({ S2425 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_723_ (
  .in1({ S2425, S2380 }),
  .out1({ S2426 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_724_ (
  .in1({ DP_AC_dout_12, S2348 }),
  .out1({ S2427 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_725_ (
  .in1({ DP_AC_dout_13, DP_LGU1_in1_0 }),
  .out1({ S2428 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_726_ (
  .in1({ S2428, S2427 }),
  .out1({ S2429 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_727_ (
  .in1({ S2429, S2327 }),
  .out1({ S2430 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_728_ (
  .in1({ DP_AC_dout_14, S2348 }),
  .out1({ S2431 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_729_ (
  .in1({ DP_AC_dout_15, DP_LGU1_in1_0 }),
  .out1({ S2432 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_730_ (
  .in1({ S2432, S2431 }),
  .out1({ S2433 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_237_ (
  .in1({ S2433 }),
  .out1({ S2434 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_731_ (
  .in1({ S2433, DP_LGU1_in1_1 }),
  .out1({ S2435 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_732_ (
  .in1({ S2435, S2430 }),
  .out1({ S2436 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_733_ (
  .in1({ S2436, DP_LGU1_in1_2 }),
  .out1({ S2437 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_734_ (
  .in1({ S2437, S2426 }),
  .out1({ S2438 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_735_ (
  .in1({ S2438, S2407 }),
  .out1({ S2439 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_736_ (
  .in1({ S2439, S2416 }),
  .out1({ S2440 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_737_ (
  .in1({ DP_AC_dout_2, S2348 }),
  .out1({ S2441 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_738_ (
  .in1({ DP_AC_dout_3, DP_LGU1_in1_0 }),
  .out1({ S1868 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_238_ (
  .in1({ S1868 }),
  .out1({ S1869 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_739_ (
  .in1({ S1868, S2441 }),
  .out1({ S1870 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_740_ (
  .in1({ S1870, DP_LGU1_in1_1 }),
  .out1({ S1871 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_741_ (
  .in1({ S2348, DP_AC_dout_0 }),
  .out1({ S1872 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_504_ (
  .in1({ S1872, DP_LGU1_in1_1 }),
  .out1({ S1873 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_239_ (
  .in1({ S1873 }),
  .out1({ S1874 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_742_ (
  .in1({ DP_LGU1_in1_0, DP_AC_dout_1 }),
  .out1({ S1875 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_743_ (
  .in1({ S1875, S1872 }),
  .out1({ S1876 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_744_ (
  .in1({ S1876, S2327 }),
  .out1({ S1877 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_745_ (
  .in1({ S1877, S1871 }),
  .out1({ S1878 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_746_ (
  .in1({ S1878, S2380 }),
  .out1({ S1879 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_505_ (
  .in1({ S2359, DP_LGU1_in1_0 }),
  .out1({ S1880 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_747_ (
  .in1({ DP_AC_dout_4, S2348 }),
  .out1({ S1881 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_748_ (
  .in1({ DP_AC_dout_5, DP_LGU1_in1_0 }),
  .out1({ S1882 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_240_ (
  .in1({ S1882 }),
  .out1({ S1883 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_506_ (
  .in1({ S1883, S1880 }),
  .out1({ S1884 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_749_ (
  .in1({ S1882, S1881 }),
  .out1({ S1885 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_507_ (
  .in1({ S1884, DP_LGU1_in1_1 }),
  .out1({ S1886 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_750_ (
  .in1({ DP_AC_dout_6, S2348 }),
  .out1({ S1887 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_751_ (
  .in1({ DP_AC_dout_7, DP_LGU1_in1_0 }),
  .out1({ S1888 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_752_ (
  .in1({ S1888, S1887 }),
  .out1({ S1889 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_753_ (
  .in1({ S1889, DP_LGU1_in1_1 }),
  .out1({ S1890 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_241_ (
  .in1({ S1890 }),
  .out1({ S1891 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_508_ (
  .in1({ S1891, S1886 }),
  .out1({ S1892 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_509_ (
  .in1({ S1892, S2380 }),
  .out1({ S1893 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_510_ (
  .in1({ S1893, DP_LGU1_in1_3 }),
  .out1({ S1894 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_754_ (
  .in1({ S1894, S1879 }),
  .out1({ S1895 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_755_ (
  .in1({ S1895, S2440 }),
  .out1({ S1896 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_756_ (
  .in1({ S1873, S2380 }),
  .out1({ S1897 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_511_ (
  .in1({ S2407, S89 }),
  .out1({ S1898 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_757_ (
  .in1({ S90, S2406 }),
  .out1({ S1899 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_512_ (
  .in1({ S1899, DP_LGU1_in1_3 }),
  .out1({ S1900 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_758_ (
  .in1({ S1898, S2317 }),
  .out1({ S1901 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_513_ (
  .in1({ S1901, S1897 }),
  .out1({ S1902 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_514_ (
  .in1({ S1902, S91 }),
  .out1({ S1903 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_759_ (
  .in1({ S1903, S1896 }),
  .out1({ S1904 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_760_ (
  .in1({ S92, DP_AC_dout_0 }),
  .out1({ S1905 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_242_ (
  .in1({ S1905 }),
  .out1({ S1906 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_515_ (
  .in1({ S1906, S93 }),
  .out1({ S1907 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_761_ (
  .in1({ S1907, S1904 }),
  .out1({ S1908 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_762_ (
  .in1({ S1908, S2414 }),
  .out1({ DP_LGU1_out_0 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_516_ (
  .in1({ S95, S94 }),
  .out1({ S1909 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_763_ (
  .in1({ S2407, S2406 }),
  .out1({ S1910 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_764_ (
  .in1({ DP_AC_dout_9, S2348 }),
  .out1({ S1911 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_765_ (
  .in1({ DP_AC_dout_10, DP_LGU1_in1_0 }),
  .out1({ S1912 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_243_ (
  .in1({ S1912 }),
  .out1({ S1913 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_766_ (
  .in1({ S1912, S1911 }),
  .out1({ S1914 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_767_ (
  .in1({ S1914, S2327 }),
  .out1({ S1915 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_517_ (
  .in1({ S2390, DP_LGU1_in1_0 }),
  .out1({ S1916 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_768_ (
  .in1({ DP_AC_dout_11, S2348 }),
  .out1({ S1917 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_769_ (
  .in1({ DP_AC_dout_12, DP_LGU1_in1_0 }),
  .out1({ S1918 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_770_ (
  .in1({ S1918, S1917 }),
  .out1({ S1919 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_244_ (
  .in1({ S1919 }),
  .out1({ S1920 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_771_ (
  .in1({ S1919, DP_LGU1_in1_1 }),
  .out1({ S1921 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_772_ (
  .in1({ S1921, S1915 }),
  .out1({ S1922 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_773_ (
  .in1({ S1922, S2380 }),
  .out1({ S1923 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_774_ (
  .in1({ DP_AC_dout_13, S2348 }),
  .out1({ S1924 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_775_ (
  .in1({ DP_AC_dout_14, DP_LGU1_in1_0 }),
  .out1({ S1925 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_245_ (
  .in1({ S1925 }),
  .out1({ S1926 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_776_ (
  .in1({ S1925, S1924 }),
  .out1({ S1927 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_777_ (
  .in1({ S1927, S2327 }),
  .out1({ S1928 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_778_ (
  .in1({ DP_AC_dout_15, DP_LGU1_in1_1 }),
  .out1({ S1929 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_779_ (
  .in1({ S1929, S1928 }),
  .out1({ S1930 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_780_ (
  .in1({ S1930, DP_LGU1_in1_2 }),
  .out1({ S1931 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_781_ (
  .in1({ S1931, S1923 }),
  .out1({ S1932 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_782_ (
  .in1({ S1932, S1909 }),
  .out1({ S1933 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_518_ (
  .in1({ S96, S2406 }),
  .out1({ S1934 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_783_ (
  .in1({ S2407, S97 }),
  .out1({ S1935 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_519_ (
  .in1({ S2401, DP_LGU1_in1_0 }),
  .out1({ S1936 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_246_ (
  .in1({ S1936 }),
  .out1({ S1937 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_784_ (
  .in1({ S1936, DP_LGU1_in1_1 }),
  .out1({ S1938 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_785_ (
  .in1({ S1938, S1928 }),
  .out1({ S1939 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_786_ (
  .in1({ S1939, DP_LGU1_in1_2 }),
  .out1({ S1940 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_787_ (
  .in1({ S1940, S1923 }),
  .out1({ S1941 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_788_ (
  .in1({ S1941, S1934 }),
  .out1({ S1942 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_789_ (
  .in1({ S1942, S1933 }),
  .out1({ S1943 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_790_ (
  .in1({ S1943, DP_LGU1_in1_3 }),
  .out1({ S1944 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_520_ (
  .in1({ DP_LGU1_in1_0, S2338 }),
  .out1({ S1945 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_791_ (
  .in1({ S2348, DP_AC_dout_1 }),
  .out1({ S1946 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_521_ (
  .in1({ S1945, S2412 }),
  .out1({ S1947 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_792_ (
  .in1({ S1946, S2413 }),
  .out1({ S1948 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_793_ (
  .in1({ S1948, S2327 }),
  .out1({ S1949 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_522_ (
  .in1({ S1949, DP_LGU1_in1_2 }),
  .out1({ S1950 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_794_ (
  .in1({ S1950, S1900 }),
  .out1({ S1951 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_795_ (
  .in1({ DP_AC_dout_2, DP_LGU1_in1_0 }),
  .out1({ S1952 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_796_ (
  .in1({ S1952, S1946 }),
  .out1({ S1953 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_797_ (
  .in1({ S1953, S2327 }),
  .out1({ S1954 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_798_ (
  .in1({ DP_AC_dout_3, S2348 }),
  .out1({ S1955 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_799_ (
  .in1({ DP_AC_dout_4, DP_LGU1_in1_0 }),
  .out1({ S1956 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_800_ (
  .in1({ S1956, S1955 }),
  .out1({ S1957 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_801_ (
  .in1({ S1957, DP_LGU1_in1_1 }),
  .out1({ S1958 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_802_ (
  .in1({ S1958, S1954 }),
  .out1({ S1959 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_803_ (
  .in1({ DP_AC_dout_5, S2348 }),
  .out1({ S1960 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_804_ (
  .in1({ DP_AC_dout_6, DP_LGU1_in1_0 }),
  .out1({ S1961 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_805_ (
  .in1({ S1961, S1960 }),
  .out1({ S1962 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_806_ (
  .in1({ S1962, S2327 }),
  .out1({ S1963 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_807_ (
  .in1({ DP_AC_dout_7, S2348 }),
  .out1({ S1964 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_808_ (
  .in1({ DP_AC_dout_8, DP_LGU1_in1_0 }),
  .out1({ S1965 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_809_ (
  .in1({ S1965, S1964 }),
  .out1({ S1966 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_810_ (
  .in1({ S1966, DP_LGU1_in1_1 }),
  .out1({ S1967 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_811_ (
  .in1({ S1967, S1963 }),
  .out1({ S1968 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_523_ (
  .in1({ S1968, S2380 }),
  .out1({ S1969 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_524_ (
  .in1({ S1959, DP_LGU1_in1_2 }),
  .out1({ S1970 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_525_ (
  .in1({ S1970, S1969 }),
  .out1({ S1971 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_812_ (
  .in1({ S1971, S2415 }),
  .out1({ S1972 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_813_ (
  .in1({ S1972, S1951 }),
  .out1({ S1973 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_526_ (
  .in1({ S1973, S98 }),
  .out1({ S1974 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_814_ (
  .in1({ S1974, S1944 }),
  .out1({ S1975 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_815_ (
  .in1({ S99, DP_AC_dout_1 }),
  .out1({ S1976 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_247_ (
  .in1({ S1976 }),
  .out1({ S1977 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_527_ (
  .in1({ S1977, S100 }),
  .out1({ S1978 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_816_ (
  .in1({ S1978, S1975 }),
  .out1({ S1979 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_528_ (
  .in1({ S2338, S2327 }),
  .out1({ S1980 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_817_ (
  .in1({ S1980, S101 }),
  .out1({ S1981 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_818_ (
  .in1({ S1981, S1979 }),
  .out1({ DP_LGU1_out_1 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_819_ (
  .in1({ DP_LGU1_in1_2, DP_AC_dout_2 }),
  .out1({ S1982 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_529_ (
  .in1({ S1982, S2409 }),
  .out1({ S1983 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_530_ (
  .in1({ S1899, DP_LGU1_in1_2 }),
  .out1({ S1984 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_820_ (
  .in1({ S1898, S2380 }),
  .out1({ S1985 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_821_ (
  .in1({ S1875, S2441 }),
  .out1({ S1986 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_822_ (
  .in1({ S1872, DP_LGU1_in1_1 }),
  .out1({ S1987 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_531_ (
  .in1({ S1986, DP_LGU1_in1_1 }),
  .out1({ S1988 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_248_ (
  .in1({ S1988 }),
  .out1({ S1989 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_823_ (
  .in1({ S1989, S1987 }),
  .out1({ S1990 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_249_ (
  .in1({ S1990 }),
  .out1({ S1991 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_532_ (
  .in1({ S1990, S1985 }),
  .out1({ S1992 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_824_ (
  .in1({ S1991, S1984 }),
  .out1({ S1993 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_533_ (
  .in1({ S1885, S2327 }),
  .out1({ S1994 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_534_ (
  .in1({ S1870, DP_LGU1_in1_1 }),
  .out1({ S1995 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_535_ (
  .in1({ S1995, S1994 }),
  .out1({ S1996 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_536_ (
  .in1({ S1996, DP_LGU1_in1_2 }),
  .out1({ S1997 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_825_ (
  .in1({ S1889, S2327 }),
  .out1({ S1998 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_826_ (
  .in1({ S2419, DP_LGU1_in1_1 }),
  .out1({ S1999 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_827_ (
  .in1({ S1999, S1998 }),
  .out1({ S2000 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_537_ (
  .in1({ S2000, S2380 }),
  .out1({ S2001 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_538_ (
  .in1({ S2001, S1997 }),
  .out1({ S2002 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_539_ (
  .in1({ S2002, DP_LGU1_in1_3 }),
  .out1({ S2003 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_540_ (
  .in1({ S2003, S102 }),
  .out1({ S2004 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_541_ (
  .in1({ S2004, S1992 }),
  .out1({ S2005 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_828_ (
  .in1({ S2423, S2327 }),
  .out1({ S2006 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_829_ (
  .in1({ S2429, DP_LGU1_in1_1 }),
  .out1({ S2007 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_830_ (
  .in1({ S2007, S2006 }),
  .out1({ S2008 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_831_ (
  .in1({ S2008, S2380 }),
  .out1({ S2009 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_542_ (
  .in1({ S2434, DP_LGU1_in1_1 }),
  .out1({ S2010 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_832_ (
  .in1({ S2433, S2327 }),
  .out1({ S2011 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_833_ (
  .in1({ S2011, S1929 }),
  .out1({ S2012 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_834_ (
  .in1({ S2012, DP_LGU1_in1_2 }),
  .out1({ S2013 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_835_ (
  .in1({ S2013, S2009 }),
  .out1({ S2014 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_836_ (
  .in1({ S2014, S1909 }),
  .out1({ S2015 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_837_ (
  .in1({ S2010, DP_LGU1_in1_2 }),
  .out1({ S2016 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_838_ (
  .in1({ S2016, S2009 }),
  .out1({ S2017 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_839_ (
  .in1({ S2017, S1934 }),
  .out1({ S2018 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_250_ (
  .in1({ S2018 }),
  .out1({ S2019 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_840_ (
  .in1({ S2015, DP_LGU1_in1_3 }),
  .out1({ S2020 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_543_ (
  .in1({ S2020, S2019 }),
  .out1({ S2021 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_544_ (
  .in1({ S2021, S2005 }),
  .out1({ S2022 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_545_ (
  .in1({ S2022, S103 }),
  .out1({ S2023 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_841_ (
  .in1({ S104, DP_AC_dout_2 }),
  .out1({ S2024 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_842_ (
  .in1({ S2024, S2409 }),
  .out1({ S2025 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_546_ (
  .in1({ S2025, S2023 }),
  .out1({ S2026 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_547_ (
  .in1({ S2026, S1983 }),
  .out1({ S2027 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_251_ (
  .in1({ S2027 }),
  .out1({ DP_LGU1_out_2 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_843_ (
  .in1({ DP_AC_dout_3, DP_LGU1_in1_3 }),
  .out1({ S2028 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_548_ (
  .in1({ S2028, S2409 }),
  .out1({ S2029 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_844_ (
  .in1({ S1955, S1952 }),
  .out1({ S2030 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_845_ (
  .in1({ S1947, DP_LGU1_in1_1 }),
  .out1({ S2031 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_252_ (
  .in1({ S2031 }),
  .out1({ S2032 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_549_ (
  .in1({ S2030, DP_LGU1_in1_1 }),
  .out1({ S2033 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_253_ (
  .in1({ S2033 }),
  .out1({ S2034 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_846_ (
  .in1({ S2034, S2031 }),
  .out1({ S2035 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_550_ (
  .in1({ S2033, S2032 }),
  .out1({ S2036 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_551_ (
  .in1({ S2035, S1985 }),
  .out1({ S2037 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_847_ (
  .in1({ S2036, S1984 }),
  .out1({ S2038 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_552_ (
  .in1({ S1962, S2327 }),
  .out1({ S2039 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_553_ (
  .in1({ S1957, DP_LGU1_in1_1 }),
  .out1({ S2040 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_554_ (
  .in1({ S2040, S2039 }),
  .out1({ S2041 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_555_ (
  .in1({ S2041, DP_LGU1_in1_2 }),
  .out1({ S2042 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_848_ (
  .in1({ S1966, S2327 }),
  .out1({ S2043 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_849_ (
  .in1({ S1914, DP_LGU1_in1_1 }),
  .out1({ S2044 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_850_ (
  .in1({ S2044, S2043 }),
  .out1({ S2045 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_556_ (
  .in1({ S2045, S2380 }),
  .out1({ S2046 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_557_ (
  .in1({ S2046, S2042 }),
  .out1({ S2047 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_558_ (
  .in1({ S2047, DP_LGU1_in1_3 }),
  .out1({ S2048 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_559_ (
  .in1({ S2048, S105 }),
  .out1({ S2049 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_560_ (
  .in1({ S2049, S2037 }),
  .out1({ S2050 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_561_ (
  .in1({ S1920, DP_LGU1_in1_1 }),
  .out1({ S2051 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_851_ (
  .in1({ S1919, S2327 }),
  .out1({ S2052 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_852_ (
  .in1({ S1927, DP_LGU1_in1_1 }),
  .out1({ S2053 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_254_ (
  .in1({ S2053 }),
  .out1({ S2054 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_562_ (
  .in1({ S2054, S2051 }),
  .out1({ S2055 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_853_ (
  .in1({ S2053, S2052 }),
  .out1({ S2056 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_854_ (
  .in1({ S2056, S2380 }),
  .out1({ S2057 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_855_ (
  .in1({ DP_AC_dout_15, DP_LGU1_in1_2 }),
  .out1({ S2058 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_856_ (
  .in1({ S2058, S2057 }),
  .out1({ S2059 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_255_ (
  .in1({ S2059 }),
  .out1({ S2060 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_563_ (
  .in1({ S2060, S1910 }),
  .out1({ S2061 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_857_ (
  .in1({ S2059, S1909 }),
  .out1({ S2062 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_564_ (
  .in1({ S1937, DP_LGU1_in1_1 }),
  .out1({ S2063 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_858_ (
  .in1({ S2063, DP_LGU1_in1_2 }),
  .out1({ S2064 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_859_ (
  .in1({ S2064, S2057 }),
  .out1({ S2065 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_860_ (
  .in1({ S2065, S1934 }),
  .out1({ S2066 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_861_ (
  .in1({ S2066, DP_LGU1_in1_3 }),
  .out1({ S2067 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_565_ (
  .in1({ S2067, S2061 }),
  .out1({ S2068 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_566_ (
  .in1({ S2068, S2050 }),
  .out1({ S2069 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_567_ (
  .in1({ S2069, S106 }),
  .out1({ S2070 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_862_ (
  .in1({ S107, DP_AC_dout_3 }),
  .out1({ S2071 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_863_ (
  .in1({ S2071, S2409 }),
  .out1({ S2072 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_568_ (
  .in1({ S2072, S2070 }),
  .out1({ S2073 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_569_ (
  .in1({ S2073, S2029 }),
  .out1({ S2074 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_256_ (
  .in1({ S2074 }),
  .out1({ DP_LGU1_out_3 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_864_ (
  .in1({ DP_LGU1_in1_4, DP_AC_dout_4 }),
  .out1({ S2075 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_865_ (
  .in1({ S2075, S108 }),
  .out1({ S2076 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_257_ (
  .in1({ S2076 }),
  .out1({ S2077 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_570_ (
  .in1({ S1880, S1869 }),
  .out1({ S2078 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_571_ (
  .in1({ S2078, DP_LGU1_in1_1 }),
  .out1({ S2079 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_866_ (
  .in1({ S1986, DP_LGU1_in1_1 }),
  .out1({ S2080 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_258_ (
  .in1({ S2080 }),
  .out1({ S2081 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_572_ (
  .in1({ S2081, S2079 }),
  .out1({ S2082 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_573_ (
  .in1({ S2082, S1985 }),
  .out1({ S2083 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_574_ (
  .in1({ S1899, S2380 }),
  .out1({ S2084 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_867_ (
  .in1({ S1898, DP_LGU1_in1_2 }),
  .out1({ S2085 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_575_ (
  .in1({ S2085, S1874 }),
  .out1({ S2086 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_576_ (
  .in1({ S2086, S2083 }),
  .out1({ S2087 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_868_ (
  .in1({ S2425, DP_LGU1_in1_2 }),
  .out1({ S2088 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_577_ (
  .in1({ S1892, DP_LGU1_in1_2 }),
  .out1({ S2089 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_578_ (
  .in1({ S2089, DP_LGU1_in1_3 }),
  .out1({ S2090 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_869_ (
  .in1({ S2090, S2088 }),
  .out1({ S2091 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_870_ (
  .in1({ S2091, S2407 }),
  .out1({ S2092 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_871_ (
  .in1({ S2092, S2087 }),
  .out1({ S2093 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_872_ (
  .in1({ S2436, S2380 }),
  .out1({ S2094 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_873_ (
  .in1({ S2094, S2058 }),
  .out1({ S2095 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_874_ (
  .in1({ S2095, S1909 }),
  .out1({ S2096 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_259_ (
  .in1({ S2096 }),
  .out1({ S2097 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_579_ (
  .in1({ S1935, DP_LGU1_in1_2 }),
  .out1({ S2098 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_875_ (
  .in1({ S2098, S2436 }),
  .out1({ S2099 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_876_ (
  .in1({ S2099, DP_LGU1_in1_3 }),
  .out1({ S2100 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_580_ (
  .in1({ S2100, S2097 }),
  .out1({ S2101 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_581_ (
  .in1({ S2101, S109 }),
  .out1({ S2102 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_877_ (
  .in1({ S2102, S2093 }),
  .out1({ S2103 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_582_ (
  .in1({ S2408, DP_AC_dout_4 }),
  .out1({ S2104 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_583_ (
  .in1({ S2104, S110 }),
  .out1({ S2105 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_878_ (
  .in1({ S2105, S2103 }),
  .out1({ S2106 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_260_ (
  .in1({ S2106 }),
  .out1({ S2107 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_584_ (
  .in1({ S2107, S2077 }),
  .out1({ DP_LGU1_out_4 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_879_ (
  .in1({ DP_LGU1_in1_5, DP_AC_dout_5 }),
  .out1({ S2108 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_880_ (
  .in1({ S2108, S111 }),
  .out1({ S2109 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_261_ (
  .in1({ S2109 }),
  .out1({ S2110 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_881_ (
  .in1({ S1960, S1956 }),
  .out1({ S2111 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_882_ (
  .in1({ S2111, S2327 }),
  .out1({ S2112 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_883_ (
  .in1({ S2030, DP_LGU1_in1_1 }),
  .out1({ S2113 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_884_ (
  .in1({ S2113, S2112 }),
  .out1({ S2114 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_885_ (
  .in1({ S2114, S1984 }),
  .out1({ S2115 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_262_ (
  .in1({ S2115 }),
  .out1({ S2116 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_585_ (
  .in1({ S2085, S1949 }),
  .out1({ S2117 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_263_ (
  .in1({ S2117 }),
  .out1({ S2118 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_586_ (
  .in1({ S2117, S2116 }),
  .out1({ S2119 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_886_ (
  .in1({ S2118, S2115 }),
  .out1({ S2120 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_887_ (
  .in1({ S1922, DP_LGU1_in1_2 }),
  .out1({ S2121 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_888_ (
  .in1({ S1968, S2380 }),
  .out1({ S2122 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_889_ (
  .in1({ S2122, S2121 }),
  .out1({ S2123 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_587_ (
  .in1({ S2123, DP_LGU1_in1_3 }),
  .out1({ S2124 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_588_ (
  .in1({ S2124, S112 }),
  .out1({ S2125 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_589_ (
  .in1({ S2125, S2120 }),
  .out1({ S2126 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_890_ (
  .in1({ S1930, S2380 }),
  .out1({ S2127 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_891_ (
  .in1({ S2127, S2058 }),
  .out1({ S2128 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_892_ (
  .in1({ S2128, S1909 }),
  .out1({ S2129 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_893_ (
  .in1({ S2098, S1939 }),
  .out1({ S2130 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_894_ (
  .in1({ S2130, DP_LGU1_in1_3 }),
  .out1({ S2131 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_264_ (
  .in1({ S2131 }),
  .out1({ S2132 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_895_ (
  .in1({ S2132, S2129 }),
  .out1({ S2133 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_896_ (
  .in1({ S2133, S2408 }),
  .out1({ S2134 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_590_ (
  .in1({ S2134, S2126 }),
  .out1({ S2135 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_897_ (
  .in1({ S113, S2369 }),
  .out1({ S2136 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_898_ (
  .in1({ S2136, S2409 }),
  .out1({ S2137 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_591_ (
  .in1({ S2137, S2135 }),
  .out1({ S2138 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_592_ (
  .in1({ S2138, S2110 }),
  .out1({ DP_LGU1_out_5 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_899_ (
  .in1({ DP_LGU1_in1_6, DP_AC_dout_6 }),
  .out1({ S2139 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_900_ (
  .in1({ S2139, S114 }),
  .out1({ S2140 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_265_ (
  .in1({ S2140 }),
  .out1({ S2141 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_901_ (
  .in1({ S1887, S1882 }),
  .out1({ S2142 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_902_ (
  .in1({ S2078, DP_LGU1_in1_1 }),
  .out1({ S2143 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_593_ (
  .in1({ S2142, DP_LGU1_in1_1 }),
  .out1({ S2144 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_266_ (
  .in1({ S2144 }),
  .out1({ S2145 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_903_ (
  .in1({ S2145, S2143 }),
  .out1({ S2146 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_594_ (
  .in1({ S2146, S1985 }),
  .out1({ S2147 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_595_ (
  .in1({ S2085, S1990 }),
  .out1({ S2148 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_596_ (
  .in1({ S2148, S2147 }),
  .out1({ S2149 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_597_ (
  .in1({ S2000, DP_LGU1_in1_2 }),
  .out1({ S2150 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_598_ (
  .in1({ S2008, S2380 }),
  .out1({ S2151 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_599_ (
  .in1({ S2151, S2150 }),
  .out1({ S2152 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_600_ (
  .in1({ S2152, DP_LGU1_in1_3 }),
  .out1({ S2153 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_601_ (
  .in1({ S2153, S115 }),
  .out1({ S2154 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_267_ (
  .in1({ S2154 }),
  .out1({ S2155 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_904_ (
  .in1({ S2155, S2149 }),
  .out1({ S2156 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_905_ (
  .in1({ S2012, S2380 }),
  .out1({ S2157 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_906_ (
  .in1({ S2157, S2058 }),
  .out1({ S2158 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_907_ (
  .in1({ S2158, S1909 }),
  .out1({ S2159 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_268_ (
  .in1({ S2159 }),
  .out1({ S2160 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_908_ (
  .in1({ S2098, S2010 }),
  .out1({ S2161 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_909_ (
  .in1({ S2161, DP_LGU1_in1_3 }),
  .out1({ S2162 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_602_ (
  .in1({ S2162, S2160 }),
  .out1({ S2163 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_603_ (
  .in1({ S2163, S116 }),
  .out1({ S2164 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_910_ (
  .in1({ S2164, S2156 }),
  .out1({ S2165 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_604_ (
  .in1({ S2408, DP_AC_dout_6 }),
  .out1({ S2166 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_605_ (
  .in1({ S2166, S117 }),
  .out1({ S2167 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_911_ (
  .in1({ S2167, S2165 }),
  .out1({ S2168 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_269_ (
  .in1({ S2168 }),
  .out1({ S2169 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_606_ (
  .in1({ S2169, S2141 }),
  .out1({ DP_LGU1_out_6 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_912_ (
  .in1({ S118, DP_AC_dout_7 }),
  .out1({ S2170 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_270_ (
  .in1({ S2170 }),
  .out1({ S2171 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_913_ (
  .in1({ S2171, DP_LGU1_in1_7 }),
  .out1({ S2172 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_607_ (
  .in1({ S2045, DP_LGU1_in1_2 }),
  .out1({ S2173 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_914_ (
  .in1({ S2055, DP_LGU1_in1_2 }),
  .out1({ S2174 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_608_ (
  .in1({ S2173, S119 }),
  .out1({ S2175 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_915_ (
  .in1({ S2175, S2174 }),
  .out1({ S2176 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_916_ (
  .in1({ S1964, S1961 }),
  .out1({ S2177 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_271_ (
  .in1({ S2177 }),
  .out1({ S2178 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_609_ (
  .in1({ S2178, DP_LGU1_in1_1 }),
  .out1({ S2179 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_917_ (
  .in1({ S2177, S2327 }),
  .out1({ S2180 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_918_ (
  .in1({ S2111, DP_LGU1_in1_1 }),
  .out1({ S2181 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_272_ (
  .in1({ S2181 }),
  .out1({ S2182 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_610_ (
  .in1({ S2182, S2179 }),
  .out1({ S2183 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_919_ (
  .in1({ S2181, S2180 }),
  .out1({ S2184 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_611_ (
  .in1({ S2183, S1985 }),
  .out1({ S2185 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_920_ (
  .in1({ S2184, S1984 }),
  .out1({ S2186 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_612_ (
  .in1({ S2085, S2035 }),
  .out1({ S2187 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_921_ (
  .in1({ S2084, S2036 }),
  .out1({ S2188 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_613_ (
  .in1({ S2187, S2185 }),
  .out1({ S2189 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_922_ (
  .in1({ S2188, S2186 }),
  .out1({ S2190 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_614_ (
  .in1({ S2190, DP_LGU1_in1_3 }),
  .out1({ S2191 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_923_ (
  .in1({ S2191, S2176 }),
  .out1({ S2192 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_924_ (
  .in1({ S2098, S2063 }),
  .out1({ S2193 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_615_ (
  .in1({ S1910, S2401 }),
  .out1({ S2194 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_616_ (
  .in1({ S2194, S2317 }),
  .out1({ S2195 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_925_ (
  .in1({ S2195, S2193 }),
  .out1({ S2196 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_926_ (
  .in1({ S2196, S2192 }),
  .out1({ S2197 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_927_ (
  .in1({ S2197, S2408 }),
  .out1({ S2198 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_928_ (
  .in1({ S120, DP_AC_dout_7 }),
  .out1({ S2199 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_273_ (
  .in1({ S2199 }),
  .out1({ S2200 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_617_ (
  .in1({ S2200, S121 }),
  .out1({ S2201 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_929_ (
  .in1({ S2201, S2198 }),
  .out1({ S2202 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_930_ (
  .in1({ S2202, S2172 }),
  .out1({ DP_LGU1_out_7 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_931_ (
  .in1({ S1888, S2417 }),
  .out1({ S2203 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_274_ (
  .in1({ S2203 }),
  .out1({ S2204 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_618_ (
  .in1({ S2204, DP_LGU1_in1_1 }),
  .out1({ S2205 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_932_ (
  .in1({ S2142, DP_LGU1_in1_1 }),
  .out1({ S2206 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_275_ (
  .in1({ S2206 }),
  .out1({ S2207 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_619_ (
  .in1({ S2207, S2205 }),
  .out1({ S2208 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_620_ (
  .in1({ S2208, S1985 }),
  .out1({ S2209 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_621_ (
  .in1({ S2085, S2082 }),
  .out1({ S2210 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_622_ (
  .in1({ S2210, S2209 }),
  .out1({ S2211 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_933_ (
  .in1({ S2211, S2439 }),
  .out1({ S2212 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_934_ (
  .in1({ S2212, S2317 }),
  .out1({ S2213 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_623_ (
  .in1({ S1899, S2317 }),
  .out1({ S2214 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_935_ (
  .in1({ S1898, DP_LGU1_in1_3 }),
  .out1({ S2215 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_624_ (
  .in1({ S2215, S1897 }),
  .out1({ S2216 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_936_ (
  .in1({ S2194, DP_LGU1_in1_3 }),
  .out1({ S2217 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_625_ (
  .in1({ S2194, S122 }),
  .out1({ S2218 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_937_ (
  .in1({ S2217, S2408 }),
  .out1({ S2219 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_276_ (
  .in1({ S2219 }),
  .out1({ S2220 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_626_ (
  .in1({ S2219, S2216 }),
  .out1({ S2221 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_938_ (
  .in1({ S2221, S2213 }),
  .out1({ S2222 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_939_ (
  .in1({ S123, DP_AC_dout_8 }),
  .out1({ S2223 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_277_ (
  .in1({ S2223 }),
  .out1({ S2224 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_627_ (
  .in1({ S2224, S124 }),
  .out1({ S2225 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_940_ (
  .in1({ S2225, S2222 }),
  .out1({ S2226 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_941_ (
  .in1({ S125, DP_AC_dout_8 }),
  .out1({ S2227 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_278_ (
  .in1({ S2227 }),
  .out1({ S2228 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_942_ (
  .in1({ S2228, DP_LGU1_in1_8 }),
  .out1({ S2229 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_943_ (
  .in1({ S2229, S2226 }),
  .out1({ DP_LGU1_out_8 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_944_ (
  .in1({ S126, DP_AC_dout_9 }),
  .out1({ S2230 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_628_ (
  .in1({ S2230, S2410 }),
  .out1({ S2231 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_945_ (
  .in1({ S1965, S1911 }),
  .out1({ S2232 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_279_ (
  .in1({ S2232 }),
  .out1({ S2233 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_629_ (
  .in1({ S2233, DP_LGU1_in1_1 }),
  .out1({ S2234 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_946_ (
  .in1({ S2232, S2327 }),
  .out1({ S2235 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_947_ (
  .in1({ S2177, DP_LGU1_in1_1 }),
  .out1({ S2236 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_280_ (
  .in1({ S2236 }),
  .out1({ S2237 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_630_ (
  .in1({ S2237, S2234 }),
  .out1({ S2238 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_948_ (
  .in1({ S2236, S2235 }),
  .out1({ S2239 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_949_ (
  .in1({ S2239, S1984 }),
  .out1({ S2240 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_950_ (
  .in1({ S2114, S2084 }),
  .out1({ S2241 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_951_ (
  .in1({ S2241, S2240 }),
  .out1({ S2242 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_631_ (
  .in1({ S2242, S1943 }),
  .out1({ S2243 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_632_ (
  .in1({ S2243, DP_LGU1_in1_3 }),
  .out1({ S2244 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_952_ (
  .in1({ S2214, S1950 }),
  .out1({ S2245 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_953_ (
  .in1({ S2245, S2220 }),
  .out1({ S2246 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_633_ (
  .in1({ S2246, S2244 }),
  .out1({ S2247 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_954_ (
  .in1({ S127, DP_AC_dout_9 }),
  .out1({ S2248 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_955_ (
  .in1({ S2248, S2409 }),
  .out1({ S2249 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_634_ (
  .in1({ S2249, S2247 }),
  .out1({ S2250 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_635_ (
  .in1({ S2250, S2231 }),
  .out1({ S2251 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_281_ (
  .in1({ S2251 }),
  .out1({ DP_LGU1_out_9 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_956_ (
  .in1({ S1993, DP_LGU1_in1_3 }),
  .out1({ S2252 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_636_ (
  .in1({ S2146, S2085 }),
  .out1({ S2253 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_957_ (
  .in1({ S2421, S2418 }),
  .out1({ S2254 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_958_ (
  .in1({ S2254, S2327 }),
  .out1({ S2255 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_959_ (
  .in1({ S2203, DP_LGU1_in1_1 }),
  .out1({ S2256 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_960_ (
  .in1({ S2256, S2255 }),
  .out1({ S2257 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_961_ (
  .in1({ S2257, S1984 }),
  .out1({ S2258 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_962_ (
  .in1({ S2258, S2215 }),
  .out1({ S2259 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_637_ (
  .in1({ S2259, S2253 }),
  .out1({ S2260 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_963_ (
  .in1({ S2260, S2018 }),
  .out1({ S2261 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_964_ (
  .in1({ S2261, S2252 }),
  .out1({ S2262 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_638_ (
  .in1({ S1910, DP_LGU1_in1_3 }),
  .out1({ S2263 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_639_ (
  .in1({ S2015, DP_LGU1_in1_3 }),
  .out1({ S2264 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_640_ (
  .in1({ S2264, S2219 }),
  .out1({ S2265 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_965_ (
  .in1({ S2265, S2262 }),
  .out1({ S2266 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_966_ (
  .in1({ S128, DP_AC_dout_10 }),
  .out1({ S2267 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_282_ (
  .in1({ S2267 }),
  .out1({ S2268 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_641_ (
  .in1({ S2268, S129 }),
  .out1({ S2269 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_967_ (
  .in1({ S2269, S2266 }),
  .out1({ S2270 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_968_ (
  .in1({ S130, DP_AC_dout_10 }),
  .out1({ S2271 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_283_ (
  .in1({ S2271 }),
  .out1({ S2272 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_969_ (
  .in1({ S2272, DP_LGU1_in1_10 }),
  .out1({ S2273 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_970_ (
  .in1({ S2273, S2270 }),
  .out1({ DP_LGU1_out_10 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_971_ (
  .in1({ S131, DP_AC_dout_11 }),
  .out1({ S2274 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_642_ (
  .in1({ S2274, S2411 }),
  .out1({ S2275 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_972_ (
  .in1({ S2038, DP_LGU1_in1_3 }),
  .out1({ S2276 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_284_ (
  .in1({ S2276 }),
  .out1({ S2277 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_973_ (
  .in1({ S2184, S2084 }),
  .out1({ S2278 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_974_ (
  .in1({ S2278, S2066 }),
  .out1({ S2279 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_643_ (
  .in1({ S2279, S2214 }),
  .out1({ S2280 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_644_ (
  .in1({ S2280, S2277 }),
  .out1({ S2281 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_645_ (
  .in1({ S1916, S1913 }),
  .out1({ S2282 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_646_ (
  .in1({ S2282, DP_LGU1_in1_1 }),
  .out1({ S2283 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_285_ (
  .in1({ S2283 }),
  .out1({ S2284 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_975_ (
  .in1({ S2232, DP_LGU1_in1_1 }),
  .out1({ S2285 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_976_ (
  .in1({ S2285, S2284 }),
  .out1({ S2286 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_977_ (
  .in1({ S2286, S1984 }),
  .out1({ S2287 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_978_ (
  .in1({ S2287, S2062 }),
  .out1({ S2288 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_979_ (
  .in1({ S2288, S2317 }),
  .out1({ S2289 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_980_ (
  .in1({ S2289, S2220 }),
  .out1({ S2290 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_647_ (
  .in1({ S2290, S2281 }),
  .out1({ S2291 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_981_ (
  .in1({ S132, DP_AC_dout_11 }),
  .out1({ S2292 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_982_ (
  .in1({ S2292, S2409 }),
  .out1({ S2293 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_648_ (
  .in1({ S2293, S2291 }),
  .out1({ S2294 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_649_ (
  .in1({ S2294, S2275 }),
  .out1({ S2295 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_286_ (
  .in1({ S2295 }),
  .out1({ DP_LGU1_out_11 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_983_ (
  .in1({ S2087, DP_LGU1_in1_3 }),
  .out1({ S2296 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_650_ (
  .in1({ S2208, S2085 }),
  .out1({ S2297 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_984_ (
  .in1({ S2254, DP_LGU1_in1_1 }),
  .out1({ S2298 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_985_ (
  .in1({ S2427, S2422 }),
  .out1({ S2299 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_287_ (
  .in1({ S2299 }),
  .out1({ S2300 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_986_ (
  .in1({ S2299, S2327 }),
  .out1({ S2301 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_987_ (
  .in1({ S2301, S2298 }),
  .out1({ S2302 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_988_ (
  .in1({ S2302, S1984 }),
  .out1({ S2303 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_989_ (
  .in1({ S2303, S2215 }),
  .out1({ S2304 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_651_ (
  .in1({ S2304, S2297 }),
  .out1({ S2305 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_990_ (
  .in1({ S2305, S2099 }),
  .out1({ S2307 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_991_ (
  .in1({ S2307, S2296 }),
  .out1({ S2308 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_652_ (
  .in1({ S2096, DP_LGU1_in1_3 }),
  .out1({ S2309 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_653_ (
  .in1({ S2309, S2219 }),
  .out1({ S2310 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_992_ (
  .in1({ S2310, S2308 }),
  .out1({ S2311 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_993_ (
  .in1({ S133, DP_AC_dout_12 }),
  .out1({ S2312 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_288_ (
  .in1({ S2312 }),
  .out1({ S2313 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_654_ (
  .in1({ S2313, S134 }),
  .out1({ S2314 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_994_ (
  .in1({ S2314, S2311 }),
  .out1({ S2315 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_995_ (
  .in1({ S135, DP_AC_dout_12 }),
  .out1({ S2316 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_289_ (
  .in1({ S2316 }),
  .out1({ S2318 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_996_ (
  .in1({ S2318, DP_LGU1_in1_12 }),
  .out1({ S2319 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_997_ (
  .in1({ S2319, S2315 }),
  .out1({ DP_LGU1_out_12 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_998_ (
  .in1({ S136, DP_AC_dout_13 }),
  .out1({ S2320 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_290_ (
  .in1({ S2320 }),
  .out1({ S2321 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_999_ (
  .in1({ S2321, DP_LGU1_in1_13 }),
  .out1({ S2322 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_655_ (
  .in1({ S2128, DP_LGU1_in1_3 }),
  .out1({ S2323 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_656_ (
  .in1({ S2263, S2194 }),
  .out1({ S2324 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_657_ (
  .in1({ S2324, S2323 }),
  .out1({ S2325 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1000_ (
  .in1({ S2119, DP_LGU1_in1_3 }),
  .out1({ S2326 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1001_ (
  .in1({ S2215, S2130 }),
  .out1({ S2328 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1002_ (
  .in1({ S1924, S1918 }),
  .out1({ S2329 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1003_ (
  .in1({ S2282, DP_LGU1_in1_1 }),
  .out1({ S2330 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_658_ (
  .in1({ S2329, DP_LGU1_in1_1 }),
  .out1({ S2331 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_659_ (
  .in1({ S2331, S1985 }),
  .out1({ S2332 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1004_ (
  .in1({ S2332, S2330 }),
  .out1({ S2333 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_660_ (
  .in1({ S2238, S2085 }),
  .out1({ S2334 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_661_ (
  .in1({ S2334, S2328 }),
  .out1({ S2335 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1005_ (
  .in1({ S2335, S2333 }),
  .out1({ S2336 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1006_ (
  .in1({ S2336, S2326 }),
  .out1({ S2337 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_662_ (
  .in1({ S2325, S137 }),
  .out1({ S2339 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1007_ (
  .in1({ S2339, S2337 }),
  .out1({ S2340 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1008_ (
  .in1({ S138, DP_AC_dout_13 }),
  .out1({ S2341 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_291_ (
  .in1({ S2341 }),
  .out1({ S2342 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_663_ (
  .in1({ S2342, S139 }),
  .out1({ S2343 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1009_ (
  .in1({ S2343, S2340 }),
  .out1({ S2344 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1010_ (
  .in1({ S2344, S2322 }),
  .out1({ DP_LGU1_out_13 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1011_ (
  .in1({ S140, DP_AC_dout_14 }),
  .out1({ S2345 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_292_ (
  .in1({ S2345 }),
  .out1({ S2346 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1012_ (
  .in1({ S2346, DP_LGU1_in1_14 }),
  .out1({ S2347 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_664_ (
  .in1({ S2158, DP_LGU1_in1_3 }),
  .out1({ S2349 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_665_ (
  .in1({ S2349, S2324 }),
  .out1({ S2350 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1013_ (
  .in1({ S2149, DP_LGU1_in1_3 }),
  .out1({ S2351 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1014_ (
  .in1({ S2257, S2084 }),
  .out1({ S2352 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1015_ (
  .in1({ S2431, S2428 }),
  .out1({ S2353 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_666_ (
  .in1({ S2353, DP_LGU1_in1_1 }),
  .out1({ S2354 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1016_ (
  .in1({ S2300, DP_LGU1_in1_1 }),
  .out1({ S2355 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1017_ (
  .in1({ S2355, S1984 }),
  .out1({ S2356 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_667_ (
  .in1({ S2356, S2354 }),
  .out1({ S2357 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1018_ (
  .in1({ S2352, S2161 }),
  .out1({ S2358 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_668_ (
  .in1({ S2358, S2357 }),
  .out1({ S2360 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1019_ (
  .in1({ S2360, S2215 }),
  .out1({ S2361 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1020_ (
  .in1({ S2361, S2351 }),
  .out1({ S2362 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_669_ (
  .in1({ S2350, S141 }),
  .out1({ S2363 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1021_ (
  .in1({ S2363, S2362 }),
  .out1({ S2364 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1022_ (
  .in1({ S142, DP_AC_dout_14 }),
  .out1({ S2365 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_293_ (
  .in1({ S2365 }),
  .out1({ S2366 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_670_ (
  .in1({ S2366, S143 }),
  .out1({ S2367 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1023_ (
  .in1({ S2367, S2364 }),
  .out1({ S2368 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1024_ (
  .in1({ S2368, S2347 }),
  .out1({ DP_LGU1_out_14 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1025_ (
  .in1({ S2189, DP_LGU1_in1_3 }),
  .out1({ S2370 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1026_ (
  .in1({ S2286, S2084 }),
  .out1({ S2371 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_671_ (
  .in1({ S1936, S1926 }),
  .out1({ S2372 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_672_ (
  .in1({ S2329, S2327 }),
  .out1({ S2373 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1027_ (
  .in1({ S2372, S2327 }),
  .out1({ S2374 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1028_ (
  .in1({ S2374, S1984 }),
  .out1({ S2375 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_673_ (
  .in1({ S2375, S2373 }),
  .out1({ S2376 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1029_ (
  .in1({ S2215, S2193 }),
  .out1({ S2377 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_674_ (
  .in1({ S2377, S2376 }),
  .out1({ S2378 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1030_ (
  .in1({ S2378, S2371 }),
  .out1({ S2379 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1031_ (
  .in1({ S2379, S2370 }),
  .out1({ S2381 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1032_ (
  .in1({ S2381, S2218 }),
  .out1({ S2382 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1033_ (
  .in1({ S144, DP_AC_dout_15 }),
  .out1({ S2383 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_294_ (
  .in1({ S2383 }),
  .out1({ S2384 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_675_ (
  .in1({ S2384, S145 }),
  .out1({ S2385 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1034_ (
  .in1({ S2385, S2382 }),
  .out1({ S2386 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1035_ (
  .in1({ S146, DP_AC_dout_15 }),
  .out1({ S2387 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_295_ (
  .in1({ S2387 }),
  .out1({ S2388 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1036_ (
  .in1({ S2388, DP_LGU1_in1_15 }),
  .out1({ S2389 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1037_ (
  .in1({ S2389, S2386 }),
  .out1({ DP_LGU1_N })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1038_ (
  .in1({ S2074, S2027 }),
  .out1({ S2391 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1039_ (
  .in1({ S2295, S2251 }),
  .out1({ S2392 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_676_ (
  .in1({ S2392, S2391 }),
  .out1({ S2393 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_677_ (
  .in1({ DP_LGU1_out_7, DP_LGU1_out_6 }),
  .out1({ S2394 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_678_ (
  .in1({ DP_LGU1_N, DP_LGU1_out_4 }),
  .out1({ S2395 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1040_ (
  .in1({ S2395, S2394 }),
  .out1({ S2396 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_679_ (
  .in1({ DP_LGU1_out_13, DP_LGU1_out_12 }),
  .out1({ S2397 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_680_ (
  .in1({ DP_LGU1_out_14, DP_LGU1_out_10 }),
  .out1({ S2398 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1041_ (
  .in1({ S2398, S2397 }),
  .out1({ S2399 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_681_ (
  .in1({ DP_LGU1_out_8, DP_LGU1_out_5 }),
  .out1({ S2400 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_682_ (
  .in1({ DP_LGU1_out_1, DP_LGU1_out_0 }),
  .out1({ S2402 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1042_ (
  .in1({ S2402, S2400 }),
  .out1({ S2403 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_683_ (
  .in1({ S2403, S2399 }),
  .out1({ S2404 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1043_ (
  .in1({ S2404, S2393 }),
  .out1({ S2405 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_684_ (
  .in1({ S2405, S2396 }),
  .out1({ DP_LGU1_Z })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_296_ (
  .in1({ S147 }),
  .out1({ S2446 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_685_ (
  .in1({ S149, S148 }),
  .out1({ S2447 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1044_ (
  .in1({ S2447, DP_IMM1_in1_0 }),
  .out1({ S2448 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_686_ (
  .in1({ S2446, S150 }),
  .out1({ S2449 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1045_ (
  .in1({ S2449, DP_OF_din_0 }),
  .out1({ S2450 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1046_ (
  .in1({ S2450, S2448 }),
  .out1({ S2442 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1047_ (
  .in1({ S2447, DP_IMM1_in1_1 }),
  .out1({ S2451 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1048_ (
  .in1({ S2449, DP_OF_din_1 }),
  .out1({ S2452 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1049_ (
  .in1({ S2452, S2451 }),
  .out1({ S2443 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1050_ (
  .in1({ S2447, DP_IMM1_in1_2 }),
  .out1({ S2453 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1051_ (
  .in1({ S2449, DP_OF_din_2 }),
  .out1({ S2454 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1052_ (
  .in1({ S2454, S2453 }),
  .out1({ S2444 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1053_ (
  .in1({ S2447, DP_IMM1_in1_3 }),
  .out1({ S2455 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1054_ (
  .in1({ S2449, DP_OF_din_3 }),
  .out1({ S2456 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1055_ (
  .in1({ S2456, S2455 }),
  .out1({ S2445 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_49_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2442 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IMM1_in1_0 }),
  .Si({ S3408 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_50_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2443 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IMM1_in1_1 }),
  .Si({ S3407 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_51_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2444 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IMM1_in1_2 }),
  .Si({ S3406 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_52_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2445 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_IMM1_in1_3 }),
  .Si({ S3427 }),
  .global_reset({ 1'b0 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_297_ (
  .in1({ S151 }),
  .out1({ S2474 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_687_ (
  .in1({ S153, S152 }),
  .out1({ S2475 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1056_ (
  .in1({ S2475, DP_INC_1_in_0 }),
  .out1({ S2476 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_688_ (
  .in1({ S2474, S154 }),
  .out1({ S2477 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1057_ (
  .in1({ S2477, DP_PC_din_0 }),
  .out1({ S2478 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1058_ (
  .in1({ S2478, S2476 }),
  .out1({ S2457 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1059_ (
  .in1({ S2475, DP_INC_1_in_1 }),
  .out1({ S2479 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1060_ (
  .in1({ S2477, DP_PC_din_1 }),
  .out1({ S2480 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1061_ (
  .in1({ S2480, S2479 }),
  .out1({ S2458 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1062_ (
  .in1({ S2475, DP_INC_1_in_2 }),
  .out1({ S2481 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1063_ (
  .in1({ S2477, DP_PC_din_2 }),
  .out1({ S2482 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1064_ (
  .in1({ S2482, S2481 }),
  .out1({ S2459 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1065_ (
  .in1({ S2475, DP_INC_1_in_3 }),
  .out1({ S2483 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1066_ (
  .in1({ S2477, DP_PC_din_3 }),
  .out1({ S2484 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1067_ (
  .in1({ S2484, S2483 }),
  .out1({ S2460 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1068_ (
  .in1({ S2475, DP_INC_1_in_4 }),
  .out1({ S2485 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1069_ (
  .in1({ S2477, DP_PC_din_4 }),
  .out1({ S2486 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1070_ (
  .in1({ S2486, S2485 }),
  .out1({ S2461 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1071_ (
  .in1({ S2475, DP_INC_1_in_5 }),
  .out1({ S2487 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1072_ (
  .in1({ S2477, DP_PC_din_5 }),
  .out1({ S2488 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1073_ (
  .in1({ S2488, S2487 }),
  .out1({ S2462 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1074_ (
  .in1({ S2475, DP_INC_1_in_6 }),
  .out1({ S2489 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1075_ (
  .in1({ S2477, DP_PC_din_6 }),
  .out1({ S2490 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1076_ (
  .in1({ S2490, S2489 }),
  .out1({ S2463 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1077_ (
  .in1({ S2475, DP_INC_1_in_7 }),
  .out1({ S2491 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1078_ (
  .in1({ S2477, DP_PC_din_7 }),
  .out1({ S2492 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1079_ (
  .in1({ S2492, S2491 }),
  .out1({ S2464 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1080_ (
  .in1({ S2475, DP_INC_1_in_8 }),
  .out1({ S2493 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1081_ (
  .in1({ S2477, DP_PC_din_8 }),
  .out1({ S2494 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1082_ (
  .in1({ S2494, S2493 }),
  .out1({ S2465 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1083_ (
  .in1({ S2475, DP_INC_1_in_9 }),
  .out1({ S2495 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1084_ (
  .in1({ S2477, DP_PC_din_9 }),
  .out1({ S2496 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1085_ (
  .in1({ S2496, S2495 }),
  .out1({ S2466 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1086_ (
  .in1({ S2475, DP_INC_1_in_10 }),
  .out1({ S2497 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1087_ (
  .in1({ S2477, DP_PC_din_10 }),
  .out1({ S2498 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1088_ (
  .in1({ S2498, S2497 }),
  .out1({ S2467 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1089_ (
  .in1({ S2475, DP_INC_1_in_11 }),
  .out1({ S2499 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1090_ (
  .in1({ S2477, DP_PC_din_11 }),
  .out1({ S2500 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1091_ (
  .in1({ S2500, S2499 }),
  .out1({ S2468 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1092_ (
  .in1({ S2475, DP_INC_1_in_12 }),
  .out1({ S2501 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1093_ (
  .in1({ S2477, DP_PC_din_12 }),
  .out1({ S2502 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1094_ (
  .in1({ S2502, S2501 }),
  .out1({ S2469 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1095_ (
  .in1({ S2475, DP_INC_1_in_13 }),
  .out1({ S2503 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1096_ (
  .in1({ S2477, DP_PC_din_13 }),
  .out1({ S2504 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1097_ (
  .in1({ S2504, S2503 }),
  .out1({ S2470 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1098_ (
  .in1({ S2475, DP_INC_1_in_14 }),
  .out1({ S2505 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1099_ (
  .in1({ S2477, DP_PC_din_14 }),
  .out1({ S2506 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1100_ (
  .in1({ S2506, S2505 }),
  .out1({ S2471 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1101_ (
  .in1({ S2475, DP_INC_1_in_15 }),
  .out1({ S2507 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1102_ (
  .in1({ S2477, DP_PC_din_15 }),
  .out1({ S2473 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1103_ (
  .in1({ S2473, S2507 }),
  .out1({ S2472 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_53_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2457 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_0 }),
  .Si({ S3423 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_54_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2458 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_1 }),
  .Si({ S3422 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_55_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2459 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_2 }),
  .Si({ S3421 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_56_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2460 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_3 }),
  .Si({ S3420 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_57_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2461 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_4 }),
  .Si({ S3419 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_58_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2462 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_5 }),
  .Si({ S3418 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_59_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2463 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_6 }),
  .Si({ S3417 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_60_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2464 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_7 }),
  .Si({ S3416 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_61_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2465 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_8 }),
  .Si({ S3415 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_62_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2466 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_9 }),
  .Si({ S3414 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_63_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2467 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_10 }),
  .Si({ S3413 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_64_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2468 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_11 }),
  .Si({ S3412 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_65_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2469 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_12 }),
  .Si({ S3411 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_66_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2470 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_13 }),
  .Si({ S3410 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_67_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2471 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_14 }),
  .Si({ S3409 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_68_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2472 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_INC_1_in_15 }),
  .Si({ S3428 }),
  .global_reset({ 1'b0 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_298_ (
  .in1({ DP_SR_C_dout }),
  .out1({ S2510 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1104_ (
  .in1({ DP_SR_C_din, S155 }),
  .out1({ S2511 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_299_ (
  .in1({ S2511 }),
  .out1({ S2512 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_689_ (
  .in1({ S2510, S156 }),
  .out1({ S2513 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_690_ (
  .in1({ S2513, S2512 }),
  .out1({ S2509 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_691_ (
  .in1({ S2509, S157 }),
  .out1({ S2508 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_69_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2508 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_SR_C_dout }),
  .Si({ S3429 }),
  .global_reset({ 1'b0 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_300_ (
  .in1({ DP_SR_N_dout }),
  .out1({ S2516 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1105_ (
  .in1({ DP_SR_N_din, S158 }),
  .out1({ S2517 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_301_ (
  .in1({ S2517 }),
  .out1({ S2518 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_692_ (
  .in1({ S2516, S159 }),
  .out1({ S2519 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_693_ (
  .in1({ S2519, S2518 }),
  .out1({ S2515 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_694_ (
  .in1({ S2515, S160 }),
  .out1({ S2514 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_70_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2514 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_SR_N_dout }),
  .Si({ S3430 }),
  .global_reset({ 1'b0 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_302_ (
  .in1({ DP_SR_V_dout }),
  .out1({ S2522 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1106_ (
  .in1({ DP_SR_V_din, S161 }),
  .out1({ S2523 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_303_ (
  .in1({ S2523 }),
  .out1({ S2524 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_695_ (
  .in1({ S2522, S162 }),
  .out1({ S2525 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_696_ (
  .in1({ S2525, S2524 }),
  .out1({ S2521 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_697_ (
  .in1({ S2521, S163 }),
  .out1({ S2520 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_71_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2520 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_SR_V_dout }),
  .Si({ S3431 }),
  .global_reset({ 1'b0 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_304_ (
  .in1({ DP_SR_Z_dout }),
  .out1({ S2528 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1107_ (
  .in1({ DP_SR_Z_din, S164 }),
  .out1({ S2529 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_305_ (
  .in1({ S2529 }),
  .out1({ S2530 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_698_ (
  .in1({ S2528, S165 }),
  .out1({ S2531 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_699_ (
  .in1({ S2531, S2530 }),
  .out1({ S2527 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_700_ (
  .in1({ S2527, S166 }),
  .out1({ S2526 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_72_ (
  .C({ CU_clk }),
  .CE({ 1'b1 }),
  .CLR({ CU_rst }),
  .D({ S2526 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ DP_SR_Z_dout }),
  .Si({ S3432 }),
  .global_reset({ 1'b0 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1108_ (
  .in1({ DP_TriBuff_in_0, S5 }),
  .out1({ S2532 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_306_ (
  .in1({ S2532 }),
  .out1({ DP_TriBuff_out_0 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1109_ (
  .in1({ DP_TriBuff_in_1, S6 }),
  .out1({ S2533 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_307_ (
  .in1({ S2533 }),
  .out1({ DP_TriBuff_out_1 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1110_ (
  .in1({ DP_TriBuff_in_2, S7 }),
  .out1({ S2534 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_308_ (
  .in1({ S2534 }),
  .out1({ DP_TriBuff_out_2 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1111_ (
  .in1({ DP_TriBuff_in_3, S8 }),
  .out1({ S2535 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_309_ (
  .in1({ S2535 }),
  .out1({ DP_TriBuff_out_3 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1112_ (
  .in1({ DP_TriBuff_in_4, S9 }),
  .out1({ S2536 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_310_ (
  .in1({ S2536 }),
  .out1({ DP_TriBuff_out_4 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1113_ (
  .in1({ DP_TriBuff_in_5, S10 }),
  .out1({ S2537 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_311_ (
  .in1({ S2537 }),
  .out1({ DP_TriBuff_out_5 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1114_ (
  .in1({ DP_TriBuff_in_6, S11 }),
  .out1({ S2538 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_312_ (
  .in1({ S2538 }),
  .out1({ DP_TriBuff_out_6 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1115_ (
  .in1({ DP_TriBuff_in_7, S12 }),
  .out1({ S2539 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_313_ (
  .in1({ S2539 }),
  .out1({ DP_TriBuff_out_7 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1116_ (
  .in1({ DP_TriBuff_in_8, S13 }),
  .out1({ S2540 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_314_ (
  .in1({ S2540 }),
  .out1({ DP_TriBuff_out_8 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1117_ (
  .in1({ DP_TriBuff_in_9, S14 }),
  .out1({ S2541 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_315_ (
  .in1({ S2541 }),
  .out1({ DP_TriBuff_out_9 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1118_ (
  .in1({ DP_TriBuff_in_10, S15 }),
  .out1({ S2542 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_316_ (
  .in1({ S2542 }),
  .out1({ DP_TriBuff_out_10 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1119_ (
  .in1({ DP_TriBuff_in_11, S16 }),
  .out1({ S2543 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_317_ (
  .in1({ S2543 }),
  .out1({ DP_TriBuff_out_11 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1120_ (
  .in1({ DP_TriBuff_in_12, S17 }),
  .out1({ S2544 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_318_ (
  .in1({ S2544 }),
  .out1({ DP_TriBuff_out_12 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1121_ (
  .in1({ DP_TriBuff_in_13, S18 }),
  .out1({ S2545 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_319_ (
  .in1({ S2545 }),
  .out1({ DP_TriBuff_out_13 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1122_ (
  .in1({ DP_TriBuff_in_14, S19 }),
  .out1({ S2546 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_320_ (
  .in1({ S2546 }),
  .out1({ DP_TriBuff_out_14 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1123_ (
  .in1({ DP_TriBuff_in_15, S20 }),
  .out1({ S2547 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_321_ (
  .in1({ S2547 }),
  .out1({ DP_TriBuff_out_15 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_322_ (
  .in1({ DP_LGU1_out_0 }),
  .out1({ S2696 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_323_ (
  .in1({ S167 }),
  .out1({ S2697 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_324_ (
  .in1({ S168 }),
  .out1({ S2698 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_325_ (
  .in1({ DP_LGU1_out_1 }),
  .out1({ S2699 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_326_ (
  .in1({ DP_LGU1_out_2 }),
  .out1({ S2700 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_327_ (
  .in1({ DP_LGU1_out_3 }),
  .out1({ S2701 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_328_ (
  .in1({ DP_LGU1_out_4 }),
  .out1({ S2702 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_329_ (
  .in1({ DP_LGU1_out_5 }),
  .out1({ S2703 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_330_ (
  .in1({ DP_LGU1_out_6 }),
  .out1({ S2704 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_331_ (
  .in1({ DP_LGU1_out_7 }),
  .out1({ S2705 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_332_ (
  .in1({ DP_LGU1_out_8 }),
  .out1({ S2706 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_333_ (
  .in1({ DP_LGU1_out_9 }),
  .out1({ S2707 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_334_ (
  .in1({ DP_LGU1_out_10 }),
  .out1({ S2708 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_335_ (
  .in1({ DP_LGU1_out_11 }),
  .out1({ S2709 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_336_ (
  .in1({ DP_LGU1_out_12 }),
  .out1({ S2710 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_337_ (
  .in1({ DP_LGU1_out_13 }),
  .out1({ S2548 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_338_ (
  .in1({ DP_LGU1_out_14 }),
  .out1({ S2549 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_339_ (
  .in1({ DP_LGU1_N }),
  .out1({ S2550 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_701_ (
  .in1({ S2698, DP_IMM1_out_0 }),
  .out1({ S2551 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1124_ (
  .in1({ S2697, S169 }),
  .out1({ S2552 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_702_ (
  .in1({ S2552, S2696 }),
  .out1({ S2553 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1125_ (
  .in1({ S170, DP_ARU1_out_0 }),
  .out1({ S2554 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_340_ (
  .in1({ S2554 }),
  .out1({ S2555 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_703_ (
  .in1({ S2555, S2553 }),
  .out1({ S2556 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_704_ (
  .in1({ S2556, S171 }),
  .out1({ S2557 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1126_ (
  .in1({ S172, DP_INC_2_in_0 }),
  .out1({ S2558 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1127_ (
  .in1({ S2558, S2698 }),
  .out1({ S2559 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_705_ (
  .in1({ S2559, S2557 }),
  .out1({ S2560 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_706_ (
  .in1({ S2560, S2551 }),
  .out1({ DP_AC_din_0 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_707_ (
  .in1({ DP_IMM1_out_1, S2698 }),
  .out1({ S2561 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_708_ (
  .in1({ S2552, S2699 }),
  .out1({ S2562 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1128_ (
  .in1({ DP_ARU1_out_1, S173 }),
  .out1({ S2563 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_341_ (
  .in1({ S2563 }),
  .out1({ S2564 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_709_ (
  .in1({ S2564, S2562 }),
  .out1({ S2565 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_710_ (
  .in1({ S2565, S174 }),
  .out1({ S2566 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1129_ (
  .in1({ DP_INC_2_in_1, S175 }),
  .out1({ S2567 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1130_ (
  .in1({ S2567, S2698 }),
  .out1({ S2568 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_711_ (
  .in1({ S2568, S2566 }),
  .out1({ S2569 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_712_ (
  .in1({ S2569, S2561 }),
  .out1({ DP_AC_din_1 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_713_ (
  .in1({ DP_IMM1_out_2, S2698 }),
  .out1({ S2570 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_714_ (
  .in1({ S2552, S2700 }),
  .out1({ S2571 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1131_ (
  .in1({ DP_ARU1_out_2, S176 }),
  .out1({ S2572 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_342_ (
  .in1({ S2572 }),
  .out1({ S2573 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_715_ (
  .in1({ S2573, S2571 }),
  .out1({ S2574 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_716_ (
  .in1({ S2574, S177 }),
  .out1({ S2575 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1132_ (
  .in1({ DP_INC_2_in_2, S178 }),
  .out1({ S2576 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1133_ (
  .in1({ S2576, S2698 }),
  .out1({ S2577 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_717_ (
  .in1({ S2577, S2575 }),
  .out1({ S2578 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_718_ (
  .in1({ S2578, S2570 }),
  .out1({ DP_AC_din_2 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_719_ (
  .in1({ DP_IMM1_out_3, S2698 }),
  .out1({ S2579 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_720_ (
  .in1({ S2552, S2701 }),
  .out1({ S2580 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1134_ (
  .in1({ DP_ARU1_out_3, S179 }),
  .out1({ S2581 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_343_ (
  .in1({ S2581 }),
  .out1({ S2582 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_721_ (
  .in1({ S2582, S2580 }),
  .out1({ S2583 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_722_ (
  .in1({ S2583, S180 }),
  .out1({ S2584 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1135_ (
  .in1({ DP_INC_2_in_3, S181 }),
  .out1({ S2585 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1136_ (
  .in1({ S2585, S2698 }),
  .out1({ S2586 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_723_ (
  .in1({ S2586, S2584 }),
  .out1({ S2587 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_724_ (
  .in1({ S2587, S2579 }),
  .out1({ DP_AC_din_3 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_725_ (
  .in1({ DP_IMM1_out_4, S2698 }),
  .out1({ S2588 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_726_ (
  .in1({ S2552, S2702 }),
  .out1({ S2589 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1137_ (
  .in1({ DP_ARU1_out_4, S182 }),
  .out1({ S2590 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_344_ (
  .in1({ S2590 }),
  .out1({ S2591 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_727_ (
  .in1({ S2591, S2589 }),
  .out1({ S2592 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_728_ (
  .in1({ S2592, S183 }),
  .out1({ S2593 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1138_ (
  .in1({ DP_INC_2_in_4, S184 }),
  .out1({ S2594 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1139_ (
  .in1({ S2594, S2698 }),
  .out1({ S2595 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_729_ (
  .in1({ S2595, S2593 }),
  .out1({ S2596 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_730_ (
  .in1({ S2596, S2588 }),
  .out1({ DP_AC_din_4 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_731_ (
  .in1({ DP_IMM1_out_5, S2698 }),
  .out1({ S2597 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_732_ (
  .in1({ S2552, S2703 }),
  .out1({ S2598 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1140_ (
  .in1({ DP_ARU1_out_5, S185 }),
  .out1({ S2599 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_345_ (
  .in1({ S2599 }),
  .out1({ S2600 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_733_ (
  .in1({ S2600, S2598 }),
  .out1({ S2601 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_734_ (
  .in1({ S2601, S186 }),
  .out1({ S2602 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1141_ (
  .in1({ DP_INC_2_in_5, S187 }),
  .out1({ S2603 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1142_ (
  .in1({ S2603, S2698 }),
  .out1({ S2604 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_735_ (
  .in1({ S2604, S2602 }),
  .out1({ S2605 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_736_ (
  .in1({ S2605, S2597 }),
  .out1({ DP_AC_din_5 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_737_ (
  .in1({ DP_IMM1_out_6, S2698 }),
  .out1({ S2606 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_738_ (
  .in1({ S2552, S2704 }),
  .out1({ S2607 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1143_ (
  .in1({ DP_ARU1_out_6, S188 }),
  .out1({ S2608 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_346_ (
  .in1({ S2608 }),
  .out1({ S2609 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_739_ (
  .in1({ S2609, S2607 }),
  .out1({ S2610 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_740_ (
  .in1({ S2610, S189 }),
  .out1({ S2611 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1144_ (
  .in1({ DP_INC_2_in_6, S190 }),
  .out1({ S2612 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1145_ (
  .in1({ S2612, S2698 }),
  .out1({ S2613 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_741_ (
  .in1({ S2613, S2611 }),
  .out1({ S2614 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_742_ (
  .in1({ S2614, S2606 }),
  .out1({ DP_AC_din_6 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_743_ (
  .in1({ DP_IMM1_out_7, S2698 }),
  .out1({ S2615 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_744_ (
  .in1({ S2552, S2705 }),
  .out1({ S2616 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1146_ (
  .in1({ DP_ARU1_out_7, S191 }),
  .out1({ S2617 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_347_ (
  .in1({ S2617 }),
  .out1({ S2618 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_745_ (
  .in1({ S2618, S2616 }),
  .out1({ S2619 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_746_ (
  .in1({ S2619, S192 }),
  .out1({ S2620 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1147_ (
  .in1({ DP_INC_2_in_7, S193 }),
  .out1({ S2621 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1148_ (
  .in1({ S2621, S2698 }),
  .out1({ S2622 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_747_ (
  .in1({ S2622, S2620 }),
  .out1({ S2623 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_748_ (
  .in1({ S2623, S2615 }),
  .out1({ DP_AC_din_7 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_749_ (
  .in1({ DP_IMM1_out_8, S2698 }),
  .out1({ S2624 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_750_ (
  .in1({ S2552, S2706 }),
  .out1({ S2625 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1149_ (
  .in1({ DP_ARU1_out_8, S194 }),
  .out1({ S2626 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_348_ (
  .in1({ S2626 }),
  .out1({ S2627 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_751_ (
  .in1({ S2627, S2625 }),
  .out1({ S2628 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_752_ (
  .in1({ S2628, S195 }),
  .out1({ S2629 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1150_ (
  .in1({ DP_INC_2_in_8, S196 }),
  .out1({ S2630 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1151_ (
  .in1({ S2630, S2698 }),
  .out1({ S2631 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_753_ (
  .in1({ S2631, S2629 }),
  .out1({ S2632 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_754_ (
  .in1({ S2632, S2624 }),
  .out1({ DP_AC_din_8 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_755_ (
  .in1({ DP_IMM1_out_9, S2698 }),
  .out1({ S2633 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_756_ (
  .in1({ S2552, S2707 }),
  .out1({ S2634 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1152_ (
  .in1({ DP_ARU1_out_9, S197 }),
  .out1({ S2635 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_349_ (
  .in1({ S2635 }),
  .out1({ S2636 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_757_ (
  .in1({ S2636, S2634 }),
  .out1({ S2637 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_758_ (
  .in1({ S2637, S198 }),
  .out1({ S2638 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1153_ (
  .in1({ DP_INC_2_in_9, S199 }),
  .out1({ S2639 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1154_ (
  .in1({ S2639, S2698 }),
  .out1({ S2640 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_759_ (
  .in1({ S2640, S2638 }),
  .out1({ S2641 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_760_ (
  .in1({ S2641, S2633 }),
  .out1({ DP_AC_din_9 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_761_ (
  .in1({ DP_IMM1_out_10, S2698 }),
  .out1({ S2642 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_762_ (
  .in1({ S2552, S2708 }),
  .out1({ S2643 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1155_ (
  .in1({ DP_ARU1_out_10, S200 }),
  .out1({ S2644 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_350_ (
  .in1({ S2644 }),
  .out1({ S2645 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_763_ (
  .in1({ S2645, S2643 }),
  .out1({ S2646 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_764_ (
  .in1({ S2646, S201 }),
  .out1({ S2647 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1156_ (
  .in1({ DP_INC_2_in_10, S202 }),
  .out1({ S2648 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1157_ (
  .in1({ S2648, S2698 }),
  .out1({ S2649 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_765_ (
  .in1({ S2649, S2647 }),
  .out1({ S2650 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_766_ (
  .in1({ S2650, S2642 }),
  .out1({ DP_AC_din_10 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_767_ (
  .in1({ DP_IMM1_out_11, S2698 }),
  .out1({ S2651 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_768_ (
  .in1({ S2552, S2709 }),
  .out1({ S2652 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1158_ (
  .in1({ DP_ARU1_out_11, S203 }),
  .out1({ S2653 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_351_ (
  .in1({ S2653 }),
  .out1({ S2654 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_769_ (
  .in1({ S2654, S2652 }),
  .out1({ S2655 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_770_ (
  .in1({ S2655, S204 }),
  .out1({ S2656 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1159_ (
  .in1({ DP_INC_2_in_11, S205 }),
  .out1({ S2657 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1160_ (
  .in1({ S2657, S2698 }),
  .out1({ S2658 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_771_ (
  .in1({ S2658, S2656 }),
  .out1({ S2659 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_772_ (
  .in1({ S2659, S2651 }),
  .out1({ DP_AC_din_11 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_773_ (
  .in1({ DP_IMM1_out_12, S2698 }),
  .out1({ S2660 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_774_ (
  .in1({ S2552, S2710 }),
  .out1({ S2661 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1161_ (
  .in1({ DP_ARU1_out_12, S206 }),
  .out1({ S2662 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_352_ (
  .in1({ S2662 }),
  .out1({ S2663 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_775_ (
  .in1({ S2663, S2661 }),
  .out1({ S2664 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_776_ (
  .in1({ S2664, S207 }),
  .out1({ S2665 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1162_ (
  .in1({ DP_INC_2_in_12, S208 }),
  .out1({ S2666 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1163_ (
  .in1({ S2666, S2698 }),
  .out1({ S2667 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_777_ (
  .in1({ S2667, S2665 }),
  .out1({ S2668 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_778_ (
  .in1({ S2668, S2660 }),
  .out1({ DP_AC_din_12 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_779_ (
  .in1({ DP_IMM1_out_13, S2698 }),
  .out1({ S2669 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_780_ (
  .in1({ S2552, S2548 }),
  .out1({ S2670 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1164_ (
  .in1({ DP_ARU1_out_13, S209 }),
  .out1({ S2671 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_353_ (
  .in1({ S2671 }),
  .out1({ S2672 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_781_ (
  .in1({ S2672, S2670 }),
  .out1({ S2673 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_782_ (
  .in1({ S2673, S210 }),
  .out1({ S2674 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1165_ (
  .in1({ DP_INC_2_in_13, S211 }),
  .out1({ S2675 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1166_ (
  .in1({ S2675, S2698 }),
  .out1({ S2676 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_783_ (
  .in1({ S2676, S2674 }),
  .out1({ S2677 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_784_ (
  .in1({ S2677, S2669 }),
  .out1({ DP_AC_din_13 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_785_ (
  .in1({ DP_IMM1_out_14, S2698 }),
  .out1({ S2678 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_786_ (
  .in1({ S2552, S2549 }),
  .out1({ S2679 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1167_ (
  .in1({ DP_ARU1_out_14, S212 }),
  .out1({ S2680 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_354_ (
  .in1({ S2680 }),
  .out1({ S2681 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_787_ (
  .in1({ S2681, S2679 }),
  .out1({ S2682 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_788_ (
  .in1({ S2682, S213 }),
  .out1({ S2683 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1168_ (
  .in1({ DP_INC_2_in_14, S214 }),
  .out1({ S2684 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1169_ (
  .in1({ S2684, S2698 }),
  .out1({ S2685 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_789_ (
  .in1({ S2685, S2683 }),
  .out1({ S2686 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_790_ (
  .in1({ S2686, S2678 }),
  .out1({ DP_AC_din_14 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_791_ (
  .in1({ DP_IMM1_out_15, S2698 }),
  .out1({ S2687 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_792_ (
  .in1({ S2552, S2550 }),
  .out1({ S2688 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1170_ (
  .in1({ DP_ARU1_N, S215 }),
  .out1({ S2689 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_355_ (
  .in1({ S2689 }),
  .out1({ S2690 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_793_ (
  .in1({ S2690, S2688 }),
  .out1({ S2691 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_794_ (
  .in1({ S2691, S216 }),
  .out1({ S2692 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1171_ (
  .in1({ DP_INC_2_in_15, S217 }),
  .out1({ S2693 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1172_ (
  .in1({ S2693, S2698 }),
  .out1({ S2694 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_795_ (
  .in1({ S2694, S2692 }),
  .out1({ S2695 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_796_ (
  .in1({ S2695, S2687 }),
  .out1({ DP_AC_din_15 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_356_ (
  .in1({ S218 }),
  .out1({ S2711 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_357_ (
  .in1({ S219 }),
  .out1({ S2712 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_358_ (
  .in1({ S220 }),
  .out1({ S2713 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_359_ (
  .in1({ S221 }),
  .out1({ S2714 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_360_ (
  .in1({ S222 }),
  .out1({ S2715 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_361_ (
  .in1({ S223 }),
  .out1({ S2716 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_797_ (
  .in1({ S2713, CU_inst_0 }),
  .out1({ S2717 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1173_ (
  .in1({ S2712, S224 }),
  .out1({ S2718 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_798_ (
  .in1({ S2718, S2711 }),
  .out1({ S2719 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1174_ (
  .in1({ S225, DP_ARU1_V }),
  .out1({ S2720 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_362_ (
  .in1({ S2720 }),
  .out1({ S2721 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_799_ (
  .in1({ S2721, S2719 }),
  .out1({ S2722 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_800_ (
  .in1({ S2722, S226 }),
  .out1({ S2723 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1175_ (
  .in1({ S228, S227 }),
  .out1({ S2724 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1176_ (
  .in1({ S2724, S2713 }),
  .out1({ S2725 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_801_ (
  .in1({ S2725, S2723 }),
  .out1({ S2726 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_802_ (
  .in1({ S2726, S2717 }),
  .out1({ DP_SR_V_din })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_803_ (
  .in1({ CU_inst_1, S2713 }),
  .out1({ S2727 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_804_ (
  .in1({ S2718, S2714 }),
  .out1({ S2728 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1177_ (
  .in1({ DP_ARU1_C, S229 }),
  .out1({ S2729 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_363_ (
  .in1({ S2729 }),
  .out1({ S2730 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_805_ (
  .in1({ S2730, S2728 }),
  .out1({ S2731 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_806_ (
  .in1({ S2731, S230 }),
  .out1({ S2732 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1178_ (
  .in1({ S232, S231 }),
  .out1({ S2733 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1179_ (
  .in1({ S2733, S2713 }),
  .out1({ S2734 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_807_ (
  .in1({ S2734, S2732 }),
  .out1({ S2735 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_808_ (
  .in1({ S2735, S2727 }),
  .out1({ DP_SR_C_din })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_809_ (
  .in1({ CU_inst_2, S2713 }),
  .out1({ S2736 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_810_ (
  .in1({ S2718, S2715 }),
  .out1({ S2737 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1180_ (
  .in1({ DP_ARU1_N, S233 }),
  .out1({ S2738 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_364_ (
  .in1({ S2738 }),
  .out1({ S2739 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_811_ (
  .in1({ S2739, S2737 }),
  .out1({ S2740 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_812_ (
  .in1({ S2740, S234 }),
  .out1({ S2741 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1181_ (
  .in1({ DP_LGU1_N, S235 }),
  .out1({ S2742 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1182_ (
  .in1({ S2742, S2713 }),
  .out1({ S2743 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_813_ (
  .in1({ S2743, S2741 }),
  .out1({ S2744 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_814_ (
  .in1({ S2744, S2736 }),
  .out1({ DP_SR_N_din })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_815_ (
  .in1({ CU_inst_3, S2713 }),
  .out1({ S2745 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_816_ (
  .in1({ S2718, S2716 }),
  .out1({ S2746 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1183_ (
  .in1({ DP_ARU1_Z, S236 }),
  .out1({ S2747 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_365_ (
  .in1({ S2747 }),
  .out1({ S2748 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_817_ (
  .in1({ S2748, S2746 }),
  .out1({ S2749 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_818_ (
  .in1({ S2749, S237 }),
  .out1({ S2750 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1184_ (
  .in1({ DP_LGU1_Z, S238 }),
  .out1({ S2751 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1185_ (
  .in1({ S2751, S2713 }),
  .out1({ S2752 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_819_ (
  .in1({ S2752, S2750 }),
  .out1({ S2753 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_820_ (
  .in1({ S2753, S2745 }),
  .out1({ DP_SR_Z_din })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_366_ (
  .in1({ S239 }),
  .out1({ S2902 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_367_ (
  .in1({ S240 }),
  .out1({ S2903 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_368_ (
  .in1({ S241 }),
  .out1({ S2904 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_369_ (
  .in1({ S242 }),
  .out1({ S2905 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_370_ (
  .in1({ S243 }),
  .out1({ S2906 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_371_ (
  .in1({ S244 }),
  .out1({ S2907 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_372_ (
  .in1({ S245 }),
  .out1({ S2908 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_373_ (
  .in1({ S246 }),
  .out1({ S2909 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_374_ (
  .in1({ S247 }),
  .out1({ S2910 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_375_ (
  .in1({ S248 }),
  .out1({ S2911 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_376_ (
  .in1({ S249 }),
  .out1({ S2912 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_377_ (
  .in1({ S250 }),
  .out1({ S2913 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_378_ (
  .in1({ S251 }),
  .out1({ S2914 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_379_ (
  .in1({ S252 }),
  .out1({ S2915 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_380_ (
  .in1({ S253 }),
  .out1({ S2916 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_381_ (
  .in1({ S254 }),
  .out1({ S2754 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_382_ (
  .in1({ S255 }),
  .out1({ S2755 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_383_ (
  .in1({ S256 }),
  .out1({ S2756 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_821_ (
  .in1({ S2904, DP_INC_1_out_0 }),
  .out1({ S2757 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1186_ (
  .in1({ S2903, S257 }),
  .out1({ S2758 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_822_ (
  .in1({ S2758, S2902 }),
  .out1({ S2759 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1187_ (
  .in1({ S258, DP_IMM1_out_0 }),
  .out1({ S2760 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_384_ (
  .in1({ S2760 }),
  .out1({ S2761 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_823_ (
  .in1({ S2761, S2759 }),
  .out1({ S2762 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_824_ (
  .in1({ S2762, S259 }),
  .out1({ S2763 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1188_ (
  .in1({ S260, DP_INC_2_in_0 }),
  .out1({ S2764 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1189_ (
  .in1({ S2764, S2904 }),
  .out1({ S2765 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_825_ (
  .in1({ S2765, S2763 }),
  .out1({ S2766 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_826_ (
  .in1({ S2766, S2757 }),
  .out1({ DP_PC_din_0 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_827_ (
  .in1({ DP_INC_1_out_1, S2904 }),
  .out1({ S2767 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_828_ (
  .in1({ S2758, S2905 }),
  .out1({ S2768 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1190_ (
  .in1({ DP_IMM1_out_1, S261 }),
  .out1({ S2769 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_385_ (
  .in1({ S2769 }),
  .out1({ S2770 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_829_ (
  .in1({ S2770, S2768 }),
  .out1({ S2771 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_830_ (
  .in1({ S2771, S262 }),
  .out1({ S2772 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1191_ (
  .in1({ DP_INC_2_in_1, S263 }),
  .out1({ S2773 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1192_ (
  .in1({ S2773, S2904 }),
  .out1({ S2774 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_831_ (
  .in1({ S2774, S2772 }),
  .out1({ S2775 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_832_ (
  .in1({ S2775, S2767 }),
  .out1({ DP_PC_din_1 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_833_ (
  .in1({ DP_INC_1_out_2, S2904 }),
  .out1({ S2776 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_834_ (
  .in1({ S2758, S2906 }),
  .out1({ S2777 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1193_ (
  .in1({ DP_IMM1_out_2, S264 }),
  .out1({ S2778 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_386_ (
  .in1({ S2778 }),
  .out1({ S2779 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_835_ (
  .in1({ S2779, S2777 }),
  .out1({ S2780 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_836_ (
  .in1({ S2780, S265 }),
  .out1({ S2781 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1194_ (
  .in1({ DP_INC_2_in_2, S266 }),
  .out1({ S2782 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1195_ (
  .in1({ S2782, S2904 }),
  .out1({ S2783 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_837_ (
  .in1({ S2783, S2781 }),
  .out1({ S2784 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_838_ (
  .in1({ S2784, S2776 }),
  .out1({ DP_PC_din_2 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_839_ (
  .in1({ DP_INC_1_out_3, S2904 }),
  .out1({ S2785 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_840_ (
  .in1({ S2758, S2907 }),
  .out1({ S2786 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1196_ (
  .in1({ DP_IMM1_out_3, S267 }),
  .out1({ S2787 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_387_ (
  .in1({ S2787 }),
  .out1({ S2788 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_841_ (
  .in1({ S2788, S2786 }),
  .out1({ S2789 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_842_ (
  .in1({ S2789, S268 }),
  .out1({ S2790 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1197_ (
  .in1({ DP_INC_2_in_3, S269 }),
  .out1({ S2791 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1198_ (
  .in1({ S2791, S2904 }),
  .out1({ S2792 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_843_ (
  .in1({ S2792, S2790 }),
  .out1({ S2793 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_844_ (
  .in1({ S2793, S2785 }),
  .out1({ DP_PC_din_3 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_845_ (
  .in1({ DP_INC_1_out_4, S2904 }),
  .out1({ S2794 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_846_ (
  .in1({ S2758, S2908 }),
  .out1({ S2795 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1199_ (
  .in1({ DP_IMM1_out_4, S270 }),
  .out1({ S2796 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_388_ (
  .in1({ S2796 }),
  .out1({ S2797 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_847_ (
  .in1({ S2797, S2795 }),
  .out1({ S2798 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_848_ (
  .in1({ S2798, S271 }),
  .out1({ S2799 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1200_ (
  .in1({ DP_INC_2_in_4, S272 }),
  .out1({ S2800 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1201_ (
  .in1({ S2800, S2904 }),
  .out1({ S2801 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_849_ (
  .in1({ S2801, S2799 }),
  .out1({ S2802 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_850_ (
  .in1({ S2802, S2794 }),
  .out1({ DP_PC_din_4 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_851_ (
  .in1({ DP_INC_1_out_5, S2904 }),
  .out1({ S2803 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_852_ (
  .in1({ S2758, S2909 }),
  .out1({ S2804 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1202_ (
  .in1({ DP_IMM1_out_5, S273 }),
  .out1({ S2805 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_389_ (
  .in1({ S2805 }),
  .out1({ S2806 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_853_ (
  .in1({ S2806, S2804 }),
  .out1({ S2807 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_854_ (
  .in1({ S2807, S274 }),
  .out1({ S2808 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1203_ (
  .in1({ DP_INC_2_in_5, S275 }),
  .out1({ S2809 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1204_ (
  .in1({ S2809, S2904 }),
  .out1({ S2810 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_855_ (
  .in1({ S2810, S2808 }),
  .out1({ S2811 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_856_ (
  .in1({ S2811, S2803 }),
  .out1({ DP_PC_din_5 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_857_ (
  .in1({ DP_INC_1_out_6, S2904 }),
  .out1({ S2812 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_858_ (
  .in1({ S2758, S2910 }),
  .out1({ S2813 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1205_ (
  .in1({ DP_IMM1_out_6, S276 }),
  .out1({ S2814 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_390_ (
  .in1({ S2814 }),
  .out1({ S2815 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_859_ (
  .in1({ S2815, S2813 }),
  .out1({ S2816 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_860_ (
  .in1({ S2816, S277 }),
  .out1({ S2817 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1206_ (
  .in1({ DP_INC_2_in_6, S278 }),
  .out1({ S2818 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1207_ (
  .in1({ S2818, S2904 }),
  .out1({ S2819 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_861_ (
  .in1({ S2819, S2817 }),
  .out1({ S2820 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_862_ (
  .in1({ S2820, S2812 }),
  .out1({ DP_PC_din_6 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_863_ (
  .in1({ DP_INC_1_out_7, S2904 }),
  .out1({ S2821 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_864_ (
  .in1({ S2758, S2911 }),
  .out1({ S2822 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1208_ (
  .in1({ DP_IMM1_out_7, S279 }),
  .out1({ S2823 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_391_ (
  .in1({ S2823 }),
  .out1({ S2824 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_865_ (
  .in1({ S2824, S2822 }),
  .out1({ S2825 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_866_ (
  .in1({ S2825, S280 }),
  .out1({ S2826 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1209_ (
  .in1({ DP_INC_2_in_7, S281 }),
  .out1({ S2827 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1210_ (
  .in1({ S2827, S2904 }),
  .out1({ S2828 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_867_ (
  .in1({ S2828, S2826 }),
  .out1({ S2829 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_868_ (
  .in1({ S2829, S2821 }),
  .out1({ DP_PC_din_7 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_869_ (
  .in1({ DP_INC_1_out_8, S2904 }),
  .out1({ S2830 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_870_ (
  .in1({ S2758, S2912 }),
  .out1({ S2831 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1211_ (
  .in1({ DP_IMM1_out_8, S282 }),
  .out1({ S2832 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_392_ (
  .in1({ S2832 }),
  .out1({ S2833 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_871_ (
  .in1({ S2833, S2831 }),
  .out1({ S2834 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_872_ (
  .in1({ S2834, S283 }),
  .out1({ S2835 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1212_ (
  .in1({ DP_INC_2_in_8, S284 }),
  .out1({ S2836 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1213_ (
  .in1({ S2836, S2904 }),
  .out1({ S2837 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_873_ (
  .in1({ S2837, S2835 }),
  .out1({ S2838 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_874_ (
  .in1({ S2838, S2830 }),
  .out1({ DP_PC_din_8 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_875_ (
  .in1({ DP_INC_1_out_9, S2904 }),
  .out1({ S2839 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_876_ (
  .in1({ S2758, S2913 }),
  .out1({ S2840 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1214_ (
  .in1({ DP_IMM1_out_9, S285 }),
  .out1({ S2841 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_393_ (
  .in1({ S2841 }),
  .out1({ S2842 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_877_ (
  .in1({ S2842, S2840 }),
  .out1({ S2843 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_878_ (
  .in1({ S2843, S286 }),
  .out1({ S2844 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1215_ (
  .in1({ DP_INC_2_in_9, S287 }),
  .out1({ S2845 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1216_ (
  .in1({ S2845, S2904 }),
  .out1({ S2846 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_879_ (
  .in1({ S2846, S2844 }),
  .out1({ S2847 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_880_ (
  .in1({ S2847, S2839 }),
  .out1({ DP_PC_din_9 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_881_ (
  .in1({ DP_INC_1_out_10, S2904 }),
  .out1({ S2848 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_882_ (
  .in1({ S2758, S2914 }),
  .out1({ S2849 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1217_ (
  .in1({ DP_IMM1_out_10, S288 }),
  .out1({ S2850 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_394_ (
  .in1({ S2850 }),
  .out1({ S2851 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_883_ (
  .in1({ S2851, S2849 }),
  .out1({ S2852 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_884_ (
  .in1({ S2852, S289 }),
  .out1({ S2853 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1218_ (
  .in1({ DP_INC_2_in_10, S290 }),
  .out1({ S2854 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1219_ (
  .in1({ S2854, S2904 }),
  .out1({ S2855 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_885_ (
  .in1({ S2855, S2853 }),
  .out1({ S2856 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_886_ (
  .in1({ S2856, S2848 }),
  .out1({ DP_PC_din_10 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_887_ (
  .in1({ DP_INC_1_out_11, S2904 }),
  .out1({ S2857 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_888_ (
  .in1({ S2758, S2915 }),
  .out1({ S2858 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1220_ (
  .in1({ DP_IMM1_out_11, S291 }),
  .out1({ S2859 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_395_ (
  .in1({ S2859 }),
  .out1({ S2860 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_889_ (
  .in1({ S2860, S2858 }),
  .out1({ S2861 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_890_ (
  .in1({ S2861, S292 }),
  .out1({ S2862 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1221_ (
  .in1({ DP_INC_2_in_11, S293 }),
  .out1({ S2863 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1222_ (
  .in1({ S2863, S2904 }),
  .out1({ S2864 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_891_ (
  .in1({ S2864, S2862 }),
  .out1({ S2865 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_892_ (
  .in1({ S2865, S2857 }),
  .out1({ DP_PC_din_11 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_893_ (
  .in1({ DP_INC_1_out_12, S2904 }),
  .out1({ S2866 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_894_ (
  .in1({ S2758, S2916 }),
  .out1({ S2867 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1223_ (
  .in1({ DP_IMM1_out_12, S294 }),
  .out1({ S2868 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_396_ (
  .in1({ S2868 }),
  .out1({ S2869 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_895_ (
  .in1({ S2869, S2867 }),
  .out1({ S2870 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_896_ (
  .in1({ S2870, S295 }),
  .out1({ S2871 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1224_ (
  .in1({ DP_INC_2_in_12, S296 }),
  .out1({ S2872 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1225_ (
  .in1({ S2872, S2904 }),
  .out1({ S2873 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_897_ (
  .in1({ S2873, S2871 }),
  .out1({ S2874 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_898_ (
  .in1({ S2874, S2866 }),
  .out1({ DP_PC_din_12 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_899_ (
  .in1({ DP_INC_1_out_13, S2904 }),
  .out1({ S2875 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_900_ (
  .in1({ S2758, S2754 }),
  .out1({ S2876 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1226_ (
  .in1({ DP_IMM1_out_13, S297 }),
  .out1({ S2877 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_397_ (
  .in1({ S2877 }),
  .out1({ S2878 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_901_ (
  .in1({ S2878, S2876 }),
  .out1({ S2879 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_902_ (
  .in1({ S2879, S298 }),
  .out1({ S2880 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1227_ (
  .in1({ DP_INC_2_in_13, S299 }),
  .out1({ S2881 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1228_ (
  .in1({ S2881, S2904 }),
  .out1({ S2882 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_903_ (
  .in1({ S2882, S2880 }),
  .out1({ S2883 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_904_ (
  .in1({ S2883, S2875 }),
  .out1({ DP_PC_din_13 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_905_ (
  .in1({ DP_INC_1_out_14, S2904 }),
  .out1({ S2884 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_906_ (
  .in1({ S2758, S2755 }),
  .out1({ S2885 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1229_ (
  .in1({ DP_IMM1_out_14, S300 }),
  .out1({ S2886 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_398_ (
  .in1({ S2886 }),
  .out1({ S2887 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_907_ (
  .in1({ S2887, S2885 }),
  .out1({ S2888 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_908_ (
  .in1({ S2888, S301 }),
  .out1({ S2889 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1230_ (
  .in1({ DP_INC_2_in_14, S302 }),
  .out1({ S2890 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1231_ (
  .in1({ S2890, S2904 }),
  .out1({ S2891 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_909_ (
  .in1({ S2891, S2889 }),
  .out1({ S2892 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_910_ (
  .in1({ S2892, S2884 }),
  .out1({ DP_PC_din_14 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_911_ (
  .in1({ DP_INC_1_out_15, S2904 }),
  .out1({ S2893 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_912_ (
  .in1({ S2758, S2756 }),
  .out1({ S2894 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1232_ (
  .in1({ DP_IMM1_out_15, S303 }),
  .out1({ S2895 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_399_ (
  .in1({ S2895 }),
  .out1({ S2896 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_913_ (
  .in1({ S2896, S2894 }),
  .out1({ S2897 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_914_ (
  .in1({ S2897, S304 }),
  .out1({ S2898 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1233_ (
  .in1({ DP_INC_2_in_15, S305 }),
  .out1({ S2899 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1234_ (
  .in1({ S2899, S2904 }),
  .out1({ S2900 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_915_ (
  .in1({ S2900, S2898 }),
  .out1({ S2901 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_916_ (
  .in1({ S2901, S2893 }),
  .out1({ DP_PC_din_15 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_400_ (
  .in1({ S306 }),
  .out1({ S2917 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_917_ (
  .in1({ S307, S2917 }),
  .out1({ S2918 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1235_ (
  .in1({ S2918, DP_INC_2_in_0 }),
  .out1({ S2919 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1236_ (
  .in1({ S308, DP_INC2_out_0 }),
  .out1({ S2920 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1237_ (
  .in1({ S2920, S2919 }),
  .out1({ DP_IN_din_0 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1238_ (
  .in1({ S2918, DP_INC_2_in_1 }),
  .out1({ S2921 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1239_ (
  .in1({ DP_INC2_out_1, S309 }),
  .out1({ S2922 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1240_ (
  .in1({ S2922, S2921 }),
  .out1({ DP_IN_din_1 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1241_ (
  .in1({ S2918, DP_INC_2_in_2 }),
  .out1({ S2923 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1242_ (
  .in1({ DP_INC2_out_2, S310 }),
  .out1({ S2924 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1243_ (
  .in1({ S2924, S2923 }),
  .out1({ DP_IN_din_2 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1244_ (
  .in1({ S2918, DP_INC_2_in_3 }),
  .out1({ S2925 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1245_ (
  .in1({ DP_INC2_out_3, S311 }),
  .out1({ S2926 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1246_ (
  .in1({ S2926, S2925 }),
  .out1({ DP_IN_din_3 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1247_ (
  .in1({ S2918, DP_INC_2_in_4 }),
  .out1({ S2927 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1248_ (
  .in1({ DP_INC2_out_4, S312 }),
  .out1({ S2928 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1249_ (
  .in1({ S2928, S2927 }),
  .out1({ DP_IN_din_4 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1250_ (
  .in1({ S2918, DP_INC_2_in_5 }),
  .out1({ S2929 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1251_ (
  .in1({ DP_INC2_out_5, S313 }),
  .out1({ S2930 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1252_ (
  .in1({ S2930, S2929 }),
  .out1({ DP_IN_din_5 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1253_ (
  .in1({ S2918, DP_INC_2_in_6 }),
  .out1({ S2931 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1254_ (
  .in1({ DP_INC2_out_6, S314 }),
  .out1({ S2932 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1255_ (
  .in1({ S2932, S2931 }),
  .out1({ DP_IN_din_6 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1256_ (
  .in1({ S2918, DP_INC_2_in_7 }),
  .out1({ S2933 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1257_ (
  .in1({ DP_INC2_out_7, S315 }),
  .out1({ S2934 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1258_ (
  .in1({ S2934, S2933 }),
  .out1({ DP_IN_din_7 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1259_ (
  .in1({ S2918, DP_INC_2_in_8 }),
  .out1({ S2935 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1260_ (
  .in1({ DP_INC2_out_8, S316 }),
  .out1({ S2936 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1261_ (
  .in1({ S2936, S2935 }),
  .out1({ DP_IN_din_8 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1262_ (
  .in1({ S2918, DP_INC_2_in_9 }),
  .out1({ S2937 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1263_ (
  .in1({ DP_INC2_out_9, S317 }),
  .out1({ S2938 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1264_ (
  .in1({ S2938, S2937 }),
  .out1({ DP_IN_din_9 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1265_ (
  .in1({ S2918, DP_INC_2_in_10 }),
  .out1({ S2939 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1266_ (
  .in1({ DP_INC2_out_10, S318 }),
  .out1({ S2940 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1267_ (
  .in1({ S2940, S2939 }),
  .out1({ DP_IN_din_10 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1268_ (
  .in1({ S2918, DP_INC_2_in_11 }),
  .out1({ S2941 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1269_ (
  .in1({ DP_INC2_out_11, S319 }),
  .out1({ S2942 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1270_ (
  .in1({ S2942, S2941 }),
  .out1({ DP_IN_din_11 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1271_ (
  .in1({ S2918, DP_INC_2_in_12 }),
  .out1({ S2943 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1272_ (
  .in1({ DP_INC2_out_12, S320 }),
  .out1({ S2944 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1273_ (
  .in1({ S2944, S2943 }),
  .out1({ DP_IN_din_12 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1274_ (
  .in1({ S2918, DP_INC_2_in_13 }),
  .out1({ S2945 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1275_ (
  .in1({ DP_INC2_out_13, S321 }),
  .out1({ S2946 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1276_ (
  .in1({ S2946, S2945 }),
  .out1({ DP_IN_din_13 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1277_ (
  .in1({ S2918, DP_INC_2_in_14 }),
  .out1({ S2947 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1278_ (
  .in1({ DP_INC2_out_14, S322 }),
  .out1({ S2948 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1279_ (
  .in1({ S2948, S2947 }),
  .out1({ DP_IN_din_14 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1280_ (
  .in1({ S2918, DP_INC_2_in_15 }),
  .out1({ S2949 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1281_ (
  .in1({ DP_INC2_out_15, S323 }),
  .out1({ S2950 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1282_ (
  .in1({ S2950, S2949 }),
  .out1({ DP_IN_din_15 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_401_ (
  .in1({ S324 }),
  .out1({ S3099 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_402_ (
  .in1({ S325 }),
  .out1({ S3100 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_403_ (
  .in1({ S326 }),
  .out1({ S3101 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_404_ (
  .in1({ S327 }),
  .out1({ S3102 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_405_ (
  .in1({ S328 }),
  .out1({ S3103 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_406_ (
  .in1({ S329 }),
  .out1({ S3104 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_407_ (
  .in1({ S330 }),
  .out1({ S3105 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_408_ (
  .in1({ S331 }),
  .out1({ S3106 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_409_ (
  .in1({ S332 }),
  .out1({ S3107 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_410_ (
  .in1({ S333 }),
  .out1({ S3108 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_411_ (
  .in1({ S334 }),
  .out1({ S3109 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_412_ (
  .in1({ S335 }),
  .out1({ S3110 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_413_ (
  .in1({ S336 }),
  .out1({ S3111 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_414_ (
  .in1({ S337 }),
  .out1({ S3112 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_415_ (
  .in1({ S338 }),
  .out1({ S3113 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_416_ (
  .in1({ S339 }),
  .out1({ S2951 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_417_ (
  .in1({ S340 }),
  .out1({ S2952 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_418_ (
  .in1({ S341 }),
  .out1({ S2953 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_918_ (
  .in1({ S3101, DP_IN_dout_0 }),
  .out1({ S2954 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1283_ (
  .in1({ S3100, S342 }),
  .out1({ S2955 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_919_ (
  .in1({ S2955, S3099 }),
  .out1({ S2956 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1284_ (
  .in1({ S343, DP_AC_dout_0 }),
  .out1({ S2957 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_419_ (
  .in1({ S2957 }),
  .out1({ S2958 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_920_ (
  .in1({ S2958, S2956 }),
  .out1({ S2959 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_921_ (
  .in1({ S2959, S344 }),
  .out1({ S2960 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1285_ (
  .in1({ S345, DP_INC_1_out_0 }),
  .out1({ S2961 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1286_ (
  .in1({ S2961, S3101 }),
  .out1({ S2962 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_922_ (
  .in1({ S2962, S2960 }),
  .out1({ S2963 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_923_ (
  .in1({ S2963, S2954 }),
  .out1({ DP_TriBuff_in_0 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_924_ (
  .in1({ DP_IN_dout_1, S3101 }),
  .out1({ S2964 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_925_ (
  .in1({ S2955, S3102 }),
  .out1({ S2965 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1287_ (
  .in1({ DP_AC_dout_1, S346 }),
  .out1({ S2966 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_420_ (
  .in1({ S2966 }),
  .out1({ S2967 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_926_ (
  .in1({ S2967, S2965 }),
  .out1({ S2968 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_927_ (
  .in1({ S2968, S347 }),
  .out1({ S2969 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1288_ (
  .in1({ DP_INC_1_out_1, S348 }),
  .out1({ S2970 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1289_ (
  .in1({ S2970, S3101 }),
  .out1({ S2971 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_928_ (
  .in1({ S2971, S2969 }),
  .out1({ S2972 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_929_ (
  .in1({ S2972, S2964 }),
  .out1({ DP_TriBuff_in_1 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_930_ (
  .in1({ DP_IN_dout_2, S3101 }),
  .out1({ S2973 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_931_ (
  .in1({ S2955, S3103 }),
  .out1({ S2974 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1290_ (
  .in1({ DP_AC_dout_2, S349 }),
  .out1({ S2975 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_421_ (
  .in1({ S2975 }),
  .out1({ S2976 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_932_ (
  .in1({ S2976, S2974 }),
  .out1({ S2977 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_933_ (
  .in1({ S2977, S350 }),
  .out1({ S2978 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1291_ (
  .in1({ DP_INC_1_out_2, S351 }),
  .out1({ S2979 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1292_ (
  .in1({ S2979, S3101 }),
  .out1({ S2980 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_934_ (
  .in1({ S2980, S2978 }),
  .out1({ S2981 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_935_ (
  .in1({ S2981, S2973 }),
  .out1({ DP_TriBuff_in_2 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_936_ (
  .in1({ DP_IN_dout_3, S3101 }),
  .out1({ S2982 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_937_ (
  .in1({ S2955, S3104 }),
  .out1({ S2983 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1293_ (
  .in1({ DP_AC_dout_3, S352 }),
  .out1({ S2984 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_422_ (
  .in1({ S2984 }),
  .out1({ S2985 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_938_ (
  .in1({ S2985, S2983 }),
  .out1({ S2986 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_939_ (
  .in1({ S2986, S353 }),
  .out1({ S2987 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1294_ (
  .in1({ DP_INC_1_out_3, S354 }),
  .out1({ S2988 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1295_ (
  .in1({ S2988, S3101 }),
  .out1({ S2989 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_940_ (
  .in1({ S2989, S2987 }),
  .out1({ S2990 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_941_ (
  .in1({ S2990, S2982 }),
  .out1({ DP_TriBuff_in_3 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_942_ (
  .in1({ DP_IN_dout_4, S3101 }),
  .out1({ S2991 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_943_ (
  .in1({ S2955, S3105 }),
  .out1({ S2992 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1296_ (
  .in1({ DP_AC_dout_4, S355 }),
  .out1({ S2993 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_423_ (
  .in1({ S2993 }),
  .out1({ S2994 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_944_ (
  .in1({ S2994, S2992 }),
  .out1({ S2995 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_945_ (
  .in1({ S2995, S356 }),
  .out1({ S2996 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1297_ (
  .in1({ DP_INC_1_out_4, S357 }),
  .out1({ S2997 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1298_ (
  .in1({ S2997, S3101 }),
  .out1({ S2998 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_946_ (
  .in1({ S2998, S2996 }),
  .out1({ S2999 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_947_ (
  .in1({ S2999, S2991 }),
  .out1({ DP_TriBuff_in_4 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_948_ (
  .in1({ DP_IN_dout_5, S3101 }),
  .out1({ S3000 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_949_ (
  .in1({ S2955, S3106 }),
  .out1({ S3001 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1299_ (
  .in1({ DP_AC_dout_5, S358 }),
  .out1({ S3002 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_424_ (
  .in1({ S3002 }),
  .out1({ S3003 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_950_ (
  .in1({ S3003, S3001 }),
  .out1({ S3004 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_951_ (
  .in1({ S3004, S359 }),
  .out1({ S3005 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1300_ (
  .in1({ DP_INC_1_out_5, S360 }),
  .out1({ S3006 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1301_ (
  .in1({ S3006, S3101 }),
  .out1({ S3007 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_952_ (
  .in1({ S3007, S3005 }),
  .out1({ S3008 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_953_ (
  .in1({ S3008, S3000 }),
  .out1({ DP_TriBuff_in_5 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_954_ (
  .in1({ DP_IN_dout_6, S3101 }),
  .out1({ S3009 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_955_ (
  .in1({ S2955, S3107 }),
  .out1({ S3010 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1302_ (
  .in1({ DP_AC_dout_6, S361 }),
  .out1({ S3011 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_425_ (
  .in1({ S3011 }),
  .out1({ S3012 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_956_ (
  .in1({ S3012, S3010 }),
  .out1({ S3013 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_957_ (
  .in1({ S3013, S362 }),
  .out1({ S3014 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1303_ (
  .in1({ DP_INC_1_out_6, S363 }),
  .out1({ S3015 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1304_ (
  .in1({ S3015, S3101 }),
  .out1({ S3016 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_958_ (
  .in1({ S3016, S3014 }),
  .out1({ S3017 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_959_ (
  .in1({ S3017, S3009 }),
  .out1({ DP_TriBuff_in_6 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_960_ (
  .in1({ DP_IN_dout_7, S3101 }),
  .out1({ S3018 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_961_ (
  .in1({ S2955, S3108 }),
  .out1({ S3019 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1305_ (
  .in1({ DP_AC_dout_7, S364 }),
  .out1({ S3020 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_426_ (
  .in1({ S3020 }),
  .out1({ S3021 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_962_ (
  .in1({ S3021, S3019 }),
  .out1({ S3022 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_963_ (
  .in1({ S3022, S365 }),
  .out1({ S3023 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1306_ (
  .in1({ DP_INC_1_out_7, S366 }),
  .out1({ S3024 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1307_ (
  .in1({ S3024, S3101 }),
  .out1({ S3025 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_964_ (
  .in1({ S3025, S3023 }),
  .out1({ S3026 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_965_ (
  .in1({ S3026, S3018 }),
  .out1({ DP_TriBuff_in_7 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_966_ (
  .in1({ DP_IN_dout_8, S3101 }),
  .out1({ S3027 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_967_ (
  .in1({ S2955, S3109 }),
  .out1({ S3028 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1308_ (
  .in1({ DP_AC_dout_8, S367 }),
  .out1({ S3029 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_427_ (
  .in1({ S3029 }),
  .out1({ S3030 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_968_ (
  .in1({ S3030, S3028 }),
  .out1({ S3031 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_969_ (
  .in1({ S3031, S368 }),
  .out1({ S3032 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1309_ (
  .in1({ DP_INC_1_out_8, S369 }),
  .out1({ S3033 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1310_ (
  .in1({ S3033, S3101 }),
  .out1({ S3034 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_970_ (
  .in1({ S3034, S3032 }),
  .out1({ S3035 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_971_ (
  .in1({ S3035, S3027 }),
  .out1({ DP_TriBuff_in_8 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_972_ (
  .in1({ DP_IN_dout_9, S3101 }),
  .out1({ S3036 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_973_ (
  .in1({ S2955, S3110 }),
  .out1({ S3037 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1311_ (
  .in1({ DP_AC_dout_9, S370 }),
  .out1({ S3038 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_428_ (
  .in1({ S3038 }),
  .out1({ S3039 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_974_ (
  .in1({ S3039, S3037 }),
  .out1({ S3040 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_975_ (
  .in1({ S3040, S371 }),
  .out1({ S3041 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1312_ (
  .in1({ DP_INC_1_out_9, S372 }),
  .out1({ S3042 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1313_ (
  .in1({ S3042, S3101 }),
  .out1({ S3043 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_976_ (
  .in1({ S3043, S3041 }),
  .out1({ S3044 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_977_ (
  .in1({ S3044, S3036 }),
  .out1({ DP_TriBuff_in_9 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_978_ (
  .in1({ DP_IN_dout_10, S3101 }),
  .out1({ S3045 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_979_ (
  .in1({ S2955, S3111 }),
  .out1({ S3046 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1314_ (
  .in1({ DP_AC_dout_10, S373 }),
  .out1({ S3047 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_429_ (
  .in1({ S3047 }),
  .out1({ S3048 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_980_ (
  .in1({ S3048, S3046 }),
  .out1({ S3049 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_981_ (
  .in1({ S3049, S374 }),
  .out1({ S3050 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1315_ (
  .in1({ DP_INC_1_out_10, S375 }),
  .out1({ S3051 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1316_ (
  .in1({ S3051, S3101 }),
  .out1({ S3052 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_982_ (
  .in1({ S3052, S3050 }),
  .out1({ S3053 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_983_ (
  .in1({ S3053, S3045 }),
  .out1({ DP_TriBuff_in_10 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_984_ (
  .in1({ DP_IN_dout_11, S3101 }),
  .out1({ S3054 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_985_ (
  .in1({ S2955, S3112 }),
  .out1({ S3055 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1317_ (
  .in1({ DP_AC_dout_11, S376 }),
  .out1({ S3056 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_430_ (
  .in1({ S3056 }),
  .out1({ S3057 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_986_ (
  .in1({ S3057, S3055 }),
  .out1({ S3058 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_987_ (
  .in1({ S3058, S377 }),
  .out1({ S3059 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1318_ (
  .in1({ DP_INC_1_out_11, S378 }),
  .out1({ S3060 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1319_ (
  .in1({ S3060, S3101 }),
  .out1({ S3061 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_988_ (
  .in1({ S3061, S3059 }),
  .out1({ S3062 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_989_ (
  .in1({ S3062, S3054 }),
  .out1({ DP_TriBuff_in_11 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_990_ (
  .in1({ DP_IN_dout_12, S3101 }),
  .out1({ S3063 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_991_ (
  .in1({ S2955, S3113 }),
  .out1({ S3064 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1320_ (
  .in1({ DP_AC_dout_12, S379 }),
  .out1({ S3065 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_431_ (
  .in1({ S3065 }),
  .out1({ S3066 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_992_ (
  .in1({ S3066, S3064 }),
  .out1({ S3067 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_993_ (
  .in1({ S3067, S380 }),
  .out1({ S3068 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1321_ (
  .in1({ DP_INC_1_out_12, S381 }),
  .out1({ S3069 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1322_ (
  .in1({ S3069, S3101 }),
  .out1({ S3070 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_994_ (
  .in1({ S3070, S3068 }),
  .out1({ S3071 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_995_ (
  .in1({ S3071, S3063 }),
  .out1({ DP_TriBuff_in_12 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_996_ (
  .in1({ DP_IN_dout_13, S3101 }),
  .out1({ S3072 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_997_ (
  .in1({ S2955, S2951 }),
  .out1({ S3073 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1323_ (
  .in1({ DP_AC_dout_13, S382 }),
  .out1({ S3074 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_432_ (
  .in1({ S3074 }),
  .out1({ S3075 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_998_ (
  .in1({ S3075, S3073 }),
  .out1({ S3076 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_999_ (
  .in1({ S3076, S383 }),
  .out1({ S3077 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1324_ (
  .in1({ DP_INC_1_out_13, S384 }),
  .out1({ S3078 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1325_ (
  .in1({ S3078, S3101 }),
  .out1({ S3079 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1000_ (
  .in1({ S3079, S3077 }),
  .out1({ S3080 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1001_ (
  .in1({ S3080, S3072 }),
  .out1({ DP_TriBuff_in_13 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1002_ (
  .in1({ DP_IN_dout_14, S3101 }),
  .out1({ S3081 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1003_ (
  .in1({ S2955, S2952 }),
  .out1({ S3082 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1326_ (
  .in1({ DP_AC_dout_14, S385 }),
  .out1({ S3083 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_433_ (
  .in1({ S3083 }),
  .out1({ S3084 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1004_ (
  .in1({ S3084, S3082 }),
  .out1({ S3085 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1005_ (
  .in1({ S3085, S386 }),
  .out1({ S3086 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1327_ (
  .in1({ DP_INC_1_out_14, S387 }),
  .out1({ S3087 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1328_ (
  .in1({ S3087, S3101 }),
  .out1({ S3088 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1006_ (
  .in1({ S3088, S3086 }),
  .out1({ S3089 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1007_ (
  .in1({ S3089, S3081 }),
  .out1({ DP_TriBuff_in_14 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1008_ (
  .in1({ DP_IN_dout_15, S3101 }),
  .out1({ S3090 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1009_ (
  .in1({ S2955, S2953 }),
  .out1({ S3091 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1329_ (
  .in1({ DP_AC_dout_15, S388 }),
  .out1({ S3092 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_434_ (
  .in1({ S3092 }),
  .out1({ S3093 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1010_ (
  .in1({ S3093, S3091 }),
  .out1({ S3094 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1011_ (
  .in1({ S3094, S389 }),
  .out1({ S3095 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1330_ (
  .in1({ DP_INC_1_out_15, S390 }),
  .out1({ S3096 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1331_ (
  .in1({ S3096, S3101 }),
  .out1({ S3097 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1012_ (
  .in1({ S3097, S3095 }),
  .out1({ S3098 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1013_ (
  .in1({ S3098, S3090 }),
  .out1({ DP_TriBuff_in_15 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_435_ (
  .in1({ S391 }),
  .out1({ S3262 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_436_ (
  .in1({ S21 }),
  .out1({ S3263 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_437_ (
  .in1({ S392 }),
  .out1({ S3264 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_438_ (
  .in1({ S393 }),
  .out1({ S3265 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_439_ (
  .in1({ S394 }),
  .out1({ S3266 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_440_ (
  .in1({ S395 }),
  .out1({ S3267 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_441_ (
  .in1({ S396 }),
  .out1({ S3268 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_442_ (
  .in1({ S397 }),
  .out1({ S3269 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_443_ (
  .in1({ S398 }),
  .out1({ S3270 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_444_ (
  .in1({ S399 }),
  .out1({ S3271 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_445_ (
  .in1({ S400 }),
  .out1({ S3272 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_446_ (
  .in1({ S401 }),
  .out1({ S3273 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_447_ (
  .in1({ S402 }),
  .out1({ S3274 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_448_ (
  .in1({ S403 }),
  .out1({ S3275 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_449_ (
  .in1({ S404 }),
  .out1({ S3276 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_450_ (
  .in1({ S405 }),
  .out1({ S3114 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_451_ (
  .in1({ S406 }),
  .out1({ S3115 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_452_ (
  .in1({ S407 }),
  .out1({ S3116 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1014_ (
  .in1({ S3264, DP_IN_dout_0 }),
  .out1({ S3117 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1332_ (
  .in1({ S3263, S408 }),
  .out1({ S3118 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1015_ (
  .in1({ S3118, S3262 }),
  .out1({ S3119 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1333_ (
  .in1({ S22, DP_INC_1_in_0 }),
  .out1({ S3120 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_453_ (
  .in1({ S3120 }),
  .out1({ S3121 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1016_ (
  .in1({ S3121, S3119 }),
  .out1({ S3122 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1017_ (
  .in1({ S3122, S409 }),
  .out1({ S3123 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1334_ (
  .in1({ S410, DP_IMM1_out_0 }),
  .out1({ S3124 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1335_ (
  .in1({ S3124, S3264 }),
  .out1({ S3125 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1018_ (
  .in1({ S3125, S3123 }),
  .out1({ S3126 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1019_ (
  .in1({ S3126, S3117 }),
  .out1({ DP_addrBus_0 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1020_ (
  .in1({ DP_IN_dout_1, S3264 }),
  .out1({ S3127 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1021_ (
  .in1({ S3118, S3265 }),
  .out1({ S3128 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1336_ (
  .in1({ DP_INC_1_in_1, S23 }),
  .out1({ S3129 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_454_ (
  .in1({ S3129 }),
  .out1({ S3130 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1022_ (
  .in1({ S3130, S3128 }),
  .out1({ S3131 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1023_ (
  .in1({ S3131, S411 }),
  .out1({ S3132 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1337_ (
  .in1({ DP_IMM1_out_1, S412 }),
  .out1({ S3133 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1338_ (
  .in1({ S3133, S3264 }),
  .out1({ S3134 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1024_ (
  .in1({ S3134, S3132 }),
  .out1({ S3135 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1025_ (
  .in1({ S3135, S3127 }),
  .out1({ DP_addrBus_1 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1026_ (
  .in1({ DP_IN_dout_2, S3264 }),
  .out1({ S3136 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1027_ (
  .in1({ S3118, S3266 }),
  .out1({ S3137 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1339_ (
  .in1({ DP_INC_1_in_2, S24 }),
  .out1({ S3138 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_455_ (
  .in1({ S3138 }),
  .out1({ S3139 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1028_ (
  .in1({ S3139, S3137 }),
  .out1({ S3140 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1029_ (
  .in1({ S3140, S413 }),
  .out1({ S3141 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1340_ (
  .in1({ DP_IMM1_out_2, S414 }),
  .out1({ S3142 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1341_ (
  .in1({ S3142, S3264 }),
  .out1({ S3143 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1030_ (
  .in1({ S3143, S3141 }),
  .out1({ S3144 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1031_ (
  .in1({ S3144, S3136 }),
  .out1({ DP_addrBus_2 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1032_ (
  .in1({ DP_IN_dout_3, S3264 }),
  .out1({ S3145 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1033_ (
  .in1({ S3118, S3267 }),
  .out1({ S3146 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1342_ (
  .in1({ DP_INC_1_in_3, S25 }),
  .out1({ S3147 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_456_ (
  .in1({ S3147 }),
  .out1({ S3148 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1034_ (
  .in1({ S3148, S3146 }),
  .out1({ S3149 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1035_ (
  .in1({ S3149, S415 }),
  .out1({ S3150 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1343_ (
  .in1({ DP_IMM1_out_3, S416 }),
  .out1({ S3151 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1344_ (
  .in1({ S3151, S3264 }),
  .out1({ S3152 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1036_ (
  .in1({ S3152, S3150 }),
  .out1({ S3153 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1037_ (
  .in1({ S3153, S3145 }),
  .out1({ DP_addrBus_3 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1038_ (
  .in1({ DP_IN_dout_4, S3264 }),
  .out1({ S3154 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1039_ (
  .in1({ S3118, S3268 }),
  .out1({ S3155 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1345_ (
  .in1({ DP_INC_1_in_4, S26 }),
  .out1({ S3156 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_457_ (
  .in1({ S3156 }),
  .out1({ S3157 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1040_ (
  .in1({ S3157, S3155 }),
  .out1({ S3158 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1041_ (
  .in1({ S3158, S417 }),
  .out1({ S3159 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1346_ (
  .in1({ DP_IMM1_out_4, S418 }),
  .out1({ S3160 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1347_ (
  .in1({ S3160, S3264 }),
  .out1({ S3161 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1042_ (
  .in1({ S3161, S3159 }),
  .out1({ S3162 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1043_ (
  .in1({ S3162, S3154 }),
  .out1({ DP_addrBus_4 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1044_ (
  .in1({ DP_IN_dout_5, S3264 }),
  .out1({ S3163 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1045_ (
  .in1({ S3118, S3269 }),
  .out1({ S3164 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1348_ (
  .in1({ DP_INC_1_in_5, S27 }),
  .out1({ S3165 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_458_ (
  .in1({ S3165 }),
  .out1({ S3166 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1046_ (
  .in1({ S3166, S3164 }),
  .out1({ S3167 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1047_ (
  .in1({ S3167, S419 }),
  .out1({ S3168 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1349_ (
  .in1({ DP_IMM1_out_5, S420 }),
  .out1({ S3169 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1350_ (
  .in1({ S3169, S3264 }),
  .out1({ S3170 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1048_ (
  .in1({ S3170, S3168 }),
  .out1({ S3171 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1049_ (
  .in1({ S3171, S3163 }),
  .out1({ DP_addrBus_5 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1050_ (
  .in1({ DP_IN_dout_6, S3264 }),
  .out1({ S3172 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1051_ (
  .in1({ S3118, S3270 }),
  .out1({ S3173 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1351_ (
  .in1({ DP_INC_1_in_6, S28 }),
  .out1({ S3174 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_459_ (
  .in1({ S3174 }),
  .out1({ S3175 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1052_ (
  .in1({ S3175, S3173 }),
  .out1({ S3176 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1053_ (
  .in1({ S3176, S421 }),
  .out1({ S3177 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1352_ (
  .in1({ DP_IMM1_out_6, S422 }),
  .out1({ S3178 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1353_ (
  .in1({ S3178, S3264 }),
  .out1({ S3179 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1054_ (
  .in1({ S3179, S3177 }),
  .out1({ S3180 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1055_ (
  .in1({ S3180, S3172 }),
  .out1({ DP_addrBus_6 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1056_ (
  .in1({ DP_IN_dout_7, S3264 }),
  .out1({ S3181 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1057_ (
  .in1({ S3118, S3271 }),
  .out1({ S3182 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1354_ (
  .in1({ DP_INC_1_in_7, S29 }),
  .out1({ S3183 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_460_ (
  .in1({ S3183 }),
  .out1({ S3184 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1058_ (
  .in1({ S3184, S3182 }),
  .out1({ S3185 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1059_ (
  .in1({ S3185, S423 }),
  .out1({ S3186 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1355_ (
  .in1({ DP_IMM1_out_7, S424 }),
  .out1({ S3187 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1356_ (
  .in1({ S3187, S3264 }),
  .out1({ S3188 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1060_ (
  .in1({ S3188, S3186 }),
  .out1({ S3189 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1061_ (
  .in1({ S3189, S3181 }),
  .out1({ DP_addrBus_7 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1062_ (
  .in1({ DP_IN_dout_8, S3264 }),
  .out1({ S3190 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1063_ (
  .in1({ S3118, S3272 }),
  .out1({ S3191 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1357_ (
  .in1({ DP_INC_1_in_8, S30 }),
  .out1({ S3192 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_461_ (
  .in1({ S3192 }),
  .out1({ S3193 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1064_ (
  .in1({ S3193, S3191 }),
  .out1({ S3194 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1065_ (
  .in1({ S3194, S425 }),
  .out1({ S3195 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1358_ (
  .in1({ DP_IMM1_out_8, S426 }),
  .out1({ S3196 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1359_ (
  .in1({ S3196, S3264 }),
  .out1({ S3197 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1066_ (
  .in1({ S3197, S3195 }),
  .out1({ S3198 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1067_ (
  .in1({ S3198, S3190 }),
  .out1({ DP_addrBus_8 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1068_ (
  .in1({ DP_IN_dout_9, S3264 }),
  .out1({ S3199 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1069_ (
  .in1({ S3118, S3273 }),
  .out1({ S3200 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1360_ (
  .in1({ DP_INC_1_in_9, S31 }),
  .out1({ S3201 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_462_ (
  .in1({ S3201 }),
  .out1({ S3202 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1070_ (
  .in1({ S3202, S3200 }),
  .out1({ S3203 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1071_ (
  .in1({ S3203, S427 }),
  .out1({ S3204 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1361_ (
  .in1({ DP_IMM1_out_9, S428 }),
  .out1({ S3205 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1362_ (
  .in1({ S3205, S3264 }),
  .out1({ S3206 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1072_ (
  .in1({ S3206, S3204 }),
  .out1({ S3207 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1073_ (
  .in1({ S3207, S3199 }),
  .out1({ DP_addrBus_9 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1074_ (
  .in1({ DP_IN_dout_10, S3264 }),
  .out1({ S3208 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1075_ (
  .in1({ S3118, S3274 }),
  .out1({ S3209 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1363_ (
  .in1({ DP_INC_1_in_10, S32 }),
  .out1({ S3210 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_463_ (
  .in1({ S3210 }),
  .out1({ S3211 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1076_ (
  .in1({ S3211, S3209 }),
  .out1({ S3212 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1077_ (
  .in1({ S3212, S429 }),
  .out1({ S3213 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1364_ (
  .in1({ DP_IMM1_out_10, S430 }),
  .out1({ S3214 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1365_ (
  .in1({ S3214, S3264 }),
  .out1({ S3215 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1078_ (
  .in1({ S3215, S3213 }),
  .out1({ S3216 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1079_ (
  .in1({ S3216, S3208 }),
  .out1({ DP_addrBus_10 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1080_ (
  .in1({ DP_IN_dout_11, S3264 }),
  .out1({ S3217 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1081_ (
  .in1({ S3118, S3275 }),
  .out1({ S3218 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1366_ (
  .in1({ DP_INC_1_in_11, S33 }),
  .out1({ S3219 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_464_ (
  .in1({ S3219 }),
  .out1({ S3220 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1082_ (
  .in1({ S3220, S3218 }),
  .out1({ S3221 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1083_ (
  .in1({ S3221, S431 }),
  .out1({ S3222 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1367_ (
  .in1({ DP_IMM1_out_11, S432 }),
  .out1({ S3223 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1368_ (
  .in1({ S3223, S3264 }),
  .out1({ S3224 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1084_ (
  .in1({ S3224, S3222 }),
  .out1({ S3225 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1085_ (
  .in1({ S3225, S3217 }),
  .out1({ DP_addrBus_11 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1086_ (
  .in1({ DP_IN_dout_12, S3264 }),
  .out1({ S3226 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1087_ (
  .in1({ S3118, S3276 }),
  .out1({ S3227 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1369_ (
  .in1({ DP_INC_1_in_12, S34 }),
  .out1({ S3228 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_465_ (
  .in1({ S3228 }),
  .out1({ S3229 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1088_ (
  .in1({ S3229, S3227 }),
  .out1({ S3230 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1089_ (
  .in1({ S3230, S433 }),
  .out1({ S3231 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1370_ (
  .in1({ DP_IMM1_out_12, S434 }),
  .out1({ S3232 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1371_ (
  .in1({ S3232, S3264 }),
  .out1({ S3233 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1090_ (
  .in1({ S3233, S3231 }),
  .out1({ S3234 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1091_ (
  .in1({ S3234, S3226 }),
  .out1({ DP_addrBus_12 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1092_ (
  .in1({ DP_IN_dout_13, S3264 }),
  .out1({ S3235 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1093_ (
  .in1({ S3118, S3114 }),
  .out1({ S3236 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1372_ (
  .in1({ DP_INC_1_in_13, S35 }),
  .out1({ S3237 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_466_ (
  .in1({ S3237 }),
  .out1({ S3238 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1094_ (
  .in1({ S3238, S3236 }),
  .out1({ S3239 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1095_ (
  .in1({ S3239, S435 }),
  .out1({ S3240 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1373_ (
  .in1({ DP_IMM1_out_13, S436 }),
  .out1({ S3241 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1374_ (
  .in1({ S3241, S3264 }),
  .out1({ S3242 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1096_ (
  .in1({ S3242, S3240 }),
  .out1({ S3243 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1097_ (
  .in1({ S3243, S3235 }),
  .out1({ DP_addrBus_13 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1098_ (
  .in1({ DP_IN_dout_14, S3264 }),
  .out1({ S3244 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1099_ (
  .in1({ S3118, S3115 }),
  .out1({ S3245 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1375_ (
  .in1({ DP_INC_1_in_14, S36 }),
  .out1({ S3246 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_467_ (
  .in1({ S3246 }),
  .out1({ S3247 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1100_ (
  .in1({ S3247, S3245 }),
  .out1({ S3248 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1101_ (
  .in1({ S3248, S437 }),
  .out1({ S3249 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1376_ (
  .in1({ DP_IMM1_out_14, S438 }),
  .out1({ S3250 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1377_ (
  .in1({ S3250, S3264 }),
  .out1({ S3251 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1102_ (
  .in1({ S3251, S3249 }),
  .out1({ S3252 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1103_ (
  .in1({ S3252, S3244 }),
  .out1({ DP_addrBus_14 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1104_ (
  .in1({ DP_IN_dout_15, S3264 }),
  .out1({ S3253 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1105_ (
  .in1({ S3118, S3116 }),
  .out1({ S3254 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1378_ (
  .in1({ DP_INC_1_in_15, S37 }),
  .out1({ S3255 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_468_ (
  .in1({ S3255 }),
  .out1({ S3256 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1106_ (
  .in1({ S3256, S3254 }),
  .out1({ S3257 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1107_ (
  .in1({ S3257, S439 }),
  .out1({ S3258 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1379_ (
  .in1({ DP_IMM1_out_15, S440 }),
  .out1({ S3259 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1380_ (
  .in1({ S3259, S3264 }),
  .out1({ S3260 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1108_ (
  .in1({ S3260, S3258 }),
  .out1({ S3261 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1109_ (
  .in1({ S3261, S3253 }),
  .out1({ DP_addrBus_15 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_469_ (
  .in1({ S441 }),
  .out1({ S3277 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1110_ (
  .in1({ S442, S3277 }),
  .out1({ S3278 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1381_ (
  .in1({ S3278, DP_INC_2_in_0 }),
  .out1({ S3279 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1382_ (
  .in1({ S443, DP_IMM1_out_0 }),
  .out1({ S3280 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1383_ (
  .in1({ S3280, S3279 }),
  .out1({ DP_LGU1_in1_0 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1384_ (
  .in1({ S3278, DP_INC_2_in_1 }),
  .out1({ S3281 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1385_ (
  .in1({ DP_IMM1_out_1, S444 }),
  .out1({ S3282 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1386_ (
  .in1({ S3282, S3281 }),
  .out1({ DP_LGU1_in1_1 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1387_ (
  .in1({ S3278, DP_INC_2_in_2 }),
  .out1({ S3283 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1388_ (
  .in1({ DP_IMM1_out_2, S445 }),
  .out1({ S3284 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1389_ (
  .in1({ S3284, S3283 }),
  .out1({ DP_LGU1_in1_2 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1390_ (
  .in1({ S3278, DP_INC_2_in_3 }),
  .out1({ S3285 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1391_ (
  .in1({ DP_IMM1_out_3, S446 }),
  .out1({ S3286 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1392_ (
  .in1({ S3286, S3285 }),
  .out1({ DP_LGU1_in1_3 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1393_ (
  .in1({ S3278, DP_INC_2_in_4 }),
  .out1({ S3287 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1394_ (
  .in1({ DP_IMM1_out_4, S447 }),
  .out1({ S3288 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1395_ (
  .in1({ S3288, S3287 }),
  .out1({ DP_LGU1_in1_4 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1396_ (
  .in1({ S3278, DP_INC_2_in_5 }),
  .out1({ S3289 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1397_ (
  .in1({ DP_IMM1_out_5, S448 }),
  .out1({ S3290 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1398_ (
  .in1({ S3290, S3289 }),
  .out1({ DP_LGU1_in1_5 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1399_ (
  .in1({ S3278, DP_INC_2_in_6 }),
  .out1({ S3291 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1400_ (
  .in1({ DP_IMM1_out_6, S449 }),
  .out1({ S3292 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1401_ (
  .in1({ S3292, S3291 }),
  .out1({ DP_LGU1_in1_6 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1402_ (
  .in1({ S3278, DP_INC_2_in_7 }),
  .out1({ S3293 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1403_ (
  .in1({ DP_IMM1_out_7, S450 }),
  .out1({ S3294 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1404_ (
  .in1({ S3294, S3293 }),
  .out1({ DP_LGU1_in1_7 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1405_ (
  .in1({ S3278, DP_INC_2_in_8 }),
  .out1({ S3295 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1406_ (
  .in1({ DP_IMM1_out_8, S451 }),
  .out1({ S3296 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1407_ (
  .in1({ S3296, S3295 }),
  .out1({ DP_LGU1_in1_8 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1408_ (
  .in1({ S3278, DP_INC_2_in_9 }),
  .out1({ S3297 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1409_ (
  .in1({ DP_IMM1_out_9, S452 }),
  .out1({ S3298 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1410_ (
  .in1({ S3298, S3297 }),
  .out1({ DP_LGU1_in1_9 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1411_ (
  .in1({ S3278, DP_INC_2_in_10 }),
  .out1({ S3299 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1412_ (
  .in1({ DP_IMM1_out_10, S453 }),
  .out1({ S3300 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1413_ (
  .in1({ S3300, S3299 }),
  .out1({ DP_LGU1_in1_10 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1414_ (
  .in1({ S3278, DP_INC_2_in_11 }),
  .out1({ S3301 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1415_ (
  .in1({ DP_IMM1_out_11, S454 }),
  .out1({ S3302 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1416_ (
  .in1({ S3302, S3301 }),
  .out1({ DP_LGU1_in1_11 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1417_ (
  .in1({ S3278, DP_INC_2_in_12 }),
  .out1({ S3303 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1418_ (
  .in1({ DP_IMM1_out_12, S455 }),
  .out1({ S3304 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1419_ (
  .in1({ S3304, S3303 }),
  .out1({ DP_LGU1_in1_12 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1420_ (
  .in1({ S3278, DP_INC_2_in_13 }),
  .out1({ S3305 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1421_ (
  .in1({ DP_IMM1_out_13, S456 }),
  .out1({ S3306 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1422_ (
  .in1({ S3306, S3305 }),
  .out1({ DP_LGU1_in1_13 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1423_ (
  .in1({ S3278, DP_INC_2_in_14 }),
  .out1({ S3307 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1424_ (
  .in1({ DP_IMM1_out_14, S457 }),
  .out1({ S3308 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1425_ (
  .in1({ S3308, S3307 }),
  .out1({ DP_LGU1_in1_14 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1426_ (
  .in1({ S3278, DP_INC_2_in_15 }),
  .out1({ S3309 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1427_ (
  .in1({ DP_IMM1_out_15, S458 }),
  .out1({ S3310 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1428_ (
  .in1({ S3310, S3309 }),
  .out1({ DP_LGU1_in1_15 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_470_ (
  .in1({ S459 }),
  .out1({ S3311 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1111_ (
  .in1({ S460, S3311 }),
  .out1({ S3312 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1429_ (
  .in1({ S3312, DP_LGU1_in1_0 }),
  .out1({ S3313 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1430_ (
  .in1({ S461, S38 }),
  .out1({ S3314 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1431_ (
  .in1({ S3314, S3313 }),
  .out1({ DP_ARU1_in1_0 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1432_ (
  .in1({ S3312, DP_LGU1_in1_1 }),
  .out1({ S3315 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1433_ (
  .in1({ S463, S462 }),
  .out1({ S3316 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1434_ (
  .in1({ S3316, S3315 }),
  .out1({ DP_ARU1_in1_1 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1435_ (
  .in1({ S3312, DP_LGU1_in1_2 }),
  .out1({ S3317 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1436_ (
  .in1({ S465, S464 }),
  .out1({ S3318 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1437_ (
  .in1({ S3318, S3317 }),
  .out1({ DP_ARU1_in1_2 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1438_ (
  .in1({ S3312, DP_LGU1_in1_3 }),
  .out1({ S3319 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1439_ (
  .in1({ S467, S466 }),
  .out1({ S3320 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1440_ (
  .in1({ S3320, S3319 }),
  .out1({ DP_ARU1_in1_3 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1441_ (
  .in1({ S3312, DP_LGU1_in1_4 }),
  .out1({ S3321 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1442_ (
  .in1({ S469, S468 }),
  .out1({ S3322 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1443_ (
  .in1({ S3322, S3321 }),
  .out1({ DP_ARU1_in1_4 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1444_ (
  .in1({ S3312, DP_LGU1_in1_5 }),
  .out1({ S3323 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1445_ (
  .in1({ S471, S470 }),
  .out1({ S3324 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1446_ (
  .in1({ S3324, S3323 }),
  .out1({ DP_ARU1_in1_5 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1447_ (
  .in1({ S3312, DP_LGU1_in1_6 }),
  .out1({ S3325 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1448_ (
  .in1({ S473, S472 }),
  .out1({ S3326 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1449_ (
  .in1({ S3326, S3325 }),
  .out1({ DP_ARU1_in1_6 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1450_ (
  .in1({ S3312, DP_LGU1_in1_7 }),
  .out1({ S3327 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1451_ (
  .in1({ S475, S474 }),
  .out1({ S3328 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1452_ (
  .in1({ S3328, S3327 }),
  .out1({ DP_ARU1_in1_7 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1453_ (
  .in1({ S3312, DP_LGU1_in1_8 }),
  .out1({ S3329 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1454_ (
  .in1({ S477, S476 }),
  .out1({ S3330 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1455_ (
  .in1({ S3330, S3329 }),
  .out1({ DP_ARU1_in1_8 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1456_ (
  .in1({ S3312, DP_LGU1_in1_9 }),
  .out1({ S3331 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1457_ (
  .in1({ S479, S478 }),
  .out1({ S3332 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1458_ (
  .in1({ S3332, S3331 }),
  .out1({ DP_ARU1_in1_9 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1459_ (
  .in1({ S3312, DP_LGU1_in1_10 }),
  .out1({ S3333 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1460_ (
  .in1({ S481, S480 }),
  .out1({ S3334 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1461_ (
  .in1({ S3334, S3333 }),
  .out1({ DP_ARU1_in1_10 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1462_ (
  .in1({ S3312, DP_LGU1_in1_11 }),
  .out1({ S3335 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1463_ (
  .in1({ S483, S482 }),
  .out1({ S3336 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1464_ (
  .in1({ S3336, S3335 }),
  .out1({ DP_ARU1_in1_11 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1465_ (
  .in1({ S3312, DP_LGU1_in1_12 }),
  .out1({ S3337 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1466_ (
  .in1({ S485, S484 }),
  .out1({ S3338 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1467_ (
  .in1({ S3338, S3337 }),
  .out1({ DP_ARU1_in1_12 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1468_ (
  .in1({ S3312, DP_LGU1_in1_13 }),
  .out1({ S3339 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1469_ (
  .in1({ S487, S486 }),
  .out1({ S3340 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1470_ (
  .in1({ S3340, S3339 }),
  .out1({ DP_ARU1_in1_13 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1471_ (
  .in1({ S3312, DP_LGU1_in1_14 }),
  .out1({ S3341 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1472_ (
  .in1({ S489, S488 }),
  .out1({ S3342 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1473_ (
  .in1({ S3342, S3341 }),
  .out1({ DP_ARU1_in1_14 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1474_ (
  .in1({ S3312, DP_LGU1_in1_15 }),
  .out1({ S3343 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1475_ (
  .in1({ S491, S490 }),
  .out1({ S3344 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1476_ (
  .in1({ S3344, S3343 }),
  .out1({ DP_ARU1_in1_15 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_471_ (
  .in1({ S492 }),
  .out1({ S3345 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1112_ (
  .in1({ S493, S3345 }),
  .out1({ S3346 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1477_ (
  .in1({ S3346, DP_IMM1_out_0 }),
  .out1({ S3347 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1478_ (
  .in1({ S494, DP_INC_1_in_12 }),
  .out1({ S3348 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1479_ (
  .in1({ S3348, S3347 }),
  .out1({ DP_OF_din_0 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1480_ (
  .in1({ S3346, DP_IMM1_out_1 }),
  .out1({ S3349 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1481_ (
  .in1({ DP_INC_1_in_13, S495 }),
  .out1({ S3350 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1482_ (
  .in1({ S3350, S3349 }),
  .out1({ DP_OF_din_1 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1483_ (
  .in1({ S3346, DP_IMM1_out_2 }),
  .out1({ S3351 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1484_ (
  .in1({ DP_INC_1_in_14, S496 }),
  .out1({ S3352 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1485_ (
  .in1({ S3352, S3351 }),
  .out1({ DP_OF_din_2 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1486_ (
  .in1({ S3346, DP_IMM1_out_3 }),
  .out1({ S3353 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1487_ (
  .in1({ DP_INC_1_in_15, S497 }),
  .out1({ S3354 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1488_ (
  .in1({ S3354, S3353 }),
  .out1({ DP_OF_din_3 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_472_ (
  .in1({ S498 }),
  .out1({ S3360 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1113_ (
  .in1({ S499, S3360 }),
  .out1({ S3355 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1489_ (
  .in1({ S3355, S39 }),
  .out1({ S3356 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1490_ (
  .in1({ S501, S500 }),
  .out1({ S3357 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1491_ (
  .in1({ S3357, S3356 }),
  .out1({ DP_INC_1_inc_value_0 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1492_ (
  .in1({ S3355, S502 }),
  .out1({ S3358 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1493_ (
  .in1({ S40, S503 }),
  .out1({ S3359 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1494_ (
  .in1({ S3359, S3358 }),
  .out1({ DP_INC_1_inc_value_1 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_506_ (
  .in1({ DP_addrBus_0 }),
  .out1({ addrBus[0] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_507_ (
  .in1({ DP_addrBus_1 }),
  .out1({ addrBus[1] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_508_ (
  .in1({ DP_addrBus_10 }),
  .out1({ addrBus[10] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_509_ (
  .in1({ DP_addrBus_11 }),
  .out1({ addrBus[11] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_510_ (
  .in1({ DP_addrBus_12 }),
  .out1({ addrBus[12] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_511_ (
  .in1({ DP_addrBus_13 }),
  .out1({ addrBus[13] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_512_ (
  .in1({ DP_addrBus_14 }),
  .out1({ addrBus[14] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_513_ (
  .in1({ DP_addrBus_15 }),
  .out1({ addrBus[15] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_514_ (
  .in1({ DP_addrBus_2 }),
  .out1({ addrBus[2] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_515_ (
  .in1({ DP_addrBus_3 }),
  .out1({ addrBus[3] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_516_ (
  .in1({ DP_addrBus_4 }),
  .out1({ addrBus[4] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_517_ (
  .in1({ DP_addrBus_5 }),
  .out1({ addrBus[5] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_518_ (
  .in1({ DP_addrBus_6 }),
  .out1({ addrBus[6] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_519_ (
  .in1({ DP_addrBus_7 }),
  .out1({ addrBus[7] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_520_ (
  .in1({ DP_addrBus_8 }),
  .out1({ addrBus[8] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_521_ (
  .in1({ DP_addrBus_9 }),
  .out1({ addrBus[9] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_522_ (
  .in1({ clk }),
  .out1({ CU_clk })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_523_ (
  .in1({ dataBus_in[0] }),
  .out1({ DP_INC_2_in_0 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_524_ (
  .in1({ dataBus_in[1] }),
  .out1({ DP_INC_2_in_1 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_525_ (
  .in1({ dataBus_in[10] }),
  .out1({ DP_INC_2_in_10 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_526_ (
  .in1({ dataBus_in[11] }),
  .out1({ DP_INC_2_in_11 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_527_ (
  .in1({ dataBus_in[12] }),
  .out1({ DP_INC_2_in_12 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_528_ (
  .in1({ dataBus_in[13] }),
  .out1({ DP_INC_2_in_13 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_529_ (
  .in1({ dataBus_in[14] }),
  .out1({ DP_INC_2_in_14 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_530_ (
  .in1({ dataBus_in[15] }),
  .out1({ DP_INC_2_in_15 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_531_ (
  .in1({ dataBus_in[2] }),
  .out1({ DP_INC_2_in_2 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_532_ (
  .in1({ dataBus_in[3] }),
  .out1({ DP_INC_2_in_3 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_533_ (
  .in1({ dataBus_in[4] }),
  .out1({ DP_INC_2_in_4 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_534_ (
  .in1({ dataBus_in[5] }),
  .out1({ DP_INC_2_in_5 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_535_ (
  .in1({ dataBus_in[6] }),
  .out1({ DP_INC_2_in_6 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_536_ (
  .in1({ dataBus_in[7] }),
  .out1({ DP_INC_2_in_7 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_537_ (
  .in1({ dataBus_in[8] }),
  .out1({ DP_INC_2_in_8 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_538_ (
  .in1({ dataBus_in[9] }),
  .out1({ DP_INC_2_in_9 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_539_ (
  .in1({ DP_TriBuff_out_0 }),
  .out1({ dataBus_out[0] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_540_ (
  .in1({ DP_TriBuff_out_1 }),
  .out1({ dataBus_out[1] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_541_ (
  .in1({ DP_TriBuff_out_10 }),
  .out1({ dataBus_out[10] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_542_ (
  .in1({ DP_TriBuff_out_11 }),
  .out1({ dataBus_out[11] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_543_ (
  .in1({ DP_TriBuff_out_12 }),
  .out1({ dataBus_out[12] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_544_ (
  .in1({ DP_TriBuff_out_13 }),
  .out1({ dataBus_out[13] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_545_ (
  .in1({ DP_TriBuff_out_14 }),
  .out1({ dataBus_out[14] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_546_ (
  .in1({ DP_TriBuff_out_15 }),
  .out1({ dataBus_out[15] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_547_ (
  .in1({ DP_TriBuff_out_2 }),
  .out1({ dataBus_out[2] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_548_ (
  .in1({ DP_TriBuff_out_3 }),
  .out1({ dataBus_out[3] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_549_ (
  .in1({ DP_TriBuff_out_4 }),
  .out1({ dataBus_out[4] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_550_ (
  .in1({ DP_TriBuff_out_5 }),
  .out1({ dataBus_out[5] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_551_ (
  .in1({ DP_TriBuff_out_6 }),
  .out1({ dataBus_out[6] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_552_ (
  .in1({ DP_TriBuff_out_7 }),
  .out1({ dataBus_out[7] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_553_ (
  .in1({ DP_TriBuff_out_8 }),
  .out1({ dataBus_out[8] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_554_ (
  .in1({ DP_TriBuff_out_9 }),
  .out1({ dataBus_out[9] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_555_ (
  .in1({ S41 }),
  .out1({ readMEM })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_556_ (
  .in1({ rst }),
  .out1({ CU_rst })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_557_ (
  .in1({ S504 }),
  .out1({ writeMEM })
);

endmodule