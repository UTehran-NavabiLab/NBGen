LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

ENTITY Circuit432 IS
    PORT (
        in4 : IN STD_LOGIC;
        in17 : IN STD_LOGIC;
        in30 : IN STD_LOGIC;
        in43 : IN STD_LOGIC;
        in56 : IN STD_LOGIC;
        in69 : IN STD_LOGIC;
        in82 : IN STD_LOGIC;
        in95 : IN STD_LOGIC;
        in108 : IN STD_LOGIC;
        in1 : IN STD_LOGIC;
        in11 : IN STD_LOGIC;
        in24 : IN STD_LOGIC;
        in37 : IN STD_LOGIC;
        in50 : IN STD_LOGIC;
        in63 : IN STD_LOGIC;
        in76 : IN STD_LOGIC;
        in89 : IN STD_LOGIC;
        in102 : IN STD_LOGIC;
        in8 : IN STD_LOGIC;
        in21 : IN STD_LOGIC;
        in34 : IN STD_LOGIC;
        in47 : IN STD_LOGIC;
        in60 : IN STD_LOGIC;
        in73 : IN STD_LOGIC;
        in86 : IN STD_LOGIC;
        in99 : IN STD_LOGIC;
        in112 : IN STD_LOGIC;
        in14 : IN STD_LOGIC;
        in27 : IN STD_LOGIC;
        in40 : IN STD_LOGIC;
        in53 : IN STD_LOGIC;
        in66 : IN STD_LOGIC;
        in79 : IN STD_LOGIC;
        in92 : IN STD_LOGIC;
        in105 : IN STD_LOGIC;
        in115 : IN STD_LOGIC;
        out223 : OUT STD_LOGIC;
        out329 : OUT STD_LOGIC;
        out370 : OUT STD_LOGIC;
        out421 : OUT STD_LOGIC;
        out430 : OUT STD_LOGIC;
        out431 : OUT STD_LOGIC;
        out432 : OUT STD_LOGIC);
END ENTITY Circuit432;

ARCHITECTURE arch OF Circuit432 IS
    SIGNAL Ckt432_I_0 : STD_LOGIC;
    SIGNAL Ckt432_I_1 : STD_LOGIC;
    SIGNAL Ckt432_I_2 : STD_LOGIC;
    SIGNAL Ckt432_I_3 : STD_LOGIC;
    SIGNAL Ckt432_I_4 : STD_LOGIC;
    SIGNAL Ckt432_I_5 : STD_LOGIC;
    SIGNAL Ckt432_I_6 : STD_LOGIC;
    SIGNAL Ckt432_I_7 : STD_LOGIC;
    SIGNAL Ckt432_I_8 : STD_LOGIC;
    SIGNAL Ckt432_M1_X1_0 : STD_LOGIC;
    SIGNAL Ckt432_M1_X1_1 : STD_LOGIC;
    SIGNAL Ckt432_M1_X1_2 : STD_LOGIC;
    SIGNAL Ckt432_M1_X1_3 : STD_LOGIC;
    SIGNAL Ckt432_M1_X1_4 : STD_LOGIC;
    SIGNAL Ckt432_M1_X1_5 : STD_LOGIC;
    SIGNAL Ckt432_M1_X1_6 : STD_LOGIC;
    SIGNAL Ckt432_M1_X1_7 : STD_LOGIC;
    SIGNAL Ckt432_M1_X1_8 : STD_LOGIC;
    SIGNAL Ckt432_M1_n1 : STD_LOGIC;
    SIGNAL Ckt432_M1_n10 : STD_LOGIC;
    SIGNAL Ckt432_M1_n11 : STD_LOGIC;
    SIGNAL Ckt432_M1_n12 : STD_LOGIC;
    SIGNAL Ckt432_M1_n13 : STD_LOGIC;
    SIGNAL Ckt432_M1_n14 : STD_LOGIC;
    SIGNAL Ckt432_M1_n15 : STD_LOGIC;
    SIGNAL Ckt432_M1_n2 : STD_LOGIC;
    SIGNAL Ckt432_M1_n3 : STD_LOGIC;
    SIGNAL Ckt432_M1_n4 : STD_LOGIC;
    SIGNAL Ckt432_M1_n5 : STD_LOGIC;
    SIGNAL Ckt432_M1_n6 : STD_LOGIC;
    SIGNAL Ckt432_M1_n7 : STD_LOGIC;
    SIGNAL Ckt432_M1_n8 : STD_LOGIC;
    SIGNAL Ckt432_M1_n9 : STD_LOGIC;
    SIGNAL Ckt432_M2_X2_0 : STD_LOGIC;
    SIGNAL Ckt432_M2_X2_1 : STD_LOGIC;
    SIGNAL Ckt432_M2_X2_2 : STD_LOGIC;
    SIGNAL Ckt432_M2_X2_3 : STD_LOGIC;
    SIGNAL Ckt432_M2_X2_4 : STD_LOGIC;
    SIGNAL Ckt432_M2_X2_5 : STD_LOGIC;
    SIGNAL Ckt432_M2_X2_6 : STD_LOGIC;
    SIGNAL Ckt432_M2_X2_7 : STD_LOGIC;
    SIGNAL Ckt432_M2_X2_8 : STD_LOGIC;
    SIGNAL Ckt432_M2_n1 : STD_LOGIC;
    SIGNAL Ckt432_M2_n10 : STD_LOGIC;
    SIGNAL Ckt432_M2_n11 : STD_LOGIC;
    SIGNAL Ckt432_M2_n12 : STD_LOGIC;
    SIGNAL Ckt432_M2_n13 : STD_LOGIC;
    SIGNAL Ckt432_M2_n14 : STD_LOGIC;
    SIGNAL Ckt432_M2_n15 : STD_LOGIC;
    SIGNAL Ckt432_M2_n16 : STD_LOGIC;
    SIGNAL Ckt432_M2_n17 : STD_LOGIC;
    SIGNAL Ckt432_M2_n18 : STD_LOGIC;
    SIGNAL Ckt432_M2_n19 : STD_LOGIC;
    SIGNAL Ckt432_M2_n2 : STD_LOGIC;
    SIGNAL Ckt432_M2_n20 : STD_LOGIC;
    SIGNAL Ckt432_M2_n3 : STD_LOGIC;
    SIGNAL Ckt432_M2_n4 : STD_LOGIC;
    SIGNAL Ckt432_M2_n5 : STD_LOGIC;
    SIGNAL Ckt432_M2_n6 : STD_LOGIC;
    SIGNAL Ckt432_M2_n7 : STD_LOGIC;
    SIGNAL Ckt432_M2_n8 : STD_LOGIC;
    SIGNAL Ckt432_M2_n9 : STD_LOGIC;
    SIGNAL Ckt432_M3_n1 : STD_LOGIC;
    SIGNAL Ckt432_M3_n10 : STD_LOGIC;
    SIGNAL Ckt432_M3_n11 : STD_LOGIC;
    SIGNAL Ckt432_M3_n12 : STD_LOGIC;
    SIGNAL Ckt432_M3_n13 : STD_LOGIC;
    SIGNAL Ckt432_M3_n14 : STD_LOGIC;
    SIGNAL Ckt432_M3_n15 : STD_LOGIC;
    SIGNAL Ckt432_M3_n16 : STD_LOGIC;
    SIGNAL Ckt432_M3_n17 : STD_LOGIC;
    SIGNAL Ckt432_M3_n18 : STD_LOGIC;
    SIGNAL Ckt432_M3_n19 : STD_LOGIC;
    SIGNAL Ckt432_M3_n2 : STD_LOGIC;
    SIGNAL Ckt432_M3_n20 : STD_LOGIC;
    SIGNAL Ckt432_M3_n3 : STD_LOGIC;
    SIGNAL Ckt432_M3_n4 : STD_LOGIC;
    SIGNAL Ckt432_M3_n5 : STD_LOGIC;
    SIGNAL Ckt432_M3_n6 : STD_LOGIC;
    SIGNAL Ckt432_M3_n7 : STD_LOGIC;
    SIGNAL Ckt432_M3_n8 : STD_LOGIC;
    SIGNAL Ckt432_M3_n9 : STD_LOGIC;
    SIGNAL Ckt432_M4_n1 : STD_LOGIC;
    SIGNAL Ckt432_M4_n10 : STD_LOGIC;
    SIGNAL Ckt432_M4_n11 : STD_LOGIC;
    SIGNAL Ckt432_M4_n12 : STD_LOGIC;
    SIGNAL Ckt432_M4_n13 : STD_LOGIC;
    SIGNAL Ckt432_M4_n14 : STD_LOGIC;
    SIGNAL Ckt432_M4_n15 : STD_LOGIC;
    SIGNAL Ckt432_M4_n16 : STD_LOGIC;
    SIGNAL Ckt432_M4_n17 : STD_LOGIC;
    SIGNAL Ckt432_M4_n18 : STD_LOGIC;
    SIGNAL Ckt432_M4_n2 : STD_LOGIC;
    SIGNAL Ckt432_M4_n3 : STD_LOGIC;
    SIGNAL Ckt432_M4_n4 : STD_LOGIC;
    SIGNAL Ckt432_M4_n5 : STD_LOGIC;
    SIGNAL Ckt432_M4_n6 : STD_LOGIC;
    SIGNAL Ckt432_M4_n7 : STD_LOGIC;
    SIGNAL Ckt432_M4_n8 : STD_LOGIC;
    SIGNAL Ckt432_M4_n9 : STD_LOGIC;
    SIGNAL Ckt432_M5_n1 : STD_LOGIC;
    SIGNAL Ckt432_M5_n2 : STD_LOGIC;
    SIGNAL Ckt432_M5_n3 : STD_LOGIC;
    SIGNAL Ckt432_M5_n4 : STD_LOGIC;
    SIGNAL Ckt432_M5_n5 : STD_LOGIC;
    SIGNAL Ckt432_M5_n6 : STD_LOGIC;
    SIGNAL Ckt432_M5_n7 : STD_LOGIC;
    SIGNAL Ckt432_M5_n8 : STD_LOGIC;
    SIGNAL Ckt432_M5_n9 : STD_LOGIC;

BEGIN
OAI21_X1_1: ENTITY WORK.OAI21_X1
    PORT MAP (
        A => out223,
        B1 => in1,
        B2 => Ckt432_M1_n1,
        ZN => Ckt432_M1_X1_8
    );
OR2_X1_1: ENTITY WORK.OR2_X1
    PORT MAP (
        A1 => Ckt432_M1_n10,
        A2 => Ckt432_M1_n11,
        ZN => out223
    );
OAI221_X1_1: ENTITY WORK.OAI221_X1
    PORT MAP (
        A => Ckt432_M1_n12,
        B1 => Ckt432_M1_n6,
        B2 => in63,
        C1 => Ckt432_M1_n5,
        C2 => in50,
        ZN => Ckt432_M1_n11
    );
INV_X1_1: ENTITY WORK.INV_X1
    PORT MAP (
        A => Ckt432_M1_n13,
        ZN => Ckt432_M1_n12
    );
OAI222_X1_1: ENTITY WORK.OAI222_X1
    PORT MAP (
        A1 => in89,
        A2 => Ckt432_M1_n8,
        B1 => in102,
        B2 => Ckt432_M1_n9,
        C1 => in76,
        C2 => Ckt432_M1_n7,
        ZN => Ckt432_M1_n13
    );
INV_X1_2: ENTITY WORK.INV_X1
    PORT MAP (
        A => in82,
        ZN => Ckt432_M1_n7
    );
INV_X1_3: ENTITY WORK.INV_X1
    PORT MAP (
        A => in108,
        ZN => Ckt432_M1_n9
    );
INV_X1_4: ENTITY WORK.INV_X1
    PORT MAP (
        A => in95,
        ZN => Ckt432_M1_n8
    );
INV_X1_5: ENTITY WORK.INV_X1
    PORT MAP (
        A => in56,
        ZN => Ckt432_M1_n5
    );
INV_X1_6: ENTITY WORK.INV_X1
    PORT MAP (
        A => in69,
        ZN => Ckt432_M1_n6
    );
OAI221_X1_2: ENTITY WORK.OAI221_X1
    PORT MAP (
        A => Ckt432_M1_n14,
        B1 => Ckt432_M1_n2,
        B2 => in11,
        C1 => Ckt432_M1_n1,
        C2 => in1,
        ZN => Ckt432_M1_n10
    );
OAI21_X1_2: ENTITY WORK.OAI21_X1
    PORT MAP (
        A => out223,
        B1 => in11,
        B2 => Ckt432_M1_n2,
        ZN => Ckt432_M1_X1_7
    );
INV_X1_7: ENTITY WORK.INV_X1
    PORT MAP (
        A => Ckt432_M1_n15,
        ZN => Ckt432_M1_n14
    );
OAI22_X1_1: ENTITY WORK.OAI22_X1
    PORT MAP (
        A1 => in24,
        A2 => Ckt432_M1_n3,
        B1 => in37,
        B2 => Ckt432_M1_n4,
        ZN => Ckt432_M1_n15
    );
INV_X1_8: ENTITY WORK.INV_X1
    PORT MAP (
        A => in43,
        ZN => Ckt432_M1_n4
    );
INV_X1_9: ENTITY WORK.INV_X1
    PORT MAP (
        A => in30,
        ZN => Ckt432_M1_n3
    );
INV_X1_10: ENTITY WORK.INV_X1
    PORT MAP (
        A => in4,
        ZN => Ckt432_M1_n1
    );
INV_X1_11: ENTITY WORK.INV_X1
    PORT MAP (
        A => in17,
        ZN => Ckt432_M1_n2
    );
OAI21_X1_3: ENTITY WORK.OAI21_X1
    PORT MAP (
        A => out223,
        B1 => in24,
        B2 => Ckt432_M1_n3,
        ZN => Ckt432_M1_X1_6
    );
OAI21_X1_4: ENTITY WORK.OAI21_X1
    PORT MAP (
        A => out223,
        B1 => in37,
        B2 => Ckt432_M1_n4,
        ZN => Ckt432_M1_X1_5
    );
OAI21_X1_5: ENTITY WORK.OAI21_X1
    PORT MAP (
        A => out223,
        B1 => in50,
        B2 => Ckt432_M1_n5,
        ZN => Ckt432_M1_X1_4
    );
OAI21_X1_6: ENTITY WORK.OAI21_X1
    PORT MAP (
        A => out223,
        B1 => in63,
        B2 => Ckt432_M1_n6,
        ZN => Ckt432_M1_X1_3
    );
OAI21_X1_7: ENTITY WORK.OAI21_X1
    PORT MAP (
        A => out223,
        B1 => in76,
        B2 => Ckt432_M1_n7,
        ZN => Ckt432_M1_X1_2
    );
OAI21_X1_8: ENTITY WORK.OAI21_X1
    PORT MAP (
        A => out223,
        B1 => in89,
        B2 => Ckt432_M1_n8,
        ZN => Ckt432_M1_X1_1
    );
OAI21_X1_9: ENTITY WORK.OAI21_X1
    PORT MAP (
        A => out223,
        B1 => in102,
        B2 => Ckt432_M1_n9,
        ZN => Ckt432_M1_X1_0
    );
NAND2_X1_1: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => out329,
        A2 => Ckt432_M2_n1,
        ZN => Ckt432_M2_X2_8
    );
NAND4_X1_1: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => Ckt432_M2_n5,
        A2 => Ckt432_M2_n4,
        A3 => Ckt432_M2_n10,
        A4 => Ckt432_M2_n11,
        ZN => out329
    );
AND4_X1_1: ENTITY WORK.AND4_X1
    PORT MAP (
        A1 => Ckt432_M2_n6,
        A2 => Ckt432_M2_n7,
        A3 => Ckt432_M2_n8,
        A4 => Ckt432_M2_n9,
        ZN => Ckt432_M2_n11
    );
NAND3_X1_1: ENTITY WORK.NAND3_X1
    PORT MAP (
        A1 => in108,
        A2 => Ckt432_M2_n12,
        A3 => Ckt432_M1_X1_0,
        ZN => Ckt432_M2_n9
    );
INV_X1_12: ENTITY WORK.INV_X1
    PORT MAP (
        A => in112,
        ZN => Ckt432_M2_n12
    );
NAND3_X1_2: ENTITY WORK.NAND3_X1
    PORT MAP (
        A1 => in95,
        A2 => Ckt432_M2_n13,
        A3 => Ckt432_M1_X1_1,
        ZN => Ckt432_M2_n8
    );
INV_X1_13: ENTITY WORK.INV_X1
    PORT MAP (
        A => in99,
        ZN => Ckt432_M2_n13
    );
NAND3_X1_3: ENTITY WORK.NAND3_X1
    PORT MAP (
        A1 => in82,
        A2 => Ckt432_M2_n14,
        A3 => Ckt432_M1_X1_2,
        ZN => Ckt432_M2_n7
    );
INV_X1_14: ENTITY WORK.INV_X1
    PORT MAP (
        A => in86,
        ZN => Ckt432_M2_n14
    );
NAND3_X1_4: ENTITY WORK.NAND3_X1
    PORT MAP (
        A1 => in69,
        A2 => Ckt432_M2_n15,
        A3 => Ckt432_M1_X1_3,
        ZN => Ckt432_M2_n6
    );
INV_X1_15: ENTITY WORK.INV_X1
    PORT MAP (
        A => in73,
        ZN => Ckt432_M2_n15
    );
NAND2_X1_2: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => out329,
        A2 => Ckt432_M2_n2,
        ZN => Ckt432_M2_X2_7
    );
AND3_X1_1: ENTITY WORK.AND3_X1
    PORT MAP (
        A1 => Ckt432_M2_n3,
        A2 => Ckt432_M2_n1,
        A3 => Ckt432_M2_n2,
        ZN => Ckt432_M2_n10
    );
NAND3_X1_5: ENTITY WORK.NAND3_X1
    PORT MAP (
        A1 => in17,
        A2 => Ckt432_M2_n16,
        A3 => Ckt432_M1_X1_7,
        ZN => Ckt432_M2_n2
    );
INV_X1_16: ENTITY WORK.INV_X1
    PORT MAP (
        A => in21,
        ZN => Ckt432_M2_n16
    );
NAND3_X1_6: ENTITY WORK.NAND3_X1
    PORT MAP (
        A1 => in4,
        A2 => Ckt432_M2_n17,
        A3 => Ckt432_M1_X1_8,
        ZN => Ckt432_M2_n1
    );
INV_X1_17: ENTITY WORK.INV_X1
    PORT MAP (
        A => in8,
        ZN => Ckt432_M2_n17
    );
NAND3_X1_7: ENTITY WORK.NAND3_X1
    PORT MAP (
        A1 => in30,
        A2 => Ckt432_M2_n18,
        A3 => Ckt432_M1_X1_6,
        ZN => Ckt432_M2_n3
    );
INV_X1_18: ENTITY WORK.INV_X1
    PORT MAP (
        A => in34,
        ZN => Ckt432_M2_n18
    );
NAND3_X1_8: ENTITY WORK.NAND3_X1
    PORT MAP (
        A1 => in43,
        A2 => Ckt432_M2_n19,
        A3 => Ckt432_M1_X1_5,
        ZN => Ckt432_M2_n4
    );
INV_X1_19: ENTITY WORK.INV_X1
    PORT MAP (
        A => in47,
        ZN => Ckt432_M2_n19
    );
NAND3_X1_9: ENTITY WORK.NAND3_X1
    PORT MAP (
        A1 => in56,
        A2 => Ckt432_M2_n20,
        A3 => Ckt432_M1_X1_4,
        ZN => Ckt432_M2_n5
    );
NAND2_X1_3: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => out329,
        A2 => Ckt432_M2_n3,
        ZN => Ckt432_M2_X2_6
    );
INV_X1_20: ENTITY WORK.INV_X1
    PORT MAP (
        A => in60,
        ZN => Ckt432_M2_n20
    );
NAND2_X1_4: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => out329,
        A2 => Ckt432_M2_n4,
        ZN => Ckt432_M2_X2_5
    );
NAND2_X1_5: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => out329,
        A2 => Ckt432_M2_n5,
        ZN => Ckt432_M2_X2_4
    );
NAND2_X1_6: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => out329,
        A2 => Ckt432_M2_n6,
        ZN => Ckt432_M2_X2_3
    );
NAND2_X1_7: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => out329,
        A2 => Ckt432_M2_n7,
        ZN => Ckt432_M2_X2_2
    );
NAND2_X1_8: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => out329,
        A2 => Ckt432_M2_n8,
        ZN => Ckt432_M2_X2_1
    );
NAND2_X1_9: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => out329,
        A2 => Ckt432_M2_n9,
        ZN => Ckt432_M2_X2_0
    );
NAND4_X1_2: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => Ckt432_M3_n1,
        A2 => Ckt432_M3_n2,
        A3 => Ckt432_M3_n3,
        A4 => Ckt432_M3_n4,
        ZN => out370
    );
INV_X1_21: ENTITY WORK.INV_X1
    PORT MAP (
        A => in14,
        ZN => Ckt432_M3_n12
    );
AND3_X1_2: ENTITY WORK.AND3_X1
    PORT MAP (
        A1 => Ckt432_M3_n13,
        A2 => Ckt432_M3_n14,
        A3 => Ckt432_M3_n15,
        ZN => Ckt432_M3_n3
    );
NAND4_X1_3: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => Ckt432_M2_X2_2,
        A2 => Ckt432_M1_X1_2,
        A3 => in82,
        A4 => Ckt432_M3_n16,
        ZN => Ckt432_M3_n15
    );
INV_X1_22: ENTITY WORK.INV_X1
    PORT MAP (
        A => in92,
        ZN => Ckt432_M3_n16
    );
NAND4_X1_4: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => Ckt432_M2_X2_0,
        A2 => Ckt432_M1_X1_0,
        A3 => in108,
        A4 => Ckt432_M3_n17,
        ZN => Ckt432_M3_n14
    );
INV_X1_23: ENTITY WORK.INV_X1
    PORT MAP (
        A => in115,
        ZN => Ckt432_M3_n17
    );
NAND4_X1_5: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => Ckt432_M2_X2_1,
        A2 => Ckt432_M1_X1_1,
        A3 => in95,
        A4 => Ckt432_M3_n18,
        ZN => Ckt432_M3_n13
    );
INV_X1_24: ENTITY WORK.INV_X1
    PORT MAP (
        A => in105,
        ZN => Ckt432_M3_n18
    );
NAND4_X1_6: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => Ckt432_M2_X2_3,
        A2 => Ckt432_M1_X1_3,
        A3 => in69,
        A4 => Ckt432_M3_n19,
        ZN => Ckt432_M3_n2
    );
INV_X1_25: ENTITY WORK.INV_X1
    PORT MAP (
        A => in79,
        ZN => Ckt432_M3_n19
    );
AND4_X1_2: ENTITY WORK.AND4_X1
    PORT MAP (
        A1 => Ckt432_M3_n5,
        A2 => Ckt432_M3_n6,
        A3 => Ckt432_M3_n7,
        A4 => Ckt432_M3_n8,
        ZN => Ckt432_M3_n4
    );
NAND4_X1_7: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => Ckt432_M2_X2_4,
        A2 => Ckt432_M1_X1_4,
        A3 => in56,
        A4 => Ckt432_M3_n20,
        ZN => Ckt432_M3_n1
    );
INV_X1_26: ENTITY WORK.INV_X1
    PORT MAP (
        A => in66,
        ZN => Ckt432_M3_n20
    );
NAND4_X1_8: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => Ckt432_M2_X2_5,
        A2 => Ckt432_M1_X1_5,
        A3 => in43,
        A4 => Ckt432_M3_n9,
        ZN => Ckt432_M3_n8
    );
INV_X1_27: ENTITY WORK.INV_X1
    PORT MAP (
        A => in53,
        ZN => Ckt432_M3_n9
    );
NAND4_X1_9: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => Ckt432_M2_X2_6,
        A2 => Ckt432_M1_X1_6,
        A3 => in30,
        A4 => Ckt432_M3_n10,
        ZN => Ckt432_M3_n7
    );
INV_X1_28: ENTITY WORK.INV_X1
    PORT MAP (
        A => in40,
        ZN => Ckt432_M3_n10
    );
NAND4_X1_10: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => Ckt432_M2_X2_7,
        A2 => Ckt432_M1_X1_7,
        A3 => in17,
        A4 => Ckt432_M3_n11,
        ZN => Ckt432_M3_n6
    );
INV_X1_29: ENTITY WORK.INV_X1
    PORT MAP (
        A => in27,
        ZN => Ckt432_M3_n11
    );
NAND4_X1_11: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => Ckt432_M2_X2_8,
        A2 => Ckt432_M1_X1_8,
        A3 => in4,
        A4 => Ckt432_M3_n12,
        ZN => Ckt432_M3_n5
    );
NAND3_X1_10: ENTITY WORK.NAND3_X1
    PORT MAP (
        A1 => in4,
        A2 => Ckt432_M4_n1,
        A3 => Ckt432_M4_n2,
        ZN => Ckt432_I_8
    );
NAND3_X1_11: ENTITY WORK.NAND3_X1
    PORT MAP (
        A1 => in43,
        A2 => Ckt432_M4_n7,
        A3 => Ckt432_M4_n8,
        ZN => Ckt432_I_5
    );
AOI22_X1_1: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => in37,
        A2 => out223,
        B1 => in47,
        B2 => out329,
        ZN => Ckt432_M4_n8
    );
NAND2_X1_10: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => in53,
        A2 => out370,
        ZN => Ckt432_M4_n7
    );
NAND3_X1_12: ENTITY WORK.NAND3_X1
    PORT MAP (
        A1 => in56,
        A2 => Ckt432_M4_n9,
        A3 => Ckt432_M4_n10,
        ZN => Ckt432_I_4
    );
AOI22_X1_2: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => in50,
        A2 => out223,
        B1 => in60,
        B2 => out329,
        ZN => Ckt432_M4_n10
    );
NAND2_X1_11: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => in66,
        A2 => out370,
        ZN => Ckt432_M4_n9
    );
NAND3_X1_13: ENTITY WORK.NAND3_X1
    PORT MAP (
        A1 => in69,
        A2 => Ckt432_M4_n11,
        A3 => Ckt432_M4_n12,
        ZN => Ckt432_I_3
    );
AOI22_X1_3: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => in63,
        A2 => out223,
        B1 => in73,
        B2 => out329,
        ZN => Ckt432_M4_n12
    );
NAND2_X1_12: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => in79,
        A2 => out370,
        ZN => Ckt432_M4_n11
    );
NAND3_X1_14: ENTITY WORK.NAND3_X1
    PORT MAP (
        A1 => in82,
        A2 => Ckt432_M4_n13,
        A3 => Ckt432_M4_n14,
        ZN => Ckt432_I_2
    );
AOI22_X1_4: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => out223,
        A2 => in1,
        B1 => out329,
        B2 => in8,
        ZN => Ckt432_M4_n2
    );
AOI22_X1_5: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => in76,
        A2 => out223,
        B1 => in86,
        B2 => out329,
        ZN => Ckt432_M4_n14
    );
NAND2_X1_13: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => in92,
        A2 => out370,
        ZN => Ckt432_M4_n13
    );
NAND3_X1_15: ENTITY WORK.NAND3_X1
    PORT MAP (
        A1 => in95,
        A2 => Ckt432_M4_n15,
        A3 => Ckt432_M4_n16,
        ZN => Ckt432_I_1
    );
AOI22_X1_6: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => in89,
        A2 => out223,
        B1 => in99,
        B2 => out329,
        ZN => Ckt432_M4_n16
    );
NAND2_X1_14: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => in105,
        A2 => out370,
        ZN => Ckt432_M4_n15
    );
NAND3_X1_16: ENTITY WORK.NAND3_X1
    PORT MAP (
        A1 => in108,
        A2 => Ckt432_M4_n17,
        A3 => Ckt432_M4_n18,
        ZN => Ckt432_I_0
    );
AOI22_X1_7: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => in102,
        A2 => out223,
        B1 => in112,
        B2 => out329,
        ZN => Ckt432_M4_n18
    );
NAND2_X1_15: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => in115,
        A2 => out370,
        ZN => Ckt432_M4_n17
    );
NAND2_X1_16: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => out370,
        A2 => in14,
        ZN => Ckt432_M4_n1
    );
NAND3_X1_17: ENTITY WORK.NAND3_X1
    PORT MAP (
        A1 => in17,
        A2 => Ckt432_M4_n3,
        A3 => Ckt432_M4_n4,
        ZN => Ckt432_I_7
    );
AOI22_X1_8: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => in11,
        A2 => out223,
        B1 => in21,
        B2 => out329,
        ZN => Ckt432_M4_n4
    );
NAND2_X1_17: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => in27,
        A2 => out370,
        ZN => Ckt432_M4_n3
    );
NAND3_X1_18: ENTITY WORK.NAND3_X1
    PORT MAP (
        A1 => in30,
        A2 => Ckt432_M4_n5,
        A3 => Ckt432_M4_n6,
        ZN => Ckt432_I_6
    );
AOI22_X1_9: ENTITY WORK.AOI22_X1
    PORT MAP (
        A1 => in24,
        A2 => out223,
        B1 => in34,
        B2 => out329,
        ZN => Ckt432_M4_n6
    );
NAND2_X1_18: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => in40,
        A2 => out370,
        ZN => Ckt432_M4_n5
    );
AND2_X1_1: ENTITY WORK.AND2_X1
    PORT MAP (
        A1 => Ckt432_I_8,
        A2 => Ckt432_M5_n1,
        ZN => out421
    );
AOI221_X1_1: ENTITY WORK.AOI221_X1
    PORT MAP (
        A => Ckt432_M5_n9,
        B1 => Ckt432_I_2,
        B2 => Ckt432_M5_n2,
        C1 => Ckt432_I_4,
        C2 => Ckt432_M5_n8,
        ZN => Ckt432_M5_n6
    );
INV_X1_30: ENTITY WORK.INV_X1
    PORT MAP (
        A => Ckt432_I_5,
        ZN => Ckt432_M5_n9
    );
INV_X1_31: ENTITY WORK.INV_X1
    PORT MAP (
        A => Ckt432_I_3,
        ZN => Ckt432_M5_n8
    );
INV_X1_32: ENTITY WORK.INV_X1
    PORT MAP (
        A => Ckt432_I_1,
        ZN => Ckt432_M5_n2
    );
OR4_X1_1: ENTITY WORK.OR4_X1
    PORT MAP (
        A1 => Ckt432_M5_n2,
        A2 => Ckt432_M5_n3,
        A3 => Ckt432_M5_n4,
        A4 => out430,
        ZN => Ckt432_M5_n1
    );
INV_X1_33: ENTITY WORK.INV_X1
    PORT MAP (
        A => Ckt432_I_0,
        ZN => Ckt432_M5_n3
    );
NAND4_X1_12: ENTITY WORK.NAND4_X1
    PORT MAP (
        A1 => Ckt432_I_7,
        A2 => Ckt432_I_6,
        A3 => Ckt432_I_5,
        A4 => Ckt432_I_4,
        ZN => out430
    );
NAND3_X1_19: ENTITY WORK.NAND3_X1
    PORT MAP (
        A1 => Ckt432_I_6,
        A2 => Ckt432_M5_n5,
        A3 => Ckt432_I_7,
        ZN => out431
    );
NAND3_X1_20: ENTITY WORK.NAND3_X1
    PORT MAP (
        A1 => Ckt432_I_4,
        A2 => Ckt432_M5_n4,
        A3 => Ckt432_I_5,
        ZN => Ckt432_M5_n5
    );
NAND2_X1_19: ENTITY WORK.NAND2_X1
    PORT MAP (
        A1 => Ckt432_I_3,
        A2 => Ckt432_I_2,
        ZN => Ckt432_M5_n4
    );
OAI21_X1_10: ENTITY WORK.OAI21_X1
    PORT MAP (
        A => Ckt432_I_7,
        B1 => Ckt432_M5_n6,
        B2 => Ckt432_M5_n7,
        ZN => out432
    );
INV_X1_34: ENTITY WORK.INV_X1
    PORT MAP (
        A => Ckt432_I_6,
        ZN => Ckt432_M5_n7
    );

END ARCHITECTURE arch;
