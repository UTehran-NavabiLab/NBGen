module counter_4bit(clk, rst, en, co, counter);

wire S0;
wire S1;
wire S2;
wire S3;
wire S4;
wire S5;
wire S6;
wire S7;
wire S8;
wire S9;
wire S10;
wire S11;
wire S12;
wire S13;
wire S14;
wire S15;
wire S16;
wire S17;
wire S18;
wire S19;
wire S20;
wire S21;
wire S22;
wire S23;
wire S24;
wire S25;
wire new_counter_reg_0;
wire new_counter_reg_1;
wire new_counter_reg_2;
wire new_counter_reg_3;
input clk;
input rst;
input en;
output co;
output [3:0] counter;
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_0_ (
  .A({ new_counter_reg_0 }),
  .Y({ S4 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1_ (
  .A({ new_counter_reg_3 }),
  .Y({ S5 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2_ (
  .A({ S20 }),
  .Y({ S6 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3_ (
  .A({ new_counter_reg_1, new_counter_reg_0 }),
  .Y({ S7 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4_ (
  .A({ new_counter_reg_2, new_counter_reg_3 }),
  .Y({ S8 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5_ (
  .A({ S8, S7 }),
  .Y({ S19 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6_ (
  .A({ S6, S4 }),
  .Y({ S9 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_7_ (
  .A({ S20, new_counter_reg_0 }),
  .Y({ S10 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_8_ (
  .A({ S10, S9 }),
  .Y({ S0 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_9_ (
  .A({ S7, S6 }),
  .Y({ S11 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_10_ (
  .A({ S9, new_counter_reg_1 }),
  .Y({ S12 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_11_ (
  .A({ S12, S11 }),
  .Y({ S1 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_12_ (
  .A({ S11, new_counter_reg_2 }),
  .Y({ S13 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_13_ (
  .A({ S13 }),
  .Y({ S14 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_14_ (
  .A({ S11, new_counter_reg_2 }),
  .Y({ S15 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_15_ (
  .A({ S15, S14 }),
  .Y({ S2 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_16_ (
  .A({ S14, new_counter_reg_3 }),
  .Y({ S16 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_17_ (
  .A({ S13, S5 }),
  .Y({ S17 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_18_ (
  .A({ S17, S16 }),
  .Y({ S3 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_19_ (
  .C({ S18 }),
  .CE({ 1'b1 }),
  .D({ S0 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_counter_reg_0 }),
  .R({ S21 }),
  .Si({ S22 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_20_ (
  .C({ S18 }),
  .CE({ 1'b1 }),
  .D({ S1 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_counter_reg_1 }),
  .R({ S21 }),
  .Si({ S23 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_21_ (
  .C({ S18 }),
  .CE({ 1'b1 }),
  .D({ S2 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_counter_reg_2 }),
  .R({ S21 }),
  .Si({ S24 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_22_ (
  .C({ S18 }),
  .CE({ 1'b1 }),
  .D({ S3 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_counter_reg_3 }),
  .R({ S21 }),
  .Si({ S25 }),
  .global_reset({ 1'b0 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_23_ (
  .I({ clk }),
  .O({ S18 })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_24_ (
  .I({ S19 }),
  .O({ co })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_25_ (
  .I({ new_counter_reg_0 }),
  .O({ counter[0] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_26_ (
  .I({ new_counter_reg_1 }),
  .O({ counter[1] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_27_ (
  .I({ new_counter_reg_2 }),
  .O({ counter[2] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_28_ (
  .I({ new_counter_reg_3 }),
  .O({ counter[3] })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_29_ (
  .I({ en }),
  .O({ S20 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_30_ (
  .I({ rst }),
  .O({ S21 })
);

endmodule