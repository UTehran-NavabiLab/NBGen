module counter(clk, rst, en, clkEn, count, co);

wire S0;
wire S1;
wire S2;
wire S3;
wire S4;
wire S5;
wire S6;
wire S7;
wire S8;
wire S9;
wire S10;
wire S11;
wire S12;
wire S13;
wire S14;
wire S15;
wire S16;
wire S17;
wire S18;
wire S19;
wire S20;
wire S21;
wire S22;
wire S23;
wire S24;
wire S25;
wire S26;
wire S27;
wire S28;
wire S29;
wire S30;
wire S31;
wire S32;
wire S33;
wire S34;
wire S35;
wire S36;
wire S37;
wire S38;
wire S39;
wire S40;
input clk;
input rst;
input en;
input clkEn;
output [3:0] count;output co;

notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_1_ (
  .in1({ S31 }),
  .out1({ S4 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_2_ (
  .in1({ S34 }),
  .out1({ S5 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_3_ (
  .in1({ S33 }),
  .out1({ S6 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_4_ (
  .in1({ S32 }),
  .out1({ S7 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_5_ (
  .in1({ S36 }),
  .out1({ S8 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1_ (
  .in1({ S34, S4 }),
  .out1({ S9 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_2_ (
  .in1({ S32, S6 }),
  .out1({ S10 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1_ (
  .in1({ S10, S9 }),
  .out1({ S30 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_3_ (
  .in1({ S35, S29 }),
  .out1({ S11 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_2_ (
  .in1({ S11, S4 }),
  .out1({ S12 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_6_ (
  .in1({ S12 }),
  .out1({ S13 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_4_ (
  .in1({ S11, S4 }),
  .out1({ S14 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_5_ (
  .in1({ S14, S8 }),
  .out1({ S15 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_3_ (
  .in1({ S15, S12 }),
  .out1({ S0 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_4_ (
  .in1({ S13, S7 }),
  .out1({ S16 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_6_ (
  .in1({ S12, S32 }),
  .out1({ S17 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_5_ (
  .in1({ S12, S32 }),
  .out1({ S18 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_6_ (
  .in1({ S18, S36 }),
  .out1({ S19 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_7_ (
  .in1({ S19, S17 }),
  .out1({ S20 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_7_ (
  .in1({ S20 }),
  .out1({ S1 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_8_ (
  .in1({ S16, S33 }),
  .out1({ S21 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_7_ (
  .in1({ S16, S33 }),
  .out1({ S22 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_8_ (
  .in1({ S22, S36 }),
  .out1({ S23 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_9_ (
  .in1({ S23, S21 }),
  .out1({ S24 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_8_ (
  .in1({ S24 }),
  .out1({ S2 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_9_ (
  .in1({ S21, S5 }),
  .out1({ S25 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_10_ (
  .in1({ S21, S5 }),
  .out1({ S26 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_11_ (
  .in1({ S26, S8 }),
  .out1({ S27 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_10_ (
  .in1({ S27, S25 }),
  .out1({ S3 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_1_ (
  .C({ S28 }),
  .CE({ 1'b1 }),
  .CLR({ 1'b0 }),
  .D({ S0 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ S31 }),
  .Si({ S37 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_2_ (
  .C({ S28 }),
  .CE({ 1'b1 }),
  .CLR({ 1'b0 }),
  .D({ S1 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ S32 }),
  .Si({ S38 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_3_ (
  .C({ S28 }),
  .CE({ 1'b1 }),
  .CLR({ 1'b0 }),
  .D({ S2 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ S33 }),
  .Si({ S39 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_4_ (
  .C({ S28 }),
  .CE({ 1'b1 }),
  .CLR({ 1'b0 }),
  .D({ S3 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ S34 }),
  .Si({ S40 }),
  .global_reset({ 1'b0 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_1_ (
  .in1({ clk }),
  .out1({ S28 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_2_ (
  .in1({ clkEn }),
  .out1({ S29 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_3_ (
  .in1({ S30 }),
  .out1({ co })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_4_ (
  .in1({ S31 }),
  .out1({ count[0] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_5_ (
  .in1({ S32 }),
  .out1({ count[1] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_6_ (
  .in1({ S33 }),
  .out1({ count[2] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_7_ (
  .in1({ S34 }),
  .out1({ count[3] })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_8_ (
  .in1({ en }),
  .out1({ S35 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_9_ (
  .in1({ rst }),
  .out1({ S36 })
);

endmodule