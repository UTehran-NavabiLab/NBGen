LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

ENTITY SAYAC_TOP IS
    PORT (
        clk : IN STD_LOGIC;
        rst : IN STD_LOGIC;
        readyMEM : IN STD_LOGIC;
        dataBusIn : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
        readMEM : OUT STD_LOGIC;
        writeMEM : OUT STD_LOGIC;
        readIO : OUT STD_LOGIC;
        writeIO : OUT STD_LOGIC;
        dataBusOut : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
        addrBus : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
        readInst : OUT STD_LOGIC;
        PCout : OUT STD_LOGIC_VECTOR (15 DOWNTO 0));
END ENTITY SAYAC_TOP;

ARCHITECTURE arch OF SAYAC_TOP IS
    SIGNAL S0 : STD_LOGIC;
    SIGNAL S1 : STD_LOGIC;
    SIGNAL S2 : STD_LOGIC;
    SIGNAL S3 : STD_LOGIC;
    SIGNAL S4 : STD_LOGIC;
    SIGNAL S5 : STD_LOGIC;
    SIGNAL S6 : STD_LOGIC;
    SIGNAL S7 : STD_LOGIC;
    SIGNAL S8 : STD_LOGIC;
    SIGNAL S9 : STD_LOGIC;
    SIGNAL S10 : STD_LOGIC;
    SIGNAL S11 : STD_LOGIC;
    SIGNAL S12 : STD_LOGIC;
    SIGNAL S13 : STD_LOGIC;
    SIGNAL S14 : STD_LOGIC;
    SIGNAL S15 : STD_LOGIC;
    SIGNAL S16 : STD_LOGIC;
    SIGNAL S17 : STD_LOGIC;
    SIGNAL S18 : STD_LOGIC;
    SIGNAL S19 : STD_LOGIC;
    SIGNAL S20 : STD_LOGIC;
    SIGNAL S21 : STD_LOGIC;
    SIGNAL S22 : STD_LOGIC;
    SIGNAL S23 : STD_LOGIC;
    SIGNAL S24 : STD_LOGIC;
    SIGNAL S25 : STD_LOGIC;
    SIGNAL S26 : STD_LOGIC;
    SIGNAL S27 : STD_LOGIC;
    SIGNAL S28 : STD_LOGIC;
    SIGNAL S29 : STD_LOGIC;
    SIGNAL S30 : STD_LOGIC;
    SIGNAL S31 : STD_LOGIC;
    SIGNAL S32 : STD_LOGIC;
    SIGNAL S33 : STD_LOGIC;
    SIGNAL S34 : STD_LOGIC;
    SIGNAL S35 : STD_LOGIC;
    SIGNAL S36 : STD_LOGIC;
    SIGNAL S37 : STD_LOGIC;
    SIGNAL S38 : STD_LOGIC;
    SIGNAL S39 : STD_LOGIC;
    SIGNAL S40 : STD_LOGIC;
    SIGNAL S41 : STD_LOGIC;
    SIGNAL S42 : STD_LOGIC;
    SIGNAL S43 : STD_LOGIC;
    SIGNAL S44 : STD_LOGIC;
    SIGNAL S45 : STD_LOGIC;
    SIGNAL S46 : STD_LOGIC;
    SIGNAL S47 : STD_LOGIC;
    SIGNAL S48 : STD_LOGIC;
    SIGNAL S49 : STD_LOGIC;
    SIGNAL S50 : STD_LOGIC;
    SIGNAL S51 : STD_LOGIC;
    SIGNAL S52 : STD_LOGIC;
    SIGNAL S53 : STD_LOGIC;
    SIGNAL S54 : STD_LOGIC;
    SIGNAL S55 : STD_LOGIC;
    SIGNAL S56 : STD_LOGIC;
    SIGNAL S57 : STD_LOGIC;
    SIGNAL S58 : STD_LOGIC;
    SIGNAL S59 : STD_LOGIC;
    SIGNAL S60 : STD_LOGIC;
    SIGNAL S61 : STD_LOGIC;
    SIGNAL S62 : STD_LOGIC;
    SIGNAL S63 : STD_LOGIC;
    SIGNAL S64 : STD_LOGIC;
    SIGNAL S65 : STD_LOGIC;
    SIGNAL S66 : STD_LOGIC;
    SIGNAL S67 : STD_LOGIC;
    SIGNAL S68 : STD_LOGIC;
    SIGNAL S69 : STD_LOGIC;
    SIGNAL S70 : STD_LOGIC;
    SIGNAL S71 : STD_LOGIC;
    SIGNAL S72 : STD_LOGIC;
    SIGNAL S73 : STD_LOGIC;
    SIGNAL S74 : STD_LOGIC;
    SIGNAL S75 : STD_LOGIC;
    SIGNAL S76 : STD_LOGIC;
    SIGNAL S77 : STD_LOGIC;
    SIGNAL S78 : STD_LOGIC;
    SIGNAL S79 : STD_LOGIC;
    SIGNAL S80 : STD_LOGIC;
    SIGNAL S81 : STD_LOGIC;
    SIGNAL S82 : STD_LOGIC;
    SIGNAL S83 : STD_LOGIC;
    SIGNAL S84 : STD_LOGIC;
    SIGNAL S85 : STD_LOGIC;
    SIGNAL S86 : STD_LOGIC;
    SIGNAL S87 : STD_LOGIC;
    SIGNAL S88 : STD_LOGIC;
    SIGNAL S89 : STD_LOGIC;
    SIGNAL S90 : STD_LOGIC;
    SIGNAL S91 : STD_LOGIC;
    SIGNAL S92 : STD_LOGIC;
    SIGNAL S93 : STD_LOGIC;
    SIGNAL S94 : STD_LOGIC;
    SIGNAL S95 : STD_LOGIC;
    SIGNAL S96 : STD_LOGIC;
    SIGNAL S97 : STD_LOGIC;
    SIGNAL S98 : STD_LOGIC;
    SIGNAL S99 : STD_LOGIC;
    SIGNAL S100 : STD_LOGIC;
    SIGNAL S101 : STD_LOGIC;
    SIGNAL S102 : STD_LOGIC;
    SIGNAL S103 : STD_LOGIC;
    SIGNAL S104 : STD_LOGIC;
    SIGNAL S105 : STD_LOGIC;
    SIGNAL S106 : STD_LOGIC;
    SIGNAL S107 : STD_LOGIC;
    SIGNAL S108 : STD_LOGIC;
    SIGNAL S109 : STD_LOGIC;
    SIGNAL S110 : STD_LOGIC;
    SIGNAL S111 : STD_LOGIC;
    SIGNAL S112 : STD_LOGIC;
    SIGNAL S113 : STD_LOGIC;
    SIGNAL S114 : STD_LOGIC;
    SIGNAL S115 : STD_LOGIC;
    SIGNAL S116 : STD_LOGIC;
    SIGNAL S117 : STD_LOGIC;
    SIGNAL S118 : STD_LOGIC;
    SIGNAL S119 : STD_LOGIC;
    SIGNAL S120 : STD_LOGIC;
    SIGNAL S121 : STD_LOGIC;
    SIGNAL S122 : STD_LOGIC;
    SIGNAL S123 : STD_LOGIC;
    SIGNAL S124 : STD_LOGIC;
    SIGNAL S125 : STD_LOGIC;
    SIGNAL S126 : STD_LOGIC;
    SIGNAL S127 : STD_LOGIC;
    SIGNAL S128 : STD_LOGIC;
    SIGNAL S129 : STD_LOGIC;
    SIGNAL S130 : STD_LOGIC;
    SIGNAL S131 : STD_LOGIC;
    SIGNAL S132 : STD_LOGIC;
    SIGNAL S133 : STD_LOGIC;
    SIGNAL S134 : STD_LOGIC;
    SIGNAL S135 : STD_LOGIC;
    SIGNAL S136 : STD_LOGIC;
    SIGNAL S137 : STD_LOGIC;
    SIGNAL S138 : STD_LOGIC;
    SIGNAL S139 : STD_LOGIC;
    SIGNAL S140 : STD_LOGIC;
    SIGNAL S141 : STD_LOGIC;
    SIGNAL S142 : STD_LOGIC;
    SIGNAL S143 : STD_LOGIC;
    SIGNAL S144 : STD_LOGIC;
    SIGNAL S145 : STD_LOGIC;
    SIGNAL S146 : STD_LOGIC;
    SIGNAL S147 : STD_LOGIC;
    SIGNAL S148 : STD_LOGIC;
    SIGNAL S149 : STD_LOGIC;
    SIGNAL S150 : STD_LOGIC;
    SIGNAL S151 : STD_LOGIC;
    SIGNAL S152 : STD_LOGIC;
    SIGNAL S153 : STD_LOGIC;
    SIGNAL S154 : STD_LOGIC;
    SIGNAL S155 : STD_LOGIC;
    SIGNAL S156 : STD_LOGIC;
    SIGNAL S157 : STD_LOGIC;
    SIGNAL S158 : STD_LOGIC;
    SIGNAL S159 : STD_LOGIC;
    SIGNAL S160 : STD_LOGIC;
    SIGNAL S161 : STD_LOGIC;
    SIGNAL S162 : STD_LOGIC;
    SIGNAL S163 : STD_LOGIC;
    SIGNAL S164 : STD_LOGIC;
    SIGNAL S165 : STD_LOGIC;
    SIGNAL S166 : STD_LOGIC;
    SIGNAL S167 : STD_LOGIC;
    SIGNAL S168 : STD_LOGIC;
    SIGNAL S169 : STD_LOGIC;
    SIGNAL S170 : STD_LOGIC;
    SIGNAL S171 : STD_LOGIC;
    SIGNAL S172 : STD_LOGIC;
    SIGNAL S173 : STD_LOGIC;
    SIGNAL S174 : STD_LOGIC;
    SIGNAL S175 : STD_LOGIC;
    SIGNAL S176 : STD_LOGIC;
    SIGNAL S177 : STD_LOGIC;
    SIGNAL S178 : STD_LOGIC;
    SIGNAL S179 : STD_LOGIC;
    SIGNAL S180 : STD_LOGIC;
    SIGNAL S181 : STD_LOGIC;
    SIGNAL S182 : STD_LOGIC;
    SIGNAL S183 : STD_LOGIC;
    SIGNAL S184 : STD_LOGIC;
    SIGNAL S185 : STD_LOGIC;
    SIGNAL S186 : STD_LOGIC;
    SIGNAL S187 : STD_LOGIC;
    SIGNAL S188 : STD_LOGIC;
    SIGNAL S189 : STD_LOGIC;
    SIGNAL S190 : STD_LOGIC;
    SIGNAL S191 : STD_LOGIC;
    SIGNAL S192 : STD_LOGIC;
    SIGNAL S193 : STD_LOGIC;
    SIGNAL S194 : STD_LOGIC;
    SIGNAL S195 : STD_LOGIC;
    SIGNAL S196 : STD_LOGIC;
    SIGNAL S197 : STD_LOGIC;
    SIGNAL S198 : STD_LOGIC;
    SIGNAL S199 : STD_LOGIC;
    SIGNAL S200 : STD_LOGIC;
    SIGNAL S201 : STD_LOGIC;
    SIGNAL S202 : STD_LOGIC;
    SIGNAL S203 : STD_LOGIC;
    SIGNAL S204 : STD_LOGIC;
    SIGNAL S205 : STD_LOGIC;
    SIGNAL S206 : STD_LOGIC;
    SIGNAL S207 : STD_LOGIC;
    SIGNAL S208 : STD_LOGIC;
    SIGNAL S209 : STD_LOGIC;
    SIGNAL S210 : STD_LOGIC;
    SIGNAL S211 : STD_LOGIC;
    SIGNAL S212 : STD_LOGIC;
    SIGNAL S213 : STD_LOGIC;
    SIGNAL S214 : STD_LOGIC;
    SIGNAL S215 : STD_LOGIC;
    SIGNAL S216 : STD_LOGIC;
    SIGNAL S217 : STD_LOGIC;
    SIGNAL S218 : STD_LOGIC;
    SIGNAL S219 : STD_LOGIC;
    SIGNAL S220 : STD_LOGIC;
    SIGNAL S221 : STD_LOGIC;
    SIGNAL S222 : STD_LOGIC;
    SIGNAL S223 : STD_LOGIC;
    SIGNAL S224 : STD_LOGIC;
    SIGNAL S225 : STD_LOGIC;
    SIGNAL S226 : STD_LOGIC;
    SIGNAL S227 : STD_LOGIC;
    SIGNAL S228 : STD_LOGIC;
    SIGNAL S229 : STD_LOGIC;
    SIGNAL S230 : STD_LOGIC;
    SIGNAL S231 : STD_LOGIC;
    SIGNAL S232 : STD_LOGIC;
    SIGNAL S233 : STD_LOGIC;
    SIGNAL S234 : STD_LOGIC;
    SIGNAL S235 : STD_LOGIC;
    SIGNAL S236 : STD_LOGIC;
    SIGNAL S237 : STD_LOGIC;
    SIGNAL S238 : STD_LOGIC;
    SIGNAL S239 : STD_LOGIC;
    SIGNAL S240 : STD_LOGIC;
    SIGNAL S241 : STD_LOGIC;
    SIGNAL S242 : STD_LOGIC;
    SIGNAL S243 : STD_LOGIC;
    SIGNAL S244 : STD_LOGIC;
    SIGNAL S245 : STD_LOGIC;
    SIGNAL S246 : STD_LOGIC;
    SIGNAL S247 : STD_LOGIC;
    SIGNAL S248 : STD_LOGIC;
    SIGNAL S249 : STD_LOGIC;
    SIGNAL S250 : STD_LOGIC;
    SIGNAL S251 : STD_LOGIC;
    SIGNAL S252 : STD_LOGIC;
    SIGNAL S253 : STD_LOGIC;
    SIGNAL S254 : STD_LOGIC;
    SIGNAL S255 : STD_LOGIC;
    SIGNAL S256 : STD_LOGIC;
    SIGNAL S257 : STD_LOGIC;
    SIGNAL S258 : STD_LOGIC;
    SIGNAL S259 : STD_LOGIC;
    SIGNAL S260 : STD_LOGIC;
    SIGNAL S261 : STD_LOGIC;
    SIGNAL S262 : STD_LOGIC;
    SIGNAL S263 : STD_LOGIC;
    SIGNAL S264 : STD_LOGIC;
    SIGNAL S265 : STD_LOGIC;
    SIGNAL S266 : STD_LOGIC;
    SIGNAL S267 : STD_LOGIC;
    SIGNAL S268 : STD_LOGIC;
    SIGNAL S269 : STD_LOGIC;
    SIGNAL S270 : STD_LOGIC;
    SIGNAL S271 : STD_LOGIC;
    SIGNAL S272 : STD_LOGIC;
    SIGNAL S273 : STD_LOGIC;
    SIGNAL S274 : STD_LOGIC;
    SIGNAL S275 : STD_LOGIC;
    SIGNAL S276 : STD_LOGIC;
    SIGNAL S277 : STD_LOGIC;
    SIGNAL S278 : STD_LOGIC;
    SIGNAL S279 : STD_LOGIC;
    SIGNAL S280 : STD_LOGIC;
    SIGNAL S281 : STD_LOGIC;
    SIGNAL S282 : STD_LOGIC;
    SIGNAL S283 : STD_LOGIC;
    SIGNAL S284 : STD_LOGIC;
    SIGNAL S285 : STD_LOGIC;
    SIGNAL S286 : STD_LOGIC;
    SIGNAL S287 : STD_LOGIC;
    SIGNAL S288 : STD_LOGIC;
    SIGNAL S289 : STD_LOGIC;
    SIGNAL S290 : STD_LOGIC;
    SIGNAL S291 : STD_LOGIC;
    SIGNAL S292 : STD_LOGIC;
    SIGNAL S293 : STD_LOGIC;
    SIGNAL S294 : STD_LOGIC;
    SIGNAL S295 : STD_LOGIC;
    SIGNAL S296 : STD_LOGIC;
    SIGNAL S297 : STD_LOGIC;
    SIGNAL S298 : STD_LOGIC;
    SIGNAL S299 : STD_LOGIC;
    SIGNAL S300 : STD_LOGIC;
    SIGNAL S301 : STD_LOGIC;
    SIGNAL S302 : STD_LOGIC;
    SIGNAL S303 : STD_LOGIC;
    SIGNAL S304 : STD_LOGIC;
    SIGNAL S305 : STD_LOGIC;
    SIGNAL S306 : STD_LOGIC;
    SIGNAL S307 : STD_LOGIC;
    SIGNAL S308 : STD_LOGIC;
    SIGNAL S309 : STD_LOGIC;
    SIGNAL S310 : STD_LOGIC;
    SIGNAL S311 : STD_LOGIC;
    SIGNAL S312 : STD_LOGIC;
    SIGNAL S313 : STD_LOGIC;
    SIGNAL S314 : STD_LOGIC;
    SIGNAL S315 : STD_LOGIC;
    SIGNAL S316 : STD_LOGIC;
    SIGNAL S317 : STD_LOGIC;
    SIGNAL S318 : STD_LOGIC;
    SIGNAL S319 : STD_LOGIC;
    SIGNAL S320 : STD_LOGIC;
    SIGNAL S321 : STD_LOGIC;
    SIGNAL S322 : STD_LOGIC;
    SIGNAL S323 : STD_LOGIC;
    SIGNAL S324 : STD_LOGIC;
    SIGNAL S325 : STD_LOGIC;
    SIGNAL S326 : STD_LOGIC;
    SIGNAL S327 : STD_LOGIC;
    SIGNAL S328 : STD_LOGIC;
    SIGNAL S329 : STD_LOGIC;
    SIGNAL S330 : STD_LOGIC;
    SIGNAL S331 : STD_LOGIC;
    SIGNAL S332 : STD_LOGIC;
    SIGNAL S333 : STD_LOGIC;
    SIGNAL S334 : STD_LOGIC;
    SIGNAL S335 : STD_LOGIC;
    SIGNAL S336 : STD_LOGIC;
    SIGNAL S337 : STD_LOGIC;
    SIGNAL S338 : STD_LOGIC;
    SIGNAL S339 : STD_LOGIC;
    SIGNAL S340 : STD_LOGIC;
    SIGNAL S341 : STD_LOGIC;
    SIGNAL S342 : STD_LOGIC;
    SIGNAL S343 : STD_LOGIC;
    SIGNAL S344 : STD_LOGIC;
    SIGNAL S345 : STD_LOGIC;
    SIGNAL S346 : STD_LOGIC;
    SIGNAL S347 : STD_LOGIC;
    SIGNAL S348 : STD_LOGIC;
    SIGNAL S349 : STD_LOGIC;
    SIGNAL S350 : STD_LOGIC;
    SIGNAL S351 : STD_LOGIC;
    SIGNAL S352 : STD_LOGIC;
    SIGNAL S353 : STD_LOGIC;
    SIGNAL S354 : STD_LOGIC;
    SIGNAL S355 : STD_LOGIC;
    SIGNAL S356 : STD_LOGIC;
    SIGNAL S357 : STD_LOGIC;
    SIGNAL S358 : STD_LOGIC;
    SIGNAL S359 : STD_LOGIC;
    SIGNAL S360 : STD_LOGIC;
    SIGNAL S361 : STD_LOGIC;
    SIGNAL S362 : STD_LOGIC;
    SIGNAL S363 : STD_LOGIC;
    SIGNAL S364 : STD_LOGIC;
    SIGNAL S365 : STD_LOGIC;
    SIGNAL S366 : STD_LOGIC;
    SIGNAL S367 : STD_LOGIC;
    SIGNAL S368 : STD_LOGIC;
    SIGNAL S369 : STD_LOGIC;
    SIGNAL S370 : STD_LOGIC;
    SIGNAL S371 : STD_LOGIC;
    SIGNAL S372 : STD_LOGIC;
    SIGNAL S373 : STD_LOGIC;
    SIGNAL S374 : STD_LOGIC;
    SIGNAL S375 : STD_LOGIC;
    SIGNAL S376 : STD_LOGIC;
    SIGNAL S377 : STD_LOGIC;
    SIGNAL S378 : STD_LOGIC;
    SIGNAL S379 : STD_LOGIC;
    SIGNAL S380 : STD_LOGIC;
    SIGNAL S381 : STD_LOGIC;
    SIGNAL S382 : STD_LOGIC;
    SIGNAL S383 : STD_LOGIC;
    SIGNAL S384 : STD_LOGIC;
    SIGNAL S385 : STD_LOGIC;
    SIGNAL S386 : STD_LOGIC;
    SIGNAL S387 : STD_LOGIC;
    SIGNAL S388 : STD_LOGIC;
    SIGNAL S389 : STD_LOGIC;
    SIGNAL S390 : STD_LOGIC;
    SIGNAL S391 : STD_LOGIC;
    SIGNAL S392 : STD_LOGIC;
    SIGNAL S393 : STD_LOGIC;
    SIGNAL S394 : STD_LOGIC;
    SIGNAL S395 : STD_LOGIC;
    SIGNAL S396 : STD_LOGIC;
    SIGNAL S397 : STD_LOGIC;
    SIGNAL S398 : STD_LOGIC;
    SIGNAL S399 : STD_LOGIC;
    SIGNAL S400 : STD_LOGIC;
    SIGNAL S401 : STD_LOGIC;
    SIGNAL S402 : STD_LOGIC;
    SIGNAL S403 : STD_LOGIC;
    SIGNAL S404 : STD_LOGIC;
    SIGNAL S405 : STD_LOGIC;
    SIGNAL S406 : STD_LOGIC;
    SIGNAL S407 : STD_LOGIC;
    SIGNAL S408 : STD_LOGIC;
    SIGNAL S409 : STD_LOGIC;
    SIGNAL S410 : STD_LOGIC;
    SIGNAL S411 : STD_LOGIC;
    SIGNAL S412 : STD_LOGIC;
    SIGNAL S413 : STD_LOGIC;
    SIGNAL S414 : STD_LOGIC;
    SIGNAL S415 : STD_LOGIC;
    SIGNAL S416 : STD_LOGIC;
    SIGNAL S417 : STD_LOGIC;
    SIGNAL S418 : STD_LOGIC;
    SIGNAL S419 : STD_LOGIC;
    SIGNAL S420 : STD_LOGIC;
    SIGNAL S421 : STD_LOGIC;
    SIGNAL S422 : STD_LOGIC;
    SIGNAL S423 : STD_LOGIC;
    SIGNAL S424 : STD_LOGIC;
    SIGNAL S425 : STD_LOGIC;
    SIGNAL S426 : STD_LOGIC;
    SIGNAL S427 : STD_LOGIC;
    SIGNAL S428 : STD_LOGIC;
    SIGNAL S429 : STD_LOGIC;
    SIGNAL S430 : STD_LOGIC;
    SIGNAL S431 : STD_LOGIC;
    SIGNAL S432 : STD_LOGIC;
    SIGNAL S433 : STD_LOGIC;
    SIGNAL S434 : STD_LOGIC;
    SIGNAL S435 : STD_LOGIC;
    SIGNAL S436 : STD_LOGIC;
    SIGNAL S437 : STD_LOGIC;
    SIGNAL S438 : STD_LOGIC;
    SIGNAL S439 : STD_LOGIC;
    SIGNAL S440 : STD_LOGIC;
    SIGNAL S441 : STD_LOGIC;
    SIGNAL S442 : STD_LOGIC;
    SIGNAL S443 : STD_LOGIC;
    SIGNAL S444 : STD_LOGIC;
    SIGNAL S445 : STD_LOGIC;
    SIGNAL S446 : STD_LOGIC;
    SIGNAL S447 : STD_LOGIC;
    SIGNAL S448 : STD_LOGIC;
    SIGNAL S449 : STD_LOGIC;
    SIGNAL S450 : STD_LOGIC;
    SIGNAL S451 : STD_LOGIC;
    SIGNAL S452 : STD_LOGIC;
    SIGNAL S453 : STD_LOGIC;
    SIGNAL S454 : STD_LOGIC;
    SIGNAL S455 : STD_LOGIC;
    SIGNAL S456 : STD_LOGIC;
    SIGNAL S457 : STD_LOGIC;
    SIGNAL S458 : STD_LOGIC;
    SIGNAL S459 : STD_LOGIC;
    SIGNAL S460 : STD_LOGIC;
    SIGNAL S461 : STD_LOGIC;
    SIGNAL S462 : STD_LOGIC;
    SIGNAL S463 : STD_LOGIC;
    SIGNAL S464 : STD_LOGIC;
    SIGNAL S465 : STD_LOGIC;
    SIGNAL S466 : STD_LOGIC;
    SIGNAL S467 : STD_LOGIC;
    SIGNAL S468 : STD_LOGIC;
    SIGNAL S469 : STD_LOGIC;
    SIGNAL S470 : STD_LOGIC;
    SIGNAL S471 : STD_LOGIC;
    SIGNAL S472 : STD_LOGIC;
    SIGNAL S473 : STD_LOGIC;
    SIGNAL S474 : STD_LOGIC;
    SIGNAL S475 : STD_LOGIC;
    SIGNAL S476 : STD_LOGIC;
    SIGNAL S477 : STD_LOGIC;
    SIGNAL S478 : STD_LOGIC;
    SIGNAL S479 : STD_LOGIC;
    SIGNAL S480 : STD_LOGIC;
    SIGNAL S481 : STD_LOGIC;
    SIGNAL S482 : STD_LOGIC;
    SIGNAL S483 : STD_LOGIC;
    SIGNAL S484 : STD_LOGIC;
    SIGNAL S485 : STD_LOGIC;
    SIGNAL S486 : STD_LOGIC;
    SIGNAL S487 : STD_LOGIC;
    SIGNAL S488 : STD_LOGIC;
    SIGNAL S489 : STD_LOGIC;
    SIGNAL S490 : STD_LOGIC;
    SIGNAL S491 : STD_LOGIC;
    SIGNAL S492 : STD_LOGIC;
    SIGNAL S493 : STD_LOGIC;
    SIGNAL S494 : STD_LOGIC;
    SIGNAL S495 : STD_LOGIC;
    SIGNAL S496 : STD_LOGIC;
    SIGNAL S497 : STD_LOGIC;
    SIGNAL S498 : STD_LOGIC;
    SIGNAL S499 : STD_LOGIC;
    SIGNAL S500 : STD_LOGIC;
    SIGNAL S501 : STD_LOGIC;
    SIGNAL S502 : STD_LOGIC;
    SIGNAL S503 : STD_LOGIC;
    SIGNAL S504 : STD_LOGIC;
    SIGNAL S505 : STD_LOGIC;
    SIGNAL S506 : STD_LOGIC;
    SIGNAL S507 : STD_LOGIC;
    SIGNAL S508 : STD_LOGIC;
    SIGNAL S509 : STD_LOGIC;
    SIGNAL S510 : STD_LOGIC;
    SIGNAL S511 : STD_LOGIC;
    SIGNAL S512 : STD_LOGIC;
    SIGNAL S513 : STD_LOGIC;
    SIGNAL S514 : STD_LOGIC;
    SIGNAL S515 : STD_LOGIC;
    SIGNAL S516 : STD_LOGIC;
    SIGNAL S517 : STD_LOGIC;
    SIGNAL S518 : STD_LOGIC;
    SIGNAL S519 : STD_LOGIC;
    SIGNAL S520 : STD_LOGIC;
    SIGNAL S521 : STD_LOGIC;
    SIGNAL S522 : STD_LOGIC;
    SIGNAL S523 : STD_LOGIC;
    SIGNAL S524 : STD_LOGIC;
    SIGNAL S525 : STD_LOGIC;
    SIGNAL S526 : STD_LOGIC;
    SIGNAL S527 : STD_LOGIC;
    SIGNAL S528 : STD_LOGIC;
    SIGNAL S529 : STD_LOGIC;
    SIGNAL S530 : STD_LOGIC;
    SIGNAL S531 : STD_LOGIC;
    SIGNAL S532 : STD_LOGIC;
    SIGNAL S533 : STD_LOGIC;
    SIGNAL S534 : STD_LOGIC;
    SIGNAL S535 : STD_LOGIC;
    SIGNAL S536 : STD_LOGIC;
    SIGNAL S537 : STD_LOGIC;
    SIGNAL S538 : STD_LOGIC;
    SIGNAL S539 : STD_LOGIC;
    SIGNAL S540 : STD_LOGIC;
    SIGNAL S541 : STD_LOGIC;
    SIGNAL S542 : STD_LOGIC;
    SIGNAL S543 : STD_LOGIC;
    SIGNAL S544 : STD_LOGIC;
    SIGNAL S545 : STD_LOGIC;
    SIGNAL S546 : STD_LOGIC;
    SIGNAL S547 : STD_LOGIC;
    SIGNAL S548 : STD_LOGIC;
    SIGNAL S549 : STD_LOGIC;
    SIGNAL S550 : STD_LOGIC;
    SIGNAL S551 : STD_LOGIC;
    SIGNAL S552 : STD_LOGIC;
    SIGNAL S553 : STD_LOGIC;
    SIGNAL S554 : STD_LOGIC;
    SIGNAL S555 : STD_LOGIC;
    SIGNAL S556 : STD_LOGIC;
    SIGNAL S557 : STD_LOGIC;
    SIGNAL S558 : STD_LOGIC;
    SIGNAL S559 : STD_LOGIC;
    SIGNAL S560 : STD_LOGIC;
    SIGNAL S561 : STD_LOGIC;
    SIGNAL S562 : STD_LOGIC;
    SIGNAL S563 : STD_LOGIC;
    SIGNAL S564 : STD_LOGIC;
    SIGNAL S565 : STD_LOGIC;
    SIGNAL S566 : STD_LOGIC;
    SIGNAL S567 : STD_LOGIC;
    SIGNAL S568 : STD_LOGIC;
    SIGNAL S569 : STD_LOGIC;
    SIGNAL S570 : STD_LOGIC;
    SIGNAL S571 : STD_LOGIC;
    SIGNAL S572 : STD_LOGIC;
    SIGNAL S573 : STD_LOGIC;
    SIGNAL S574 : STD_LOGIC;
    SIGNAL S575 : STD_LOGIC;
    SIGNAL S576 : STD_LOGIC;
    SIGNAL S577 : STD_LOGIC;
    SIGNAL S578 : STD_LOGIC;
    SIGNAL S579 : STD_LOGIC;
    SIGNAL S580 : STD_LOGIC;
    SIGNAL S581 : STD_LOGIC;
    SIGNAL S582 : STD_LOGIC;
    SIGNAL S583 : STD_LOGIC;
    SIGNAL S584 : STD_LOGIC;
    SIGNAL S585 : STD_LOGIC;
    SIGNAL S586 : STD_LOGIC;
    SIGNAL S587 : STD_LOGIC;
    SIGNAL S588 : STD_LOGIC;
    SIGNAL S589 : STD_LOGIC;
    SIGNAL S590 : STD_LOGIC;
    SIGNAL S591 : STD_LOGIC;
    SIGNAL S592 : STD_LOGIC;
    SIGNAL S593 : STD_LOGIC;
    SIGNAL S594 : STD_LOGIC;
    SIGNAL S595 : STD_LOGIC;
    SIGNAL S596 : STD_LOGIC;
    SIGNAL S597 : STD_LOGIC;
    SIGNAL S598 : STD_LOGIC;
    SIGNAL S599 : STD_LOGIC;
    SIGNAL S600 : STD_LOGIC;
    SIGNAL S601 : STD_LOGIC;
    SIGNAL S602 : STD_LOGIC;
    SIGNAL S603 : STD_LOGIC;
    SIGNAL S604 : STD_LOGIC;
    SIGNAL S605 : STD_LOGIC;
    SIGNAL S606 : STD_LOGIC;
    SIGNAL S607 : STD_LOGIC;
    SIGNAL S608 : STD_LOGIC;
    SIGNAL S609 : STD_LOGIC;
    SIGNAL S610 : STD_LOGIC;
    SIGNAL S611 : STD_LOGIC;
    SIGNAL S612 : STD_LOGIC;
    SIGNAL S613 : STD_LOGIC;
    SIGNAL S614 : STD_LOGIC;
    SIGNAL S615 : STD_LOGIC;
    SIGNAL S616 : STD_LOGIC;
    SIGNAL S617 : STD_LOGIC;
    SIGNAL S618 : STD_LOGIC;
    SIGNAL S619 : STD_LOGIC;
    SIGNAL S620 : STD_LOGIC;
    SIGNAL S621 : STD_LOGIC;
    SIGNAL S622 : STD_LOGIC;
    SIGNAL S623 : STD_LOGIC;
    SIGNAL S624 : STD_LOGIC;
    SIGNAL S625 : STD_LOGIC;
    SIGNAL S626 : STD_LOGIC;
    SIGNAL S627 : STD_LOGIC;
    SIGNAL S628 : STD_LOGIC;
    SIGNAL S629 : STD_LOGIC;
    SIGNAL S630 : STD_LOGIC;
    SIGNAL S631 : STD_LOGIC;
    SIGNAL S632 : STD_LOGIC;
    SIGNAL S633 : STD_LOGIC;
    SIGNAL S634 : STD_LOGIC;
    SIGNAL S635 : STD_LOGIC;
    SIGNAL S636 : STD_LOGIC;
    SIGNAL S637 : STD_LOGIC;
    SIGNAL S638 : STD_LOGIC;
    SIGNAL S639 : STD_LOGIC;
    SIGNAL S640 : STD_LOGIC;
    SIGNAL S641 : STD_LOGIC;
    SIGNAL S642 : STD_LOGIC;
    SIGNAL S643 : STD_LOGIC;
    SIGNAL S644 : STD_LOGIC;
    SIGNAL S645 : STD_LOGIC;
    SIGNAL S646 : STD_LOGIC;
    SIGNAL S647 : STD_LOGIC;
    SIGNAL S648 : STD_LOGIC;
    SIGNAL S649 : STD_LOGIC;
    SIGNAL S650 : STD_LOGIC;
    SIGNAL S651 : STD_LOGIC;
    SIGNAL S652 : STD_LOGIC;
    SIGNAL S653 : STD_LOGIC;
    SIGNAL S654 : STD_LOGIC;
    SIGNAL S655 : STD_LOGIC;
    SIGNAL S656 : STD_LOGIC;
    SIGNAL S657 : STD_LOGIC;
    SIGNAL S658 : STD_LOGIC;
    SIGNAL S659 : STD_LOGIC;
    SIGNAL S660 : STD_LOGIC;
    SIGNAL S661 : STD_LOGIC;
    SIGNAL S662 : STD_LOGIC;
    SIGNAL S663 : STD_LOGIC;
    SIGNAL S664 : STD_LOGIC;
    SIGNAL S665 : STD_LOGIC;
    SIGNAL S666 : STD_LOGIC;
    SIGNAL S667 : STD_LOGIC;
    SIGNAL S668 : STD_LOGIC;
    SIGNAL S669 : STD_LOGIC;
    SIGNAL S670 : STD_LOGIC;
    SIGNAL S671 : STD_LOGIC;
    SIGNAL S672 : STD_LOGIC;
    SIGNAL S673 : STD_LOGIC;
    SIGNAL S674 : STD_LOGIC;
    SIGNAL S675 : STD_LOGIC;
    SIGNAL S676 : STD_LOGIC;
    SIGNAL S677 : STD_LOGIC;
    SIGNAL S678 : STD_LOGIC;
    SIGNAL S679 : STD_LOGIC;
    SIGNAL S680 : STD_LOGIC;
    SIGNAL S681 : STD_LOGIC;
    SIGNAL S682 : STD_LOGIC;
    SIGNAL S683 : STD_LOGIC;
    SIGNAL S684 : STD_LOGIC;
    SIGNAL S685 : STD_LOGIC;
    SIGNAL S686 : STD_LOGIC;
    SIGNAL S687 : STD_LOGIC;
    SIGNAL S688 : STD_LOGIC;
    SIGNAL S689 : STD_LOGIC;
    SIGNAL S690 : STD_LOGIC;
    SIGNAL S691 : STD_LOGIC;
    SIGNAL S692 : STD_LOGIC;
    SIGNAL S693 : STD_LOGIC;
    SIGNAL S694 : STD_LOGIC;
    SIGNAL S695 : STD_LOGIC;
    SIGNAL S696 : STD_LOGIC;
    SIGNAL S697 : STD_LOGIC;
    SIGNAL S698 : STD_LOGIC;
    SIGNAL S699 : STD_LOGIC;
    SIGNAL S700 : STD_LOGIC;
    SIGNAL S701 : STD_LOGIC;
    SIGNAL S702 : STD_LOGIC;
    SIGNAL S703 : STD_LOGIC;
    SIGNAL S704 : STD_LOGIC;
    SIGNAL S705 : STD_LOGIC;
    SIGNAL S706 : STD_LOGIC;
    SIGNAL S707 : STD_LOGIC;
    SIGNAL S708 : STD_LOGIC;
    SIGNAL S709 : STD_LOGIC;
    SIGNAL S710 : STD_LOGIC;
    SIGNAL S711 : STD_LOGIC;
    SIGNAL S712 : STD_LOGIC;
    SIGNAL S713 : STD_LOGIC;
    SIGNAL S714 : STD_LOGIC;
    SIGNAL S715 : STD_LOGIC;
    SIGNAL S716 : STD_LOGIC;
    SIGNAL S717 : STD_LOGIC;
    SIGNAL S718 : STD_LOGIC;
    SIGNAL S719 : STD_LOGIC;
    SIGNAL S720 : STD_LOGIC;
    SIGNAL S721 : STD_LOGIC;
    SIGNAL S722 : STD_LOGIC;
    SIGNAL S723 : STD_LOGIC;
    SIGNAL S724 : STD_LOGIC;
    SIGNAL S725 : STD_LOGIC;
    SIGNAL S726 : STD_LOGIC;
    SIGNAL S727 : STD_LOGIC;
    SIGNAL S728 : STD_LOGIC;
    SIGNAL S729 : STD_LOGIC;
    SIGNAL S730 : STD_LOGIC;
    SIGNAL S731 : STD_LOGIC;
    SIGNAL S732 : STD_LOGIC;
    SIGNAL S733 : STD_LOGIC;
    SIGNAL S734 : STD_LOGIC;
    SIGNAL S735 : STD_LOGIC;
    SIGNAL S736 : STD_LOGIC;
    SIGNAL S737 : STD_LOGIC;
    SIGNAL S738 : STD_LOGIC;
    SIGNAL S739 : STD_LOGIC;
    SIGNAL S740 : STD_LOGIC;
    SIGNAL S741 : STD_LOGIC;
    SIGNAL S742 : STD_LOGIC;
    SIGNAL S743 : STD_LOGIC;
    SIGNAL S744 : STD_LOGIC;
    SIGNAL S745 : STD_LOGIC;
    SIGNAL S746 : STD_LOGIC;
    SIGNAL S747 : STD_LOGIC;
    SIGNAL S748 : STD_LOGIC;
    SIGNAL S749 : STD_LOGIC;
    SIGNAL S750 : STD_LOGIC;
    SIGNAL S751 : STD_LOGIC;
    SIGNAL S752 : STD_LOGIC;
    SIGNAL S753 : STD_LOGIC;
    SIGNAL S754 : STD_LOGIC;
    SIGNAL S755 : STD_LOGIC;
    SIGNAL S756 : STD_LOGIC;
    SIGNAL S757 : STD_LOGIC;
    SIGNAL S758 : STD_LOGIC;
    SIGNAL S759 : STD_LOGIC;
    SIGNAL S760 : STD_LOGIC;
    SIGNAL S761 : STD_LOGIC;
    SIGNAL S762 : STD_LOGIC;
    SIGNAL S763 : STD_LOGIC;
    SIGNAL S764 : STD_LOGIC;
    SIGNAL S765 : STD_LOGIC;
    SIGNAL S766 : STD_LOGIC;
    SIGNAL S767 : STD_LOGIC;
    SIGNAL S768 : STD_LOGIC;
    SIGNAL S769 : STD_LOGIC;
    SIGNAL S770 : STD_LOGIC;
    SIGNAL S771 : STD_LOGIC;
    SIGNAL S772 : STD_LOGIC;
    SIGNAL S773 : STD_LOGIC;
    SIGNAL S774 : STD_LOGIC;
    SIGNAL S775 : STD_LOGIC;
    SIGNAL S776 : STD_LOGIC;
    SIGNAL S777 : STD_LOGIC;
    SIGNAL S778 : STD_LOGIC;
    SIGNAL S779 : STD_LOGIC;
    SIGNAL S780 : STD_LOGIC;
    SIGNAL S781 : STD_LOGIC;
    SIGNAL S782 : STD_LOGIC;
    SIGNAL S783 : STD_LOGIC;
    SIGNAL S784 : STD_LOGIC;
    SIGNAL S785 : STD_LOGIC;
    SIGNAL S786 : STD_LOGIC;
    SIGNAL S787 : STD_LOGIC;
    SIGNAL S788 : STD_LOGIC;
    SIGNAL S789 : STD_LOGIC;
    SIGNAL S790 : STD_LOGIC;
    SIGNAL S791 : STD_LOGIC;
    SIGNAL S792 : STD_LOGIC;
    SIGNAL S793 : STD_LOGIC;
    SIGNAL S794 : STD_LOGIC;
    SIGNAL S795 : STD_LOGIC;
    SIGNAL S796 : STD_LOGIC;
    SIGNAL S797 : STD_LOGIC;
    SIGNAL S798 : STD_LOGIC;
    SIGNAL S799 : STD_LOGIC;
    SIGNAL S800 : STD_LOGIC;
    SIGNAL S801 : STD_LOGIC;
    SIGNAL S802 : STD_LOGIC;
    SIGNAL S803 : STD_LOGIC;
    SIGNAL S804 : STD_LOGIC;
    SIGNAL S805 : STD_LOGIC;
    SIGNAL S806 : STD_LOGIC;
    SIGNAL S807 : STD_LOGIC;
    SIGNAL S808 : STD_LOGIC;
    SIGNAL S809 : STD_LOGIC;
    SIGNAL S810 : STD_LOGIC;
    SIGNAL S811 : STD_LOGIC;
    SIGNAL S812 : STD_LOGIC;
    SIGNAL S813 : STD_LOGIC;
    SIGNAL S814 : STD_LOGIC;
    SIGNAL S815 : STD_LOGIC;
    SIGNAL S816 : STD_LOGIC;
    SIGNAL S817 : STD_LOGIC;
    SIGNAL S818 : STD_LOGIC;
    SIGNAL S819 : STD_LOGIC;
    SIGNAL S820 : STD_LOGIC;
    SIGNAL S821 : STD_LOGIC;
    SIGNAL S822 : STD_LOGIC;
    SIGNAL S823 : STD_LOGIC;
    SIGNAL S824 : STD_LOGIC;
    SIGNAL S825 : STD_LOGIC;
    SIGNAL S826 : STD_LOGIC;
    SIGNAL S827 : STD_LOGIC;
    SIGNAL S828 : STD_LOGIC;
    SIGNAL S829 : STD_LOGIC;
    SIGNAL S830 : STD_LOGIC;
    SIGNAL S831 : STD_LOGIC;
    SIGNAL S832 : STD_LOGIC;
    SIGNAL S833 : STD_LOGIC;
    SIGNAL S834 : STD_LOGIC;
    SIGNAL S835 : STD_LOGIC;
    SIGNAL S836 : STD_LOGIC;
    SIGNAL S837 : STD_LOGIC;
    SIGNAL S838 : STD_LOGIC;
    SIGNAL S839 : STD_LOGIC;
    SIGNAL S840 : STD_LOGIC;
    SIGNAL S841 : STD_LOGIC;
    SIGNAL S842 : STD_LOGIC;
    SIGNAL S843 : STD_LOGIC;
    SIGNAL S844 : STD_LOGIC;
    SIGNAL S845 : STD_LOGIC;
    SIGNAL S846 : STD_LOGIC;
    SIGNAL S847 : STD_LOGIC;
    SIGNAL S848 : STD_LOGIC;
    SIGNAL S849 : STD_LOGIC;
    SIGNAL S850 : STD_LOGIC;
    SIGNAL S851 : STD_LOGIC;
    SIGNAL S852 : STD_LOGIC;
    SIGNAL S853 : STD_LOGIC;
    SIGNAL S854 : STD_LOGIC;
    SIGNAL S855 : STD_LOGIC;
    SIGNAL S856 : STD_LOGIC;
    SIGNAL S857 : STD_LOGIC;
    SIGNAL S858 : STD_LOGIC;
    SIGNAL S859 : STD_LOGIC;
    SIGNAL S860 : STD_LOGIC;
    SIGNAL S861 : STD_LOGIC;
    SIGNAL S862 : STD_LOGIC;
    SIGNAL S863 : STD_LOGIC;
    SIGNAL S864 : STD_LOGIC;
    SIGNAL S865 : STD_LOGIC;
    SIGNAL S866 : STD_LOGIC;
    SIGNAL S867 : STD_LOGIC;
    SIGNAL S868 : STD_LOGIC;
    SIGNAL S869 : STD_LOGIC;
    SIGNAL S870 : STD_LOGIC;
    SIGNAL S871 : STD_LOGIC;
    SIGNAL S872 : STD_LOGIC;
    SIGNAL S873 : STD_LOGIC;
    SIGNAL S874 : STD_LOGIC;
    SIGNAL S875 : STD_LOGIC;
    SIGNAL S876 : STD_LOGIC;
    SIGNAL S877 : STD_LOGIC;
    SIGNAL S878 : STD_LOGIC;
    SIGNAL S879 : STD_LOGIC;
    SIGNAL S880 : STD_LOGIC;
    SIGNAL S881 : STD_LOGIC;
    SIGNAL S882 : STD_LOGIC;
    SIGNAL S883 : STD_LOGIC;
    SIGNAL S884 : STD_LOGIC;
    SIGNAL S885 : STD_LOGIC;
    SIGNAL S886 : STD_LOGIC;
    SIGNAL S887 : STD_LOGIC;
    SIGNAL S888 : STD_LOGIC;
    SIGNAL S889 : STD_LOGIC;
    SIGNAL S890 : STD_LOGIC;
    SIGNAL S891 : STD_LOGIC;
    SIGNAL S892 : STD_LOGIC;
    SIGNAL S893 : STD_LOGIC;
    SIGNAL S894 : STD_LOGIC;
    SIGNAL S895 : STD_LOGIC;
    SIGNAL S896 : STD_LOGIC;
    SIGNAL S897 : STD_LOGIC;
    SIGNAL S898 : STD_LOGIC;
    SIGNAL S899 : STD_LOGIC;
    SIGNAL S900 : STD_LOGIC;
    SIGNAL S901 : STD_LOGIC;
    SIGNAL S902 : STD_LOGIC;
    SIGNAL S903 : STD_LOGIC;
    SIGNAL S904 : STD_LOGIC;
    SIGNAL S905 : STD_LOGIC;
    SIGNAL S906 : STD_LOGIC;
    SIGNAL S907 : STD_LOGIC;
    SIGNAL S908 : STD_LOGIC;
    SIGNAL S909 : STD_LOGIC;
    SIGNAL S910 : STD_LOGIC;
    SIGNAL S911 : STD_LOGIC;
    SIGNAL S912 : STD_LOGIC;
    SIGNAL S913 : STD_LOGIC;
    SIGNAL S914 : STD_LOGIC;
    SIGNAL S915 : STD_LOGIC;
    SIGNAL S916 : STD_LOGIC;
    SIGNAL S917 : STD_LOGIC;
    SIGNAL S918 : STD_LOGIC;
    SIGNAL S919 : STD_LOGIC;
    SIGNAL S920 : STD_LOGIC;
    SIGNAL S921 : STD_LOGIC;
    SIGNAL S922 : STD_LOGIC;
    SIGNAL S923 : STD_LOGIC;
    SIGNAL S924 : STD_LOGIC;
    SIGNAL S925 : STD_LOGIC;
    SIGNAL S926 : STD_LOGIC;
    SIGNAL S927 : STD_LOGIC;
    SIGNAL S928 : STD_LOGIC;
    SIGNAL S929 : STD_LOGIC;
    SIGNAL S930 : STD_LOGIC;
    SIGNAL S931 : STD_LOGIC;
    SIGNAL S932 : STD_LOGIC;
    SIGNAL S933 : STD_LOGIC;
    SIGNAL S934 : STD_LOGIC;
    SIGNAL S935 : STD_LOGIC;
    SIGNAL S936 : STD_LOGIC;
    SIGNAL S937 : STD_LOGIC;
    SIGNAL S938 : STD_LOGIC;
    SIGNAL S939 : STD_LOGIC;
    SIGNAL S940 : STD_LOGIC;
    SIGNAL S941 : STD_LOGIC;
    SIGNAL S942 : STD_LOGIC;
    SIGNAL S943 : STD_LOGIC;
    SIGNAL S944 : STD_LOGIC;
    SIGNAL S945 : STD_LOGIC;
    SIGNAL S946 : STD_LOGIC;
    SIGNAL S947 : STD_LOGIC;
    SIGNAL S948 : STD_LOGIC;
    SIGNAL S949 : STD_LOGIC;
    SIGNAL S950 : STD_LOGIC;
    SIGNAL S951 : STD_LOGIC;
    SIGNAL S952 : STD_LOGIC;
    SIGNAL S953 : STD_LOGIC;
    SIGNAL S954 : STD_LOGIC;
    SIGNAL S955 : STD_LOGIC;
    SIGNAL S956 : STD_LOGIC;
    SIGNAL S957 : STD_LOGIC;
    SIGNAL S958 : STD_LOGIC;
    SIGNAL S959 : STD_LOGIC;
    SIGNAL S960 : STD_LOGIC;
    SIGNAL S961 : STD_LOGIC;
    SIGNAL S962 : STD_LOGIC;
    SIGNAL S963 : STD_LOGIC;
    SIGNAL S964 : STD_LOGIC;
    SIGNAL S965 : STD_LOGIC;
    SIGNAL S966 : STD_LOGIC;
    SIGNAL S967 : STD_LOGIC;
    SIGNAL S968 : STD_LOGIC;
    SIGNAL S969 : STD_LOGIC;
    SIGNAL S970 : STD_LOGIC;
    SIGNAL S971 : STD_LOGIC;
    SIGNAL S972 : STD_LOGIC;
    SIGNAL S973 : STD_LOGIC;
    SIGNAL S974 : STD_LOGIC;
    SIGNAL S975 : STD_LOGIC;
    SIGNAL S976 : STD_LOGIC;
    SIGNAL S977 : STD_LOGIC;
    SIGNAL S978 : STD_LOGIC;
    SIGNAL S979 : STD_LOGIC;
    SIGNAL S980 : STD_LOGIC;
    SIGNAL S981 : STD_LOGIC;
    SIGNAL S982 : STD_LOGIC;
    SIGNAL S983 : STD_LOGIC;
    SIGNAL S984 : STD_LOGIC;
    SIGNAL S985 : STD_LOGIC;
    SIGNAL S986 : STD_LOGIC;
    SIGNAL S987 : STD_LOGIC;
    SIGNAL S988 : STD_LOGIC;
    SIGNAL S989 : STD_LOGIC;
    SIGNAL S990 : STD_LOGIC;
    SIGNAL S991 : STD_LOGIC;
    SIGNAL S992 : STD_LOGIC;
    SIGNAL S993 : STD_LOGIC;
    SIGNAL S994 : STD_LOGIC;
    SIGNAL S995 : STD_LOGIC;
    SIGNAL S996 : STD_LOGIC;
    SIGNAL S997 : STD_LOGIC;
    SIGNAL S998 : STD_LOGIC;
    SIGNAL S999 : STD_LOGIC;
    SIGNAL S1000 : STD_LOGIC;
    SIGNAL S1001 : STD_LOGIC;
    SIGNAL S1002 : STD_LOGIC;
    SIGNAL S1003 : STD_LOGIC;
    SIGNAL S1004 : STD_LOGIC;
    SIGNAL S1005 : STD_LOGIC;
    SIGNAL S1006 : STD_LOGIC;
    SIGNAL S1007 : STD_LOGIC;
    SIGNAL S1008 : STD_LOGIC;
    SIGNAL S1009 : STD_LOGIC;
    SIGNAL S1010 : STD_LOGIC;
    SIGNAL S1011 : STD_LOGIC;
    SIGNAL S1012 : STD_LOGIC;
    SIGNAL S1013 : STD_LOGIC;
    SIGNAL S1014 : STD_LOGIC;
    SIGNAL S1015 : STD_LOGIC;
    SIGNAL S1016 : STD_LOGIC;
    SIGNAL S1017 : STD_LOGIC;
    SIGNAL S1018 : STD_LOGIC;
    SIGNAL S1019 : STD_LOGIC;
    SIGNAL S1020 : STD_LOGIC;
    SIGNAL S1021 : STD_LOGIC;
    SIGNAL S1022 : STD_LOGIC;
    SIGNAL S1023 : STD_LOGIC;
    SIGNAL S1024 : STD_LOGIC;
    SIGNAL S1025 : STD_LOGIC;
    SIGNAL S1026 : STD_LOGIC;
    SIGNAL S1027 : STD_LOGIC;
    SIGNAL S1028 : STD_LOGIC;
    SIGNAL S1029 : STD_LOGIC;
    SIGNAL S1030 : STD_LOGIC;
    SIGNAL S1031 : STD_LOGIC;
    SIGNAL S1032 : STD_LOGIC;
    SIGNAL S1033 : STD_LOGIC;
    SIGNAL S1034 : STD_LOGIC;
    SIGNAL S1035 : STD_LOGIC;
    SIGNAL S1036 : STD_LOGIC;
    SIGNAL S1037 : STD_LOGIC;
    SIGNAL S1038 : STD_LOGIC;
    SIGNAL S1039 : STD_LOGIC;
    SIGNAL S1040 : STD_LOGIC;
    SIGNAL S1041 : STD_LOGIC;
    SIGNAL S1042 : STD_LOGIC;
    SIGNAL S1043 : STD_LOGIC;
    SIGNAL S1044 : STD_LOGIC;
    SIGNAL S1045 : STD_LOGIC;
    SIGNAL S1046 : STD_LOGIC;
    SIGNAL S1047 : STD_LOGIC;
    SIGNAL S1048 : STD_LOGIC;
    SIGNAL S1049 : STD_LOGIC;
    SIGNAL S1050 : STD_LOGIC;
    SIGNAL S1051 : STD_LOGIC;
    SIGNAL S1052 : STD_LOGIC;
    SIGNAL S1053 : STD_LOGIC;
    SIGNAL S1054 : STD_LOGIC;
    SIGNAL S1055 : STD_LOGIC;
    SIGNAL S1056 : STD_LOGIC;
    SIGNAL S1057 : STD_LOGIC;
    SIGNAL S1058 : STD_LOGIC;
    SIGNAL S1059 : STD_LOGIC;
    SIGNAL S1060 : STD_LOGIC;
    SIGNAL S1061 : STD_LOGIC;
    SIGNAL S1062 : STD_LOGIC;
    SIGNAL S1063 : STD_LOGIC;
    SIGNAL S1064 : STD_LOGIC;
    SIGNAL S1065 : STD_LOGIC;
    SIGNAL S1066 : STD_LOGIC;
    SIGNAL S1067 : STD_LOGIC;
    SIGNAL S1068 : STD_LOGIC;
    SIGNAL S1069 : STD_LOGIC;
    SIGNAL S1070 : STD_LOGIC;
    SIGNAL S1071 : STD_LOGIC;
    SIGNAL S1072 : STD_LOGIC;
    SIGNAL S1073 : STD_LOGIC;
    SIGNAL S1074 : STD_LOGIC;
    SIGNAL S1075 : STD_LOGIC;
    SIGNAL S1076 : STD_LOGIC;
    SIGNAL S1077 : STD_LOGIC;
    SIGNAL S1078 : STD_LOGIC;
    SIGNAL S1079 : STD_LOGIC;
    SIGNAL S1080 : STD_LOGIC;
    SIGNAL S1081 : STD_LOGIC;
    SIGNAL S1082 : STD_LOGIC;
    SIGNAL S1083 : STD_LOGIC;
    SIGNAL S1084 : STD_LOGIC;
    SIGNAL S1085 : STD_LOGIC;
    SIGNAL S1086 : STD_LOGIC;
    SIGNAL S1087 : STD_LOGIC;
    SIGNAL S1088 : STD_LOGIC;
    SIGNAL S1089 : STD_LOGIC;
    SIGNAL S1090 : STD_LOGIC;
    SIGNAL S1091 : STD_LOGIC;
    SIGNAL S1092 : STD_LOGIC;
    SIGNAL S1093 : STD_LOGIC;
    SIGNAL S1094 : STD_LOGIC;
    SIGNAL S1095 : STD_LOGIC;
    SIGNAL S1096 : STD_LOGIC;
    SIGNAL S1097 : STD_LOGIC;
    SIGNAL S1098 : STD_LOGIC;
    SIGNAL S1099 : STD_LOGIC;
    SIGNAL S1100 : STD_LOGIC;
    SIGNAL S1101 : STD_LOGIC;
    SIGNAL S1102 : STD_LOGIC;
    SIGNAL S1103 : STD_LOGIC;
    SIGNAL S1104 : STD_LOGIC;
    SIGNAL S1105 : STD_LOGIC;
    SIGNAL S1106 : STD_LOGIC;
    SIGNAL S1107 : STD_LOGIC;
    SIGNAL S1108 : STD_LOGIC;
    SIGNAL S1109 : STD_LOGIC;
    SIGNAL S1110 : STD_LOGIC;
    SIGNAL S1111 : STD_LOGIC;
    SIGNAL S1112 : STD_LOGIC;
    SIGNAL S1113 : STD_LOGIC;
    SIGNAL S1114 : STD_LOGIC;
    SIGNAL S1115 : STD_LOGIC;
    SIGNAL S1116 : STD_LOGIC;
    SIGNAL S1117 : STD_LOGIC;
    SIGNAL S1118 : STD_LOGIC;
    SIGNAL S1119 : STD_LOGIC;
    SIGNAL S1120 : STD_LOGIC;
    SIGNAL S1121 : STD_LOGIC;
    SIGNAL S1122 : STD_LOGIC;
    SIGNAL S1123 : STD_LOGIC;
    SIGNAL S1124 : STD_LOGIC;
    SIGNAL S1125 : STD_LOGIC;
    SIGNAL S1126 : STD_LOGIC;
    SIGNAL S1127 : STD_LOGIC;
    SIGNAL S1128 : STD_LOGIC;
    SIGNAL S1129 : STD_LOGIC;
    SIGNAL S1130 : STD_LOGIC;
    SIGNAL S1131 : STD_LOGIC;
    SIGNAL S1132 : STD_LOGIC;
    SIGNAL S1133 : STD_LOGIC;
    SIGNAL S1134 : STD_LOGIC;
    SIGNAL S1135 : STD_LOGIC;
    SIGNAL S1136 : STD_LOGIC;
    SIGNAL S1137 : STD_LOGIC;
    SIGNAL S1138 : STD_LOGIC;
    SIGNAL S1139 : STD_LOGIC;
    SIGNAL S1140 : STD_LOGIC;
    SIGNAL S1141 : STD_LOGIC;
    SIGNAL S1142 : STD_LOGIC;
    SIGNAL S1143 : STD_LOGIC;
    SIGNAL S1144 : STD_LOGIC;
    SIGNAL S1145 : STD_LOGIC;
    SIGNAL S1146 : STD_LOGIC;
    SIGNAL S1147 : STD_LOGIC;
    SIGNAL S1148 : STD_LOGIC;
    SIGNAL S1149 : STD_LOGIC;
    SIGNAL S1150 : STD_LOGIC;
    SIGNAL S1151 : STD_LOGIC;
    SIGNAL S1152 : STD_LOGIC;
    SIGNAL S1153 : STD_LOGIC;
    SIGNAL S1154 : STD_LOGIC;
    SIGNAL S1155 : STD_LOGIC;
    SIGNAL S1156 : STD_LOGIC;
    SIGNAL S1157 : STD_LOGIC;
    SIGNAL S1158 : STD_LOGIC;
    SIGNAL S1159 : STD_LOGIC;
    SIGNAL S1160 : STD_LOGIC;
    SIGNAL S1161 : STD_LOGIC;
    SIGNAL S1162 : STD_LOGIC;
    SIGNAL S1163 : STD_LOGIC;
    SIGNAL S1164 : STD_LOGIC;
    SIGNAL S1165 : STD_LOGIC;
    SIGNAL S1166 : STD_LOGIC;
    SIGNAL S1167 : STD_LOGIC;
    SIGNAL S1168 : STD_LOGIC;
    SIGNAL S1169 : STD_LOGIC;
    SIGNAL S1170 : STD_LOGIC;
    SIGNAL S1171 : STD_LOGIC;
    SIGNAL S1172 : STD_LOGIC;
    SIGNAL S1173 : STD_LOGIC;
    SIGNAL S1174 : STD_LOGIC;
    SIGNAL S1175 : STD_LOGIC;
    SIGNAL S1176 : STD_LOGIC;
    SIGNAL S1177 : STD_LOGIC;
    SIGNAL S1178 : STD_LOGIC;
    SIGNAL S1179 : STD_LOGIC;
    SIGNAL S1180 : STD_LOGIC;
    SIGNAL S1181 : STD_LOGIC;
    SIGNAL S1182 : STD_LOGIC;
    SIGNAL S1183 : STD_LOGIC;
    SIGNAL S1184 : STD_LOGIC;
    SIGNAL S1185 : STD_LOGIC;
    SIGNAL S1186 : STD_LOGIC;
    SIGNAL S1187 : STD_LOGIC;
    SIGNAL S1188 : STD_LOGIC;
    SIGNAL S1189 : STD_LOGIC;
    SIGNAL S1190 : STD_LOGIC;
    SIGNAL S1191 : STD_LOGIC;
    SIGNAL S1192 : STD_LOGIC;
    SIGNAL S1193 : STD_LOGIC;
    SIGNAL S1194 : STD_LOGIC;
    SIGNAL S1195 : STD_LOGIC;
    SIGNAL S1196 : STD_LOGIC;
    SIGNAL S1197 : STD_LOGIC;
    SIGNAL S1198 : STD_LOGIC;
    SIGNAL S1199 : STD_LOGIC;
    SIGNAL S1200 : STD_LOGIC;
    SIGNAL S1201 : STD_LOGIC;
    SIGNAL S1202 : STD_LOGIC;
    SIGNAL S1203 : STD_LOGIC;
    SIGNAL S1204 : STD_LOGIC;
    SIGNAL S1205 : STD_LOGIC;
    SIGNAL S1206 : STD_LOGIC;
    SIGNAL S1207 : STD_LOGIC;
    SIGNAL S1208 : STD_LOGIC;
    SIGNAL S1209 : STD_LOGIC;
    SIGNAL S1210 : STD_LOGIC;
    SIGNAL S1211 : STD_LOGIC;
    SIGNAL S1212 : STD_LOGIC;
    SIGNAL S1213 : STD_LOGIC;
    SIGNAL S1214 : STD_LOGIC;
    SIGNAL S1215 : STD_LOGIC;
    SIGNAL S1216 : STD_LOGIC;
    SIGNAL S1217 : STD_LOGIC;
    SIGNAL S1218 : STD_LOGIC;
    SIGNAL S1219 : STD_LOGIC;
    SIGNAL S1220 : STD_LOGIC;
    SIGNAL S1221 : STD_LOGIC;
    SIGNAL S1222 : STD_LOGIC;
    SIGNAL S1223 : STD_LOGIC;
    SIGNAL S1224 : STD_LOGIC;
    SIGNAL S1225 : STD_LOGIC;
    SIGNAL S1226 : STD_LOGIC;
    SIGNAL S1227 : STD_LOGIC;
    SIGNAL S1228 : STD_LOGIC;
    SIGNAL S1229 : STD_LOGIC;
    SIGNAL S1230 : STD_LOGIC;
    SIGNAL S1231 : STD_LOGIC;
    SIGNAL S1232 : STD_LOGIC;
    SIGNAL S1233 : STD_LOGIC;
    SIGNAL S1234 : STD_LOGIC;
    SIGNAL S1235 : STD_LOGIC;
    SIGNAL S1236 : STD_LOGIC;
    SIGNAL S1237 : STD_LOGIC;
    SIGNAL S1238 : STD_LOGIC;
    SIGNAL S1239 : STD_LOGIC;
    SIGNAL S1240 : STD_LOGIC;
    SIGNAL S1241 : STD_LOGIC;
    SIGNAL S1242 : STD_LOGIC;
    SIGNAL S1243 : STD_LOGIC;
    SIGNAL S1244 : STD_LOGIC;
    SIGNAL S1245 : STD_LOGIC;
    SIGNAL S1246 : STD_LOGIC;
    SIGNAL S1247 : STD_LOGIC;
    SIGNAL S1248 : STD_LOGIC;
    SIGNAL S1249 : STD_LOGIC;
    SIGNAL S1250 : STD_LOGIC;
    SIGNAL S1251 : STD_LOGIC;
    SIGNAL S1252 : STD_LOGIC;
    SIGNAL S1253 : STD_LOGIC;
    SIGNAL S1254 : STD_LOGIC;
    SIGNAL S1255 : STD_LOGIC;
    SIGNAL S1256 : STD_LOGIC;
    SIGNAL S1257 : STD_LOGIC;
    SIGNAL S1258 : STD_LOGIC;
    SIGNAL S1259 : STD_LOGIC;
    SIGNAL S1260 : STD_LOGIC;
    SIGNAL S1261 : STD_LOGIC;
    SIGNAL S1262 : STD_LOGIC;
    SIGNAL S1263 : STD_LOGIC;
    SIGNAL S1264 : STD_LOGIC;
    SIGNAL S1265 : STD_LOGIC;
    SIGNAL S1266 : STD_LOGIC;
    SIGNAL S1267 : STD_LOGIC;
    SIGNAL S1268 : STD_LOGIC;
    SIGNAL S1269 : STD_LOGIC;
    SIGNAL S1270 : STD_LOGIC;
    SIGNAL S1271 : STD_LOGIC;
    SIGNAL S1272 : STD_LOGIC;
    SIGNAL S1273 : STD_LOGIC;
    SIGNAL S1274 : STD_LOGIC;
    SIGNAL S1275 : STD_LOGIC;
    SIGNAL S1276 : STD_LOGIC;
    SIGNAL S1277 : STD_LOGIC;
    SIGNAL S1278 : STD_LOGIC;
    SIGNAL S1279 : STD_LOGIC;
    SIGNAL S1280 : STD_LOGIC;
    SIGNAL S1281 : STD_LOGIC;
    SIGNAL S1282 : STD_LOGIC;
    SIGNAL S1283 : STD_LOGIC;
    SIGNAL S1284 : STD_LOGIC;
    SIGNAL S1285 : STD_LOGIC;
    SIGNAL S1286 : STD_LOGIC;
    SIGNAL S1287 : STD_LOGIC;
    SIGNAL S1288 : STD_LOGIC;
    SIGNAL S1289 : STD_LOGIC;
    SIGNAL S1290 : STD_LOGIC;
    SIGNAL S1291 : STD_LOGIC;
    SIGNAL S1292 : STD_LOGIC;
    SIGNAL S1293 : STD_LOGIC;
    SIGNAL S1294 : STD_LOGIC;
    SIGNAL S1295 : STD_LOGIC;
    SIGNAL S1296 : STD_LOGIC;
    SIGNAL S1297 : STD_LOGIC;
    SIGNAL S1298 : STD_LOGIC;
    SIGNAL S1299 : STD_LOGIC;
    SIGNAL S1300 : STD_LOGIC;
    SIGNAL S1301 : STD_LOGIC;
    SIGNAL S1302 : STD_LOGIC;
    SIGNAL S1303 : STD_LOGIC;
    SIGNAL S1304 : STD_LOGIC;
    SIGNAL S1305 : STD_LOGIC;
    SIGNAL S1306 : STD_LOGIC;
    SIGNAL S1307 : STD_LOGIC;
    SIGNAL S1308 : STD_LOGIC;
    SIGNAL S1309 : STD_LOGIC;
    SIGNAL S1310 : STD_LOGIC;
    SIGNAL S1311 : STD_LOGIC;
    SIGNAL S1312 : STD_LOGIC;
    SIGNAL S1313 : STD_LOGIC;
    SIGNAL S1314 : STD_LOGIC;
    SIGNAL S1315 : STD_LOGIC;
    SIGNAL S1316 : STD_LOGIC;
    SIGNAL S1317 : STD_LOGIC;
    SIGNAL S1318 : STD_LOGIC;
    SIGNAL S1319 : STD_LOGIC;
    SIGNAL S1320 : STD_LOGIC;
    SIGNAL S1321 : STD_LOGIC;
    SIGNAL S1322 : STD_LOGIC;
    SIGNAL S1323 : STD_LOGIC;
    SIGNAL S1324 : STD_LOGIC;
    SIGNAL S1325 : STD_LOGIC;
    SIGNAL S1326 : STD_LOGIC;
    SIGNAL S1327 : STD_LOGIC;
    SIGNAL S1328 : STD_LOGIC;
    SIGNAL S1329 : STD_LOGIC;
    SIGNAL S1330 : STD_LOGIC;
    SIGNAL S1331 : STD_LOGIC;
    SIGNAL S1332 : STD_LOGIC;
    SIGNAL S1333 : STD_LOGIC;
    SIGNAL S1334 : STD_LOGIC;
    SIGNAL S1335 : STD_LOGIC;
    SIGNAL S1336 : STD_LOGIC;
    SIGNAL S1337 : STD_LOGIC;
    SIGNAL S1338 : STD_LOGIC;
    SIGNAL S1339 : STD_LOGIC;
    SIGNAL S1340 : STD_LOGIC;
    SIGNAL S1341 : STD_LOGIC;
    SIGNAL S1342 : STD_LOGIC;
    SIGNAL S1343 : STD_LOGIC;
    SIGNAL S1344 : STD_LOGIC;
    SIGNAL S1345 : STD_LOGIC;
    SIGNAL S1346 : STD_LOGIC;
    SIGNAL S1347 : STD_LOGIC;
    SIGNAL S1348 : STD_LOGIC;
    SIGNAL S1349 : STD_LOGIC;
    SIGNAL S1350 : STD_LOGIC;
    SIGNAL S1351 : STD_LOGIC;
    SIGNAL S1352 : STD_LOGIC;
    SIGNAL S1353 : STD_LOGIC;
    SIGNAL S1354 : STD_LOGIC;
    SIGNAL S1355 : STD_LOGIC;
    SIGNAL S1356 : STD_LOGIC;
    SIGNAL S1357 : STD_LOGIC;
    SIGNAL S1358 : STD_LOGIC;
    SIGNAL S1359 : STD_LOGIC;
    SIGNAL S1360 : STD_LOGIC;
    SIGNAL S1361 : STD_LOGIC;
    SIGNAL S1362 : STD_LOGIC;
    SIGNAL S1363 : STD_LOGIC;
    SIGNAL S1364 : STD_LOGIC;
    SIGNAL S1365 : STD_LOGIC;
    SIGNAL S1366 : STD_LOGIC;
    SIGNAL S1367 : STD_LOGIC;
    SIGNAL S1368 : STD_LOGIC;
    SIGNAL S1369 : STD_LOGIC;
    SIGNAL S1370 : STD_LOGIC;
    SIGNAL S1371 : STD_LOGIC;
    SIGNAL S1372 : STD_LOGIC;
    SIGNAL S1373 : STD_LOGIC;
    SIGNAL S1374 : STD_LOGIC;
    SIGNAL S1375 : STD_LOGIC;
    SIGNAL S1376 : STD_LOGIC;
    SIGNAL S1377 : STD_LOGIC;
    SIGNAL S1378 : STD_LOGIC;
    SIGNAL S1379 : STD_LOGIC;
    SIGNAL S1380 : STD_LOGIC;
    SIGNAL S1381 : STD_LOGIC;
    SIGNAL S1382 : STD_LOGIC;
    SIGNAL S1383 : STD_LOGIC;
    SIGNAL S1384 : STD_LOGIC;
    SIGNAL S1385 : STD_LOGIC;
    SIGNAL S1386 : STD_LOGIC;
    SIGNAL S1387 : STD_LOGIC;
    SIGNAL S1388 : STD_LOGIC;
    SIGNAL S1389 : STD_LOGIC;
    SIGNAL S1390 : STD_LOGIC;
    SIGNAL S1391 : STD_LOGIC;
    SIGNAL S1392 : STD_LOGIC;
    SIGNAL S1393 : STD_LOGIC;
    SIGNAL S1394 : STD_LOGIC;
    SIGNAL S1395 : STD_LOGIC;
    SIGNAL S1396 : STD_LOGIC;
    SIGNAL S1397 : STD_LOGIC;
    SIGNAL S1398 : STD_LOGIC;
    SIGNAL S1399 : STD_LOGIC;
    SIGNAL S1400 : STD_LOGIC;
    SIGNAL S1401 : STD_LOGIC;
    SIGNAL S1402 : STD_LOGIC;
    SIGNAL S1403 : STD_LOGIC;
    SIGNAL S1404 : STD_LOGIC;
    SIGNAL S1405 : STD_LOGIC;
    SIGNAL S1406 : STD_LOGIC;
    SIGNAL S1407 : STD_LOGIC;
    SIGNAL S1408 : STD_LOGIC;
    SIGNAL S1409 : STD_LOGIC;
    SIGNAL S1410 : STD_LOGIC;
    SIGNAL S1411 : STD_LOGIC;
    SIGNAL S1412 : STD_LOGIC;
    SIGNAL S1413 : STD_LOGIC;
    SIGNAL S1414 : STD_LOGIC;
    SIGNAL S1415 : STD_LOGIC;
    SIGNAL S1416 : STD_LOGIC;
    SIGNAL S1417 : STD_LOGIC;
    SIGNAL S1418 : STD_LOGIC;
    SIGNAL S1419 : STD_LOGIC;
    SIGNAL S1420 : STD_LOGIC;
    SIGNAL S1421 : STD_LOGIC;
    SIGNAL S1422 : STD_LOGIC;
    SIGNAL S1423 : STD_LOGIC;
    SIGNAL S1424 : STD_LOGIC;
    SIGNAL S1425 : STD_LOGIC;
    SIGNAL S1426 : STD_LOGIC;
    SIGNAL S1427 : STD_LOGIC;
    SIGNAL S1428 : STD_LOGIC;
    SIGNAL S1429 : STD_LOGIC;
    SIGNAL S1430 : STD_LOGIC;
    SIGNAL S1431 : STD_LOGIC;
    SIGNAL S1432 : STD_LOGIC;
    SIGNAL S1433 : STD_LOGIC;
    SIGNAL S1434 : STD_LOGIC;
    SIGNAL S1435 : STD_LOGIC;
    SIGNAL S1436 : STD_LOGIC;
    SIGNAL S1437 : STD_LOGIC;
    SIGNAL S1438 : STD_LOGIC;
    SIGNAL S1439 : STD_LOGIC;
    SIGNAL S1440 : STD_LOGIC;
    SIGNAL S1441 : STD_LOGIC;
    SIGNAL S1442 : STD_LOGIC;
    SIGNAL S1443 : STD_LOGIC;
    SIGNAL S1444 : STD_LOGIC;
    SIGNAL S1445 : STD_LOGIC;
    SIGNAL S1446 : STD_LOGIC;
    SIGNAL S1447 : STD_LOGIC;
    SIGNAL S1448 : STD_LOGIC;
    SIGNAL S1449 : STD_LOGIC;
    SIGNAL S1450 : STD_LOGIC;
    SIGNAL S1451 : STD_LOGIC;
    SIGNAL S1452 : STD_LOGIC;
    SIGNAL S1453 : STD_LOGIC;
    SIGNAL S1454 : STD_LOGIC;
    SIGNAL S1455 : STD_LOGIC;
    SIGNAL S1456 : STD_LOGIC;
    SIGNAL S1457 : STD_LOGIC;
    SIGNAL S1458 : STD_LOGIC;
    SIGNAL S1459 : STD_LOGIC;
    SIGNAL S1460 : STD_LOGIC;
    SIGNAL S1461 : STD_LOGIC;
    SIGNAL S1462 : STD_LOGIC;
    SIGNAL S1463 : STD_LOGIC;
    SIGNAL S1464 : STD_LOGIC;
    SIGNAL S1465 : STD_LOGIC;
    SIGNAL S1466 : STD_LOGIC;
    SIGNAL S1467 : STD_LOGIC;
    SIGNAL S1468 : STD_LOGIC;
    SIGNAL S1469 : STD_LOGIC;
    SIGNAL S1470 : STD_LOGIC;
    SIGNAL S1471 : STD_LOGIC;
    SIGNAL S1472 : STD_LOGIC;
    SIGNAL S1473 : STD_LOGIC;
    SIGNAL S1474 : STD_LOGIC;
    SIGNAL S1475 : STD_LOGIC;
    SIGNAL S1476 : STD_LOGIC;
    SIGNAL S1477 : STD_LOGIC;
    SIGNAL S1478 : STD_LOGIC;
    SIGNAL S1479 : STD_LOGIC;
    SIGNAL S1480 : STD_LOGIC;
    SIGNAL S1481 : STD_LOGIC;
    SIGNAL S1482 : STD_LOGIC;
    SIGNAL S1483 : STD_LOGIC;
    SIGNAL S1484 : STD_LOGIC;
    SIGNAL S1485 : STD_LOGIC;
    SIGNAL S1486 : STD_LOGIC;
    SIGNAL S1487 : STD_LOGIC;
    SIGNAL S1488 : STD_LOGIC;
    SIGNAL S1489 : STD_LOGIC;
    SIGNAL S1490 : STD_LOGIC;
    SIGNAL S1491 : STD_LOGIC;
    SIGNAL S1492 : STD_LOGIC;
    SIGNAL S1493 : STD_LOGIC;
    SIGNAL S1494 : STD_LOGIC;
    SIGNAL S1495 : STD_LOGIC;
    SIGNAL S1496 : STD_LOGIC;
    SIGNAL S1497 : STD_LOGIC;
    SIGNAL S1498 : STD_LOGIC;
    SIGNAL S1499 : STD_LOGIC;
    SIGNAL S1500 : STD_LOGIC;
    SIGNAL S1501 : STD_LOGIC;
    SIGNAL S1502 : STD_LOGIC;
    SIGNAL S1503 : STD_LOGIC;
    SIGNAL S1504 : STD_LOGIC;
    SIGNAL S1505 : STD_LOGIC;
    SIGNAL S1506 : STD_LOGIC;
    SIGNAL S1507 : STD_LOGIC;
    SIGNAL S1508 : STD_LOGIC;
    SIGNAL S1509 : STD_LOGIC;
    SIGNAL S1510 : STD_LOGIC;
    SIGNAL S1511 : STD_LOGIC;
    SIGNAL S1512 : STD_LOGIC;
    SIGNAL S1513 : STD_LOGIC;
    SIGNAL S1514 : STD_LOGIC;
    SIGNAL S1515 : STD_LOGIC;
    SIGNAL S1516 : STD_LOGIC;
    SIGNAL S1517 : STD_LOGIC;
    SIGNAL S1518 : STD_LOGIC;
    SIGNAL S1519 : STD_LOGIC;
    SIGNAL S1520 : STD_LOGIC;
    SIGNAL S1521 : STD_LOGIC;
    SIGNAL S1522 : STD_LOGIC;
    SIGNAL S1523 : STD_LOGIC;
    SIGNAL S1524 : STD_LOGIC;
    SIGNAL S1525 : STD_LOGIC;
    SIGNAL S1526 : STD_LOGIC;
    SIGNAL S1527 : STD_LOGIC;
    SIGNAL S1528 : STD_LOGIC;
    SIGNAL S1529 : STD_LOGIC;
    SIGNAL S1530 : STD_LOGIC;
    SIGNAL S1531 : STD_LOGIC;
    SIGNAL S1532 : STD_LOGIC;
    SIGNAL S1533 : STD_LOGIC;
    SIGNAL S1534 : STD_LOGIC;
    SIGNAL S1535 : STD_LOGIC;
    SIGNAL S1536 : STD_LOGIC;
    SIGNAL S1537 : STD_LOGIC;
    SIGNAL S1538 : STD_LOGIC;
    SIGNAL S1539 : STD_LOGIC;
    SIGNAL S1540 : STD_LOGIC;
    SIGNAL S1541 : STD_LOGIC;
    SIGNAL S1542 : STD_LOGIC;
    SIGNAL S1543 : STD_LOGIC;
    SIGNAL S1544 : STD_LOGIC;
    SIGNAL S1545 : STD_LOGIC;
    SIGNAL S1546 : STD_LOGIC;
    SIGNAL S1547 : STD_LOGIC;
    SIGNAL S1548 : STD_LOGIC;
    SIGNAL S1549 : STD_LOGIC;
    SIGNAL S1550 : STD_LOGIC;
    SIGNAL S1551 : STD_LOGIC;
    SIGNAL S1552 : STD_LOGIC;
    SIGNAL S1553 : STD_LOGIC;
    SIGNAL S1554 : STD_LOGIC;
    SIGNAL S1555 : STD_LOGIC;
    SIGNAL S1556 : STD_LOGIC;
    SIGNAL S1557 : STD_LOGIC;
    SIGNAL S1558 : STD_LOGIC;
    SIGNAL S1559 : STD_LOGIC;
    SIGNAL S1560 : STD_LOGIC;
    SIGNAL S1561 : STD_LOGIC;
    SIGNAL S1562 : STD_LOGIC;
    SIGNAL S1563 : STD_LOGIC;
    SIGNAL S1564 : STD_LOGIC;
    SIGNAL S1565 : STD_LOGIC;
    SIGNAL S1566 : STD_LOGIC;
    SIGNAL S1567 : STD_LOGIC;
    SIGNAL S1568 : STD_LOGIC;
    SIGNAL S1569 : STD_LOGIC;
    SIGNAL S1570 : STD_LOGIC;
    SIGNAL S1571 : STD_LOGIC;
    SIGNAL S1572 : STD_LOGIC;
    SIGNAL S1573 : STD_LOGIC;
    SIGNAL S1574 : STD_LOGIC;
    SIGNAL S1575 : STD_LOGIC;
    SIGNAL S1576 : STD_LOGIC;
    SIGNAL S1577 : STD_LOGIC;
    SIGNAL S1578 : STD_LOGIC;
    SIGNAL S1579 : STD_LOGIC;
    SIGNAL S1580 : STD_LOGIC;
    SIGNAL S1581 : STD_LOGIC;
    SIGNAL S1582 : STD_LOGIC;
    SIGNAL S1583 : STD_LOGIC;
    SIGNAL S1584 : STD_LOGIC;
    SIGNAL S1585 : STD_LOGIC;
    SIGNAL S1586 : STD_LOGIC;
    SIGNAL S1587 : STD_LOGIC;
    SIGNAL S1588 : STD_LOGIC;
    SIGNAL S1589 : STD_LOGIC;
    SIGNAL S1590 : STD_LOGIC;
    SIGNAL S1591 : STD_LOGIC;
    SIGNAL S1592 : STD_LOGIC;
    SIGNAL S1593 : STD_LOGIC;
    SIGNAL S1594 : STD_LOGIC;
    SIGNAL S1595 : STD_LOGIC;
    SIGNAL S1596 : STD_LOGIC;
    SIGNAL S1597 : STD_LOGIC;
    SIGNAL S1598 : STD_LOGIC;
    SIGNAL S1599 : STD_LOGIC;
    SIGNAL S1600 : STD_LOGIC;
    SIGNAL S1601 : STD_LOGIC;
    SIGNAL S1602 : STD_LOGIC;
    SIGNAL S1603 : STD_LOGIC;
    SIGNAL S1604 : STD_LOGIC;
    SIGNAL S1605 : STD_LOGIC;
    SIGNAL S1606 : STD_LOGIC;
    SIGNAL S1607 : STD_LOGIC;
    SIGNAL S1608 : STD_LOGIC;
    SIGNAL S1609 : STD_LOGIC;
    SIGNAL S1610 : STD_LOGIC;
    SIGNAL S1611 : STD_LOGIC;
    SIGNAL S1612 : STD_LOGIC;
    SIGNAL S1613 : STD_LOGIC;
    SIGNAL S1614 : STD_LOGIC;
    SIGNAL S1615 : STD_LOGIC;
    SIGNAL S1616 : STD_LOGIC;
    SIGNAL S1617 : STD_LOGIC;
    SIGNAL S1618 : STD_LOGIC;
    SIGNAL S1619 : STD_LOGIC;
    SIGNAL S1620 : STD_LOGIC;
    SIGNAL S1621 : STD_LOGIC;
    SIGNAL S1622 : STD_LOGIC;
    SIGNAL S1623 : STD_LOGIC;
    SIGNAL S1624 : STD_LOGIC;
    SIGNAL S1625 : STD_LOGIC;
    SIGNAL S1626 : STD_LOGIC;
    SIGNAL S1627 : STD_LOGIC;
    SIGNAL S1628 : STD_LOGIC;
    SIGNAL S1629 : STD_LOGIC;
    SIGNAL S1630 : STD_LOGIC;
    SIGNAL S1631 : STD_LOGIC;
    SIGNAL S1632 : STD_LOGIC;
    SIGNAL S1633 : STD_LOGIC;
    SIGNAL S1634 : STD_LOGIC;
    SIGNAL S1635 : STD_LOGIC;
    SIGNAL S1636 : STD_LOGIC;
    SIGNAL S1637 : STD_LOGIC;
    SIGNAL S1638 : STD_LOGIC;
    SIGNAL S1639 : STD_LOGIC;
    SIGNAL S1640 : STD_LOGIC;
    SIGNAL S1641 : STD_LOGIC;
    SIGNAL S1642 : STD_LOGIC;
    SIGNAL S1643 : STD_LOGIC;
    SIGNAL S1644 : STD_LOGIC;
    SIGNAL S1645 : STD_LOGIC;
    SIGNAL S1646 : STD_LOGIC;
    SIGNAL S1647 : STD_LOGIC;
    SIGNAL S1648 : STD_LOGIC;
    SIGNAL S1649 : STD_LOGIC;
    SIGNAL S1650 : STD_LOGIC;
    SIGNAL S1651 : STD_LOGIC;
    SIGNAL S1652 : STD_LOGIC;
    SIGNAL S1653 : STD_LOGIC;
    SIGNAL S1654 : STD_LOGIC;
    SIGNAL S1655 : STD_LOGIC;
    SIGNAL S1656 : STD_LOGIC;
    SIGNAL S1657 : STD_LOGIC;
    SIGNAL S1658 : STD_LOGIC;
    SIGNAL S1659 : STD_LOGIC;
    SIGNAL S1660 : STD_LOGIC;
    SIGNAL S1661 : STD_LOGIC;
    SIGNAL S1662 : STD_LOGIC;
    SIGNAL S1663 : STD_LOGIC;
    SIGNAL S1664 : STD_LOGIC;
    SIGNAL S1665 : STD_LOGIC;
    SIGNAL S1666 : STD_LOGIC;
    SIGNAL S1667 : STD_LOGIC;
    SIGNAL S1668 : STD_LOGIC;
    SIGNAL S1669 : STD_LOGIC;
    SIGNAL S1670 : STD_LOGIC;
    SIGNAL S1671 : STD_LOGIC;
    SIGNAL S1672 : STD_LOGIC;
    SIGNAL S1673 : STD_LOGIC;
    SIGNAL S1674 : STD_LOGIC;
    SIGNAL S1675 : STD_LOGIC;
    SIGNAL S1676 : STD_LOGIC;
    SIGNAL S1677 : STD_LOGIC;
    SIGNAL S1678 : STD_LOGIC;
    SIGNAL S1679 : STD_LOGIC;
    SIGNAL S1680 : STD_LOGIC;
    SIGNAL S1681 : STD_LOGIC;
    SIGNAL S1682 : STD_LOGIC;
    SIGNAL S1683 : STD_LOGIC;
    SIGNAL S1684 : STD_LOGIC;
    SIGNAL S1685 : STD_LOGIC;
    SIGNAL S1686 : STD_LOGIC;
    SIGNAL S1687 : STD_LOGIC;
    SIGNAL S1688 : STD_LOGIC;
    SIGNAL S1689 : STD_LOGIC;
    SIGNAL S1690 : STD_LOGIC;
    SIGNAL S1691 : STD_LOGIC;
    SIGNAL S1692 : STD_LOGIC;
    SIGNAL S1693 : STD_LOGIC;
    SIGNAL S1694 : STD_LOGIC;
    SIGNAL S1695 : STD_LOGIC;
    SIGNAL S1696 : STD_LOGIC;
    SIGNAL S1697 : STD_LOGIC;
    SIGNAL S1698 : STD_LOGIC;
    SIGNAL S1699 : STD_LOGIC;
    SIGNAL S1700 : STD_LOGIC;
    SIGNAL S1701 : STD_LOGIC;
    SIGNAL S1702 : STD_LOGIC;
    SIGNAL S1703 : STD_LOGIC;
    SIGNAL S1704 : STD_LOGIC;
    SIGNAL S1705 : STD_LOGIC;
    SIGNAL S1706 : STD_LOGIC;
    SIGNAL S1707 : STD_LOGIC;
    SIGNAL S1708 : STD_LOGIC;
    SIGNAL S1709 : STD_LOGIC;
    SIGNAL S1710 : STD_LOGIC;
    SIGNAL S1711 : STD_LOGIC;
    SIGNAL S1712 : STD_LOGIC;
    SIGNAL S1713 : STD_LOGIC;
    SIGNAL S1714 : STD_LOGIC;
    SIGNAL S1715 : STD_LOGIC;
    SIGNAL S1716 : STD_LOGIC;
    SIGNAL S1717 : STD_LOGIC;
    SIGNAL S1718 : STD_LOGIC;
    SIGNAL S1719 : STD_LOGIC;
    SIGNAL S1720 : STD_LOGIC;
    SIGNAL S1721 : STD_LOGIC;
    SIGNAL S1722 : STD_LOGIC;
    SIGNAL S1723 : STD_LOGIC;
    SIGNAL S1724 : STD_LOGIC;
    SIGNAL S1725 : STD_LOGIC;
    SIGNAL S1726 : STD_LOGIC;
    SIGNAL S1727 : STD_LOGIC;
    SIGNAL S1728 : STD_LOGIC;
    SIGNAL S1729 : STD_LOGIC;
    SIGNAL S1730 : STD_LOGIC;
    SIGNAL S1731 : STD_LOGIC;
    SIGNAL S1732 : STD_LOGIC;
    SIGNAL S1733 : STD_LOGIC;
    SIGNAL S1734 : STD_LOGIC;
    SIGNAL S1735 : STD_LOGIC;
    SIGNAL S1736 : STD_LOGIC;
    SIGNAL S1737 : STD_LOGIC;
    SIGNAL S1738 : STD_LOGIC;
    SIGNAL S1739 : STD_LOGIC;
    SIGNAL S1740 : STD_LOGIC;
    SIGNAL S1741 : STD_LOGIC;
    SIGNAL S1742 : STD_LOGIC;
    SIGNAL S1743 : STD_LOGIC;
    SIGNAL S1744 : STD_LOGIC;
    SIGNAL S1745 : STD_LOGIC;
    SIGNAL S1746 : STD_LOGIC;
    SIGNAL S1747 : STD_LOGIC;
    SIGNAL S1748 : STD_LOGIC;
    SIGNAL S1749 : STD_LOGIC;
    SIGNAL S1750 : STD_LOGIC;
    SIGNAL S1751 : STD_LOGIC;
    SIGNAL S1752 : STD_LOGIC;
    SIGNAL S1753 : STD_LOGIC;
    SIGNAL S1754 : STD_LOGIC;
    SIGNAL S1755 : STD_LOGIC;
    SIGNAL S1756 : STD_LOGIC;
    SIGNAL S1757 : STD_LOGIC;
    SIGNAL S1758 : STD_LOGIC;
    SIGNAL S1759 : STD_LOGIC;
    SIGNAL S1760 : STD_LOGIC;
    SIGNAL S1761 : STD_LOGIC;
    SIGNAL S1762 : STD_LOGIC;
    SIGNAL S1763 : STD_LOGIC;
    SIGNAL S1764 : STD_LOGIC;
    SIGNAL S1765 : STD_LOGIC;
    SIGNAL S1766 : STD_LOGIC;
    SIGNAL S1767 : STD_LOGIC;
    SIGNAL S1768 : STD_LOGIC;
    SIGNAL S1769 : STD_LOGIC;
    SIGNAL S1770 : STD_LOGIC;
    SIGNAL S1771 : STD_LOGIC;
    SIGNAL S1772 : STD_LOGIC;
    SIGNAL S1773 : STD_LOGIC;
    SIGNAL S1774 : STD_LOGIC;
    SIGNAL S1775 : STD_LOGIC;
    SIGNAL S1776 : STD_LOGIC;
    SIGNAL S1777 : STD_LOGIC;
    SIGNAL S1778 : STD_LOGIC;
    SIGNAL S1779 : STD_LOGIC;
    SIGNAL S1780 : STD_LOGIC;
    SIGNAL S1781 : STD_LOGIC;
    SIGNAL S1782 : STD_LOGIC;
    SIGNAL S1783 : STD_LOGIC;
    SIGNAL S1784 : STD_LOGIC;
    SIGNAL S1785 : STD_LOGIC;
    SIGNAL S1786 : STD_LOGIC;
    SIGNAL S1787 : STD_LOGIC;
    SIGNAL S1788 : STD_LOGIC;
    SIGNAL S1789 : STD_LOGIC;
    SIGNAL S1790 : STD_LOGIC;
    SIGNAL S1791 : STD_LOGIC;
    SIGNAL S1792 : STD_LOGIC;
    SIGNAL S1793 : STD_LOGIC;
    SIGNAL S1794 : STD_LOGIC;
    SIGNAL S1795 : STD_LOGIC;
    SIGNAL S1796 : STD_LOGIC;
    SIGNAL S1797 : STD_LOGIC;
    SIGNAL S1798 : STD_LOGIC;
    SIGNAL S1799 : STD_LOGIC;
    SIGNAL S1800 : STD_LOGIC;
    SIGNAL S1801 : STD_LOGIC;
    SIGNAL S1802 : STD_LOGIC;
    SIGNAL S1803 : STD_LOGIC;
    SIGNAL S1804 : STD_LOGIC;
    SIGNAL S1805 : STD_LOGIC;
    SIGNAL S1806 : STD_LOGIC;
    SIGNAL S1807 : STD_LOGIC;
    SIGNAL S1808 : STD_LOGIC;
    SIGNAL S1809 : STD_LOGIC;
    SIGNAL S1810 : STD_LOGIC;
    SIGNAL S1811 : STD_LOGIC;
    SIGNAL S1812 : STD_LOGIC;
    SIGNAL S1813 : STD_LOGIC;
    SIGNAL S1814 : STD_LOGIC;
    SIGNAL S1815 : STD_LOGIC;
    SIGNAL S1816 : STD_LOGIC;
    SIGNAL S1817 : STD_LOGIC;
    SIGNAL S1818 : STD_LOGIC;
    SIGNAL S1819 : STD_LOGIC;
    SIGNAL S1820 : STD_LOGIC;
    SIGNAL S1821 : STD_LOGIC;
    SIGNAL S1822 : STD_LOGIC;
    SIGNAL S1823 : STD_LOGIC;
    SIGNAL S1824 : STD_LOGIC;
    SIGNAL S1825 : STD_LOGIC;
    SIGNAL S1826 : STD_LOGIC;
    SIGNAL S1827 : STD_LOGIC;
    SIGNAL S1828 : STD_LOGIC;
    SIGNAL S1829 : STD_LOGIC;
    SIGNAL S1830 : STD_LOGIC;
    SIGNAL S1831 : STD_LOGIC;
    SIGNAL S1832 : STD_LOGIC;
    SIGNAL S1833 : STD_LOGIC;
    SIGNAL S1834 : STD_LOGIC;
    SIGNAL S1835 : STD_LOGIC;
    SIGNAL S1836 : STD_LOGIC;
    SIGNAL S1837 : STD_LOGIC;
    SIGNAL S1838 : STD_LOGIC;
    SIGNAL S1839 : STD_LOGIC;
    SIGNAL S1840 : STD_LOGIC;
    SIGNAL S1841 : STD_LOGIC;
    SIGNAL S1842 : STD_LOGIC;
    SIGNAL S1843 : STD_LOGIC;
    SIGNAL S1844 : STD_LOGIC;
    SIGNAL S1845 : STD_LOGIC;
    SIGNAL S1846 : STD_LOGIC;
    SIGNAL S1847 : STD_LOGIC;
    SIGNAL S1848 : STD_LOGIC;
    SIGNAL S1849 : STD_LOGIC;
    SIGNAL S1850 : STD_LOGIC;
    SIGNAL S1851 : STD_LOGIC;
    SIGNAL S1852 : STD_LOGIC;
    SIGNAL S1853 : STD_LOGIC;
    SIGNAL S1854 : STD_LOGIC;
    SIGNAL S1855 : STD_LOGIC;
    SIGNAL S1856 : STD_LOGIC;
    SIGNAL S1857 : STD_LOGIC;
    SIGNAL S1858 : STD_LOGIC;
    SIGNAL S1859 : STD_LOGIC;
    SIGNAL S1860 : STD_LOGIC;
    SIGNAL S1861 : STD_LOGIC;
    SIGNAL S1862 : STD_LOGIC;
    SIGNAL S1863 : STD_LOGIC;
    SIGNAL S1864 : STD_LOGIC;
    SIGNAL S1865 : STD_LOGIC;
    SIGNAL S1866 : STD_LOGIC;
    SIGNAL S1867 : STD_LOGIC;
    SIGNAL S1868 : STD_LOGIC;
    SIGNAL S1869 : STD_LOGIC;
    SIGNAL S1870 : STD_LOGIC;
    SIGNAL S1871 : STD_LOGIC;
    SIGNAL S1872 : STD_LOGIC;
    SIGNAL S1873 : STD_LOGIC;
    SIGNAL S1874 : STD_LOGIC;
    SIGNAL S1875 : STD_LOGIC;
    SIGNAL S1876 : STD_LOGIC;
    SIGNAL S1877 : STD_LOGIC;
    SIGNAL S1878 : STD_LOGIC;
    SIGNAL S1879 : STD_LOGIC;
    SIGNAL S1880 : STD_LOGIC;
    SIGNAL S1881 : STD_LOGIC;
    SIGNAL S1882 : STD_LOGIC;
    SIGNAL S1883 : STD_LOGIC;
    SIGNAL S1884 : STD_LOGIC;
    SIGNAL S1885 : STD_LOGIC;
    SIGNAL S1886 : STD_LOGIC;
    SIGNAL S1887 : STD_LOGIC;
    SIGNAL S1888 : STD_LOGIC;
    SIGNAL S1889 : STD_LOGIC;
    SIGNAL S1890 : STD_LOGIC;
    SIGNAL S1891 : STD_LOGIC;
    SIGNAL S1892 : STD_LOGIC;
    SIGNAL S1893 : STD_LOGIC;
    SIGNAL S1894 : STD_LOGIC;
    SIGNAL S1895 : STD_LOGIC;
    SIGNAL S1896 : STD_LOGIC;
    SIGNAL S1897 : STD_LOGIC;
    SIGNAL S1898 : STD_LOGIC;
    SIGNAL S1899 : STD_LOGIC;
    SIGNAL S1900 : STD_LOGIC;
    SIGNAL S1901 : STD_LOGIC;
    SIGNAL S1902 : STD_LOGIC;
    SIGNAL S1903 : STD_LOGIC;
    SIGNAL S1904 : STD_LOGIC;
    SIGNAL S1905 : STD_LOGIC;
    SIGNAL S1906 : STD_LOGIC;
    SIGNAL S1907 : STD_LOGIC;
    SIGNAL S1908 : STD_LOGIC;
    SIGNAL S1909 : STD_LOGIC;
    SIGNAL S1910 : STD_LOGIC;
    SIGNAL S1911 : STD_LOGIC;
    SIGNAL S1912 : STD_LOGIC;
    SIGNAL S1913 : STD_LOGIC;
    SIGNAL S1914 : STD_LOGIC;
    SIGNAL S1915 : STD_LOGIC;
    SIGNAL S1916 : STD_LOGIC;
    SIGNAL S1917 : STD_LOGIC;
    SIGNAL S1918 : STD_LOGIC;
    SIGNAL S1919 : STD_LOGIC;
    SIGNAL S1920 : STD_LOGIC;
    SIGNAL S1921 : STD_LOGIC;
    SIGNAL S1922 : STD_LOGIC;
    SIGNAL S1923 : STD_LOGIC;
    SIGNAL S1924 : STD_LOGIC;
    SIGNAL S1925 : STD_LOGIC;
    SIGNAL S1926 : STD_LOGIC;
    SIGNAL S1927 : STD_LOGIC;
    SIGNAL S1928 : STD_LOGIC;
    SIGNAL S1929 : STD_LOGIC;
    SIGNAL S1930 : STD_LOGIC;
    SIGNAL S1931 : STD_LOGIC;
    SIGNAL S1932 : STD_LOGIC;
    SIGNAL S1933 : STD_LOGIC;
    SIGNAL S1934 : STD_LOGIC;
    SIGNAL S1935 : STD_LOGIC;
    SIGNAL S1936 : STD_LOGIC;
    SIGNAL S1937 : STD_LOGIC;
    SIGNAL S1938 : STD_LOGIC;
    SIGNAL S1939 : STD_LOGIC;
    SIGNAL S1940 : STD_LOGIC;
    SIGNAL S1941 : STD_LOGIC;
    SIGNAL S1942 : STD_LOGIC;
    SIGNAL S1943 : STD_LOGIC;
    SIGNAL S1944 : STD_LOGIC;
    SIGNAL S1945 : STD_LOGIC;
    SIGNAL S1946 : STD_LOGIC;
    SIGNAL S1947 : STD_LOGIC;
    SIGNAL S1948 : STD_LOGIC;
    SIGNAL S1949 : STD_LOGIC;
    SIGNAL S1950 : STD_LOGIC;
    SIGNAL S1951 : STD_LOGIC;
    SIGNAL S1952 : STD_LOGIC;
    SIGNAL S1953 : STD_LOGIC;
    SIGNAL S1954 : STD_LOGIC;
    SIGNAL S1955 : STD_LOGIC;
    SIGNAL S1956 : STD_LOGIC;
    SIGNAL S1957 : STD_LOGIC;
    SIGNAL S1958 : STD_LOGIC;
    SIGNAL S1959 : STD_LOGIC;
    SIGNAL S1960 : STD_LOGIC;
    SIGNAL S1961 : STD_LOGIC;
    SIGNAL S1962 : STD_LOGIC;
    SIGNAL S1963 : STD_LOGIC;
    SIGNAL S1964 : STD_LOGIC;
    SIGNAL S1965 : STD_LOGIC;
    SIGNAL S1966 : STD_LOGIC;
    SIGNAL S1967 : STD_LOGIC;
    SIGNAL S1968 : STD_LOGIC;
    SIGNAL S1969 : STD_LOGIC;
    SIGNAL S1970 : STD_LOGIC;
    SIGNAL S1971 : STD_LOGIC;
    SIGNAL S1972 : STD_LOGIC;
    SIGNAL S1973 : STD_LOGIC;
    SIGNAL S1974 : STD_LOGIC;
    SIGNAL S1975 : STD_LOGIC;
    SIGNAL S1976 : STD_LOGIC;
    SIGNAL S1977 : STD_LOGIC;
    SIGNAL S1978 : STD_LOGIC;
    SIGNAL S1979 : STD_LOGIC;
    SIGNAL S1980 : STD_LOGIC;
    SIGNAL S1981 : STD_LOGIC;
    SIGNAL S1982 : STD_LOGIC;
    SIGNAL S1983 : STD_LOGIC;
    SIGNAL S1984 : STD_LOGIC;
    SIGNAL S1985 : STD_LOGIC;
    SIGNAL S1986 : STD_LOGIC;
    SIGNAL S1987 : STD_LOGIC;
    SIGNAL S1988 : STD_LOGIC;
    SIGNAL S1989 : STD_LOGIC;
    SIGNAL S1990 : STD_LOGIC;
    SIGNAL S1991 : STD_LOGIC;
    SIGNAL S1992 : STD_LOGIC;
    SIGNAL S1993 : STD_LOGIC;
    SIGNAL S1994 : STD_LOGIC;
    SIGNAL S1995 : STD_LOGIC;
    SIGNAL S1996 : STD_LOGIC;
    SIGNAL S1997 : STD_LOGIC;
    SIGNAL S1998 : STD_LOGIC;
    SIGNAL S1999 : STD_LOGIC;
    SIGNAL S2000 : STD_LOGIC;
    SIGNAL S2001 : STD_LOGIC;
    SIGNAL S2002 : STD_LOGIC;
    SIGNAL S2003 : STD_LOGIC;
    SIGNAL S2004 : STD_LOGIC;
    SIGNAL S2005 : STD_LOGIC;
    SIGNAL S2006 : STD_LOGIC;
    SIGNAL S2007 : STD_LOGIC;
    SIGNAL S2008 : STD_LOGIC;
    SIGNAL S2009 : STD_LOGIC;
    SIGNAL S2010 : STD_LOGIC;
    SIGNAL S2011 : STD_LOGIC;
    SIGNAL S2012 : STD_LOGIC;
    SIGNAL S2013 : STD_LOGIC;
    SIGNAL S2014 : STD_LOGIC;
    SIGNAL S2015 : STD_LOGIC;
    SIGNAL S2016 : STD_LOGIC;
    SIGNAL S2017 : STD_LOGIC;
    SIGNAL S2018 : STD_LOGIC;
    SIGNAL S2019 : STD_LOGIC;
    SIGNAL S2020 : STD_LOGIC;
    SIGNAL S2021 : STD_LOGIC;
    SIGNAL S2022 : STD_LOGIC;
    SIGNAL S2023 : STD_LOGIC;
    SIGNAL S2024 : STD_LOGIC;
    SIGNAL S2025 : STD_LOGIC;
    SIGNAL S2026 : STD_LOGIC;
    SIGNAL S2027 : STD_LOGIC;
    SIGNAL S2028 : STD_LOGIC;
    SIGNAL S2029 : STD_LOGIC;
    SIGNAL S2030 : STD_LOGIC;
    SIGNAL S2031 : STD_LOGIC;
    SIGNAL S2032 : STD_LOGIC;
    SIGNAL S2033 : STD_LOGIC;
    SIGNAL S2034 : STD_LOGIC;
    SIGNAL S2035 : STD_LOGIC;
    SIGNAL S2036 : STD_LOGIC;
    SIGNAL S2037 : STD_LOGIC;
    SIGNAL S2038 : STD_LOGIC;
    SIGNAL S2039 : STD_LOGIC;
    SIGNAL S2040 : STD_LOGIC;
    SIGNAL S2041 : STD_LOGIC;
    SIGNAL S2042 : STD_LOGIC;
    SIGNAL S2043 : STD_LOGIC;
    SIGNAL S2044 : STD_LOGIC;
    SIGNAL S2045 : STD_LOGIC;
    SIGNAL S2046 : STD_LOGIC;
    SIGNAL S2047 : STD_LOGIC;
    SIGNAL S2048 : STD_LOGIC;
    SIGNAL S2049 : STD_LOGIC;
    SIGNAL S2050 : STD_LOGIC;
    SIGNAL S2051 : STD_LOGIC;
    SIGNAL S2052 : STD_LOGIC;
    SIGNAL S2053 : STD_LOGIC;
    SIGNAL S2054 : STD_LOGIC;
    SIGNAL S2055 : STD_LOGIC;
    SIGNAL S2056 : STD_LOGIC;
    SIGNAL S2057 : STD_LOGIC;
    SIGNAL S2058 : STD_LOGIC;
    SIGNAL S2059 : STD_LOGIC;
    SIGNAL S2060 : STD_LOGIC;
    SIGNAL S2061 : STD_LOGIC;
    SIGNAL S2062 : STD_LOGIC;
    SIGNAL S2063 : STD_LOGIC;
    SIGNAL S2064 : STD_LOGIC;
    SIGNAL S2065 : STD_LOGIC;
    SIGNAL S2066 : STD_LOGIC;
    SIGNAL S2067 : STD_LOGIC;
    SIGNAL S2068 : STD_LOGIC;
    SIGNAL S2069 : STD_LOGIC;
    SIGNAL S2070 : STD_LOGIC;
    SIGNAL S2071 : STD_LOGIC;
    SIGNAL S2072 : STD_LOGIC;
    SIGNAL S2073 : STD_LOGIC;
    SIGNAL S2074 : STD_LOGIC;
    SIGNAL S2075 : STD_LOGIC;
    SIGNAL S2076 : STD_LOGIC;
    SIGNAL S2077 : STD_LOGIC;
    SIGNAL S2078 : STD_LOGIC;
    SIGNAL S2079 : STD_LOGIC;
    SIGNAL S2080 : STD_LOGIC;
    SIGNAL S2081 : STD_LOGIC;
    SIGNAL S2082 : STD_LOGIC;
    SIGNAL S2083 : STD_LOGIC;
    SIGNAL S2084 : STD_LOGIC;
    SIGNAL S2085 : STD_LOGIC;
    SIGNAL S2086 : STD_LOGIC;
    SIGNAL S2087 : STD_LOGIC;
    SIGNAL S2088 : STD_LOGIC;
    SIGNAL S2089 : STD_LOGIC;
    SIGNAL S2090 : STD_LOGIC;
    SIGNAL S2091 : STD_LOGIC;
    SIGNAL S2092 : STD_LOGIC;
    SIGNAL S2093 : STD_LOGIC;
    SIGNAL S2094 : STD_LOGIC;
    SIGNAL S2095 : STD_LOGIC;
    SIGNAL S2096 : STD_LOGIC;
    SIGNAL S2097 : STD_LOGIC;
    SIGNAL S2098 : STD_LOGIC;
    SIGNAL S2099 : STD_LOGIC;
    SIGNAL S2100 : STD_LOGIC;
    SIGNAL S2101 : STD_LOGIC;
    SIGNAL S2102 : STD_LOGIC;
    SIGNAL S2103 : STD_LOGIC;
    SIGNAL S2104 : STD_LOGIC;
    SIGNAL S2105 : STD_LOGIC;
    SIGNAL S2106 : STD_LOGIC;
    SIGNAL S2107 : STD_LOGIC;
    SIGNAL S2108 : STD_LOGIC;
    SIGNAL S2109 : STD_LOGIC;
    SIGNAL S2110 : STD_LOGIC;
    SIGNAL S2111 : STD_LOGIC;
    SIGNAL S2112 : STD_LOGIC;
    SIGNAL S2113 : STD_LOGIC;
    SIGNAL S2114 : STD_LOGIC;
    SIGNAL S2115 : STD_LOGIC;
    SIGNAL S2116 : STD_LOGIC;
    SIGNAL S2117 : STD_LOGIC;
    SIGNAL S2118 : STD_LOGIC;
    SIGNAL S2119 : STD_LOGIC;
    SIGNAL S2120 : STD_LOGIC;
    SIGNAL S2121 : STD_LOGIC;
    SIGNAL S2122 : STD_LOGIC;
    SIGNAL S2123 : STD_LOGIC;
    SIGNAL S2124 : STD_LOGIC;
    SIGNAL S2125 : STD_LOGIC;
    SIGNAL S2126 : STD_LOGIC;
    SIGNAL S2127 : STD_LOGIC;
    SIGNAL S2128 : STD_LOGIC;
    SIGNAL S2129 : STD_LOGIC;
    SIGNAL S2130 : STD_LOGIC;
    SIGNAL S2131 : STD_LOGIC;
    SIGNAL S2132 : STD_LOGIC;
    SIGNAL S2133 : STD_LOGIC;
    SIGNAL S2134 : STD_LOGIC;
    SIGNAL S2135 : STD_LOGIC;
    SIGNAL S2136 : STD_LOGIC;
    SIGNAL S2137 : STD_LOGIC;
    SIGNAL S2138 : STD_LOGIC;
    SIGNAL S2139 : STD_LOGIC;
    SIGNAL S2140 : STD_LOGIC;
    SIGNAL S2141 : STD_LOGIC;
    SIGNAL S2142 : STD_LOGIC;
    SIGNAL S2143 : STD_LOGIC;
    SIGNAL S2144 : STD_LOGIC;
    SIGNAL S2145 : STD_LOGIC;
    SIGNAL S2146 : STD_LOGIC;
    SIGNAL S2147 : STD_LOGIC;
    SIGNAL S2148 : STD_LOGIC;
    SIGNAL S2149 : STD_LOGIC;
    SIGNAL S2150 : STD_LOGIC;
    SIGNAL S2151 : STD_LOGIC;
    SIGNAL S2152 : STD_LOGIC;
    SIGNAL S2153 : STD_LOGIC;
    SIGNAL S2154 : STD_LOGIC;
    SIGNAL S2155 : STD_LOGIC;
    SIGNAL S2156 : STD_LOGIC;
    SIGNAL S2157 : STD_LOGIC;
    SIGNAL S2158 : STD_LOGIC;
    SIGNAL S2159 : STD_LOGIC;
    SIGNAL S2160 : STD_LOGIC;
    SIGNAL S2161 : STD_LOGIC;
    SIGNAL S2162 : STD_LOGIC;
    SIGNAL S2163 : STD_LOGIC;
    SIGNAL S2164 : STD_LOGIC;
    SIGNAL S2165 : STD_LOGIC;
    SIGNAL S2166 : STD_LOGIC;
    SIGNAL S2167 : STD_LOGIC;
    SIGNAL S2168 : STD_LOGIC;
    SIGNAL S2169 : STD_LOGIC;
    SIGNAL S2170 : STD_LOGIC;
    SIGNAL S2171 : STD_LOGIC;
    SIGNAL S2172 : STD_LOGIC;
    SIGNAL S2173 : STD_LOGIC;
    SIGNAL S2174 : STD_LOGIC;
    SIGNAL S2175 : STD_LOGIC;
    SIGNAL S2176 : STD_LOGIC;
    SIGNAL S2177 : STD_LOGIC;
    SIGNAL S2178 : STD_LOGIC;
    SIGNAL S2179 : STD_LOGIC;
    SIGNAL S2180 : STD_LOGIC;
    SIGNAL S2181 : STD_LOGIC;
    SIGNAL S2182 : STD_LOGIC;
    SIGNAL S2183 : STD_LOGIC;
    SIGNAL S2184 : STD_LOGIC;
    SIGNAL S2185 : STD_LOGIC;
    SIGNAL S2186 : STD_LOGIC;
    SIGNAL S2187 : STD_LOGIC;
    SIGNAL S2188 : STD_LOGIC;
    SIGNAL S2189 : STD_LOGIC;
    SIGNAL S2190 : STD_LOGIC;
    SIGNAL S2191 : STD_LOGIC;
    SIGNAL S2192 : STD_LOGIC;
    SIGNAL S2193 : STD_LOGIC;
    SIGNAL S2194 : STD_LOGIC;
    SIGNAL S2195 : STD_LOGIC;
    SIGNAL S2196 : STD_LOGIC;
    SIGNAL S2197 : STD_LOGIC;
    SIGNAL S2198 : STD_LOGIC;
    SIGNAL S2199 : STD_LOGIC;
    SIGNAL S2200 : STD_LOGIC;
    SIGNAL S2201 : STD_LOGIC;
    SIGNAL S2202 : STD_LOGIC;
    SIGNAL S2203 : STD_LOGIC;
    SIGNAL S2204 : STD_LOGIC;
    SIGNAL S2205 : STD_LOGIC;
    SIGNAL S2206 : STD_LOGIC;
    SIGNAL S2207 : STD_LOGIC;
    SIGNAL S2208 : STD_LOGIC;
    SIGNAL S2209 : STD_LOGIC;
    SIGNAL S2210 : STD_LOGIC;
    SIGNAL S2211 : STD_LOGIC;
    SIGNAL S2212 : STD_LOGIC;
    SIGNAL S2213 : STD_LOGIC;
    SIGNAL S2214 : STD_LOGIC;
    SIGNAL S2215 : STD_LOGIC;
    SIGNAL S2216 : STD_LOGIC;
    SIGNAL S2217 : STD_LOGIC;
    SIGNAL S2218 : STD_LOGIC;
    SIGNAL S2219 : STD_LOGIC;
    SIGNAL S2220 : STD_LOGIC;
    SIGNAL S2221 : STD_LOGIC;
    SIGNAL S2222 : STD_LOGIC;
    SIGNAL S2223 : STD_LOGIC;
    SIGNAL S2224 : STD_LOGIC;
    SIGNAL S2225 : STD_LOGIC;
    SIGNAL S2226 : STD_LOGIC;
    SIGNAL S2227 : STD_LOGIC;
    SIGNAL S2228 : STD_LOGIC;
    SIGNAL S2229 : STD_LOGIC;
    SIGNAL S2230 : STD_LOGIC;
    SIGNAL S2231 : STD_LOGIC;
    SIGNAL S2232 : STD_LOGIC;
    SIGNAL S2233 : STD_LOGIC;
    SIGNAL S2234 : STD_LOGIC;
    SIGNAL S2235 : STD_LOGIC;
    SIGNAL S2236 : STD_LOGIC;
    SIGNAL S2237 : STD_LOGIC;
    SIGNAL S2238 : STD_LOGIC;
    SIGNAL S2239 : STD_LOGIC;
    SIGNAL S2240 : STD_LOGIC;
    SIGNAL S2241 : STD_LOGIC;
    SIGNAL S2242 : STD_LOGIC;
    SIGNAL S2243 : STD_LOGIC;
    SIGNAL S2244 : STD_LOGIC;
    SIGNAL S2245 : STD_LOGIC;
    SIGNAL S2246 : STD_LOGIC;
    SIGNAL S2247 : STD_LOGIC;
    SIGNAL S2248 : STD_LOGIC;
    SIGNAL S2249 : STD_LOGIC;
    SIGNAL S2250 : STD_LOGIC;
    SIGNAL S2251 : STD_LOGIC;
    SIGNAL S2252 : STD_LOGIC;
    SIGNAL S2253 : STD_LOGIC;
    SIGNAL S2254 : STD_LOGIC;
    SIGNAL S2255 : STD_LOGIC;
    SIGNAL S2256 : STD_LOGIC;
    SIGNAL S2257 : STD_LOGIC;
    SIGNAL S2258 : STD_LOGIC;
    SIGNAL S2259 : STD_LOGIC;
    SIGNAL S2260 : STD_LOGIC;
    SIGNAL S2261 : STD_LOGIC;
    SIGNAL S2262 : STD_LOGIC;
    SIGNAL S2263 : STD_LOGIC;
    SIGNAL S2264 : STD_LOGIC;
    SIGNAL S2265 : STD_LOGIC;
    SIGNAL S2266 : STD_LOGIC;
    SIGNAL S2267 : STD_LOGIC;
    SIGNAL S2268 : STD_LOGIC;
    SIGNAL S2269 : STD_LOGIC;
    SIGNAL S2270 : STD_LOGIC;
    SIGNAL S2271 : STD_LOGIC;
    SIGNAL S2272 : STD_LOGIC;
    SIGNAL S2273 : STD_LOGIC;
    SIGNAL S2274 : STD_LOGIC;
    SIGNAL S2275 : STD_LOGIC;
    SIGNAL S2276 : STD_LOGIC;
    SIGNAL S2277 : STD_LOGIC;
    SIGNAL S2278 : STD_LOGIC;
    SIGNAL S2279 : STD_LOGIC;
    SIGNAL S2280 : STD_LOGIC;
    SIGNAL S2281 : STD_LOGIC;
    SIGNAL S2282 : STD_LOGIC;
    SIGNAL S2283 : STD_LOGIC;
    SIGNAL S2284 : STD_LOGIC;
    SIGNAL S2285 : STD_LOGIC;
    SIGNAL S2286 : STD_LOGIC;
    SIGNAL S2287 : STD_LOGIC;
    SIGNAL S2288 : STD_LOGIC;
    SIGNAL S2289 : STD_LOGIC;
    SIGNAL S2290 : STD_LOGIC;
    SIGNAL S2291 : STD_LOGIC;
    SIGNAL S2292 : STD_LOGIC;
    SIGNAL S2293 : STD_LOGIC;
    SIGNAL S2294 : STD_LOGIC;
    SIGNAL S2295 : STD_LOGIC;
    SIGNAL S2296 : STD_LOGIC;
    SIGNAL S2297 : STD_LOGIC;
    SIGNAL S2298 : STD_LOGIC;
    SIGNAL S2299 : STD_LOGIC;
    SIGNAL S2300 : STD_LOGIC;
    SIGNAL S2301 : STD_LOGIC;
    SIGNAL S2302 : STD_LOGIC;
    SIGNAL S2303 : STD_LOGIC;
    SIGNAL S2304 : STD_LOGIC;
    SIGNAL S2305 : STD_LOGIC;
    SIGNAL S2306 : STD_LOGIC;
    SIGNAL S2307 : STD_LOGIC;
    SIGNAL S2308 : STD_LOGIC;
    SIGNAL S2309 : STD_LOGIC;
    SIGNAL S2310 : STD_LOGIC;
    SIGNAL S2311 : STD_LOGIC;
    SIGNAL S2312 : STD_LOGIC;
    SIGNAL S2313 : STD_LOGIC;
    SIGNAL S2314 : STD_LOGIC;
    SIGNAL S2315 : STD_LOGIC;
    SIGNAL S2316 : STD_LOGIC;
    SIGNAL S2317 : STD_LOGIC;
    SIGNAL S2318 : STD_LOGIC;
    SIGNAL S2319 : STD_LOGIC;
    SIGNAL S2320 : STD_LOGIC;
    SIGNAL S2321 : STD_LOGIC;
    SIGNAL S2322 : STD_LOGIC;
    SIGNAL S2323 : STD_LOGIC;
    SIGNAL S2324 : STD_LOGIC;
    SIGNAL S2325 : STD_LOGIC;
    SIGNAL S2326 : STD_LOGIC;
    SIGNAL S2327 : STD_LOGIC;
    SIGNAL S2328 : STD_LOGIC;
    SIGNAL S2329 : STD_LOGIC;
    SIGNAL S2330 : STD_LOGIC;
    SIGNAL S2331 : STD_LOGIC;
    SIGNAL S2332 : STD_LOGIC;
    SIGNAL S2333 : STD_LOGIC;
    SIGNAL S2334 : STD_LOGIC;
    SIGNAL S2335 : STD_LOGIC;
    SIGNAL S2336 : STD_LOGIC;
    SIGNAL S2337 : STD_LOGIC;
    SIGNAL S2338 : STD_LOGIC;
    SIGNAL S2339 : STD_LOGIC;
    SIGNAL S2340 : STD_LOGIC;
    SIGNAL S2341 : STD_LOGIC;
    SIGNAL S2342 : STD_LOGIC;
    SIGNAL S2343 : STD_LOGIC;
    SIGNAL S2344 : STD_LOGIC;
    SIGNAL S2345 : STD_LOGIC;
    SIGNAL S2346 : STD_LOGIC;
    SIGNAL S2347 : STD_LOGIC;
    SIGNAL S2348 : STD_LOGIC;
    SIGNAL S2349 : STD_LOGIC;
    SIGNAL S2350 : STD_LOGIC;
    SIGNAL S2351 : STD_LOGIC;
    SIGNAL S2352 : STD_LOGIC;
    SIGNAL S2353 : STD_LOGIC;
    SIGNAL S2354 : STD_LOGIC;
    SIGNAL S2355 : STD_LOGIC;
    SIGNAL S2356 : STD_LOGIC;
    SIGNAL S2357 : STD_LOGIC;
    SIGNAL S2358 : STD_LOGIC;
    SIGNAL S2359 : STD_LOGIC;
    SIGNAL S2360 : STD_LOGIC;
    SIGNAL S2361 : STD_LOGIC;
    SIGNAL S2362 : STD_LOGIC;
    SIGNAL S2363 : STD_LOGIC;
    SIGNAL S2364 : STD_LOGIC;
    SIGNAL S2365 : STD_LOGIC;
    SIGNAL S2366 : STD_LOGIC;
    SIGNAL S2367 : STD_LOGIC;
    SIGNAL S2368 : STD_LOGIC;
    SIGNAL S2369 : STD_LOGIC;
    SIGNAL S2370 : STD_LOGIC;
    SIGNAL S2371 : STD_LOGIC;
    SIGNAL S2372 : STD_LOGIC;
    SIGNAL S2373 : STD_LOGIC;
    SIGNAL S2374 : STD_LOGIC;
    SIGNAL S2375 : STD_LOGIC;
    SIGNAL S2376 : STD_LOGIC;
    SIGNAL S2377 : STD_LOGIC;
    SIGNAL S2378 : STD_LOGIC;
    SIGNAL S2379 : STD_LOGIC;
    SIGNAL S2380 : STD_LOGIC;
    SIGNAL S2381 : STD_LOGIC;
    SIGNAL S2382 : STD_LOGIC;
    SIGNAL S2383 : STD_LOGIC;
    SIGNAL S2384 : STD_LOGIC;
    SIGNAL S2385 : STD_LOGIC;
    SIGNAL S2386 : STD_LOGIC;
    SIGNAL S2387 : STD_LOGIC;
    SIGNAL S2388 : STD_LOGIC;
    SIGNAL S2389 : STD_LOGIC;
    SIGNAL S2390 : STD_LOGIC;
    SIGNAL S2391 : STD_LOGIC;
    SIGNAL S2392 : STD_LOGIC;
    SIGNAL S2393 : STD_LOGIC;
    SIGNAL S2394 : STD_LOGIC;
    SIGNAL S2395 : STD_LOGIC;
    SIGNAL S2396 : STD_LOGIC;
    SIGNAL S2397 : STD_LOGIC;
    SIGNAL S2398 : STD_LOGIC;
    SIGNAL S2399 : STD_LOGIC;
    SIGNAL S2400 : STD_LOGIC;
    SIGNAL S2401 : STD_LOGIC;
    SIGNAL S2402 : STD_LOGIC;
    SIGNAL S2403 : STD_LOGIC;
    SIGNAL S2404 : STD_LOGIC;
    SIGNAL S2405 : STD_LOGIC;
    SIGNAL S2406 : STD_LOGIC;
    SIGNAL S2407 : STD_LOGIC;
    SIGNAL S2408 : STD_LOGIC;
    SIGNAL S2409 : STD_LOGIC;
    SIGNAL S2410 : STD_LOGIC;
    SIGNAL S2411 : STD_LOGIC;
    SIGNAL S2412 : STD_LOGIC;
    SIGNAL S2413 : STD_LOGIC;
    SIGNAL S2414 : STD_LOGIC;
    SIGNAL S2415 : STD_LOGIC;
    SIGNAL S2416 : STD_LOGIC;
    SIGNAL S2417 : STD_LOGIC;
    SIGNAL S2418 : STD_LOGIC;
    SIGNAL S2419 : STD_LOGIC;
    SIGNAL S2420 : STD_LOGIC;
    SIGNAL S2421 : STD_LOGIC;
    SIGNAL S2422 : STD_LOGIC;
    SIGNAL S2423 : STD_LOGIC;
    SIGNAL S2424 : STD_LOGIC;
    SIGNAL S2425 : STD_LOGIC;
    SIGNAL S2426 : STD_LOGIC;
    SIGNAL S2427 : STD_LOGIC;
    SIGNAL S2428 : STD_LOGIC;
    SIGNAL S2429 : STD_LOGIC;
    SIGNAL S2430 : STD_LOGIC;
    SIGNAL S2431 : STD_LOGIC;
    SIGNAL S2432 : STD_LOGIC;
    SIGNAL S2433 : STD_LOGIC;
    SIGNAL S2434 : STD_LOGIC;
    SIGNAL S2435 : STD_LOGIC;
    SIGNAL S2436 : STD_LOGIC;
    SIGNAL S2437 : STD_LOGIC;
    SIGNAL S2438 : STD_LOGIC;
    SIGNAL S2439 : STD_LOGIC;
    SIGNAL S2440 : STD_LOGIC;
    SIGNAL S2441 : STD_LOGIC;
    SIGNAL S2442 : STD_LOGIC;
    SIGNAL S2443 : STD_LOGIC;
    SIGNAL S2444 : STD_LOGIC;
    SIGNAL S2445 : STD_LOGIC;
    SIGNAL S2446 : STD_LOGIC;
    SIGNAL S2447 : STD_LOGIC;
    SIGNAL S2448 : STD_LOGIC;
    SIGNAL S2449 : STD_LOGIC;
    SIGNAL S2450 : STD_LOGIC;
    SIGNAL S2451 : STD_LOGIC;
    SIGNAL S2452 : STD_LOGIC;
    SIGNAL S2453 : STD_LOGIC;
    SIGNAL S2454 : STD_LOGIC;
    SIGNAL S2455 : STD_LOGIC;
    SIGNAL S2456 : STD_LOGIC;
    SIGNAL S2457 : STD_LOGIC;
    SIGNAL S2458 : STD_LOGIC;
    SIGNAL S2459 : STD_LOGIC;
    SIGNAL S2460 : STD_LOGIC;
    SIGNAL S2461 : STD_LOGIC;
    SIGNAL S2462 : STD_LOGIC;
    SIGNAL S2463 : STD_LOGIC;
    SIGNAL S2464 : STD_LOGIC;
    SIGNAL S2465 : STD_LOGIC;
    SIGNAL S2466 : STD_LOGIC;
    SIGNAL S2467 : STD_LOGIC;
    SIGNAL S2468 : STD_LOGIC;
    SIGNAL S2469 : STD_LOGIC;
    SIGNAL S2470 : STD_LOGIC;
    SIGNAL S2471 : STD_LOGIC;
    SIGNAL S2472 : STD_LOGIC;
    SIGNAL S2473 : STD_LOGIC;
    SIGNAL S2474 : STD_LOGIC;
    SIGNAL S2475 : STD_LOGIC;
    SIGNAL S2476 : STD_LOGIC;
    SIGNAL S2477 : STD_LOGIC;
    SIGNAL S2478 : STD_LOGIC;
    SIGNAL S2479 : STD_LOGIC;
    SIGNAL S2480 : STD_LOGIC;
    SIGNAL S2481 : STD_LOGIC;
    SIGNAL S2482 : STD_LOGIC;
    SIGNAL S2483 : STD_LOGIC;
    SIGNAL S2484 : STD_LOGIC;
    SIGNAL S2485 : STD_LOGIC;
    SIGNAL S2486 : STD_LOGIC;
    SIGNAL S2487 : STD_LOGIC;
    SIGNAL S2488 : STD_LOGIC;
    SIGNAL S2489 : STD_LOGIC;
    SIGNAL S2490 : STD_LOGIC;
    SIGNAL S2491 : STD_LOGIC;
    SIGNAL S2492 : STD_LOGIC;
    SIGNAL S2493 : STD_LOGIC;
    SIGNAL S2494 : STD_LOGIC;
    SIGNAL S2495 : STD_LOGIC;
    SIGNAL S2496 : STD_LOGIC;
    SIGNAL S2497 : STD_LOGIC;
    SIGNAL S2498 : STD_LOGIC;
    SIGNAL S2499 : STD_LOGIC;
    SIGNAL S2500 : STD_LOGIC;
    SIGNAL S2501 : STD_LOGIC;
    SIGNAL S2502 : STD_LOGIC;
    SIGNAL S2503 : STD_LOGIC;
    SIGNAL S2504 : STD_LOGIC;
    SIGNAL S2505 : STD_LOGIC;
    SIGNAL S2506 : STD_LOGIC;
    SIGNAL S2507 : STD_LOGIC;
    SIGNAL S2508 : STD_LOGIC;
    SIGNAL S2509 : STD_LOGIC;
    SIGNAL S2510 : STD_LOGIC;
    SIGNAL S2511 : STD_LOGIC;
    SIGNAL S2512 : STD_LOGIC;
    SIGNAL S2513 : STD_LOGIC;
    SIGNAL S2514 : STD_LOGIC;
    SIGNAL S2515 : STD_LOGIC;
    SIGNAL S2516 : STD_LOGIC;
    SIGNAL S2517 : STD_LOGIC;
    SIGNAL S2518 : STD_LOGIC;
    SIGNAL S2519 : STD_LOGIC;
    SIGNAL S2520 : STD_LOGIC;
    SIGNAL S2521 : STD_LOGIC;
    SIGNAL S2522 : STD_LOGIC;
    SIGNAL S2523 : STD_LOGIC;
    SIGNAL S2524 : STD_LOGIC;
    SIGNAL S2525 : STD_LOGIC;
    SIGNAL S2526 : STD_LOGIC;
    SIGNAL S2527 : STD_LOGIC;
    SIGNAL S2528 : STD_LOGIC;
    SIGNAL S2529 : STD_LOGIC;
    SIGNAL S2530 : STD_LOGIC;
    SIGNAL S2531 : STD_LOGIC;
    SIGNAL S2532 : STD_LOGIC;
    SIGNAL S2533 : STD_LOGIC;
    SIGNAL S2534 : STD_LOGIC;
    SIGNAL S2535 : STD_LOGIC;
    SIGNAL S2536 : STD_LOGIC;
    SIGNAL S2537 : STD_LOGIC;
    SIGNAL S2538 : STD_LOGIC;
    SIGNAL S2539 : STD_LOGIC;
    SIGNAL S2540 : STD_LOGIC;
    SIGNAL S2541 : STD_LOGIC;
    SIGNAL S2542 : STD_LOGIC;
    SIGNAL S2543 : STD_LOGIC;
    SIGNAL S2544 : STD_LOGIC;
    SIGNAL S2545 : STD_LOGIC;
    SIGNAL S2546 : STD_LOGIC;
    SIGNAL S2547 : STD_LOGIC;
    SIGNAL S2548 : STD_LOGIC;
    SIGNAL S2549 : STD_LOGIC;
    SIGNAL S2550 : STD_LOGIC;
    SIGNAL S2551 : STD_LOGIC;
    SIGNAL S2552 : STD_LOGIC;
    SIGNAL S2553 : STD_LOGIC;
    SIGNAL S2554 : STD_LOGIC;
    SIGNAL S2555 : STD_LOGIC;
    SIGNAL S2556 : STD_LOGIC;
    SIGNAL S2557 : STD_LOGIC;
    SIGNAL S2558 : STD_LOGIC;
    SIGNAL S2559 : STD_LOGIC;
    SIGNAL S2560 : STD_LOGIC;
    SIGNAL S2561 : STD_LOGIC;
    SIGNAL S2562 : STD_LOGIC;
    SIGNAL S2563 : STD_LOGIC;
    SIGNAL S2564 : STD_LOGIC;
    SIGNAL S2565 : STD_LOGIC;
    SIGNAL S2566 : STD_LOGIC;
    SIGNAL S2567 : STD_LOGIC;
    SIGNAL S2568 : STD_LOGIC;
    SIGNAL S2569 : STD_LOGIC;
    SIGNAL S2570 : STD_LOGIC;
    SIGNAL S2571 : STD_LOGIC;
    SIGNAL S2572 : STD_LOGIC;
    SIGNAL S2573 : STD_LOGIC;
    SIGNAL S2574 : STD_LOGIC;
    SIGNAL S2575 : STD_LOGIC;
    SIGNAL S2576 : STD_LOGIC;
    SIGNAL S2577 : STD_LOGIC;
    SIGNAL S2578 : STD_LOGIC;
    SIGNAL S2579 : STD_LOGIC;
    SIGNAL S2580 : STD_LOGIC;
    SIGNAL S2581 : STD_LOGIC;
    SIGNAL S2582 : STD_LOGIC;
    SIGNAL S2583 : STD_LOGIC;
    SIGNAL S2584 : STD_LOGIC;
    SIGNAL S2585 : STD_LOGIC;
    SIGNAL S2586 : STD_LOGIC;
    SIGNAL S2587 : STD_LOGIC;
    SIGNAL S2588 : STD_LOGIC;
    SIGNAL S2589 : STD_LOGIC;
    SIGNAL S2590 : STD_LOGIC;
    SIGNAL S2591 : STD_LOGIC;
    SIGNAL S2592 : STD_LOGIC;
    SIGNAL S2593 : STD_LOGIC;
    SIGNAL S2594 : STD_LOGIC;
    SIGNAL S2595 : STD_LOGIC;
    SIGNAL S2596 : STD_LOGIC;
    SIGNAL S2597 : STD_LOGIC;
    SIGNAL S2598 : STD_LOGIC;
    SIGNAL S2599 : STD_LOGIC;
    SIGNAL S2600 : STD_LOGIC;
    SIGNAL S2601 : STD_LOGIC;
    SIGNAL S2602 : STD_LOGIC;
    SIGNAL S2603 : STD_LOGIC;
    SIGNAL S2604 : STD_LOGIC;
    SIGNAL S2605 : STD_LOGIC;
    SIGNAL S2606 : STD_LOGIC;
    SIGNAL S2607 : STD_LOGIC;
    SIGNAL S2608 : STD_LOGIC;
    SIGNAL S2609 : STD_LOGIC;
    SIGNAL S2610 : STD_LOGIC;
    SIGNAL S2611 : STD_LOGIC;
    SIGNAL S2612 : STD_LOGIC;
    SIGNAL S2613 : STD_LOGIC;
    SIGNAL S2614 : STD_LOGIC;
    SIGNAL S2615 : STD_LOGIC;
    SIGNAL S2616 : STD_LOGIC;
    SIGNAL S2617 : STD_LOGIC;
    SIGNAL S2618 : STD_LOGIC;
    SIGNAL S2619 : STD_LOGIC;
    SIGNAL S2620 : STD_LOGIC;
    SIGNAL S2621 : STD_LOGIC;
    SIGNAL S2622 : STD_LOGIC;
    SIGNAL S2623 : STD_LOGIC;
    SIGNAL S2624 : STD_LOGIC;
    SIGNAL S2625 : STD_LOGIC;
    SIGNAL S2626 : STD_LOGIC;
    SIGNAL S2627 : STD_LOGIC;
    SIGNAL S2628 : STD_LOGIC;
    SIGNAL S2629 : STD_LOGIC;
    SIGNAL S2630 : STD_LOGIC;
    SIGNAL S2631 : STD_LOGIC;
    SIGNAL S2632 : STD_LOGIC;
    SIGNAL S2633 : STD_LOGIC;
    SIGNAL S2634 : STD_LOGIC;
    SIGNAL S2635 : STD_LOGIC;
    SIGNAL S2636 : STD_LOGIC;
    SIGNAL S2637 : STD_LOGIC;
    SIGNAL S2638 : STD_LOGIC;
    SIGNAL S2639 : STD_LOGIC;
    SIGNAL S2640 : STD_LOGIC;
    SIGNAL S2641 : STD_LOGIC;
    SIGNAL S2642 : STD_LOGIC;
    SIGNAL S2643 : STD_LOGIC;
    SIGNAL S2644 : STD_LOGIC;
    SIGNAL S2645 : STD_LOGIC;
    SIGNAL S2646 : STD_LOGIC;
    SIGNAL S2647 : STD_LOGIC;
    SIGNAL S2648 : STD_LOGIC;
    SIGNAL S2649 : STD_LOGIC;
    SIGNAL S2650 : STD_LOGIC;
    SIGNAL S2651 : STD_LOGIC;
    SIGNAL S2652 : STD_LOGIC;
    SIGNAL S2653 : STD_LOGIC;
    SIGNAL S2654 : STD_LOGIC;
    SIGNAL S2655 : STD_LOGIC;
    SIGNAL S2656 : STD_LOGIC;
    SIGNAL S2657 : STD_LOGIC;
    SIGNAL S2658 : STD_LOGIC;
    SIGNAL S2659 : STD_LOGIC;
    SIGNAL S2660 : STD_LOGIC;
    SIGNAL S2661 : STD_LOGIC;
    SIGNAL S2662 : STD_LOGIC;
    SIGNAL S2663 : STD_LOGIC;
    SIGNAL S2664 : STD_LOGIC;
    SIGNAL S2665 : STD_LOGIC;
    SIGNAL S2666 : STD_LOGIC;
    SIGNAL S2667 : STD_LOGIC;
    SIGNAL S2668 : STD_LOGIC;
    SIGNAL S2669 : STD_LOGIC;
    SIGNAL S2670 : STD_LOGIC;
    SIGNAL S2671 : STD_LOGIC;
    SIGNAL S2672 : STD_LOGIC;
    SIGNAL S2673 : STD_LOGIC;
    SIGNAL S2674 : STD_LOGIC;
    SIGNAL S2675 : STD_LOGIC;
    SIGNAL S2676 : STD_LOGIC;
    SIGNAL S2677 : STD_LOGIC;
    SIGNAL S2678 : STD_LOGIC;
    SIGNAL S2679 : STD_LOGIC;
    SIGNAL S2680 : STD_LOGIC;
    SIGNAL S2681 : STD_LOGIC;
    SIGNAL S2682 : STD_LOGIC;
    SIGNAL S2683 : STD_LOGIC;
    SIGNAL S2684 : STD_LOGIC;
    SIGNAL S2685 : STD_LOGIC;
    SIGNAL S2686 : STD_LOGIC;
    SIGNAL S2687 : STD_LOGIC;
    SIGNAL S2688 : STD_LOGIC;
    SIGNAL S2689 : STD_LOGIC;
    SIGNAL S2690 : STD_LOGIC;
    SIGNAL S2691 : STD_LOGIC;
    SIGNAL S2692 : STD_LOGIC;
    SIGNAL S2693 : STD_LOGIC;
    SIGNAL S2694 : STD_LOGIC;
    SIGNAL S2695 : STD_LOGIC;
    SIGNAL S2696 : STD_LOGIC;
    SIGNAL S2697 : STD_LOGIC;
    SIGNAL S2698 : STD_LOGIC;
    SIGNAL S2699 : STD_LOGIC;
    SIGNAL S2700 : STD_LOGIC;
    SIGNAL S2701 : STD_LOGIC;
    SIGNAL S2702 : STD_LOGIC;
    SIGNAL S2703 : STD_LOGIC;
    SIGNAL S2704 : STD_LOGIC;
    SIGNAL S2705 : STD_LOGIC;
    SIGNAL S2706 : STD_LOGIC;
    SIGNAL S2707 : STD_LOGIC;
    SIGNAL S2708 : STD_LOGIC;
    SIGNAL S2709 : STD_LOGIC;
    SIGNAL S2710 : STD_LOGIC;
    SIGNAL S2711 : STD_LOGIC;
    SIGNAL S2712 : STD_LOGIC;
    SIGNAL S2713 : STD_LOGIC;
    SIGNAL S2714 : STD_LOGIC;
    SIGNAL S2715 : STD_LOGIC;
    SIGNAL S2716 : STD_LOGIC;
    SIGNAL S2717 : STD_LOGIC;
    SIGNAL S2718 : STD_LOGIC;
    SIGNAL S2719 : STD_LOGIC;
    SIGNAL S2720 : STD_LOGIC;
    SIGNAL S2721 : STD_LOGIC;
    SIGNAL S2722 : STD_LOGIC;
    SIGNAL S2723 : STD_LOGIC;
    SIGNAL S2724 : STD_LOGIC;
    SIGNAL S2725 : STD_LOGIC;
    SIGNAL S2726 : STD_LOGIC;
    SIGNAL S2727 : STD_LOGIC;
    SIGNAL S2728 : STD_LOGIC;
    SIGNAL S2729 : STD_LOGIC;
    SIGNAL S2730 : STD_LOGIC;
    SIGNAL S2731 : STD_LOGIC;
    SIGNAL S2732 : STD_LOGIC;
    SIGNAL S2733 : STD_LOGIC;
    SIGNAL S2734 : STD_LOGIC;
    SIGNAL S2735 : STD_LOGIC;
    SIGNAL S2736 : STD_LOGIC;
    SIGNAL S2737 : STD_LOGIC;
    SIGNAL S2738 : STD_LOGIC;
    SIGNAL S2739 : STD_LOGIC;
    SIGNAL S2740 : STD_LOGIC;
    SIGNAL S2741 : STD_LOGIC;
    SIGNAL S2742 : STD_LOGIC;
    SIGNAL S2743 : STD_LOGIC;
    SIGNAL S2744 : STD_LOGIC;
    SIGNAL S2745 : STD_LOGIC;
    SIGNAL S2746 : STD_LOGIC;
    SIGNAL S2747 : STD_LOGIC;
    SIGNAL S2748 : STD_LOGIC;
    SIGNAL S2749 : STD_LOGIC;
    SIGNAL S2750 : STD_LOGIC;
    SIGNAL S2751 : STD_LOGIC;
    SIGNAL S2752 : STD_LOGIC;
    SIGNAL S2753 : STD_LOGIC;
    SIGNAL S2754 : STD_LOGIC;
    SIGNAL S2755 : STD_LOGIC;
    SIGNAL S2756 : STD_LOGIC;
    SIGNAL S2757 : STD_LOGIC;
    SIGNAL S2758 : STD_LOGIC;
    SIGNAL S2759 : STD_LOGIC;
    SIGNAL S2760 : STD_LOGIC;
    SIGNAL S2761 : STD_LOGIC;
    SIGNAL S2762 : STD_LOGIC;
    SIGNAL S2763 : STD_LOGIC;
    SIGNAL S2764 : STD_LOGIC;
    SIGNAL S2765 : STD_LOGIC;
    SIGNAL S2766 : STD_LOGIC;
    SIGNAL S2767 : STD_LOGIC;
    SIGNAL S2768 : STD_LOGIC;
    SIGNAL S2769 : STD_LOGIC;
    SIGNAL S2770 : STD_LOGIC;
    SIGNAL S2771 : STD_LOGIC;
    SIGNAL S2772 : STD_LOGIC;
    SIGNAL S2773 : STD_LOGIC;
    SIGNAL S2774 : STD_LOGIC;
    SIGNAL S2775 : STD_LOGIC;
    SIGNAL S2776 : STD_LOGIC;
    SIGNAL S2777 : STD_LOGIC;
    SIGNAL S2778 : STD_LOGIC;
    SIGNAL S2779 : STD_LOGIC;
    SIGNAL S2780 : STD_LOGIC;
    SIGNAL S2781 : STD_LOGIC;
    SIGNAL S2782 : STD_LOGIC;
    SIGNAL S2783 : STD_LOGIC;
    SIGNAL S2784 : STD_LOGIC;
    SIGNAL S2785 : STD_LOGIC;
    SIGNAL S2786 : STD_LOGIC;
    SIGNAL S2787 : STD_LOGIC;
    SIGNAL S2788 : STD_LOGIC;
    SIGNAL S2789 : STD_LOGIC;
    SIGNAL S2790 : STD_LOGIC;
    SIGNAL S2791 : STD_LOGIC;
    SIGNAL S2792 : STD_LOGIC;
    SIGNAL S2793 : STD_LOGIC;
    SIGNAL S2794 : STD_LOGIC;
    SIGNAL S2795 : STD_LOGIC;
    SIGNAL S2796 : STD_LOGIC;
    SIGNAL S2797 : STD_LOGIC;
    SIGNAL S2798 : STD_LOGIC;
    SIGNAL S2799 : STD_LOGIC;
    SIGNAL S2800 : STD_LOGIC;
    SIGNAL S2801 : STD_LOGIC;
    SIGNAL S2802 : STD_LOGIC;
    SIGNAL S2803 : STD_LOGIC;
    SIGNAL S2804 : STD_LOGIC;
    SIGNAL S2805 : STD_LOGIC;
    SIGNAL S2806 : STD_LOGIC;
    SIGNAL S2807 : STD_LOGIC;
    SIGNAL S2808 : STD_LOGIC;
    SIGNAL S2809 : STD_LOGIC;
    SIGNAL S2810 : STD_LOGIC;
    SIGNAL S2811 : STD_LOGIC;
    SIGNAL S2812 : STD_LOGIC;
    SIGNAL S2813 : STD_LOGIC;
    SIGNAL S2814 : STD_LOGIC;
    SIGNAL S2815 : STD_LOGIC;
    SIGNAL S2816 : STD_LOGIC;
    SIGNAL S2817 : STD_LOGIC;
    SIGNAL S2818 : STD_LOGIC;
    SIGNAL S2819 : STD_LOGIC;
    SIGNAL S2820 : STD_LOGIC;
    SIGNAL S2821 : STD_LOGIC;
    SIGNAL S2822 : STD_LOGIC;
    SIGNAL S2823 : STD_LOGIC;
    SIGNAL S2824 : STD_LOGIC;
    SIGNAL S2825 : STD_LOGIC;
    SIGNAL S2826 : STD_LOGIC;
    SIGNAL S2827 : STD_LOGIC;
    SIGNAL S2828 : STD_LOGIC;
    SIGNAL S2829 : STD_LOGIC;
    SIGNAL S2830 : STD_LOGIC;
    SIGNAL S2831 : STD_LOGIC;
    SIGNAL S2832 : STD_LOGIC;
    SIGNAL S2833 : STD_LOGIC;
    SIGNAL S2834 : STD_LOGIC;
    SIGNAL S2835 : STD_LOGIC;
    SIGNAL S2836 : STD_LOGIC;
    SIGNAL S2837 : STD_LOGIC;
    SIGNAL S2838 : STD_LOGIC;
    SIGNAL S2839 : STD_LOGIC;
    SIGNAL S2840 : STD_LOGIC;
    SIGNAL S2841 : STD_LOGIC;
    SIGNAL S2842 : STD_LOGIC;
    SIGNAL S2843 : STD_LOGIC;
    SIGNAL S2844 : STD_LOGIC;
    SIGNAL S2845 : STD_LOGIC;
    SIGNAL S2846 : STD_LOGIC;
    SIGNAL S2847 : STD_LOGIC;
    SIGNAL S2848 : STD_LOGIC;
    SIGNAL S2849 : STD_LOGIC;
    SIGNAL S2850 : STD_LOGIC;
    SIGNAL S2851 : STD_LOGIC;
    SIGNAL S2852 : STD_LOGIC;
    SIGNAL S2853 : STD_LOGIC;
    SIGNAL S2854 : STD_LOGIC;
    SIGNAL S2855 : STD_LOGIC;
    SIGNAL S2856 : STD_LOGIC;
    SIGNAL S2857 : STD_LOGIC;
    SIGNAL S2858 : STD_LOGIC;
    SIGNAL S2859 : STD_LOGIC;
    SIGNAL S2860 : STD_LOGIC;
    SIGNAL S2861 : STD_LOGIC;
    SIGNAL S2862 : STD_LOGIC;
    SIGNAL S2863 : STD_LOGIC;
    SIGNAL S2864 : STD_LOGIC;
    SIGNAL S2865 : STD_LOGIC;
    SIGNAL S2866 : STD_LOGIC;
    SIGNAL S2867 : STD_LOGIC;
    SIGNAL S2868 : STD_LOGIC;
    SIGNAL S2869 : STD_LOGIC;
    SIGNAL S2870 : STD_LOGIC;
    SIGNAL S2871 : STD_LOGIC;
    SIGNAL S2872 : STD_LOGIC;
    SIGNAL S2873 : STD_LOGIC;
    SIGNAL S2874 : STD_LOGIC;
    SIGNAL S2875 : STD_LOGIC;
    SIGNAL S2876 : STD_LOGIC;
    SIGNAL S2877 : STD_LOGIC;
    SIGNAL S2878 : STD_LOGIC;
    SIGNAL S2879 : STD_LOGIC;
    SIGNAL S2880 : STD_LOGIC;
    SIGNAL S2881 : STD_LOGIC;
    SIGNAL S2882 : STD_LOGIC;
    SIGNAL S2883 : STD_LOGIC;
    SIGNAL S2884 : STD_LOGIC;
    SIGNAL S2885 : STD_LOGIC;
    SIGNAL S2886 : STD_LOGIC;
    SIGNAL S2887 : STD_LOGIC;
    SIGNAL S2888 : STD_LOGIC;
    SIGNAL S2889 : STD_LOGIC;
    SIGNAL S2890 : STD_LOGIC;
    SIGNAL S2891 : STD_LOGIC;
    SIGNAL S2892 : STD_LOGIC;
    SIGNAL S2893 : STD_LOGIC;
    SIGNAL S2894 : STD_LOGIC;
    SIGNAL S2895 : STD_LOGIC;
    SIGNAL S2896 : STD_LOGIC;
    SIGNAL S2897 : STD_LOGIC;
    SIGNAL S2898 : STD_LOGIC;
    SIGNAL S2899 : STD_LOGIC;
    SIGNAL S2900 : STD_LOGIC;
    SIGNAL S2901 : STD_LOGIC;
    SIGNAL S2902 : STD_LOGIC;
    SIGNAL S2903 : STD_LOGIC;
    SIGNAL S2904 : STD_LOGIC;
    SIGNAL S2905 : STD_LOGIC;
    SIGNAL S2906 : STD_LOGIC;
    SIGNAL S2907 : STD_LOGIC;
    SIGNAL S2908 : STD_LOGIC;
    SIGNAL S2909 : STD_LOGIC;
    SIGNAL S2910 : STD_LOGIC;
    SIGNAL S2911 : STD_LOGIC;
    SIGNAL S2912 : STD_LOGIC;
    SIGNAL S2913 : STD_LOGIC;
    SIGNAL S2914 : STD_LOGIC;
    SIGNAL S2915 : STD_LOGIC;
    SIGNAL S2916 : STD_LOGIC;
    SIGNAL S2917 : STD_LOGIC;
    SIGNAL S2918 : STD_LOGIC;
    SIGNAL S2919 : STD_LOGIC;
    SIGNAL S2920 : STD_LOGIC;
    SIGNAL S2921 : STD_LOGIC;
    SIGNAL S2922 : STD_LOGIC;
    SIGNAL S2923 : STD_LOGIC;
    SIGNAL S2924 : STD_LOGIC;
    SIGNAL S2925 : STD_LOGIC;
    SIGNAL S2926 : STD_LOGIC;
    SIGNAL S2927 : STD_LOGIC;
    SIGNAL S2928 : STD_LOGIC;
    SIGNAL S2929 : STD_LOGIC;
    SIGNAL S2930 : STD_LOGIC;
    SIGNAL S2931 : STD_LOGIC;
    SIGNAL S2932 : STD_LOGIC;
    SIGNAL S2933 : STD_LOGIC;
    SIGNAL S2934 : STD_LOGIC;
    SIGNAL S2935 : STD_LOGIC;
    SIGNAL S2936 : STD_LOGIC;
    SIGNAL S2937 : STD_LOGIC;
    SIGNAL S2938 : STD_LOGIC;
    SIGNAL S2939 : STD_LOGIC;
    SIGNAL S2940 : STD_LOGIC;
    SIGNAL S2941 : STD_LOGIC;
    SIGNAL S2942 : STD_LOGIC;
    SIGNAL S2943 : STD_LOGIC;
    SIGNAL S2944 : STD_LOGIC;
    SIGNAL S2945 : STD_LOGIC;
    SIGNAL S2946 : STD_LOGIC;
    SIGNAL S2947 : STD_LOGIC;
    SIGNAL S2948 : STD_LOGIC;
    SIGNAL S2949 : STD_LOGIC;
    SIGNAL S2950 : STD_LOGIC;
    SIGNAL S2951 : STD_LOGIC;
    SIGNAL S2952 : STD_LOGIC;
    SIGNAL S2953 : STD_LOGIC;
    SIGNAL S2954 : STD_LOGIC;
    SIGNAL S2955 : STD_LOGIC;
    SIGNAL S2956 : STD_LOGIC;
    SIGNAL S2957 : STD_LOGIC;
    SIGNAL S2958 : STD_LOGIC;
    SIGNAL S2959 : STD_LOGIC;
    SIGNAL S2960 : STD_LOGIC;
    SIGNAL S2961 : STD_LOGIC;
    SIGNAL S2962 : STD_LOGIC;
    SIGNAL S2963 : STD_LOGIC;
    SIGNAL S2964 : STD_LOGIC;
    SIGNAL S2965 : STD_LOGIC;
    SIGNAL S2966 : STD_LOGIC;
    SIGNAL S2967 : STD_LOGIC;
    SIGNAL S2968 : STD_LOGIC;
    SIGNAL S2969 : STD_LOGIC;
    SIGNAL S2970 : STD_LOGIC;
    SIGNAL S2971 : STD_LOGIC;
    SIGNAL S2972 : STD_LOGIC;
    SIGNAL S2973 : STD_LOGIC;
    SIGNAL S2974 : STD_LOGIC;
    SIGNAL S2975 : STD_LOGIC;
    SIGNAL S2976 : STD_LOGIC;
    SIGNAL S2977 : STD_LOGIC;
    SIGNAL S2978 : STD_LOGIC;
    SIGNAL S2979 : STD_LOGIC;
    SIGNAL S2980 : STD_LOGIC;
    SIGNAL S2981 : STD_LOGIC;
    SIGNAL S2982 : STD_LOGIC;
    SIGNAL S2983 : STD_LOGIC;
    SIGNAL S2984 : STD_LOGIC;
    SIGNAL S2985 : STD_LOGIC;
    SIGNAL S2986 : STD_LOGIC;
    SIGNAL S2987 : STD_LOGIC;
    SIGNAL S2988 : STD_LOGIC;
    SIGNAL S2989 : STD_LOGIC;
    SIGNAL S2990 : STD_LOGIC;
    SIGNAL S2991 : STD_LOGIC;
    SIGNAL S2992 : STD_LOGIC;
    SIGNAL S2993 : STD_LOGIC;
    SIGNAL S2994 : STD_LOGIC;
    SIGNAL S2995 : STD_LOGIC;
    SIGNAL S2996 : STD_LOGIC;
    SIGNAL S2997 : STD_LOGIC;
    SIGNAL S2998 : STD_LOGIC;
    SIGNAL S2999 : STD_LOGIC;
    SIGNAL S3000 : STD_LOGIC;
    SIGNAL S3001 : STD_LOGIC;
    SIGNAL S3002 : STD_LOGIC;
    SIGNAL S3003 : STD_LOGIC;
    SIGNAL S3004 : STD_LOGIC;
    SIGNAL S3005 : STD_LOGIC;
    SIGNAL S3006 : STD_LOGIC;
    SIGNAL S3007 : STD_LOGIC;
    SIGNAL S3008 : STD_LOGIC;
    SIGNAL S3009 : STD_LOGIC;
    SIGNAL S3010 : STD_LOGIC;
    SIGNAL S3011 : STD_LOGIC;
    SIGNAL S3012 : STD_LOGIC;
    SIGNAL S3013 : STD_LOGIC;
    SIGNAL S3014 : STD_LOGIC;
    SIGNAL S3015 : STD_LOGIC;
    SIGNAL S3016 : STD_LOGIC;
    SIGNAL S3017 : STD_LOGIC;
    SIGNAL S3018 : STD_LOGIC;
    SIGNAL S3019 : STD_LOGIC;
    SIGNAL S3020 : STD_LOGIC;
    SIGNAL S3021 : STD_LOGIC;
    SIGNAL S3022 : STD_LOGIC;
    SIGNAL S3023 : STD_LOGIC;
    SIGNAL S3024 : STD_LOGIC;
    SIGNAL S3025 : STD_LOGIC;
    SIGNAL S3026 : STD_LOGIC;
    SIGNAL S3027 : STD_LOGIC;
    SIGNAL S3028 : STD_LOGIC;
    SIGNAL S3029 : STD_LOGIC;
    SIGNAL S3030 : STD_LOGIC;
    SIGNAL S3031 : STD_LOGIC;
    SIGNAL S3032 : STD_LOGIC;
    SIGNAL S3033 : STD_LOGIC;
    SIGNAL S3034 : STD_LOGIC;
    SIGNAL S3035 : STD_LOGIC;
    SIGNAL S3036 : STD_LOGIC;
    SIGNAL S3037 : STD_LOGIC;
    SIGNAL S3038 : STD_LOGIC;
    SIGNAL S3039 : STD_LOGIC;
    SIGNAL S3040 : STD_LOGIC;
    SIGNAL S3041 : STD_LOGIC;
    SIGNAL S3042 : STD_LOGIC;
    SIGNAL S3043 : STD_LOGIC;
    SIGNAL S3044 : STD_LOGIC;
    SIGNAL S3045 : STD_LOGIC;
    SIGNAL S3046 : STD_LOGIC;
    SIGNAL S3047 : STD_LOGIC;
    SIGNAL S3048 : STD_LOGIC;
    SIGNAL S3049 : STD_LOGIC;
    SIGNAL S3050 : STD_LOGIC;
    SIGNAL S3051 : STD_LOGIC;
    SIGNAL S3052 : STD_LOGIC;
    SIGNAL S3053 : STD_LOGIC;
    SIGNAL S3054 : STD_LOGIC;
    SIGNAL S3055 : STD_LOGIC;
    SIGNAL S3056 : STD_LOGIC;
    SIGNAL S3057 : STD_LOGIC;
    SIGNAL S3058 : STD_LOGIC;
    SIGNAL S3059 : STD_LOGIC;
    SIGNAL S3060 : STD_LOGIC;
    SIGNAL S3061 : STD_LOGIC;
    SIGNAL S3062 : STD_LOGIC;
    SIGNAL S3063 : STD_LOGIC;
    SIGNAL S3064 : STD_LOGIC;
    SIGNAL S3065 : STD_LOGIC;
    SIGNAL S3066 : STD_LOGIC;
    SIGNAL S3067 : STD_LOGIC;
    SIGNAL S3068 : STD_LOGIC;
    SIGNAL S3069 : STD_LOGIC;
    SIGNAL S3070 : STD_LOGIC;
    SIGNAL S3071 : STD_LOGIC;
    SIGNAL S3072 : STD_LOGIC;
    SIGNAL S3073 : STD_LOGIC;
    SIGNAL S3074 : STD_LOGIC;
    SIGNAL S3075 : STD_LOGIC;
    SIGNAL S3076 : STD_LOGIC;
    SIGNAL S3077 : STD_LOGIC;
    SIGNAL S3078 : STD_LOGIC;
    SIGNAL S3079 : STD_LOGIC;
    SIGNAL S3080 : STD_LOGIC;
    SIGNAL S3081 : STD_LOGIC;
    SIGNAL S3082 : STD_LOGIC;
    SIGNAL S3083 : STD_LOGIC;
    SIGNAL S3084 : STD_LOGIC;
    SIGNAL S3085 : STD_LOGIC;
    SIGNAL S3086 : STD_LOGIC;
    SIGNAL S3087 : STD_LOGIC;
    SIGNAL S3088 : STD_LOGIC;
    SIGNAL S3089 : STD_LOGIC;
    SIGNAL S3090 : STD_LOGIC;
    SIGNAL S3091 : STD_LOGIC;
    SIGNAL S3092 : STD_LOGIC;
    SIGNAL S3093 : STD_LOGIC;
    SIGNAL S3094 : STD_LOGIC;
    SIGNAL S3095 : STD_LOGIC;
    SIGNAL S3096 : STD_LOGIC;
    SIGNAL S3097 : STD_LOGIC;
    SIGNAL S3098 : STD_LOGIC;
    SIGNAL S3099 : STD_LOGIC;
    SIGNAL S3100 : STD_LOGIC;
    SIGNAL S3101 : STD_LOGIC;
    SIGNAL S3102 : STD_LOGIC;
    SIGNAL S3103 : STD_LOGIC;
    SIGNAL S3104 : STD_LOGIC;
    SIGNAL S3105 : STD_LOGIC;
    SIGNAL S3106 : STD_LOGIC;
    SIGNAL S3107 : STD_LOGIC;
    SIGNAL S3108 : STD_LOGIC;
    SIGNAL S3109 : STD_LOGIC;
    SIGNAL S3110 : STD_LOGIC;
    SIGNAL S3111 : STD_LOGIC;
    SIGNAL S3112 : STD_LOGIC;
    SIGNAL S3113 : STD_LOGIC;
    SIGNAL S3114 : STD_LOGIC;
    SIGNAL S3115 : STD_LOGIC;
    SIGNAL S3116 : STD_LOGIC;
    SIGNAL S3117 : STD_LOGIC;
    SIGNAL S3118 : STD_LOGIC;
    SIGNAL S3119 : STD_LOGIC;
    SIGNAL S3120 : STD_LOGIC;
    SIGNAL S3121 : STD_LOGIC;
    SIGNAL S3122 : STD_LOGIC;
    SIGNAL S3123 : STD_LOGIC;
    SIGNAL S3124 : STD_LOGIC;
    SIGNAL S3125 : STD_LOGIC;
    SIGNAL S3126 : STD_LOGIC;
    SIGNAL S3127 : STD_LOGIC;
    SIGNAL S3128 : STD_LOGIC;
    SIGNAL S3129 : STD_LOGIC;
    SIGNAL S3130 : STD_LOGIC;
    SIGNAL S3131 : STD_LOGIC;
    SIGNAL S3132 : STD_LOGIC;
    SIGNAL S3133 : STD_LOGIC;
    SIGNAL S3134 : STD_LOGIC;
    SIGNAL S3135 : STD_LOGIC;
    SIGNAL S3136 : STD_LOGIC;
    SIGNAL S3137 : STD_LOGIC;
    SIGNAL S3138 : STD_LOGIC;
    SIGNAL S3139 : STD_LOGIC;
    SIGNAL S3140 : STD_LOGIC;
    SIGNAL S3141 : STD_LOGIC;
    SIGNAL S3142 : STD_LOGIC;
    SIGNAL S3143 : STD_LOGIC;
    SIGNAL S3144 : STD_LOGIC;
    SIGNAL S3145 : STD_LOGIC;
    SIGNAL S3146 : STD_LOGIC;
    SIGNAL S3147 : STD_LOGIC;
    SIGNAL S3148 : STD_LOGIC;
    SIGNAL S3149 : STD_LOGIC;
    SIGNAL S3150 : STD_LOGIC;
    SIGNAL S3151 : STD_LOGIC;
    SIGNAL S3152 : STD_LOGIC;
    SIGNAL S3153 : STD_LOGIC;
    SIGNAL S3154 : STD_LOGIC;
    SIGNAL S3155 : STD_LOGIC;
    SIGNAL S3156 : STD_LOGIC;
    SIGNAL S3157 : STD_LOGIC;
    SIGNAL S3158 : STD_LOGIC;
    SIGNAL S3159 : STD_LOGIC;
    SIGNAL S3160 : STD_LOGIC;
    SIGNAL S3161 : STD_LOGIC;
    SIGNAL S3162 : STD_LOGIC;
    SIGNAL S3163 : STD_LOGIC;
    SIGNAL S3164 : STD_LOGIC;
    SIGNAL S3165 : STD_LOGIC;
    SIGNAL S3166 : STD_LOGIC;
    SIGNAL S3167 : STD_LOGIC;
    SIGNAL S3168 : STD_LOGIC;
    SIGNAL S3169 : STD_LOGIC;
    SIGNAL S3170 : STD_LOGIC;
    SIGNAL S3171 : STD_LOGIC;
    SIGNAL S3172 : STD_LOGIC;
    SIGNAL S3173 : STD_LOGIC;
    SIGNAL S3174 : STD_LOGIC;
    SIGNAL S3175 : STD_LOGIC;
    SIGNAL S3176 : STD_LOGIC;
    SIGNAL S3177 : STD_LOGIC;
    SIGNAL S3178 : STD_LOGIC;
    SIGNAL S3179 : STD_LOGIC;
    SIGNAL S3180 : STD_LOGIC;
    SIGNAL S3181 : STD_LOGIC;
    SIGNAL S3182 : STD_LOGIC;
    SIGNAL S3183 : STD_LOGIC;
    SIGNAL S3184 : STD_LOGIC;
    SIGNAL S3185 : STD_LOGIC;
    SIGNAL S3186 : STD_LOGIC;
    SIGNAL S3187 : STD_LOGIC;
    SIGNAL S3188 : STD_LOGIC;
    SIGNAL S3189 : STD_LOGIC;
    SIGNAL S3190 : STD_LOGIC;
    SIGNAL S3191 : STD_LOGIC;
    SIGNAL S3192 : STD_LOGIC;
    SIGNAL S3193 : STD_LOGIC;
    SIGNAL S3194 : STD_LOGIC;
    SIGNAL S3195 : STD_LOGIC;
    SIGNAL S3196 : STD_LOGIC;
    SIGNAL S3197 : STD_LOGIC;
    SIGNAL S3198 : STD_LOGIC;
    SIGNAL S3199 : STD_LOGIC;
    SIGNAL S3200 : STD_LOGIC;
    SIGNAL S3201 : STD_LOGIC;
    SIGNAL S3202 : STD_LOGIC;
    SIGNAL S3203 : STD_LOGIC;
    SIGNAL S3204 : STD_LOGIC;
    SIGNAL S3205 : STD_LOGIC;
    SIGNAL S3206 : STD_LOGIC;
    SIGNAL S3207 : STD_LOGIC;
    SIGNAL S3208 : STD_LOGIC;
    SIGNAL S3209 : STD_LOGIC;
    SIGNAL S3210 : STD_LOGIC;
    SIGNAL S3211 : STD_LOGIC;
    SIGNAL S3212 : STD_LOGIC;
    SIGNAL S3213 : STD_LOGIC;
    SIGNAL S3214 : STD_LOGIC;
    SIGNAL S3215 : STD_LOGIC;
    SIGNAL S3216 : STD_LOGIC;
    SIGNAL S3217 : STD_LOGIC;
    SIGNAL S3218 : STD_LOGIC;
    SIGNAL S3219 : STD_LOGIC;
    SIGNAL S3220 : STD_LOGIC;
    SIGNAL S3221 : STD_LOGIC;
    SIGNAL S3222 : STD_LOGIC;
    SIGNAL S3223 : STD_LOGIC;
    SIGNAL S3224 : STD_LOGIC;
    SIGNAL S3225 : STD_LOGIC;
    SIGNAL S3226 : STD_LOGIC;
    SIGNAL S3227 : STD_LOGIC;
    SIGNAL S3228 : STD_LOGIC;
    SIGNAL S3229 : STD_LOGIC;
    SIGNAL S3230 : STD_LOGIC;
    SIGNAL S3231 : STD_LOGIC;
    SIGNAL S3232 : STD_LOGIC;
    SIGNAL S3233 : STD_LOGIC;
    SIGNAL S3234 : STD_LOGIC;
    SIGNAL S3235 : STD_LOGIC;
    SIGNAL S3236 : STD_LOGIC;
    SIGNAL S3237 : STD_LOGIC;
    SIGNAL S3238 : STD_LOGIC;
    SIGNAL S3239 : STD_LOGIC;
    SIGNAL S3240 : STD_LOGIC;
    SIGNAL S3241 : STD_LOGIC;
    SIGNAL S3242 : STD_LOGIC;
    SIGNAL S3243 : STD_LOGIC;
    SIGNAL S3244 : STD_LOGIC;
    SIGNAL S3245 : STD_LOGIC;
    SIGNAL S3246 : STD_LOGIC;
    SIGNAL S3247 : STD_LOGIC;
    SIGNAL S3248 : STD_LOGIC;
    SIGNAL S3249 : STD_LOGIC;
    SIGNAL S3250 : STD_LOGIC;
    SIGNAL S3251 : STD_LOGIC;
    SIGNAL S3252 : STD_LOGIC;
    SIGNAL S3253 : STD_LOGIC;
    SIGNAL S3254 : STD_LOGIC;
    SIGNAL S3255 : STD_LOGIC;
    SIGNAL S3256 : STD_LOGIC;
    SIGNAL S3257 : STD_LOGIC;
    SIGNAL S3258 : STD_LOGIC;
    SIGNAL S3259 : STD_LOGIC;
    SIGNAL S3260 : STD_LOGIC;
    SIGNAL S3261 : STD_LOGIC;
    SIGNAL S3262 : STD_LOGIC;
    SIGNAL S3263 : STD_LOGIC;
    SIGNAL S3264 : STD_LOGIC;
    SIGNAL S3265 : STD_LOGIC;
    SIGNAL S3266 : STD_LOGIC;
    SIGNAL S3267 : STD_LOGIC;
    SIGNAL S3268 : STD_LOGIC;
    SIGNAL S3269 : STD_LOGIC;
    SIGNAL S3270 : STD_LOGIC;
    SIGNAL S3271 : STD_LOGIC;
    SIGNAL S3272 : STD_LOGIC;
    SIGNAL S3273 : STD_LOGIC;
    SIGNAL S3274 : STD_LOGIC;
    SIGNAL S3275 : STD_LOGIC;
    SIGNAL S3276 : STD_LOGIC;
    SIGNAL S3277 : STD_LOGIC;
    SIGNAL S3278 : STD_LOGIC;
    SIGNAL S3279 : STD_LOGIC;
    SIGNAL S3280 : STD_LOGIC;
    SIGNAL S3281 : STD_LOGIC;
    SIGNAL S3282 : STD_LOGIC;
    SIGNAL S3283 : STD_LOGIC;
    SIGNAL S3284 : STD_LOGIC;
    SIGNAL S3285 : STD_LOGIC;
    SIGNAL S3286 : STD_LOGIC;
    SIGNAL S3287 : STD_LOGIC;
    SIGNAL S3288 : STD_LOGIC;
    SIGNAL S3289 : STD_LOGIC;
    SIGNAL S3290 : STD_LOGIC;
    SIGNAL S3291 : STD_LOGIC;
    SIGNAL S3292 : STD_LOGIC;
    SIGNAL S3293 : STD_LOGIC;
    SIGNAL S3294 : STD_LOGIC;
    SIGNAL S3295 : STD_LOGIC;
    SIGNAL S3296 : STD_LOGIC;
    SIGNAL S3297 : STD_LOGIC;
    SIGNAL S3298 : STD_LOGIC;
    SIGNAL S3299 : STD_LOGIC;
    SIGNAL S3300 : STD_LOGIC;
    SIGNAL S3301 : STD_LOGIC;
    SIGNAL S3302 : STD_LOGIC;
    SIGNAL S3303 : STD_LOGIC;
    SIGNAL S3304 : STD_LOGIC;
    SIGNAL S3305 : STD_LOGIC;
    SIGNAL S3306 : STD_LOGIC;
    SIGNAL S3307 : STD_LOGIC;
    SIGNAL S3308 : STD_LOGIC;
    SIGNAL S3309 : STD_LOGIC;
    SIGNAL S3310 : STD_LOGIC;
    SIGNAL S3311 : STD_LOGIC;
    SIGNAL S3312 : STD_LOGIC;
    SIGNAL S3313 : STD_LOGIC;
    SIGNAL S3314 : STD_LOGIC;
    SIGNAL S3315 : STD_LOGIC;
    SIGNAL S3316 : STD_LOGIC;
    SIGNAL S3317 : STD_LOGIC;
    SIGNAL S3318 : STD_LOGIC;
    SIGNAL S3319 : STD_LOGIC;
    SIGNAL S3320 : STD_LOGIC;
    SIGNAL S3321 : STD_LOGIC;
    SIGNAL S3322 : STD_LOGIC;
    SIGNAL S3323 : STD_LOGIC;
    SIGNAL S3324 : STD_LOGIC;
    SIGNAL S3325 : STD_LOGIC;
    SIGNAL S3326 : STD_LOGIC;
    SIGNAL S3327 : STD_LOGIC;
    SIGNAL S3328 : STD_LOGIC;
    SIGNAL S3329 : STD_LOGIC;
    SIGNAL S3330 : STD_LOGIC;
    SIGNAL S3331 : STD_LOGIC;
    SIGNAL S3332 : STD_LOGIC;
    SIGNAL S3333 : STD_LOGIC;
    SIGNAL S3334 : STD_LOGIC;
    SIGNAL S3335 : STD_LOGIC;
    SIGNAL S3336 : STD_LOGIC;
    SIGNAL S3337 : STD_LOGIC;
    SIGNAL S3338 : STD_LOGIC;
    SIGNAL S3339 : STD_LOGIC;
    SIGNAL S3340 : STD_LOGIC;
    SIGNAL S3341 : STD_LOGIC;
    SIGNAL S3342 : STD_LOGIC;
    SIGNAL S3343 : STD_LOGIC;
    SIGNAL S3344 : STD_LOGIC;
    SIGNAL S3345 : STD_LOGIC;
    SIGNAL S3346 : STD_LOGIC;
    SIGNAL S3347 : STD_LOGIC;
    SIGNAL S3348 : STD_LOGIC;
    SIGNAL S3349 : STD_LOGIC;
    SIGNAL S3350 : STD_LOGIC;
    SIGNAL S3351 : STD_LOGIC;
    SIGNAL S3352 : STD_LOGIC;
    SIGNAL S3353 : STD_LOGIC;
    SIGNAL S3354 : STD_LOGIC;
    SIGNAL S3355 : STD_LOGIC;
    SIGNAL S3356 : STD_LOGIC;
    SIGNAL S3357 : STD_LOGIC;
    SIGNAL S3358 : STD_LOGIC;
    SIGNAL S3359 : STD_LOGIC;
    SIGNAL S3360 : STD_LOGIC;
    SIGNAL S3361 : STD_LOGIC;
    SIGNAL S3362 : STD_LOGIC;
    SIGNAL S3363 : STD_LOGIC;
    SIGNAL S3364 : STD_LOGIC;
    SIGNAL S3365 : STD_LOGIC;
    SIGNAL S3366 : STD_LOGIC;
    SIGNAL S3367 : STD_LOGIC;
    SIGNAL S3368 : STD_LOGIC;
    SIGNAL S3369 : STD_LOGIC;
    SIGNAL S3370 : STD_LOGIC;
    SIGNAL S3371 : STD_LOGIC;
    SIGNAL S3372 : STD_LOGIC;
    SIGNAL S3373 : STD_LOGIC;
    SIGNAL S3374 : STD_LOGIC;
    SIGNAL S3375 : STD_LOGIC;
    SIGNAL S3376 : STD_LOGIC;
    SIGNAL S3377 : STD_LOGIC;
    SIGNAL S3378 : STD_LOGIC;
    SIGNAL S3379 : STD_LOGIC;
    SIGNAL S3380 : STD_LOGIC;
    SIGNAL S3381 : STD_LOGIC;
    SIGNAL S3382 : STD_LOGIC;
    SIGNAL S3383 : STD_LOGIC;
    SIGNAL S3384 : STD_LOGIC;
    SIGNAL S3385 : STD_LOGIC;
    SIGNAL S3386 : STD_LOGIC;
    SIGNAL S3387 : STD_LOGIC;
    SIGNAL S3388 : STD_LOGIC;
    SIGNAL S3389 : STD_LOGIC;
    SIGNAL S3390 : STD_LOGIC;
    SIGNAL S3391 : STD_LOGIC;
    SIGNAL S3392 : STD_LOGIC;
    SIGNAL S3393 : STD_LOGIC;
    SIGNAL S3394 : STD_LOGIC;
    SIGNAL S3395 : STD_LOGIC;
    SIGNAL S3396 : STD_LOGIC;
    SIGNAL S3397 : STD_LOGIC;
    SIGNAL S3398 : STD_LOGIC;
    SIGNAL S3399 : STD_LOGIC;
    SIGNAL S3400 : STD_LOGIC;
    SIGNAL S3401 : STD_LOGIC;
    SIGNAL S3402 : STD_LOGIC;
    SIGNAL S3403 : STD_LOGIC;
    SIGNAL S3404 : STD_LOGIC;
    SIGNAL S3405 : STD_LOGIC;
    SIGNAL S3406 : STD_LOGIC;
    SIGNAL S3407 : STD_LOGIC;
    SIGNAL S3408 : STD_LOGIC;
    SIGNAL S3409 : STD_LOGIC;
    SIGNAL S3410 : STD_LOGIC;
    SIGNAL S3411 : STD_LOGIC;
    SIGNAL S3412 : STD_LOGIC;
    SIGNAL S3413 : STD_LOGIC;
    SIGNAL S3414 : STD_LOGIC;
    SIGNAL S3415 : STD_LOGIC;
    SIGNAL S3416 : STD_LOGIC;
    SIGNAL S3417 : STD_LOGIC;
    SIGNAL S3418 : STD_LOGIC;
    SIGNAL S3419 : STD_LOGIC;
    SIGNAL S3420 : STD_LOGIC;
    SIGNAL S3421 : STD_LOGIC;
    SIGNAL S3422 : STD_LOGIC;
    SIGNAL S3423 : STD_LOGIC;
    SIGNAL S3424 : STD_LOGIC;
    SIGNAL S3425 : STD_LOGIC;
    SIGNAL S3426 : STD_LOGIC;
    SIGNAL S3427 : STD_LOGIC;
    SIGNAL S3428 : STD_LOGIC;
    SIGNAL S3429 : STD_LOGIC;
    SIGNAL S3430 : STD_LOGIC;
    SIGNAL S3431 : STD_LOGIC;
    SIGNAL S3432 : STD_LOGIC;
    SIGNAL S3433 : STD_LOGIC;
    SIGNAL S3434 : STD_LOGIC;
    SIGNAL S3435 : STD_LOGIC;
    SIGNAL S3436 : STD_LOGIC;
    SIGNAL S3437 : STD_LOGIC;
    SIGNAL S3438 : STD_LOGIC;
    SIGNAL S3439 : STD_LOGIC;
    SIGNAL S3440 : STD_LOGIC;
    SIGNAL S3441 : STD_LOGIC;
    SIGNAL S3442 : STD_LOGIC;
    SIGNAL S3443 : STD_LOGIC;
    SIGNAL S3444 : STD_LOGIC;
    SIGNAL S3445 : STD_LOGIC;
    SIGNAL S3446 : STD_LOGIC;
    SIGNAL S3447 : STD_LOGIC;
    SIGNAL S3448 : STD_LOGIC;
    SIGNAL S3449 : STD_LOGIC;
    SIGNAL S3450 : STD_LOGIC;
    SIGNAL S3451 : STD_LOGIC;
    SIGNAL S3452 : STD_LOGIC;
    SIGNAL S3453 : STD_LOGIC;
    SIGNAL S3454 : STD_LOGIC;
    SIGNAL S3455 : STD_LOGIC;
    SIGNAL S3456 : STD_LOGIC;
    SIGNAL S3457 : STD_LOGIC;
    SIGNAL S3458 : STD_LOGIC;
    SIGNAL S3459 : STD_LOGIC;
    SIGNAL S3460 : STD_LOGIC;
    SIGNAL S3461 : STD_LOGIC;
    SIGNAL S3462 : STD_LOGIC;
    SIGNAL S3463 : STD_LOGIC;
    SIGNAL S3464 : STD_LOGIC;
    SIGNAL S3465 : STD_LOGIC;
    SIGNAL S3466 : STD_LOGIC;
    SIGNAL S3467 : STD_LOGIC;
    SIGNAL S3468 : STD_LOGIC;
    SIGNAL S3469 : STD_LOGIC;
    SIGNAL S3470 : STD_LOGIC;
    SIGNAL S3471 : STD_LOGIC;
    SIGNAL S3472 : STD_LOGIC;
    SIGNAL S3473 : STD_LOGIC;
    SIGNAL S3474 : STD_LOGIC;
    SIGNAL S3475 : STD_LOGIC;
    SIGNAL S3476 : STD_LOGIC;
    SIGNAL S3477 : STD_LOGIC;
    SIGNAL S3478 : STD_LOGIC;
    SIGNAL S3479 : STD_LOGIC;
    SIGNAL S3480 : STD_LOGIC;
    SIGNAL S3481 : STD_LOGIC;
    SIGNAL S3482 : STD_LOGIC;
    SIGNAL S3483 : STD_LOGIC;
    SIGNAL S3484 : STD_LOGIC;
    SIGNAL S3485 : STD_LOGIC;
    SIGNAL S3486 : STD_LOGIC;
    SIGNAL S3487 : STD_LOGIC;
    SIGNAL S3488 : STD_LOGIC;
    SIGNAL S3489 : STD_LOGIC;
    SIGNAL S3490 : STD_LOGIC;
    SIGNAL S3491 : STD_LOGIC;
    SIGNAL S3492 : STD_LOGIC;
    SIGNAL S3493 : STD_LOGIC;
    SIGNAL S3494 : STD_LOGIC;
    SIGNAL S3495 : STD_LOGIC;
    SIGNAL S3496 : STD_LOGIC;
    SIGNAL S3497 : STD_LOGIC;
    SIGNAL S3498 : STD_LOGIC;
    SIGNAL S3499 : STD_LOGIC;
    SIGNAL S3500 : STD_LOGIC;
    SIGNAL S3501 : STD_LOGIC;
    SIGNAL S3502 : STD_LOGIC;
    SIGNAL S3503 : STD_LOGIC;
    SIGNAL S3504 : STD_LOGIC;
    SIGNAL S3505 : STD_LOGIC;
    SIGNAL S3506 : STD_LOGIC;
    SIGNAL S3507 : STD_LOGIC;
    SIGNAL S3508 : STD_LOGIC;
    SIGNAL S3509 : STD_LOGIC;
    SIGNAL S3510 : STD_LOGIC;
    SIGNAL S3511 : STD_LOGIC;
    SIGNAL S3512 : STD_LOGIC;
    SIGNAL S3513 : STD_LOGIC;
    SIGNAL S3514 : STD_LOGIC;
    SIGNAL S3515 : STD_LOGIC;
    SIGNAL S3516 : STD_LOGIC;
    SIGNAL S3517 : STD_LOGIC;
    SIGNAL S3518 : STD_LOGIC;
    SIGNAL S3519 : STD_LOGIC;
    SIGNAL S3520 : STD_LOGIC;
    SIGNAL S3521 : STD_LOGIC;
    SIGNAL S3522 : STD_LOGIC;
    SIGNAL S3523 : STD_LOGIC;
    SIGNAL S3524 : STD_LOGIC;
    SIGNAL S3525 : STD_LOGIC;
    SIGNAL S3526 : STD_LOGIC;
    SIGNAL S3527 : STD_LOGIC;
    SIGNAL S3528 : STD_LOGIC;
    SIGNAL S3529 : STD_LOGIC;
    SIGNAL S3530 : STD_LOGIC;
    SIGNAL S3531 : STD_LOGIC;
    SIGNAL S3532 : STD_LOGIC;
    SIGNAL S3533 : STD_LOGIC;
    SIGNAL S3534 : STD_LOGIC;
    SIGNAL S3535 : STD_LOGIC;
    SIGNAL S3536 : STD_LOGIC;
    SIGNAL S3537 : STD_LOGIC;
    SIGNAL S3538 : STD_LOGIC;
    SIGNAL S3539 : STD_LOGIC;
    SIGNAL S3540 : STD_LOGIC;
    SIGNAL S3541 : STD_LOGIC;
    SIGNAL S3542 : STD_LOGIC;
    SIGNAL S3543 : STD_LOGIC;
    SIGNAL S3544 : STD_LOGIC;
    SIGNAL S3545 : STD_LOGIC;
    SIGNAL S3546 : STD_LOGIC;
    SIGNAL S3547 : STD_LOGIC;
    SIGNAL S3548 : STD_LOGIC;
    SIGNAL S3549 : STD_LOGIC;
    SIGNAL S3550 : STD_LOGIC;
    SIGNAL S3551 : STD_LOGIC;
    SIGNAL S3552 : STD_LOGIC;
    SIGNAL S3553 : STD_LOGIC;
    SIGNAL S3554 : STD_LOGIC;
    SIGNAL S3555 : STD_LOGIC;
    SIGNAL S3556 : STD_LOGIC;
    SIGNAL S3557 : STD_LOGIC;
    SIGNAL S3558 : STD_LOGIC;
    SIGNAL S3559 : STD_LOGIC;
    SIGNAL S3560 : STD_LOGIC;
    SIGNAL S3561 : STD_LOGIC;
    SIGNAL S3562 : STD_LOGIC;
    SIGNAL S3563 : STD_LOGIC;
    SIGNAL S3564 : STD_LOGIC;
    SIGNAL S3565 : STD_LOGIC;
    SIGNAL S3566 : STD_LOGIC;
    SIGNAL S3567 : STD_LOGIC;
    SIGNAL S3568 : STD_LOGIC;
    SIGNAL S3569 : STD_LOGIC;
    SIGNAL S3570 : STD_LOGIC;
    SIGNAL S3571 : STD_LOGIC;
    SIGNAL S3572 : STD_LOGIC;
    SIGNAL S3573 : STD_LOGIC;
    SIGNAL S3574 : STD_LOGIC;
    SIGNAL S3575 : STD_LOGIC;
    SIGNAL S3576 : STD_LOGIC;
    SIGNAL S3577 : STD_LOGIC;
    SIGNAL S3578 : STD_LOGIC;
    SIGNAL S3579 : STD_LOGIC;
    SIGNAL S3580 : STD_LOGIC;
    SIGNAL S3581 : STD_LOGIC;
    SIGNAL S3582 : STD_LOGIC;
    SIGNAL S3583 : STD_LOGIC;
    SIGNAL S3584 : STD_LOGIC;
    SIGNAL S3585 : STD_LOGIC;
    SIGNAL S3586 : STD_LOGIC;
    SIGNAL S3587 : STD_LOGIC;
    SIGNAL S3588 : STD_LOGIC;
    SIGNAL S3589 : STD_LOGIC;
    SIGNAL S3590 : STD_LOGIC;
    SIGNAL S3591 : STD_LOGIC;
    SIGNAL S3592 : STD_LOGIC;
    SIGNAL S3593 : STD_LOGIC;
    SIGNAL S3594 : STD_LOGIC;
    SIGNAL S3595 : STD_LOGIC;
    SIGNAL S3596 : STD_LOGIC;
    SIGNAL S3597 : STD_LOGIC;
    SIGNAL S3598 : STD_LOGIC;
    SIGNAL S3599 : STD_LOGIC;
    SIGNAL S3600 : STD_LOGIC;
    SIGNAL S3601 : STD_LOGIC;
    SIGNAL S3602 : STD_LOGIC;
    SIGNAL S3603 : STD_LOGIC;
    SIGNAL S3604 : STD_LOGIC;
    SIGNAL S3605 : STD_LOGIC;
    SIGNAL S3606 : STD_LOGIC;
    SIGNAL S3607 : STD_LOGIC;
    SIGNAL S3608 : STD_LOGIC;
    SIGNAL S3609 : STD_LOGIC;
    SIGNAL S3610 : STD_LOGIC;
    SIGNAL S3611 : STD_LOGIC;
    SIGNAL S3612 : STD_LOGIC;
    SIGNAL S3613 : STD_LOGIC;
    SIGNAL S3614 : STD_LOGIC;
    SIGNAL S3615 : STD_LOGIC;
    SIGNAL S3616 : STD_LOGIC;
    SIGNAL S3617 : STD_LOGIC;
    SIGNAL S3618 : STD_LOGIC;
    SIGNAL S3619 : STD_LOGIC;
    SIGNAL S3620 : STD_LOGIC;
    SIGNAL S3621 : STD_LOGIC;
    SIGNAL S3622 : STD_LOGIC;
    SIGNAL S3623 : STD_LOGIC;
    SIGNAL S3624 : STD_LOGIC;
    SIGNAL S3625 : STD_LOGIC;
    SIGNAL S3626 : STD_LOGIC;
    SIGNAL S3627 : STD_LOGIC;
    SIGNAL S3628 : STD_LOGIC;
    SIGNAL S3629 : STD_LOGIC;
    SIGNAL S3630 : STD_LOGIC;
    SIGNAL S3631 : STD_LOGIC;
    SIGNAL S3632 : STD_LOGIC;
    SIGNAL S3633 : STD_LOGIC;
    SIGNAL S3634 : STD_LOGIC;
    SIGNAL S3635 : STD_LOGIC;
    SIGNAL S3636 : STD_LOGIC;
    SIGNAL S3637 : STD_LOGIC;
    SIGNAL S3638 : STD_LOGIC;
    SIGNAL S3639 : STD_LOGIC;
    SIGNAL S3640 : STD_LOGIC;
    SIGNAL S3641 : STD_LOGIC;
    SIGNAL S3642 : STD_LOGIC;
    SIGNAL S3643 : STD_LOGIC;
    SIGNAL S3644 : STD_LOGIC;
    SIGNAL S3645 : STD_LOGIC;
    SIGNAL S3646 : STD_LOGIC;
    SIGNAL S3647 : STD_LOGIC;
    SIGNAL S3648 : STD_LOGIC;
    SIGNAL S3649 : STD_LOGIC;
    SIGNAL S3650 : STD_LOGIC;
    SIGNAL S3651 : STD_LOGIC;
    SIGNAL S3652 : STD_LOGIC;
    SIGNAL S3653 : STD_LOGIC;
    SIGNAL S3654 : STD_LOGIC;
    SIGNAL S3655 : STD_LOGIC;
    SIGNAL S3656 : STD_LOGIC;
    SIGNAL S3657 : STD_LOGIC;
    SIGNAL S3658 : STD_LOGIC;
    SIGNAL S3659 : STD_LOGIC;
    SIGNAL S3660 : STD_LOGIC;
    SIGNAL S3661 : STD_LOGIC;
    SIGNAL S3662 : STD_LOGIC;
    SIGNAL S3663 : STD_LOGIC;
    SIGNAL S3664 : STD_LOGIC;
    SIGNAL S3665 : STD_LOGIC;
    SIGNAL S3666 : STD_LOGIC;
    SIGNAL S3667 : STD_LOGIC;
    SIGNAL S3668 : STD_LOGIC;
    SIGNAL S3669 : STD_LOGIC;
    SIGNAL S3670 : STD_LOGIC;
    SIGNAL S3671 : STD_LOGIC;
    SIGNAL S3672 : STD_LOGIC;
    SIGNAL S3673 : STD_LOGIC;
    SIGNAL S3674 : STD_LOGIC;
    SIGNAL S3675 : STD_LOGIC;
    SIGNAL S3676 : STD_LOGIC;
    SIGNAL S3677 : STD_LOGIC;
    SIGNAL S3678 : STD_LOGIC;
    SIGNAL S3679 : STD_LOGIC;
    SIGNAL S3680 : STD_LOGIC;
    SIGNAL S3681 : STD_LOGIC;
    SIGNAL S3682 : STD_LOGIC;
    SIGNAL S3683 : STD_LOGIC;
    SIGNAL S3684 : STD_LOGIC;
    SIGNAL S3685 : STD_LOGIC;
    SIGNAL S3686 : STD_LOGIC;
    SIGNAL S3687 : STD_LOGIC;
    SIGNAL S3688 : STD_LOGIC;
    SIGNAL S3689 : STD_LOGIC;
    SIGNAL S3690 : STD_LOGIC;
    SIGNAL S3691 : STD_LOGIC;
    SIGNAL S3692 : STD_LOGIC;
    SIGNAL S3693 : STD_LOGIC;
    SIGNAL S3694 : STD_LOGIC;
    SIGNAL S3695 : STD_LOGIC;
    SIGNAL S3696 : STD_LOGIC;
    SIGNAL S3697 : STD_LOGIC;
    SIGNAL S3698 : STD_LOGIC;
    SIGNAL S3699 : STD_LOGIC;
    SIGNAL S3700 : STD_LOGIC;
    SIGNAL S3701 : STD_LOGIC;
    SIGNAL S3702 : STD_LOGIC;
    SIGNAL S3703 : STD_LOGIC;
    SIGNAL S3704 : STD_LOGIC;
    SIGNAL S3705 : STD_LOGIC;
    SIGNAL S3706 : STD_LOGIC;
    SIGNAL S3707 : STD_LOGIC;
    SIGNAL S3708 : STD_LOGIC;
    SIGNAL S3709 : STD_LOGIC;
    SIGNAL S3710 : STD_LOGIC;
    SIGNAL S3711 : STD_LOGIC;
    SIGNAL S3712 : STD_LOGIC;
    SIGNAL S3713 : STD_LOGIC;
    SIGNAL S3714 : STD_LOGIC;
    SIGNAL S3715 : STD_LOGIC;
    SIGNAL S3716 : STD_LOGIC;
    SIGNAL S3717 : STD_LOGIC;
    SIGNAL S3718 : STD_LOGIC;
    SIGNAL S3719 : STD_LOGIC;
    SIGNAL S3720 : STD_LOGIC;
    SIGNAL S3721 : STD_LOGIC;
    SIGNAL S3722 : STD_LOGIC;
    SIGNAL S3723 : STD_LOGIC;
    SIGNAL S3724 : STD_LOGIC;
    SIGNAL S3725 : STD_LOGIC;
    SIGNAL S3726 : STD_LOGIC;
    SIGNAL S3727 : STD_LOGIC;
    SIGNAL S3728 : STD_LOGIC;
    SIGNAL S3729 : STD_LOGIC;
    SIGNAL S3730 : STD_LOGIC;
    SIGNAL S3731 : STD_LOGIC;
    SIGNAL S3732 : STD_LOGIC;
    SIGNAL S3733 : STD_LOGIC;
    SIGNAL S3734 : STD_LOGIC;
    SIGNAL S3735 : STD_LOGIC;
    SIGNAL S3736 : STD_LOGIC;
    SIGNAL S3737 : STD_LOGIC;
    SIGNAL S3738 : STD_LOGIC;
    SIGNAL S3739 : STD_LOGIC;
    SIGNAL S3740 : STD_LOGIC;
    SIGNAL S3741 : STD_LOGIC;
    SIGNAL S3742 : STD_LOGIC;
    SIGNAL S3743 : STD_LOGIC;
    SIGNAL S3744 : STD_LOGIC;
    SIGNAL S3745 : STD_LOGIC;
    SIGNAL S3746 : STD_LOGIC;
    SIGNAL S3747 : STD_LOGIC;
    SIGNAL S3748 : STD_LOGIC;
    SIGNAL S3749 : STD_LOGIC;
    SIGNAL S3750 : STD_LOGIC;
    SIGNAL S3751 : STD_LOGIC;
    SIGNAL S3752 : STD_LOGIC;
    SIGNAL S3753 : STD_LOGIC;
    SIGNAL S3754 : STD_LOGIC;
    SIGNAL S3755 : STD_LOGIC;
    SIGNAL S3756 : STD_LOGIC;
    SIGNAL S3757 : STD_LOGIC;
    SIGNAL S3758 : STD_LOGIC;
    SIGNAL S3759 : STD_LOGIC;
    SIGNAL S3760 : STD_LOGIC;
    SIGNAL S3761 : STD_LOGIC;
    SIGNAL S3762 : STD_LOGIC;
    SIGNAL S3763 : STD_LOGIC;
    SIGNAL S3764 : STD_LOGIC;
    SIGNAL S3765 : STD_LOGIC;
    SIGNAL S3766 : STD_LOGIC;
    SIGNAL S3767 : STD_LOGIC;
    SIGNAL S3768 : STD_LOGIC;
    SIGNAL S3769 : STD_LOGIC;
    SIGNAL S3770 : STD_LOGIC;
    SIGNAL S3771 : STD_LOGIC;
    SIGNAL S3772 : STD_LOGIC;
    SIGNAL S3773 : STD_LOGIC;
    SIGNAL S3774 : STD_LOGIC;
    SIGNAL S3775 : STD_LOGIC;
    SIGNAL S3776 : STD_LOGIC;
    SIGNAL S3777 : STD_LOGIC;
    SIGNAL S3778 : STD_LOGIC;
    SIGNAL S3779 : STD_LOGIC;
    SIGNAL S3780 : STD_LOGIC;
    SIGNAL S3781 : STD_LOGIC;
    SIGNAL S3782 : STD_LOGIC;
    SIGNAL S3783 : STD_LOGIC;
    SIGNAL S3784 : STD_LOGIC;
    SIGNAL S3785 : STD_LOGIC;
    SIGNAL S3786 : STD_LOGIC;
    SIGNAL S3787 : STD_LOGIC;
    SIGNAL S3788 : STD_LOGIC;
    SIGNAL S3789 : STD_LOGIC;
    SIGNAL S3790 : STD_LOGIC;
    SIGNAL S3791 : STD_LOGIC;
    SIGNAL S3792 : STD_LOGIC;
    SIGNAL S3793 : STD_LOGIC;
    SIGNAL S3794 : STD_LOGIC;
    SIGNAL S3795 : STD_LOGIC;
    SIGNAL S3796 : STD_LOGIC;
    SIGNAL S3797 : STD_LOGIC;
    SIGNAL S3798 : STD_LOGIC;
    SIGNAL S3799 : STD_LOGIC;
    SIGNAL S3800 : STD_LOGIC;
    SIGNAL S3801 : STD_LOGIC;
    SIGNAL S3802 : STD_LOGIC;
    SIGNAL S3803 : STD_LOGIC;
    SIGNAL S3804 : STD_LOGIC;
    SIGNAL S3805 : STD_LOGIC;
    SIGNAL S3806 : STD_LOGIC;
    SIGNAL S3807 : STD_LOGIC;
    SIGNAL S3808 : STD_LOGIC;
    SIGNAL S3809 : STD_LOGIC;
    SIGNAL S3810 : STD_LOGIC;
    SIGNAL S3811 : STD_LOGIC;
    SIGNAL S3812 : STD_LOGIC;
    SIGNAL S3813 : STD_LOGIC;
    SIGNAL S3814 : STD_LOGIC;
    SIGNAL S3815 : STD_LOGIC;
    SIGNAL S3816 : STD_LOGIC;
    SIGNAL S3817 : STD_LOGIC;
    SIGNAL S3818 : STD_LOGIC;
    SIGNAL S3819 : STD_LOGIC;
    SIGNAL S3820 : STD_LOGIC;
    SIGNAL S3821 : STD_LOGIC;
    SIGNAL S3822 : STD_LOGIC;
    SIGNAL S3823 : STD_LOGIC;
    SIGNAL S3824 : STD_LOGIC;
    SIGNAL S3825 : STD_LOGIC;
    SIGNAL S3826 : STD_LOGIC;
    SIGNAL S3827 : STD_LOGIC;
    SIGNAL S3828 : STD_LOGIC;
    SIGNAL S3829 : STD_LOGIC;
    SIGNAL S3830 : STD_LOGIC;
    SIGNAL S3831 : STD_LOGIC;
    SIGNAL S3832 : STD_LOGIC;
    SIGNAL S3833 : STD_LOGIC;
    SIGNAL S3834 : STD_LOGIC;
    SIGNAL S3835 : STD_LOGIC;
    SIGNAL S3836 : STD_LOGIC;
    SIGNAL S3837 : STD_LOGIC;
    SIGNAL S3838 : STD_LOGIC;
    SIGNAL S3839 : STD_LOGIC;
    SIGNAL S3840 : STD_LOGIC;
    SIGNAL S3841 : STD_LOGIC;
    SIGNAL S3842 : STD_LOGIC;
    SIGNAL S3843 : STD_LOGIC;
    SIGNAL S3844 : STD_LOGIC;
    SIGNAL S3845 : STD_LOGIC;
    SIGNAL S3846 : STD_LOGIC;
    SIGNAL S3847 : STD_LOGIC;
    SIGNAL S3848 : STD_LOGIC;
    SIGNAL S3849 : STD_LOGIC;
    SIGNAL S3850 : STD_LOGIC;
    SIGNAL S3851 : STD_LOGIC;
    SIGNAL S3852 : STD_LOGIC;
    SIGNAL S3853 : STD_LOGIC;
    SIGNAL S3854 : STD_LOGIC;
    SIGNAL S3855 : STD_LOGIC;
    SIGNAL S3856 : STD_LOGIC;
    SIGNAL S3857 : STD_LOGIC;
    SIGNAL S3858 : STD_LOGIC;
    SIGNAL S3859 : STD_LOGIC;
    SIGNAL S3860 : STD_LOGIC;
    SIGNAL S3861 : STD_LOGIC;
    SIGNAL S3862 : STD_LOGIC;
    SIGNAL S3863 : STD_LOGIC;
    SIGNAL S3864 : STD_LOGIC;
    SIGNAL S3865 : STD_LOGIC;
    SIGNAL S3866 : STD_LOGIC;
    SIGNAL S3867 : STD_LOGIC;
    SIGNAL S3868 : STD_LOGIC;
    SIGNAL S3869 : STD_LOGIC;
    SIGNAL S3870 : STD_LOGIC;
    SIGNAL S3871 : STD_LOGIC;
    SIGNAL S3872 : STD_LOGIC;
    SIGNAL S3873 : STD_LOGIC;
    SIGNAL S3874 : STD_LOGIC;
    SIGNAL S3875 : STD_LOGIC;
    SIGNAL S3876 : STD_LOGIC;
    SIGNAL S3877 : STD_LOGIC;
    SIGNAL S3878 : STD_LOGIC;
    SIGNAL S3879 : STD_LOGIC;
    SIGNAL S3880 : STD_LOGIC;
    SIGNAL S3881 : STD_LOGIC;
    SIGNAL S3882 : STD_LOGIC;
    SIGNAL S3883 : STD_LOGIC;
    SIGNAL S3884 : STD_LOGIC;
    SIGNAL S3885 : STD_LOGIC;
    SIGNAL S3886 : STD_LOGIC;
    SIGNAL S3887 : STD_LOGIC;
    SIGNAL S3888 : STD_LOGIC;
    SIGNAL S3889 : STD_LOGIC;
    SIGNAL S3890 : STD_LOGIC;
    SIGNAL S3891 : STD_LOGIC;
    SIGNAL S3892 : STD_LOGIC;
    SIGNAL S3893 : STD_LOGIC;
    SIGNAL S3894 : STD_LOGIC;
    SIGNAL S3895 : STD_LOGIC;
    SIGNAL S3896 : STD_LOGIC;
    SIGNAL S3897 : STD_LOGIC;
    SIGNAL S3898 : STD_LOGIC;
    SIGNAL S3899 : STD_LOGIC;
    SIGNAL S3900 : STD_LOGIC;
    SIGNAL S3901 : STD_LOGIC;
    SIGNAL S3902 : STD_LOGIC;
    SIGNAL S3903 : STD_LOGIC;
    SIGNAL S3904 : STD_LOGIC;
    SIGNAL S3905 : STD_LOGIC;
    SIGNAL S3906 : STD_LOGIC;
    SIGNAL S3907 : STD_LOGIC;
    SIGNAL S3908 : STD_LOGIC;
    SIGNAL S3909 : STD_LOGIC;
    SIGNAL S3910 : STD_LOGIC;
    SIGNAL S3911 : STD_LOGIC;
    SIGNAL S3912 : STD_LOGIC;
    SIGNAL S3913 : STD_LOGIC;
    SIGNAL S3914 : STD_LOGIC;
    SIGNAL S3915 : STD_LOGIC;
    SIGNAL S3916 : STD_LOGIC;
    SIGNAL S3917 : STD_LOGIC;
    SIGNAL S3918 : STD_LOGIC;
    SIGNAL S3919 : STD_LOGIC;
    SIGNAL S3920 : STD_LOGIC;
    SIGNAL S3921 : STD_LOGIC;
    SIGNAL S3922 : STD_LOGIC;
    SIGNAL S3923 : STD_LOGIC;
    SIGNAL S3924 : STD_LOGIC;
    SIGNAL S3925 : STD_LOGIC;
    SIGNAL S3926 : STD_LOGIC;
    SIGNAL S3927 : STD_LOGIC;
    SIGNAL S3928 : STD_LOGIC;
    SIGNAL S3929 : STD_LOGIC;
    SIGNAL S3930 : STD_LOGIC;
    SIGNAL S3931 : STD_LOGIC;
    SIGNAL S3932 : STD_LOGIC;
    SIGNAL S3933 : STD_LOGIC;
    SIGNAL S3934 : STD_LOGIC;
    SIGNAL S3935 : STD_LOGIC;
    SIGNAL S3936 : STD_LOGIC;
    SIGNAL S3937 : STD_LOGIC;
    SIGNAL S3938 : STD_LOGIC;
    SIGNAL S3939 : STD_LOGIC;
    SIGNAL S3940 : STD_LOGIC;
    SIGNAL S3941 : STD_LOGIC;
    SIGNAL S3942 : STD_LOGIC;
    SIGNAL S3943 : STD_LOGIC;
    SIGNAL S3944 : STD_LOGIC;
    SIGNAL S3945 : STD_LOGIC;
    SIGNAL S3946 : STD_LOGIC;
    SIGNAL S3947 : STD_LOGIC;
    SIGNAL S3948 : STD_LOGIC;
    SIGNAL S3949 : STD_LOGIC;
    SIGNAL S3950 : STD_LOGIC;
    SIGNAL S3951 : STD_LOGIC;
    SIGNAL S3952 : STD_LOGIC;
    SIGNAL S3953 : STD_LOGIC;
    SIGNAL S3954 : STD_LOGIC;
    SIGNAL S3955 : STD_LOGIC;
    SIGNAL S3956 : STD_LOGIC;
    SIGNAL S3957 : STD_LOGIC;
    SIGNAL S3958 : STD_LOGIC;
    SIGNAL S3959 : STD_LOGIC;
    SIGNAL S3960 : STD_LOGIC;
    SIGNAL S3961 : STD_LOGIC;
    SIGNAL S3962 : STD_LOGIC;
    SIGNAL S3963 : STD_LOGIC;
    SIGNAL S3964 : STD_LOGIC;
    SIGNAL S3965 : STD_LOGIC;
    SIGNAL S3966 : STD_LOGIC;
    SIGNAL S3967 : STD_LOGIC;
    SIGNAL S3968 : STD_LOGIC;
    SIGNAL S3969 : STD_LOGIC;
    SIGNAL S3970 : STD_LOGIC;
    SIGNAL S3971 : STD_LOGIC;
    SIGNAL S3972 : STD_LOGIC;
    SIGNAL S3973 : STD_LOGIC;
    SIGNAL S3974 : STD_LOGIC;
    SIGNAL S3975 : STD_LOGIC;
    SIGNAL S3976 : STD_LOGIC;
    SIGNAL S3977 : STD_LOGIC;
    SIGNAL S3978 : STD_LOGIC;
    SIGNAL S3979 : STD_LOGIC;
    SIGNAL S3980 : STD_LOGIC;
    SIGNAL S3981 : STD_LOGIC;
    SIGNAL S3982 : STD_LOGIC;
    SIGNAL S3983 : STD_LOGIC;
    SIGNAL S3984 : STD_LOGIC;
    SIGNAL S3985 : STD_LOGIC;
    SIGNAL S3986 : STD_LOGIC;
    SIGNAL S3987 : STD_LOGIC;
    SIGNAL S3988 : STD_LOGIC;
    SIGNAL S3989 : STD_LOGIC;
    SIGNAL S3990 : STD_LOGIC;
    SIGNAL S3991 : STD_LOGIC;
    SIGNAL S3992 : STD_LOGIC;
    SIGNAL S3993 : STD_LOGIC;
    SIGNAL S3994 : STD_LOGIC;
    SIGNAL S3995 : STD_LOGIC;
    SIGNAL S3996 : STD_LOGIC;
    SIGNAL S3997 : STD_LOGIC;
    SIGNAL S3998 : STD_LOGIC;
    SIGNAL S3999 : STD_LOGIC;
    SIGNAL S4000 : STD_LOGIC;
    SIGNAL S4001 : STD_LOGIC;
    SIGNAL S4002 : STD_LOGIC;
    SIGNAL S4003 : STD_LOGIC;
    SIGNAL S4004 : STD_LOGIC;
    SIGNAL S4005 : STD_LOGIC;
    SIGNAL S4006 : STD_LOGIC;
    SIGNAL S4007 : STD_LOGIC;
    SIGNAL S4008 : STD_LOGIC;
    SIGNAL S4009 : STD_LOGIC;
    SIGNAL S4010 : STD_LOGIC;
    SIGNAL S4011 : STD_LOGIC;
    SIGNAL S4012 : STD_LOGIC;
    SIGNAL S4013 : STD_LOGIC;
    SIGNAL S4014 : STD_LOGIC;
    SIGNAL S4015 : STD_LOGIC;
    SIGNAL S4016 : STD_LOGIC;
    SIGNAL S4017 : STD_LOGIC;
    SIGNAL S4018 : STD_LOGIC;
    SIGNAL S4019 : STD_LOGIC;
    SIGNAL S4020 : STD_LOGIC;
    SIGNAL S4021 : STD_LOGIC;
    SIGNAL S4022 : STD_LOGIC;
    SIGNAL S4023 : STD_LOGIC;
    SIGNAL S4024 : STD_LOGIC;
    SIGNAL S4025 : STD_LOGIC;
    SIGNAL S4026 : STD_LOGIC;
    SIGNAL S4027 : STD_LOGIC;
    SIGNAL S4028 : STD_LOGIC;
    SIGNAL S4029 : STD_LOGIC;
    SIGNAL S4030 : STD_LOGIC;
    SIGNAL S4031 : STD_LOGIC;
    SIGNAL S4032 : STD_LOGIC;
    SIGNAL S4033 : STD_LOGIC;
    SIGNAL S4034 : STD_LOGIC;
    SIGNAL S4035 : STD_LOGIC;
    SIGNAL S4036 : STD_LOGIC;
    SIGNAL S4037 : STD_LOGIC;
    SIGNAL S4038 : STD_LOGIC;
    SIGNAL S4039 : STD_LOGIC;
    SIGNAL S4040 : STD_LOGIC;
    SIGNAL S4041 : STD_LOGIC;
    SIGNAL S4042 : STD_LOGIC;
    SIGNAL S4043 : STD_LOGIC;
    SIGNAL S4044 : STD_LOGIC;
    SIGNAL S4045 : STD_LOGIC;
    SIGNAL S4046 : STD_LOGIC;
    SIGNAL S4047 : STD_LOGIC;
    SIGNAL S4048 : STD_LOGIC;
    SIGNAL S4049 : STD_LOGIC;
    SIGNAL S4050 : STD_LOGIC;
    SIGNAL S4051 : STD_LOGIC;
    SIGNAL S4052 : STD_LOGIC;
    SIGNAL S4053 : STD_LOGIC;
    SIGNAL S4054 : STD_LOGIC;
    SIGNAL S4055 : STD_LOGIC;
    SIGNAL S4056 : STD_LOGIC;
    SIGNAL S4057 : STD_LOGIC;
    SIGNAL S4058 : STD_LOGIC;
    SIGNAL S4059 : STD_LOGIC;
    SIGNAL S4060 : STD_LOGIC;
    SIGNAL S4061 : STD_LOGIC;
    SIGNAL S4062 : STD_LOGIC;
    SIGNAL S4063 : STD_LOGIC;
    SIGNAL S4064 : STD_LOGIC;
    SIGNAL S4065 : STD_LOGIC;
    SIGNAL S4066 : STD_LOGIC;
    SIGNAL S4067 : STD_LOGIC;
    SIGNAL S4068 : STD_LOGIC;
    SIGNAL S4069 : STD_LOGIC;
    SIGNAL S4070 : STD_LOGIC;
    SIGNAL S4071 : STD_LOGIC;
    SIGNAL S4072 : STD_LOGIC;
    SIGNAL S4073 : STD_LOGIC;
    SIGNAL S4074 : STD_LOGIC;
    SIGNAL S4075 : STD_LOGIC;
    SIGNAL S4076 : STD_LOGIC;
    SIGNAL S4077 : STD_LOGIC;
    SIGNAL S4078 : STD_LOGIC;
    SIGNAL S4079 : STD_LOGIC;
    SIGNAL S4080 : STD_LOGIC;
    SIGNAL S4081 : STD_LOGIC;
    SIGNAL S4082 : STD_LOGIC;
    SIGNAL S4083 : STD_LOGIC;
    SIGNAL S4084 : STD_LOGIC;
    SIGNAL S4085 : STD_LOGIC;
    SIGNAL S4086 : STD_LOGIC;
    SIGNAL S4087 : STD_LOGIC;
    SIGNAL S4088 : STD_LOGIC;
    SIGNAL S4089 : STD_LOGIC;
    SIGNAL S4090 : STD_LOGIC;
    SIGNAL S4091 : STD_LOGIC;
    SIGNAL S4092 : STD_LOGIC;
    SIGNAL S4093 : STD_LOGIC;
    SIGNAL S4094 : STD_LOGIC;
    SIGNAL S4095 : STD_LOGIC;
    SIGNAL S4096 : STD_LOGIC;
    SIGNAL S4097 : STD_LOGIC;
    SIGNAL S4098 : STD_LOGIC;
    SIGNAL S4099 : STD_LOGIC;
    SIGNAL S4100 : STD_LOGIC;
    SIGNAL S4101 : STD_LOGIC;
    SIGNAL S4102 : STD_LOGIC;
    SIGNAL S4103 : STD_LOGIC;
    SIGNAL S4104 : STD_LOGIC;
    SIGNAL S4105 : STD_LOGIC;
    SIGNAL S4106 : STD_LOGIC;
    SIGNAL S4107 : STD_LOGIC;
    SIGNAL S4108 : STD_LOGIC;
    SIGNAL S4109 : STD_LOGIC;
    SIGNAL S4110 : STD_LOGIC;
    SIGNAL S4111 : STD_LOGIC;
    SIGNAL S4112 : STD_LOGIC;
    SIGNAL S4113 : STD_LOGIC;
    SIGNAL S4114 : STD_LOGIC;
    SIGNAL S4115 : STD_LOGIC;
    SIGNAL S4116 : STD_LOGIC;
    SIGNAL S4117 : STD_LOGIC;
    SIGNAL S4118 : STD_LOGIC;
    SIGNAL S4119 : STD_LOGIC;
    SIGNAL S4120 : STD_LOGIC;
    SIGNAL S4121 : STD_LOGIC;
    SIGNAL S4122 : STD_LOGIC;
    SIGNAL S4123 : STD_LOGIC;
    SIGNAL S4124 : STD_LOGIC;
    SIGNAL S4125 : STD_LOGIC;
    SIGNAL S4126 : STD_LOGIC;
    SIGNAL S4127 : STD_LOGIC;
    SIGNAL S4128 : STD_LOGIC;
    SIGNAL S4129 : STD_LOGIC;
    SIGNAL S4130 : STD_LOGIC;
    SIGNAL S4131 : STD_LOGIC;
    SIGNAL S4132 : STD_LOGIC;
    SIGNAL S4133 : STD_LOGIC;
    SIGNAL S4134 : STD_LOGIC;
    SIGNAL S4135 : STD_LOGIC;
    SIGNAL S4136 : STD_LOGIC;
    SIGNAL S4137 : STD_LOGIC;
    SIGNAL S4138 : STD_LOGIC;
    SIGNAL S4139 : STD_LOGIC;
    SIGNAL S4140 : STD_LOGIC;
    SIGNAL S4141 : STD_LOGIC;
    SIGNAL S4142 : STD_LOGIC;
    SIGNAL S4143 : STD_LOGIC;
    SIGNAL S4144 : STD_LOGIC;
    SIGNAL S4145 : STD_LOGIC;
    SIGNAL S4146 : STD_LOGIC;
    SIGNAL S4147 : STD_LOGIC;
    SIGNAL S4148 : STD_LOGIC;
    SIGNAL S4149 : STD_LOGIC;
    SIGNAL S4150 : STD_LOGIC;
    SIGNAL S4151 : STD_LOGIC;
    SIGNAL S4152 : STD_LOGIC;
    SIGNAL S4153 : STD_LOGIC;
    SIGNAL S4154 : STD_LOGIC;
    SIGNAL S4155 : STD_LOGIC;
    SIGNAL S4156 : STD_LOGIC;
    SIGNAL S4157 : STD_LOGIC;
    SIGNAL S4158 : STD_LOGIC;
    SIGNAL S4159 : STD_LOGIC;
    SIGNAL S4160 : STD_LOGIC;
    SIGNAL S4161 : STD_LOGIC;
    SIGNAL S4162 : STD_LOGIC;
    SIGNAL S4163 : STD_LOGIC;
    SIGNAL S4164 : STD_LOGIC;
    SIGNAL S4165 : STD_LOGIC;
    SIGNAL S4166 : STD_LOGIC;
    SIGNAL S4167 : STD_LOGIC;
    SIGNAL S4168 : STD_LOGIC;
    SIGNAL S4169 : STD_LOGIC;
    SIGNAL S4170 : STD_LOGIC;
    SIGNAL S4171 : STD_LOGIC;
    SIGNAL S4172 : STD_LOGIC;
    SIGNAL S4173 : STD_LOGIC;
    SIGNAL S4174 : STD_LOGIC;
    SIGNAL S4175 : STD_LOGIC;
    SIGNAL S4176 : STD_LOGIC;
    SIGNAL S4177 : STD_LOGIC;
    SIGNAL S4178 : STD_LOGIC;
    SIGNAL S4179 : STD_LOGIC;
    SIGNAL S4180 : STD_LOGIC;
    SIGNAL S4181 : STD_LOGIC;
    SIGNAL S4182 : STD_LOGIC;
    SIGNAL S4183 : STD_LOGIC;
    SIGNAL S4184 : STD_LOGIC;
    SIGNAL S4185 : STD_LOGIC;
    SIGNAL S4186 : STD_LOGIC;
    SIGNAL S4187 : STD_LOGIC;
    SIGNAL S4188 : STD_LOGIC;
    SIGNAL S4189 : STD_LOGIC;
    SIGNAL S4190 : STD_LOGIC;
    SIGNAL S4191 : STD_LOGIC;
    SIGNAL S4192 : STD_LOGIC;
    SIGNAL S4193 : STD_LOGIC;
    SIGNAL S4194 : STD_LOGIC;
    SIGNAL S4195 : STD_LOGIC;
    SIGNAL S4196 : STD_LOGIC;
    SIGNAL S4197 : STD_LOGIC;
    SIGNAL S4198 : STD_LOGIC;
    SIGNAL S4199 : STD_LOGIC;
    SIGNAL S4200 : STD_LOGIC;
    SIGNAL S4201 : STD_LOGIC;
    SIGNAL S4202 : STD_LOGIC;
    SIGNAL S4203 : STD_LOGIC;
    SIGNAL S4204 : STD_LOGIC;
    SIGNAL S4205 : STD_LOGIC;
    SIGNAL S4206 : STD_LOGIC;
    SIGNAL S4207 : STD_LOGIC;
    SIGNAL S4208 : STD_LOGIC;
    SIGNAL S4209 : STD_LOGIC;
    SIGNAL S4210 : STD_LOGIC;
    SIGNAL S4211 : STD_LOGIC;
    SIGNAL S4212 : STD_LOGIC;
    SIGNAL S4213 : STD_LOGIC;
    SIGNAL S4214 : STD_LOGIC;
    SIGNAL S4215 : STD_LOGIC;
    SIGNAL S4216 : STD_LOGIC;
    SIGNAL S4217 : STD_LOGIC;
    SIGNAL S4218 : STD_LOGIC;
    SIGNAL S4219 : STD_LOGIC;
    SIGNAL S4220 : STD_LOGIC;
    SIGNAL S4221 : STD_LOGIC;
    SIGNAL S4222 : STD_LOGIC;
    SIGNAL S4223 : STD_LOGIC;
    SIGNAL S4224 : STD_LOGIC;
    SIGNAL S4225 : STD_LOGIC;
    SIGNAL S4226 : STD_LOGIC;
    SIGNAL S4227 : STD_LOGIC;
    SIGNAL S4228 : STD_LOGIC;
    SIGNAL S4229 : STD_LOGIC;
    SIGNAL S4230 : STD_LOGIC;
    SIGNAL S4231 : STD_LOGIC;
    SIGNAL S4232 : STD_LOGIC;
    SIGNAL S4233 : STD_LOGIC;
    SIGNAL S4234 : STD_LOGIC;
    SIGNAL S4235 : STD_LOGIC;
    SIGNAL S4236 : STD_LOGIC;
    SIGNAL S4237 : STD_LOGIC;
    SIGNAL S4238 : STD_LOGIC;
    SIGNAL S4239 : STD_LOGIC;
    SIGNAL S4240 : STD_LOGIC;
    SIGNAL S4241 : STD_LOGIC;
    SIGNAL S4242 : STD_LOGIC;
    SIGNAL S4243 : STD_LOGIC;
    SIGNAL S4244 : STD_LOGIC;
    SIGNAL S4245 : STD_LOGIC;
    SIGNAL S4246 : STD_LOGIC;
    SIGNAL S4247 : STD_LOGIC;
    SIGNAL S4248 : STD_LOGIC;
    SIGNAL S4249 : STD_LOGIC;
    SIGNAL S4250 : STD_LOGIC;
    SIGNAL S4251 : STD_LOGIC;
    SIGNAL S4252 : STD_LOGIC;
    SIGNAL S4253 : STD_LOGIC;
    SIGNAL S4254 : STD_LOGIC;
    SIGNAL S4255 : STD_LOGIC;
    SIGNAL S4256 : STD_LOGIC;
    SIGNAL S4257 : STD_LOGIC;
    SIGNAL S4258 : STD_LOGIC;
    SIGNAL S4259 : STD_LOGIC;
    SIGNAL S4260 : STD_LOGIC;
    SIGNAL S4261 : STD_LOGIC;
    SIGNAL S4262 : STD_LOGIC;
    SIGNAL S4263 : STD_LOGIC;
    SIGNAL S4264 : STD_LOGIC;
    SIGNAL S4265 : STD_LOGIC;
    SIGNAL S4266 : STD_LOGIC;
    SIGNAL S4267 : STD_LOGIC;
    SIGNAL S4268 : STD_LOGIC;
    SIGNAL S4269 : STD_LOGIC;
    SIGNAL S4270 : STD_LOGIC;
    SIGNAL S4271 : STD_LOGIC;
    SIGNAL S4272 : STD_LOGIC;
    SIGNAL S4273 : STD_LOGIC;
    SIGNAL S4274 : STD_LOGIC;
    SIGNAL S4275 : STD_LOGIC;
    SIGNAL S4276 : STD_LOGIC;
    SIGNAL S4277 : STD_LOGIC;
    SIGNAL S4278 : STD_LOGIC;
    SIGNAL S4279 : STD_LOGIC;
    SIGNAL S4280 : STD_LOGIC;
    SIGNAL S4281 : STD_LOGIC;
    SIGNAL S4282 : STD_LOGIC;
    SIGNAL S4283 : STD_LOGIC;
    SIGNAL S4284 : STD_LOGIC;
    SIGNAL S4285 : STD_LOGIC;
    SIGNAL S4286 : STD_LOGIC;
    SIGNAL S4287 : STD_LOGIC;
    SIGNAL S4288 : STD_LOGIC;
    SIGNAL S4289 : STD_LOGIC;
    SIGNAL S4290 : STD_LOGIC;
    SIGNAL S4291 : STD_LOGIC;
    SIGNAL S4292 : STD_LOGIC;
    SIGNAL S4293 : STD_LOGIC;
    SIGNAL S4294 : STD_LOGIC;
    SIGNAL S4295 : STD_LOGIC;
    SIGNAL S4296 : STD_LOGIC;
    SIGNAL S4297 : STD_LOGIC;
    SIGNAL S4298 : STD_LOGIC;
    SIGNAL S4299 : STD_LOGIC;
    SIGNAL S4300 : STD_LOGIC;
    SIGNAL S4301 : STD_LOGIC;
    SIGNAL S4302 : STD_LOGIC;
    SIGNAL S4303 : STD_LOGIC;
    SIGNAL S4304 : STD_LOGIC;
    SIGNAL S4305 : STD_LOGIC;
    SIGNAL S4306 : STD_LOGIC;
    SIGNAL S4307 : STD_LOGIC;
    SIGNAL S4308 : STD_LOGIC;
    SIGNAL S4309 : STD_LOGIC;
    SIGNAL S4310 : STD_LOGIC;
    SIGNAL S4311 : STD_LOGIC;
    SIGNAL S4312 : STD_LOGIC;
    SIGNAL S4313 : STD_LOGIC;
    SIGNAL S4314 : STD_LOGIC;
    SIGNAL S4315 : STD_LOGIC;
    SIGNAL S4316 : STD_LOGIC;
    SIGNAL S4317 : STD_LOGIC;
    SIGNAL S4318 : STD_LOGIC;
    SIGNAL S4319 : STD_LOGIC;
    SIGNAL S4320 : STD_LOGIC;
    SIGNAL S4321 : STD_LOGIC;
    SIGNAL S4322 : STD_LOGIC;
    SIGNAL S4323 : STD_LOGIC;
    SIGNAL S4324 : STD_LOGIC;
    SIGNAL S4325 : STD_LOGIC;
    SIGNAL S4326 : STD_LOGIC;
    SIGNAL S4327 : STD_LOGIC;
    SIGNAL S4328 : STD_LOGIC;
    SIGNAL S4329 : STD_LOGIC;
    SIGNAL S4330 : STD_LOGIC;
    SIGNAL S4331 : STD_LOGIC;
    SIGNAL S4332 : STD_LOGIC;
    SIGNAL S4333 : STD_LOGIC;
    SIGNAL S4334 : STD_LOGIC;
    SIGNAL S4335 : STD_LOGIC;
    SIGNAL S4336 : STD_LOGIC;
    SIGNAL S4337 : STD_LOGIC;
    SIGNAL S4338 : STD_LOGIC;
    SIGNAL S4339 : STD_LOGIC;
    SIGNAL S4340 : STD_LOGIC;
    SIGNAL S4341 : STD_LOGIC;
    SIGNAL S4342 : STD_LOGIC;
    SIGNAL S4343 : STD_LOGIC;
    SIGNAL S4344 : STD_LOGIC;
    SIGNAL S4345 : STD_LOGIC;
    SIGNAL S4346 : STD_LOGIC;
    SIGNAL S4347 : STD_LOGIC;
    SIGNAL S4348 : STD_LOGIC;
    SIGNAL S4349 : STD_LOGIC;
    SIGNAL S4350 : STD_LOGIC;
    SIGNAL S4351 : STD_LOGIC;
    SIGNAL S4352 : STD_LOGIC;
    SIGNAL S4353 : STD_LOGIC;
    SIGNAL S4354 : STD_LOGIC;
    SIGNAL S4355 : STD_LOGIC;
    SIGNAL S4356 : STD_LOGIC;
    SIGNAL S4357 : STD_LOGIC;
    SIGNAL S4358 : STD_LOGIC;
    SIGNAL S4359 : STD_LOGIC;
    SIGNAL S4360 : STD_LOGIC;
    SIGNAL S4361 : STD_LOGIC;
    SIGNAL S4362 : STD_LOGIC;
    SIGNAL S4363 : STD_LOGIC;
    SIGNAL S4364 : STD_LOGIC;
    SIGNAL S4365 : STD_LOGIC;
    SIGNAL S4366 : STD_LOGIC;
    SIGNAL S4367 : STD_LOGIC;
    SIGNAL S4368 : STD_LOGIC;
    SIGNAL S4369 : STD_LOGIC;
    SIGNAL S4370 : STD_LOGIC;
    SIGNAL S4371 : STD_LOGIC;
    SIGNAL S4372 : STD_LOGIC;
    SIGNAL S4373 : STD_LOGIC;
    SIGNAL S4374 : STD_LOGIC;
    SIGNAL S4375 : STD_LOGIC;
    SIGNAL S4376 : STD_LOGIC;
    SIGNAL S4377 : STD_LOGIC;
    SIGNAL S4378 : STD_LOGIC;
    SIGNAL S4379 : STD_LOGIC;
    SIGNAL S4380 : STD_LOGIC;
    SIGNAL S4381 : STD_LOGIC;
    SIGNAL S4382 : STD_LOGIC;
    SIGNAL S4383 : STD_LOGIC;
    SIGNAL S4384 : STD_LOGIC;
    SIGNAL S4385 : STD_LOGIC;
    SIGNAL S4386 : STD_LOGIC;
    SIGNAL S4387 : STD_LOGIC;
    SIGNAL S4388 : STD_LOGIC;
    SIGNAL S4389 : STD_LOGIC;
    SIGNAL S4390 : STD_LOGIC;
    SIGNAL S4391 : STD_LOGIC;
    SIGNAL S4392 : STD_LOGIC;
    SIGNAL S4393 : STD_LOGIC;
    SIGNAL S4394 : STD_LOGIC;
    SIGNAL S4395 : STD_LOGIC;
    SIGNAL S4396 : STD_LOGIC;
    SIGNAL S4397 : STD_LOGIC;
    SIGNAL S4398 : STD_LOGIC;
    SIGNAL S4399 : STD_LOGIC;
    SIGNAL S4400 : STD_LOGIC;
    SIGNAL S4401 : STD_LOGIC;
    SIGNAL S4402 : STD_LOGIC;
    SIGNAL S4403 : STD_LOGIC;
    SIGNAL S4404 : STD_LOGIC;
    SIGNAL S4405 : STD_LOGIC;
    SIGNAL S4406 : STD_LOGIC;
    SIGNAL S4407 : STD_LOGIC;
    SIGNAL S4408 : STD_LOGIC;
    SIGNAL S4409 : STD_LOGIC;
    SIGNAL S4410 : STD_LOGIC;
    SIGNAL S4411 : STD_LOGIC;
    SIGNAL S4412 : STD_LOGIC;
    SIGNAL S4413 : STD_LOGIC;
    SIGNAL S4414 : STD_LOGIC;
    SIGNAL S4415 : STD_LOGIC;
    SIGNAL S4416 : STD_LOGIC;
    SIGNAL S4417 : STD_LOGIC;
    SIGNAL S4418 : STD_LOGIC;
    SIGNAL S4419 : STD_LOGIC;
    SIGNAL S4420 : STD_LOGIC;
    SIGNAL S4421 : STD_LOGIC;
    SIGNAL S4422 : STD_LOGIC;
    SIGNAL S4423 : STD_LOGIC;
    SIGNAL S4424 : STD_LOGIC;
    SIGNAL S4425 : STD_LOGIC;
    SIGNAL S4426 : STD_LOGIC;
    SIGNAL S4427 : STD_LOGIC;
    SIGNAL S4428 : STD_LOGIC;
    SIGNAL S4429 : STD_LOGIC;
    SIGNAL S4430 : STD_LOGIC;
    SIGNAL S4431 : STD_LOGIC;
    SIGNAL S4432 : STD_LOGIC;
    SIGNAL S4433 : STD_LOGIC;
    SIGNAL S4434 : STD_LOGIC;
    SIGNAL S4435 : STD_LOGIC;
    SIGNAL S4436 : STD_LOGIC;
    SIGNAL S4437 : STD_LOGIC;
    SIGNAL S4438 : STD_LOGIC;
    SIGNAL S4439 : STD_LOGIC;
    SIGNAL S4440 : STD_LOGIC;
    SIGNAL S4441 : STD_LOGIC;
    SIGNAL S4442 : STD_LOGIC;
    SIGNAL S4443 : STD_LOGIC;
    SIGNAL S4444 : STD_LOGIC;
    SIGNAL S4445 : STD_LOGIC;
    SIGNAL S4446 : STD_LOGIC;
    SIGNAL S4447 : STD_LOGIC;
    SIGNAL S4448 : STD_LOGIC;
    SIGNAL S4449 : STD_LOGIC;
    SIGNAL S4450 : STD_LOGIC;
    SIGNAL S4451 : STD_LOGIC;
    SIGNAL S4452 : STD_LOGIC;
    SIGNAL S4453 : STD_LOGIC;
    SIGNAL S4454 : STD_LOGIC;
    SIGNAL S4455 : STD_LOGIC;
    SIGNAL S4456 : STD_LOGIC;
    SIGNAL S4457 : STD_LOGIC;
    SIGNAL S4458 : STD_LOGIC;
    SIGNAL S4459 : STD_LOGIC;
    SIGNAL S4460 : STD_LOGIC;
    SIGNAL S4461 : STD_LOGIC;
    SIGNAL S4462 : STD_LOGIC;
    SIGNAL S4463 : STD_LOGIC;
    SIGNAL S4464 : STD_LOGIC;
    SIGNAL S4465 : STD_LOGIC;
    SIGNAL S4466 : STD_LOGIC;
    SIGNAL S4467 : STD_LOGIC;
    SIGNAL S4468 : STD_LOGIC;
    SIGNAL S4469 : STD_LOGIC;
    SIGNAL S4470 : STD_LOGIC;
    SIGNAL S4471 : STD_LOGIC;
    SIGNAL S4472 : STD_LOGIC;
    SIGNAL S4473 : STD_LOGIC;
    SIGNAL S4474 : STD_LOGIC;
    SIGNAL S4475 : STD_LOGIC;
    SIGNAL S4476 : STD_LOGIC;
    SIGNAL S4477 : STD_LOGIC;
    SIGNAL S4478 : STD_LOGIC;
    SIGNAL S4479 : STD_LOGIC;
    SIGNAL S4480 : STD_LOGIC;
    SIGNAL S4481 : STD_LOGIC;
    SIGNAL S4482 : STD_LOGIC;
    SIGNAL S4483 : STD_LOGIC;
    SIGNAL S4484 : STD_LOGIC;
    SIGNAL S4485 : STD_LOGIC;
    SIGNAL S4486 : STD_LOGIC;
    SIGNAL S4487 : STD_LOGIC;
    SIGNAL S4488 : STD_LOGIC;
    SIGNAL S4489 : STD_LOGIC;
    SIGNAL S4490 : STD_LOGIC;
    SIGNAL S4491 : STD_LOGIC;
    SIGNAL S4492 : STD_LOGIC;
    SIGNAL S4493 : STD_LOGIC;
    SIGNAL S4494 : STD_LOGIC;
    SIGNAL S4495 : STD_LOGIC;
    SIGNAL S4496 : STD_LOGIC;
    SIGNAL S4497 : STD_LOGIC;
    SIGNAL S4498 : STD_LOGIC;
    SIGNAL S4499 : STD_LOGIC;
    SIGNAL S4500 : STD_LOGIC;
    SIGNAL S4501 : STD_LOGIC;
    SIGNAL S4502 : STD_LOGIC;
    SIGNAL S4503 : STD_LOGIC;
    SIGNAL S4504 : STD_LOGIC;
    SIGNAL S4505 : STD_LOGIC;
    SIGNAL S4506 : STD_LOGIC;
    SIGNAL S4507 : STD_LOGIC;
    SIGNAL S4508 : STD_LOGIC;
    SIGNAL S4509 : STD_LOGIC;
    SIGNAL S4510 : STD_LOGIC;
    SIGNAL S4511 : STD_LOGIC;
    SIGNAL S4512 : STD_LOGIC;
    SIGNAL S4513 : STD_LOGIC;
    SIGNAL S4514 : STD_LOGIC;
    SIGNAL S4515 : STD_LOGIC;
    SIGNAL S4516 : STD_LOGIC;
    SIGNAL S4517 : STD_LOGIC;
    SIGNAL S4518 : STD_LOGIC;
    SIGNAL S4519 : STD_LOGIC;
    SIGNAL S4520 : STD_LOGIC;
    SIGNAL S4521 : STD_LOGIC;
    SIGNAL S4522 : STD_LOGIC;
    SIGNAL S4523 : STD_LOGIC;
    SIGNAL S4524 : STD_LOGIC;
    SIGNAL S4525 : STD_LOGIC;
    SIGNAL S4526 : STD_LOGIC;
    SIGNAL S4527 : STD_LOGIC;
    SIGNAL S4528 : STD_LOGIC;
    SIGNAL S4529 : STD_LOGIC;
    SIGNAL S4530 : STD_LOGIC;
    SIGNAL S4531 : STD_LOGIC;
    SIGNAL S4532 : STD_LOGIC;
    SIGNAL S4533 : STD_LOGIC;
    SIGNAL S4534 : STD_LOGIC;
    SIGNAL S4535 : STD_LOGIC;
    SIGNAL S4536 : STD_LOGIC;
    SIGNAL S4537 : STD_LOGIC;
    SIGNAL S4538 : STD_LOGIC;
    SIGNAL S4539 : STD_LOGIC;
    SIGNAL S4540 : STD_LOGIC;
    SIGNAL S4541 : STD_LOGIC;
    SIGNAL S4542 : STD_LOGIC;
    SIGNAL S4543 : STD_LOGIC;
    SIGNAL S4544 : STD_LOGIC;
    SIGNAL S4545 : STD_LOGIC;
    SIGNAL S4546 : STD_LOGIC;
    SIGNAL S4547 : STD_LOGIC;
    SIGNAL S4548 : STD_LOGIC;
    SIGNAL S4549 : STD_LOGIC;
    SIGNAL S4550 : STD_LOGIC;
    SIGNAL S4551 : STD_LOGIC;
    SIGNAL S4552 : STD_LOGIC;
    SIGNAL S4553 : STD_LOGIC;
    SIGNAL S4554 : STD_LOGIC;
    SIGNAL S4555 : STD_LOGIC;
    SIGNAL S4556 : STD_LOGIC;
    SIGNAL S4557 : STD_LOGIC;
    SIGNAL S4558 : STD_LOGIC;
    SIGNAL S4559 : STD_LOGIC;
    SIGNAL S4560 : STD_LOGIC;
    SIGNAL S4561 : STD_LOGIC;
    SIGNAL S4562 : STD_LOGIC;
    SIGNAL S4563 : STD_LOGIC;
    SIGNAL S4564 : STD_LOGIC;
    SIGNAL S4565 : STD_LOGIC;
    SIGNAL S4566 : STD_LOGIC;
    SIGNAL S4567 : STD_LOGIC;
    SIGNAL S4568 : STD_LOGIC;
    SIGNAL S4569 : STD_LOGIC;
    SIGNAL S4570 : STD_LOGIC;
    SIGNAL S4571 : STD_LOGIC;
    SIGNAL S4572 : STD_LOGIC;
    SIGNAL S4573 : STD_LOGIC;
    SIGNAL S4574 : STD_LOGIC;
    SIGNAL S4575 : STD_LOGIC;
    SIGNAL S4576 : STD_LOGIC;
    SIGNAL S4577 : STD_LOGIC;
    SIGNAL S4578 : STD_LOGIC;
    SIGNAL S4579 : STD_LOGIC;
    SIGNAL S4580 : STD_LOGIC;
    SIGNAL S4581 : STD_LOGIC;
    SIGNAL S4582 : STD_LOGIC;
    SIGNAL S4583 : STD_LOGIC;
    SIGNAL S4584 : STD_LOGIC;
    SIGNAL S4585 : STD_LOGIC;
    SIGNAL S4586 : STD_LOGIC;
    SIGNAL S4587 : STD_LOGIC;
    SIGNAL S4588 : STD_LOGIC;
    SIGNAL S4589 : STD_LOGIC;
    SIGNAL S4590 : STD_LOGIC;
    SIGNAL S4591 : STD_LOGIC;
    SIGNAL S4592 : STD_LOGIC;
    SIGNAL S4593 : STD_LOGIC;
    SIGNAL S4594 : STD_LOGIC;
    SIGNAL S4595 : STD_LOGIC;
    SIGNAL S4596 : STD_LOGIC;
    SIGNAL S4597 : STD_LOGIC;
    SIGNAL S4598 : STD_LOGIC;
    SIGNAL S4599 : STD_LOGIC;
    SIGNAL S4600 : STD_LOGIC;
    SIGNAL S4601 : STD_LOGIC;
    SIGNAL S4602 : STD_LOGIC;
    SIGNAL S4603 : STD_LOGIC;
    SIGNAL S4604 : STD_LOGIC;
    SIGNAL S4605 : STD_LOGIC;
    SIGNAL S4606 : STD_LOGIC;
    SIGNAL S4607 : STD_LOGIC;
    SIGNAL S4608 : STD_LOGIC;
    SIGNAL S4609 : STD_LOGIC;
    SIGNAL S4610 : STD_LOGIC;
    SIGNAL S4611 : STD_LOGIC;
    SIGNAL S4612 : STD_LOGIC;
    SIGNAL S4613 : STD_LOGIC;
    SIGNAL S4614 : STD_LOGIC;
    SIGNAL S4615 : STD_LOGIC;
    SIGNAL S4616 : STD_LOGIC;
    SIGNAL S4617 : STD_LOGIC;
    SIGNAL S4618 : STD_LOGIC;
    SIGNAL S4619 : STD_LOGIC;
    SIGNAL S4620 : STD_LOGIC;
    SIGNAL S4621 : STD_LOGIC;
    SIGNAL S4622 : STD_LOGIC;
    SIGNAL S4623 : STD_LOGIC;
    SIGNAL S4624 : STD_LOGIC;
    SIGNAL S4625 : STD_LOGIC;
    SIGNAL S4626 : STD_LOGIC;
    SIGNAL S4627 : STD_LOGIC;
    SIGNAL S4628 : STD_LOGIC;
    SIGNAL S4629 : STD_LOGIC;
    SIGNAL S4630 : STD_LOGIC;
    SIGNAL S4631 : STD_LOGIC;
    SIGNAL S4632 : STD_LOGIC;
    SIGNAL S4633 : STD_LOGIC;
    SIGNAL S4634 : STD_LOGIC;
    SIGNAL S4635 : STD_LOGIC;
    SIGNAL S4636 : STD_LOGIC;
    SIGNAL S4637 : STD_LOGIC;
    SIGNAL S4638 : STD_LOGIC;
    SIGNAL S4639 : STD_LOGIC;
    SIGNAL S4640 : STD_LOGIC;
    SIGNAL S4641 : STD_LOGIC;
    SIGNAL S4642 : STD_LOGIC;
    SIGNAL S4643 : STD_LOGIC;
    SIGNAL S4644 : STD_LOGIC;
    SIGNAL S4645 : STD_LOGIC;
    SIGNAL S4646 : STD_LOGIC;
    SIGNAL S4647 : STD_LOGIC;
    SIGNAL S4648 : STD_LOGIC;
    SIGNAL S4649 : STD_LOGIC;
    SIGNAL S4650 : STD_LOGIC;
    SIGNAL S4651 : STD_LOGIC;
    SIGNAL S4652 : STD_LOGIC;
    SIGNAL S4653 : STD_LOGIC;
    SIGNAL S4654 : STD_LOGIC;
    SIGNAL S4655 : STD_LOGIC;
    SIGNAL S4656 : STD_LOGIC;
    SIGNAL S4657 : STD_LOGIC;
    SIGNAL S4658 : STD_LOGIC;
    SIGNAL S4659 : STD_LOGIC;
    SIGNAL S4660 : STD_LOGIC;
    SIGNAL S4661 : STD_LOGIC;
    SIGNAL S4662 : STD_LOGIC;
    SIGNAL S4663 : STD_LOGIC;
    SIGNAL S4664 : STD_LOGIC;
    SIGNAL S4665 : STD_LOGIC;
    SIGNAL S4666 : STD_LOGIC;
    SIGNAL S4667 : STD_LOGIC;
    SIGNAL S4668 : STD_LOGIC;
    SIGNAL S4669 : STD_LOGIC;
    SIGNAL S4670 : STD_LOGIC;
    SIGNAL S4671 : STD_LOGIC;
    SIGNAL S4672 : STD_LOGIC;
    SIGNAL S4673 : STD_LOGIC;
    SIGNAL S4674 : STD_LOGIC;
    SIGNAL S4675 : STD_LOGIC;
    SIGNAL S4676 : STD_LOGIC;
    SIGNAL S4677 : STD_LOGIC;
    SIGNAL S4678 : STD_LOGIC;
    SIGNAL S4679 : STD_LOGIC;
    SIGNAL S4680 : STD_LOGIC;
    SIGNAL S4681 : STD_LOGIC;
    SIGNAL S4682 : STD_LOGIC;
    SIGNAL S4683 : STD_LOGIC;
    SIGNAL S4684 : STD_LOGIC;
    SIGNAL S4685 : STD_LOGIC;
    SIGNAL S4686 : STD_LOGIC;
    SIGNAL S4687 : STD_LOGIC;
    SIGNAL S4688 : STD_LOGIC;
    SIGNAL S4689 : STD_LOGIC;
    SIGNAL S4690 : STD_LOGIC;
    SIGNAL S4691 : STD_LOGIC;
    SIGNAL S4692 : STD_LOGIC;
    SIGNAL S4693 : STD_LOGIC;
    SIGNAL S4694 : STD_LOGIC;
    SIGNAL S4695 : STD_LOGIC;
    SIGNAL S4696 : STD_LOGIC;
    SIGNAL S4697 : STD_LOGIC;
    SIGNAL S4698 : STD_LOGIC;
    SIGNAL S4699 : STD_LOGIC;
    SIGNAL S4700 : STD_LOGIC;
    SIGNAL S4701 : STD_LOGIC;
    SIGNAL S4702 : STD_LOGIC;
    SIGNAL S4703 : STD_LOGIC;
    SIGNAL S4704 : STD_LOGIC;
    SIGNAL S4705 : STD_LOGIC;
    SIGNAL S4706 : STD_LOGIC;
    SIGNAL S4707 : STD_LOGIC;
    SIGNAL S4708 : STD_LOGIC;
    SIGNAL S4709 : STD_LOGIC;
    SIGNAL S4710 : STD_LOGIC;
    SIGNAL S4711 : STD_LOGIC;
    SIGNAL S4712 : STD_LOGIC;
    SIGNAL S4713 : STD_LOGIC;
    SIGNAL S4714 : STD_LOGIC;
    SIGNAL S4715 : STD_LOGIC;
    SIGNAL S4716 : STD_LOGIC;
    SIGNAL S4717 : STD_LOGIC;
    SIGNAL S4718 : STD_LOGIC;
    SIGNAL S4719 : STD_LOGIC;
    SIGNAL S4720 : STD_LOGIC;
    SIGNAL S4721 : STD_LOGIC;
    SIGNAL S4722 : STD_LOGIC;
    SIGNAL S4723 : STD_LOGIC;
    SIGNAL S4724 : STD_LOGIC;
    SIGNAL S4725 : STD_LOGIC;
    SIGNAL S4726 : STD_LOGIC;
    SIGNAL S4727 : STD_LOGIC;
    SIGNAL S4728 : STD_LOGIC;
    SIGNAL S4729 : STD_LOGIC;
    SIGNAL S4730 : STD_LOGIC;
    SIGNAL S4731 : STD_LOGIC;
    SIGNAL S4732 : STD_LOGIC;
    SIGNAL S4733 : STD_LOGIC;
    SIGNAL S4734 : STD_LOGIC;
    SIGNAL S4735 : STD_LOGIC;
    SIGNAL S4736 : STD_LOGIC;
    SIGNAL S4737 : STD_LOGIC;
    SIGNAL S4738 : STD_LOGIC;
    SIGNAL S4739 : STD_LOGIC;
    SIGNAL S4740 : STD_LOGIC;
    SIGNAL S4741 : STD_LOGIC;
    SIGNAL S4742 : STD_LOGIC;
    SIGNAL S4743 : STD_LOGIC;
    SIGNAL S4744 : STD_LOGIC;
    SIGNAL S4745 : STD_LOGIC;
    SIGNAL S4746 : STD_LOGIC;
    SIGNAL S4747 : STD_LOGIC;
    SIGNAL S4748 : STD_LOGIC;
    SIGNAL S4749 : STD_LOGIC;
    SIGNAL S4750 : STD_LOGIC;
    SIGNAL S4751 : STD_LOGIC;
    SIGNAL S4752 : STD_LOGIC;
    SIGNAL S4753 : STD_LOGIC;
    SIGNAL S4754 : STD_LOGIC;
    SIGNAL S4755 : STD_LOGIC;
    SIGNAL S4756 : STD_LOGIC;
    SIGNAL S4757 : STD_LOGIC;
    SIGNAL S4758 : STD_LOGIC;
    SIGNAL S4759 : STD_LOGIC;
    SIGNAL S4760 : STD_LOGIC;
    SIGNAL S4761 : STD_LOGIC;
    SIGNAL S4762 : STD_LOGIC;
    SIGNAL S4763 : STD_LOGIC;
    SIGNAL S4764 : STD_LOGIC;
    SIGNAL S4765 : STD_LOGIC;
    SIGNAL S4766 : STD_LOGIC;
    SIGNAL S4767 : STD_LOGIC;
    SIGNAL S4768 : STD_LOGIC;
    SIGNAL S4769 : STD_LOGIC;
    SIGNAL S4770 : STD_LOGIC;
    SIGNAL S4771 : STD_LOGIC;
    SIGNAL S4772 : STD_LOGIC;
    SIGNAL S4773 : STD_LOGIC;
    SIGNAL S4774 : STD_LOGIC;
    SIGNAL S4775 : STD_LOGIC;
    SIGNAL S4776 : STD_LOGIC;
    SIGNAL S4777 : STD_LOGIC;
    SIGNAL S4778 : STD_LOGIC;
    SIGNAL S4779 : STD_LOGIC;
    SIGNAL S4780 : STD_LOGIC;
    SIGNAL S4781 : STD_LOGIC;
    SIGNAL S4782 : STD_LOGIC;
    SIGNAL S4783 : STD_LOGIC;
    SIGNAL S4784 : STD_LOGIC;
    SIGNAL S4785 : STD_LOGIC;
    SIGNAL S4786 : STD_LOGIC;
    SIGNAL S4787 : STD_LOGIC;
    SIGNAL S4788 : STD_LOGIC;
    SIGNAL S4789 : STD_LOGIC;
    SIGNAL S4790 : STD_LOGIC;
    SIGNAL S4791 : STD_LOGIC;
    SIGNAL S4792 : STD_LOGIC;
    SIGNAL S4793 : STD_LOGIC;
    SIGNAL S4794 : STD_LOGIC;
    SIGNAL S4795 : STD_LOGIC;
    SIGNAL S4796 : STD_LOGIC;
    SIGNAL S4797 : STD_LOGIC;
    SIGNAL S4798 : STD_LOGIC;
    SIGNAL S4799 : STD_LOGIC;
    SIGNAL S4800 : STD_LOGIC;
    SIGNAL S4801 : STD_LOGIC;
    SIGNAL S4802 : STD_LOGIC;
    SIGNAL S4803 : STD_LOGIC;
    SIGNAL S4804 : STD_LOGIC;
    SIGNAL S4805 : STD_LOGIC;
    SIGNAL S4806 : STD_LOGIC;
    SIGNAL S4807 : STD_LOGIC;
    SIGNAL S4808 : STD_LOGIC;
    SIGNAL S4809 : STD_LOGIC;
    SIGNAL S4810 : STD_LOGIC;
    SIGNAL S4811 : STD_LOGIC;
    SIGNAL S4812 : STD_LOGIC;
    SIGNAL S4813 : STD_LOGIC;
    SIGNAL S4814 : STD_LOGIC;
    SIGNAL S4815 : STD_LOGIC;
    SIGNAL S4816 : STD_LOGIC;
    SIGNAL S4817 : STD_LOGIC;
    SIGNAL S4818 : STD_LOGIC;
    SIGNAL S4819 : STD_LOGIC;
    SIGNAL S4820 : STD_LOGIC;
    SIGNAL S4821 : STD_LOGIC;
    SIGNAL S4822 : STD_LOGIC;
    SIGNAL S4823 : STD_LOGIC;
    SIGNAL S4824 : STD_LOGIC;
    SIGNAL S4825 : STD_LOGIC;
    SIGNAL S4826 : STD_LOGIC;
    SIGNAL S4827 : STD_LOGIC;
    SIGNAL S4828 : STD_LOGIC;
    SIGNAL S4829 : STD_LOGIC;
    SIGNAL S4830 : STD_LOGIC;
    SIGNAL S4831 : STD_LOGIC;
    SIGNAL S4832 : STD_LOGIC;
    SIGNAL S4833 : STD_LOGIC;
    SIGNAL S4834 : STD_LOGIC;
    SIGNAL S4835 : STD_LOGIC;
    SIGNAL S4836 : STD_LOGIC;
    SIGNAL S4837 : STD_LOGIC;
    SIGNAL S4838 : STD_LOGIC;
    SIGNAL S4839 : STD_LOGIC;
    SIGNAL S4840 : STD_LOGIC;
    SIGNAL S4841 : STD_LOGIC;
    SIGNAL S4842 : STD_LOGIC;
    SIGNAL S4843 : STD_LOGIC;
    SIGNAL S4844 : STD_LOGIC;
    SIGNAL S4845 : STD_LOGIC;
    SIGNAL S4846 : STD_LOGIC;
    SIGNAL S4847 : STD_LOGIC;
    SIGNAL S4848 : STD_LOGIC;
    SIGNAL S4849 : STD_LOGIC;
    SIGNAL S4850 : STD_LOGIC;
    SIGNAL S4851 : STD_LOGIC;
    SIGNAL S4852 : STD_LOGIC;
    SIGNAL S4853 : STD_LOGIC;
    SIGNAL S4854 : STD_LOGIC;
    SIGNAL S4855 : STD_LOGIC;
    SIGNAL S4856 : STD_LOGIC;
    SIGNAL S4857 : STD_LOGIC;
    SIGNAL S4858 : STD_LOGIC;
    SIGNAL S4859 : STD_LOGIC;
    SIGNAL S4860 : STD_LOGIC;
    SIGNAL S4861 : STD_LOGIC;
    SIGNAL S4862 : STD_LOGIC;
    SIGNAL S4863 : STD_LOGIC;
    SIGNAL S4864 : STD_LOGIC;
    SIGNAL S4865 : STD_LOGIC;
    SIGNAL S4866 : STD_LOGIC;
    SIGNAL S4867 : STD_LOGIC;
    SIGNAL S4868 : STD_LOGIC;
    SIGNAL S4869 : STD_LOGIC;
    SIGNAL S4870 : STD_LOGIC;
    SIGNAL S4871 : STD_LOGIC;
    SIGNAL S4872 : STD_LOGIC;
    SIGNAL S4873 : STD_LOGIC;
    SIGNAL S4874 : STD_LOGIC;
    SIGNAL S4875 : STD_LOGIC;
    SIGNAL S4876 : STD_LOGIC;
    SIGNAL S4877 : STD_LOGIC;
    SIGNAL S4878 : STD_LOGIC;
    SIGNAL S4879 : STD_LOGIC;
    SIGNAL S4880 : STD_LOGIC;
    SIGNAL S4881 : STD_LOGIC;
    SIGNAL S4882 : STD_LOGIC;
    SIGNAL S4883 : STD_LOGIC;
    SIGNAL S4884 : STD_LOGIC;
    SIGNAL S4885 : STD_LOGIC;
    SIGNAL S4886 : STD_LOGIC;
    SIGNAL S4887 : STD_LOGIC;
    SIGNAL S4888 : STD_LOGIC;
    SIGNAL S4889 : STD_LOGIC;
    SIGNAL S4890 : STD_LOGIC;
    SIGNAL S4891 : STD_LOGIC;
    SIGNAL S4892 : STD_LOGIC;
    SIGNAL S4893 : STD_LOGIC;
    SIGNAL S4894 : STD_LOGIC;
    SIGNAL S4895 : STD_LOGIC;
    SIGNAL S4896 : STD_LOGIC;
    SIGNAL S4897 : STD_LOGIC;
    SIGNAL S4898 : STD_LOGIC;
    SIGNAL S4899 : STD_LOGIC;
    SIGNAL S4900 : STD_LOGIC;
    SIGNAL S4901 : STD_LOGIC;
    SIGNAL S4902 : STD_LOGIC;
    SIGNAL S4903 : STD_LOGIC;
    SIGNAL S4904 : STD_LOGIC;
    SIGNAL S4905 : STD_LOGIC;
    SIGNAL S4906 : STD_LOGIC;
    SIGNAL S4907 : STD_LOGIC;
    SIGNAL S4908 : STD_LOGIC;
    SIGNAL S4909 : STD_LOGIC;
    SIGNAL S4910 : STD_LOGIC;
    SIGNAL S4911 : STD_LOGIC;
    SIGNAL S4912 : STD_LOGIC;
    SIGNAL S4913 : STD_LOGIC;
    SIGNAL S4914 : STD_LOGIC;
    SIGNAL S4915 : STD_LOGIC;
    SIGNAL S4916 : STD_LOGIC;
    SIGNAL S4917 : STD_LOGIC;
    SIGNAL S4918 : STD_LOGIC;
    SIGNAL S4919 : STD_LOGIC;
    SIGNAL S4920 : STD_LOGIC;
    SIGNAL S4921 : STD_LOGIC;
    SIGNAL S4922 : STD_LOGIC;
    SIGNAL S4923 : STD_LOGIC;
    SIGNAL S4924 : STD_LOGIC;
    SIGNAL S4925 : STD_LOGIC;
    SIGNAL S4926 : STD_LOGIC;
    SIGNAL S4927 : STD_LOGIC;
    SIGNAL S4928 : STD_LOGIC;
    SIGNAL S4929 : STD_LOGIC;
    SIGNAL S4930 : STD_LOGIC;
    SIGNAL S4931 : STD_LOGIC;
    SIGNAL S4932 : STD_LOGIC;
    SIGNAL S4933 : STD_LOGIC;
    SIGNAL S4934 : STD_LOGIC;
    SIGNAL S4935 : STD_LOGIC;
    SIGNAL S4936 : STD_LOGIC;
    SIGNAL S4937 : STD_LOGIC;
    SIGNAL S4938 : STD_LOGIC;
    SIGNAL S4939 : STD_LOGIC;
    SIGNAL S4940 : STD_LOGIC;
    SIGNAL S4941 : STD_LOGIC;
    SIGNAL S4942 : STD_LOGIC;
    SIGNAL S4943 : STD_LOGIC;
    SIGNAL S4944 : STD_LOGIC;
    SIGNAL S4945 : STD_LOGIC;
    SIGNAL S4946 : STD_LOGIC;
    SIGNAL S4947 : STD_LOGIC;
    SIGNAL S4948 : STD_LOGIC;
    SIGNAL S4949 : STD_LOGIC;
    SIGNAL S4950 : STD_LOGIC;
    SIGNAL S4951 : STD_LOGIC;
    SIGNAL S4952 : STD_LOGIC;
    SIGNAL S4953 : STD_LOGIC;
    SIGNAL S4954 : STD_LOGIC;
    SIGNAL S4955 : STD_LOGIC;
    SIGNAL S4956 : STD_LOGIC;
    SIGNAL S4957 : STD_LOGIC;
    SIGNAL S4958 : STD_LOGIC;
    SIGNAL S4959 : STD_LOGIC;
    SIGNAL S4960 : STD_LOGIC;
    SIGNAL S4961 : STD_LOGIC;
    SIGNAL S4962 : STD_LOGIC;
    SIGNAL S4963 : STD_LOGIC;
    SIGNAL S4964 : STD_LOGIC;
    SIGNAL S4965 : STD_LOGIC;
    SIGNAL S4966 : STD_LOGIC;
    SIGNAL S4967 : STD_LOGIC;
    SIGNAL S4968 : STD_LOGIC;
    SIGNAL S4969 : STD_LOGIC;
    SIGNAL S4970 : STD_LOGIC;
    SIGNAL S4971 : STD_LOGIC;
    SIGNAL S4972 : STD_LOGIC;
    SIGNAL S4973 : STD_LOGIC;
    SIGNAL S4974 : STD_LOGIC;
    SIGNAL S4975 : STD_LOGIC;
    SIGNAL S4976 : STD_LOGIC;
    SIGNAL S4977 : STD_LOGIC;
    SIGNAL S4978 : STD_LOGIC;
    SIGNAL S4979 : STD_LOGIC;
    SIGNAL S4980 : STD_LOGIC;
    SIGNAL S4981 : STD_LOGIC;
    SIGNAL S4982 : STD_LOGIC;
    SIGNAL S4983 : STD_LOGIC;
    SIGNAL S4984 : STD_LOGIC;
    SIGNAL S4985 : STD_LOGIC;
    SIGNAL S4986 : STD_LOGIC;
    SIGNAL S4987 : STD_LOGIC;
    SIGNAL S4988 : STD_LOGIC;
    SIGNAL S4989 : STD_LOGIC;
    SIGNAL S4990 : STD_LOGIC;
    SIGNAL S4991 : STD_LOGIC;
    SIGNAL S4992 : STD_LOGIC;
    SIGNAL S4993 : STD_LOGIC;
    SIGNAL S4994 : STD_LOGIC;
    SIGNAL S4995 : STD_LOGIC;
    SIGNAL S4996 : STD_LOGIC;
    SIGNAL S4997 : STD_LOGIC;
    SIGNAL S4998 : STD_LOGIC;
    SIGNAL S4999 : STD_LOGIC;
    SIGNAL S5000 : STD_LOGIC;
    SIGNAL S5001 : STD_LOGIC;
    SIGNAL S5002 : STD_LOGIC;
    SIGNAL S5003 : STD_LOGIC;
    SIGNAL S5004 : STD_LOGIC;
    SIGNAL S5005 : STD_LOGIC;
    SIGNAL S5006 : STD_LOGIC;
    SIGNAL S5007 : STD_LOGIC;
    SIGNAL S5008 : STD_LOGIC;
    SIGNAL S5009 : STD_LOGIC;
    SIGNAL S5010 : STD_LOGIC;
    SIGNAL S5011 : STD_LOGIC;
    SIGNAL S5012 : STD_LOGIC;
    SIGNAL S5013 : STD_LOGIC;
    SIGNAL S5014 : STD_LOGIC;
    SIGNAL S5015 : STD_LOGIC;
    SIGNAL S5016 : STD_LOGIC;
    SIGNAL S5017 : STD_LOGIC;
    SIGNAL S5018 : STD_LOGIC;
    SIGNAL S5019 : STD_LOGIC;
    SIGNAL S5020 : STD_LOGIC;
    SIGNAL S5021 : STD_LOGIC;
    SIGNAL S5022 : STD_LOGIC;
    SIGNAL S5023 : STD_LOGIC;
    SIGNAL S5024 : STD_LOGIC;
    SIGNAL S5025 : STD_LOGIC;
    SIGNAL S5026 : STD_LOGIC;
    SIGNAL S5027 : STD_LOGIC;
    SIGNAL S5028 : STD_LOGIC;
    SIGNAL S5029 : STD_LOGIC;
    SIGNAL S5030 : STD_LOGIC;
    SIGNAL S5031 : STD_LOGIC;
    SIGNAL S5032 : STD_LOGIC;
    SIGNAL S5033 : STD_LOGIC;
    SIGNAL S5034 : STD_LOGIC;
    SIGNAL S5035 : STD_LOGIC;
    SIGNAL S5036 : STD_LOGIC;
    SIGNAL S5037 : STD_LOGIC;
    SIGNAL S5038 : STD_LOGIC;
    SIGNAL S5039 : STD_LOGIC;
    SIGNAL S5040 : STD_LOGIC;
    SIGNAL S5041 : STD_LOGIC;
    SIGNAL S5042 : STD_LOGIC;
    SIGNAL S5043 : STD_LOGIC;
    SIGNAL S5044 : STD_LOGIC;
    SIGNAL S5045 : STD_LOGIC;
    SIGNAL S5046 : STD_LOGIC;
    SIGNAL S5047 : STD_LOGIC;
    SIGNAL S5048 : STD_LOGIC;
    SIGNAL S5049 : STD_LOGIC;
    SIGNAL S5050 : STD_LOGIC;
    SIGNAL S5051 : STD_LOGIC;
    SIGNAL S5052 : STD_LOGIC;
    SIGNAL S5053 : STD_LOGIC;
    SIGNAL S5054 : STD_LOGIC;
    SIGNAL S5055 : STD_LOGIC;
    SIGNAL S5056 : STD_LOGIC;
    SIGNAL S5057 : STD_LOGIC;
    SIGNAL S5058 : STD_LOGIC;
    SIGNAL S5059 : STD_LOGIC;
    SIGNAL S5060 : STD_LOGIC;
    SIGNAL S5061 : STD_LOGIC;
    SIGNAL S5062 : STD_LOGIC;
    SIGNAL S5063 : STD_LOGIC;
    SIGNAL S5064 : STD_LOGIC;
    SIGNAL S5065 : STD_LOGIC;
    SIGNAL S5066 : STD_LOGIC;
    SIGNAL S5067 : STD_LOGIC;
    SIGNAL S5068 : STD_LOGIC;
    SIGNAL S5069 : STD_LOGIC;
    SIGNAL S5070 : STD_LOGIC;
    SIGNAL S5071 : STD_LOGIC;
    SIGNAL S5072 : STD_LOGIC;
    SIGNAL S5073 : STD_LOGIC;
    SIGNAL S5074 : STD_LOGIC;
    SIGNAL S5075 : STD_LOGIC;
    SIGNAL S5076 : STD_LOGIC;
    SIGNAL S5077 : STD_LOGIC;
    SIGNAL S5078 : STD_LOGIC;
    SIGNAL S5079 : STD_LOGIC;
    SIGNAL S5080 : STD_LOGIC;
    SIGNAL S5081 : STD_LOGIC;
    SIGNAL S5082 : STD_LOGIC;
    SIGNAL S5083 : STD_LOGIC;
    SIGNAL S5084 : STD_LOGIC;
    SIGNAL S5085 : STD_LOGIC;
    SIGNAL S5086 : STD_LOGIC;
    SIGNAL S5087 : STD_LOGIC;
    SIGNAL S5088 : STD_LOGIC;
    SIGNAL S5089 : STD_LOGIC;
    SIGNAL S5090 : STD_LOGIC;
    SIGNAL S5091 : STD_LOGIC;
    SIGNAL S5092 : STD_LOGIC;
    SIGNAL S5093 : STD_LOGIC;
    SIGNAL S5094 : STD_LOGIC;
    SIGNAL S5095 : STD_LOGIC;
    SIGNAL S5096 : STD_LOGIC;
    SIGNAL S5097 : STD_LOGIC;
    SIGNAL S5098 : STD_LOGIC;
    SIGNAL S5099 : STD_LOGIC;
    SIGNAL S5100 : STD_LOGIC;
    SIGNAL S5101 : STD_LOGIC;
    SIGNAL S5102 : STD_LOGIC;
    SIGNAL S5103 : STD_LOGIC;
    SIGNAL S5104 : STD_LOGIC;
    SIGNAL S5105 : STD_LOGIC;
    SIGNAL S5106 : STD_LOGIC;
    SIGNAL S5107 : STD_LOGIC;
    SIGNAL S5108 : STD_LOGIC;
    SIGNAL S5109 : STD_LOGIC;
    SIGNAL S5110 : STD_LOGIC;
    SIGNAL S5111 : STD_LOGIC;
    SIGNAL S5112 : STD_LOGIC;
    SIGNAL S5113 : STD_LOGIC;
    SIGNAL S5114 : STD_LOGIC;
    SIGNAL S5115 : STD_LOGIC;
    SIGNAL S5116 : STD_LOGIC;
    SIGNAL S5117 : STD_LOGIC;
    SIGNAL S5118 : STD_LOGIC;
    SIGNAL S5119 : STD_LOGIC;
    SIGNAL S5120 : STD_LOGIC;
    SIGNAL S5121 : STD_LOGIC;
    SIGNAL S5122 : STD_LOGIC;
    SIGNAL S5123 : STD_LOGIC;
    SIGNAL S5124 : STD_LOGIC;
    SIGNAL S5125 : STD_LOGIC;
    SIGNAL S5126 : STD_LOGIC;
    SIGNAL S5127 : STD_LOGIC;
    SIGNAL S5128 : STD_LOGIC;
    SIGNAL S5129 : STD_LOGIC;
    SIGNAL S5130 : STD_LOGIC;
    SIGNAL S5131 : STD_LOGIC;
    SIGNAL S5132 : STD_LOGIC;
    SIGNAL S5133 : STD_LOGIC;
    SIGNAL S5134 : STD_LOGIC;
    SIGNAL S5135 : STD_LOGIC;
    SIGNAL S5136 : STD_LOGIC;
    SIGNAL S5137 : STD_LOGIC;
    SIGNAL S5138 : STD_LOGIC;
    SIGNAL S5139 : STD_LOGIC;
    SIGNAL S5140 : STD_LOGIC;
    SIGNAL S5141 : STD_LOGIC;
    SIGNAL S5142 : STD_LOGIC;
    SIGNAL S5143 : STD_LOGIC;
    SIGNAL S5144 : STD_LOGIC;
    SIGNAL S5145 : STD_LOGIC;
    SIGNAL S5146 : STD_LOGIC;
    SIGNAL S5147 : STD_LOGIC;
    SIGNAL S5148 : STD_LOGIC;
    SIGNAL S5149 : STD_LOGIC;
    SIGNAL S5150 : STD_LOGIC;
    SIGNAL S5151 : STD_LOGIC;
    SIGNAL S5152 : STD_LOGIC;
    SIGNAL S5153 : STD_LOGIC;
    SIGNAL S5154 : STD_LOGIC;
    SIGNAL S5155 : STD_LOGIC;
    SIGNAL S5156 : STD_LOGIC;
    SIGNAL S5157 : STD_LOGIC;
    SIGNAL S5158 : STD_LOGIC;
    SIGNAL S5159 : STD_LOGIC;
    SIGNAL S5160 : STD_LOGIC;
    SIGNAL S5161 : STD_LOGIC;
    SIGNAL S5162 : STD_LOGIC;
    SIGNAL S5163 : STD_LOGIC;
    SIGNAL S5164 : STD_LOGIC;
    SIGNAL S5165 : STD_LOGIC;
    SIGNAL S5166 : STD_LOGIC;
    SIGNAL S5167 : STD_LOGIC;
    SIGNAL S5168 : STD_LOGIC;
    SIGNAL S5169 : STD_LOGIC;
    SIGNAL S5170 : STD_LOGIC;
    SIGNAL S5171 : STD_LOGIC;
    SIGNAL S5172 : STD_LOGIC;
    SIGNAL S5173 : STD_LOGIC;
    SIGNAL S5174 : STD_LOGIC;
    SIGNAL S5175 : STD_LOGIC;
    SIGNAL S5176 : STD_LOGIC;
    SIGNAL S5177 : STD_LOGIC;
    SIGNAL S5178 : STD_LOGIC;
    SIGNAL S5179 : STD_LOGIC;
    SIGNAL S5180 : STD_LOGIC;
    SIGNAL S5181 : STD_LOGIC;
    SIGNAL S5182 : STD_LOGIC;
    SIGNAL S5183 : STD_LOGIC;
    SIGNAL S5184 : STD_LOGIC;
    SIGNAL S5185 : STD_LOGIC;
    SIGNAL S5186 : STD_LOGIC;
    SIGNAL S5187 : STD_LOGIC;
    SIGNAL S5188 : STD_LOGIC;
    SIGNAL S5189 : STD_LOGIC;
    SIGNAL S5190 : STD_LOGIC;
    SIGNAL S5191 : STD_LOGIC;
    SIGNAL S5192 : STD_LOGIC;
    SIGNAL S5193 : STD_LOGIC;
    SIGNAL S5194 : STD_LOGIC;
    SIGNAL S5195 : STD_LOGIC;
    SIGNAL S5196 : STD_LOGIC;
    SIGNAL S5197 : STD_LOGIC;
    SIGNAL S5198 : STD_LOGIC;
    SIGNAL S5199 : STD_LOGIC;
    SIGNAL S5200 : STD_LOGIC;
    SIGNAL S5201 : STD_LOGIC;
    SIGNAL S5202 : STD_LOGIC;
    SIGNAL S5203 : STD_LOGIC;
    SIGNAL S5204 : STD_LOGIC;
    SIGNAL S5205 : STD_LOGIC;
    SIGNAL S5206 : STD_LOGIC;
    SIGNAL S5207 : STD_LOGIC;
    SIGNAL S5208 : STD_LOGIC;
    SIGNAL S5209 : STD_LOGIC;
    SIGNAL S5210 : STD_LOGIC;
    SIGNAL S5211 : STD_LOGIC;
    SIGNAL S5212 : STD_LOGIC;
    SIGNAL S5213 : STD_LOGIC;
    SIGNAL S5214 : STD_LOGIC;
    SIGNAL S5215 : STD_LOGIC;
    SIGNAL S5216 : STD_LOGIC;
    SIGNAL S5217 : STD_LOGIC;
    SIGNAL S5218 : STD_LOGIC;
    SIGNAL S5219 : STD_LOGIC;
    SIGNAL S5220 : STD_LOGIC;
    SIGNAL S5221 : STD_LOGIC;
    SIGNAL S5222 : STD_LOGIC;
    SIGNAL S5223 : STD_LOGIC;
    SIGNAL S5224 : STD_LOGIC;
    SIGNAL S5225 : STD_LOGIC;
    SIGNAL S5226 : STD_LOGIC;
    SIGNAL S5227 : STD_LOGIC;
    SIGNAL S5228 : STD_LOGIC;
    SIGNAL S5229 : STD_LOGIC;
    SIGNAL S5230 : STD_LOGIC;
    SIGNAL S5231 : STD_LOGIC;
    SIGNAL S5232 : STD_LOGIC;
    SIGNAL S5233 : STD_LOGIC;
    SIGNAL S5234 : STD_LOGIC;
    SIGNAL S5235 : STD_LOGIC;
    SIGNAL S5236 : STD_LOGIC;
    SIGNAL S5237 : STD_LOGIC;
    SIGNAL S5238 : STD_LOGIC;
    SIGNAL S5239 : STD_LOGIC;
    SIGNAL S5240 : STD_LOGIC;
    SIGNAL S5241 : STD_LOGIC;
    SIGNAL S5242 : STD_LOGIC;
    SIGNAL S5243 : STD_LOGIC;
    SIGNAL S5244 : STD_LOGIC;
    SIGNAL S5245 : STD_LOGIC;
    SIGNAL S5246 : STD_LOGIC;
    SIGNAL S5247 : STD_LOGIC;
    SIGNAL S5248 : STD_LOGIC;
    SIGNAL S5249 : STD_LOGIC;
    SIGNAL S5250 : STD_LOGIC;
    SIGNAL S5251 : STD_LOGIC;
    SIGNAL S5252 : STD_LOGIC;
    SIGNAL S5253 : STD_LOGIC;
    SIGNAL S5254 : STD_LOGIC;
    SIGNAL S5255 : STD_LOGIC;
    SIGNAL S5256 : STD_LOGIC;
    SIGNAL S5257 : STD_LOGIC;
    SIGNAL S5258 : STD_LOGIC;
    SIGNAL S5259 : STD_LOGIC;
    SIGNAL S5260 : STD_LOGIC;
    SIGNAL S5261 : STD_LOGIC;
    SIGNAL S5262 : STD_LOGIC;
    SIGNAL S5263 : STD_LOGIC;
    SIGNAL S5264 : STD_LOGIC;
    SIGNAL S5265 : STD_LOGIC;
    SIGNAL S5266 : STD_LOGIC;
    SIGNAL S5267 : STD_LOGIC;
    SIGNAL S5268 : STD_LOGIC;
    SIGNAL S5269 : STD_LOGIC;
    SIGNAL S5270 : STD_LOGIC;
    SIGNAL S5271 : STD_LOGIC;
    SIGNAL S5272 : STD_LOGIC;
    SIGNAL S5273 : STD_LOGIC;
    SIGNAL S5274 : STD_LOGIC;
    SIGNAL S5275 : STD_LOGIC;
    SIGNAL S5276 : STD_LOGIC;
    SIGNAL S5277 : STD_LOGIC;
    SIGNAL S5278 : STD_LOGIC;
    SIGNAL S5279 : STD_LOGIC;
    SIGNAL S5280 : STD_LOGIC;
    SIGNAL S5281 : STD_LOGIC;
    SIGNAL S5282 : STD_LOGIC;
    SIGNAL S5283 : STD_LOGIC;
    SIGNAL S5284 : STD_LOGIC;
    SIGNAL S5285 : STD_LOGIC;
    SIGNAL S5286 : STD_LOGIC;
    SIGNAL S5287 : STD_LOGIC;
    SIGNAL S5288 : STD_LOGIC;
    SIGNAL S5289 : STD_LOGIC;
    SIGNAL S5290 : STD_LOGIC;
    SIGNAL S5291 : STD_LOGIC;
    SIGNAL S5292 : STD_LOGIC;
    SIGNAL S5293 : STD_LOGIC;
    SIGNAL S5294 : STD_LOGIC;
    SIGNAL S5295 : STD_LOGIC;
    SIGNAL S5296 : STD_LOGIC;
    SIGNAL S5297 : STD_LOGIC;
    SIGNAL S5298 : STD_LOGIC;
    SIGNAL S5299 : STD_LOGIC;
    SIGNAL S5300 : STD_LOGIC;
    SIGNAL S5301 : STD_LOGIC;
    SIGNAL S5302 : STD_LOGIC;
    SIGNAL S5303 : STD_LOGIC;
    SIGNAL S5304 : STD_LOGIC;
    SIGNAL S5305 : STD_LOGIC;
    SIGNAL S5306 : STD_LOGIC;
    SIGNAL S5307 : STD_LOGIC;
    SIGNAL S5308 : STD_LOGIC;
    SIGNAL S5309 : STD_LOGIC;
    SIGNAL S5310 : STD_LOGIC;
    SIGNAL S5311 : STD_LOGIC;
    SIGNAL S5312 : STD_LOGIC;
    SIGNAL S5313 : STD_LOGIC;
    SIGNAL S5314 : STD_LOGIC;
    SIGNAL S5315 : STD_LOGIC;
    SIGNAL S5316 : STD_LOGIC;
    SIGNAL S5317 : STD_LOGIC;
    SIGNAL S5318 : STD_LOGIC;
    SIGNAL S5319 : STD_LOGIC;
    SIGNAL S5320 : STD_LOGIC;
    SIGNAL S5321 : STD_LOGIC;
    SIGNAL S5322 : STD_LOGIC;
    SIGNAL S5323 : STD_LOGIC;
    SIGNAL S5324 : STD_LOGIC;
    SIGNAL S5325 : STD_LOGIC;
    SIGNAL S5326 : STD_LOGIC;
    SIGNAL S5327 : STD_LOGIC;
    SIGNAL S5328 : STD_LOGIC;
    SIGNAL S5329 : STD_LOGIC;
    SIGNAL S5330 : STD_LOGIC;
    SIGNAL S5331 : STD_LOGIC;
    SIGNAL S5332 : STD_LOGIC;
    SIGNAL S5333 : STD_LOGIC;
    SIGNAL S5334 : STD_LOGIC;
    SIGNAL S5335 : STD_LOGIC;
    SIGNAL S5336 : STD_LOGIC;
    SIGNAL S5337 : STD_LOGIC;
    SIGNAL S5338 : STD_LOGIC;
    SIGNAL S5339 : STD_LOGIC;
    SIGNAL S5340 : STD_LOGIC;
    SIGNAL S5341 : STD_LOGIC;
    SIGNAL S5342 : STD_LOGIC;
    SIGNAL S5343 : STD_LOGIC;
    SIGNAL S5344 : STD_LOGIC;
    SIGNAL S5345 : STD_LOGIC;
    SIGNAL S5346 : STD_LOGIC;
    SIGNAL S5347 : STD_LOGIC;
    SIGNAL S5348 : STD_LOGIC;
    SIGNAL S5349 : STD_LOGIC;
    SIGNAL S5350 : STD_LOGIC;
    SIGNAL S5351 : STD_LOGIC;
    SIGNAL S5352 : STD_LOGIC;
    SIGNAL S5353 : STD_LOGIC;
    SIGNAL S5354 : STD_LOGIC;
    SIGNAL S5355 : STD_LOGIC;
    SIGNAL S5356 : STD_LOGIC;
    SIGNAL S5357 : STD_LOGIC;
    SIGNAL S5358 : STD_LOGIC;
    SIGNAL S5359 : STD_LOGIC;
    SIGNAL S5360 : STD_LOGIC;
    SIGNAL S5361 : STD_LOGIC;
    SIGNAL S5362 : STD_LOGIC;
    SIGNAL S5363 : STD_LOGIC;
    SIGNAL S5364 : STD_LOGIC;
    SIGNAL S5365 : STD_LOGIC;
    SIGNAL S5366 : STD_LOGIC;
    SIGNAL S5367 : STD_LOGIC;
    SIGNAL S5368 : STD_LOGIC;
    SIGNAL S5369 : STD_LOGIC;
    SIGNAL S5370 : STD_LOGIC;
    SIGNAL S5371 : STD_LOGIC;
    SIGNAL S5372 : STD_LOGIC;
    SIGNAL S5373 : STD_LOGIC;
    SIGNAL S5374 : STD_LOGIC;
    SIGNAL S5375 : STD_LOGIC;
    SIGNAL S5376 : STD_LOGIC;
    SIGNAL S5377 : STD_LOGIC;
    SIGNAL S5378 : STD_LOGIC;
    SIGNAL S5379 : STD_LOGIC;
    SIGNAL S5380 : STD_LOGIC;
    SIGNAL S5381 : STD_LOGIC;
    SIGNAL S5382 : STD_LOGIC;
    SIGNAL S5383 : STD_LOGIC;
    SIGNAL S5384 : STD_LOGIC;
    SIGNAL S5385 : STD_LOGIC;
    SIGNAL S5386 : STD_LOGIC;
    SIGNAL S5387 : STD_LOGIC;
    SIGNAL S5388 : STD_LOGIC;
    SIGNAL S5389 : STD_LOGIC;
    SIGNAL S5390 : STD_LOGIC;
    SIGNAL S5391 : STD_LOGIC;
    SIGNAL S5392 : STD_LOGIC;
    SIGNAL S5393 : STD_LOGIC;
    SIGNAL S5394 : STD_LOGIC;
    SIGNAL S5395 : STD_LOGIC;
    SIGNAL S5396 : STD_LOGIC;
    SIGNAL S5397 : STD_LOGIC;
    SIGNAL S5398 : STD_LOGIC;
    SIGNAL S5399 : STD_LOGIC;
    SIGNAL S5400 : STD_LOGIC;
    SIGNAL S5401 : STD_LOGIC;
    SIGNAL S5402 : STD_LOGIC;
    SIGNAL S5403 : STD_LOGIC;
    SIGNAL S5404 : STD_LOGIC;
    SIGNAL S5405 : STD_LOGIC;
    SIGNAL S5406 : STD_LOGIC;
    SIGNAL S5407 : STD_LOGIC;
    SIGNAL S5408 : STD_LOGIC;
    SIGNAL S5409 : STD_LOGIC;
    SIGNAL S5410 : STD_LOGIC;
    SIGNAL S5411 : STD_LOGIC;
    SIGNAL S5412 : STD_LOGIC;
    SIGNAL S5413 : STD_LOGIC;
    SIGNAL S5414 : STD_LOGIC;
    SIGNAL S5415 : STD_LOGIC;
    SIGNAL S5416 : STD_LOGIC;
    SIGNAL S5417 : STD_LOGIC;
    SIGNAL S5418 : STD_LOGIC;
    SIGNAL S5419 : STD_LOGIC;
    SIGNAL S5420 : STD_LOGIC;
    SIGNAL S5421 : STD_LOGIC;
    SIGNAL S5422 : STD_LOGIC;
    SIGNAL S5423 : STD_LOGIC;
    SIGNAL S5424 : STD_LOGIC;
    SIGNAL S5425 : STD_LOGIC;
    SIGNAL S5426 : STD_LOGIC;
    SIGNAL S5427 : STD_LOGIC;
    SIGNAL S5428 : STD_LOGIC;
    SIGNAL S5429 : STD_LOGIC;
    SIGNAL S5430 : STD_LOGIC;
    SIGNAL S5431 : STD_LOGIC;
    SIGNAL S5432 : STD_LOGIC;
    SIGNAL S5433 : STD_LOGIC;
    SIGNAL S5434 : STD_LOGIC;
    SIGNAL S5435 : STD_LOGIC;
    SIGNAL S5436 : STD_LOGIC;
    SIGNAL S5437 : STD_LOGIC;
    SIGNAL S5438 : STD_LOGIC;
    SIGNAL S5439 : STD_LOGIC;
    SIGNAL S5440 : STD_LOGIC;
    SIGNAL S5441 : STD_LOGIC;
    SIGNAL S5442 : STD_LOGIC;
    SIGNAL S5443 : STD_LOGIC;
    SIGNAL S5444 : STD_LOGIC;
    SIGNAL S5445 : STD_LOGIC;
    SIGNAL S5446 : STD_LOGIC;
    SIGNAL S5447 : STD_LOGIC;
    SIGNAL S5448 : STD_LOGIC;
    SIGNAL S5449 : STD_LOGIC;
    SIGNAL S5450 : STD_LOGIC;
    SIGNAL S5451 : STD_LOGIC;
    SIGNAL S5452 : STD_LOGIC;
    SIGNAL S5453 : STD_LOGIC;
    SIGNAL S5454 : STD_LOGIC;
    SIGNAL S5455 : STD_LOGIC;
    SIGNAL S5456 : STD_LOGIC;
    SIGNAL S5457 : STD_LOGIC;
    SIGNAL S5458 : STD_LOGIC;
    SIGNAL S5459 : STD_LOGIC;
    SIGNAL S5460 : STD_LOGIC;
    SIGNAL S5461 : STD_LOGIC;
    SIGNAL S5462 : STD_LOGIC;
    SIGNAL S5463 : STD_LOGIC;
    SIGNAL S5464 : STD_LOGIC;
    SIGNAL S5465 : STD_LOGIC;
    SIGNAL S5466 : STD_LOGIC;
    SIGNAL S5467 : STD_LOGIC;
    SIGNAL S5468 : STD_LOGIC;
    SIGNAL S5469 : STD_LOGIC;
    SIGNAL S5470 : STD_LOGIC;
    SIGNAL S5471 : STD_LOGIC;
    SIGNAL S5472 : STD_LOGIC;
    SIGNAL S5473 : STD_LOGIC;
    SIGNAL S5474 : STD_LOGIC;
    SIGNAL S5475 : STD_LOGIC;
    SIGNAL S5476 : STD_LOGIC;
    SIGNAL S5477 : STD_LOGIC;
    SIGNAL S5478 : STD_LOGIC;
    SIGNAL S5479 : STD_LOGIC;
    SIGNAL S5480 : STD_LOGIC;
    SIGNAL S5481 : STD_LOGIC;
    SIGNAL S5482 : STD_LOGIC;
    SIGNAL S5483 : STD_LOGIC;
    SIGNAL S5484 : STD_LOGIC;
    SIGNAL S5485 : STD_LOGIC;
    SIGNAL S5486 : STD_LOGIC;
    SIGNAL S5487 : STD_LOGIC;
    SIGNAL S5488 : STD_LOGIC;
    SIGNAL S5489 : STD_LOGIC;
    SIGNAL S5490 : STD_LOGIC;
    SIGNAL S5491 : STD_LOGIC;
    SIGNAL S5492 : STD_LOGIC;
    SIGNAL S5493 : STD_LOGIC;
    SIGNAL S5494 : STD_LOGIC;
    SIGNAL S5495 : STD_LOGIC;
    SIGNAL S5496 : STD_LOGIC;
    SIGNAL S5497 : STD_LOGIC;
    SIGNAL S5498 : STD_LOGIC;
    SIGNAL S5499 : STD_LOGIC;
    SIGNAL S5500 : STD_LOGIC;
    SIGNAL S5501 : STD_LOGIC;
    SIGNAL S5502 : STD_LOGIC;
    SIGNAL S5503 : STD_LOGIC;
    SIGNAL S5504 : STD_LOGIC;
    SIGNAL S5505 : STD_LOGIC;
    SIGNAL S5506 : STD_LOGIC;
    SIGNAL S5507 : STD_LOGIC;
    SIGNAL S5508 : STD_LOGIC;
    SIGNAL S5509 : STD_LOGIC;
    SIGNAL S5510 : STD_LOGIC;
    SIGNAL S5511 : STD_LOGIC;
    SIGNAL S5512 : STD_LOGIC;
    SIGNAL S5513 : STD_LOGIC;
    SIGNAL S5514 : STD_LOGIC;
    SIGNAL S5515 : STD_LOGIC;
    SIGNAL S5516 : STD_LOGIC;
    SIGNAL S5517 : STD_LOGIC;
    SIGNAL S5518 : STD_LOGIC;
    SIGNAL S5519 : STD_LOGIC;
    SIGNAL S5520 : STD_LOGIC;
    SIGNAL S5521 : STD_LOGIC;
    SIGNAL S5522 : STD_LOGIC;
    SIGNAL S5523 : STD_LOGIC;
    SIGNAL S5524 : STD_LOGIC;
    SIGNAL S5525 : STD_LOGIC;
    SIGNAL S5526 : STD_LOGIC;
    SIGNAL S5527 : STD_LOGIC;
    SIGNAL S5528 : STD_LOGIC;
    SIGNAL S5529 : STD_LOGIC;
    SIGNAL S5530 : STD_LOGIC;
    SIGNAL S5531 : STD_LOGIC;
    SIGNAL S5532 : STD_LOGIC;
    SIGNAL S5533 : STD_LOGIC;
    SIGNAL S5534 : STD_LOGIC;
    SIGNAL S5535 : STD_LOGIC;
    SIGNAL S5536 : STD_LOGIC;
    SIGNAL S5537 : STD_LOGIC;
    SIGNAL S5538 : STD_LOGIC;
    SIGNAL S5539 : STD_LOGIC;
    SIGNAL S5540 : STD_LOGIC;
    SIGNAL S5541 : STD_LOGIC;
    SIGNAL S5542 : STD_LOGIC;
    SIGNAL S5543 : STD_LOGIC;
    SIGNAL S5544 : STD_LOGIC;
    SIGNAL S5545 : STD_LOGIC;
    SIGNAL S5546 : STD_LOGIC;
    SIGNAL S5547 : STD_LOGIC;
    SIGNAL S5548 : STD_LOGIC;
    SIGNAL S5549 : STD_LOGIC;
    SIGNAL S5550 : STD_LOGIC;
    SIGNAL S5551 : STD_LOGIC;
    SIGNAL S5552 : STD_LOGIC;
    SIGNAL S5553 : STD_LOGIC;
    SIGNAL S5554 : STD_LOGIC;
    SIGNAL S5555 : STD_LOGIC;
    SIGNAL S5556 : STD_LOGIC;
    SIGNAL S5557 : STD_LOGIC;
    SIGNAL S5558 : STD_LOGIC;
    SIGNAL S5559 : STD_LOGIC;
    SIGNAL S5560 : STD_LOGIC;
    SIGNAL S5561 : STD_LOGIC;
    SIGNAL S5562 : STD_LOGIC;
    SIGNAL S5563 : STD_LOGIC;
    SIGNAL S5564 : STD_LOGIC;
    SIGNAL S5565 : STD_LOGIC;
    SIGNAL S5566 : STD_LOGIC;
    SIGNAL S5567 : STD_LOGIC;
    SIGNAL S5568 : STD_LOGIC;
    SIGNAL S5569 : STD_LOGIC;
    SIGNAL S5570 : STD_LOGIC;
    SIGNAL S5571 : STD_LOGIC;
    SIGNAL S5572 : STD_LOGIC;
    SIGNAL S5573 : STD_LOGIC;
    SIGNAL S5574 : STD_LOGIC;
    SIGNAL S5575 : STD_LOGIC;
    SIGNAL S5576 : STD_LOGIC;
    SIGNAL S5577 : STD_LOGIC;
    SIGNAL S5578 : STD_LOGIC;
    SIGNAL S5579 : STD_LOGIC;
    SIGNAL S5580 : STD_LOGIC;
    SIGNAL S5581 : STD_LOGIC;
    SIGNAL S5582 : STD_LOGIC;
    SIGNAL S5583 : STD_LOGIC;
    SIGNAL S5584 : STD_LOGIC;
    SIGNAL S5585 : STD_LOGIC;
    SIGNAL S5586 : STD_LOGIC;
    SIGNAL S5587 : STD_LOGIC;
    SIGNAL S5588 : STD_LOGIC;
    SIGNAL S5589 : STD_LOGIC;
    SIGNAL S5590 : STD_LOGIC;
    SIGNAL S5591 : STD_LOGIC;
    SIGNAL S5592 : STD_LOGIC;
    SIGNAL S5593 : STD_LOGIC;
    SIGNAL S5594 : STD_LOGIC;
    SIGNAL S5595 : STD_LOGIC;
    SIGNAL S5596 : STD_LOGIC;
    SIGNAL S5597 : STD_LOGIC;
    SIGNAL S5598 : STD_LOGIC;
    SIGNAL S5599 : STD_LOGIC;
    SIGNAL S5600 : STD_LOGIC;
    SIGNAL S5601 : STD_LOGIC;
    SIGNAL S5602 : STD_LOGIC;
    SIGNAL S5603 : STD_LOGIC;
    SIGNAL S5604 : STD_LOGIC;
    SIGNAL S5605 : STD_LOGIC;
    SIGNAL S5606 : STD_LOGIC;
    SIGNAL S5607 : STD_LOGIC;
    SIGNAL S5608 : STD_LOGIC;
    SIGNAL S5609 : STD_LOGIC;
    SIGNAL S5610 : STD_LOGIC;
    SIGNAL S5611 : STD_LOGIC;
    SIGNAL S5612 : STD_LOGIC;
    SIGNAL S5613 : STD_LOGIC;
    SIGNAL S5614 : STD_LOGIC;
    SIGNAL S5615 : STD_LOGIC;
    SIGNAL S5616 : STD_LOGIC;
    SIGNAL S5617 : STD_LOGIC;
    SIGNAL S5618 : STD_LOGIC;
    SIGNAL S5619 : STD_LOGIC;
    SIGNAL S5620 : STD_LOGIC;
    SIGNAL S5621 : STD_LOGIC;
    SIGNAL S5622 : STD_LOGIC;
    SIGNAL S5623 : STD_LOGIC;
    SIGNAL S5624 : STD_LOGIC;
    SIGNAL S5625 : STD_LOGIC;
    SIGNAL S5626 : STD_LOGIC;
    SIGNAL S5627 : STD_LOGIC;
    SIGNAL S5628 : STD_LOGIC;
    SIGNAL S5629 : STD_LOGIC;
    SIGNAL S5630 : STD_LOGIC;
    SIGNAL S5631 : STD_LOGIC;
    SIGNAL S5632 : STD_LOGIC;
    SIGNAL S5633 : STD_LOGIC;
    SIGNAL S5634 : STD_LOGIC;
    SIGNAL S5635 : STD_LOGIC;
    SIGNAL S5636 : STD_LOGIC;
    SIGNAL S5637 : STD_LOGIC;
    SIGNAL S5638 : STD_LOGIC;
    SIGNAL S5639 : STD_LOGIC;
    SIGNAL S5640 : STD_LOGIC;
    SIGNAL S5641 : STD_LOGIC;
    SIGNAL S5642 : STD_LOGIC;
    SIGNAL S5643 : STD_LOGIC;
    SIGNAL S5644 : STD_LOGIC;
    SIGNAL S5645 : STD_LOGIC;
    SIGNAL S5646 : STD_LOGIC;
    SIGNAL S5647 : STD_LOGIC;
    SIGNAL S5648 : STD_LOGIC;
    SIGNAL S5649 : STD_LOGIC;
    SIGNAL S5650 : STD_LOGIC;
    SIGNAL S5651 : STD_LOGIC;
    SIGNAL S5652 : STD_LOGIC;
    SIGNAL S5653 : STD_LOGIC;
    SIGNAL S5654 : STD_LOGIC;
    SIGNAL S5655 : STD_LOGIC;
    SIGNAL S5656 : STD_LOGIC;
    SIGNAL S5657 : STD_LOGIC;
    SIGNAL S5658 : STD_LOGIC;
    SIGNAL S5659 : STD_LOGIC;
    SIGNAL S5660 : STD_LOGIC;
    SIGNAL S5661 : STD_LOGIC;
    SIGNAL S5662 : STD_LOGIC;
    SIGNAL S5663 : STD_LOGIC;
    SIGNAL S5664 : STD_LOGIC;
    SIGNAL S5665 : STD_LOGIC;
    SIGNAL S5666 : STD_LOGIC;
    SIGNAL S5667 : STD_LOGIC;
    SIGNAL S5668 : STD_LOGIC;
    SIGNAL S5669 : STD_LOGIC;
    SIGNAL S5670 : STD_LOGIC;
    SIGNAL S5671 : STD_LOGIC;
    SIGNAL S5672 : STD_LOGIC;
    SIGNAL S5673 : STD_LOGIC;
    SIGNAL S5674 : STD_LOGIC;
    SIGNAL S5675 : STD_LOGIC;
    SIGNAL S5676 : STD_LOGIC;
    SIGNAL S5677 : STD_LOGIC;
    SIGNAL S5678 : STD_LOGIC;
    SIGNAL S5679 : STD_LOGIC;
    SIGNAL S5680 : STD_LOGIC;
    SIGNAL S5681 : STD_LOGIC;
    SIGNAL S5682 : STD_LOGIC;
    SIGNAL S5683 : STD_LOGIC;
    SIGNAL S5684 : STD_LOGIC;
    SIGNAL S5685 : STD_LOGIC;
    SIGNAL S5686 : STD_LOGIC;
    SIGNAL S5687 : STD_LOGIC;
    SIGNAL S5688 : STD_LOGIC;
    SIGNAL S5689 : STD_LOGIC;
    SIGNAL S5690 : STD_LOGIC;
    SIGNAL S5691 : STD_LOGIC;
    SIGNAL S5692 : STD_LOGIC;
    SIGNAL S5693 : STD_LOGIC;
    SIGNAL S5694 : STD_LOGIC;
    SIGNAL S5695 : STD_LOGIC;
    SIGNAL S5696 : STD_LOGIC;
    SIGNAL S5697 : STD_LOGIC;
    SIGNAL S5698 : STD_LOGIC;
    SIGNAL S5699 : STD_LOGIC;
    SIGNAL S5700 : STD_LOGIC;
    SIGNAL S5701 : STD_LOGIC;
    SIGNAL S5702 : STD_LOGIC;
    SIGNAL S5703 : STD_LOGIC;
    SIGNAL S5704 : STD_LOGIC;
    SIGNAL S5705 : STD_LOGIC;
    SIGNAL S5706 : STD_LOGIC;
    SIGNAL S5707 : STD_LOGIC;
    SIGNAL S5708 : STD_LOGIC;
    SIGNAL S5709 : STD_LOGIC;
    SIGNAL S5710 : STD_LOGIC;
    SIGNAL S5711 : STD_LOGIC;
    SIGNAL S5712 : STD_LOGIC;
    SIGNAL S5713 : STD_LOGIC;
    SIGNAL S5714 : STD_LOGIC;
    SIGNAL S5715 : STD_LOGIC;
    SIGNAL S5716 : STD_LOGIC;
    SIGNAL S5717 : STD_LOGIC;
    SIGNAL S5718 : STD_LOGIC;
    SIGNAL S5719 : STD_LOGIC;
    SIGNAL S5720 : STD_LOGIC;
    SIGNAL S5721 : STD_LOGIC;
    SIGNAL S5722 : STD_LOGIC;
    SIGNAL S5723 : STD_LOGIC;
    SIGNAL S5724 : STD_LOGIC;
    SIGNAL S5725 : STD_LOGIC;
    SIGNAL S5726 : STD_LOGIC;
    SIGNAL S5727 : STD_LOGIC;
    SIGNAL S5728 : STD_LOGIC;
    SIGNAL S5729 : STD_LOGIC;
    SIGNAL S5730 : STD_LOGIC;
    SIGNAL S5731 : STD_LOGIC;
    SIGNAL S5732 : STD_LOGIC;
    SIGNAL S5733 : STD_LOGIC;
    SIGNAL S5734 : STD_LOGIC;
    SIGNAL S5735 : STD_LOGIC;
    SIGNAL S5736 : STD_LOGIC;
    SIGNAL S5737 : STD_LOGIC;
    SIGNAL S5738 : STD_LOGIC;
    SIGNAL S5739 : STD_LOGIC;
    SIGNAL S5740 : STD_LOGIC;
    SIGNAL S5741 : STD_LOGIC;
    SIGNAL S5742 : STD_LOGIC;
    SIGNAL S5743 : STD_LOGIC;
    SIGNAL S5744 : STD_LOGIC;
    SIGNAL S5745 : STD_LOGIC;
    SIGNAL S5746 : STD_LOGIC;
    SIGNAL S5747 : STD_LOGIC;
    SIGNAL S5748 : STD_LOGIC;
    SIGNAL S5749 : STD_LOGIC;
    SIGNAL S5750 : STD_LOGIC;
    SIGNAL S5751 : STD_LOGIC;
    SIGNAL S5752 : STD_LOGIC;
    SIGNAL S5753 : STD_LOGIC;
    SIGNAL S5754 : STD_LOGIC;
    SIGNAL S5755 : STD_LOGIC;
    SIGNAL S5756 : STD_LOGIC;
    SIGNAL S5757 : STD_LOGIC;
    SIGNAL S5758 : STD_LOGIC;
    SIGNAL S5759 : STD_LOGIC;
    SIGNAL S5760 : STD_LOGIC;
    SIGNAL S5761 : STD_LOGIC;
    SIGNAL S5762 : STD_LOGIC;
    SIGNAL S5763 : STD_LOGIC;
    SIGNAL S5764 : STD_LOGIC;
    SIGNAL S5765 : STD_LOGIC;
    SIGNAL S5766 : STD_LOGIC;
    SIGNAL S5767 : STD_LOGIC;
    SIGNAL S5768 : STD_LOGIC;
    SIGNAL S5769 : STD_LOGIC;
    SIGNAL S5770 : STD_LOGIC;
    SIGNAL S5771 : STD_LOGIC;
    SIGNAL S5772 : STD_LOGIC;
    SIGNAL S5773 : STD_LOGIC;
    SIGNAL S5774 : STD_LOGIC;
    SIGNAL S5775 : STD_LOGIC;
    SIGNAL S5776 : STD_LOGIC;
    SIGNAL S5777 : STD_LOGIC;
    SIGNAL S5778 : STD_LOGIC;
    SIGNAL S5779 : STD_LOGIC;
    SIGNAL S5780 : STD_LOGIC;
    SIGNAL S5781 : STD_LOGIC;
    SIGNAL S5782 : STD_LOGIC;
    SIGNAL S5783 : STD_LOGIC;
    SIGNAL S5784 : STD_LOGIC;
    SIGNAL S5785 : STD_LOGIC;
    SIGNAL S5786 : STD_LOGIC;
    SIGNAL S5787 : STD_LOGIC;
    SIGNAL S5788 : STD_LOGIC;
    SIGNAL S5789 : STD_LOGIC;
    SIGNAL S5790 : STD_LOGIC;
    SIGNAL S5791 : STD_LOGIC;
    SIGNAL S5792 : STD_LOGIC;
    SIGNAL S5793 : STD_LOGIC;
    SIGNAL S5794 : STD_LOGIC;
    SIGNAL S5795 : STD_LOGIC;
    SIGNAL S5796 : STD_LOGIC;
    SIGNAL S5797 : STD_LOGIC;
    SIGNAL S5798 : STD_LOGIC;
    SIGNAL S5799 : STD_LOGIC;
    SIGNAL S5800 : STD_LOGIC;
    SIGNAL S5801 : STD_LOGIC;
    SIGNAL S5802 : STD_LOGIC;
    SIGNAL S5803 : STD_LOGIC;
    SIGNAL S5804 : STD_LOGIC;
    SIGNAL S5805 : STD_LOGIC;
    SIGNAL S5806 : STD_LOGIC;
    SIGNAL S5807 : STD_LOGIC;
    SIGNAL S5808 : STD_LOGIC;
    SIGNAL S5809 : STD_LOGIC;
    SIGNAL S5810 : STD_LOGIC;
    SIGNAL S5811 : STD_LOGIC;
    SIGNAL S5812 : STD_LOGIC;
    SIGNAL S5813 : STD_LOGIC;
    SIGNAL S5814 : STD_LOGIC;
    SIGNAL S5815 : STD_LOGIC;
    SIGNAL S5816 : STD_LOGIC;
    SIGNAL S5817 : STD_LOGIC;
    SIGNAL S5818 : STD_LOGIC;
    SIGNAL S5819 : STD_LOGIC;
    SIGNAL S5820 : STD_LOGIC;
    SIGNAL S5821 : STD_LOGIC;
    SIGNAL S5822 : STD_LOGIC;
    SIGNAL S5823 : STD_LOGIC;
    SIGNAL S5824 : STD_LOGIC;
    SIGNAL S5825 : STD_LOGIC;
    SIGNAL S5826 : STD_LOGIC;
    SIGNAL S5827 : STD_LOGIC;
    SIGNAL S5828 : STD_LOGIC;
    SIGNAL S5829 : STD_LOGIC;
    SIGNAL S5830 : STD_LOGIC;
    SIGNAL S5831 : STD_LOGIC;
    SIGNAL S5832 : STD_LOGIC;
    SIGNAL S5833 : STD_LOGIC;
    SIGNAL S5834 : STD_LOGIC;
    SIGNAL S5835 : STD_LOGIC;
    SIGNAL S5836 : STD_LOGIC;
    SIGNAL S5837 : STD_LOGIC;
    SIGNAL S5838 : STD_LOGIC;
    SIGNAL S5839 : STD_LOGIC;
    SIGNAL S5840 : STD_LOGIC;
    SIGNAL S5841 : STD_LOGIC;
    SIGNAL S5842 : STD_LOGIC;
    SIGNAL S5843 : STD_LOGIC;
    SIGNAL S5844 : STD_LOGIC;
    SIGNAL S5845 : STD_LOGIC;
    SIGNAL S5846 : STD_LOGIC;
    SIGNAL S5847 : STD_LOGIC;
    SIGNAL S5848 : STD_LOGIC;
    SIGNAL S5849 : STD_LOGIC;
    SIGNAL S5850 : STD_LOGIC;
    SIGNAL S5851 : STD_LOGIC;
    SIGNAL S5852 : STD_LOGIC;
    SIGNAL S5853 : STD_LOGIC;
    SIGNAL S5854 : STD_LOGIC;
    SIGNAL S5855 : STD_LOGIC;
    SIGNAL S5856 : STD_LOGIC;
    SIGNAL S5857 : STD_LOGIC;
    SIGNAL S5858 : STD_LOGIC;
    SIGNAL S5859 : STD_LOGIC;
    SIGNAL S5860 : STD_LOGIC;
    SIGNAL S5861 : STD_LOGIC;
    SIGNAL S5862 : STD_LOGIC;
    SIGNAL S5863 : STD_LOGIC;
    SIGNAL S5864 : STD_LOGIC;
    SIGNAL S5865 : STD_LOGIC;
    SIGNAL S5866 : STD_LOGIC;
    SIGNAL S5867 : STD_LOGIC;
    SIGNAL S5868 : STD_LOGIC;
    SIGNAL S5869 : STD_LOGIC;
    SIGNAL S5870 : STD_LOGIC;
    SIGNAL S5871 : STD_LOGIC;
    SIGNAL S5872 : STD_LOGIC;
    SIGNAL S5873 : STD_LOGIC;
    SIGNAL S5874 : STD_LOGIC;
    SIGNAL S5875 : STD_LOGIC;
    SIGNAL S5876 : STD_LOGIC;
    SIGNAL S5877 : STD_LOGIC;
    SIGNAL S5878 : STD_LOGIC;
    SIGNAL S5879 : STD_LOGIC;
    SIGNAL S5880 : STD_LOGIC;
    SIGNAL S5881 : STD_LOGIC;
    SIGNAL S5882 : STD_LOGIC;
    SIGNAL S5883 : STD_LOGIC;
    SIGNAL S5884 : STD_LOGIC;
    SIGNAL S5885 : STD_LOGIC;
    SIGNAL S5886 : STD_LOGIC;
    SIGNAL S5887 : STD_LOGIC;
    SIGNAL S5888 : STD_LOGIC;
    SIGNAL S5889 : STD_LOGIC;
    SIGNAL S5890 : STD_LOGIC;
    SIGNAL S5891 : STD_LOGIC;
    SIGNAL S5892 : STD_LOGIC;
    SIGNAL S5893 : STD_LOGIC;
    SIGNAL S5894 : STD_LOGIC;
    SIGNAL S5895 : STD_LOGIC;
    SIGNAL S5896 : STD_LOGIC;
    SIGNAL S5897 : STD_LOGIC;
    SIGNAL S5898 : STD_LOGIC;
    SIGNAL S5899 : STD_LOGIC;
    SIGNAL S5900 : STD_LOGIC;
    SIGNAL S5901 : STD_LOGIC;
    SIGNAL S5902 : STD_LOGIC;
    SIGNAL S5903 : STD_LOGIC;
    SIGNAL S5904 : STD_LOGIC;
    SIGNAL S5905 : STD_LOGIC;
    SIGNAL S5906 : STD_LOGIC;
    SIGNAL S5907 : STD_LOGIC;
    SIGNAL S5908 : STD_LOGIC;
    SIGNAL S5909 : STD_LOGIC;
    SIGNAL S5910 : STD_LOGIC;
    SIGNAL S5911 : STD_LOGIC;
    SIGNAL S5912 : STD_LOGIC;
    SIGNAL S5913 : STD_LOGIC;
    SIGNAL S5914 : STD_LOGIC;
    SIGNAL S5915 : STD_LOGIC;
    SIGNAL S5916 : STD_LOGIC;
    SIGNAL S5917 : STD_LOGIC;
    SIGNAL S5918 : STD_LOGIC;
    SIGNAL S5919 : STD_LOGIC;
    SIGNAL S5920 : STD_LOGIC;
    SIGNAL S5921 : STD_LOGIC;
    SIGNAL S5922 : STD_LOGIC;
    SIGNAL S5923 : STD_LOGIC;
    SIGNAL S5924 : STD_LOGIC;
    SIGNAL S5925 : STD_LOGIC;
    SIGNAL S5926 : STD_LOGIC;
    SIGNAL S5927 : STD_LOGIC;
    SIGNAL S5928 : STD_LOGIC;
    SIGNAL S5929 : STD_LOGIC;
    SIGNAL S5930 : STD_LOGIC;
    SIGNAL S5931 : STD_LOGIC;
    SIGNAL S5932 : STD_LOGIC;
    SIGNAL S5933 : STD_LOGIC;
    SIGNAL S5934 : STD_LOGIC;
    SIGNAL S5935 : STD_LOGIC;
    SIGNAL S5936 : STD_LOGIC;
    SIGNAL S5937 : STD_LOGIC;
    SIGNAL S5938 : STD_LOGIC;
    SIGNAL S5939 : STD_LOGIC;
    SIGNAL S5940 : STD_LOGIC;
    SIGNAL S5941 : STD_LOGIC;
    SIGNAL S5942 : STD_LOGIC;
    SIGNAL S5943 : STD_LOGIC;
    SIGNAL S5944 : STD_LOGIC;
    SIGNAL S5945 : STD_LOGIC;
    SIGNAL S5946 : STD_LOGIC;
    SIGNAL S5947 : STD_LOGIC;
    SIGNAL S5948 : STD_LOGIC;
    SIGNAL S5949 : STD_LOGIC;
    SIGNAL S5950 : STD_LOGIC;
    SIGNAL S5951 : STD_LOGIC;
    SIGNAL S5952 : STD_LOGIC;
    SIGNAL S5953 : STD_LOGIC;
    SIGNAL S5954 : STD_LOGIC;
    SIGNAL S5955 : STD_LOGIC;
    SIGNAL S5956 : STD_LOGIC;
    SIGNAL S5957 : STD_LOGIC;
    SIGNAL S5958 : STD_LOGIC;
    SIGNAL S5959 : STD_LOGIC;
    SIGNAL S5960 : STD_LOGIC;
    SIGNAL S5961 : STD_LOGIC;
    SIGNAL S5962 : STD_LOGIC;
    SIGNAL S5963 : STD_LOGIC;
    SIGNAL S5964 : STD_LOGIC;
    SIGNAL S5965 : STD_LOGIC;
    SIGNAL S5966 : STD_LOGIC;
    SIGNAL S5967 : STD_LOGIC;
    SIGNAL S5968 : STD_LOGIC;
    SIGNAL S5969 : STD_LOGIC;
    SIGNAL S5970 : STD_LOGIC;
    SIGNAL S5971 : STD_LOGIC;
    SIGNAL S5972 : STD_LOGIC;
    SIGNAL S5973 : STD_LOGIC;
    SIGNAL S5974 : STD_LOGIC;
    SIGNAL S5975 : STD_LOGIC;
    SIGNAL S5976 : STD_LOGIC;
    SIGNAL S5977 : STD_LOGIC;
    SIGNAL S5978 : STD_LOGIC;
    SIGNAL S5979 : STD_LOGIC;
    SIGNAL S5980 : STD_LOGIC;
    SIGNAL S5981 : STD_LOGIC;
    SIGNAL S5982 : STD_LOGIC;
    SIGNAL S5983 : STD_LOGIC;
    SIGNAL S5984 : STD_LOGIC;
    SIGNAL S5985 : STD_LOGIC;
    SIGNAL S5986 : STD_LOGIC;
    SIGNAL S5987 : STD_LOGIC;
    SIGNAL S5988 : STD_LOGIC;
    SIGNAL S5989 : STD_LOGIC;
    SIGNAL S5990 : STD_LOGIC;
    SIGNAL S5991 : STD_LOGIC;
    SIGNAL S5992 : STD_LOGIC;
    SIGNAL S5993 : STD_LOGIC;
    SIGNAL S5994 : STD_LOGIC;
    SIGNAL S5995 : STD_LOGIC;
    SIGNAL S5996 : STD_LOGIC;
    SIGNAL S5997 : STD_LOGIC;
    SIGNAL S5998 : STD_LOGIC;
    SIGNAL S5999 : STD_LOGIC;
    SIGNAL S6000 : STD_LOGIC;
    SIGNAL S6001 : STD_LOGIC;
    SIGNAL S6002 : STD_LOGIC;
    SIGNAL S6003 : STD_LOGIC;
    SIGNAL S6004 : STD_LOGIC;
    SIGNAL S6005 : STD_LOGIC;
    SIGNAL S6006 : STD_LOGIC;
    SIGNAL S6007 : STD_LOGIC;
    SIGNAL S6008 : STD_LOGIC;
    SIGNAL S6009 : STD_LOGIC;
    SIGNAL S6010 : STD_LOGIC;
    SIGNAL S6011 : STD_LOGIC;
    SIGNAL S6012 : STD_LOGIC;
    SIGNAL S6013 : STD_LOGIC;
    SIGNAL S6014 : STD_LOGIC;
    SIGNAL S6015 : STD_LOGIC;
    SIGNAL S6016 : STD_LOGIC;
    SIGNAL S6017 : STD_LOGIC;
    SIGNAL S6018 : STD_LOGIC;
    SIGNAL S6019 : STD_LOGIC;
    SIGNAL S6020 : STD_LOGIC;
    SIGNAL S6021 : STD_LOGIC;
    SIGNAL S6022 : STD_LOGIC;
    SIGNAL S6023 : STD_LOGIC;
    SIGNAL S6024 : STD_LOGIC;
    SIGNAL S6025 : STD_LOGIC;
    SIGNAL S6026 : STD_LOGIC;
    SIGNAL S6027 : STD_LOGIC;
    SIGNAL S6028 : STD_LOGIC;
    SIGNAL S6029 : STD_LOGIC;
    SIGNAL S6030 : STD_LOGIC;
    SIGNAL S6031 : STD_LOGIC;
    SIGNAL S6032 : STD_LOGIC;
    SIGNAL S6033 : STD_LOGIC;
    SIGNAL S6034 : STD_LOGIC;
    SIGNAL S6035 : STD_LOGIC;
    SIGNAL S6036 : STD_LOGIC;
    SIGNAL S6037 : STD_LOGIC;
    SIGNAL S6038 : STD_LOGIC;
    SIGNAL S6039 : STD_LOGIC;
    SIGNAL S6040 : STD_LOGIC;
    SIGNAL S6041 : STD_LOGIC;
    SIGNAL S6042 : STD_LOGIC;
    SIGNAL S6043 : STD_LOGIC;
    SIGNAL S6044 : STD_LOGIC;
    SIGNAL S6045 : STD_LOGIC;
    SIGNAL S6046 : STD_LOGIC;
    SIGNAL S6047 : STD_LOGIC;
    SIGNAL S6048 : STD_LOGIC;
    SIGNAL S6049 : STD_LOGIC;
    SIGNAL S6050 : STD_LOGIC;
    SIGNAL S6051 : STD_LOGIC;
    SIGNAL S6052 : STD_LOGIC;
    SIGNAL S6053 : STD_LOGIC;
    SIGNAL S6054 : STD_LOGIC;
    SIGNAL S6055 : STD_LOGIC;
    SIGNAL S6056 : STD_LOGIC;
    SIGNAL S6057 : STD_LOGIC;
    SIGNAL S6058 : STD_LOGIC;
    SIGNAL S6059 : STD_LOGIC;
    SIGNAL S6060 : STD_LOGIC;
    SIGNAL S6061 : STD_LOGIC;
    SIGNAL S6062 : STD_LOGIC;
    SIGNAL S6063 : STD_LOGIC;
    SIGNAL S6064 : STD_LOGIC;
    SIGNAL S6065 : STD_LOGIC;
    SIGNAL S6066 : STD_LOGIC;
    SIGNAL S6067 : STD_LOGIC;
    SIGNAL S6068 : STD_LOGIC;
    SIGNAL S6069 : STD_LOGIC;
    SIGNAL S6070 : STD_LOGIC;
    SIGNAL S6071 : STD_LOGIC;
    SIGNAL S6072 : STD_LOGIC;
    SIGNAL S6073 : STD_LOGIC;
    SIGNAL S6074 : STD_LOGIC;
    SIGNAL S6075 : STD_LOGIC;
    SIGNAL S6076 : STD_LOGIC;
    SIGNAL S6077 : STD_LOGIC;
    SIGNAL S6078 : STD_LOGIC;
    SIGNAL S6079 : STD_LOGIC;
    SIGNAL S6080 : STD_LOGIC;
    SIGNAL S6081 : STD_LOGIC;
    SIGNAL S6082 : STD_LOGIC;
    SIGNAL S6083 : STD_LOGIC;
    SIGNAL S6084 : STD_LOGIC;
    SIGNAL S6085 : STD_LOGIC;
    SIGNAL S6086 : STD_LOGIC;
    SIGNAL S6087 : STD_LOGIC;
    SIGNAL S6088 : STD_LOGIC;
    SIGNAL S6089 : STD_LOGIC;
    SIGNAL S6090 : STD_LOGIC;
    SIGNAL S6091 : STD_LOGIC;
    SIGNAL S6092 : STD_LOGIC;
    SIGNAL S6093 : STD_LOGIC;
    SIGNAL S6094 : STD_LOGIC;
    SIGNAL S6095 : STD_LOGIC;
    SIGNAL S6096 : STD_LOGIC;
    SIGNAL S6097 : STD_LOGIC;
    SIGNAL S6098 : STD_LOGIC;
    SIGNAL S6099 : STD_LOGIC;
    SIGNAL S6100 : STD_LOGIC;
    SIGNAL S6101 : STD_LOGIC;
    SIGNAL S6102 : STD_LOGIC;
    SIGNAL S6103 : STD_LOGIC;
    SIGNAL S6104 : STD_LOGIC;
    SIGNAL S6105 : STD_LOGIC;
    SIGNAL S6106 : STD_LOGIC;
    SIGNAL S6107 : STD_LOGIC;
    SIGNAL S6108 : STD_LOGIC;
    SIGNAL S6109 : STD_LOGIC;
    SIGNAL S6110 : STD_LOGIC;
    SIGNAL S6111 : STD_LOGIC;
    SIGNAL S6112 : STD_LOGIC;
    SIGNAL S6113 : STD_LOGIC;
    SIGNAL S6114 : STD_LOGIC;
    SIGNAL S6115 : STD_LOGIC;
    SIGNAL S6116 : STD_LOGIC;
    SIGNAL S6117 : STD_LOGIC;
    SIGNAL S6118 : STD_LOGIC;
    SIGNAL S6119 : STD_LOGIC;
    SIGNAL S6120 : STD_LOGIC;
    SIGNAL S6121 : STD_LOGIC;
    SIGNAL S6122 : STD_LOGIC;
    SIGNAL S6123 : STD_LOGIC;
    SIGNAL S6124 : STD_LOGIC;
    SIGNAL S6125 : STD_LOGIC;
    SIGNAL S6126 : STD_LOGIC;
    SIGNAL S6127 : STD_LOGIC;
    SIGNAL S6128 : STD_LOGIC;
    SIGNAL S6129 : STD_LOGIC;
    SIGNAL S6130 : STD_LOGIC;
    SIGNAL S6131 : STD_LOGIC;
    SIGNAL S6132 : STD_LOGIC;
    SIGNAL S6133 : STD_LOGIC;
    SIGNAL S6134 : STD_LOGIC;
    SIGNAL S6135 : STD_LOGIC;
    SIGNAL S6136 : STD_LOGIC;
    SIGNAL S6137 : STD_LOGIC;
    SIGNAL S6138 : STD_LOGIC;
    SIGNAL S6139 : STD_LOGIC;
    SIGNAL S6140 : STD_LOGIC;
    SIGNAL S6141 : STD_LOGIC;
    SIGNAL S6142 : STD_LOGIC;
    SIGNAL S6143 : STD_LOGIC;
    SIGNAL S6144 : STD_LOGIC;
    SIGNAL S6145 : STD_LOGIC;
    SIGNAL S6146 : STD_LOGIC;
    SIGNAL S6147 : STD_LOGIC;
    SIGNAL S6148 : STD_LOGIC;
    SIGNAL S6149 : STD_LOGIC;
    SIGNAL S6150 : STD_LOGIC;
    SIGNAL S6151 : STD_LOGIC;
    SIGNAL S6152 : STD_LOGIC;
    SIGNAL S6153 : STD_LOGIC;
    SIGNAL S6154 : STD_LOGIC;
    SIGNAL S6155 : STD_LOGIC;
    SIGNAL S6156 : STD_LOGIC;
    SIGNAL S6157 : STD_LOGIC;
    SIGNAL S6158 : STD_LOGIC;
    SIGNAL S6159 : STD_LOGIC;
    SIGNAL S6160 : STD_LOGIC;
    SIGNAL S6161 : STD_LOGIC;
    SIGNAL S6162 : STD_LOGIC;
    SIGNAL S6163 : STD_LOGIC;
    SIGNAL S6164 : STD_LOGIC;
    SIGNAL S6165 : STD_LOGIC;
    SIGNAL S6166 : STD_LOGIC;
    SIGNAL S6167 : STD_LOGIC;
    SIGNAL S6168 : STD_LOGIC;
    SIGNAL S6169 : STD_LOGIC;
    SIGNAL S6170 : STD_LOGIC;
    SIGNAL S6171 : STD_LOGIC;
    SIGNAL S6172 : STD_LOGIC;
    SIGNAL S6173 : STD_LOGIC;
    SIGNAL S6174 : STD_LOGIC;
    SIGNAL S6175 : STD_LOGIC;
    SIGNAL S6176 : STD_LOGIC;
    SIGNAL S6177 : STD_LOGIC;
    SIGNAL S6178 : STD_LOGIC;
    SIGNAL S6179 : STD_LOGIC;
    SIGNAL S6180 : STD_LOGIC;
    SIGNAL S6181 : STD_LOGIC;
    SIGNAL S6182 : STD_LOGIC;
    SIGNAL S6183 : STD_LOGIC;
    SIGNAL S6184 : STD_LOGIC;
    SIGNAL S6185 : STD_LOGIC;
    SIGNAL S6186 : STD_LOGIC;
    SIGNAL S6187 : STD_LOGIC;
    SIGNAL S6188 : STD_LOGIC;
    SIGNAL S6189 : STD_LOGIC;
    SIGNAL S6190 : STD_LOGIC;
    SIGNAL S6191 : STD_LOGIC;
    SIGNAL S6192 : STD_LOGIC;
    SIGNAL S6193 : STD_LOGIC;
    SIGNAL S6194 : STD_LOGIC;
    SIGNAL S6195 : STD_LOGIC;
    SIGNAL S6196 : STD_LOGIC;
    SIGNAL S6197 : STD_LOGIC;
    SIGNAL S6198 : STD_LOGIC;
    SIGNAL S6199 : STD_LOGIC;
    SIGNAL S6200 : STD_LOGIC;
    SIGNAL S6201 : STD_LOGIC;
    SIGNAL S6202 : STD_LOGIC;
    SIGNAL S6203 : STD_LOGIC;
    SIGNAL S6204 : STD_LOGIC;
    SIGNAL S6205 : STD_LOGIC;
    SIGNAL S6206 : STD_LOGIC;
    SIGNAL S6207 : STD_LOGIC;
    SIGNAL S6208 : STD_LOGIC;
    SIGNAL S6209 : STD_LOGIC;
    SIGNAL S6210 : STD_LOGIC;
    SIGNAL S6211 : STD_LOGIC;
    SIGNAL S6212 : STD_LOGIC;
    SIGNAL S6213 : STD_LOGIC;
    SIGNAL S6214 : STD_LOGIC;
    SIGNAL S6215 : STD_LOGIC;
    SIGNAL S6216 : STD_LOGIC;
    SIGNAL S6217 : STD_LOGIC;
    SIGNAL S6218 : STD_LOGIC;
    SIGNAL S6219 : STD_LOGIC;
    SIGNAL S6220 : STD_LOGIC;
    SIGNAL S6221 : STD_LOGIC;
    SIGNAL S6222 : STD_LOGIC;
    SIGNAL S6223 : STD_LOGIC;
    SIGNAL S6224 : STD_LOGIC;
    SIGNAL S6225 : STD_LOGIC;
    SIGNAL S6226 : STD_LOGIC;
    SIGNAL S6227 : STD_LOGIC;
    SIGNAL S6228 : STD_LOGIC;
    SIGNAL S6229 : STD_LOGIC;
    SIGNAL S6230 : STD_LOGIC;
    SIGNAL S6231 : STD_LOGIC;
    SIGNAL S6232 : STD_LOGIC;
    SIGNAL S6233 : STD_LOGIC;
    SIGNAL S6234 : STD_LOGIC;
    SIGNAL S6235 : STD_LOGIC;
    SIGNAL S6236 : STD_LOGIC;
    SIGNAL S6237 : STD_LOGIC;
    SIGNAL S6238 : STD_LOGIC;
    SIGNAL S6239 : STD_LOGIC;
    SIGNAL S6240 : STD_LOGIC;
    SIGNAL S6241 : STD_LOGIC;
    SIGNAL S6242 : STD_LOGIC;
    SIGNAL S6243 : STD_LOGIC;
    SIGNAL S6244 : STD_LOGIC;
    SIGNAL S6245 : STD_LOGIC;
    SIGNAL S6246 : STD_LOGIC;
    SIGNAL S6247 : STD_LOGIC;
    SIGNAL S6248 : STD_LOGIC;
    SIGNAL S6249 : STD_LOGIC;
    SIGNAL S6250 : STD_LOGIC;
    SIGNAL S6251 : STD_LOGIC;
    SIGNAL S6252 : STD_LOGIC;
    SIGNAL S6253 : STD_LOGIC;
    SIGNAL S6254 : STD_LOGIC;
    SIGNAL S6255 : STD_LOGIC;
    SIGNAL S6256 : STD_LOGIC;
    SIGNAL S6257 : STD_LOGIC;
    SIGNAL S6258 : STD_LOGIC;
    SIGNAL S6259 : STD_LOGIC;
    SIGNAL S6260 : STD_LOGIC;
    SIGNAL S6261 : STD_LOGIC;
    SIGNAL S6262 : STD_LOGIC;
    SIGNAL S6263 : STD_LOGIC;
    SIGNAL S6264 : STD_LOGIC;
    SIGNAL S6265 : STD_LOGIC;
    SIGNAL S6266 : STD_LOGIC;
    SIGNAL S6267 : STD_LOGIC;
    SIGNAL S6268 : STD_LOGIC;
    SIGNAL S6269 : STD_LOGIC;
    SIGNAL S6270 : STD_LOGIC;
    SIGNAL S6271 : STD_LOGIC;
    SIGNAL S6272 : STD_LOGIC;
    SIGNAL S6273 : STD_LOGIC;
    SIGNAL S6274 : STD_LOGIC;
    SIGNAL S6275 : STD_LOGIC;
    SIGNAL S6276 : STD_LOGIC;
    SIGNAL S6277 : STD_LOGIC;
    SIGNAL S6278 : STD_LOGIC;
    SIGNAL S6279 : STD_LOGIC;
    SIGNAL S6280 : STD_LOGIC;
    SIGNAL S6281 : STD_LOGIC;
    SIGNAL S6282 : STD_LOGIC;
    SIGNAL S6283 : STD_LOGIC;
    SIGNAL S6284 : STD_LOGIC;
    SIGNAL S6285 : STD_LOGIC;
    SIGNAL S6286 : STD_LOGIC;
    SIGNAL S6287 : STD_LOGIC;
    SIGNAL S6288 : STD_LOGIC;
    SIGNAL S6289 : STD_LOGIC;
    SIGNAL S6290 : STD_LOGIC;
    SIGNAL S6291 : STD_LOGIC;
    SIGNAL S6292 : STD_LOGIC;
    SIGNAL S6293 : STD_LOGIC;
    SIGNAL S6294 : STD_LOGIC;
    SIGNAL S6295 : STD_LOGIC;
    SIGNAL S6296 : STD_LOGIC;
    SIGNAL S6297 : STD_LOGIC;
    SIGNAL S6298 : STD_LOGIC;
    SIGNAL S6299 : STD_LOGIC;
    SIGNAL S6300 : STD_LOGIC;
    SIGNAL S6301 : STD_LOGIC;
    SIGNAL S6302 : STD_LOGIC;
    SIGNAL S6303 : STD_LOGIC;
    SIGNAL S6304 : STD_LOGIC;
    SIGNAL S6305 : STD_LOGIC;
    SIGNAL S6306 : STD_LOGIC;
    SIGNAL S6307 : STD_LOGIC;
    SIGNAL S6308 : STD_LOGIC;
    SIGNAL S6309 : STD_LOGIC;
    SIGNAL S6310 : STD_LOGIC;
    SIGNAL S6311 : STD_LOGIC;
    SIGNAL S6312 : STD_LOGIC;
    SIGNAL S6313 : STD_LOGIC;
    SIGNAL S6314 : STD_LOGIC;
    SIGNAL S6315 : STD_LOGIC;
    SIGNAL S6316 : STD_LOGIC;
    SIGNAL S6317 : STD_LOGIC;
    SIGNAL S6318 : STD_LOGIC;
    SIGNAL S6319 : STD_LOGIC;
    SIGNAL S6320 : STD_LOGIC;
    SIGNAL S6321 : STD_LOGIC;
    SIGNAL S6322 : STD_LOGIC;
    SIGNAL S6323 : STD_LOGIC;
    SIGNAL S6324 : STD_LOGIC;
    SIGNAL S6325 : STD_LOGIC;
    SIGNAL S6326 : STD_LOGIC;
    SIGNAL S6327 : STD_LOGIC;
    SIGNAL S6328 : STD_LOGIC;
    SIGNAL S6329 : STD_LOGIC;
    SIGNAL S6330 : STD_LOGIC;
    SIGNAL S6331 : STD_LOGIC;
    SIGNAL S6332 : STD_LOGIC;
    SIGNAL S6333 : STD_LOGIC;
    SIGNAL S6334 : STD_LOGIC;
    SIGNAL S6335 : STD_LOGIC;
    SIGNAL S6336 : STD_LOGIC;
    SIGNAL S6337 : STD_LOGIC;
    SIGNAL S6338 : STD_LOGIC;
    SIGNAL S6339 : STD_LOGIC;
    SIGNAL S6340 : STD_LOGIC;
    SIGNAL S6341 : STD_LOGIC;
    SIGNAL S6342 : STD_LOGIC;
    SIGNAL S6343 : STD_LOGIC;
    SIGNAL S6344 : STD_LOGIC;
    SIGNAL S6345 : STD_LOGIC;
    SIGNAL S6346 : STD_LOGIC;
    SIGNAL S6347 : STD_LOGIC;
    SIGNAL S6348 : STD_LOGIC;
    SIGNAL S6349 : STD_LOGIC;
    SIGNAL S6350 : STD_LOGIC;
    SIGNAL S6351 : STD_LOGIC;
    SIGNAL S6352 : STD_LOGIC;
    SIGNAL S6353 : STD_LOGIC;
    SIGNAL S6354 : STD_LOGIC;
    SIGNAL S6355 : STD_LOGIC;
    SIGNAL S6356 : STD_LOGIC;
    SIGNAL S6357 : STD_LOGIC;
    SIGNAL S6358 : STD_LOGIC;
    SIGNAL S6359 : STD_LOGIC;
    SIGNAL S6360 : STD_LOGIC;
    SIGNAL S6361 : STD_LOGIC;
    SIGNAL S6362 : STD_LOGIC;
    SIGNAL S6363 : STD_LOGIC;
    SIGNAL S6364 : STD_LOGIC;
    SIGNAL S6365 : STD_LOGIC;
    SIGNAL S6366 : STD_LOGIC;
    SIGNAL S6367 : STD_LOGIC;
    SIGNAL S6368 : STD_LOGIC;
    SIGNAL S6369 : STD_LOGIC;
    SIGNAL S6370 : STD_LOGIC;
    SIGNAL S6371 : STD_LOGIC;
    SIGNAL S6372 : STD_LOGIC;
    SIGNAL S6373 : STD_LOGIC;
    SIGNAL S6374 : STD_LOGIC;
    SIGNAL S6375 : STD_LOGIC;
    SIGNAL S6376 : STD_LOGIC;
    SIGNAL S6377 : STD_LOGIC;
    SIGNAL S6378 : STD_LOGIC;
    SIGNAL S6379 : STD_LOGIC;
    SIGNAL S6380 : STD_LOGIC;
    SIGNAL S6381 : STD_LOGIC;
    SIGNAL S6382 : STD_LOGIC;
    SIGNAL S6383 : STD_LOGIC;
    SIGNAL S6384 : STD_LOGIC;
    SIGNAL S6385 : STD_LOGIC;
    SIGNAL S6386 : STD_LOGIC;
    SIGNAL S6387 : STD_LOGIC;
    SIGNAL S6388 : STD_LOGIC;
    SIGNAL S6389 : STD_LOGIC;
    SIGNAL S6390 : STD_LOGIC;
    SIGNAL S6391 : STD_LOGIC;
    SIGNAL S6392 : STD_LOGIC;
    SIGNAL S6393 : STD_LOGIC;
    SIGNAL S6394 : STD_LOGIC;
    SIGNAL S6395 : STD_LOGIC;
    SIGNAL S6396 : STD_LOGIC;
    SIGNAL S6397 : STD_LOGIC;
    SIGNAL S6398 : STD_LOGIC;
    SIGNAL S6399 : STD_LOGIC;
    SIGNAL S6400 : STD_LOGIC;
    SIGNAL S6401 : STD_LOGIC;
    SIGNAL S6402 : STD_LOGIC;
    SIGNAL S6403 : STD_LOGIC;
    SIGNAL S6404 : STD_LOGIC;
    SIGNAL S6405 : STD_LOGIC;
    SIGNAL S6406 : STD_LOGIC;
    SIGNAL S6407 : STD_LOGIC;
    SIGNAL S6408 : STD_LOGIC;
    SIGNAL S6409 : STD_LOGIC;
    SIGNAL S6410 : STD_LOGIC;
    SIGNAL S6411 : STD_LOGIC;
    SIGNAL S6412 : STD_LOGIC;
    SIGNAL S6413 : STD_LOGIC;
    SIGNAL S6414 : STD_LOGIC;
    SIGNAL S6415 : STD_LOGIC;
    SIGNAL S6416 : STD_LOGIC;
    SIGNAL S6417 : STD_LOGIC;
    SIGNAL S6418 : STD_LOGIC;
    SIGNAL S6419 : STD_LOGIC;
    SIGNAL S6420 : STD_LOGIC;
    SIGNAL S6421 : STD_LOGIC;
    SIGNAL S6422 : STD_LOGIC;
    SIGNAL S6423 : STD_LOGIC;
    SIGNAL S6424 : STD_LOGIC;
    SIGNAL S6425 : STD_LOGIC;
    SIGNAL S6426 : STD_LOGIC;
    SIGNAL S6427 : STD_LOGIC;
    SIGNAL S6428 : STD_LOGIC;
    SIGNAL S6429 : STD_LOGIC;
    SIGNAL S6430 : STD_LOGIC;
    SIGNAL S6431 : STD_LOGIC;
    SIGNAL S6432 : STD_LOGIC;
    SIGNAL S6433 : STD_LOGIC;
    SIGNAL S6434 : STD_LOGIC;
    SIGNAL S6435 : STD_LOGIC;
    SIGNAL S6436 : STD_LOGIC;
    SIGNAL S6437 : STD_LOGIC;
    SIGNAL S6438 : STD_LOGIC;
    SIGNAL S6439 : STD_LOGIC;
    SIGNAL S6440 : STD_LOGIC;
    SIGNAL S6441 : STD_LOGIC;
    SIGNAL S6442 : STD_LOGIC;
    SIGNAL S6443 : STD_LOGIC;
    SIGNAL S6444 : STD_LOGIC;
    SIGNAL S6445 : STD_LOGIC;
    SIGNAL S6446 : STD_LOGIC;
    SIGNAL S6447 : STD_LOGIC;
    SIGNAL S6448 : STD_LOGIC;
    SIGNAL S6449 : STD_LOGIC;
    SIGNAL S6450 : STD_LOGIC;
    SIGNAL S6451 : STD_LOGIC;
    SIGNAL S6452 : STD_LOGIC;
    SIGNAL S6453 : STD_LOGIC;
    SIGNAL S6454 : STD_LOGIC;
    SIGNAL S6455 : STD_LOGIC;
    SIGNAL S6456 : STD_LOGIC;
    SIGNAL S6457 : STD_LOGIC;
    SIGNAL S6458 : STD_LOGIC;
    SIGNAL S6459 : STD_LOGIC;
    SIGNAL S6460 : STD_LOGIC;
    SIGNAL S6461 : STD_LOGIC;
    SIGNAL S6462 : STD_LOGIC;
    SIGNAL S6463 : STD_LOGIC;
    SIGNAL S6464 : STD_LOGIC;
    SIGNAL S6465 : STD_LOGIC;
    SIGNAL S6466 : STD_LOGIC;
    SIGNAL S6467 : STD_LOGIC;
    SIGNAL S6468 : STD_LOGIC;
    SIGNAL S6469 : STD_LOGIC;
    SIGNAL S6470 : STD_LOGIC;
    SIGNAL S6471 : STD_LOGIC;
    SIGNAL S6472 : STD_LOGIC;
    SIGNAL S6473 : STD_LOGIC;
    SIGNAL S6474 : STD_LOGIC;
    SIGNAL S6475 : STD_LOGIC;
    SIGNAL S6476 : STD_LOGIC;
    SIGNAL S6477 : STD_LOGIC;
    SIGNAL S6478 : STD_LOGIC;
    SIGNAL S6479 : STD_LOGIC;
    SIGNAL S6480 : STD_LOGIC;
    SIGNAL S6481 : STD_LOGIC;
    SIGNAL S6482 : STD_LOGIC;
    SIGNAL S6483 : STD_LOGIC;
    SIGNAL S6484 : STD_LOGIC;
    SIGNAL S6485 : STD_LOGIC;
    SIGNAL S6486 : STD_LOGIC;
    SIGNAL S6487 : STD_LOGIC;
    SIGNAL S6488 : STD_LOGIC;
    SIGNAL S6489 : STD_LOGIC;
    SIGNAL S6490 : STD_LOGIC;
    SIGNAL S6491 : STD_LOGIC;
    SIGNAL S6492 : STD_LOGIC;
    SIGNAL S6493 : STD_LOGIC;
    SIGNAL S6494 : STD_LOGIC;
    SIGNAL S6495 : STD_LOGIC;
    SIGNAL S6496 : STD_LOGIC;
    SIGNAL S6497 : STD_LOGIC;
    SIGNAL S6498 : STD_LOGIC;
    SIGNAL S6499 : STD_LOGIC;
    SIGNAL S6500 : STD_LOGIC;
    SIGNAL S6501 : STD_LOGIC;
    SIGNAL S6502 : STD_LOGIC;
    SIGNAL S6503 : STD_LOGIC;
    SIGNAL S6504 : STD_LOGIC;
    SIGNAL S6505 : STD_LOGIC;
    SIGNAL S6506 : STD_LOGIC;
    SIGNAL S6507 : STD_LOGIC;
    SIGNAL S6508 : STD_LOGIC;
    SIGNAL S6509 : STD_LOGIC;
    SIGNAL S6510 : STD_LOGIC;
    SIGNAL S6511 : STD_LOGIC;
    SIGNAL S6512 : STD_LOGIC;
    SIGNAL S6513 : STD_LOGIC;
    SIGNAL S6514 : STD_LOGIC;
    SIGNAL S6515 : STD_LOGIC;
    SIGNAL S6516 : STD_LOGIC;
    SIGNAL S6517 : STD_LOGIC;
    SIGNAL S6518 : STD_LOGIC;
    SIGNAL S6519 : STD_LOGIC;
    SIGNAL S6520 : STD_LOGIC;
    SIGNAL S6521 : STD_LOGIC;
    SIGNAL S6522 : STD_LOGIC;
    SIGNAL S6523 : STD_LOGIC;
    SIGNAL S6524 : STD_LOGIC;
    SIGNAL S6525 : STD_LOGIC;
    SIGNAL S6526 : STD_LOGIC;
    SIGNAL S6527 : STD_LOGIC;
    SIGNAL S6528 : STD_LOGIC;
    SIGNAL S6529 : STD_LOGIC;
    SIGNAL S6530 : STD_LOGIC;
    SIGNAL S6531 : STD_LOGIC;
    SIGNAL S6532 : STD_LOGIC;
    SIGNAL S6533 : STD_LOGIC;
    SIGNAL S6534 : STD_LOGIC;
    SIGNAL S6535 : STD_LOGIC;
    SIGNAL S6536 : STD_LOGIC;
    SIGNAL S6537 : STD_LOGIC;
    SIGNAL S6538 : STD_LOGIC;
    SIGNAL S6539 : STD_LOGIC;
    SIGNAL S6540 : STD_LOGIC;
    SIGNAL S6541 : STD_LOGIC;
    SIGNAL S6542 : STD_LOGIC;
    SIGNAL S6543 : STD_LOGIC;
    SIGNAL S6544 : STD_LOGIC;
    SIGNAL S6545 : STD_LOGIC;
    SIGNAL S6546 : STD_LOGIC;
    SIGNAL S6547 : STD_LOGIC;
    SIGNAL S6548 : STD_LOGIC;
    SIGNAL S6549 : STD_LOGIC;
    SIGNAL S6550 : STD_LOGIC;
    SIGNAL S6551 : STD_LOGIC;
    SIGNAL S6552 : STD_LOGIC;
    SIGNAL S6553 : STD_LOGIC;
    SIGNAL S6554 : STD_LOGIC;
    SIGNAL S6555 : STD_LOGIC;
    SIGNAL S6556 : STD_LOGIC;
    SIGNAL S6557 : STD_LOGIC;
    SIGNAL S6558 : STD_LOGIC;
    SIGNAL S6559 : STD_LOGIC;
    SIGNAL S6560 : STD_LOGIC;
    SIGNAL S6561 : STD_LOGIC;
    SIGNAL S6562 : STD_LOGIC;
    SIGNAL S6563 : STD_LOGIC;
    SIGNAL S6564 : STD_LOGIC;
    SIGNAL S6565 : STD_LOGIC;
    SIGNAL S6566 : STD_LOGIC;
    SIGNAL S6567 : STD_LOGIC;
    SIGNAL S6568 : STD_LOGIC;
    SIGNAL S6569 : STD_LOGIC;
    SIGNAL S6570 : STD_LOGIC;
    SIGNAL S6571 : STD_LOGIC;
    SIGNAL S6572 : STD_LOGIC;
    SIGNAL S6573 : STD_LOGIC;
    SIGNAL S6574 : STD_LOGIC;
    SIGNAL S6575 : STD_LOGIC;
    SIGNAL S6576 : STD_LOGIC;
    SIGNAL S6577 : STD_LOGIC;
    SIGNAL S6578 : STD_LOGIC;
    SIGNAL S6579 : STD_LOGIC;
    SIGNAL S6580 : STD_LOGIC;
    SIGNAL S6581 : STD_LOGIC;
    SIGNAL S6582 : STD_LOGIC;
    SIGNAL S6583 : STD_LOGIC;
    SIGNAL S6584 : STD_LOGIC;
    SIGNAL S6585 : STD_LOGIC;
    SIGNAL S6586 : STD_LOGIC;
    SIGNAL S6587 : STD_LOGIC;
    SIGNAL S6588 : STD_LOGIC;
    SIGNAL S6589 : STD_LOGIC;
    SIGNAL S6590 : STD_LOGIC;
    SIGNAL S6591 : STD_LOGIC;
    SIGNAL S6592 : STD_LOGIC;
    SIGNAL S6593 : STD_LOGIC;
    SIGNAL S6594 : STD_LOGIC;
    SIGNAL S6595 : STD_LOGIC;
    SIGNAL S6596 : STD_LOGIC;
    SIGNAL S6597 : STD_LOGIC;
    SIGNAL S6598 : STD_LOGIC;
    SIGNAL S6599 : STD_LOGIC;
    SIGNAL S6600 : STD_LOGIC;
    SIGNAL S6601 : STD_LOGIC;
    SIGNAL S6602 : STD_LOGIC;
    SIGNAL S6603 : STD_LOGIC;
    SIGNAL S6604 : STD_LOGIC;
    SIGNAL S6605 : STD_LOGIC;
    SIGNAL S6606 : STD_LOGIC;
    SIGNAL S6607 : STD_LOGIC;
    SIGNAL S6608 : STD_LOGIC;
    SIGNAL S6609 : STD_LOGIC;
    SIGNAL S6610 : STD_LOGIC;
    SIGNAL S6611 : STD_LOGIC;
    SIGNAL S6612 : STD_LOGIC;
    SIGNAL S6613 : STD_LOGIC;
    SIGNAL S6614 : STD_LOGIC;
    SIGNAL S6615 : STD_LOGIC;
    SIGNAL S6616 : STD_LOGIC;
    SIGNAL S6617 : STD_LOGIC;
    SIGNAL S6618 : STD_LOGIC;
    SIGNAL S6619 : STD_LOGIC;
    SIGNAL S6620 : STD_LOGIC;
    SIGNAL S6621 : STD_LOGIC;
    SIGNAL S6622 : STD_LOGIC;
    SIGNAL S6623 : STD_LOGIC;
    SIGNAL S6624 : STD_LOGIC;
    SIGNAL S6625 : STD_LOGIC;
    SIGNAL S6626 : STD_LOGIC;
    SIGNAL S6627 : STD_LOGIC;
    SIGNAL S6628 : STD_LOGIC;
    SIGNAL S6629 : STD_LOGIC;
    SIGNAL S6630 : STD_LOGIC;
    SIGNAL S6631 : STD_LOGIC;
    SIGNAL S6632 : STD_LOGIC;
    SIGNAL S6633 : STD_LOGIC;
    SIGNAL S6634 : STD_LOGIC;
    SIGNAL S6635 : STD_LOGIC;
    SIGNAL S6636 : STD_LOGIC;
    SIGNAL S6637 : STD_LOGIC;
    SIGNAL S6638 : STD_LOGIC;
    SIGNAL S6639 : STD_LOGIC;
    SIGNAL S6640 : STD_LOGIC;
    SIGNAL S6641 : STD_LOGIC;
    SIGNAL S6642 : STD_LOGIC;
    SIGNAL S6643 : STD_LOGIC;
    SIGNAL S6644 : STD_LOGIC;
    SIGNAL S6645 : STD_LOGIC;
    SIGNAL S6646 : STD_LOGIC;
    SIGNAL S6647 : STD_LOGIC;
    SIGNAL S6648 : STD_LOGIC;
    SIGNAL S6649 : STD_LOGIC;
    SIGNAL S6650 : STD_LOGIC;
    SIGNAL S6651 : STD_LOGIC;
    SIGNAL S6652 : STD_LOGIC;
    SIGNAL S6653 : STD_LOGIC;
    SIGNAL S6654 : STD_LOGIC;
    SIGNAL S6655 : STD_LOGIC;
    SIGNAL S6656 : STD_LOGIC;
    SIGNAL S6657 : STD_LOGIC;
    SIGNAL S6658 : STD_LOGIC;
    SIGNAL S6659 : STD_LOGIC;
    SIGNAL S6660 : STD_LOGIC;
    SIGNAL S6661 : STD_LOGIC;
    SIGNAL S6662 : STD_LOGIC;
    SIGNAL S6663 : STD_LOGIC;
    SIGNAL S6664 : STD_LOGIC;
    SIGNAL S6665 : STD_LOGIC;
    SIGNAL S6666 : STD_LOGIC;
    SIGNAL S6667 : STD_LOGIC;
    SIGNAL S6668 : STD_LOGIC;
    SIGNAL S6669 : STD_LOGIC;
    SIGNAL S6670 : STD_LOGIC;
    SIGNAL S6671 : STD_LOGIC;
    SIGNAL S6672 : STD_LOGIC;
    SIGNAL S6673 : STD_LOGIC;
    SIGNAL S6674 : STD_LOGIC;
    SIGNAL S6675 : STD_LOGIC;
    SIGNAL S6676 : STD_LOGIC;
    SIGNAL S6677 : STD_LOGIC;
    SIGNAL S6678 : STD_LOGIC;
    SIGNAL S6679 : STD_LOGIC;
    SIGNAL S6680 : STD_LOGIC;
    SIGNAL S6681 : STD_LOGIC;
    SIGNAL S6682 : STD_LOGIC;
    SIGNAL S6683 : STD_LOGIC;
    SIGNAL S6684 : STD_LOGIC;
    SIGNAL S6685 : STD_LOGIC;
    SIGNAL S6686 : STD_LOGIC;
    SIGNAL S6687 : STD_LOGIC;
    SIGNAL S6688 : STD_LOGIC;
    SIGNAL S6689 : STD_LOGIC;
    SIGNAL S6690 : STD_LOGIC;
    SIGNAL S6691 : STD_LOGIC;
    SIGNAL S6692 : STD_LOGIC;
    SIGNAL S6693 : STD_LOGIC;
    SIGNAL S6694 : STD_LOGIC;
    SIGNAL S6695 : STD_LOGIC;
    SIGNAL S6696 : STD_LOGIC;
    SIGNAL S6697 : STD_LOGIC;
    SIGNAL S6698 : STD_LOGIC;
    SIGNAL S6699 : STD_LOGIC;
    SIGNAL S6700 : STD_LOGIC;
    SIGNAL S6701 : STD_LOGIC;
    SIGNAL S6702 : STD_LOGIC;
    SIGNAL S6703 : STD_LOGIC;
    SIGNAL S6704 : STD_LOGIC;
    SIGNAL S6705 : STD_LOGIC;
    SIGNAL S6706 : STD_LOGIC;
    SIGNAL S6707 : STD_LOGIC;
    SIGNAL S6708 : STD_LOGIC;
    SIGNAL S6709 : STD_LOGIC;
    SIGNAL S6710 : STD_LOGIC;
    SIGNAL S6711 : STD_LOGIC;
    SIGNAL S6712 : STD_LOGIC;
    SIGNAL S6713 : STD_LOGIC;
    SIGNAL S6714 : STD_LOGIC;
    SIGNAL S6715 : STD_LOGIC;
    SIGNAL S6716 : STD_LOGIC;
    SIGNAL S6717 : STD_LOGIC;
    SIGNAL S6718 : STD_LOGIC;
    SIGNAL S6719 : STD_LOGIC;
    SIGNAL S6720 : STD_LOGIC;
    SIGNAL S6721 : STD_LOGIC;
    SIGNAL S6722 : STD_LOGIC;
    SIGNAL S6723 : STD_LOGIC;
    SIGNAL S6724 : STD_LOGIC;
    SIGNAL S6725 : STD_LOGIC;
    SIGNAL S6726 : STD_LOGIC;
    SIGNAL S6727 : STD_LOGIC;
    SIGNAL S6728 : STD_LOGIC;
    SIGNAL S6729 : STD_LOGIC;
    SIGNAL S6730 : STD_LOGIC;
    SIGNAL S6731 : STD_LOGIC;
    SIGNAL S6732 : STD_LOGIC;
    SIGNAL S6733 : STD_LOGIC;
    SIGNAL S6734 : STD_LOGIC;
    SIGNAL S6735 : STD_LOGIC;
    SIGNAL S6736 : STD_LOGIC;
    SIGNAL S6737 : STD_LOGIC;
    SIGNAL S6738 : STD_LOGIC;
    SIGNAL S6739 : STD_LOGIC;
    SIGNAL S6740 : STD_LOGIC;
    SIGNAL S6741 : STD_LOGIC;
    SIGNAL S6742 : STD_LOGIC;
    SIGNAL S6743 : STD_LOGIC;
    SIGNAL S6744 : STD_LOGIC;
    SIGNAL S6745 : STD_LOGIC;
    SIGNAL S6746 : STD_LOGIC;
    SIGNAL S6747 : STD_LOGIC;
    SIGNAL S6748 : STD_LOGIC;
    SIGNAL S6749 : STD_LOGIC;
    SIGNAL S6750 : STD_LOGIC;
    SIGNAL S6751 : STD_LOGIC;
    SIGNAL S6752 : STD_LOGIC;
    SIGNAL S6753 : STD_LOGIC;
    SIGNAL S6754 : STD_LOGIC;
    SIGNAL S6755 : STD_LOGIC;
    SIGNAL S6756 : STD_LOGIC;
    SIGNAL S6757 : STD_LOGIC;
    SIGNAL S6758 : STD_LOGIC;
    SIGNAL S6759 : STD_LOGIC;
    SIGNAL S6760 : STD_LOGIC;
    SIGNAL S6761 : STD_LOGIC;
    SIGNAL S6762 : STD_LOGIC;
    SIGNAL S6763 : STD_LOGIC;
    SIGNAL S6764 : STD_LOGIC;
    SIGNAL S6765 : STD_LOGIC;
    SIGNAL S6766 : STD_LOGIC;
    SIGNAL S6767 : STD_LOGIC;
    SIGNAL S6768 : STD_LOGIC;
    SIGNAL S6769 : STD_LOGIC;
    SIGNAL S6770 : STD_LOGIC;
    SIGNAL S6771 : STD_LOGIC;
    SIGNAL S6772 : STD_LOGIC;
    SIGNAL S6773 : STD_LOGIC;
    SIGNAL S6774 : STD_LOGIC;
    SIGNAL S6775 : STD_LOGIC;
    SIGNAL S6776 : STD_LOGIC;
    SIGNAL S6777 : STD_LOGIC;
    SIGNAL S6778 : STD_LOGIC;
    SIGNAL S6779 : STD_LOGIC;
    SIGNAL S6780 : STD_LOGIC;
    SIGNAL S6781 : STD_LOGIC;
    SIGNAL S6782 : STD_LOGIC;
    SIGNAL S6783 : STD_LOGIC;
    SIGNAL S6784 : STD_LOGIC;
    SIGNAL S6785 : STD_LOGIC;
    SIGNAL S6786 : STD_LOGIC;
    SIGNAL S6787 : STD_LOGIC;
    SIGNAL S6788 : STD_LOGIC;
    SIGNAL S6789 : STD_LOGIC;
    SIGNAL S6790 : STD_LOGIC;
    SIGNAL S6791 : STD_LOGIC;
    SIGNAL S6792 : STD_LOGIC;
    SIGNAL S6793 : STD_LOGIC;
    SIGNAL S6794 : STD_LOGIC;
    SIGNAL S6795 : STD_LOGIC;
    SIGNAL S6796 : STD_LOGIC;
    SIGNAL S6797 : STD_LOGIC;
    SIGNAL S6798 : STD_LOGIC;
    SIGNAL S6799 : STD_LOGIC;
    SIGNAL S6800 : STD_LOGIC;
    SIGNAL S6801 : STD_LOGIC;
    SIGNAL S6802 : STD_LOGIC;
    SIGNAL S6803 : STD_LOGIC;
    SIGNAL S6804 : STD_LOGIC;
    SIGNAL S6805 : STD_LOGIC;
    SIGNAL S6806 : STD_LOGIC;
    SIGNAL S6807 : STD_LOGIC;
    SIGNAL S6808 : STD_LOGIC;
    SIGNAL S6809 : STD_LOGIC;
    SIGNAL S6810 : STD_LOGIC;
    SIGNAL S6811 : STD_LOGIC;
    SIGNAL S6812 : STD_LOGIC;
    SIGNAL S6813 : STD_LOGIC;
    SIGNAL S6814 : STD_LOGIC;
    SIGNAL S6815 : STD_LOGIC;
    SIGNAL S6816 : STD_LOGIC;
    SIGNAL S6817 : STD_LOGIC;
    SIGNAL S6818 : STD_LOGIC;
    SIGNAL S6819 : STD_LOGIC;
    SIGNAL S6820 : STD_LOGIC;
    SIGNAL S6821 : STD_LOGIC;
    SIGNAL S6822 : STD_LOGIC;
    SIGNAL S6823 : STD_LOGIC;
    SIGNAL S6824 : STD_LOGIC;
    SIGNAL S6825 : STD_LOGIC;
    SIGNAL S6826 : STD_LOGIC;
    SIGNAL S6827 : STD_LOGIC;
    SIGNAL S6828 : STD_LOGIC;
    SIGNAL S6829 : STD_LOGIC;
    SIGNAL S6830 : STD_LOGIC;
    SIGNAL S6831 : STD_LOGIC;
    SIGNAL S6832 : STD_LOGIC;
    SIGNAL S6833 : STD_LOGIC;
    SIGNAL S6834 : STD_LOGIC;
    SIGNAL S6835 : STD_LOGIC;
    SIGNAL S6836 : STD_LOGIC;
    SIGNAL S6837 : STD_LOGIC;
    SIGNAL S6838 : STD_LOGIC;
    SIGNAL S6839 : STD_LOGIC;
    SIGNAL S6840 : STD_LOGIC;
    SIGNAL S6841 : STD_LOGIC;
    SIGNAL S6842 : STD_LOGIC;
    SIGNAL S6843 : STD_LOGIC;
    SIGNAL S6844 : STD_LOGIC;
    SIGNAL S6845 : STD_LOGIC;
    SIGNAL S6846 : STD_LOGIC;
    SIGNAL S6847 : STD_LOGIC;
    SIGNAL S6848 : STD_LOGIC;
    SIGNAL S6849 : STD_LOGIC;
    SIGNAL S6850 : STD_LOGIC;
    SIGNAL S6851 : STD_LOGIC;
    SIGNAL S6852 : STD_LOGIC;
    SIGNAL S6853 : STD_LOGIC;
    SIGNAL S6854 : STD_LOGIC;
    SIGNAL S6855 : STD_LOGIC;
    SIGNAL S6856 : STD_LOGIC;
    SIGNAL S6857 : STD_LOGIC;
    SIGNAL S6858 : STD_LOGIC;
    SIGNAL S6859 : STD_LOGIC;
    SIGNAL S6860 : STD_LOGIC;
    SIGNAL S6861 : STD_LOGIC;
    SIGNAL S6862 : STD_LOGIC;
    SIGNAL S6863 : STD_LOGIC;
    SIGNAL S6864 : STD_LOGIC;
    SIGNAL S6865 : STD_LOGIC;
    SIGNAL S6866 : STD_LOGIC;
    SIGNAL S6867 : STD_LOGIC;
    SIGNAL S6868 : STD_LOGIC;
    SIGNAL S6869 : STD_LOGIC;
    SIGNAL S6870 : STD_LOGIC;
    SIGNAL S6871 : STD_LOGIC;
    SIGNAL S6872 : STD_LOGIC;
    SIGNAL S6873 : STD_LOGIC;
    SIGNAL S6874 : STD_LOGIC;
    SIGNAL S6875 : STD_LOGIC;
    SIGNAL S6876 : STD_LOGIC;
    SIGNAL S6877 : STD_LOGIC;
    SIGNAL S6878 : STD_LOGIC;
    SIGNAL S6879 : STD_LOGIC;
    SIGNAL S6880 : STD_LOGIC;
    SIGNAL S6881 : STD_LOGIC;
    SIGNAL S6882 : STD_LOGIC;
    SIGNAL S6883 : STD_LOGIC;
    SIGNAL S6884 : STD_LOGIC;
    SIGNAL S6885 : STD_LOGIC;
    SIGNAL S6886 : STD_LOGIC;
    SIGNAL S6887 : STD_LOGIC;
    SIGNAL S6888 : STD_LOGIC;
    SIGNAL S6889 : STD_LOGIC;
    SIGNAL S6890 : STD_LOGIC;
    SIGNAL S6891 : STD_LOGIC;
    SIGNAL S6892 : STD_LOGIC;
    SIGNAL S6893 : STD_LOGIC;
    SIGNAL S6894 : STD_LOGIC;
    SIGNAL S6895 : STD_LOGIC;
    SIGNAL S6896 : STD_LOGIC;
    SIGNAL S6897 : STD_LOGIC;
    SIGNAL S6898 : STD_LOGIC;
    SIGNAL S6899 : STD_LOGIC;
    SIGNAL S6900 : STD_LOGIC;
    SIGNAL S6901 : STD_LOGIC;
    SIGNAL S6902 : STD_LOGIC;
    SIGNAL S6903 : STD_LOGIC;
    SIGNAL S6904 : STD_LOGIC;
    SIGNAL S6905 : STD_LOGIC;
    SIGNAL S6906 : STD_LOGIC;
    SIGNAL S6907 : STD_LOGIC;
    SIGNAL S6908 : STD_LOGIC;
    SIGNAL S6909 : STD_LOGIC;
    SIGNAL S6910 : STD_LOGIC;
    SIGNAL S6911 : STD_LOGIC;
    SIGNAL S6912 : STD_LOGIC;
    SIGNAL S6913 : STD_LOGIC;
    SIGNAL S6914 : STD_LOGIC;
    SIGNAL S6915 : STD_LOGIC;
    SIGNAL S6916 : STD_LOGIC;
    SIGNAL S6917 : STD_LOGIC;
    SIGNAL S6918 : STD_LOGIC;
    SIGNAL S6919 : STD_LOGIC;
    SIGNAL S6920 : STD_LOGIC;
    SIGNAL S6921 : STD_LOGIC;
    SIGNAL S6922 : STD_LOGIC;
    SIGNAL S6923 : STD_LOGIC;
    SIGNAL S6924 : STD_LOGIC;
    SIGNAL S6925 : STD_LOGIC;
    SIGNAL S6926 : STD_LOGIC;
    SIGNAL S6927 : STD_LOGIC;
    SIGNAL S6928 : STD_LOGIC;
    SIGNAL S6929 : STD_LOGIC;
    SIGNAL S6930 : STD_LOGIC;
    SIGNAL S6931 : STD_LOGIC;
    SIGNAL S6932 : STD_LOGIC;
    SIGNAL S6933 : STD_LOGIC;
    SIGNAL S6934 : STD_LOGIC;
    SIGNAL S6935 : STD_LOGIC;
    SIGNAL S6936 : STD_LOGIC;
    SIGNAL S6937 : STD_LOGIC;
    SIGNAL S6938 : STD_LOGIC;
    SIGNAL S6939 : STD_LOGIC;
    SIGNAL S6940 : STD_LOGIC;
    SIGNAL S6941 : STD_LOGIC;
    SIGNAL S6942 : STD_LOGIC;
    SIGNAL S6943 : STD_LOGIC;
    SIGNAL S6944 : STD_LOGIC;
    SIGNAL S6945 : STD_LOGIC;
    SIGNAL S6946 : STD_LOGIC;
    SIGNAL S6947 : STD_LOGIC;
    SIGNAL S6948 : STD_LOGIC;
    SIGNAL S6949 : STD_LOGIC;
    SIGNAL S6950 : STD_LOGIC;
    SIGNAL S6951 : STD_LOGIC;
    SIGNAL S6952 : STD_LOGIC;
    SIGNAL S6953 : STD_LOGIC;
    SIGNAL S6954 : STD_LOGIC;
    SIGNAL S6955 : STD_LOGIC;
    SIGNAL S6956 : STD_LOGIC;
    SIGNAL S6957 : STD_LOGIC;
    SIGNAL S6958 : STD_LOGIC;
    SIGNAL S6959 : STD_LOGIC;
    SIGNAL S6960 : STD_LOGIC;
    SIGNAL S6961 : STD_LOGIC;
    SIGNAL S6962 : STD_LOGIC;
    SIGNAL S6963 : STD_LOGIC;
    SIGNAL S6964 : STD_LOGIC;
    SIGNAL S6965 : STD_LOGIC;
    SIGNAL S6966 : STD_LOGIC;
    SIGNAL S6967 : STD_LOGIC;
    SIGNAL S6968 : STD_LOGIC;
    SIGNAL S6969 : STD_LOGIC;
    SIGNAL S6970 : STD_LOGIC;
    SIGNAL S6971 : STD_LOGIC;
    SIGNAL S6972 : STD_LOGIC;
    SIGNAL S6973 : STD_LOGIC;
    SIGNAL S6974 : STD_LOGIC;
    SIGNAL S6975 : STD_LOGIC;
    SIGNAL S6976 : STD_LOGIC;
    SIGNAL S6977 : STD_LOGIC;
    SIGNAL S6978 : STD_LOGIC;
    SIGNAL S6979 : STD_LOGIC;
    SIGNAL S6980 : STD_LOGIC;
    SIGNAL S6981 : STD_LOGIC;
    SIGNAL S6982 : STD_LOGIC;
    SIGNAL S6983 : STD_LOGIC;
    SIGNAL S6984 : STD_LOGIC;
    SIGNAL S6985 : STD_LOGIC;
    SIGNAL S6986 : STD_LOGIC;
    SIGNAL S6987 : STD_LOGIC;
    SIGNAL S6988 : STD_LOGIC;
    SIGNAL S6989 : STD_LOGIC;
    SIGNAL S6990 : STD_LOGIC;
    SIGNAL S6991 : STD_LOGIC;
    SIGNAL S6992 : STD_LOGIC;
    SIGNAL S6993 : STD_LOGIC;
    SIGNAL S6994 : STD_LOGIC;
    SIGNAL S6995 : STD_LOGIC;
    SIGNAL S6996 : STD_LOGIC;
    SIGNAL S6997 : STD_LOGIC;
    SIGNAL S6998 : STD_LOGIC;
    SIGNAL S6999 : STD_LOGIC;
    SIGNAL S7000 : STD_LOGIC;
    SIGNAL S7001 : STD_LOGIC;
    SIGNAL S7002 : STD_LOGIC;
    SIGNAL S7003 : STD_LOGIC;
    SIGNAL S7004 : STD_LOGIC;
    SIGNAL S7005 : STD_LOGIC;
    SIGNAL S7006 : STD_LOGIC;
    SIGNAL S7007 : STD_LOGIC;
    SIGNAL S7008 : STD_LOGIC;
    SIGNAL S7009 : STD_LOGIC;
    SIGNAL S7010 : STD_LOGIC;
    SIGNAL S7011 : STD_LOGIC;
    SIGNAL S7012 : STD_LOGIC;
    SIGNAL S7013 : STD_LOGIC;
    SIGNAL S7014 : STD_LOGIC;
    SIGNAL S7015 : STD_LOGIC;
    SIGNAL S7016 : STD_LOGIC;
    SIGNAL S7017 : STD_LOGIC;
    SIGNAL S7018 : STD_LOGIC;
    SIGNAL S7019 : STD_LOGIC;
    SIGNAL S7020 : STD_LOGIC;
    SIGNAL S7021 : STD_LOGIC;
    SIGNAL S7022 : STD_LOGIC;
    SIGNAL S7023 : STD_LOGIC;
    SIGNAL S7024 : STD_LOGIC;
    SIGNAL S7025 : STD_LOGIC;
    SIGNAL S7026 : STD_LOGIC;
    SIGNAL S7027 : STD_LOGIC;
    SIGNAL S7028 : STD_LOGIC;
    SIGNAL S7029 : STD_LOGIC;
    SIGNAL S7030 : STD_LOGIC;
    SIGNAL S7031 : STD_LOGIC;
    SIGNAL S7032 : STD_LOGIC;
    SIGNAL S7033 : STD_LOGIC;
    SIGNAL S7034 : STD_LOGIC;
    SIGNAL S7035 : STD_LOGIC;
    SIGNAL S7036 : STD_LOGIC;
    SIGNAL S7037 : STD_LOGIC;
    SIGNAL S7038 : STD_LOGIC;
    SIGNAL S7039 : STD_LOGIC;
    SIGNAL S7040 : STD_LOGIC;
    SIGNAL S7041 : STD_LOGIC;
    SIGNAL S7042 : STD_LOGIC;
    SIGNAL S7043 : STD_LOGIC;
    SIGNAL S7044 : STD_LOGIC;
    SIGNAL S7045 : STD_LOGIC;
    SIGNAL S7046 : STD_LOGIC;
    SIGNAL S7047 : STD_LOGIC;
    SIGNAL S7048 : STD_LOGIC;
    SIGNAL S7049 : STD_LOGIC;
    SIGNAL S7050 : STD_LOGIC;
    SIGNAL S7051 : STD_LOGIC;
    SIGNAL S7052 : STD_LOGIC;
    SIGNAL S7053 : STD_LOGIC;
    SIGNAL S7054 : STD_LOGIC;
    SIGNAL S7055 : STD_LOGIC;
    SIGNAL S7056 : STD_LOGIC;
    SIGNAL S7057 : STD_LOGIC;
    SIGNAL S7058 : STD_LOGIC;
    SIGNAL S7059 : STD_LOGIC;
    SIGNAL S7060 : STD_LOGIC;
    SIGNAL S7061 : STD_LOGIC;
    SIGNAL S7062 : STD_LOGIC;
    SIGNAL S7063 : STD_LOGIC;
    SIGNAL S7064 : STD_LOGIC;
    SIGNAL S7065 : STD_LOGIC;
    SIGNAL S7066 : STD_LOGIC;
    SIGNAL S7067 : STD_LOGIC;
    SIGNAL S7068 : STD_LOGIC;
    SIGNAL S7069 : STD_LOGIC;
    SIGNAL S7070 : STD_LOGIC;
    SIGNAL S7071 : STD_LOGIC;
    SIGNAL S7072 : STD_LOGIC;
    SIGNAL S7073 : STD_LOGIC;
    SIGNAL S7074 : STD_LOGIC;
    SIGNAL S7075 : STD_LOGIC;
    SIGNAL S7076 : STD_LOGIC;
    SIGNAL S7077 : STD_LOGIC;
    SIGNAL S7078 : STD_LOGIC;
    SIGNAL S7079 : STD_LOGIC;
    SIGNAL S7080 : STD_LOGIC;
    SIGNAL S7081 : STD_LOGIC;
    SIGNAL S7082 : STD_LOGIC;
    SIGNAL S7083 : STD_LOGIC;
    SIGNAL S7084 : STD_LOGIC;
    SIGNAL S7085 : STD_LOGIC;
    SIGNAL S7086 : STD_LOGIC;
    SIGNAL S7087 : STD_LOGIC;
    SIGNAL S7088 : STD_LOGIC;
    SIGNAL S7089 : STD_LOGIC;
    SIGNAL S7090 : STD_LOGIC;
    SIGNAL S7091 : STD_LOGIC;
    SIGNAL S7092 : STD_LOGIC;
    SIGNAL S7093 : STD_LOGIC;
    SIGNAL S7094 : STD_LOGIC;
    SIGNAL S7095 : STD_LOGIC;
    SIGNAL S7096 : STD_LOGIC;
    SIGNAL S7097 : STD_LOGIC;
    SIGNAL S7098 : STD_LOGIC;
    SIGNAL S7099 : STD_LOGIC;
    SIGNAL S7100 : STD_LOGIC;
    SIGNAL S7101 : STD_LOGIC;
    SIGNAL S7102 : STD_LOGIC;
    SIGNAL S7103 : STD_LOGIC;
    SIGNAL S7104 : STD_LOGIC;
    SIGNAL S7105 : STD_LOGIC;
    SIGNAL S7106 : STD_LOGIC;
    SIGNAL S7107 : STD_LOGIC;
    SIGNAL S7108 : STD_LOGIC;
    SIGNAL S7109 : STD_LOGIC;
    SIGNAL S7110 : STD_LOGIC;
    SIGNAL S7111 : STD_LOGIC;
    SIGNAL S7112 : STD_LOGIC;
    SIGNAL S7113 : STD_LOGIC;
    SIGNAL S7114 : STD_LOGIC;
    SIGNAL S7115 : STD_LOGIC;
    SIGNAL S7116 : STD_LOGIC;
    SIGNAL S7117 : STD_LOGIC;
    SIGNAL S7118 : STD_LOGIC;
    SIGNAL S7119 : STD_LOGIC;
    SIGNAL S7120 : STD_LOGIC;
    SIGNAL S7121 : STD_LOGIC;
    SIGNAL S7122 : STD_LOGIC;
    SIGNAL S7123 : STD_LOGIC;
    SIGNAL S7124 : STD_LOGIC;
    SIGNAL S7125 : STD_LOGIC;
    SIGNAL S7126 : STD_LOGIC;
    SIGNAL S7127 : STD_LOGIC;
    SIGNAL S7128 : STD_LOGIC;
    SIGNAL S7129 : STD_LOGIC;
    SIGNAL S7130 : STD_LOGIC;
    SIGNAL S7131 : STD_LOGIC;
    SIGNAL S7132 : STD_LOGIC;
    SIGNAL S7133 : STD_LOGIC;
    SIGNAL S7134 : STD_LOGIC;
    SIGNAL S7135 : STD_LOGIC;
    SIGNAL S7136 : STD_LOGIC;
    SIGNAL S7137 : STD_LOGIC;
    SIGNAL S7138 : STD_LOGIC;
    SIGNAL S7139 : STD_LOGIC;
    SIGNAL S7140 : STD_LOGIC;
    SIGNAL S7141 : STD_LOGIC;
    SIGNAL S7142 : STD_LOGIC;
    SIGNAL S7143 : STD_LOGIC;
    SIGNAL S7144 : STD_LOGIC;
    SIGNAL S7145 : STD_LOGIC;
    SIGNAL S7146 : STD_LOGIC;
    SIGNAL S7147 : STD_LOGIC;
    SIGNAL S7148 : STD_LOGIC;
    SIGNAL S7149 : STD_LOGIC;
    SIGNAL S7150 : STD_LOGIC;
    SIGNAL S7151 : STD_LOGIC;
    SIGNAL S7152 : STD_LOGIC;
    SIGNAL S7153 : STD_LOGIC;
    SIGNAL S7154 : STD_LOGIC;
    SIGNAL S7155 : STD_LOGIC;
    SIGNAL S7156 : STD_LOGIC;
    SIGNAL S7157 : STD_LOGIC;
    SIGNAL S7158 : STD_LOGIC;
    SIGNAL S7159 : STD_LOGIC;
    SIGNAL S7160 : STD_LOGIC;
    SIGNAL S7161 : STD_LOGIC;
    SIGNAL S7162 : STD_LOGIC;
    SIGNAL S7163 : STD_LOGIC;
    SIGNAL S7164 : STD_LOGIC;
    SIGNAL S7165 : STD_LOGIC;
    SIGNAL S7166 : STD_LOGIC;
    SIGNAL S7167 : STD_LOGIC;
    SIGNAL S7168 : STD_LOGIC;
    SIGNAL S7169 : STD_LOGIC;
    SIGNAL S7170 : STD_LOGIC;
    SIGNAL S7171 : STD_LOGIC;
    SIGNAL S7172 : STD_LOGIC;
    SIGNAL S7173 : STD_LOGIC;
    SIGNAL S7174 : STD_LOGIC;
    SIGNAL S7175 : STD_LOGIC;
    SIGNAL S7176 : STD_LOGIC;
    SIGNAL S7177 : STD_LOGIC;
    SIGNAL S7178 : STD_LOGIC;
    SIGNAL S7179 : STD_LOGIC;
    SIGNAL S7180 : STD_LOGIC;
    SIGNAL S7181 : STD_LOGIC;
    SIGNAL S7182 : STD_LOGIC;
    SIGNAL S7183 : STD_LOGIC;
    SIGNAL S7184 : STD_LOGIC;
    SIGNAL S7185 : STD_LOGIC;
    SIGNAL S7186 : STD_LOGIC;
    SIGNAL S7187 : STD_LOGIC;
    SIGNAL S7188 : STD_LOGIC;
    SIGNAL S7189 : STD_LOGIC;
    SIGNAL S7190 : STD_LOGIC;
    SIGNAL S7191 : STD_LOGIC;
    SIGNAL S7192 : STD_LOGIC;
    SIGNAL S7193 : STD_LOGIC;
    SIGNAL S7194 : STD_LOGIC;
    SIGNAL S7195 : STD_LOGIC;
    SIGNAL S7196 : STD_LOGIC;
    SIGNAL S7197 : STD_LOGIC;
    SIGNAL S7198 : STD_LOGIC;
    SIGNAL S7199 : STD_LOGIC;
    SIGNAL S7200 : STD_LOGIC;
    SIGNAL S7201 : STD_LOGIC;
    SIGNAL S7202 : STD_LOGIC;
    SIGNAL S7203 : STD_LOGIC;
    SIGNAL S7204 : STD_LOGIC;
    SIGNAL S7205 : STD_LOGIC;
    SIGNAL S7206 : STD_LOGIC;
    SIGNAL S7207 : STD_LOGIC;
    SIGNAL S7208 : STD_LOGIC;
    SIGNAL S7209 : STD_LOGIC;
    SIGNAL S7210 : STD_LOGIC;
    SIGNAL S7211 : STD_LOGIC;
    SIGNAL S7212 : STD_LOGIC;
    SIGNAL S7213 : STD_LOGIC;
    SIGNAL S7214 : STD_LOGIC;
    SIGNAL S7215 : STD_LOGIC;
    SIGNAL S7216 : STD_LOGIC;
    SIGNAL S7217 : STD_LOGIC;
    SIGNAL S7218 : STD_LOGIC;
    SIGNAL S7219 : STD_LOGIC;
    SIGNAL S7220 : STD_LOGIC;
    SIGNAL S7221 : STD_LOGIC;
    SIGNAL S7222 : STD_LOGIC;
    SIGNAL S7223 : STD_LOGIC;
    SIGNAL S7224 : STD_LOGIC;
    SIGNAL S7225 : STD_LOGIC;
    SIGNAL S7226 : STD_LOGIC;
    SIGNAL S7227 : STD_LOGIC;
    SIGNAL S7228 : STD_LOGIC;
    SIGNAL S7229 : STD_LOGIC;
    SIGNAL S7230 : STD_LOGIC;
    SIGNAL S7231 : STD_LOGIC;
    SIGNAL S7232 : STD_LOGIC;
    SIGNAL S7233 : STD_LOGIC;
    SIGNAL S7234 : STD_LOGIC;
    SIGNAL S7235 : STD_LOGIC;
    SIGNAL S7236 : STD_LOGIC;
    SIGNAL S7237 : STD_LOGIC;
    SIGNAL S7238 : STD_LOGIC;
    SIGNAL S7239 : STD_LOGIC;
    SIGNAL S7240 : STD_LOGIC;
    SIGNAL S7241 : STD_LOGIC;
    SIGNAL S7242 : STD_LOGIC;
    SIGNAL S7243 : STD_LOGIC;
    SIGNAL S7244 : STD_LOGIC;
    SIGNAL S7245 : STD_LOGIC;
    SIGNAL S7246 : STD_LOGIC;
    SIGNAL S7247 : STD_LOGIC;
    SIGNAL S7248 : STD_LOGIC;
    SIGNAL S7249 : STD_LOGIC;
    SIGNAL S7250 : STD_LOGIC;
    SIGNAL S7251 : STD_LOGIC;
    SIGNAL S7252 : STD_LOGIC;
    SIGNAL S7253 : STD_LOGIC;
    SIGNAL S7254 : STD_LOGIC;
    SIGNAL S7255 : STD_LOGIC;
    SIGNAL S7256 : STD_LOGIC;
    SIGNAL S7257 : STD_LOGIC;
    SIGNAL S7258 : STD_LOGIC;
    SIGNAL S7259 : STD_LOGIC;
    SIGNAL S7260 : STD_LOGIC;
    SIGNAL S7261 : STD_LOGIC;
    SIGNAL S7262 : STD_LOGIC;
    SIGNAL S7263 : STD_LOGIC;
    SIGNAL S7264 : STD_LOGIC;
    SIGNAL S7265 : STD_LOGIC;
    SIGNAL S7266 : STD_LOGIC;
    SIGNAL S7267 : STD_LOGIC;
    SIGNAL S7268 : STD_LOGIC;
    SIGNAL S7269 : STD_LOGIC;
    SIGNAL S7270 : STD_LOGIC;
    SIGNAL S7271 : STD_LOGIC;
    SIGNAL S7272 : STD_LOGIC;
    SIGNAL S7273 : STD_LOGIC;
    SIGNAL S7274 : STD_LOGIC;
    SIGNAL S7275 : STD_LOGIC;
    SIGNAL S7276 : STD_LOGIC;
    SIGNAL S7277 : STD_LOGIC;
    SIGNAL S7278 : STD_LOGIC;
    SIGNAL S7279 : STD_LOGIC;
    SIGNAL S7280 : STD_LOGIC;
    SIGNAL S7281 : STD_LOGIC;
    SIGNAL S7282 : STD_LOGIC;
    SIGNAL S7283 : STD_LOGIC;
    SIGNAL S7284 : STD_LOGIC;
    SIGNAL S7285 : STD_LOGIC;
    SIGNAL S7286 : STD_LOGIC;
    SIGNAL S7287 : STD_LOGIC;
    SIGNAL S7288 : STD_LOGIC;
    SIGNAL S7289 : STD_LOGIC;
    SIGNAL S7290 : STD_LOGIC;
    SIGNAL S7291 : STD_LOGIC;
    SIGNAL S7292 : STD_LOGIC;
    SIGNAL S7293 : STD_LOGIC;
    SIGNAL S7294 : STD_LOGIC;
    SIGNAL S7295 : STD_LOGIC;
    SIGNAL S7296 : STD_LOGIC;
    SIGNAL S7297 : STD_LOGIC;
    SIGNAL S7298 : STD_LOGIC;
    SIGNAL S7299 : STD_LOGIC;
    SIGNAL S7300 : STD_LOGIC;
    SIGNAL S7301 : STD_LOGIC;
    SIGNAL S7302 : STD_LOGIC;
    SIGNAL S7303 : STD_LOGIC;
    SIGNAL S7304 : STD_LOGIC;
    SIGNAL S7305 : STD_LOGIC;
    SIGNAL S7306 : STD_LOGIC;
    SIGNAL S7307 : STD_LOGIC;
    SIGNAL S7308 : STD_LOGIC;
    SIGNAL S7309 : STD_LOGIC;
    SIGNAL S7310 : STD_LOGIC;
    SIGNAL S7311 : STD_LOGIC;
    SIGNAL S7312 : STD_LOGIC;
    SIGNAL S7313 : STD_LOGIC;
    SIGNAL S7314 : STD_LOGIC;
    SIGNAL S7315 : STD_LOGIC;
    SIGNAL S7316 : STD_LOGIC;
    SIGNAL S7317 : STD_LOGIC;
    SIGNAL S7318 : STD_LOGIC;
    SIGNAL S7319 : STD_LOGIC;
    SIGNAL S7320 : STD_LOGIC;
    SIGNAL S7321 : STD_LOGIC;
    SIGNAL S7322 : STD_LOGIC;
    SIGNAL S7323 : STD_LOGIC;
    SIGNAL S7324 : STD_LOGIC;
    SIGNAL S7325 : STD_LOGIC;
    SIGNAL S7326 : STD_LOGIC;
    SIGNAL S7327 : STD_LOGIC;
    SIGNAL S7328 : STD_LOGIC;
    SIGNAL S7329 : STD_LOGIC;
    SIGNAL S7330 : STD_LOGIC;
    SIGNAL S7331 : STD_LOGIC;
    SIGNAL S7332 : STD_LOGIC;
    SIGNAL S7333 : STD_LOGIC;
    SIGNAL S7334 : STD_LOGIC;
    SIGNAL S7335 : STD_LOGIC;
    SIGNAL S7336 : STD_LOGIC;
    SIGNAL S7337 : STD_LOGIC;
    SIGNAL S7338 : STD_LOGIC;
    SIGNAL S7339 : STD_LOGIC;
    SIGNAL S7340 : STD_LOGIC;
    SIGNAL S7341 : STD_LOGIC;
    SIGNAL S7342 : STD_LOGIC;
    SIGNAL S7343 : STD_LOGIC;
    SIGNAL S7344 : STD_LOGIC;
    SIGNAL S7345 : STD_LOGIC;
    SIGNAL S7346 : STD_LOGIC;
    SIGNAL S7347 : STD_LOGIC;
    SIGNAL S7348 : STD_LOGIC;
    SIGNAL S7349 : STD_LOGIC;
    SIGNAL S7350 : STD_LOGIC;
    SIGNAL S7351 : STD_LOGIC;
    SIGNAL S7352 : STD_LOGIC;
    SIGNAL S7353 : STD_LOGIC;
    SIGNAL S7354 : STD_LOGIC;
    SIGNAL S7355 : STD_LOGIC;
    SIGNAL S7356 : STD_LOGIC;
    SIGNAL S7357 : STD_LOGIC;
    SIGNAL S7358 : STD_LOGIC;
    SIGNAL S7359 : STD_LOGIC;
    SIGNAL S7360 : STD_LOGIC;
    SIGNAL S7361 : STD_LOGIC;
    SIGNAL S7362 : STD_LOGIC;
    SIGNAL S7363 : STD_LOGIC;
    SIGNAL S7364 : STD_LOGIC;
    SIGNAL S7365 : STD_LOGIC;
    SIGNAL S7366 : STD_LOGIC;
    SIGNAL S7367 : STD_LOGIC;
    SIGNAL S7368 : STD_LOGIC;
    SIGNAL S7369 : STD_LOGIC;
    SIGNAL S7370 : STD_LOGIC;
    SIGNAL S7371 : STD_LOGIC;
    SIGNAL S7372 : STD_LOGIC;
    SIGNAL S7373 : STD_LOGIC;
    SIGNAL S7374 : STD_LOGIC;
    SIGNAL S7375 : STD_LOGIC;
    SIGNAL S7376 : STD_LOGIC;
    SIGNAL S7377 : STD_LOGIC;
    SIGNAL S7378 : STD_LOGIC;
    SIGNAL S7379 : STD_LOGIC;
    SIGNAL S7380 : STD_LOGIC;
    SIGNAL S7381 : STD_LOGIC;
    SIGNAL S7382 : STD_LOGIC;
    SIGNAL S7383 : STD_LOGIC;
    SIGNAL S7384 : STD_LOGIC;
    SIGNAL S7385 : STD_LOGIC;
    SIGNAL S7386 : STD_LOGIC;
    SIGNAL S7387 : STD_LOGIC;
    SIGNAL S7388 : STD_LOGIC;
    SIGNAL S7389 : STD_LOGIC;
    SIGNAL S7390 : STD_LOGIC;
    SIGNAL S7391 : STD_LOGIC;
    SIGNAL S7392 : STD_LOGIC;
    SIGNAL S7393 : STD_LOGIC;
    SIGNAL S7394 : STD_LOGIC;
    SIGNAL S7395 : STD_LOGIC;
    SIGNAL S7396 : STD_LOGIC;
    SIGNAL S7397 : STD_LOGIC;
    SIGNAL S7398 : STD_LOGIC;
    SIGNAL S7399 : STD_LOGIC;
    SIGNAL S7400 : STD_LOGIC;
    SIGNAL S7401 : STD_LOGIC;
    SIGNAL S7402 : STD_LOGIC;
    SIGNAL S7403 : STD_LOGIC;
    SIGNAL S7404 : STD_LOGIC;
    SIGNAL S7405 : STD_LOGIC;
    SIGNAL S7406 : STD_LOGIC;
    SIGNAL S7407 : STD_LOGIC;
    SIGNAL S7408 : STD_LOGIC;
    SIGNAL S7409 : STD_LOGIC;
    SIGNAL S7410 : STD_LOGIC;
    SIGNAL S7411 : STD_LOGIC;
    SIGNAL S7412 : STD_LOGIC;
    SIGNAL S7413 : STD_LOGIC;
    SIGNAL S7414 : STD_LOGIC;
    SIGNAL S7415 : STD_LOGIC;
    SIGNAL S7416 : STD_LOGIC;
    SIGNAL S7417 : STD_LOGIC;
    SIGNAL S7418 : STD_LOGIC;
    SIGNAL S7419 : STD_LOGIC;
    SIGNAL S7420 : STD_LOGIC;
    SIGNAL S7421 : STD_LOGIC;
    SIGNAL S7422 : STD_LOGIC;
    SIGNAL S7423 : STD_LOGIC;
    SIGNAL S7424 : STD_LOGIC;
    SIGNAL S7425 : STD_LOGIC;
    SIGNAL S7426 : STD_LOGIC;
    SIGNAL S7427 : STD_LOGIC;
    SIGNAL S7428 : STD_LOGIC;
    SIGNAL S7429 : STD_LOGIC;
    SIGNAL S7430 : STD_LOGIC;
    SIGNAL S7431 : STD_LOGIC;
    SIGNAL S7432 : STD_LOGIC;
    SIGNAL S7433 : STD_LOGIC;
    SIGNAL S7434 : STD_LOGIC;
    SIGNAL S7435 : STD_LOGIC;
    SIGNAL S7436 : STD_LOGIC;
    SIGNAL S7437 : STD_LOGIC;
    SIGNAL S7438 : STD_LOGIC;
    SIGNAL S7439 : STD_LOGIC;
    SIGNAL S7440 : STD_LOGIC;
    SIGNAL S7441 : STD_LOGIC;
    SIGNAL S7442 : STD_LOGIC;
    SIGNAL S7443 : STD_LOGIC;
    SIGNAL S7444 : STD_LOGIC;
    SIGNAL S7445 : STD_LOGIC;
    SIGNAL S7446 : STD_LOGIC;
    SIGNAL S7447 : STD_LOGIC;
    SIGNAL S7448 : STD_LOGIC;
    SIGNAL S7449 : STD_LOGIC;
    SIGNAL S7450 : STD_LOGIC;
    SIGNAL S7451 : STD_LOGIC;
    SIGNAL S7452 : STD_LOGIC;
    SIGNAL S7453 : STD_LOGIC;
    SIGNAL S7454 : STD_LOGIC;
    SIGNAL S7455 : STD_LOGIC;
    SIGNAL S7456 : STD_LOGIC;
    SIGNAL S7457 : STD_LOGIC;
    SIGNAL S7458 : STD_LOGIC;
    SIGNAL S7459 : STD_LOGIC;
    SIGNAL S7460 : STD_LOGIC;
    SIGNAL S7461 : STD_LOGIC;
    SIGNAL S7462 : STD_LOGIC;
    SIGNAL S7463 : STD_LOGIC;
    SIGNAL S7464 : STD_LOGIC;
    SIGNAL S7465 : STD_LOGIC;
    SIGNAL S7466 : STD_LOGIC;
    SIGNAL S7467 : STD_LOGIC;
    SIGNAL S7468 : STD_LOGIC;
    SIGNAL S7469 : STD_LOGIC;
    SIGNAL S7470 : STD_LOGIC;
    SIGNAL S7471 : STD_LOGIC;
    SIGNAL S7472 : STD_LOGIC;
    SIGNAL S7473 : STD_LOGIC;
    SIGNAL S7474 : STD_LOGIC;
    SIGNAL S7475 : STD_LOGIC;
    SIGNAL S7476 : STD_LOGIC;
    SIGNAL S7477 : STD_LOGIC;
    SIGNAL S7478 : STD_LOGIC;
    SIGNAL S7479 : STD_LOGIC;
    SIGNAL S7480 : STD_LOGIC;
    SIGNAL S7481 : STD_LOGIC;
    SIGNAL S7482 : STD_LOGIC;
    SIGNAL S7483 : STD_LOGIC;
    SIGNAL S7484 : STD_LOGIC;
    SIGNAL S7485 : STD_LOGIC;
    SIGNAL S7486 : STD_LOGIC;
    SIGNAL S7487 : STD_LOGIC;
    SIGNAL S7488 : STD_LOGIC;
    SIGNAL S7489 : STD_LOGIC;
    SIGNAL S7490 : STD_LOGIC;
    SIGNAL S7491 : STD_LOGIC;
    SIGNAL S7492 : STD_LOGIC;
    SIGNAL S7493 : STD_LOGIC;
    SIGNAL S7494 : STD_LOGIC;
    SIGNAL S7495 : STD_LOGIC;
    SIGNAL S7496 : STD_LOGIC;
    SIGNAL S7497 : STD_LOGIC;
    SIGNAL S7498 : STD_LOGIC;
    SIGNAL S7499 : STD_LOGIC;
    SIGNAL S7500 : STD_LOGIC;
    SIGNAL S7501 : STD_LOGIC;
    SIGNAL S7502 : STD_LOGIC;
    SIGNAL S7503 : STD_LOGIC;
    SIGNAL S7504 : STD_LOGIC;
    SIGNAL S7505 : STD_LOGIC;
    SIGNAL S7506 : STD_LOGIC;
    SIGNAL S7507 : STD_LOGIC;
    SIGNAL S7508 : STD_LOGIC;
    SIGNAL S7509 : STD_LOGIC;
    SIGNAL S7510 : STD_LOGIC;
    SIGNAL S7511 : STD_LOGIC;
    SIGNAL S7512 : STD_LOGIC;
    SIGNAL S7513 : STD_LOGIC;
    SIGNAL S7514 : STD_LOGIC;
    SIGNAL S7515 : STD_LOGIC;
    SIGNAL S7516 : STD_LOGIC;
    SIGNAL S7517 : STD_LOGIC;
    SIGNAL S7518 : STD_LOGIC;
    SIGNAL S7519 : STD_LOGIC;
    SIGNAL S7520 : STD_LOGIC;
    SIGNAL S7521 : STD_LOGIC;
    SIGNAL S7522 : STD_LOGIC;
    SIGNAL S7523 : STD_LOGIC;
    SIGNAL S7524 : STD_LOGIC;
    SIGNAL S7525 : STD_LOGIC;
    SIGNAL S7526 : STD_LOGIC;
    SIGNAL S7527 : STD_LOGIC;
    SIGNAL S7528 : STD_LOGIC;
    SIGNAL S7529 : STD_LOGIC;
    SIGNAL S7530 : STD_LOGIC;
    SIGNAL S7531 : STD_LOGIC;
    SIGNAL S7532 : STD_LOGIC;
    SIGNAL S7533 : STD_LOGIC;
    SIGNAL S7534 : STD_LOGIC;
    SIGNAL S7535 : STD_LOGIC;
    SIGNAL S7536 : STD_LOGIC;
    SIGNAL S7537 : STD_LOGIC;
    SIGNAL S7538 : STD_LOGIC;
    SIGNAL S7539 : STD_LOGIC;
    SIGNAL S7540 : STD_LOGIC;
    SIGNAL S7541 : STD_LOGIC;
    SIGNAL S7542 : STD_LOGIC;
    SIGNAL S7543 : STD_LOGIC;
    SIGNAL S7544 : STD_LOGIC;
    SIGNAL S7545 : STD_LOGIC;
    SIGNAL S7546 : STD_LOGIC;
    SIGNAL S7547 : STD_LOGIC;
    SIGNAL S7548 : STD_LOGIC;
    SIGNAL S7549 : STD_LOGIC;
    SIGNAL S7550 : STD_LOGIC;
    SIGNAL S7551 : STD_LOGIC;
    SIGNAL S7552 : STD_LOGIC;
    SIGNAL S7553 : STD_LOGIC;
    SIGNAL S7554 : STD_LOGIC;
    SIGNAL S7555 : STD_LOGIC;
    SIGNAL S7556 : STD_LOGIC;
    SIGNAL S7557 : STD_LOGIC;
    SIGNAL S7558 : STD_LOGIC;
    SIGNAL S7559 : STD_LOGIC;
    SIGNAL S7560 : STD_LOGIC;
    SIGNAL S7561 : STD_LOGIC;
    SIGNAL S7562 : STD_LOGIC;
    SIGNAL S7563 : STD_LOGIC;
    SIGNAL S7564 : STD_LOGIC;
    SIGNAL S7565 : STD_LOGIC;
    SIGNAL S7566 : STD_LOGIC;
    SIGNAL S7567 : STD_LOGIC;
    SIGNAL S7568 : STD_LOGIC;
    SIGNAL S7569 : STD_LOGIC;
    SIGNAL S7570 : STD_LOGIC;
    SIGNAL S7571 : STD_LOGIC;
    SIGNAL S7572 : STD_LOGIC;
    SIGNAL S7573 : STD_LOGIC;
    SIGNAL S7574 : STD_LOGIC;
    SIGNAL S7575 : STD_LOGIC;
    SIGNAL S7576 : STD_LOGIC;
    SIGNAL S7577 : STD_LOGIC;
    SIGNAL S7578 : STD_LOGIC;
    SIGNAL S7579 : STD_LOGIC;
    SIGNAL S7580 : STD_LOGIC;
    SIGNAL S7581 : STD_LOGIC;
    SIGNAL S7582 : STD_LOGIC;
    SIGNAL S7583 : STD_LOGIC;
    SIGNAL S7584 : STD_LOGIC;
    SIGNAL S7585 : STD_LOGIC;
    SIGNAL S7586 : STD_LOGIC;
    SIGNAL S7587 : STD_LOGIC;
    SIGNAL S7588 : STD_LOGIC;
    SIGNAL S7589 : STD_LOGIC;
    SIGNAL S7590 : STD_LOGIC;
    SIGNAL S7591 : STD_LOGIC;
    SIGNAL S7592 : STD_LOGIC;
    SIGNAL S7593 : STD_LOGIC;
    SIGNAL S7594 : STD_LOGIC;
    SIGNAL S7595 : STD_LOGIC;
    SIGNAL S7596 : STD_LOGIC;
    SIGNAL S7597 : STD_LOGIC;
    SIGNAL S7598 : STD_LOGIC;
    SIGNAL S7599 : STD_LOGIC;
    SIGNAL S7600 : STD_LOGIC;
    SIGNAL S7601 : STD_LOGIC;
    SIGNAL S7602 : STD_LOGIC;
    SIGNAL S7603 : STD_LOGIC;
    SIGNAL S7604 : STD_LOGIC;
    SIGNAL S7605 : STD_LOGIC;
    SIGNAL S7606 : STD_LOGIC;
    SIGNAL S7607 : STD_LOGIC;
    SIGNAL S7608 : STD_LOGIC;
    SIGNAL S7609 : STD_LOGIC;
    SIGNAL S7610 : STD_LOGIC;
    SIGNAL S7611 : STD_LOGIC;
    SIGNAL S7612 : STD_LOGIC;
    SIGNAL S7613 : STD_LOGIC;
    SIGNAL S7614 : STD_LOGIC;
    SIGNAL S7615 : STD_LOGIC;
    SIGNAL S7616 : STD_LOGIC;
    SIGNAL S7617 : STD_LOGIC;
    SIGNAL S7618 : STD_LOGIC;
    SIGNAL S7619 : STD_LOGIC;
    SIGNAL S7620 : STD_LOGIC;
    SIGNAL S7621 : STD_LOGIC;
    SIGNAL S7622 : STD_LOGIC;
    SIGNAL S7623 : STD_LOGIC;
    SIGNAL S7624 : STD_LOGIC;
    SIGNAL S7625 : STD_LOGIC;
    SIGNAL S7626 : STD_LOGIC;
    SIGNAL S7627 : STD_LOGIC;
    SIGNAL S7628 : STD_LOGIC;
    SIGNAL S7629 : STD_LOGIC;
    SIGNAL S7630 : STD_LOGIC;
    SIGNAL S7631 : STD_LOGIC;
    SIGNAL S7632 : STD_LOGIC;
    SIGNAL S7633 : STD_LOGIC;
    SIGNAL S7634 : STD_LOGIC;
    SIGNAL S7635 : STD_LOGIC;
    SIGNAL S7636 : STD_LOGIC;
    SIGNAL S7637 : STD_LOGIC;
    SIGNAL S7638 : STD_LOGIC;
    SIGNAL S7639 : STD_LOGIC;
    SIGNAL S7640 : STD_LOGIC;
    SIGNAL S7641 : STD_LOGIC;
    SIGNAL S7642 : STD_LOGIC;
    SIGNAL S7643 : STD_LOGIC;
    SIGNAL S7644 : STD_LOGIC;
    SIGNAL S7645 : STD_LOGIC;
    SIGNAL S7646 : STD_LOGIC;
    SIGNAL S7647 : STD_LOGIC;
    SIGNAL S7648 : STD_LOGIC;
    SIGNAL S7649 : STD_LOGIC;
    SIGNAL S7650 : STD_LOGIC;
    SIGNAL S7651 : STD_LOGIC;
    SIGNAL S7652 : STD_LOGIC;
    SIGNAL S7653 : STD_LOGIC;
    SIGNAL S7654 : STD_LOGIC;
    SIGNAL S7655 : STD_LOGIC;
    SIGNAL S7656 : STD_LOGIC;
    SIGNAL S7657 : STD_LOGIC;
    SIGNAL S7658 : STD_LOGIC;
    SIGNAL S7659 : STD_LOGIC;
    SIGNAL S7660 : STD_LOGIC;
    SIGNAL S7661 : STD_LOGIC;
    SIGNAL S7662 : STD_LOGIC;
    SIGNAL S7663 : STD_LOGIC;
    SIGNAL S7664 : STD_LOGIC;
    SIGNAL S7665 : STD_LOGIC;
    SIGNAL S7666 : STD_LOGIC;
    SIGNAL S7667 : STD_LOGIC;
    SIGNAL S7668 : STD_LOGIC;
    SIGNAL S7669 : STD_LOGIC;
    SIGNAL S7670 : STD_LOGIC;
    SIGNAL S7671 : STD_LOGIC;
    SIGNAL S7672 : STD_LOGIC;
    SIGNAL S7673 : STD_LOGIC;
    SIGNAL S7674 : STD_LOGIC;
    SIGNAL S7675 : STD_LOGIC;
    SIGNAL S7676 : STD_LOGIC;
    SIGNAL S7677 : STD_LOGIC;
    SIGNAL S7678 : STD_LOGIC;
    SIGNAL S7679 : STD_LOGIC;
    SIGNAL S7680 : STD_LOGIC;
    SIGNAL S7681 : STD_LOGIC;
    SIGNAL S7682 : STD_LOGIC;
    SIGNAL S7683 : STD_LOGIC;
    SIGNAL S7684 : STD_LOGIC;
    SIGNAL S7685 : STD_LOGIC;
    SIGNAL S7686 : STD_LOGIC;
    SIGNAL S7687 : STD_LOGIC;
    SIGNAL S7688 : STD_LOGIC;
    SIGNAL S7689 : STD_LOGIC;
    SIGNAL S7690 : STD_LOGIC;
    SIGNAL S7691 : STD_LOGIC;
    SIGNAL S7692 : STD_LOGIC;
    SIGNAL S7693 : STD_LOGIC;
    SIGNAL S7694 : STD_LOGIC;
    SIGNAL S7695 : STD_LOGIC;
    SIGNAL S7696 : STD_LOGIC;
    SIGNAL S7697 : STD_LOGIC;
    SIGNAL S7698 : STD_LOGIC;
    SIGNAL S7699 : STD_LOGIC;
    SIGNAL S7700 : STD_LOGIC;
    SIGNAL S7701 : STD_LOGIC;
    SIGNAL S7702 : STD_LOGIC;
    SIGNAL S7703 : STD_LOGIC;
    SIGNAL S7704 : STD_LOGIC;
    SIGNAL S7705 : STD_LOGIC;
    SIGNAL S7706 : STD_LOGIC;
    SIGNAL S7707 : STD_LOGIC;
    SIGNAL S7708 : STD_LOGIC;
    SIGNAL S7709 : STD_LOGIC;
    SIGNAL S7710 : STD_LOGIC;
    SIGNAL S7711 : STD_LOGIC;
    SIGNAL S7712 : STD_LOGIC;
    SIGNAL S7713 : STD_LOGIC;
    SIGNAL S7714 : STD_LOGIC;
    SIGNAL S7715 : STD_LOGIC;
    SIGNAL S7716 : STD_LOGIC;
    SIGNAL S7717 : STD_LOGIC;
    SIGNAL S7718 : STD_LOGIC;
    SIGNAL S7719 : STD_LOGIC;
    SIGNAL S7720 : STD_LOGIC;
    SIGNAL S7721 : STD_LOGIC;
    SIGNAL S7722 : STD_LOGIC;
    SIGNAL S7723 : STD_LOGIC;
    SIGNAL S7724 : STD_LOGIC;
    SIGNAL S7725 : STD_LOGIC;
    SIGNAL S7726 : STD_LOGIC;
    SIGNAL S7727 : STD_LOGIC;
    SIGNAL S7728 : STD_LOGIC;
    SIGNAL S7729 : STD_LOGIC;
    SIGNAL S7730 : STD_LOGIC;
    SIGNAL S7731 : STD_LOGIC;
    SIGNAL S7732 : STD_LOGIC;
    SIGNAL S7733 : STD_LOGIC;
    SIGNAL S7734 : STD_LOGIC;
    SIGNAL S7735 : STD_LOGIC;
    SIGNAL S7736 : STD_LOGIC;
    SIGNAL S7737 : STD_LOGIC;
    SIGNAL S7738 : STD_LOGIC;
    SIGNAL S7739 : STD_LOGIC;
    SIGNAL S7740 : STD_LOGIC;
    SIGNAL S7741 : STD_LOGIC;
    SIGNAL S7742 : STD_LOGIC;
    SIGNAL S7743 : STD_LOGIC;
    SIGNAL S7744 : STD_LOGIC;
    SIGNAL S7745 : STD_LOGIC;
    SIGNAL S7746 : STD_LOGIC;
    SIGNAL S7747 : STD_LOGIC;
    SIGNAL S7748 : STD_LOGIC;
    SIGNAL S7749 : STD_LOGIC;
    SIGNAL S7750 : STD_LOGIC;
    SIGNAL S7751 : STD_LOGIC;
    SIGNAL S7752 : STD_LOGIC;
    SIGNAL S7753 : STD_LOGIC;
    SIGNAL S7754 : STD_LOGIC;
    SIGNAL S7755 : STD_LOGIC;
    SIGNAL S7756 : STD_LOGIC;
    SIGNAL S7757 : STD_LOGIC;
    SIGNAL S7758 : STD_LOGIC;
    SIGNAL S7759 : STD_LOGIC;
    SIGNAL S7760 : STD_LOGIC;
    SIGNAL S7761 : STD_LOGIC;
    SIGNAL S7762 : STD_LOGIC;
    SIGNAL S7763 : STD_LOGIC;
    SIGNAL S7764 : STD_LOGIC;
    SIGNAL S7765 : STD_LOGIC;
    SIGNAL S7766 : STD_LOGIC;
    SIGNAL S7767 : STD_LOGIC;
    SIGNAL S7768 : STD_LOGIC;
    SIGNAL S7769 : STD_LOGIC;
    SIGNAL S7770 : STD_LOGIC;
    SIGNAL S7771 : STD_LOGIC;
    SIGNAL S7772 : STD_LOGIC;
    SIGNAL S7773 : STD_LOGIC;
    SIGNAL S7774 : STD_LOGIC;
    SIGNAL S7775 : STD_LOGIC;
    SIGNAL S7776 : STD_LOGIC;
    SIGNAL S7777 : STD_LOGIC;
    SIGNAL S7778 : STD_LOGIC;
    SIGNAL S7779 : STD_LOGIC;
    SIGNAL S7780 : STD_LOGIC;
    SIGNAL S7781 : STD_LOGIC;
    SIGNAL S7782 : STD_LOGIC;
    SIGNAL S7783 : STD_LOGIC;
    SIGNAL S7784 : STD_LOGIC;
    SIGNAL S7785 : STD_LOGIC;
    SIGNAL S7786 : STD_LOGIC;
    SIGNAL S7787 : STD_LOGIC;
    SIGNAL S7788 : STD_LOGIC;
    SIGNAL S7789 : STD_LOGIC;
    SIGNAL S7790 : STD_LOGIC;
    SIGNAL S7791 : STD_LOGIC;
    SIGNAL S7792 : STD_LOGIC;
    SIGNAL S7793 : STD_LOGIC;
    SIGNAL S7794 : STD_LOGIC;
    SIGNAL S7795 : STD_LOGIC;
    SIGNAL S7796 : STD_LOGIC;
    SIGNAL S7797 : STD_LOGIC;
    SIGNAL S7798 : STD_LOGIC;
    SIGNAL S7799 : STD_LOGIC;
    SIGNAL S7800 : STD_LOGIC;
    SIGNAL S7801 : STD_LOGIC;
    SIGNAL S7802 : STD_LOGIC;
    SIGNAL S7803 : STD_LOGIC;
    SIGNAL S7804 : STD_LOGIC;
    SIGNAL S7805 : STD_LOGIC;
    SIGNAL S7806 : STD_LOGIC;
    SIGNAL S7807 : STD_LOGIC;
    SIGNAL S7808 : STD_LOGIC;
    SIGNAL S7809 : STD_LOGIC;
    SIGNAL S7810 : STD_LOGIC;
    SIGNAL S7811 : STD_LOGIC;
    SIGNAL S7812 : STD_LOGIC;
    SIGNAL S7813 : STD_LOGIC;
    SIGNAL S7814 : STD_LOGIC;
    SIGNAL S7815 : STD_LOGIC;
    SIGNAL S7816 : STD_LOGIC;
    SIGNAL S7817 : STD_LOGIC;
    SIGNAL S7818 : STD_LOGIC;
    SIGNAL S7819 : STD_LOGIC;
    SIGNAL S7820 : STD_LOGIC;
    SIGNAL S7821 : STD_LOGIC;
    SIGNAL S7822 : STD_LOGIC;
    SIGNAL S7823 : STD_LOGIC;
    SIGNAL S7824 : STD_LOGIC;
    SIGNAL S7825 : STD_LOGIC;
    SIGNAL S7826 : STD_LOGIC;
    SIGNAL S7827 : STD_LOGIC;
    SIGNAL S7828 : STD_LOGIC;
    SIGNAL S7829 : STD_LOGIC;
    SIGNAL S7830 : STD_LOGIC;
    SIGNAL S7831 : STD_LOGIC;
    SIGNAL S7832 : STD_LOGIC;
    SIGNAL S7833 : STD_LOGIC;
    SIGNAL S7834 : STD_LOGIC;
    SIGNAL S7835 : STD_LOGIC;
    SIGNAL S7836 : STD_LOGIC;
    SIGNAL S7837 : STD_LOGIC;
    SIGNAL S7838 : STD_LOGIC;
    SIGNAL S7839 : STD_LOGIC;
    SIGNAL S7840 : STD_LOGIC;
    SIGNAL S7841 : STD_LOGIC;
    SIGNAL S7842 : STD_LOGIC;
    SIGNAL S7843 : STD_LOGIC;
    SIGNAL S7844 : STD_LOGIC;
    SIGNAL S7845 : STD_LOGIC;
    SIGNAL S7846 : STD_LOGIC;
    SIGNAL S7847 : STD_LOGIC;
    SIGNAL S7848 : STD_LOGIC;
    SIGNAL S7849 : STD_LOGIC;
    SIGNAL S7850 : STD_LOGIC;
    SIGNAL S7851 : STD_LOGIC;
    SIGNAL S7852 : STD_LOGIC;
    SIGNAL S7853 : STD_LOGIC;
    SIGNAL S7854 : STD_LOGIC;
    SIGNAL S7855 : STD_LOGIC;
    SIGNAL S7856 : STD_LOGIC;
    SIGNAL S7857 : STD_LOGIC;
    SIGNAL S7858 : STD_LOGIC;
    SIGNAL S7859 : STD_LOGIC;
    SIGNAL S7860 : STD_LOGIC;
    SIGNAL S7861 : STD_LOGIC;
    SIGNAL S7862 : STD_LOGIC;
    SIGNAL S7863 : STD_LOGIC;
    SIGNAL S7864 : STD_LOGIC;
    SIGNAL S7865 : STD_LOGIC;
    SIGNAL S7866 : STD_LOGIC;
    SIGNAL S7867 : STD_LOGIC;
    SIGNAL S7868 : STD_LOGIC;
    SIGNAL S7869 : STD_LOGIC;
    SIGNAL S7870 : STD_LOGIC;
    SIGNAL S7871 : STD_LOGIC;
    SIGNAL S7872 : STD_LOGIC;
    SIGNAL S7873 : STD_LOGIC;
    SIGNAL S7874 : STD_LOGIC;
    SIGNAL S7875 : STD_LOGIC;
    SIGNAL S7876 : STD_LOGIC;
    SIGNAL S7877 : STD_LOGIC;
    SIGNAL S7878 : STD_LOGIC;
    SIGNAL S7879 : STD_LOGIC;
    SIGNAL S7880 : STD_LOGIC;
    SIGNAL S7881 : STD_LOGIC;
    SIGNAL S7882 : STD_LOGIC;
    SIGNAL S7883 : STD_LOGIC;
    SIGNAL S7884 : STD_LOGIC;
    SIGNAL S7885 : STD_LOGIC;
    SIGNAL S7886 : STD_LOGIC;
    SIGNAL S7887 : STD_LOGIC;
    SIGNAL S7888 : STD_LOGIC;
    SIGNAL S7889 : STD_LOGIC;
    SIGNAL S7890 : STD_LOGIC;
    SIGNAL S7891 : STD_LOGIC;
    SIGNAL S7892 : STD_LOGIC;
    SIGNAL S7893 : STD_LOGIC;
    SIGNAL S7894 : STD_LOGIC;
    SIGNAL S7895 : STD_LOGIC;
    SIGNAL S7896 : STD_LOGIC;
    SIGNAL S7897 : STD_LOGIC;
    SIGNAL S7898 : STD_LOGIC;
    SIGNAL S7899 : STD_LOGIC;
    SIGNAL S7900 : STD_LOGIC;
    SIGNAL S7901 : STD_LOGIC;
    SIGNAL S7902 : STD_LOGIC;
    SIGNAL S7903 : STD_LOGIC;
    SIGNAL S7904 : STD_LOGIC;
    SIGNAL S7905 : STD_LOGIC;
    SIGNAL S7906 : STD_LOGIC;
    SIGNAL S7907 : STD_LOGIC;
    SIGNAL S7908 : STD_LOGIC;
    SIGNAL S7909 : STD_LOGIC;
    SIGNAL S7910 : STD_LOGIC;
    SIGNAL S7911 : STD_LOGIC;
    SIGNAL S7912 : STD_LOGIC;
    SIGNAL S7913 : STD_LOGIC;
    SIGNAL S7914 : STD_LOGIC;
    SIGNAL S7915 : STD_LOGIC;
    SIGNAL S7916 : STD_LOGIC;
    SIGNAL S7917 : STD_LOGIC;
    SIGNAL S7918 : STD_LOGIC;
    SIGNAL S7919 : STD_LOGIC;
    SIGNAL S7920 : STD_LOGIC;
    SIGNAL S7921 : STD_LOGIC;
    SIGNAL S7922 : STD_LOGIC;
    SIGNAL S7923 : STD_LOGIC;
    SIGNAL S7924 : STD_LOGIC;
    SIGNAL S7925 : STD_LOGIC;
    SIGNAL S7926 : STD_LOGIC;
    SIGNAL S7927 : STD_LOGIC;
    SIGNAL S7928 : STD_LOGIC;
    SIGNAL S7929 : STD_LOGIC;
    SIGNAL S7930 : STD_LOGIC;
    SIGNAL S7931 : STD_LOGIC;
    SIGNAL S7932 : STD_LOGIC;
    SIGNAL S7933 : STD_LOGIC;
    SIGNAL S7934 : STD_LOGIC;
    SIGNAL S7935 : STD_LOGIC;
    SIGNAL S7936 : STD_LOGIC;
    SIGNAL S7937 : STD_LOGIC;
    SIGNAL S7938 : STD_LOGIC;
    SIGNAL S7939 : STD_LOGIC;
    SIGNAL S7940 : STD_LOGIC;
    SIGNAL S7941 : STD_LOGIC;
    SIGNAL S7942 : STD_LOGIC;
    SIGNAL S7943 : STD_LOGIC;
    SIGNAL S7944 : STD_LOGIC;
    SIGNAL S7945 : STD_LOGIC;
    SIGNAL S7946 : STD_LOGIC;
    SIGNAL S7947 : STD_LOGIC;
    SIGNAL S7948 : STD_LOGIC;
    SIGNAL S7949 : STD_LOGIC;
    SIGNAL S7950 : STD_LOGIC;
    SIGNAL S7951 : STD_LOGIC;
    SIGNAL S7952 : STD_LOGIC;
    SIGNAL S7953 : STD_LOGIC;
    SIGNAL S7954 : STD_LOGIC;
    SIGNAL S7955 : STD_LOGIC;
    SIGNAL S7956 : STD_LOGIC;
    SIGNAL S7957 : STD_LOGIC;
    SIGNAL S7958 : STD_LOGIC;
    SIGNAL S7959 : STD_LOGIC;
    SIGNAL S7960 : STD_LOGIC;
    SIGNAL S7961 : STD_LOGIC;
    SIGNAL S7962 : STD_LOGIC;
    SIGNAL S7963 : STD_LOGIC;
    SIGNAL S7964 : STD_LOGIC;
    SIGNAL S7965 : STD_LOGIC;
    SIGNAL S7966 : STD_LOGIC;
    SIGNAL S7967 : STD_LOGIC;
    SIGNAL S7968 : STD_LOGIC;
    SIGNAL S7969 : STD_LOGIC;
    SIGNAL S7970 : STD_LOGIC;
    SIGNAL S7971 : STD_LOGIC;
    SIGNAL S7972 : STD_LOGIC;
    SIGNAL S7973 : STD_LOGIC;
    SIGNAL S7974 : STD_LOGIC;
    SIGNAL S7975 : STD_LOGIC;
    SIGNAL S7976 : STD_LOGIC;
    SIGNAL S7977 : STD_LOGIC;
    SIGNAL S7978 : STD_LOGIC;
    SIGNAL S7979 : STD_LOGIC;
    SIGNAL S7980 : STD_LOGIC;
    SIGNAL S7981 : STD_LOGIC;
    SIGNAL S7982 : STD_LOGIC;
    SIGNAL S7983 : STD_LOGIC;
    SIGNAL S7984 : STD_LOGIC;
    SIGNAL S7985 : STD_LOGIC;
    SIGNAL S7986 : STD_LOGIC;
    SIGNAL S7987 : STD_LOGIC;
    SIGNAL S7988 : STD_LOGIC;
    SIGNAL S7989 : STD_LOGIC;
    SIGNAL S7990 : STD_LOGIC;
    SIGNAL S7991 : STD_LOGIC;
    SIGNAL S7992 : STD_LOGIC;
    SIGNAL S7993 : STD_LOGIC;
    SIGNAL S7994 : STD_LOGIC;
    SIGNAL S7995 : STD_LOGIC;
    SIGNAL S7996 : STD_LOGIC;
    SIGNAL S7997 : STD_LOGIC;
    SIGNAL S7998 : STD_LOGIC;
    SIGNAL S7999 : STD_LOGIC;
    SIGNAL S8000 : STD_LOGIC;
    SIGNAL S8001 : STD_LOGIC;
    SIGNAL S8002 : STD_LOGIC;
    SIGNAL S8003 : STD_LOGIC;
    SIGNAL S8004 : STD_LOGIC;
    SIGNAL S8005 : STD_LOGIC;
    SIGNAL S8006 : STD_LOGIC;
    SIGNAL S8007 : STD_LOGIC;
    SIGNAL S8008 : STD_LOGIC;
    SIGNAL S8009 : STD_LOGIC;
    SIGNAL S8010 : STD_LOGIC;
    SIGNAL S8011 : STD_LOGIC;
    SIGNAL S8012 : STD_LOGIC;
    SIGNAL S8013 : STD_LOGIC;
    SIGNAL S8014 : STD_LOGIC;
    SIGNAL S8015 : STD_LOGIC;
    SIGNAL S8016 : STD_LOGIC;
    SIGNAL S8017 : STD_LOGIC;
    SIGNAL S8018 : STD_LOGIC;
    SIGNAL S8019 : STD_LOGIC;
    SIGNAL S8020 : STD_LOGIC;
    SIGNAL S8021 : STD_LOGIC;
    SIGNAL S8022 : STD_LOGIC;
    SIGNAL S8023 : STD_LOGIC;
    SIGNAL S8024 : STD_LOGIC;
    SIGNAL S8025 : STD_LOGIC;
    SIGNAL S8026 : STD_LOGIC;
    SIGNAL S8027 : STD_LOGIC;
    SIGNAL S8028 : STD_LOGIC;
    SIGNAL S8029 : STD_LOGIC;
    SIGNAL S8030 : STD_LOGIC;
    SIGNAL S8031 : STD_LOGIC;
    SIGNAL S8032 : STD_LOGIC;
    SIGNAL S8033 : STD_LOGIC;
    SIGNAL S8034 : STD_LOGIC;
    SIGNAL S8035 : STD_LOGIC;
    SIGNAL S8036 : STD_LOGIC;
    SIGNAL S8037 : STD_LOGIC;
    SIGNAL S8038 : STD_LOGIC;
    SIGNAL S8039 : STD_LOGIC;
    SIGNAL S8040 : STD_LOGIC;
    SIGNAL S8041 : STD_LOGIC;
    SIGNAL S8042 : STD_LOGIC;
    SIGNAL S8043 : STD_LOGIC;
    SIGNAL S8044 : STD_LOGIC;
    SIGNAL S8045 : STD_LOGIC;
    SIGNAL S8046 : STD_LOGIC;
    SIGNAL S8047 : STD_LOGIC;
    SIGNAL S8048 : STD_LOGIC;
    SIGNAL S8049 : STD_LOGIC;
    SIGNAL S8050 : STD_LOGIC;
    SIGNAL S8051 : STD_LOGIC;
    SIGNAL S8052 : STD_LOGIC;
    SIGNAL S8053 : STD_LOGIC;
    SIGNAL S8054 : STD_LOGIC;
    SIGNAL S8055 : STD_LOGIC;
    SIGNAL S8056 : STD_LOGIC;
    SIGNAL S8057 : STD_LOGIC;
    SIGNAL S8058 : STD_LOGIC;
    SIGNAL S8059 : STD_LOGIC;
    SIGNAL S8060 : STD_LOGIC;
    SIGNAL S8061 : STD_LOGIC;
    SIGNAL S8062 : STD_LOGIC;
    SIGNAL S8063 : STD_LOGIC;
    SIGNAL S8064 : STD_LOGIC;
    SIGNAL S8065 : STD_LOGIC;
    SIGNAL S8066 : STD_LOGIC;
    SIGNAL S8067 : STD_LOGIC;
    SIGNAL S8068 : STD_LOGIC;
    SIGNAL S8069 : STD_LOGIC;
    SIGNAL S8070 : STD_LOGIC;
    SIGNAL S8071 : STD_LOGIC;
    SIGNAL S8072 : STD_LOGIC;
    SIGNAL S8073 : STD_LOGIC;
    SIGNAL S8074 : STD_LOGIC;
    SIGNAL S8075 : STD_LOGIC;
    SIGNAL S8076 : STD_LOGIC;
    SIGNAL S8077 : STD_LOGIC;
    SIGNAL S8078 : STD_LOGIC;
    SIGNAL S8079 : STD_LOGIC;
    SIGNAL S8080 : STD_LOGIC;
    SIGNAL S8081 : STD_LOGIC;
    SIGNAL S8082 : STD_LOGIC;
    SIGNAL S8083 : STD_LOGIC;
    SIGNAL S8084 : STD_LOGIC;
    SIGNAL S8085 : STD_LOGIC;
    SIGNAL S8086 : STD_LOGIC;
    SIGNAL S8087 : STD_LOGIC;
    SIGNAL S8088 : STD_LOGIC;
    SIGNAL S8089 : STD_LOGIC;
    SIGNAL S8090 : STD_LOGIC;
    SIGNAL S8091 : STD_LOGIC;
    SIGNAL S8092 : STD_LOGIC;
    SIGNAL S8093 : STD_LOGIC;
    SIGNAL S8094 : STD_LOGIC;
    SIGNAL S8095 : STD_LOGIC;
    SIGNAL S8096 : STD_LOGIC;
    SIGNAL S8097 : STD_LOGIC;
    SIGNAL S8098 : STD_LOGIC;
    SIGNAL S8099 : STD_LOGIC;
    SIGNAL S8100 : STD_LOGIC;
    SIGNAL S8101 : STD_LOGIC;
    SIGNAL S8102 : STD_LOGIC;
    SIGNAL S8103 : STD_LOGIC;
    SIGNAL S8104 : STD_LOGIC;
    SIGNAL S8105 : STD_LOGIC;
    SIGNAL S8106 : STD_LOGIC;
    SIGNAL S8107 : STD_LOGIC;
    SIGNAL S8108 : STD_LOGIC;
    SIGNAL S8109 : STD_LOGIC;
    SIGNAL S8110 : STD_LOGIC;
    SIGNAL S8111 : STD_LOGIC;
    SIGNAL S8112 : STD_LOGIC;
    SIGNAL S8113 : STD_LOGIC;
    SIGNAL S8114 : STD_LOGIC;
    SIGNAL S8115 : STD_LOGIC;
    SIGNAL S8116 : STD_LOGIC;
    SIGNAL S8117 : STD_LOGIC;
    SIGNAL S8118 : STD_LOGIC;
    SIGNAL S8119 : STD_LOGIC;
    SIGNAL S8120 : STD_LOGIC;
    SIGNAL S8121 : STD_LOGIC;
    SIGNAL S8122 : STD_LOGIC;
    SIGNAL S8123 : STD_LOGIC;
    SIGNAL S8124 : STD_LOGIC;
    SIGNAL S8125 : STD_LOGIC;
    SIGNAL S8126 : STD_LOGIC;
    SIGNAL S8127 : STD_LOGIC;
    SIGNAL S8128 : STD_LOGIC;
    SIGNAL S8129 : STD_LOGIC;
    SIGNAL S8130 : STD_LOGIC;
    SIGNAL S8131 : STD_LOGIC;
    SIGNAL S8132 : STD_LOGIC;
    SIGNAL S8133 : STD_LOGIC;
    SIGNAL S8134 : STD_LOGIC;
    SIGNAL S8135 : STD_LOGIC;
    SIGNAL S8136 : STD_LOGIC;
    SIGNAL S8137 : STD_LOGIC;
    SIGNAL S8138 : STD_LOGIC;
    SIGNAL S8139 : STD_LOGIC;
    SIGNAL S8140 : STD_LOGIC;
    SIGNAL S8141 : STD_LOGIC;
    SIGNAL S8142 : STD_LOGIC;
    SIGNAL S8143 : STD_LOGIC;
    SIGNAL S8144 : STD_LOGIC;
    SIGNAL S8145 : STD_LOGIC;
    SIGNAL S8146 : STD_LOGIC;
    SIGNAL S8147 : STD_LOGIC;
    SIGNAL S8148 : STD_LOGIC;
    SIGNAL S8149 : STD_LOGIC;
    SIGNAL S8150 : STD_LOGIC;
    SIGNAL S8151 : STD_LOGIC;
    SIGNAL S8152 : STD_LOGIC;
    SIGNAL S8153 : STD_LOGIC;
    SIGNAL S8154 : STD_LOGIC;
    SIGNAL S8155 : STD_LOGIC;
    SIGNAL S8156 : STD_LOGIC;
    SIGNAL S8157 : STD_LOGIC;
    SIGNAL S8158 : STD_LOGIC;
    SIGNAL S8159 : STD_LOGIC;
    SIGNAL S8160 : STD_LOGIC;
    SIGNAL S8161 : STD_LOGIC;
    SIGNAL S8162 : STD_LOGIC;
    SIGNAL S8163 : STD_LOGIC;
    SIGNAL S8164 : STD_LOGIC;
    SIGNAL S8165 : STD_LOGIC;
    SIGNAL S8166 : STD_LOGIC;
    SIGNAL S8167 : STD_LOGIC;
    SIGNAL S8168 : STD_LOGIC;
    SIGNAL S8169 : STD_LOGIC;
    SIGNAL S8170 : STD_LOGIC;
    SIGNAL S8171 : STD_LOGIC;
    SIGNAL S8172 : STD_LOGIC;
    SIGNAL S8173 : STD_LOGIC;
    SIGNAL S8174 : STD_LOGIC;
    SIGNAL S8175 : STD_LOGIC;
    SIGNAL S8176 : STD_LOGIC;
    SIGNAL S8177 : STD_LOGIC;
    SIGNAL S8178 : STD_LOGIC;
    SIGNAL S8179 : STD_LOGIC;
    SIGNAL S8180 : STD_LOGIC;
    SIGNAL S8181 : STD_LOGIC;
    SIGNAL S8182 : STD_LOGIC;
    SIGNAL S8183 : STD_LOGIC;
    SIGNAL S8184 : STD_LOGIC;
    SIGNAL S8185 : STD_LOGIC;
    SIGNAL S8186 : STD_LOGIC;
    SIGNAL S8187 : STD_LOGIC;
    SIGNAL S8188 : STD_LOGIC;
    SIGNAL S8189 : STD_LOGIC;
    SIGNAL S8190 : STD_LOGIC;
    SIGNAL S8191 : STD_LOGIC;
    SIGNAL S8192 : STD_LOGIC;
    SIGNAL S8193 : STD_LOGIC;
    SIGNAL S8194 : STD_LOGIC;
    SIGNAL S8195 : STD_LOGIC;
    SIGNAL S8196 : STD_LOGIC;
    SIGNAL S8197 : STD_LOGIC;
    SIGNAL S8198 : STD_LOGIC;
    SIGNAL S8199 : STD_LOGIC;
    SIGNAL S8200 : STD_LOGIC;
    SIGNAL S8201 : STD_LOGIC;
    SIGNAL S8202 : STD_LOGIC;
    SIGNAL S8203 : STD_LOGIC;
    SIGNAL S8204 : STD_LOGIC;
    SIGNAL S8205 : STD_LOGIC;
    SIGNAL S8206 : STD_LOGIC;
    SIGNAL S8207 : STD_LOGIC;
    SIGNAL S8208 : STD_LOGIC;
    SIGNAL S8209 : STD_LOGIC;
    SIGNAL S8210 : STD_LOGIC;
    SIGNAL S8211 : STD_LOGIC;
    SIGNAL S8212 : STD_LOGIC;
    SIGNAL S8213 : STD_LOGIC;
    SIGNAL S8214 : STD_LOGIC;
    SIGNAL S8215 : STD_LOGIC;
    SIGNAL S8216 : STD_LOGIC;
    SIGNAL S8217 : STD_LOGIC;
    SIGNAL S8218 : STD_LOGIC;
    SIGNAL S8219 : STD_LOGIC;
    SIGNAL S8220 : STD_LOGIC;
    SIGNAL S8221 : STD_LOGIC;
    SIGNAL S8222 : STD_LOGIC;
    SIGNAL S8223 : STD_LOGIC;
    SIGNAL S8224 : STD_LOGIC;
    SIGNAL S8225 : STD_LOGIC;
    SIGNAL S8226 : STD_LOGIC;
    SIGNAL S8227 : STD_LOGIC;
    SIGNAL S8228 : STD_LOGIC;
    SIGNAL S8229 : STD_LOGIC;
    SIGNAL S8230 : STD_LOGIC;
    SIGNAL S8231 : STD_LOGIC;
    SIGNAL S8232 : STD_LOGIC;
    SIGNAL S8233 : STD_LOGIC;
    SIGNAL S8234 : STD_LOGIC;
    SIGNAL S8235 : STD_LOGIC;
    SIGNAL S8236 : STD_LOGIC;
    SIGNAL S8237 : STD_LOGIC;
    SIGNAL S8238 : STD_LOGIC;
    SIGNAL S8239 : STD_LOGIC;
    SIGNAL S8240 : STD_LOGIC;
    SIGNAL S8241 : STD_LOGIC;
    SIGNAL S8242 : STD_LOGIC;
    SIGNAL S8243 : STD_LOGIC;
    SIGNAL S8244 : STD_LOGIC;
    SIGNAL S8245 : STD_LOGIC;
    SIGNAL S8246 : STD_LOGIC;
    SIGNAL S8247 : STD_LOGIC;
    SIGNAL S8248 : STD_LOGIC;
    SIGNAL S8249 : STD_LOGIC;
    SIGNAL S8250 : STD_LOGIC;
    SIGNAL S8251 : STD_LOGIC;
    SIGNAL S8252 : STD_LOGIC;
    SIGNAL S8253 : STD_LOGIC;
    SIGNAL S8254 : STD_LOGIC;
    SIGNAL S8255 : STD_LOGIC;
    SIGNAL S8256 : STD_LOGIC;
    SIGNAL S8257 : STD_LOGIC;
    SIGNAL S8258 : STD_LOGIC;
    SIGNAL S8259 : STD_LOGIC;
    SIGNAL S8260 : STD_LOGIC;
    SIGNAL S8261 : STD_LOGIC;
    SIGNAL S8262 : STD_LOGIC;
    SIGNAL S8263 : STD_LOGIC;
    SIGNAL S8264 : STD_LOGIC;
    SIGNAL S8265 : STD_LOGIC;
    SIGNAL S8266 : STD_LOGIC;
    SIGNAL S8267 : STD_LOGIC;
    SIGNAL S8268 : STD_LOGIC;
    SIGNAL S8269 : STD_LOGIC;
    SIGNAL S8270 : STD_LOGIC;
    SIGNAL S8271 : STD_LOGIC;
    SIGNAL S8272 : STD_LOGIC;
    SIGNAL S8273 : STD_LOGIC;
    SIGNAL S8274 : STD_LOGIC;
    SIGNAL S8275 : STD_LOGIC;
    SIGNAL S8276 : STD_LOGIC;
    SIGNAL S8277 : STD_LOGIC;
    SIGNAL S8278 : STD_LOGIC;
    SIGNAL S8279 : STD_LOGIC;
    SIGNAL S8280 : STD_LOGIC;
    SIGNAL S8281 : STD_LOGIC;
    SIGNAL S8282 : STD_LOGIC;
    SIGNAL S8283 : STD_LOGIC;
    SIGNAL S8284 : STD_LOGIC;
    SIGNAL S8285 : STD_LOGIC;
    SIGNAL S8286 : STD_LOGIC;
    SIGNAL S8287 : STD_LOGIC;
    SIGNAL S8288 : STD_LOGIC;
    SIGNAL S8289 : STD_LOGIC;
    SIGNAL S8290 : STD_LOGIC;
    SIGNAL S8291 : STD_LOGIC;
    SIGNAL S8292 : STD_LOGIC;
    SIGNAL S8293 : STD_LOGIC;
    SIGNAL S8294 : STD_LOGIC;
    SIGNAL S8295 : STD_LOGIC;
    SIGNAL S8296 : STD_LOGIC;
    SIGNAL S8297 : STD_LOGIC;
    SIGNAL S8298 : STD_LOGIC;
    SIGNAL S8299 : STD_LOGIC;
    SIGNAL S8300 : STD_LOGIC;
    SIGNAL S8301 : STD_LOGIC;
    SIGNAL S8302 : STD_LOGIC;
    SIGNAL S8303 : STD_LOGIC;
    SIGNAL S8304 : STD_LOGIC;
    SIGNAL S8305 : STD_LOGIC;
    SIGNAL S8306 : STD_LOGIC;
    SIGNAL S8307 : STD_LOGIC;
    SIGNAL S8308 : STD_LOGIC;
    SIGNAL S8309 : STD_LOGIC;
    SIGNAL S8310 : STD_LOGIC;
    SIGNAL S8311 : STD_LOGIC;
    SIGNAL S8312 : STD_LOGIC;
    SIGNAL S8313 : STD_LOGIC;
    SIGNAL S8314 : STD_LOGIC;
    SIGNAL S8315 : STD_LOGIC;
    SIGNAL S8316 : STD_LOGIC;
    SIGNAL S8317 : STD_LOGIC;
    SIGNAL S8318 : STD_LOGIC;
    SIGNAL S8319 : STD_LOGIC;
    SIGNAL S8320 : STD_LOGIC;
    SIGNAL S8321 : STD_LOGIC;
    SIGNAL S8322 : STD_LOGIC;
    SIGNAL S8323 : STD_LOGIC;
    SIGNAL S8324 : STD_LOGIC;
    SIGNAL S8325 : STD_LOGIC;
    SIGNAL S8326 : STD_LOGIC;
    SIGNAL S8327 : STD_LOGIC;
    SIGNAL S8328 : STD_LOGIC;
    SIGNAL S8329 : STD_LOGIC;
    SIGNAL S8330 : STD_LOGIC;
    SIGNAL S8331 : STD_LOGIC;
    SIGNAL S8332 : STD_LOGIC;
    SIGNAL S8333 : STD_LOGIC;
    SIGNAL S8334 : STD_LOGIC;
    SIGNAL S8335 : STD_LOGIC;
    SIGNAL S8336 : STD_LOGIC;
    SIGNAL S8337 : STD_LOGIC;
    SIGNAL S8338 : STD_LOGIC;
    SIGNAL S8339 : STD_LOGIC;
    SIGNAL S8340 : STD_LOGIC;
    SIGNAL S8341 : STD_LOGIC;
    SIGNAL S8342 : STD_LOGIC;
    SIGNAL S8343 : STD_LOGIC;
    SIGNAL S8344 : STD_LOGIC;
    SIGNAL S8345 : STD_LOGIC;
    SIGNAL S8346 : STD_LOGIC;
    SIGNAL S8347 : STD_LOGIC;
    SIGNAL S8348 : STD_LOGIC;
    SIGNAL S8349 : STD_LOGIC;
    SIGNAL S8350 : STD_LOGIC;
    SIGNAL S8351 : STD_LOGIC;
    SIGNAL S8352 : STD_LOGIC;
    SIGNAL S8353 : STD_LOGIC;
    SIGNAL S8354 : STD_LOGIC;
    SIGNAL S8355 : STD_LOGIC;
    SIGNAL S8356 : STD_LOGIC;
    SIGNAL S8357 : STD_LOGIC;
    SIGNAL S8358 : STD_LOGIC;
    SIGNAL S8359 : STD_LOGIC;
    SIGNAL S8360 : STD_LOGIC;
    SIGNAL S8361 : STD_LOGIC;
    SIGNAL S8362 : STD_LOGIC;
    SIGNAL S8363 : STD_LOGIC;
    SIGNAL S8364 : STD_LOGIC;
    SIGNAL S8365 : STD_LOGIC;
    SIGNAL S8366 : STD_LOGIC;
    SIGNAL S8367 : STD_LOGIC;
    SIGNAL S8368 : STD_LOGIC;
    SIGNAL S8369 : STD_LOGIC;
    SIGNAL S8370 : STD_LOGIC;
    SIGNAL S8371 : STD_LOGIC;
    SIGNAL S8372 : STD_LOGIC;
    SIGNAL S8373 : STD_LOGIC;
    SIGNAL S8374 : STD_LOGIC;
    SIGNAL S8375 : STD_LOGIC;
    SIGNAL S8376 : STD_LOGIC;
    SIGNAL S8377 : STD_LOGIC;
    SIGNAL S8378 : STD_LOGIC;
    SIGNAL S8379 : STD_LOGIC;
    SIGNAL S8380 : STD_LOGIC;
    SIGNAL S8381 : STD_LOGIC;
    SIGNAL S8382 : STD_LOGIC;
    SIGNAL S8383 : STD_LOGIC;
    SIGNAL S8384 : STD_LOGIC;
    SIGNAL S8385 : STD_LOGIC;
    SIGNAL S8386 : STD_LOGIC;
    SIGNAL S8387 : STD_LOGIC;
    SIGNAL S8388 : STD_LOGIC;
    SIGNAL S8389 : STD_LOGIC;
    SIGNAL S8390 : STD_LOGIC;
    SIGNAL S8391 : STD_LOGIC;
    SIGNAL S8392 : STD_LOGIC;
    SIGNAL S8393 : STD_LOGIC;
    SIGNAL S8394 : STD_LOGIC;
    SIGNAL S8395 : STD_LOGIC;
    SIGNAL S8396 : STD_LOGIC;
    SIGNAL S8397 : STD_LOGIC;
    SIGNAL S8398 : STD_LOGIC;
    SIGNAL S8399 : STD_LOGIC;
    SIGNAL S8400 : STD_LOGIC;
    SIGNAL S8401 : STD_LOGIC;
    SIGNAL S8402 : STD_LOGIC;
    SIGNAL S8403 : STD_LOGIC;
    SIGNAL S8404 : STD_LOGIC;
    SIGNAL S8405 : STD_LOGIC;
    SIGNAL S8406 : STD_LOGIC;
    SIGNAL S8407 : STD_LOGIC;
    SIGNAL S8408 : STD_LOGIC;
    SIGNAL S8409 : STD_LOGIC;
    SIGNAL S8410 : STD_LOGIC;
    SIGNAL S8411 : STD_LOGIC;
    SIGNAL S8412 : STD_LOGIC;
    SIGNAL S8413 : STD_LOGIC;
    SIGNAL S8414 : STD_LOGIC;
    SIGNAL S8415 : STD_LOGIC;
    SIGNAL S8416 : STD_LOGIC;
    SIGNAL S8417 : STD_LOGIC;
    SIGNAL S8418 : STD_LOGIC;
    SIGNAL S8419 : STD_LOGIC;
    SIGNAL S8420 : STD_LOGIC;
    SIGNAL S8421 : STD_LOGIC;
    SIGNAL S8422 : STD_LOGIC;
    SIGNAL S8423 : STD_LOGIC;
    SIGNAL S8424 : STD_LOGIC;
    SIGNAL S8425 : STD_LOGIC;
    SIGNAL S8426 : STD_LOGIC;
    SIGNAL S8427 : STD_LOGIC;
    SIGNAL S8428 : STD_LOGIC;
    SIGNAL S8429 : STD_LOGIC;
    SIGNAL S8430 : STD_LOGIC;
    SIGNAL S8431 : STD_LOGIC;
    SIGNAL S8432 : STD_LOGIC;
    SIGNAL S8433 : STD_LOGIC;
    SIGNAL S8434 : STD_LOGIC;
    SIGNAL S8435 : STD_LOGIC;
    SIGNAL S8436 : STD_LOGIC;
    SIGNAL S8437 : STD_LOGIC;
    SIGNAL S8438 : STD_LOGIC;
    SIGNAL S8439 : STD_LOGIC;
    SIGNAL S8440 : STD_LOGIC;
    SIGNAL S8441 : STD_LOGIC;
    SIGNAL S8442 : STD_LOGIC;
    SIGNAL S8443 : STD_LOGIC;
    SIGNAL S8444 : STD_LOGIC;
    SIGNAL S8445 : STD_LOGIC;
    SIGNAL S8446 : STD_LOGIC;
    SIGNAL S8447 : STD_LOGIC;
    SIGNAL S8448 : STD_LOGIC;
    SIGNAL S8449 : STD_LOGIC;
    SIGNAL S8450 : STD_LOGIC;
    SIGNAL S8451 : STD_LOGIC;
    SIGNAL S8452 : STD_LOGIC;
    SIGNAL S8453 : STD_LOGIC;
    SIGNAL S8454 : STD_LOGIC;
    SIGNAL S8455 : STD_LOGIC;
    SIGNAL S8456 : STD_LOGIC;
    SIGNAL S8457 : STD_LOGIC;
    SIGNAL S8458 : STD_LOGIC;
    SIGNAL S8459 : STD_LOGIC;
    SIGNAL S8460 : STD_LOGIC;
    SIGNAL S8461 : STD_LOGIC;
    SIGNAL S8462 : STD_LOGIC;
    SIGNAL S8463 : STD_LOGIC;
    SIGNAL S8464 : STD_LOGIC;
    SIGNAL S8465 : STD_LOGIC;
    SIGNAL S8466 : STD_LOGIC;
    SIGNAL S8467 : STD_LOGIC;
    SIGNAL S8468 : STD_LOGIC;
    SIGNAL S8469 : STD_LOGIC;
    SIGNAL S8470 : STD_LOGIC;
    SIGNAL S8471 : STD_LOGIC;
    SIGNAL S8472 : STD_LOGIC;
    SIGNAL S8473 : STD_LOGIC;
    SIGNAL S8474 : STD_LOGIC;
    SIGNAL S8475 : STD_LOGIC;
    SIGNAL S8476 : STD_LOGIC;
    SIGNAL S8477 : STD_LOGIC;
    SIGNAL S8478 : STD_LOGIC;
    SIGNAL S8479 : STD_LOGIC;
    SIGNAL S8480 : STD_LOGIC;
    SIGNAL S8481 : STD_LOGIC;
    SIGNAL S8482 : STD_LOGIC;
    SIGNAL S8483 : STD_LOGIC;
    SIGNAL S8484 : STD_LOGIC;
    SIGNAL S8485 : STD_LOGIC;
    SIGNAL S8486 : STD_LOGIC;
    SIGNAL S8487 : STD_LOGIC;
    SIGNAL S8488 : STD_LOGIC;
    SIGNAL S8489 : STD_LOGIC;
    SIGNAL S8490 : STD_LOGIC;
    SIGNAL S8491 : STD_LOGIC;
    SIGNAL S8492 : STD_LOGIC;
    SIGNAL S8493 : STD_LOGIC;
    SIGNAL S8494 : STD_LOGIC;
    SIGNAL S8495 : STD_LOGIC;
    SIGNAL S8496 : STD_LOGIC;
    SIGNAL S8497 : STD_LOGIC;
    SIGNAL S8498 : STD_LOGIC;
    SIGNAL S8499 : STD_LOGIC;
    SIGNAL S8500 : STD_LOGIC;
    SIGNAL S8501 : STD_LOGIC;
    SIGNAL S8502 : STD_LOGIC;
    SIGNAL S8503 : STD_LOGIC;
    SIGNAL S8504 : STD_LOGIC;
    SIGNAL S8505 : STD_LOGIC;
    SIGNAL S8506 : STD_LOGIC;
    SIGNAL S8507 : STD_LOGIC;
    SIGNAL S8508 : STD_LOGIC;
    SIGNAL S8509 : STD_LOGIC;
    SIGNAL S8510 : STD_LOGIC;
    SIGNAL S8511 : STD_LOGIC;
    SIGNAL S8512 : STD_LOGIC;
    SIGNAL S8513 : STD_LOGIC;
    SIGNAL S8514 : STD_LOGIC;
    SIGNAL S8515 : STD_LOGIC;
    SIGNAL S8516 : STD_LOGIC;
    SIGNAL S8517 : STD_LOGIC;
    SIGNAL S8518 : STD_LOGIC;
    SIGNAL S8519 : STD_LOGIC;
    SIGNAL S8520 : STD_LOGIC;
    SIGNAL S8521 : STD_LOGIC;
    SIGNAL S8522 : STD_LOGIC;
    SIGNAL S8523 : STD_LOGIC;
    SIGNAL S8524 : STD_LOGIC;
    SIGNAL S8525 : STD_LOGIC;
    SIGNAL S8526 : STD_LOGIC;
    SIGNAL S8527 : STD_LOGIC;
    SIGNAL S8528 : STD_LOGIC;
    SIGNAL S8529 : STD_LOGIC;
    SIGNAL S8530 : STD_LOGIC;
    SIGNAL S8531 : STD_LOGIC;
    SIGNAL S8532 : STD_LOGIC;
    SIGNAL S8533 : STD_LOGIC;
    SIGNAL S8534 : STD_LOGIC;
    SIGNAL S8535 : STD_LOGIC;
    SIGNAL S8536 : STD_LOGIC;
    SIGNAL S8537 : STD_LOGIC;
    SIGNAL S8538 : STD_LOGIC;
    SIGNAL S8539 : STD_LOGIC;
    SIGNAL S8540 : STD_LOGIC;
    SIGNAL S8541 : STD_LOGIC;
    SIGNAL S8542 : STD_LOGIC;
    SIGNAL S8543 : STD_LOGIC;
    SIGNAL S8544 : STD_LOGIC;
    SIGNAL S8545 : STD_LOGIC;
    SIGNAL S8546 : STD_LOGIC;
    SIGNAL S8547 : STD_LOGIC;
    SIGNAL S8548 : STD_LOGIC;
    SIGNAL S8549 : STD_LOGIC;
    SIGNAL S8550 : STD_LOGIC;
    SIGNAL S8551 : STD_LOGIC;
    SIGNAL S8552 : STD_LOGIC;
    SIGNAL S8553 : STD_LOGIC;
    SIGNAL S8554 : STD_LOGIC;
    SIGNAL S8555 : STD_LOGIC;
    SIGNAL S8556 : STD_LOGIC;
    SIGNAL S8557 : STD_LOGIC;
    SIGNAL S8558 : STD_LOGIC;
    SIGNAL S8559 : STD_LOGIC;
    SIGNAL S8560 : STD_LOGIC;
    SIGNAL S8561 : STD_LOGIC;
    SIGNAL S8562 : STD_LOGIC;
    SIGNAL S8563 : STD_LOGIC;
    SIGNAL S8564 : STD_LOGIC;
    SIGNAL S8565 : STD_LOGIC;
    SIGNAL S8566 : STD_LOGIC;
    SIGNAL S8567 : STD_LOGIC;
    SIGNAL S8568 : STD_LOGIC;
    SIGNAL S8569 : STD_LOGIC;
    SIGNAL S8570 : STD_LOGIC;
    SIGNAL S8571 : STD_LOGIC;
    SIGNAL S8572 : STD_LOGIC;
    SIGNAL S8573 : STD_LOGIC;
    SIGNAL S8574 : STD_LOGIC;
    SIGNAL S8575 : STD_LOGIC;
    SIGNAL S8576 : STD_LOGIC;
    SIGNAL S8577 : STD_LOGIC;
    SIGNAL S8578 : STD_LOGIC;
    SIGNAL S8579 : STD_LOGIC;
    SIGNAL S8580 : STD_LOGIC;
    SIGNAL S8581 : STD_LOGIC;
    SIGNAL S8582 : STD_LOGIC;
    SIGNAL S8583 : STD_LOGIC;
    SIGNAL S8584 : STD_LOGIC;
    SIGNAL S8585 : STD_LOGIC;
    SIGNAL S8586 : STD_LOGIC;
    SIGNAL S8587 : STD_LOGIC;
    SIGNAL S8588 : STD_LOGIC;
    SIGNAL S8589 : STD_LOGIC;
    SIGNAL S8590 : STD_LOGIC;
    SIGNAL S8591 : STD_LOGIC;
    SIGNAL controller_1115_S_0 : STD_LOGIC;
    SIGNAL controller_1405_Y_0 : STD_LOGIC;
    SIGNAL controller_1405_Y_1 : STD_LOGIC;
    SIGNAL controller_216_B_0 : STD_LOGIC;
    SIGNAL controller_389_B_0 : STD_LOGIC;
    SIGNAL controller_389_B_2 : STD_LOGIC;
    SIGNAL controller_clk : STD_LOGIC;
    SIGNAL controller_fib_0 : STD_LOGIC;
    SIGNAL controller_fib_1 : STD_LOGIC;
    SIGNAL controller_fib_2 : STD_LOGIC;
    SIGNAL controller_fib_3 : STD_LOGIC;
    SIGNAL controller_fib_4 : STD_LOGIC;
    SIGNAL controller_opcode_2 : STD_LOGIC;
    SIGNAL controller_opcode_3 : STD_LOGIC;
    SIGNAL controller_opcode_4 : STD_LOGIC;
    SIGNAL controller_opcode_5 : STD_LOGIC;
    SIGNAL controller_opcode_6 : STD_LOGIC;
    SIGNAL controller_opcode_7 : STD_LOGIC;
    SIGNAL controller_outflag_0 : STD_LOGIC;
    SIGNAL controller_outflag_1 : STD_LOGIC;
    SIGNAL controller_outflag_2 : STD_LOGIC;
    SIGNAL controller_outflag_3 : STD_LOGIC;
    SIGNAL controller_outflag_6 : STD_LOGIC;
    SIGNAL controller_outflag_7 : STD_LOGIC;
    SIGNAL controller_pstate_0 : STD_LOGIC;
    SIGNAL controller_pstate_1 : STD_LOGIC;
    SIGNAL controller_readio : STD_LOGIC;
    SIGNAL controller_readmem : STD_LOGIC;
    SIGNAL controller_readymem : STD_LOGIC;
    SIGNAL controller_rst : STD_LOGIC;
    SIGNAL controller_writeio : STD_LOGIC;
    SIGNAL controller_writemem : STD_LOGIC;
    SIGNAL datapath_addrbus_0 : STD_LOGIC;
    SIGNAL datapath_addrbus_10 : STD_LOGIC;
    SIGNAL datapath_addrbus_11 : STD_LOGIC;
    SIGNAL datapath_addrbus_12 : STD_LOGIC;
    SIGNAL datapath_addrbus_13 : STD_LOGIC;
    SIGNAL datapath_addrbus_14 : STD_LOGIC;
    SIGNAL datapath_addrbus_15 : STD_LOGIC;
    SIGNAL datapath_addrbus_1 : STD_LOGIC;
    SIGNAL datapath_addrbus_2 : STD_LOGIC;
    SIGNAL datapath_addrbus_3 : STD_LOGIC;
    SIGNAL datapath_addrbus_4 : STD_LOGIC;
    SIGNAL datapath_addrbus_5 : STD_LOGIC;
    SIGNAL datapath_addrbus_6 : STD_LOGIC;
    SIGNAL datapath_addrbus_7 : STD_LOGIC;
    SIGNAL datapath_addrbus_8 : STD_LOGIC;
    SIGNAL datapath_addrbus_9 : STD_LOGIC;
    SIGNAL datapath_addsubunit_in1_0 : STD_LOGIC;
    SIGNAL datapath_addsubunit_in1_10 : STD_LOGIC;
    SIGNAL datapath_addsubunit_in1_11 : STD_LOGIC;
    SIGNAL datapath_addsubunit_in1_12 : STD_LOGIC;
    SIGNAL datapath_addsubunit_in1_13 : STD_LOGIC;
    SIGNAL datapath_addsubunit_in1_14 : STD_LOGIC;
    SIGNAL datapath_addsubunit_in1_15 : STD_LOGIC;
    SIGNAL datapath_addsubunit_in1_1 : STD_LOGIC;
    SIGNAL datapath_addsubunit_in1_2 : STD_LOGIC;
    SIGNAL datapath_addsubunit_in1_3 : STD_LOGIC;
    SIGNAL datapath_addsubunit_in1_4 : STD_LOGIC;
    SIGNAL datapath_addsubunit_in1_5 : STD_LOGIC;
    SIGNAL datapath_addsubunit_in1_6 : STD_LOGIC;
    SIGNAL datapath_addsubunit_in1_7 : STD_LOGIC;
    SIGNAL datapath_addsubunit_in1_8 : STD_LOGIC;
    SIGNAL datapath_addsubunit_in1_9 : STD_LOGIC;
    SIGNAL datapath_adr_outreg_0 : STD_LOGIC;
    SIGNAL datapath_adr_outreg_10 : STD_LOGIC;
    SIGNAL datapath_adr_outreg_11 : STD_LOGIC;
    SIGNAL datapath_adr_outreg_12 : STD_LOGIC;
    SIGNAL datapath_adr_outreg_13 : STD_LOGIC;
    SIGNAL datapath_adr_outreg_14 : STD_LOGIC;
    SIGNAL datapath_adr_outreg_15 : STD_LOGIC;
    SIGNAL datapath_adr_outreg_1 : STD_LOGIC;
    SIGNAL datapath_adr_outreg_2 : STD_LOGIC;
    SIGNAL datapath_adr_outreg_3 : STD_LOGIC;
    SIGNAL datapath_adr_outreg_4 : STD_LOGIC;
    SIGNAL datapath_adr_outreg_5 : STD_LOGIC;
    SIGNAL datapath_adr_outreg_6 : STD_LOGIC;
    SIGNAL datapath_adr_outreg_7 : STD_LOGIC;
    SIGNAL datapath_adr_outreg_8 : STD_LOGIC;
    SIGNAL datapath_adr_outreg_9 : STD_LOGIC;
    SIGNAL datapath_databusin_0 : STD_LOGIC;
    SIGNAL datapath_databusin_10 : STD_LOGIC;
    SIGNAL datapath_databusin_11 : STD_LOGIC;
    SIGNAL datapath_databusin_12 : STD_LOGIC;
    SIGNAL datapath_databusin_13 : STD_LOGIC;
    SIGNAL datapath_databusin_14 : STD_LOGIC;
    SIGNAL datapath_databusin_15 : STD_LOGIC;
    SIGNAL datapath_databusin_1 : STD_LOGIC;
    SIGNAL datapath_databusin_2 : STD_LOGIC;
    SIGNAL datapath_databusin_3 : STD_LOGIC;
    SIGNAL datapath_databusin_4 : STD_LOGIC;
    SIGNAL datapath_databusin_5 : STD_LOGIC;
    SIGNAL datapath_databusin_6 : STD_LOGIC;
    SIGNAL datapath_databusin_7 : STD_LOGIC;
    SIGNAL datapath_databusin_8 : STD_LOGIC;
    SIGNAL datapath_databusin_9 : STD_LOGIC;
    SIGNAL datapath_indatatrf_0 : STD_LOGIC;
    SIGNAL datapath_indatatrf_10 : STD_LOGIC;
    SIGNAL datapath_indatatrf_11 : STD_LOGIC;
    SIGNAL datapath_indatatrf_12 : STD_LOGIC;
    SIGNAL datapath_indatatrf_13 : STD_LOGIC;
    SIGNAL datapath_indatatrf_14 : STD_LOGIC;
    SIGNAL datapath_indatatrf_15 : STD_LOGIC;
    SIGNAL datapath_indatatrf_1 : STD_LOGIC;
    SIGNAL datapath_indatatrf_2 : STD_LOGIC;
    SIGNAL datapath_indatatrf_3 : STD_LOGIC;
    SIGNAL datapath_indatatrf_4 : STD_LOGIC;
    SIGNAL datapath_indatatrf_5 : STD_LOGIC;
    SIGNAL datapath_indatatrf_6 : STD_LOGIC;
    SIGNAL datapath_indatatrf_7 : STD_LOGIC;
    SIGNAL datapath_indatatrf_8 : STD_LOGIC;
    SIGNAL datapath_indatatrf_9 : STD_LOGIC;
    SIGNAL datapath_instruction_0 : STD_LOGIC;
    SIGNAL datapath_instruction_1 : STD_LOGIC;
    SIGNAL datapath_instruction_2 : STD_LOGIC;
    SIGNAL datapath_instruction_3 : STD_LOGIC;
    SIGNAL datapath_multdivunit_outmdu1_0 : STD_LOGIC;
    SIGNAL datapath_multdivunit_outmdu1_10 : STD_LOGIC;
    SIGNAL datapath_multdivunit_outmdu1_11 : STD_LOGIC;
    SIGNAL datapath_multdivunit_outmdu1_12 : STD_LOGIC;
    SIGNAL datapath_multdivunit_outmdu1_13 : STD_LOGIC;
    SIGNAL datapath_multdivunit_outmdu1_14 : STD_LOGIC;
    SIGNAL datapath_multdivunit_outmdu1_15 : STD_LOGIC;
    SIGNAL datapath_multdivunit_outmdu1_1 : STD_LOGIC;
    SIGNAL datapath_multdivunit_outmdu1_2 : STD_LOGIC;
    SIGNAL datapath_multdivunit_outmdu1_3 : STD_LOGIC;
    SIGNAL datapath_multdivunit_outmdu1_4 : STD_LOGIC;
    SIGNAL datapath_multdivunit_outmdu1_5 : STD_LOGIC;
    SIGNAL datapath_multdivunit_outmdu1_6 : STD_LOGIC;
    SIGNAL datapath_multdivunit_outmdu1_7 : STD_LOGIC;
    SIGNAL datapath_multdivunit_outmdu1_8 : STD_LOGIC;
    SIGNAL datapath_multdivunit_outmdu1_9 : STD_LOGIC;
    SIGNAL datapath_multdivunit_outmdu2_0 : STD_LOGIC;
    SIGNAL datapath_multdivunit_outmdu2_10 : STD_LOGIC;
    SIGNAL datapath_multdivunit_outmdu2_11 : STD_LOGIC;
    SIGNAL datapath_multdivunit_outmdu2_12 : STD_LOGIC;
    SIGNAL datapath_multdivunit_outmdu2_13 : STD_LOGIC;
    SIGNAL datapath_multdivunit_outmdu2_14 : STD_LOGIC;
    SIGNAL datapath_multdivunit_outmdu2_15 : STD_LOGIC;
    SIGNAL datapath_multdivunit_outmdu2_1 : STD_LOGIC;
    SIGNAL datapath_multdivunit_outmdu2_2 : STD_LOGIC;
    SIGNAL datapath_multdivunit_outmdu2_3 : STD_LOGIC;
    SIGNAL datapath_multdivunit_outmdu2_4 : STD_LOGIC;
    SIGNAL datapath_multdivunit_outmdu2_5 : STD_LOGIC;
    SIGNAL datapath_multdivunit_outmdu2_6 : STD_LOGIC;
    SIGNAL datapath_multdivunit_outmdu2_7 : STD_LOGIC;
    SIGNAL datapath_multdivunit_outmdu2_8 : STD_LOGIC;
    SIGNAL datapath_multdivunit_outmdu2_9 : STD_LOGIC;
    SIGNAL datapath_muxmem_in2_0 : STD_LOGIC;
    SIGNAL datapath_muxmem_in2_10 : STD_LOGIC;
    SIGNAL datapath_muxmem_in2_11 : STD_LOGIC;
    SIGNAL datapath_muxmem_in2_12 : STD_LOGIC;
    SIGNAL datapath_muxmem_in2_13 : STD_LOGIC;
    SIGNAL datapath_muxmem_in2_14 : STD_LOGIC;
    SIGNAL datapath_muxmem_in2_15 : STD_LOGIC;
    SIGNAL datapath_muxmem_in2_1 : STD_LOGIC;
    SIGNAL datapath_muxmem_in2_2 : STD_LOGIC;
    SIGNAL datapath_muxmem_in2_3 : STD_LOGIC;
    SIGNAL datapath_muxmem_in2_4 : STD_LOGIC;
    SIGNAL datapath_muxmem_in2_5 : STD_LOGIC;
    SIGNAL datapath_muxmem_in2_6 : STD_LOGIC;
    SIGNAL datapath_muxmem_in2_7 : STD_LOGIC;
    SIGNAL datapath_muxmem_in2_8 : STD_LOGIC;
    SIGNAL datapath_muxmem_in2_9 : STD_LOGIC;
    SIGNAL datapath_shiftunit_2135_A : STD_LOGIC;
    SIGNAL datapath_shiftunit_2153_A : STD_LOGIC;
    SIGNAL datapath_shiftunit_2171_A : STD_LOGIC;
    SIGNAL datapath_shiftunit_2189_A : STD_LOGIC;
    SIGNAL datapath_shiftunit_2207_A : STD_LOGIC;
    SIGNAL datapath_shiftunit_2225_A : STD_LOGIC;
    SIGNAL datapath_shiftunit_2243_A : STD_LOGIC;
    SIGNAL datapath_shiftunit_2261_A : STD_LOGIC;
    SIGNAL datapath_shiftunit_2279_A : STD_LOGIC;
    SIGNAL datapath_shiftunit_2297_A : STD_LOGIC;
    SIGNAL datapath_shiftunit_2315_A : STD_LOGIC;
    SIGNAL datapath_shiftunit_2333_A : STD_LOGIC;
    SIGNAL datapath_shiftunit_2351_A : STD_LOGIC;
    SIGNAL datapath_shiftunit_2369_A : STD_LOGIC;
    SIGNAL datapath_shiftunit_2387_A : STD_LOGIC;
    SIGNAL datapath_shiftunit_2405_A : STD_LOGIC;
    SIGNAL datapath_shiftunit_2439_A : STD_LOGIC;
    SIGNAL datapath_shiftunit_2457_A : STD_LOGIC;
    SIGNAL datapath_shiftunit_2475_A : STD_LOGIC;
    SIGNAL datapath_shiftunit_2493_A : STD_LOGIC;
    SIGNAL datapath_shiftunit_2511_A : STD_LOGIC;
    SIGNAL datapath_shiftunit_2529_A : STD_LOGIC;
    SIGNAL datapath_shiftunit_2547_A : STD_LOGIC;
    SIGNAL datapath_shiftunit_2565_A : STD_LOGIC;
    SIGNAL datapath_shiftunit_2583_A : STD_LOGIC;
    SIGNAL datapath_shiftunit_2601_A : STD_LOGIC;
    SIGNAL datapath_shiftunit_2619_A : STD_LOGIC;
    SIGNAL datapath_shiftunit_2637_A : STD_LOGIC;
    SIGNAL datapath_shiftunit_2655_A : STD_LOGIC;
    SIGNAL datapath_shiftunit_2673_A : STD_LOGIC;
    SIGNAL datapath_shiftunit_2691_A : STD_LOGIC;
    SIGNAL datapath_shiftunit_2708_A : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_0 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_100 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_101 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_102 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_103 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_104 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_105 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_106 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_107 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_108 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_109 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_10 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_110 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_111 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_112 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_113 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_114 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_115 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_116 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_117 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_118 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_119 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_11 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_120 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_121 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_122 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_123 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_124 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_125 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_126 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_127 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_128 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_129 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_12 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_130 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_131 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_132 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_133 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_134 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_135 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_136 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_137 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_138 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_139 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_13 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_140 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_141 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_142 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_143 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_144 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_145 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_146 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_147 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_148 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_149 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_14 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_150 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_151 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_152 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_153 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_154 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_155 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_156 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_157 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_158 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_159 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_15 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_160 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_161 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_162 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_163 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_164 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_165 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_166 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_167 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_168 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_169 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_16 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_170 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_171 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_172 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_173 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_174 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_175 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_176 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_177 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_178 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_179 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_17 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_180 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_181 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_182 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_183 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_184 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_185 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_186 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_187 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_188 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_189 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_18 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_190 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_191 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_192 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_193 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_194 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_195 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_196 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_197 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_198 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_199 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_19 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_1 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_200 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_201 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_202 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_203 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_204 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_205 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_206 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_207 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_208 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_209 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_20 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_210 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_211 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_212 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_213 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_214 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_215 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_216 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_217 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_218 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_219 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_21 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_220 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_221 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_222 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_223 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_224 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_225 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_226 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_227 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_228 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_229 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_22 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_230 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_231 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_232 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_233 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_234 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_235 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_236 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_237 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_238 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_239 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_23 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_240 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_241 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_242 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_243 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_244 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_245 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_246 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_247 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_248 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_249 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_24 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_250 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_251 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_252 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_253 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_254 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_255 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_25 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_26 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_27 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_28 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_29 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_2 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_30 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_31 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_32 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_33 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_34 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_35 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_36 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_37 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_38 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_39 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_3 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_40 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_41 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_42 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_43 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_44 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_45 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_46 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_47 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_48 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_49 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_4 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_50 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_51 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_52 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_53 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_54 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_55 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_56 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_57 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_58 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_59 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_5 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_60 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_61 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_62 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_63 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_64 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_65 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_66 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_67 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_68 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_69 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_6 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_70 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_71 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_72 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_73 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_74 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_75 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_76 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_77 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_78 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_79 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_7 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_80 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_81 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_82 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_83 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_84 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_85 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_86 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_87 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_88 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_89 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_8 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_90 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_91 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_92 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_93 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_94 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_95 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_96 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_97 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_98 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_99 : STD_LOGIC;
    SIGNAL datapath_theregisterfile_memtrf_9 : STD_LOGIC;

BEGIN
NOT_1: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_multdivunit_outmdu2_15,
        Y => S7476
    );
NOT_2: ENTITY WORK.NOT
    PORT MAP (
        A => controller_opcode_7,
        Y => S7487
    );
NOT_3: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_theregisterfile_memtrf_78,
        Y => S7498
    );
NOT_4: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_theregisterfile_memtrf_62,
        Y => S7509
    );
NOT_5: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_theregisterfile_memtrf_96,
        Y => S7520
    );
NOT_6: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_theregisterfile_memtrf_97,
        Y => S7531
    );
NOT_7: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_theregisterfile_memtrf_14,
        Y => S7542
    );
NOT_8: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_theregisterfile_memtrf_157,
        Y => S7553
    );
NOT_9: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_theregisterfile_memtrf_158,
        Y => S7564
    );
NOT_10: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_theregisterfile_memtrf_175,
        Y => S7574
    );
NOT_11: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_theregisterfile_memtrf_179,
        Y => S7585
    );
NOT_12: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_theregisterfile_memtrf_180,
        Y => S7596
    );
NOT_13: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_theregisterfile_memtrf_184,
        Y => S7607
    );
NOT_14: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_theregisterfile_memtrf_185,
        Y => S7618
    );
NOT_15: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_theregisterfile_memtrf_186,
        Y => S7629
    );
NOT_16: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_theregisterfile_memtrf_187,
        Y => S7640
    );
NOT_17: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_theregisterfile_memtrf_188,
        Y => S7651
    );
NOT_18: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_theregisterfile_memtrf_191,
        Y => S7662
    );
NOT_19: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_theregisterfile_memtrf_192,
        Y => S7673
    );
NOT_20: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_theregisterfile_memtrf_193,
        Y => S7684
    );
NOT_21: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_theregisterfile_memtrf_195,
        Y => S7695
    );
NOT_22: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_theregisterfile_memtrf_197,
        Y => S7706
    );
NOT_23: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_theregisterfile_memtrf_198,
        Y => S7717
    );
NOT_24: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_theregisterfile_memtrf_199,
        Y => S7728
    );
NOT_25: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_theregisterfile_memtrf_200,
        Y => S7739
    );
NOT_26: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_theregisterfile_memtrf_204,
        Y => S7750
    );
NOT_27: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_theregisterfile_memtrf_205,
        Y => S7761
    );
NOT_28: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_theregisterfile_memtrf_206,
        Y => S7772
    );
NOT_29: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_theregisterfile_memtrf_224,
        Y => S7783
    );
NOT_30: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_theregisterfile_memtrf_225,
        Y => S7794
    );
NOT_31: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_theregisterfile_memtrf_226,
        Y => S7805
    );
NOT_32: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_theregisterfile_memtrf_228,
        Y => S7816
    );
NOT_33: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_theregisterfile_memtrf_229,
        Y => S7822
    );
NOT_34: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_theregisterfile_memtrf_230,
        Y => S7823
    );
NOT_35: ENTITY WORK.NOT
    PORT MAP (
        A => controller_outflag_0,
        Y => S7830
    );
NOT_36: ENTITY WORK.NOT
    PORT MAP (
        A => controller_outflag_1,
        Y => S7838
    );
NOT_37: ENTITY WORK.NOT
    PORT MAP (
        A => controller_outflag_2,
        Y => S7846
    );
NOT_38: ENTITY WORK.NOT
    PORT MAP (
        A => controller_outflag_3,
        Y => S7853
    );
NOT_39: ENTITY WORK.NOT
    PORT MAP (
        A => controller_389_B_0,
        Y => S7861
    );
NOT_40: ENTITY WORK.NOT
    PORT MAP (
        A => controller_389_B_2,
        Y => S7869
    );
NOT_41: ENTITY WORK.NOT
    PORT MAP (
        A => controller_outflag_6,
        Y => S7876
    );
NOT_42: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_muxmem_in2_0,
        Y => S7884
    );
NOT_43: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_muxmem_in2_1,
        Y => S7892
    );
NOT_44: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_muxmem_in2_2,
        Y => S7897
    );
NOT_45: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_muxmem_in2_3,
        Y => S7905
    );
NOT_46: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_muxmem_in2_4,
        Y => S7913
    );
NOT_47: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_muxmem_in2_5,
        Y => S7920
    );
NOT_48: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_muxmem_in2_6,
        Y => S7928
    );
NOT_49: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_muxmem_in2_7,
        Y => S7936
    );
NOT_50: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_muxmem_in2_8,
        Y => S7946
    );
NOT_51: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_muxmem_in2_9,
        Y => S7957
    );
NOT_52: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_muxmem_in2_10,
        Y => S7968
    );
NOT_53: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_muxmem_in2_11,
        Y => S7978
    );
NOT_54: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_muxmem_in2_12,
        Y => S7989
    );
NOT_55: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_muxmem_in2_13,
        Y => S8000
    );
NOT_56: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_multdivunit_outmdu1_2,
        Y => S8011
    );
NOT_57: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_multdivunit_outmdu1_6,
        Y => S8022
    );
NOT_58: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_multdivunit_outmdu2_0,
        Y => S8033
    );
NOT_59: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_multdivunit_outmdu2_1,
        Y => S8044
    );
NOT_60: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_multdivunit_outmdu2_2,
        Y => S8054
    );
NOT_61: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_multdivunit_outmdu2_3,
        Y => S8065
    );
NOT_62: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_multdivunit_outmdu2_4,
        Y => S8076
    );
NOT_63: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_multdivunit_outmdu2_5,
        Y => S8087
    );
NOT_64: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_multdivunit_outmdu2_6,
        Y => S8097
    );
NOT_65: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_multdivunit_outmdu2_7,
        Y => S8108
    );
NOT_66: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_multdivunit_outmdu2_8,
        Y => S8119
    );
NOT_67: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_multdivunit_outmdu2_9,
        Y => S8129
    );
NOT_68: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_multdivunit_outmdu2_10,
        Y => S8140
    );
NOT_69: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_multdivunit_outmdu2_11,
        Y => S8151
    );
NOT_70: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_multdivunit_outmdu2_12,
        Y => S8161
    );
NOT_71: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_multdivunit_outmdu2_13,
        Y => S8172
    );
NOT_72: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_multdivunit_outmdu2_14,
        Y => S8183
    );
NOT_73: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_instruction_2,
        Y => S8193
    );
NOT_74: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_instruction_3,
        Y => S8204
    );
NOT_75: ENTITY WORK.NOT
    PORT MAP (
        A => controller_fib_0,
        Y => S8215
    );
NOT_76: ENTITY WORK.NOT
    PORT MAP (
        A => controller_fib_1,
        Y => S8225
    );
NOT_77: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_databusin_5,
        Y => S8236
    );
NOT_78: ENTITY WORK.NOT
    PORT MAP (
        A => controller_fib_2,
        Y => S8246
    );
NOT_79: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_databusin_6,
        Y => S8257
    );
NOT_80: ENTITY WORK.NOT
    PORT MAP (
        A => controller_fib_4,
        Y => S8267
    );
NOT_81: ENTITY WORK.NOT
    PORT MAP (
        A => controller_216_B_0,
        Y => S8278
    );
NOT_82: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_databusin_9,
        Y => S8288
    );
NOT_83: ENTITY WORK.NOT
    PORT MAP (
        A => controller_opcode_2,
        Y => S8299
    );
NOT_84: ENTITY WORK.NOT
    PORT MAP (
        A => controller_opcode_3,
        Y => S8309
    );
NOT_85: ENTITY WORK.NOT
    PORT MAP (
        A => controller_opcode_4,
        Y => S8319
    );
NOT_86: ENTITY WORK.NOT
    PORT MAP (
        A => controller_opcode_5,
        Y => S8329
    );
NOT_87: ENTITY WORK.NOT
    PORT MAP (
        A => controller_opcode_6,
        Y => S8339
    );
NOT_88: ENTITY WORK.NOT
    PORT MAP (
        A => controller_outflag_7,
        Y => S8349
    );
NOT_89: ENTITY WORK.NOT
    PORT MAP (
        A => controller_pstate_1,
        Y => S8356
    );
NOT_90: ENTITY WORK.NOT
    PORT MAP (
        A => controller_pstate_0,
        Y => S8365
    );
NOR_1: ENTITY WORK.NOR
    PORT MAP (
        A => controller_pstate_1,
        B => S8365,
        Y => S8375
    );
NAND_1: ENTITY WORK.NAND
    PORT MAP (
        A => S8356,
        B => controller_pstate_0,
        Y => S8385
    );
NOR_2: ENTITY WORK.NOR
    PORT MAP (
        A => S7487,
        B => S8339,
        Y => S8395
    );
NAND_2: ENTITY WORK.NAND
    PORT MAP (
        A => controller_opcode_7,
        B => controller_opcode_6,
        Y => S8405
    );
NOR_3: ENTITY WORK.NOR
    PORT MAP (
        A => controller_opcode_4,
        B => controller_opcode_5,
        Y => S8416
    );
NAND_3: ENTITY WORK.NAND
    PORT MAP (
        A => S8319,
        B => S8329,
        Y => S8426
    );
NOR_4: ENTITY WORK.NOR
    PORT MAP (
        A => S8405,
        B => S8416,
        Y => S8436
    );
NOT_91: ENTITY WORK.NOT
    PORT MAP (
        A => S8436,
        Y => S8447
    );
NOR_5: ENTITY WORK.NOR
    PORT MAP (
        A => S8319,
        B => S8329,
        Y => S8457
    );
NAND_4: ENTITY WORK.NAND
    PORT MAP (
        A => controller_opcode_4,
        B => controller_opcode_5,
        Y => S8468
    );
NOR_6: ENTITY WORK.NOR
    PORT MAP (
        A => controller_opcode_7,
        B => controller_opcode_6,
        Y => S8478
    );
NAND_5: ENTITY WORK.NAND
    PORT MAP (
        A => S7487,
        B => S8339,
        Y => S8489
    );
NAND_6: ENTITY WORK.NAND
    PORT MAP (
        A => S8468,
        B => S8478,
        Y => S8499
    );
NAND_7: ENTITY WORK.NAND
    PORT MAP (
        A => S8447,
        B => S8499,
        Y => S8510
    );
NOT_92: ENTITY WORK.NOT
    PORT MAP (
        A => S8510,
        Y => S8520
    );
NOR_7: ENTITY WORK.NOR
    PORT MAP (
        A => controller_opcode_5,
        B => S8489,
        Y => S8531
    );
NOR_8: ENTITY WORK.NOR
    PORT MAP (
        A => controller_opcode_2,
        B => S8309,
        Y => S8541
    );
NAND_8: ENTITY WORK.NAND
    PORT MAP (
        A => S8299,
        B => controller_opcode_3,
        Y => S8542
    );
NOR_9: ENTITY WORK.NOR
    PORT MAP (
        A => S8405,
        B => S8468,
        Y => S8543
    );
NAND_9: ENTITY WORK.NAND
    PORT MAP (
        A => S8395,
        B => S8457,
        Y => S8544
    );
NAND_10: ENTITY WORK.NAND
    PORT MAP (
        A => S8541,
        B => S8543,
        Y => S8545
    );
NOT_93: ENTITY WORK.NOT
    PORT MAP (
        A => S8545,
        Y => S8546
    );
NAND_11: ENTITY WORK.NAND
    PORT MAP (
        A => S8510,
        B => S8545,
        Y => S8547
    );
NOR_10: ENTITY WORK.NOR
    PORT MAP (
        A => S8531,
        B => S8547,
        Y => S8548
    );
NOT_94: ENTITY WORK.NOT
    PORT MAP (
        A => S8548,
        Y => S8549
    );
NOR_11: ENTITY WORK.NOR
    PORT MAP (
        A => S8299,
        B => controller_opcode_3,
        Y => S8550
    );
NAND_12: ENTITY WORK.NAND
    PORT MAP (
        A => controller_opcode_2,
        B => S8309,
        Y => S8551
    );
NAND_13: ENTITY WORK.NAND
    PORT MAP (
        A => controller_fib_1,
        B => controller_fib_2,
        Y => S8552
    );
NOR_12: ENTITY WORK.NOR
    PORT MAP (
        A => S8551,
        B => S8552,
        Y => S8553
    );
NAND_14: ENTITY WORK.NAND
    PORT MAP (
        A => S8542,
        B => S8543,
        Y => S8554
    );
NOR_13: ENTITY WORK.NOR
    PORT MAP (
        A => S8553,
        B => S8554,
        Y => S8555
    );
NOR_14: ENTITY WORK.NOR
    PORT MAP (
        A => controller_opcode_4,
        B => S8329,
        Y => S8556
    );
NAND_15: ENTITY WORK.NAND
    PORT MAP (
        A => S8319,
        B => controller_opcode_5,
        Y => S8557
    );
NOR_15: ENTITY WORK.NOR
    PORT MAP (
        A => S8489,
        B => S8557,
        Y => S8558
    );
NAND_16: ENTITY WORK.NAND
    PORT MAP (
        A => S8478,
        B => S8556,
        Y => S8559
    );
NAND_17: ENTITY WORK.NAND
    PORT MAP (
        A => controller_opcode_3,
        B => S8558,
        Y => S8560
    );
NAND_18: ENTITY WORK.NAND
    PORT MAP (
        A => S8548,
        B => S8560,
        Y => S8561
    );
NOR_16: ENTITY WORK.NOR
    PORT MAP (
        A => S8555,
        B => S8561,
        Y => S8562
    );
NOR_17: ENTITY WORK.NOR
    PORT MAP (
        A => S8385,
        B => S8562,
        Y => S8563
    );
NOR_18: ENTITY WORK.NOR
    PORT MAP (
        A => S8416,
        B => S8457,
        Y => S8564
    );
NAND_19: ENTITY WORK.NAND
    PORT MAP (
        A => S8426,
        B => S8468,
        Y => S8565
    );
NAND_20: ENTITY WORK.NAND
    PORT MAP (
        A => controller_pstate_1,
        B => S8436,
        Y => S8566
    );
NOT_95: ENTITY WORK.NOT
    PORT MAP (
        A => S8566,
        Y => S8567
    );
NOR_19: ENTITY WORK.NOR
    PORT MAP (
        A => S8457,
        B => S8566,
        Y => S8568
    );
NAND_21: ENTITY WORK.NAND
    PORT MAP (
        A => S8468,
        B => S8567,
        Y => S8569
    );
NOR_20: ENTITY WORK.NOR
    PORT MAP (
        A => S8365,
        B => S8569,
        Y => S8570
    );
NAND_22: ENTITY WORK.NAND
    PORT MAP (
        A => controller_pstate_0,
        B => S8568,
        Y => S8571
    );
NOR_21: ENTITY WORK.NOR
    PORT MAP (
        A => controller_216_B_0,
        B => controller_readymem,
        Y => S8572
    );
NOT_96: ENTITY WORK.NOT
    PORT MAP (
        A => S8572,
        Y => S8573
    );
NOR_22: ENTITY WORK.NOR
    PORT MAP (
        A => controller_opcode_3,
        B => S8356,
        Y => S8574
    );
NAND_23: ENTITY WORK.NAND
    PORT MAP (
        A => S8365,
        B => S8574,
        Y => S8575
    );
NOR_23: ENTITY WORK.NOR
    PORT MAP (
        A => S8559,
        B => S8575,
        Y => S8576
    );
NOT_97: ENTITY WORK.NOT
    PORT MAP (
        A => S8576,
        Y => S8577
    );
NAND_24: ENTITY WORK.NAND
    PORT MAP (
        A => S8573,
        B => S8576,
        Y => S8578
    );
NAND_25: ENTITY WORK.NAND
    PORT MAP (
        A => S8571,
        B => S8578,
        Y => S8579
    );
NOR_24: ENTITY WORK.NOR
    PORT MAP (
        A => S8563,
        B => S8579,
        Y => S8580
    );
NAND_26: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_15,
        B => S8580,
        Y => S8581
    );
NAND_27: ENTITY WORK.NAND
    PORT MAP (
        A => controller_216_B_0,
        B => S8543,
        Y => S8582
    );
NAND_28: ENTITY WORK.NAND
    PORT MAP (
        A => controller_fib_0,
        B => controller_fib_2,
        Y => S8583
    );
NOR_25: ENTITY WORK.NOR
    PORT MAP (
        A => controller_fib_1,
        B => S8583,
        Y => S8584
    );
NAND_29: ENTITY WORK.NAND
    PORT MAP (
        A => S7861,
        B => S8584,
        Y => S8585
    );
NOR_26: ENTITY WORK.NOR
    PORT MAP (
        A => S8225,
        B => controller_fib_2,
        Y => S8586
    );
NOR_27: ENTITY WORK.NOR
    PORT MAP (
        A => controller_389_B_0,
        B => controller_389_B_2,
        Y => S8587
    );
NOR_28: ENTITY WORK.NOR
    PORT MAP (
        A => controller_389_B_2,
        B => controller_fib_0,
        Y => S8588
    );
NOT_98: ENTITY WORK.NOT
    PORT MAP (
        A => S8588,
        Y => S8589
    );
NAND_30: ENTITY WORK.NAND
    PORT MAP (
        A => S8586,
        B => S8589,
        Y => S8590
    );
NOR_29: ENTITY WORK.NOR
    PORT MAP (
        A => S8587,
        B => S8590,
        Y => S8591
    );
NOR_30: ENTITY WORK.NOR
    PORT MAP (
        A => S8215,
        B => controller_fib_2,
        Y => S344
    );
NAND_31: ENTITY WORK.NAND
    PORT MAP (
        A => controller_fib_0,
        B => S8246,
        Y => S345
    );
NOR_31: ENTITY WORK.NOR
    PORT MAP (
        A => controller_fib_1,
        B => S345,
        Y => S346
    );
NOR_32: ENTITY WORK.NOR
    PORT MAP (
        A => controller_fib_0,
        B => controller_fib_1,
        Y => S347
    );
NAND_32: ENTITY WORK.NAND
    PORT MAP (
        A => controller_fib_2,
        B => S347,
        Y => S348
    );
NOT_99: ENTITY WORK.NOT
    PORT MAP (
        A => S348,
        Y => S349
    );
NOR_33: ENTITY WORK.NOR
    PORT MAP (
        A => S346,
        B => S349,
        Y => S350
    );
NOR_34: ENTITY WORK.NOR
    PORT MAP (
        A => controller_389_B_2,
        B => S350,
        Y => S351
    );
NOR_35: ENTITY WORK.NOR
    PORT MAP (
        A => controller_389_B_0,
        B => S351,
        Y => S352
    );
NAND_33: ENTITY WORK.NAND
    PORT MAP (
        A => S8246,
        B => S347,
        Y => S353
    );
NOR_36: ENTITY WORK.NOR
    PORT MAP (
        A => S7861,
        B => S347,
        Y => S354
    );
NOR_37: ENTITY WORK.NOR
    PORT MAP (
        A => S352,
        B => S354,
        Y => S355
    );
NOR_38: ENTITY WORK.NOR
    PORT MAP (
        A => S8591,
        B => S355,
        Y => S356
    );
NAND_34: ENTITY WORK.NAND
    PORT MAP (
        A => S8585,
        B => S356,
        Y => S357
    );
NAND_35: ENTITY WORK.NAND
    PORT MAP (
        A => S8550,
        B => S357,
        Y => S358
    );
NOT_100: ENTITY WORK.NOT
    PORT MAP (
        A => S358,
        Y => S359
    );
NOR_39: ENTITY WORK.NOR
    PORT MAP (
        A => S8551,
        B => S8582,
        Y => S360
    );
NOT_101: ENTITY WORK.NOT
    PORT MAP (
        A => S360,
        Y => S361
    );
NAND_36: ENTITY WORK.NAND
    PORT MAP (
        A => S357,
        B => S360,
        Y => S362
    );
NAND_37: ENTITY WORK.NAND
    PORT MAP (
        A => S8560,
        B => S362,
        Y => S363
    );
NAND_38: ENTITY WORK.NAND
    PORT MAP (
        A => S8375,
        B => S363,
        Y => S364
    );
NOT_102: ENTITY WORK.NOT
    PORT MAP (
        A => S364,
        Y => S365
    );
NAND_39: ENTITY WORK.NAND
    PORT MAP (
        A => controller_opcode_2,
        B => controller_opcode_3,
        Y => S366
    );
NOT_103: ENTITY WORK.NOT
    PORT MAP (
        A => S366,
        Y => S367
    );
NOR_40: ENTITY WORK.NOR
    PORT MAP (
        A => S8385,
        B => S8559,
        Y => S368
    );
NAND_40: ENTITY WORK.NAND
    PORT MAP (
        A => S8375,
        B => S8558,
        Y => S369
    );
NOR_41: ENTITY WORK.NOR
    PORT MAP (
        A => S366,
        B => S369,
        Y => S370
    );
NOT_104: ENTITY WORK.NOT
    PORT MAP (
        A => S370,
        Y => S371
    );
NAND_41: ENTITY WORK.NAND
    PORT MAP (
        A => controller_216_B_0,
        B => S370,
        Y => S372
    );
NOR_42: ENTITY WORK.NOR
    PORT MAP (
        A => S8541,
        B => S8550,
        Y => S373
    );
NAND_42: ENTITY WORK.NAND
    PORT MAP (
        A => controller_216_B_0,
        B => S373,
        Y => S374
    );
NAND_43: ENTITY WORK.NAND
    PORT MAP (
        A => S358,
        B => S374,
        Y => S375
    );
NOR_43: ENTITY WORK.NOR
    PORT MAP (
        A => S8385,
        B => S8405,
        Y => S376
    );
NAND_44: ENTITY WORK.NAND
    PORT MAP (
        A => S8375,
        B => S8395,
        Y => S377
    );
NAND_45: ENTITY WORK.NAND
    PORT MAP (
        A => controller_opcode_4,
        B => S8375,
        Y => S378
    );
NOR_44: ENTITY WORK.NOR
    PORT MAP (
        A => S8385,
        B => S8544,
        Y => S379
    );
NAND_46: ENTITY WORK.NAND
    PORT MAP (
        A => S8375,
        B => S8543,
        Y => S380
    );
NAND_47: ENTITY WORK.NAND
    PORT MAP (
        A => S375,
        B => S379,
        Y => S381
    );
NOR_45: ENTITY WORK.NOR
    PORT MAP (
        A => controller_opcode_7,
        B => S8339,
        Y => S382
    );
NAND_48: ENTITY WORK.NAND
    PORT MAP (
        A => S7487,
        B => controller_opcode_6,
        Y => S383
    );
NOR_46: ENTITY WORK.NOR
    PORT MAP (
        A => S8557,
        B => S383,
        Y => S384
    );
NOR_47: ENTITY WORK.NOR
    PORT MAP (
        A => S8546,
        B => S384,
        Y => S385
    );
NOR_48: ENTITY WORK.NOR
    PORT MAP (
        A => S8551,
        B => S8559,
        Y => S386
    );
NAND_49: ENTITY WORK.NAND
    PORT MAP (
        A => controller_opcode_7,
        B => S8339,
        Y => S387
    );
NOR_49: ENTITY WORK.NOR
    PORT MAP (
        A => S8319,
        B => S387,
        Y => S388
    );
NOR_50: ENTITY WORK.NOR
    PORT MAP (
        A => S8468,
        B => S387,
        Y => S389
    );
NOT_105: ENTITY WORK.NOT
    PORT MAP (
        A => S389,
        Y => S390
    );
NAND_50: ENTITY WORK.NAND
    PORT MAP (
        A => controller_opcode_6,
        B => S8416,
        Y => S391
    );
NAND_51: ENTITY WORK.NAND
    PORT MAP (
        A => S390,
        B => S391,
        Y => S392
    );
NOR_51: ENTITY WORK.NOR
    PORT MAP (
        A => S386,
        B => S392,
        Y => S393
    );
NAND_52: ENTITY WORK.NAND
    PORT MAP (
        A => S385,
        B => S393,
        Y => S394
    );
NAND_53: ENTITY WORK.NAND
    PORT MAP (
        A => S8375,
        B => S394,
        Y => S395
    );
NAND_54: ENTITY WORK.NAND
    PORT MAP (
        A => S381,
        B => S395,
        Y => S396
    );
NAND_55: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_instruction_2,
        B => S396,
        Y => S397
    );
NOT_106: ENTITY WORK.NOT
    PORT MAP (
        A => S397,
        Y => S398
    );
NOR_52: ENTITY WORK.NOR
    PORT MAP (
        A => controller_opcode_2,
        B => S8559,
        Y => S399
    );
NOR_53: ENTITY WORK.NOR
    PORT MAP (
        A => controller_216_B_0,
        B => S8544,
        Y => S400
    );
NAND_56: ENTITY WORK.NAND
    PORT MAP (
        A => S8278,
        B => S8543,
        Y => S401
    );
NAND_57: ENTITY WORK.NAND
    PORT MAP (
        A => S373,
        B => S400,
        Y => S402
    );
NAND_58: ENTITY WORK.NAND
    PORT MAP (
        A => controller_opcode_2,
        B => S8576,
        Y => S403
    );
NOR_54: ENTITY WORK.NOR
    PORT MAP (
        A => controller_opcode_7,
        B => S8468,
        Y => S404
    );
NOT_107: ENTITY WORK.NOT
    PORT MAP (
        A => S404,
        Y => S405
    );
NAND_59: ENTITY WORK.NAND
    PORT MAP (
        A => controller_opcode_7,
        B => S8468,
        Y => S406
    );
NOT_108: ENTITY WORK.NOT
    PORT MAP (
        A => S406,
        Y => S407
    );
NOR_55: ENTITY WORK.NOR
    PORT MAP (
        A => S404,
        B => S407,
        Y => S408
    );
NOR_56: ENTITY WORK.NOR
    PORT MAP (
        A => S8405,
        B => S8426,
        Y => S409
    );
NAND_60: ENTITY WORK.NAND
    PORT MAP (
        A => S8395,
        B => S8416,
        Y => S410
    );
NAND_61: ENTITY WORK.NAND
    PORT MAP (
        A => S8375,
        B => S410,
        Y => S411
    );
NAND_62: ENTITY WORK.NAND
    PORT MAP (
        A => S391,
        B => S407,
        Y => S412
    );
NAND_63: ENTITY WORK.NAND
    PORT MAP (
        A => S405,
        B => S412,
        Y => S413
    );
NOR_57: ENTITY WORK.NOR
    PORT MAP (
        A => S408,
        B => S411,
        Y => S414
    );
NAND_64: ENTITY WORK.NAND
    PORT MAP (
        A => S8375,
        B => S413,
        Y => S415
    );
NOR_58: ENTITY WORK.NOR
    PORT MAP (
        A => S399,
        B => S413,
        Y => S416
    );
NAND_65: ENTITY WORK.NAND
    PORT MAP (
        A => S402,
        B => S416,
        Y => S417
    );
NAND_66: ENTITY WORK.NAND
    PORT MAP (
        A => S8375,
        B => S417,
        Y => S418
    );
NAND_67: ENTITY WORK.NAND
    PORT MAP (
        A => S403,
        B => S418,
        Y => S419
    );
NAND_68: ENTITY WORK.NAND
    PORT MAP (
        A => controller_fib_2,
        B => S419,
        Y => S420
    );
NOT_109: ENTITY WORK.NOT
    PORT MAP (
        A => S420,
        Y => S421
    );
NOR_59: ENTITY WORK.NOR
    PORT MAP (
        A => S398,
        B => S421,
        Y => S422
    );
NAND_69: ENTITY WORK.NAND
    PORT MAP (
        A => S397,
        B => S420,
        Y => S423
    );
NAND_70: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_instruction_3,
        B => S396,
        Y => S424
    );
NOT_110: ENTITY WORK.NOT
    PORT MAP (
        A => S424,
        Y => S425
    );
NAND_71: ENTITY WORK.NAND
    PORT MAP (
        A => controller_fib_3,
        B => S419,
        Y => S426
    );
NOT_111: ENTITY WORK.NOT
    PORT MAP (
        A => S426,
        Y => S427
    );
NOR_60: ENTITY WORK.NOR
    PORT MAP (
        A => S425,
        B => S427,
        Y => S428
    );
NOR_61: ENTITY WORK.NOR
    PORT MAP (
        A => S422,
        B => S428,
        Y => S429
    );
NOT_112: ENTITY WORK.NOT
    PORT MAP (
        A => S429,
        Y => S430
    );
NAND_72: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_instruction_0,
        B => S396,
        Y => S431
    );
NOT_113: ENTITY WORK.NOT
    PORT MAP (
        A => S431,
        Y => S432
    );
NAND_73: ENTITY WORK.NAND
    PORT MAP (
        A => controller_fib_0,
        B => S419,
        Y => S433
    );
NOT_114: ENTITY WORK.NOT
    PORT MAP (
        A => S433,
        Y => S434
    );
NOR_62: ENTITY WORK.NOR
    PORT MAP (
        A => S432,
        B => S434,
        Y => S435
    );
NAND_74: ENTITY WORK.NAND
    PORT MAP (
        A => S431,
        B => S433,
        Y => S436
    );
NAND_75: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_instruction_1,
        B => S396,
        Y => S437
    );
NOT_115: ENTITY WORK.NOT
    PORT MAP (
        A => S437,
        Y => S438
    );
NAND_76: ENTITY WORK.NAND
    PORT MAP (
        A => controller_fib_1,
        B => S419,
        Y => S439
    );
NOT_116: ENTITY WORK.NOT
    PORT MAP (
        A => S439,
        Y => S440
    );
NOR_63: ENTITY WORK.NOR
    PORT MAP (
        A => S438,
        B => S440,
        Y => S441
    );
NAND_77: ENTITY WORK.NAND
    PORT MAP (
        A => S437,
        B => S439,
        Y => S442
    );
NOR_64: ENTITY WORK.NOR
    PORT MAP (
        A => S435,
        B => S441,
        Y => S443
    );
NAND_78: ENTITY WORK.NAND
    PORT MAP (
        A => S429,
        B => S442,
        Y => S444
    );
NOR_65: ENTITY WORK.NOR
    PORT MAP (
        A => S435,
        B => S444,
        Y => S445
    );
NAND_79: ENTITY WORK.NAND
    PORT MAP (
        A => S429,
        B => S443,
        Y => S446
    );
NAND_80: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_238,
        B => S436,
        Y => S447
    );
NAND_81: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_254,
        B => S435,
        Y => S448
    );
NAND_82: ENTITY WORK.NAND
    PORT MAP (
        A => S447,
        B => S448,
        Y => S449
    );
NAND_83: ENTITY WORK.NAND
    PORT MAP (
        A => S422,
        B => S449,
        Y => S450
    );
NAND_84: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_174,
        B => S436,
        Y => S451
    );
NAND_85: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_190,
        B => S435,
        Y => S452
    );
NAND_86: ENTITY WORK.NAND
    PORT MAP (
        A => S451,
        B => S452,
        Y => S453
    );
NAND_87: ENTITY WORK.NAND
    PORT MAP (
        A => S423,
        B => S453,
        Y => S454
    );
NAND_88: ENTITY WORK.NAND
    PORT MAP (
        A => S450,
        B => S454,
        Y => S455
    );
NOR_66: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_222,
        B => S423,
        Y => S456
    );
NAND_89: ENTITY WORK.NAND
    PORT MAP (
        A => S7564,
        B => S423,
        Y => S457
    );
NAND_90: ENTITY WORK.NAND
    PORT MAP (
        A => S435,
        B => S457,
        Y => S458
    );
NOR_67: ENTITY WORK.NOR
    PORT MAP (
        A => S456,
        B => S458,
        Y => S459
    );
NOR_68: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_142,
        B => S422,
        Y => S460
    );
NAND_91: ENTITY WORK.NAND
    PORT MAP (
        A => S7772,
        B => S422,
        Y => S461
    );
NAND_92: ENTITY WORK.NAND
    PORT MAP (
        A => S436,
        B => S461,
        Y => S462
    );
NOR_69: ENTITY WORK.NOR
    PORT MAP (
        A => S460,
        B => S462,
        Y => S463
    );
NOR_70: ENTITY WORK.NOR
    PORT MAP (
        A => S459,
        B => S463,
        Y => S464
    );
NAND_93: ENTITY WORK.NAND
    PORT MAP (
        A => S442,
        B => S464,
        Y => S465
    );
NOR_71: ENTITY WORK.NOR
    PORT MAP (
        A => S442,
        B => S455,
        Y => S466
    );
NAND_94: ENTITY WORK.NAND
    PORT MAP (
        A => S428,
        B => S465,
        Y => S467
    );
NOR_72: ENTITY WORK.NOR
    PORT MAP (
        A => S466,
        B => S467,
        Y => S468
    );
NAND_95: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_62,
        B => S435,
        Y => S469
    );
NAND_96: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_46,
        B => S436,
        Y => S470
    );
NAND_97: ENTITY WORK.NAND
    PORT MAP (
        A => S469,
        B => S470,
        Y => S471
    );
NAND_98: ENTITY WORK.NAND
    PORT MAP (
        A => S441,
        B => S471,
        Y => S472
    );
NAND_99: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_30,
        B => S435,
        Y => S473
    );
NAND_100: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_14,
        B => S436,
        Y => S474
    );
NAND_101: ENTITY WORK.NAND
    PORT MAP (
        A => S473,
        B => S474,
        Y => S475
    );
NAND_102: ENTITY WORK.NAND
    PORT MAP (
        A => S442,
        B => S475,
        Y => S476
    );
NAND_103: ENTITY WORK.NAND
    PORT MAP (
        A => S472,
        B => S476,
        Y => S477
    );
NAND_104: ENTITY WORK.NAND
    PORT MAP (
        A => S429,
        B => S477,
        Y => S478
    );
NOR_73: ENTITY WORK.NOR
    PORT MAP (
        A => S423,
        B => S428,
        Y => S479
    );
NAND_105: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_126,
        B => S435,
        Y => S480
    );
NAND_106: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_110,
        B => S436,
        Y => S481
    );
NAND_107: ENTITY WORK.NAND
    PORT MAP (
        A => S480,
        B => S481,
        Y => S482
    );
NAND_108: ENTITY WORK.NAND
    PORT MAP (
        A => S441,
        B => S482,
        Y => S483
    );
NAND_109: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_94,
        B => S435,
        Y => S484
    );
NAND_110: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_78,
        B => S436,
        Y => S485
    );
NAND_111: ENTITY WORK.NAND
    PORT MAP (
        A => S484,
        B => S485,
        Y => S486
    );
NAND_112: ENTITY WORK.NAND
    PORT MAP (
        A => S442,
        B => S486,
        Y => S487
    );
NAND_113: ENTITY WORK.NAND
    PORT MAP (
        A => S483,
        B => S487,
        Y => S488
    );
NAND_114: ENTITY WORK.NAND
    PORT MAP (
        A => S479,
        B => S488,
        Y => S489
    );
NAND_115: ENTITY WORK.NAND
    PORT MAP (
        A => S478,
        B => S489,
        Y => S490
    );
NOR_74: ENTITY WORK.NOR
    PORT MAP (
        A => S468,
        B => S490,
        Y => S491
    );
NOR_75: ENTITY WORK.NOR
    PORT MAP (
        A => S445,
        B => S491,
        Y => datapath_addsubunit_in1_14
    );
NOT_117: ENTITY WORK.NOT
    PORT MAP (
        A => datapath_addsubunit_in1_14,
        Y => S492
    );
NAND_116: ENTITY WORK.NAND
    PORT MAP (
        A => S366,
        B => S368,
        Y => S493
    );
NOR_76: ENTITY WORK.NOR
    PORT MAP (
        A => S356,
        B => S361,
        Y => S494
    );
NAND_117: ENTITY WORK.NAND
    PORT MAP (
        A => S8375,
        B => S494,
        Y => S495
    );
NAND_118: ENTITY WORK.NAND
    PORT MAP (
        A => S493,
        B => S495,
        Y => S496
    );
NAND_119: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_14,
        B => S496,
        Y => S497
    );
NAND_120: ENTITY WORK.NAND
    PORT MAP (
        A => S372,
        B => S497,
        Y => S498
    );
NAND_121: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_14,
        B => S498,
        Y => S499
    );
NOT_118: ENTITY WORK.NOT
    PORT MAP (
        A => S499,
        Y => S500
    );
NOR_77: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_muxmem_in2_14,
        B => S498,
        Y => S501
    );
NOR_78: ENTITY WORK.NOR
    PORT MAP (
        A => S500,
        B => S501,
        Y => S502
    );
NAND_122: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_237,
        B => S436,
        Y => S503
    );
NAND_123: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_253,
        B => S435,
        Y => S504
    );
NAND_124: ENTITY WORK.NAND
    PORT MAP (
        A => S503,
        B => S504,
        Y => S505
    );
NAND_125: ENTITY WORK.NAND
    PORT MAP (
        A => S422,
        B => S505,
        Y => S506
    );
NAND_126: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_173,
        B => S436,
        Y => S507
    );
NAND_127: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_189,
        B => S435,
        Y => S508
    );
NAND_128: ENTITY WORK.NAND
    PORT MAP (
        A => S507,
        B => S508,
        Y => S509
    );
NAND_129: ENTITY WORK.NAND
    PORT MAP (
        A => S423,
        B => S509,
        Y => S510
    );
NAND_130: ENTITY WORK.NAND
    PORT MAP (
        A => S506,
        B => S510,
        Y => S511
    );
NOR_79: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_221,
        B => S423,
        Y => S512
    );
NAND_131: ENTITY WORK.NAND
    PORT MAP (
        A => S7553,
        B => S423,
        Y => S513
    );
NAND_132: ENTITY WORK.NAND
    PORT MAP (
        A => S435,
        B => S513,
        Y => S514
    );
NOR_80: ENTITY WORK.NOR
    PORT MAP (
        A => S512,
        B => S514,
        Y => S515
    );
NOR_81: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_141,
        B => S422,
        Y => S516
    );
NAND_133: ENTITY WORK.NAND
    PORT MAP (
        A => S7761,
        B => S422,
        Y => S517
    );
NAND_134: ENTITY WORK.NAND
    PORT MAP (
        A => S436,
        B => S517,
        Y => S518
    );
NOR_82: ENTITY WORK.NOR
    PORT MAP (
        A => S516,
        B => S518,
        Y => S519
    );
NOR_83: ENTITY WORK.NOR
    PORT MAP (
        A => S515,
        B => S519,
        Y => S520
    );
NAND_135: ENTITY WORK.NAND
    PORT MAP (
        A => S442,
        B => S520,
        Y => S521
    );
NOR_84: ENTITY WORK.NOR
    PORT MAP (
        A => S442,
        B => S511,
        Y => S522
    );
NAND_136: ENTITY WORK.NAND
    PORT MAP (
        A => S428,
        B => S521,
        Y => S523
    );
NOR_85: ENTITY WORK.NOR
    PORT MAP (
        A => S522,
        B => S523,
        Y => S524
    );
NAND_137: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_61,
        B => S435,
        Y => S525
    );
NAND_138: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_45,
        B => S436,
        Y => S526
    );
NAND_139: ENTITY WORK.NAND
    PORT MAP (
        A => S525,
        B => S526,
        Y => S527
    );
NAND_140: ENTITY WORK.NAND
    PORT MAP (
        A => S441,
        B => S527,
        Y => S528
    );
NAND_141: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_29,
        B => S435,
        Y => S529
    );
NAND_142: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_13,
        B => S436,
        Y => S530
    );
NAND_143: ENTITY WORK.NAND
    PORT MAP (
        A => S529,
        B => S530,
        Y => S531
    );
NAND_144: ENTITY WORK.NAND
    PORT MAP (
        A => S442,
        B => S531,
        Y => S532
    );
NAND_145: ENTITY WORK.NAND
    PORT MAP (
        A => S528,
        B => S532,
        Y => S533
    );
NAND_146: ENTITY WORK.NAND
    PORT MAP (
        A => S429,
        B => S533,
        Y => S534
    );
NAND_147: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_125,
        B => S435,
        Y => S535
    );
NAND_148: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_109,
        B => S436,
        Y => S536
    );
NAND_149: ENTITY WORK.NAND
    PORT MAP (
        A => S535,
        B => S536,
        Y => S537
    );
NAND_150: ENTITY WORK.NAND
    PORT MAP (
        A => S441,
        B => S537,
        Y => S538
    );
NAND_151: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_93,
        B => S435,
        Y => S539
    );
NAND_152: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_77,
        B => S436,
        Y => S540
    );
NAND_153: ENTITY WORK.NAND
    PORT MAP (
        A => S539,
        B => S540,
        Y => S541
    );
NAND_154: ENTITY WORK.NAND
    PORT MAP (
        A => S442,
        B => S541,
        Y => S542
    );
NAND_155: ENTITY WORK.NAND
    PORT MAP (
        A => S538,
        B => S542,
        Y => S543
    );
NAND_156: ENTITY WORK.NAND
    PORT MAP (
        A => S479,
        B => S543,
        Y => S544
    );
NOT_119: ENTITY WORK.NOT
    PORT MAP (
        A => S544,
        Y => S545
    );
NOR_86: ENTITY WORK.NOR
    PORT MAP (
        A => S524,
        B => S545,
        Y => S546
    );
NAND_157: ENTITY WORK.NAND
    PORT MAP (
        A => S534,
        B => S546,
        Y => S547
    );
NAND_158: ENTITY WORK.NAND
    PORT MAP (
        A => S446,
        B => S547,
        Y => S548
    );
NOT_120: ENTITY WORK.NOT
    PORT MAP (
        A => S548,
        Y => datapath_addsubunit_in1_13
    );
NAND_159: ENTITY WORK.NAND
    PORT MAP (
        A => S496,
        B => datapath_addsubunit_in1_13,
        Y => S549
    );
NAND_160: ENTITY WORK.NAND
    PORT MAP (
        A => S372,
        B => S549,
        Y => S550
    );
NOT_121: ENTITY WORK.NOT
    PORT MAP (
        A => S550,
        Y => S551
    );
NOR_87: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_muxmem_in2_13,
        B => S550,
        Y => S552
    );
NOR_88: ENTITY WORK.NOR
    PORT MAP (
        A => S8000,
        B => S551,
        Y => S553
    );
NOR_89: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_172,
        B => S422,
        Y => S554
    );
NOR_90: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_236,
        B => S423,
        Y => S555
    );
NOR_91: ENTITY WORK.NOR
    PORT MAP (
        A => S554,
        B => S555,
        Y => S556
    );
NAND_161: ENTITY WORK.NAND
    PORT MAP (
        A => S436,
        B => S556,
        Y => S557
    );
NOR_92: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_252,
        B => S423,
        Y => S558
    );
NAND_162: ENTITY WORK.NAND
    PORT MAP (
        A => S7651,
        B => S423,
        Y => S559
    );
NAND_163: ENTITY WORK.NAND
    PORT MAP (
        A => S435,
        B => S559,
        Y => S560
    );
NOR_93: ENTITY WORK.NOR
    PORT MAP (
        A => S558,
        B => S560,
        Y => S561
    );
NAND_164: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_204,
        B => S436,
        Y => S562
    );
NAND_165: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_220,
        B => S435,
        Y => S563
    );
NAND_166: ENTITY WORK.NAND
    PORT MAP (
        A => S562,
        B => S563,
        Y => S564
    );
NAND_167: ENTITY WORK.NAND
    PORT MAP (
        A => S422,
        B => S564,
        Y => S565
    );
NAND_168: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_140,
        B => S436,
        Y => S566
    );
NAND_169: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_156,
        B => S435,
        Y => S567
    );
NAND_170: ENTITY WORK.NAND
    PORT MAP (
        A => S566,
        B => S567,
        Y => S568
    );
NAND_171: ENTITY WORK.NAND
    PORT MAP (
        A => S423,
        B => S568,
        Y => S569
    );
NAND_172: ENTITY WORK.NAND
    PORT MAP (
        A => S565,
        B => S569,
        Y => S570
    );
NOR_94: ENTITY WORK.NOR
    PORT MAP (
        A => S441,
        B => S570,
        Y => S571
    );
NOR_95: ENTITY WORK.NOR
    PORT MAP (
        A => S442,
        B => S561,
        Y => S572
    );
NAND_173: ENTITY WORK.NAND
    PORT MAP (
        A => S557,
        B => S572,
        Y => S573
    );
NAND_174: ENTITY WORK.NAND
    PORT MAP (
        A => S428,
        B => S573,
        Y => S574
    );
NOR_96: ENTITY WORK.NOR
    PORT MAP (
        A => S571,
        B => S574,
        Y => S575
    );
NAND_175: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_124,
        B => S435,
        Y => S576
    );
NAND_176: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_108,
        B => S436,
        Y => S577
    );
NAND_177: ENTITY WORK.NAND
    PORT MAP (
        A => S576,
        B => S577,
        Y => S578
    );
NAND_178: ENTITY WORK.NAND
    PORT MAP (
        A => S441,
        B => S578,
        Y => S579
    );
NAND_179: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_92,
        B => S435,
        Y => S580
    );
NAND_180: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_76,
        B => S436,
        Y => S581
    );
NAND_181: ENTITY WORK.NAND
    PORT MAP (
        A => S580,
        B => S581,
        Y => S582
    );
NAND_182: ENTITY WORK.NAND
    PORT MAP (
        A => S442,
        B => S582,
        Y => S583
    );
NAND_183: ENTITY WORK.NAND
    PORT MAP (
        A => S579,
        B => S583,
        Y => S584
    );
NAND_184: ENTITY WORK.NAND
    PORT MAP (
        A => S479,
        B => S584,
        Y => S585
    );
NAND_185: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_60,
        B => S435,
        Y => S586
    );
NAND_186: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_44,
        B => S436,
        Y => S587
    );
NAND_187: ENTITY WORK.NAND
    PORT MAP (
        A => S586,
        B => S587,
        Y => S588
    );
NAND_188: ENTITY WORK.NAND
    PORT MAP (
        A => S441,
        B => S588,
        Y => S589
    );
NAND_189: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_28,
        B => S435,
        Y => S590
    );
NAND_190: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_12,
        B => S436,
        Y => S591
    );
NAND_191: ENTITY WORK.NAND
    PORT MAP (
        A => S590,
        B => S591,
        Y => S592
    );
NAND_192: ENTITY WORK.NAND
    PORT MAP (
        A => S442,
        B => S592,
        Y => S593
    );
NAND_193: ENTITY WORK.NAND
    PORT MAP (
        A => S589,
        B => S593,
        Y => S594
    );
NAND_194: ENTITY WORK.NAND
    PORT MAP (
        A => S429,
        B => S594,
        Y => S595
    );
NOT_122: ENTITY WORK.NOT
    PORT MAP (
        A => S595,
        Y => S596
    );
NOR_97: ENTITY WORK.NOR
    PORT MAP (
        A => S575,
        B => S596,
        Y => S597
    );
NAND_195: ENTITY WORK.NAND
    PORT MAP (
        A => S585,
        B => S597,
        Y => S598
    );
NAND_196: ENTITY WORK.NAND
    PORT MAP (
        A => S446,
        B => S598,
        Y => S599
    );
NOT_123: ENTITY WORK.NOT
    PORT MAP (
        A => S599,
        Y => datapath_addsubunit_in1_12
    );
NAND_197: ENTITY WORK.NAND
    PORT MAP (
        A => S496,
        B => datapath_addsubunit_in1_12,
        Y => S600
    );
NAND_198: ENTITY WORK.NAND
    PORT MAP (
        A => S372,
        B => S600,
        Y => S601
    );
NAND_199: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_12,
        B => S601,
        Y => S602
    );
NOT_124: ENTITY WORK.NOT
    PORT MAP (
        A => S602,
        Y => S603
    );
NOR_98: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_muxmem_in2_12,
        B => S601,
        Y => S604
    );
NOR_99: ENTITY WORK.NOR
    PORT MAP (
        A => S603,
        B => S604,
        Y => S605
    );
NOR_100: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_171,
        B => S422,
        Y => S606
    );
NOR_101: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_235,
        B => S423,
        Y => S607
    );
NOR_102: ENTITY WORK.NOR
    PORT MAP (
        A => S606,
        B => S607,
        Y => S608
    );
NAND_200: ENTITY WORK.NAND
    PORT MAP (
        A => S436,
        B => S608,
        Y => S609
    );
NOR_103: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_251,
        B => S423,
        Y => S610
    );
NAND_201: ENTITY WORK.NAND
    PORT MAP (
        A => S7640,
        B => S423,
        Y => S611
    );
NAND_202: ENTITY WORK.NAND
    PORT MAP (
        A => S435,
        B => S611,
        Y => S612
    );
NOR_104: ENTITY WORK.NOR
    PORT MAP (
        A => S610,
        B => S612,
        Y => S613
    );
NAND_203: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_203,
        B => S436,
        Y => S614
    );
NAND_204: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_219,
        B => S435,
        Y => S615
    );
NAND_205: ENTITY WORK.NAND
    PORT MAP (
        A => S614,
        B => S615,
        Y => S616
    );
NAND_206: ENTITY WORK.NAND
    PORT MAP (
        A => S422,
        B => S616,
        Y => S617
    );
NAND_207: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_139,
        B => S436,
        Y => S618
    );
NAND_208: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_155,
        B => S435,
        Y => S619
    );
NAND_209: ENTITY WORK.NAND
    PORT MAP (
        A => S618,
        B => S619,
        Y => S620
    );
NAND_210: ENTITY WORK.NAND
    PORT MAP (
        A => S423,
        B => S620,
        Y => S621
    );
NAND_211: ENTITY WORK.NAND
    PORT MAP (
        A => S617,
        B => S621,
        Y => S622
    );
NOR_105: ENTITY WORK.NOR
    PORT MAP (
        A => S441,
        B => S622,
        Y => S623
    );
NOR_106: ENTITY WORK.NOR
    PORT MAP (
        A => S442,
        B => S613,
        Y => S624
    );
NAND_212: ENTITY WORK.NAND
    PORT MAP (
        A => S609,
        B => S624,
        Y => S625
    );
NAND_213: ENTITY WORK.NAND
    PORT MAP (
        A => S428,
        B => S625,
        Y => S626
    );
NOR_107: ENTITY WORK.NOR
    PORT MAP (
        A => S623,
        B => S626,
        Y => S627
    );
NAND_214: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_59,
        B => S435,
        Y => S628
    );
NAND_215: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_43,
        B => S436,
        Y => S629
    );
NAND_216: ENTITY WORK.NAND
    PORT MAP (
        A => S628,
        B => S629,
        Y => S630
    );
NAND_217: ENTITY WORK.NAND
    PORT MAP (
        A => S441,
        B => S630,
        Y => S631
    );
NAND_218: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_27,
        B => S435,
        Y => S632
    );
NAND_219: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_11,
        B => S436,
        Y => S633
    );
NAND_220: ENTITY WORK.NAND
    PORT MAP (
        A => S632,
        B => S633,
        Y => S634
    );
NAND_221: ENTITY WORK.NAND
    PORT MAP (
        A => S442,
        B => S634,
        Y => S635
    );
NAND_222: ENTITY WORK.NAND
    PORT MAP (
        A => S631,
        B => S635,
        Y => S636
    );
NAND_223: ENTITY WORK.NAND
    PORT MAP (
        A => S429,
        B => S636,
        Y => S637
    );
NAND_224: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_123,
        B => S435,
        Y => S638
    );
NAND_225: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_107,
        B => S436,
        Y => S639
    );
NAND_226: ENTITY WORK.NAND
    PORT MAP (
        A => S638,
        B => S639,
        Y => S640
    );
NAND_227: ENTITY WORK.NAND
    PORT MAP (
        A => S441,
        B => S640,
        Y => S641
    );
NAND_228: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_91,
        B => S435,
        Y => S642
    );
NAND_229: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_75,
        B => S436,
        Y => S643
    );
NAND_230: ENTITY WORK.NAND
    PORT MAP (
        A => S642,
        B => S643,
        Y => S644
    );
NAND_231: ENTITY WORK.NAND
    PORT MAP (
        A => S442,
        B => S644,
        Y => S645
    );
NAND_232: ENTITY WORK.NAND
    PORT MAP (
        A => S641,
        B => S645,
        Y => S646
    );
NAND_233: ENTITY WORK.NAND
    PORT MAP (
        A => S479,
        B => S646,
        Y => S647
    );
NOT_125: ENTITY WORK.NOT
    PORT MAP (
        A => S647,
        Y => S648
    );
NOR_108: ENTITY WORK.NOR
    PORT MAP (
        A => S627,
        B => S648,
        Y => S649
    );
NAND_234: ENTITY WORK.NAND
    PORT MAP (
        A => S637,
        B => S649,
        Y => S650
    );
NAND_235: ENTITY WORK.NAND
    PORT MAP (
        A => S446,
        B => S650,
        Y => S651
    );
NOT_126: ENTITY WORK.NOT
    PORT MAP (
        A => S651,
        Y => datapath_addsubunit_in1_11
    );
NAND_236: ENTITY WORK.NAND
    PORT MAP (
        A => S496,
        B => datapath_addsubunit_in1_11,
        Y => S652
    );
NAND_237: ENTITY WORK.NAND
    PORT MAP (
        A => S372,
        B => S652,
        Y => S653
    );
NOT_127: ENTITY WORK.NOT
    PORT MAP (
        A => S653,
        Y => S654
    );
NOR_109: ENTITY WORK.NOR
    PORT MAP (
        A => S7978,
        B => S654,
        Y => S655
    );
NOR_110: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_muxmem_in2_11,
        B => S653,
        Y => S656
    );
NOR_111: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_170,
        B => S422,
        Y => S657
    );
NOR_112: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_234,
        B => S423,
        Y => S658
    );
NOR_113: ENTITY WORK.NOR
    PORT MAP (
        A => S657,
        B => S658,
        Y => S659
    );
NAND_238: ENTITY WORK.NAND
    PORT MAP (
        A => S436,
        B => S659,
        Y => S660
    );
NOR_114: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_250,
        B => S423,
        Y => S661
    );
NAND_239: ENTITY WORK.NAND
    PORT MAP (
        A => S7629,
        B => S423,
        Y => S662
    );
NAND_240: ENTITY WORK.NAND
    PORT MAP (
        A => S435,
        B => S662,
        Y => S663
    );
NOR_115: ENTITY WORK.NOR
    PORT MAP (
        A => S661,
        B => S663,
        Y => S664
    );
NAND_241: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_202,
        B => S436,
        Y => S665
    );
NAND_242: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_218,
        B => S435,
        Y => S666
    );
NAND_243: ENTITY WORK.NAND
    PORT MAP (
        A => S665,
        B => S666,
        Y => S667
    );
NAND_244: ENTITY WORK.NAND
    PORT MAP (
        A => S422,
        B => S667,
        Y => S668
    );
NAND_245: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_138,
        B => S436,
        Y => S669
    );
NAND_246: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_154,
        B => S435,
        Y => S670
    );
NAND_247: ENTITY WORK.NAND
    PORT MAP (
        A => S669,
        B => S670,
        Y => S671
    );
NAND_248: ENTITY WORK.NAND
    PORT MAP (
        A => S423,
        B => S671,
        Y => S672
    );
NAND_249: ENTITY WORK.NAND
    PORT MAP (
        A => S668,
        B => S672,
        Y => S673
    );
NOR_116: ENTITY WORK.NOR
    PORT MAP (
        A => S441,
        B => S673,
        Y => S674
    );
NOR_117: ENTITY WORK.NOR
    PORT MAP (
        A => S442,
        B => S664,
        Y => S675
    );
NAND_250: ENTITY WORK.NAND
    PORT MAP (
        A => S660,
        B => S675,
        Y => S676
    );
NAND_251: ENTITY WORK.NAND
    PORT MAP (
        A => S428,
        B => S676,
        Y => S677
    );
NOR_118: ENTITY WORK.NOR
    PORT MAP (
        A => S674,
        B => S677,
        Y => S678
    );
NAND_252: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_122,
        B => S435,
        Y => S679
    );
NAND_253: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_106,
        B => S436,
        Y => S680
    );
NAND_254: ENTITY WORK.NAND
    PORT MAP (
        A => S679,
        B => S680,
        Y => S681
    );
NAND_255: ENTITY WORK.NAND
    PORT MAP (
        A => S441,
        B => S681,
        Y => S682
    );
NAND_256: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_90,
        B => S435,
        Y => S683
    );
NAND_257: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_74,
        B => S436,
        Y => S684
    );
NAND_258: ENTITY WORK.NAND
    PORT MAP (
        A => S683,
        B => S684,
        Y => S685
    );
NAND_259: ENTITY WORK.NAND
    PORT MAP (
        A => S442,
        B => S685,
        Y => S686
    );
NAND_260: ENTITY WORK.NAND
    PORT MAP (
        A => S682,
        B => S686,
        Y => S687
    );
NAND_261: ENTITY WORK.NAND
    PORT MAP (
        A => S479,
        B => S687,
        Y => S688
    );
NAND_262: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_58,
        B => S435,
        Y => S689
    );
NAND_263: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_42,
        B => S436,
        Y => S690
    );
NAND_264: ENTITY WORK.NAND
    PORT MAP (
        A => S689,
        B => S690,
        Y => S691
    );
NAND_265: ENTITY WORK.NAND
    PORT MAP (
        A => S441,
        B => S691,
        Y => S692
    );
NAND_266: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_26,
        B => S435,
        Y => S693
    );
NAND_267: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_10,
        B => S436,
        Y => S694
    );
NAND_268: ENTITY WORK.NAND
    PORT MAP (
        A => S693,
        B => S694,
        Y => S695
    );
NAND_269: ENTITY WORK.NAND
    PORT MAP (
        A => S442,
        B => S695,
        Y => S696
    );
NAND_270: ENTITY WORK.NAND
    PORT MAP (
        A => S692,
        B => S696,
        Y => S697
    );
NAND_271: ENTITY WORK.NAND
    PORT MAP (
        A => S429,
        B => S697,
        Y => S698
    );
NOT_128: ENTITY WORK.NOT
    PORT MAP (
        A => S698,
        Y => S699
    );
NOR_119: ENTITY WORK.NOR
    PORT MAP (
        A => S678,
        B => S699,
        Y => S700
    );
NAND_272: ENTITY WORK.NAND
    PORT MAP (
        A => S688,
        B => S700,
        Y => S701
    );
NAND_273: ENTITY WORK.NAND
    PORT MAP (
        A => S446,
        B => S701,
        Y => S702
    );
NOT_129: ENTITY WORK.NOT
    PORT MAP (
        A => S702,
        Y => datapath_addsubunit_in1_10
    );
NAND_274: ENTITY WORK.NAND
    PORT MAP (
        A => S496,
        B => datapath_addsubunit_in1_10,
        Y => S703
    );
NAND_275: ENTITY WORK.NAND
    PORT MAP (
        A => S372,
        B => S703,
        Y => S704
    );
NAND_276: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_10,
        B => S704,
        Y => S705
    );
NOT_130: ENTITY WORK.NOT
    PORT MAP (
        A => S705,
        Y => S706
    );
NOR_120: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_muxmem_in2_10,
        B => S704,
        Y => S707
    );
NOR_121: ENTITY WORK.NOR
    PORT MAP (
        A => S706,
        B => S707,
        Y => S708
    );
NOR_122: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_169,
        B => S422,
        Y => S709
    );
NOR_123: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_233,
        B => S423,
        Y => S710
    );
NOR_124: ENTITY WORK.NOR
    PORT MAP (
        A => S709,
        B => S710,
        Y => S711
    );
NAND_277: ENTITY WORK.NAND
    PORT MAP (
        A => S436,
        B => S711,
        Y => S712
    );
NOR_125: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_249,
        B => S423,
        Y => S713
    );
NAND_278: ENTITY WORK.NAND
    PORT MAP (
        A => S7618,
        B => S423,
        Y => S714
    );
NAND_279: ENTITY WORK.NAND
    PORT MAP (
        A => S435,
        B => S714,
        Y => S715
    );
NOR_126: ENTITY WORK.NOR
    PORT MAP (
        A => S713,
        B => S715,
        Y => S716
    );
NAND_280: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_201,
        B => S436,
        Y => S717
    );
NAND_281: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_217,
        B => S435,
        Y => S718
    );
NAND_282: ENTITY WORK.NAND
    PORT MAP (
        A => S717,
        B => S718,
        Y => S719
    );
NAND_283: ENTITY WORK.NAND
    PORT MAP (
        A => S422,
        B => S719,
        Y => S720
    );
NAND_284: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_137,
        B => S436,
        Y => S721
    );
NAND_285: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_153,
        B => S435,
        Y => S722
    );
NAND_286: ENTITY WORK.NAND
    PORT MAP (
        A => S721,
        B => S722,
        Y => S723
    );
NAND_287: ENTITY WORK.NAND
    PORT MAP (
        A => S423,
        B => S723,
        Y => S724
    );
NAND_288: ENTITY WORK.NAND
    PORT MAP (
        A => S720,
        B => S724,
        Y => S725
    );
NOR_127: ENTITY WORK.NOR
    PORT MAP (
        A => S441,
        B => S725,
        Y => S726
    );
NOR_128: ENTITY WORK.NOR
    PORT MAP (
        A => S442,
        B => S716,
        Y => S727
    );
NAND_289: ENTITY WORK.NAND
    PORT MAP (
        A => S712,
        B => S727,
        Y => S728
    );
NAND_290: ENTITY WORK.NAND
    PORT MAP (
        A => S428,
        B => S728,
        Y => S729
    );
NOR_129: ENTITY WORK.NOR
    PORT MAP (
        A => S726,
        B => S729,
        Y => S730
    );
NAND_291: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_121,
        B => S435,
        Y => S731
    );
NAND_292: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_105,
        B => S436,
        Y => S732
    );
NAND_293: ENTITY WORK.NAND
    PORT MAP (
        A => S731,
        B => S732,
        Y => S733
    );
NAND_294: ENTITY WORK.NAND
    PORT MAP (
        A => S441,
        B => S733,
        Y => S734
    );
NAND_295: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_89,
        B => S435,
        Y => S735
    );
NAND_296: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_73,
        B => S436,
        Y => S736
    );
NAND_297: ENTITY WORK.NAND
    PORT MAP (
        A => S735,
        B => S736,
        Y => S737
    );
NAND_298: ENTITY WORK.NAND
    PORT MAP (
        A => S442,
        B => S737,
        Y => S738
    );
NAND_299: ENTITY WORK.NAND
    PORT MAP (
        A => S734,
        B => S738,
        Y => S739
    );
NAND_300: ENTITY WORK.NAND
    PORT MAP (
        A => S479,
        B => S739,
        Y => S740
    );
NAND_301: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_57,
        B => S435,
        Y => S741
    );
NAND_302: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_41,
        B => S436,
        Y => S742
    );
NAND_303: ENTITY WORK.NAND
    PORT MAP (
        A => S741,
        B => S742,
        Y => S743
    );
NAND_304: ENTITY WORK.NAND
    PORT MAP (
        A => S441,
        B => S743,
        Y => S744
    );
NAND_305: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_25,
        B => S435,
        Y => S745
    );
NAND_306: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_9,
        B => S436,
        Y => S746
    );
NAND_307: ENTITY WORK.NAND
    PORT MAP (
        A => S745,
        B => S746,
        Y => S747
    );
NAND_308: ENTITY WORK.NAND
    PORT MAP (
        A => S442,
        B => S747,
        Y => S748
    );
NAND_309: ENTITY WORK.NAND
    PORT MAP (
        A => S744,
        B => S748,
        Y => S749
    );
NAND_310: ENTITY WORK.NAND
    PORT MAP (
        A => S429,
        B => S749,
        Y => S750
    );
NOT_131: ENTITY WORK.NOT
    PORT MAP (
        A => S750,
        Y => S751
    );
NOR_130: ENTITY WORK.NOR
    PORT MAP (
        A => S730,
        B => S751,
        Y => S752
    );
NAND_311: ENTITY WORK.NAND
    PORT MAP (
        A => S740,
        B => S752,
        Y => S753
    );
NAND_312: ENTITY WORK.NAND
    PORT MAP (
        A => S446,
        B => S753,
        Y => S754
    );
NOT_132: ENTITY WORK.NOT
    PORT MAP (
        A => S754,
        Y => datapath_addsubunit_in1_9
    );
NAND_313: ENTITY WORK.NAND
    PORT MAP (
        A => S496,
        B => datapath_addsubunit_in1_9,
        Y => S755
    );
NAND_314: ENTITY WORK.NAND
    PORT MAP (
        A => S372,
        B => S755,
        Y => S756
    );
NOT_133: ENTITY WORK.NOT
    PORT MAP (
        A => S756,
        Y => S757
    );
NOR_131: ENTITY WORK.NOR
    PORT MAP (
        A => S7957,
        B => S757,
        Y => S758
    );
NOR_132: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_muxmem_in2_9,
        B => S756,
        Y => S759
    );
NOR_133: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_168,
        B => S422,
        Y => S760
    );
NOR_134: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_232,
        B => S423,
        Y => S761
    );
NOR_135: ENTITY WORK.NOR
    PORT MAP (
        A => S760,
        B => S761,
        Y => S762
    );
NAND_315: ENTITY WORK.NAND
    PORT MAP (
        A => S436,
        B => S762,
        Y => S763
    );
NOR_136: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_248,
        B => S423,
        Y => S764
    );
NAND_316: ENTITY WORK.NAND
    PORT MAP (
        A => S7607,
        B => S423,
        Y => S765
    );
NAND_317: ENTITY WORK.NAND
    PORT MAP (
        A => S435,
        B => S765,
        Y => S766
    );
NOR_137: ENTITY WORK.NOR
    PORT MAP (
        A => S764,
        B => S766,
        Y => S767
    );
NAND_318: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_200,
        B => S436,
        Y => S768
    );
NAND_319: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_216,
        B => S435,
        Y => S769
    );
NAND_320: ENTITY WORK.NAND
    PORT MAP (
        A => S768,
        B => S769,
        Y => S770
    );
NAND_321: ENTITY WORK.NAND
    PORT MAP (
        A => S422,
        B => S770,
        Y => S771
    );
NAND_322: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_136,
        B => S436,
        Y => S772
    );
NAND_323: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_152,
        B => S435,
        Y => S773
    );
NAND_324: ENTITY WORK.NAND
    PORT MAP (
        A => S772,
        B => S773,
        Y => S774
    );
NAND_325: ENTITY WORK.NAND
    PORT MAP (
        A => S423,
        B => S774,
        Y => S775
    );
NAND_326: ENTITY WORK.NAND
    PORT MAP (
        A => S771,
        B => S775,
        Y => S776
    );
NOR_138: ENTITY WORK.NOR
    PORT MAP (
        A => S441,
        B => S776,
        Y => S777
    );
NOR_139: ENTITY WORK.NOR
    PORT MAP (
        A => S442,
        B => S767,
        Y => S778
    );
NAND_327: ENTITY WORK.NAND
    PORT MAP (
        A => S763,
        B => S778,
        Y => S779
    );
NAND_328: ENTITY WORK.NAND
    PORT MAP (
        A => S428,
        B => S779,
        Y => S780
    );
NOR_140: ENTITY WORK.NOR
    PORT MAP (
        A => S777,
        B => S780,
        Y => S781
    );
NAND_329: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_120,
        B => S435,
        Y => S782
    );
NAND_330: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_104,
        B => S436,
        Y => S783
    );
NAND_331: ENTITY WORK.NAND
    PORT MAP (
        A => S782,
        B => S783,
        Y => S784
    );
NAND_332: ENTITY WORK.NAND
    PORT MAP (
        A => S441,
        B => S784,
        Y => S785
    );
NAND_333: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_88,
        B => S435,
        Y => S786
    );
NAND_334: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_72,
        B => S436,
        Y => S787
    );
NAND_335: ENTITY WORK.NAND
    PORT MAP (
        A => S786,
        B => S787,
        Y => S788
    );
NAND_336: ENTITY WORK.NAND
    PORT MAP (
        A => S442,
        B => S788,
        Y => S789
    );
NAND_337: ENTITY WORK.NAND
    PORT MAP (
        A => S785,
        B => S789,
        Y => S790
    );
NAND_338: ENTITY WORK.NAND
    PORT MAP (
        A => S479,
        B => S790,
        Y => S791
    );
NAND_339: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_56,
        B => S435,
        Y => S792
    );
NAND_340: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_40,
        B => S436,
        Y => S793
    );
NAND_341: ENTITY WORK.NAND
    PORT MAP (
        A => S792,
        B => S793,
        Y => S794
    );
NAND_342: ENTITY WORK.NAND
    PORT MAP (
        A => S441,
        B => S794,
        Y => S795
    );
NAND_343: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_24,
        B => S435,
        Y => S796
    );
NAND_344: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_8,
        B => S436,
        Y => S797
    );
NAND_345: ENTITY WORK.NAND
    PORT MAP (
        A => S796,
        B => S797,
        Y => S798
    );
NAND_346: ENTITY WORK.NAND
    PORT MAP (
        A => S442,
        B => S798,
        Y => S799
    );
NAND_347: ENTITY WORK.NAND
    PORT MAP (
        A => S795,
        B => S799,
        Y => S800
    );
NAND_348: ENTITY WORK.NAND
    PORT MAP (
        A => S429,
        B => S800,
        Y => S801
    );
NOT_134: ENTITY WORK.NOT
    PORT MAP (
        A => S801,
        Y => S802
    );
NOR_141: ENTITY WORK.NOR
    PORT MAP (
        A => S781,
        B => S802,
        Y => S803
    );
NAND_349: ENTITY WORK.NAND
    PORT MAP (
        A => S791,
        B => S803,
        Y => S804
    );
NAND_350: ENTITY WORK.NAND
    PORT MAP (
        A => S446,
        B => S804,
        Y => S805
    );
NOT_135: ENTITY WORK.NOT
    PORT MAP (
        A => S805,
        Y => datapath_addsubunit_in1_8
    );
NAND_351: ENTITY WORK.NAND
    PORT MAP (
        A => S496,
        B => datapath_addsubunit_in1_8,
        Y => S806
    );
NAND_352: ENTITY WORK.NAND
    PORT MAP (
        A => S372,
        B => S806,
        Y => S807
    );
NAND_353: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_8,
        B => S807,
        Y => S808
    );
NOT_136: ENTITY WORK.NOT
    PORT MAP (
        A => S808,
        Y => S809
    );
NOR_142: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_muxmem_in2_8,
        B => S807,
        Y => S810
    );
NOR_143: ENTITY WORK.NOR
    PORT MAP (
        A => S809,
        B => S810,
        Y => S811
    );
NAND_354: ENTITY WORK.NAND
    PORT MAP (
        A => S8349,
        B => S445,
        Y => S812
    );
NAND_355: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_183,
        B => S423,
        Y => S813
    );
NAND_356: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_247,
        B => S422,
        Y => S814
    );
NAND_357: ENTITY WORK.NAND
    PORT MAP (
        A => S813,
        B => S814,
        Y => S815
    );
NAND_358: ENTITY WORK.NAND
    PORT MAP (
        A => S435,
        B => S815,
        Y => S816
    );
NOR_144: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_167,
        B => S422,
        Y => S817
    );
NOR_145: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_231,
        B => S423,
        Y => S818
    );
NOR_146: ENTITY WORK.NOR
    PORT MAP (
        A => S817,
        B => S818,
        Y => S819
    );
NAND_359: ENTITY WORK.NAND
    PORT MAP (
        A => S436,
        B => S819,
        Y => S820
    );
NAND_360: ENTITY WORK.NAND
    PORT MAP (
        A => S816,
        B => S820,
        Y => S821
    );
NAND_361: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_215,
        B => S422,
        Y => S822
    );
NAND_362: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_151,
        B => S423,
        Y => S823
    );
NAND_363: ENTITY WORK.NAND
    PORT MAP (
        A => S822,
        B => S823,
        Y => S824
    );
NAND_364: ENTITY WORK.NAND
    PORT MAP (
        A => S435,
        B => S824,
        Y => S825
    );
NOR_147: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_135,
        B => S422,
        Y => S826
    );
NAND_365: ENTITY WORK.NAND
    PORT MAP (
        A => S7728,
        B => S422,
        Y => S827
    );
NAND_366: ENTITY WORK.NAND
    PORT MAP (
        A => S436,
        B => S827,
        Y => S828
    );
NOR_148: ENTITY WORK.NOR
    PORT MAP (
        A => S826,
        B => S828,
        Y => S829
    );
NOR_149: ENTITY WORK.NOR
    PORT MAP (
        A => S442,
        B => S821,
        Y => S830
    );
NOR_150: ENTITY WORK.NOR
    PORT MAP (
        A => S441,
        B => S829,
        Y => S831
    );
NAND_367: ENTITY WORK.NAND
    PORT MAP (
        A => S825,
        B => S831,
        Y => S832
    );
NAND_368: ENTITY WORK.NAND
    PORT MAP (
        A => S428,
        B => S832,
        Y => S833
    );
NOR_151: ENTITY WORK.NOR
    PORT MAP (
        A => S830,
        B => S833,
        Y => S834
    );
NAND_369: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_55,
        B => S435,
        Y => S835
    );
NAND_370: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_39,
        B => S436,
        Y => S836
    );
NAND_371: ENTITY WORK.NAND
    PORT MAP (
        A => S835,
        B => S836,
        Y => S837
    );
NAND_372: ENTITY WORK.NAND
    PORT MAP (
        A => S441,
        B => S837,
        Y => S838
    );
NAND_373: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_7,
        B => S436,
        Y => S839
    );
NAND_374: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_23,
        B => S435,
        Y => S840
    );
NAND_375: ENTITY WORK.NAND
    PORT MAP (
        A => S839,
        B => S840,
        Y => S841
    );
NAND_376: ENTITY WORK.NAND
    PORT MAP (
        A => S442,
        B => S841,
        Y => S842
    );
NAND_377: ENTITY WORK.NAND
    PORT MAP (
        A => S838,
        B => S842,
        Y => S843
    );
NAND_378: ENTITY WORK.NAND
    PORT MAP (
        A => S429,
        B => S843,
        Y => S844
    );
NAND_379: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_119,
        B => S435,
        Y => S845
    );
NAND_380: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_103,
        B => S436,
        Y => S846
    );
NAND_381: ENTITY WORK.NAND
    PORT MAP (
        A => S845,
        B => S846,
        Y => S847
    );
NAND_382: ENTITY WORK.NAND
    PORT MAP (
        A => S441,
        B => S847,
        Y => S848
    );
NAND_383: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_87,
        B => S435,
        Y => S849
    );
NAND_384: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_71,
        B => S436,
        Y => S850
    );
NAND_385: ENTITY WORK.NAND
    PORT MAP (
        A => S849,
        B => S850,
        Y => S851
    );
NAND_386: ENTITY WORK.NAND
    PORT MAP (
        A => S442,
        B => S851,
        Y => S852
    );
NAND_387: ENTITY WORK.NAND
    PORT MAP (
        A => S848,
        B => S852,
        Y => S853
    );
NAND_388: ENTITY WORK.NAND
    PORT MAP (
        A => S479,
        B => S853,
        Y => S854
    );
NAND_389: ENTITY WORK.NAND
    PORT MAP (
        A => S844,
        B => S854,
        Y => S855
    );
NOR_152: ENTITY WORK.NOR
    PORT MAP (
        A => S834,
        B => S855,
        Y => S856
    );
NAND_390: ENTITY WORK.NAND
    PORT MAP (
        A => S446,
        B => S856,
        Y => S857
    );
NAND_391: ENTITY WORK.NAND
    PORT MAP (
        A => S812,
        B => S857,
        Y => S858
    );
NOT_137: ENTITY WORK.NOT
    PORT MAP (
        A => S858,
        Y => datapath_addsubunit_in1_7
    );
NAND_392: ENTITY WORK.NAND
    PORT MAP (
        A => S496,
        B => datapath_addsubunit_in1_7,
        Y => S859
    );
NAND_393: ENTITY WORK.NAND
    PORT MAP (
        A => S372,
        B => S859,
        Y => S860
    );
NOT_138: ENTITY WORK.NOT
    PORT MAP (
        A => S860,
        Y => S861
    );
NOR_153: ENTITY WORK.NOR
    PORT MAP (
        A => S7936,
        B => S861,
        Y => S862
    );
NOR_154: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_muxmem_in2_7,
        B => S860,
        Y => S863
    );
NAND_394: ENTITY WORK.NAND
    PORT MAP (
        A => S7876,
        B => S445,
        Y => S864
    );
NAND_395: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_182,
        B => S423,
        Y => S865
    );
NAND_396: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_246,
        B => S422,
        Y => S866
    );
NAND_397: ENTITY WORK.NAND
    PORT MAP (
        A => S865,
        B => S866,
        Y => S867
    );
NAND_398: ENTITY WORK.NAND
    PORT MAP (
        A => S435,
        B => S867,
        Y => S868
    );
NOR_155: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_166,
        B => S422,
        Y => S869
    );
NOR_156: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_230,
        B => S423,
        Y => S870
    );
NOR_157: ENTITY WORK.NOR
    PORT MAP (
        A => S869,
        B => S870,
        Y => S871
    );
NAND_399: ENTITY WORK.NAND
    PORT MAP (
        A => S436,
        B => S871,
        Y => S872
    );
NAND_400: ENTITY WORK.NAND
    PORT MAP (
        A => S868,
        B => S872,
        Y => S873
    );
NAND_401: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_214,
        B => S422,
        Y => S874
    );
NAND_402: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_150,
        B => S423,
        Y => S875
    );
NAND_403: ENTITY WORK.NAND
    PORT MAP (
        A => S874,
        B => S875,
        Y => S876
    );
NAND_404: ENTITY WORK.NAND
    PORT MAP (
        A => S435,
        B => S876,
        Y => S877
    );
NOR_158: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_134,
        B => S422,
        Y => S878
    );
NAND_405: ENTITY WORK.NAND
    PORT MAP (
        A => S7717,
        B => S422,
        Y => S879
    );
NAND_406: ENTITY WORK.NAND
    PORT MAP (
        A => S436,
        B => S879,
        Y => S880
    );
NOR_159: ENTITY WORK.NOR
    PORT MAP (
        A => S878,
        B => S880,
        Y => S881
    );
NOR_160: ENTITY WORK.NOR
    PORT MAP (
        A => S442,
        B => S873,
        Y => S882
    );
NOR_161: ENTITY WORK.NOR
    PORT MAP (
        A => S441,
        B => S881,
        Y => S883
    );
NAND_407: ENTITY WORK.NAND
    PORT MAP (
        A => S877,
        B => S883,
        Y => S884
    );
NAND_408: ENTITY WORK.NAND
    PORT MAP (
        A => S428,
        B => S884,
        Y => S885
    );
NOR_162: ENTITY WORK.NOR
    PORT MAP (
        A => S882,
        B => S885,
        Y => S886
    );
NAND_409: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_54,
        B => S435,
        Y => S887
    );
NAND_410: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_38,
        B => S436,
        Y => S888
    );
NAND_411: ENTITY WORK.NAND
    PORT MAP (
        A => S887,
        B => S888,
        Y => S889
    );
NAND_412: ENTITY WORK.NAND
    PORT MAP (
        A => S441,
        B => S889,
        Y => S890
    );
NAND_413: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_6,
        B => S436,
        Y => S891
    );
NAND_414: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_22,
        B => S435,
        Y => S892
    );
NAND_415: ENTITY WORK.NAND
    PORT MAP (
        A => S891,
        B => S892,
        Y => S893
    );
NAND_416: ENTITY WORK.NAND
    PORT MAP (
        A => S442,
        B => S893,
        Y => S894
    );
NAND_417: ENTITY WORK.NAND
    PORT MAP (
        A => S890,
        B => S894,
        Y => S895
    );
NAND_418: ENTITY WORK.NAND
    PORT MAP (
        A => S429,
        B => S895,
        Y => S896
    );
NAND_419: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_118,
        B => S435,
        Y => S897
    );
NAND_420: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_102,
        B => S436,
        Y => S898
    );
NAND_421: ENTITY WORK.NAND
    PORT MAP (
        A => S897,
        B => S898,
        Y => S899
    );
NAND_422: ENTITY WORK.NAND
    PORT MAP (
        A => S441,
        B => S899,
        Y => S900
    );
NAND_423: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_86,
        B => S435,
        Y => S901
    );
NAND_424: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_70,
        B => S436,
        Y => S902
    );
NAND_425: ENTITY WORK.NAND
    PORT MAP (
        A => S901,
        B => S902,
        Y => S903
    );
NAND_426: ENTITY WORK.NAND
    PORT MAP (
        A => S442,
        B => S903,
        Y => S904
    );
NAND_427: ENTITY WORK.NAND
    PORT MAP (
        A => S900,
        B => S904,
        Y => S905
    );
NAND_428: ENTITY WORK.NAND
    PORT MAP (
        A => S479,
        B => S905,
        Y => S906
    );
NAND_429: ENTITY WORK.NAND
    PORT MAP (
        A => S446,
        B => S906,
        Y => S907
    );
NOR_163: ENTITY WORK.NOR
    PORT MAP (
        A => S886,
        B => S907,
        Y => S908
    );
NAND_430: ENTITY WORK.NAND
    PORT MAP (
        A => S896,
        B => S908,
        Y => S909
    );
NAND_431: ENTITY WORK.NAND
    PORT MAP (
        A => S864,
        B => S909,
        Y => S910
    );
NOT_139: ENTITY WORK.NOT
    PORT MAP (
        A => S910,
        Y => datapath_addsubunit_in1_6
    );
NAND_432: ENTITY WORK.NAND
    PORT MAP (
        A => S496,
        B => datapath_addsubunit_in1_6,
        Y => S911
    );
NAND_433: ENTITY WORK.NAND
    PORT MAP (
        A => S372,
        B => S911,
        Y => S912
    );
NAND_434: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_6,
        B => S912,
        Y => S913
    );
NOT_140: ENTITY WORK.NOT
    PORT MAP (
        A => S913,
        Y => S914
    );
NOR_164: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_muxmem_in2_6,
        B => S912,
        Y => S915
    );
NOR_165: ENTITY WORK.NOR
    PORT MAP (
        A => S914,
        B => S915,
        Y => S916
    );
NAND_435: ENTITY WORK.NAND
    PORT MAP (
        A => S7869,
        B => S445,
        Y => S917
    );
NAND_436: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_181,
        B => S423,
        Y => S918
    );
NAND_437: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_245,
        B => S422,
        Y => S919
    );
NAND_438: ENTITY WORK.NAND
    PORT MAP (
        A => S918,
        B => S919,
        Y => S920
    );
NAND_439: ENTITY WORK.NAND
    PORT MAP (
        A => S435,
        B => S920,
        Y => S921
    );
NOR_166: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_165,
        B => S422,
        Y => S922
    );
NOR_167: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_229,
        B => S423,
        Y => S923
    );
NOR_168: ENTITY WORK.NOR
    PORT MAP (
        A => S922,
        B => S923,
        Y => S924
    );
NAND_440: ENTITY WORK.NAND
    PORT MAP (
        A => S436,
        B => S924,
        Y => S925
    );
NAND_441: ENTITY WORK.NAND
    PORT MAP (
        A => S921,
        B => S925,
        Y => S926
    );
NAND_442: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_213,
        B => S422,
        Y => S927
    );
NAND_443: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_149,
        B => S423,
        Y => S928
    );
NAND_444: ENTITY WORK.NAND
    PORT MAP (
        A => S927,
        B => S928,
        Y => S929
    );
NAND_445: ENTITY WORK.NAND
    PORT MAP (
        A => S435,
        B => S929,
        Y => S930
    );
NOR_169: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_133,
        B => S422,
        Y => S931
    );
NAND_446: ENTITY WORK.NAND
    PORT MAP (
        A => S7706,
        B => S422,
        Y => S932
    );
NAND_447: ENTITY WORK.NAND
    PORT MAP (
        A => S436,
        B => S932,
        Y => S933
    );
NOR_170: ENTITY WORK.NOR
    PORT MAP (
        A => S931,
        B => S933,
        Y => S934
    );
NOR_171: ENTITY WORK.NOR
    PORT MAP (
        A => S442,
        B => S926,
        Y => S935
    );
NOR_172: ENTITY WORK.NOR
    PORT MAP (
        A => S441,
        B => S934,
        Y => S936
    );
NAND_448: ENTITY WORK.NAND
    PORT MAP (
        A => S930,
        B => S936,
        Y => S937
    );
NAND_449: ENTITY WORK.NAND
    PORT MAP (
        A => S428,
        B => S937,
        Y => S938
    );
NOR_173: ENTITY WORK.NOR
    PORT MAP (
        A => S935,
        B => S938,
        Y => S939
    );
NAND_450: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_53,
        B => S435,
        Y => S940
    );
NAND_451: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_37,
        B => S436,
        Y => S941
    );
NAND_452: ENTITY WORK.NAND
    PORT MAP (
        A => S940,
        B => S941,
        Y => S942
    );
NAND_453: ENTITY WORK.NAND
    PORT MAP (
        A => S441,
        B => S942,
        Y => S943
    );
NAND_454: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_5,
        B => S436,
        Y => S944
    );
NAND_455: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_21,
        B => S435,
        Y => S945
    );
NAND_456: ENTITY WORK.NAND
    PORT MAP (
        A => S944,
        B => S945,
        Y => S946
    );
NAND_457: ENTITY WORK.NAND
    PORT MAP (
        A => S442,
        B => S946,
        Y => S947
    );
NAND_458: ENTITY WORK.NAND
    PORT MAP (
        A => S943,
        B => S947,
        Y => S948
    );
NAND_459: ENTITY WORK.NAND
    PORT MAP (
        A => S429,
        B => S948,
        Y => S949
    );
NAND_460: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_117,
        B => S435,
        Y => S950
    );
NAND_461: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_101,
        B => S436,
        Y => S951
    );
NAND_462: ENTITY WORK.NAND
    PORT MAP (
        A => S950,
        B => S951,
        Y => S952
    );
NAND_463: ENTITY WORK.NAND
    PORT MAP (
        A => S441,
        B => S952,
        Y => S953
    );
NAND_464: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_85,
        B => S435,
        Y => S954
    );
NAND_465: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_69,
        B => S436,
        Y => S955
    );
NAND_466: ENTITY WORK.NAND
    PORT MAP (
        A => S954,
        B => S955,
        Y => S956
    );
NAND_467: ENTITY WORK.NAND
    PORT MAP (
        A => S442,
        B => S956,
        Y => S957
    );
NAND_468: ENTITY WORK.NAND
    PORT MAP (
        A => S953,
        B => S957,
        Y => S958
    );
NAND_469: ENTITY WORK.NAND
    PORT MAP (
        A => S479,
        B => S958,
        Y => S959
    );
NAND_470: ENTITY WORK.NAND
    PORT MAP (
        A => S949,
        B => S959,
        Y => S960
    );
NOR_174: ENTITY WORK.NOR
    PORT MAP (
        A => S939,
        B => S960,
        Y => S961
    );
NAND_471: ENTITY WORK.NAND
    PORT MAP (
        A => S446,
        B => S961,
        Y => S962
    );
NAND_472: ENTITY WORK.NAND
    PORT MAP (
        A => S917,
        B => S962,
        Y => S963
    );
NOT_141: ENTITY WORK.NOT
    PORT MAP (
        A => S963,
        Y => datapath_addsubunit_in1_5
    );
NAND_473: ENTITY WORK.NAND
    PORT MAP (
        A => S496,
        B => datapath_addsubunit_in1_5,
        Y => S964
    );
NAND_474: ENTITY WORK.NAND
    PORT MAP (
        A => S372,
        B => S964,
        Y => S965
    );
NOT_142: ENTITY WORK.NOT
    PORT MAP (
        A => S965,
        Y => S966
    );
NOR_175: ENTITY WORK.NOR
    PORT MAP (
        A => S7920,
        B => S966,
        Y => S967
    );
NOR_176: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_muxmem_in2_5,
        B => S965,
        Y => S968
    );
NAND_475: ENTITY WORK.NAND
    PORT MAP (
        A => controller_fib_4,
        B => S370,
        Y => S969
    );
NAND_476: ENTITY WORK.NAND
    PORT MAP (
        A => S7861,
        B => S445,
        Y => S970
    );
NOR_177: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_164,
        B => S422,
        Y => S971
    );
NOR_178: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_228,
        B => S423,
        Y => S972
    );
NOR_179: ENTITY WORK.NOR
    PORT MAP (
        A => S971,
        B => S972,
        Y => S973
    );
NAND_477: ENTITY WORK.NAND
    PORT MAP (
        A => S436,
        B => S973,
        Y => S974
    );
NOR_180: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_244,
        B => S423,
        Y => S975
    );
NAND_478: ENTITY WORK.NAND
    PORT MAP (
        A => S7596,
        B => S423,
        Y => S976
    );
NAND_479: ENTITY WORK.NAND
    PORT MAP (
        A => S435,
        B => S976,
        Y => S977
    );
NOR_181: ENTITY WORK.NOR
    PORT MAP (
        A => S975,
        B => S977,
        Y => S978
    );
NAND_480: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_196,
        B => S436,
        Y => S979
    );
NAND_481: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_212,
        B => S435,
        Y => S980
    );
NAND_482: ENTITY WORK.NAND
    PORT MAP (
        A => S979,
        B => S980,
        Y => S981
    );
NAND_483: ENTITY WORK.NAND
    PORT MAP (
        A => S422,
        B => S981,
        Y => S982
    );
NAND_484: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_132,
        B => S436,
        Y => S983
    );
NAND_485: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_148,
        B => S435,
        Y => S984
    );
NAND_486: ENTITY WORK.NAND
    PORT MAP (
        A => S983,
        B => S984,
        Y => S985
    );
NAND_487: ENTITY WORK.NAND
    PORT MAP (
        A => S423,
        B => S985,
        Y => S986
    );
NAND_488: ENTITY WORK.NAND
    PORT MAP (
        A => S982,
        B => S986,
        Y => S987
    );
NOR_182: ENTITY WORK.NOR
    PORT MAP (
        A => S441,
        B => S987,
        Y => S988
    );
NOR_183: ENTITY WORK.NOR
    PORT MAP (
        A => S442,
        B => S978,
        Y => S989
    );
NAND_489: ENTITY WORK.NAND
    PORT MAP (
        A => S974,
        B => S989,
        Y => S990
    );
NAND_490: ENTITY WORK.NAND
    PORT MAP (
        A => S428,
        B => S990,
        Y => S991
    );
NOR_184: ENTITY WORK.NOR
    PORT MAP (
        A => S988,
        B => S991,
        Y => S992
    );
NAND_491: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_116,
        B => S435,
        Y => S993
    );
NAND_492: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_100,
        B => S436,
        Y => S994
    );
NAND_493: ENTITY WORK.NAND
    PORT MAP (
        A => S993,
        B => S994,
        Y => S995
    );
NAND_494: ENTITY WORK.NAND
    PORT MAP (
        A => S441,
        B => S995,
        Y => S996
    );
NAND_495: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_84,
        B => S435,
        Y => S997
    );
NAND_496: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_68,
        B => S436,
        Y => S998
    );
NAND_497: ENTITY WORK.NAND
    PORT MAP (
        A => S997,
        B => S998,
        Y => S999
    );
NAND_498: ENTITY WORK.NAND
    PORT MAP (
        A => S442,
        B => S999,
        Y => S1000
    );
NAND_499: ENTITY WORK.NAND
    PORT MAP (
        A => S996,
        B => S1000,
        Y => S1001
    );
NAND_500: ENTITY WORK.NAND
    PORT MAP (
        A => S479,
        B => S1001,
        Y => S1002
    );
NOR_185: ENTITY WORK.NOR
    PORT MAP (
        A => S436,
        B => S442,
        Y => S1003
    );
NAND_501: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_52,
        B => S1003,
        Y => S1004
    );
NOR_186: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_20,
        B => S436,
        Y => S1005
    );
NOR_187: ENTITY WORK.NOR
    PORT MAP (
        A => S441,
        B => S1005,
        Y => S1006
    );
NAND_502: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_36,
        B => S436,
        Y => S1007
    );
NAND_503: ENTITY WORK.NAND
    PORT MAP (
        A => S1004,
        B => S1007,
        Y => S1008
    );
NOR_188: ENTITY WORK.NOR
    PORT MAP (
        A => S1006,
        B => S1008,
        Y => S1009
    );
NOR_189: ENTITY WORK.NOR
    PORT MAP (
        A => S430,
        B => S1009,
        Y => S1010
    );
NOR_190: ENTITY WORK.NOR
    PORT MAP (
        A => S992,
        B => S1010,
        Y => S1011
    );
NAND_504: ENTITY WORK.NAND
    PORT MAP (
        A => S1002,
        B => S1011,
        Y => S1012
    );
NAND_505: ENTITY WORK.NAND
    PORT MAP (
        A => S970,
        B => S1012,
        Y => S1013
    );
NOT_143: ENTITY WORK.NOT
    PORT MAP (
        A => S1013,
        Y => datapath_addsubunit_in1_4
    );
NAND_506: ENTITY WORK.NAND
    PORT MAP (
        A => S496,
        B => datapath_addsubunit_in1_4,
        Y => S1014
    );
NAND_507: ENTITY WORK.NAND
    PORT MAP (
        A => S969,
        B => S1014,
        Y => S1015
    );
NAND_508: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_4,
        B => S1015,
        Y => S1016
    );
NOT_144: ENTITY WORK.NOT
    PORT MAP (
        A => S1016,
        Y => S1017
    );
NOR_191: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_muxmem_in2_4,
        B => S1015,
        Y => S1018
    );
NOR_192: ENTITY WORK.NOR
    PORT MAP (
        A => S1017,
        B => S1018,
        Y => S1019
    );
NAND_509: ENTITY WORK.NAND
    PORT MAP (
        A => controller_fib_3,
        B => S370,
        Y => S1020
    );
NAND_510: ENTITY WORK.NAND
    PORT MAP (
        A => S7853,
        B => S445,
        Y => S1021
    );
NOR_193: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_163,
        B => S422,
        Y => S1022
    );
NOR_194: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_227,
        B => S423,
        Y => S1023
    );
NOR_195: ENTITY WORK.NOR
    PORT MAP (
        A => S1022,
        B => S1023,
        Y => S1024
    );
NAND_511: ENTITY WORK.NAND
    PORT MAP (
        A => S436,
        B => S1024,
        Y => S1025
    );
NOR_196: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_243,
        B => S423,
        Y => S1026
    );
NAND_512: ENTITY WORK.NAND
    PORT MAP (
        A => S7585,
        B => S423,
        Y => S1027
    );
NAND_513: ENTITY WORK.NAND
    PORT MAP (
        A => S435,
        B => S1027,
        Y => S1028
    );
NOR_197: ENTITY WORK.NOR
    PORT MAP (
        A => S1026,
        B => S1028,
        Y => S1029
    );
NAND_514: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_195,
        B => S436,
        Y => S1030
    );
NAND_515: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_211,
        B => S435,
        Y => S1031
    );
NAND_516: ENTITY WORK.NAND
    PORT MAP (
        A => S1030,
        B => S1031,
        Y => S1032
    );
NAND_517: ENTITY WORK.NAND
    PORT MAP (
        A => S422,
        B => S1032,
        Y => S1033
    );
NAND_518: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_131,
        B => S436,
        Y => S1034
    );
NAND_519: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_147,
        B => S435,
        Y => S1035
    );
NAND_520: ENTITY WORK.NAND
    PORT MAP (
        A => S1034,
        B => S1035,
        Y => S1036
    );
NAND_521: ENTITY WORK.NAND
    PORT MAP (
        A => S423,
        B => S1036,
        Y => S1037
    );
NAND_522: ENTITY WORK.NAND
    PORT MAP (
        A => S1033,
        B => S1037,
        Y => S1038
    );
NOR_198: ENTITY WORK.NOR
    PORT MAP (
        A => S441,
        B => S1038,
        Y => S1039
    );
NOR_199: ENTITY WORK.NOR
    PORT MAP (
        A => S442,
        B => S1029,
        Y => S1040
    );
NAND_523: ENTITY WORK.NAND
    PORT MAP (
        A => S1025,
        B => S1040,
        Y => S1041
    );
NAND_524: ENTITY WORK.NAND
    PORT MAP (
        A => S428,
        B => S1041,
        Y => S1042
    );
NOR_200: ENTITY WORK.NOR
    PORT MAP (
        A => S1039,
        B => S1042,
        Y => S1043
    );
NAND_525: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_83,
        B => S442,
        Y => S1044
    );
NAND_526: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_115,
        B => S441,
        Y => S1045
    );
NAND_527: ENTITY WORK.NAND
    PORT MAP (
        A => S1044,
        B => S1045,
        Y => S1046
    );
NAND_528: ENTITY WORK.NAND
    PORT MAP (
        A => S435,
        B => S1046,
        Y => S1047
    );
NAND_529: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_99,
        B => S441,
        Y => S1048
    );
NAND_530: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_67,
        B => S442,
        Y => S1049
    );
NAND_531: ENTITY WORK.NAND
    PORT MAP (
        A => S1048,
        B => S1049,
        Y => S1050
    );
NAND_532: ENTITY WORK.NAND
    PORT MAP (
        A => S436,
        B => S1050,
        Y => S1051
    );
NAND_533: ENTITY WORK.NAND
    PORT MAP (
        A => S1047,
        B => S1051,
        Y => S1052
    );
NAND_534: ENTITY WORK.NAND
    PORT MAP (
        A => S479,
        B => S1052,
        Y => S1053
    );
NAND_535: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_51,
        B => S1003,
        Y => S1054
    );
NAND_536: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_35,
        B => S436,
        Y => S1055
    );
NOT_145: ENTITY WORK.NOT
    PORT MAP (
        A => S1055,
        Y => S1056
    );
NOR_201: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_19,
        B => S436,
        Y => S1057
    );
NOR_202: ENTITY WORK.NOR
    PORT MAP (
        A => S441,
        B => S1057,
        Y => S1058
    );
NOR_203: ENTITY WORK.NOR
    PORT MAP (
        A => S1056,
        B => S1058,
        Y => S1059
    );
NAND_537: ENTITY WORK.NAND
    PORT MAP (
        A => S1054,
        B => S1059,
        Y => S1060
    );
NAND_538: ENTITY WORK.NAND
    PORT MAP (
        A => S429,
        B => S1060,
        Y => S1061
    );
NOT_146: ENTITY WORK.NOT
    PORT MAP (
        A => S1061,
        Y => S1062
    );
NOR_204: ENTITY WORK.NOR
    PORT MAP (
        A => S1043,
        B => S1062,
        Y => S1063
    );
NAND_539: ENTITY WORK.NAND
    PORT MAP (
        A => S1053,
        B => S1063,
        Y => S1064
    );
NAND_540: ENTITY WORK.NAND
    PORT MAP (
        A => S1021,
        B => S1064,
        Y => S1065
    );
NOT_147: ENTITY WORK.NOT
    PORT MAP (
        A => S1065,
        Y => datapath_addsubunit_in1_3
    );
NAND_541: ENTITY WORK.NAND
    PORT MAP (
        A => S496,
        B => datapath_addsubunit_in1_3,
        Y => S1066
    );
NAND_542: ENTITY WORK.NAND
    PORT MAP (
        A => S1020,
        B => S1066,
        Y => S1067
    );
NAND_543: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_3,
        B => S1067,
        Y => S1068
    );
NOT_148: ENTITY WORK.NOT
    PORT MAP (
        A => S1068,
        Y => S1069
    );
NOR_205: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_muxmem_in2_3,
        B => S1067,
        Y => S1070
    );
NAND_544: ENTITY WORK.NAND
    PORT MAP (
        A => controller_fib_2,
        B => S370,
        Y => S1071
    );
NAND_545: ENTITY WORK.NAND
    PORT MAP (
        A => S7846,
        B => S445,
        Y => S1072
    );
NAND_546: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_178,
        B => S423,
        Y => S1073
    );
NAND_547: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_242,
        B => S422,
        Y => S1074
    );
NAND_548: ENTITY WORK.NAND
    PORT MAP (
        A => S1073,
        B => S1074,
        Y => S1075
    );
NAND_549: ENTITY WORK.NAND
    PORT MAP (
        A => S435,
        B => S1075,
        Y => S1076
    );
NOR_206: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_162,
        B => S422,
        Y => S1077
    );
NOR_207: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_226,
        B => S423,
        Y => S1078
    );
NOR_208: ENTITY WORK.NOR
    PORT MAP (
        A => S1077,
        B => S1078,
        Y => S1079
    );
NAND_550: ENTITY WORK.NAND
    PORT MAP (
        A => S436,
        B => S1079,
        Y => S1080
    );
NAND_551: ENTITY WORK.NAND
    PORT MAP (
        A => S1076,
        B => S1080,
        Y => S1081
    );
NAND_552: ENTITY WORK.NAND
    PORT MAP (
        A => S441,
        B => S1081,
        Y => S1082
    );
NAND_553: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_210,
        B => S422,
        Y => S1083
    );
NAND_554: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_146,
        B => S423,
        Y => S1084
    );
NAND_555: ENTITY WORK.NAND
    PORT MAP (
        A => S1083,
        B => S1084,
        Y => S1085
    );
NAND_556: ENTITY WORK.NAND
    PORT MAP (
        A => S435,
        B => S1085,
        Y => S1086
    );
NOR_209: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_130,
        B => S422,
        Y => S1087
    );
NOR_210: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_194,
        B => S423,
        Y => S1088
    );
NOR_211: ENTITY WORK.NOR
    PORT MAP (
        A => S1087,
        B => S1088,
        Y => S1089
    );
NAND_557: ENTITY WORK.NAND
    PORT MAP (
        A => S436,
        B => S1089,
        Y => S1090
    );
NAND_558: ENTITY WORK.NAND
    PORT MAP (
        A => S1086,
        B => S1090,
        Y => S1091
    );
NAND_559: ENTITY WORK.NAND
    PORT MAP (
        A => S442,
        B => S1091,
        Y => S1092
    );
NAND_560: ENTITY WORK.NAND
    PORT MAP (
        A => S1082,
        B => S1092,
        Y => S1093
    );
NAND_561: ENTITY WORK.NAND
    PORT MAP (
        A => S428,
        B => S1093,
        Y => S1094
    );
NAND_562: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_114,
        B => S435,
        Y => S1095
    );
NAND_563: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_98,
        B => S436,
        Y => S1096
    );
NAND_564: ENTITY WORK.NAND
    PORT MAP (
        A => S1095,
        B => S1096,
        Y => S1097
    );
NAND_565: ENTITY WORK.NAND
    PORT MAP (
        A => S441,
        B => S1097,
        Y => S1098
    );
NAND_566: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_82,
        B => S435,
        Y => S1099
    );
NAND_567: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_66,
        B => S436,
        Y => S1100
    );
NAND_568: ENTITY WORK.NAND
    PORT MAP (
        A => S1099,
        B => S1100,
        Y => S1101
    );
NAND_569: ENTITY WORK.NAND
    PORT MAP (
        A => S442,
        B => S1101,
        Y => S1102
    );
NAND_570: ENTITY WORK.NAND
    PORT MAP (
        A => S1098,
        B => S1102,
        Y => S1103
    );
NAND_571: ENTITY WORK.NAND
    PORT MAP (
        A => S479,
        B => S1103,
        Y => S1104
    );
NOT_149: ENTITY WORK.NOT
    PORT MAP (
        A => S1104,
        Y => S1105
    );
NOR_212: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_18,
        B => S441,
        Y => S1106
    );
NOR_213: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_50,
        B => S442,
        Y => S1107
    );
NOR_214: ENTITY WORK.NOR
    PORT MAP (
        A => S1106,
        B => S1107,
        Y => S1108
    );
NOR_215: ENTITY WORK.NOR
    PORT MAP (
        A => S436,
        B => S1108,
        Y => S1109
    );
NOR_216: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_34,
        B => S442,
        Y => S1110
    );
NAND_572: ENTITY WORK.NAND
    PORT MAP (
        A => S436,
        B => S1110,
        Y => S1111
    );
NAND_573: ENTITY WORK.NAND
    PORT MAP (
        A => S429,
        B => S1111,
        Y => S1112
    );
NOR_217: ENTITY WORK.NOR
    PORT MAP (
        A => S1109,
        B => S1112,
        Y => S1113
    );
NOR_218: ENTITY WORK.NOR
    PORT MAP (
        A => S1105,
        B => S1113,
        Y => S1114
    );
NAND_574: ENTITY WORK.NAND
    PORT MAP (
        A => S1094,
        B => S1114,
        Y => S1115
    );
NAND_575: ENTITY WORK.NAND
    PORT MAP (
        A => S1072,
        B => S1115,
        Y => S1116
    );
NOT_150: ENTITY WORK.NOT
    PORT MAP (
        A => S1116,
        Y => datapath_addsubunit_in1_2
    );
NAND_576: ENTITY WORK.NAND
    PORT MAP (
        A => S496,
        B => datapath_addsubunit_in1_2,
        Y => S1117
    );
NAND_577: ENTITY WORK.NAND
    PORT MAP (
        A => S1071,
        B => S1117,
        Y => S1118
    );
NAND_578: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_2,
        B => S1118,
        Y => S1119
    );
NOT_151: ENTITY WORK.NOT
    PORT MAP (
        A => S1119,
        Y => S1120
    );
NAND_579: ENTITY WORK.NAND
    PORT MAP (
        A => controller_fib_1,
        B => S370,
        Y => S1121
    );
NAND_580: ENTITY WORK.NAND
    PORT MAP (
        A => S7838,
        B => S445,
        Y => S1122
    );
NAND_581: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_177,
        B => S423,
        Y => S1123
    );
NAND_582: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_241,
        B => S422,
        Y => S1124
    );
NAND_583: ENTITY WORK.NAND
    PORT MAP (
        A => S1123,
        B => S1124,
        Y => S1125
    );
NAND_584: ENTITY WORK.NAND
    PORT MAP (
        A => S435,
        B => S1125,
        Y => S1126
    );
NOR_219: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_161,
        B => S422,
        Y => S1127
    );
NOR_220: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_225,
        B => S423,
        Y => S1128
    );
NOR_221: ENTITY WORK.NOR
    PORT MAP (
        A => S1127,
        B => S1128,
        Y => S1129
    );
NAND_585: ENTITY WORK.NAND
    PORT MAP (
        A => S436,
        B => S1129,
        Y => S1130
    );
NAND_586: ENTITY WORK.NAND
    PORT MAP (
        A => S1126,
        B => S1130,
        Y => S1131
    );
NAND_587: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_209,
        B => S422,
        Y => S1132
    );
NAND_588: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_145,
        B => S423,
        Y => S1133
    );
NAND_589: ENTITY WORK.NAND
    PORT MAP (
        A => S1132,
        B => S1133,
        Y => S1134
    );
NAND_590: ENTITY WORK.NAND
    PORT MAP (
        A => S435,
        B => S1134,
        Y => S1135
    );
NOR_222: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_129,
        B => S422,
        Y => S1136
    );
NAND_591: ENTITY WORK.NAND
    PORT MAP (
        A => S7684,
        B => S422,
        Y => S1137
    );
NAND_592: ENTITY WORK.NAND
    PORT MAP (
        A => S436,
        B => S1137,
        Y => S1138
    );
NOR_223: ENTITY WORK.NOR
    PORT MAP (
        A => S1136,
        B => S1138,
        Y => S1139
    );
NOR_224: ENTITY WORK.NOR
    PORT MAP (
        A => S442,
        B => S1131,
        Y => S1140
    );
NOR_225: ENTITY WORK.NOR
    PORT MAP (
        A => S441,
        B => S1139,
        Y => S1141
    );
NAND_593: ENTITY WORK.NAND
    PORT MAP (
        A => S1135,
        B => S1141,
        Y => S1142
    );
NAND_594: ENTITY WORK.NAND
    PORT MAP (
        A => S428,
        B => S1142,
        Y => S1143
    );
NOR_226: ENTITY WORK.NOR
    PORT MAP (
        A => S1140,
        B => S1143,
        Y => S1144
    );
NAND_595: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_17,
        B => S442,
        Y => S1145
    );
NAND_596: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_49,
        B => S441,
        Y => S1146
    );
NAND_597: ENTITY WORK.NAND
    PORT MAP (
        A => S1145,
        B => S1146,
        Y => S1147
    );
NAND_598: ENTITY WORK.NAND
    PORT MAP (
        A => S435,
        B => S1147,
        Y => S1148
    );
NAND_599: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_1,
        B => S442,
        Y => S1149
    );
NAND_600: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_33,
        B => S441,
        Y => S1150
    );
NAND_601: ENTITY WORK.NAND
    PORT MAP (
        A => S1149,
        B => S1150,
        Y => S1151
    );
NAND_602: ENTITY WORK.NAND
    PORT MAP (
        A => S436,
        B => S1151,
        Y => S1152
    );
NAND_603: ENTITY WORK.NAND
    PORT MAP (
        A => S1148,
        B => S1152,
        Y => S1153
    );
NAND_604: ENTITY WORK.NAND
    PORT MAP (
        A => S429,
        B => S1153,
        Y => S1154
    );
NAND_605: ENTITY WORK.NAND
    PORT MAP (
        A => S7531,
        B => S436,
        Y => S1155
    );
NOR_227: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_113,
        B => S436,
        Y => S1156
    );
NOR_228: ENTITY WORK.NOR
    PORT MAP (
        A => S442,
        B => S1156,
        Y => S1157
    );
NAND_606: ENTITY WORK.NAND
    PORT MAP (
        A => S1155,
        B => S1157,
        Y => S1158
    );
NOR_229: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_65,
        B => S435,
        Y => S1159
    );
NOR_230: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_81,
        B => S436,
        Y => S1160
    );
NOR_231: ENTITY WORK.NOR
    PORT MAP (
        A => S1159,
        B => S1160,
        Y => S1161
    );
NAND_607: ENTITY WORK.NAND
    PORT MAP (
        A => S442,
        B => S1161,
        Y => S1162
    );
NAND_608: ENTITY WORK.NAND
    PORT MAP (
        A => S1158,
        B => S1162,
        Y => S1163
    );
NAND_609: ENTITY WORK.NAND
    PORT MAP (
        A => S479,
        B => S1163,
        Y => S1164
    );
NAND_610: ENTITY WORK.NAND
    PORT MAP (
        A => S1154,
        B => S1164,
        Y => S1165
    );
NOR_232: ENTITY WORK.NOR
    PORT MAP (
        A => S1144,
        B => S1165,
        Y => S1166
    );
NAND_611: ENTITY WORK.NAND
    PORT MAP (
        A => S446,
        B => S1166,
        Y => S1167
    );
NAND_612: ENTITY WORK.NAND
    PORT MAP (
        A => S1122,
        B => S1167,
        Y => S1168
    );
NOT_152: ENTITY WORK.NOT
    PORT MAP (
        A => S1168,
        Y => datapath_addsubunit_in1_1
    );
NAND_613: ENTITY WORK.NAND
    PORT MAP (
        A => S496,
        B => datapath_addsubunit_in1_1,
        Y => S1169
    );
NAND_614: ENTITY WORK.NAND
    PORT MAP (
        A => S1121,
        B => S1169,
        Y => S1170
    );
NAND_615: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_1,
        B => S1170,
        Y => S1171
    );
NOT_153: ENTITY WORK.NOT
    PORT MAP (
        A => S1171,
        Y => S1172
    );
NAND_616: ENTITY WORK.NAND
    PORT MAP (
        A => controller_fib_0,
        B => S370,
        Y => S1173
    );
NAND_617: ENTITY WORK.NAND
    PORT MAP (
        A => S7830,
        B => S445,
        Y => S1174
    );
NAND_618: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_176,
        B => S423,
        Y => S1175
    );
NAND_619: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_240,
        B => S422,
        Y => S1176
    );
NAND_620: ENTITY WORK.NAND
    PORT MAP (
        A => S1175,
        B => S1176,
        Y => S1177
    );
NAND_621: ENTITY WORK.NAND
    PORT MAP (
        A => S435,
        B => S1177,
        Y => S1178
    );
NOR_233: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_160,
        B => S422,
        Y => S1179
    );
NOR_234: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_224,
        B => S423,
        Y => S1180
    );
NOR_235: ENTITY WORK.NOR
    PORT MAP (
        A => S1179,
        B => S1180,
        Y => S1181
    );
NAND_622: ENTITY WORK.NAND
    PORT MAP (
        A => S436,
        B => S1181,
        Y => S1182
    );
NAND_623: ENTITY WORK.NAND
    PORT MAP (
        A => S1178,
        B => S1182,
        Y => S1183
    );
NAND_624: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_208,
        B => S422,
        Y => S1184
    );
NAND_625: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_144,
        B => S423,
        Y => S1185
    );
NAND_626: ENTITY WORK.NAND
    PORT MAP (
        A => S1184,
        B => S1185,
        Y => S1186
    );
NAND_627: ENTITY WORK.NAND
    PORT MAP (
        A => S435,
        B => S1186,
        Y => S1187
    );
NOR_236: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_128,
        B => S422,
        Y => S1188
    );
NAND_628: ENTITY WORK.NAND
    PORT MAP (
        A => S7673,
        B => S422,
        Y => S1189
    );
NAND_629: ENTITY WORK.NAND
    PORT MAP (
        A => S436,
        B => S1189,
        Y => S1190
    );
NOR_237: ENTITY WORK.NOR
    PORT MAP (
        A => S1188,
        B => S1190,
        Y => S1191
    );
NOR_238: ENTITY WORK.NOR
    PORT MAP (
        A => S442,
        B => S1183,
        Y => S1192
    );
NOR_239: ENTITY WORK.NOR
    PORT MAP (
        A => S441,
        B => S1191,
        Y => S1193
    );
NAND_630: ENTITY WORK.NAND
    PORT MAP (
        A => S1187,
        B => S1193,
        Y => S1194
    );
NAND_631: ENTITY WORK.NAND
    PORT MAP (
        A => S428,
        B => S1194,
        Y => S1195
    );
NOR_240: ENTITY WORK.NOR
    PORT MAP (
        A => S1192,
        B => S1195,
        Y => S1196
    );
NAND_632: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_16,
        B => S442,
        Y => S1197
    );
NAND_633: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_48,
        B => S441,
        Y => S1198
    );
NAND_634: ENTITY WORK.NAND
    PORT MAP (
        A => S1197,
        B => S1198,
        Y => S1199
    );
NAND_635: ENTITY WORK.NAND
    PORT MAP (
        A => S435,
        B => S1199,
        Y => S1200
    );
NAND_636: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_0,
        B => S442,
        Y => S1201
    );
NAND_637: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_32,
        B => S441,
        Y => S1202
    );
NAND_638: ENTITY WORK.NAND
    PORT MAP (
        A => S1201,
        B => S1202,
        Y => S1203
    );
NAND_639: ENTITY WORK.NAND
    PORT MAP (
        A => S436,
        B => S1203,
        Y => S1204
    );
NAND_640: ENTITY WORK.NAND
    PORT MAP (
        A => S1200,
        B => S1204,
        Y => S1205
    );
NAND_641: ENTITY WORK.NAND
    PORT MAP (
        A => S429,
        B => S1205,
        Y => S1206
    );
NAND_642: ENTITY WORK.NAND
    PORT MAP (
        A => S7520,
        B => S436,
        Y => S1207
    );
NOR_241: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_112,
        B => S436,
        Y => S1208
    );
NOR_242: ENTITY WORK.NOR
    PORT MAP (
        A => S442,
        B => S1208,
        Y => S1209
    );
NAND_643: ENTITY WORK.NAND
    PORT MAP (
        A => S1207,
        B => S1209,
        Y => S1210
    );
NOR_243: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_64,
        B => S435,
        Y => S1211
    );
NOR_244: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_80,
        B => S436,
        Y => S1212
    );
NOR_245: ENTITY WORK.NOR
    PORT MAP (
        A => S1211,
        B => S1212,
        Y => S1213
    );
NAND_644: ENTITY WORK.NAND
    PORT MAP (
        A => S442,
        B => S1213,
        Y => S1214
    );
NAND_645: ENTITY WORK.NAND
    PORT MAP (
        A => S1210,
        B => S1214,
        Y => S1215
    );
NAND_646: ENTITY WORK.NAND
    PORT MAP (
        A => S479,
        B => S1215,
        Y => S1216
    );
NAND_647: ENTITY WORK.NAND
    PORT MAP (
        A => S1206,
        B => S1216,
        Y => S1217
    );
NOR_246: ENTITY WORK.NOR
    PORT MAP (
        A => S1196,
        B => S1217,
        Y => S1218
    );
NAND_648: ENTITY WORK.NAND
    PORT MAP (
        A => S446,
        B => S1218,
        Y => S1219
    );
NAND_649: ENTITY WORK.NAND
    PORT MAP (
        A => S1174,
        B => S1219,
        Y => S1220
    );
NOT_154: ENTITY WORK.NOT
    PORT MAP (
        A => S1220,
        Y => datapath_addsubunit_in1_0
    );
NAND_650: ENTITY WORK.NAND
    PORT MAP (
        A => S496,
        B => datapath_addsubunit_in1_0,
        Y => S1221
    );
NAND_651: ENTITY WORK.NAND
    PORT MAP (
        A => S1173,
        B => S1221,
        Y => S1222
    );
NAND_652: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_0,
        B => S1222,
        Y => S1223
    );
NOT_155: ENTITY WORK.NOT
    PORT MAP (
        A => S1223,
        Y => S1224
    );
NOR_247: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_muxmem_in2_1,
        B => S1170,
        Y => S1225
    );
NOR_248: ENTITY WORK.NOR
    PORT MAP (
        A => S1172,
        B => S1225,
        Y => S1226
    );
NAND_653: ENTITY WORK.NAND
    PORT MAP (
        A => S1224,
        B => S1226,
        Y => S1227
    );
NOT_156: ENTITY WORK.NOT
    PORT MAP (
        A => S1227,
        Y => S1228
    );
NAND_654: ENTITY WORK.NAND
    PORT MAP (
        A => S1171,
        B => S1227,
        Y => S1229
    );
NOR_249: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_muxmem_in2_2,
        B => S1118,
        Y => S1230
    );
NOR_250: ENTITY WORK.NOR
    PORT MAP (
        A => S1120,
        B => S1230,
        Y => S1231
    );
NAND_655: ENTITY WORK.NAND
    PORT MAP (
        A => S1229,
        B => S1231,
        Y => S1232
    );
NAND_656: ENTITY WORK.NAND
    PORT MAP (
        A => S1119,
        B => S1232,
        Y => S1233
    );
NOR_251: ENTITY WORK.NOR
    PORT MAP (
        A => S1069,
        B => S1233,
        Y => S1234
    );
NOR_252: ENTITY WORK.NOR
    PORT MAP (
        A => S1070,
        B => S1234,
        Y => S1235
    );
NAND_657: ENTITY WORK.NAND
    PORT MAP (
        A => S1019,
        B => S1235,
        Y => S1236
    );
NAND_658: ENTITY WORK.NAND
    PORT MAP (
        A => S1016,
        B => S1236,
        Y => S1237
    );
NOR_253: ENTITY WORK.NOR
    PORT MAP (
        A => S967,
        B => S1237,
        Y => S1238
    );
NOR_254: ENTITY WORK.NOR
    PORT MAP (
        A => S968,
        B => S1238,
        Y => S1239
    );
NAND_659: ENTITY WORK.NAND
    PORT MAP (
        A => S916,
        B => S1239,
        Y => S1240
    );
NAND_660: ENTITY WORK.NAND
    PORT MAP (
        A => S913,
        B => S1240,
        Y => S1241
    );
NOR_255: ENTITY WORK.NOR
    PORT MAP (
        A => S862,
        B => S1241,
        Y => S1242
    );
NOR_256: ENTITY WORK.NOR
    PORT MAP (
        A => S863,
        B => S1242,
        Y => S1243
    );
NAND_661: ENTITY WORK.NAND
    PORT MAP (
        A => S811,
        B => S1243,
        Y => S1244
    );
NAND_662: ENTITY WORK.NAND
    PORT MAP (
        A => S808,
        B => S1244,
        Y => S1245
    );
NOR_257: ENTITY WORK.NOR
    PORT MAP (
        A => S758,
        B => S1245,
        Y => S1246
    );
NOR_258: ENTITY WORK.NOR
    PORT MAP (
        A => S759,
        B => S1246,
        Y => S1247
    );
NAND_663: ENTITY WORK.NAND
    PORT MAP (
        A => S708,
        B => S1247,
        Y => S1248
    );
NAND_664: ENTITY WORK.NAND
    PORT MAP (
        A => S705,
        B => S1248,
        Y => S1249
    );
NOR_259: ENTITY WORK.NOR
    PORT MAP (
        A => S655,
        B => S1249,
        Y => S1250
    );
NOR_260: ENTITY WORK.NOR
    PORT MAP (
        A => S656,
        B => S1250,
        Y => S1251
    );
NAND_665: ENTITY WORK.NAND
    PORT MAP (
        A => S605,
        B => S1251,
        Y => S1252
    );
NAND_666: ENTITY WORK.NAND
    PORT MAP (
        A => S602,
        B => S1252,
        Y => S1253
    );
NOR_261: ENTITY WORK.NOR
    PORT MAP (
        A => S553,
        B => S1253,
        Y => S1254
    );
NOR_262: ENTITY WORK.NOR
    PORT MAP (
        A => S552,
        B => S1254,
        Y => S1255
    );
NAND_667: ENTITY WORK.NAND
    PORT MAP (
        A => S502,
        B => S1255,
        Y => S1256
    );
NAND_668: ENTITY WORK.NAND
    PORT MAP (
        A => S499,
        B => S1256,
        Y => S1257
    );
NOT_157: ENTITY WORK.NOT
    PORT MAP (
        A => S1257,
        Y => S1258
    );
NAND_669: ENTITY WORK.NAND
    PORT MAP (
        A => S7574,
        B => S423,
        Y => S1259
    );
NOR_263: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_239,
        B => S423,
        Y => S1260
    );
NOR_264: ENTITY WORK.NOR
    PORT MAP (
        A => S435,
        B => S1260,
        Y => S1261
    );
NAND_670: ENTITY WORK.NAND
    PORT MAP (
        A => S1259,
        B => S1261,
        Y => S1262
    );
NOR_265: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_255,
        B => S423,
        Y => S1263
    );
NAND_671: ENTITY WORK.NAND
    PORT MAP (
        A => S7662,
        B => S423,
        Y => S1264
    );
NAND_672: ENTITY WORK.NAND
    PORT MAP (
        A => S435,
        B => S1264,
        Y => S1265
    );
NOR_266: ENTITY WORK.NOR
    PORT MAP (
        A => S1263,
        B => S1265,
        Y => S1266
    );
NAND_673: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_207,
        B => S436,
        Y => S1267
    );
NAND_674: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_223,
        B => S435,
        Y => S1268
    );
NAND_675: ENTITY WORK.NAND
    PORT MAP (
        A => S1267,
        B => S1268,
        Y => S1269
    );
NAND_676: ENTITY WORK.NAND
    PORT MAP (
        A => S422,
        B => S1269,
        Y => S1270
    );
NAND_677: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_143,
        B => S436,
        Y => S1271
    );
NAND_678: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_159,
        B => S435,
        Y => S1272
    );
NAND_679: ENTITY WORK.NAND
    PORT MAP (
        A => S1271,
        B => S1272,
        Y => S1273
    );
NAND_680: ENTITY WORK.NAND
    PORT MAP (
        A => S423,
        B => S1273,
        Y => S1274
    );
NAND_681: ENTITY WORK.NAND
    PORT MAP (
        A => S1270,
        B => S1274,
        Y => S1275
    );
NOR_267: ENTITY WORK.NOR
    PORT MAP (
        A => S441,
        B => S1275,
        Y => S1276
    );
NOR_268: ENTITY WORK.NOR
    PORT MAP (
        A => S442,
        B => S1266,
        Y => S1277
    );
NAND_682: ENTITY WORK.NAND
    PORT MAP (
        A => S1262,
        B => S1277,
        Y => S1278
    );
NAND_683: ENTITY WORK.NAND
    PORT MAP (
        A => S428,
        B => S1278,
        Y => S1279
    );
NOR_269: ENTITY WORK.NOR
    PORT MAP (
        A => S1276,
        B => S1279,
        Y => S1280
    );
NAND_684: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_127,
        B => S435,
        Y => S1281
    );
NAND_685: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_111,
        B => S436,
        Y => S1282
    );
NAND_686: ENTITY WORK.NAND
    PORT MAP (
        A => S1281,
        B => S1282,
        Y => S1283
    );
NAND_687: ENTITY WORK.NAND
    PORT MAP (
        A => S441,
        B => S1283,
        Y => S1284
    );
NAND_688: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_95,
        B => S435,
        Y => S1285
    );
NAND_689: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_79,
        B => S436,
        Y => S1286
    );
NAND_690: ENTITY WORK.NAND
    PORT MAP (
        A => S1285,
        B => S1286,
        Y => S1287
    );
NAND_691: ENTITY WORK.NAND
    PORT MAP (
        A => S442,
        B => S1287,
        Y => S1288
    );
NAND_692: ENTITY WORK.NAND
    PORT MAP (
        A => S1284,
        B => S1288,
        Y => S1289
    );
NAND_693: ENTITY WORK.NAND
    PORT MAP (
        A => S479,
        B => S1289,
        Y => S1290
    );
NAND_694: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_63,
        B => S435,
        Y => S1291
    );
NAND_695: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_47,
        B => S436,
        Y => S1292
    );
NAND_696: ENTITY WORK.NAND
    PORT MAP (
        A => S1291,
        B => S1292,
        Y => S1293
    );
NAND_697: ENTITY WORK.NAND
    PORT MAP (
        A => S441,
        B => S1293,
        Y => S1294
    );
NAND_698: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_31,
        B => S435,
        Y => S1295
    );
NAND_699: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_15,
        B => S436,
        Y => S1296
    );
NAND_700: ENTITY WORK.NAND
    PORT MAP (
        A => S1295,
        B => S1296,
        Y => S1297
    );
NAND_701: ENTITY WORK.NAND
    PORT MAP (
        A => S442,
        B => S1297,
        Y => S1298
    );
NAND_702: ENTITY WORK.NAND
    PORT MAP (
        A => S1294,
        B => S1298,
        Y => S1299
    );
NAND_703: ENTITY WORK.NAND
    PORT MAP (
        A => S429,
        B => S1299,
        Y => S1300
    );
NOT_158: ENTITY WORK.NOT
    PORT MAP (
        A => S1300,
        Y => S1301
    );
NOR_270: ENTITY WORK.NOR
    PORT MAP (
        A => S1280,
        B => S1301,
        Y => S1302
    );
NAND_704: ENTITY WORK.NAND
    PORT MAP (
        A => S1290,
        B => S1302,
        Y => S1303
    );
NAND_705: ENTITY WORK.NAND
    PORT MAP (
        A => S446,
        B => S1303,
        Y => S1304
    );
NOT_159: ENTITY WORK.NOT
    PORT MAP (
        A => S1304,
        Y => datapath_addsubunit_in1_15
    );
NAND_706: ENTITY WORK.NAND
    PORT MAP (
        A => S496,
        B => datapath_addsubunit_in1_15,
        Y => S1305
    );
NAND_707: ENTITY WORK.NAND
    PORT MAP (
        A => S372,
        B => S1305,
        Y => S1306
    );
NAND_708: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_15,
        B => S1306,
        Y => S1307
    );
NOT_160: ENTITY WORK.NOT
    PORT MAP (
        A => S1307,
        Y => S1308
    );
NOR_271: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_muxmem_in2_15,
        B => S1306,
        Y => S1309
    );
NOT_161: ENTITY WORK.NOT
    PORT MAP (
        A => S1309,
        Y => S1310
    );
NOR_272: ENTITY WORK.NOR
    PORT MAP (
        A => S1308,
        B => S1309,
        Y => S1311
    );
NAND_709: ENTITY WORK.NAND
    PORT MAP (
        A => S1307,
        B => S1310,
        Y => S1312
    );
NAND_710: ENTITY WORK.NAND
    PORT MAP (
        A => S1258,
        B => S1311,
        Y => S1313
    );
NAND_711: ENTITY WORK.NAND
    PORT MAP (
        A => S1257,
        B => S1312,
        Y => S1314
    );
NAND_712: ENTITY WORK.NAND
    PORT MAP (
        A => S1313,
        B => S1314,
        Y => S1315
    );
NAND_713: ENTITY WORK.NAND
    PORT MAP (
        A => S365,
        B => S1315,
        Y => S1316
    );
NOR_273: ENTITY WORK.NOR
    PORT MAP (
        A => controller_389_B_0,
        B => S348,
        Y => S1317
    );
NOR_274: ENTITY WORK.NOR
    PORT MAP (
        A => S346,
        B => S1317,
        Y => S1318
    );
NOR_275: ENTITY WORK.NOR
    PORT MAP (
        A => S8587,
        B => S1318,
        Y => S1319
    );
NAND_714: ENTITY WORK.NAND
    PORT MAP (
        A => S8587,
        B => S344,
        Y => S1320
    );
NOR_276: ENTITY WORK.NOR
    PORT MAP (
        A => S8225,
        B => S1320,
        Y => S1321
    );
NAND_715: ENTITY WORK.NAND
    PORT MAP (
        A => S8586,
        B => S8588,
        Y => S1322
    );
NOR_277: ENTITY WORK.NOR
    PORT MAP (
        A => controller_389_B_0,
        B => S353,
        Y => S1323
    );
NAND_716: ENTITY WORK.NAND
    PORT MAP (
        A => controller_389_B_0,
        B => S8584,
        Y => S1324
    );
NOR_278: ENTITY WORK.NOR
    PORT MAP (
        A => S1321,
        B => S1323,
        Y => S1325
    );
NAND_717: ENTITY WORK.NAND
    PORT MAP (
        A => S1322,
        B => S1324,
        Y => S1326
    );
NOR_279: ENTITY WORK.NOR
    PORT MAP (
        A => S8551,
        B => S1326,
        Y => S1327
    );
NAND_718: ENTITY WORK.NAND
    PORT MAP (
        A => S1325,
        B => S1327,
        Y => S1328
    );
NOR_280: ENTITY WORK.NOR
    PORT MAP (
        A => S1319,
        B => S1328,
        Y => S1329
    );
NOR_281: ENTITY WORK.NOR
    PORT MAP (
        A => S8554,
        B => S1329,
        Y => S1330
    );
NOR_282: ENTITY WORK.NOR
    PORT MAP (
        A => S8549,
        B => S1330,
        Y => S1331
    );
NOR_283: ENTITY WORK.NOR
    PORT MAP (
        A => S8385,
        B => S1331,
        Y => S1332
    );
NAND_719: ENTITY WORK.NAND
    PORT MAP (
        A => S8571,
        B => S8577,
        Y => S1333
    );
NOR_284: ENTITY WORK.NOR
    PORT MAP (
        A => S1332,
        B => S1333,
        Y => S1334
    );
NOR_285: ENTITY WORK.NOR
    PORT MAP (
        A => S7884,
        B => S7892,
        Y => S1335
    );
NAND_720: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_0,
        B => datapath_muxmem_in2_1,
        Y => S1336
    );
NOR_286: ENTITY WORK.NOR
    PORT MAP (
        A => S7897,
        B => S1336,
        Y => S1337
    );
NAND_721: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_2,
        B => S1335,
        Y => S1338
    );
NOR_287: ENTITY WORK.NOR
    PORT MAP (
        A => S7905,
        B => S1338,
        Y => S1339
    );
NAND_722: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_3,
        B => S1337,
        Y => S1340
    );
NAND_723: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_4,
        B => S1339,
        Y => S1341
    );
NOT_162: ENTITY WORK.NOT
    PORT MAP (
        A => S1341,
        Y => S1342
    );
NOR_288: ENTITY WORK.NOR
    PORT MAP (
        A => S7920,
        B => S1341,
        Y => S1343
    );
NAND_724: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_5,
        B => S1342,
        Y => S1344
    );
NOR_289: ENTITY WORK.NOR
    PORT MAP (
        A => S7928,
        B => S1344,
        Y => S1345
    );
NAND_725: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_6,
        B => S1343,
        Y => S1346
    );
NAND_726: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_7,
        B => S1345,
        Y => S1347
    );
NOT_163: ENTITY WORK.NOT
    PORT MAP (
        A => S1347,
        Y => S1348
    );
NOR_290: ENTITY WORK.NOR
    PORT MAP (
        A => S7946,
        B => S1347,
        Y => S1349
    );
NAND_727: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_8,
        B => S1348,
        Y => S1350
    );
NOR_291: ENTITY WORK.NOR
    PORT MAP (
        A => S7957,
        B => S1350,
        Y => S1351
    );
NAND_728: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_9,
        B => S1349,
        Y => S1352
    );
NOR_292: ENTITY WORK.NOR
    PORT MAP (
        A => S7968,
        B => S1352,
        Y => S1353
    );
NAND_729: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_10,
        B => S1351,
        Y => S1354
    );
NOR_293: ENTITY WORK.NOR
    PORT MAP (
        A => S7978,
        B => S1354,
        Y => S1355
    );
NAND_730: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_11,
        B => S1353,
        Y => S1356
    );
NOR_294: ENTITY WORK.NOR
    PORT MAP (
        A => S7989,
        B => S1356,
        Y => S1357
    );
NAND_731: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_12,
        B => S1355,
        Y => S1358
    );
NOR_295: ENTITY WORK.NOR
    PORT MAP (
        A => S8000,
        B => S1358,
        Y => S1359
    );
NAND_732: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_14,
        B => S1359,
        Y => S1360
    );
NAND_733: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_15,
        B => S1360,
        Y => S1361
    );
NOR_296: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_muxmem_in2_15,
        B => S1360,
        Y => S1362
    );
NOT_164: ENTITY WORK.NOT
    PORT MAP (
        A => S1362,
        Y => S1363
    );
NAND_734: ENTITY WORK.NAND
    PORT MAP (
        A => S1361,
        B => S1363,
        Y => S1364
    );
NOT_165: ENTITY WORK.NOT
    PORT MAP (
        A => S1364,
        Y => S1365
    );
NOR_297: ENTITY WORK.NOR
    PORT MAP (
        A => S1334,
        B => S1365,
        Y => S1366
    );
NAND_735: ENTITY WORK.NAND
    PORT MAP (
        A => controller_216_B_0,
        B => S8585,
        Y => S1367
    );
NAND_736: ENTITY WORK.NAND
    PORT MAP (
        A => S379,
        B => S1367,
        Y => S1368
    );
NOT_166: ENTITY WORK.NOT
    PORT MAP (
        A => S1368,
        Y => S1369
    );
NOR_298: ENTITY WORK.NOR
    PORT MAP (
        A => S358,
        B => S1368,
        Y => S1370
    );
NAND_737: ENTITY WORK.NAND
    PORT MAP (
        A => S359,
        B => S1369,
        Y => S1371
    );
NOR_299: ENTITY WORK.NOR
    PORT MAP (
        A => S1366,
        B => S1370,
        Y => S1372
    );
NAND_738: ENTITY WORK.NAND
    PORT MAP (
        A => S1316,
        B => S1372,
        Y => S1373
    );
NOR_300: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_15,
        B => S1371,
        Y => S1374
    );
NOR_301: ENTITY WORK.NOR
    PORT MAP (
        A => S8580,
        B => S1374,
        Y => S1375
    );
NAND_739: ENTITY WORK.NAND
    PORT MAP (
        A => S1373,
        B => S1375,
        Y => S1376
    );
NAND_740: ENTITY WORK.NAND
    PORT MAP (
        A => S8581,
        B => S1376,
        Y => S0
    );
NOR_302: ENTITY WORK.NOR
    PORT MAP (
        A => controller_pstate_0,
        B => S8569,
        Y => S1377
    );
NAND_741: ENTITY WORK.NAND
    PORT MAP (
        A => S8365,
        B => S8568,
        Y => S1378
    );
NOR_303: ENTITY WORK.NOR
    PORT MAP (
        A => S7476,
        B => S1377,
        Y => S1
    );
NAND_742: ENTITY WORK.NAND
    PORT MAP (
        A => S8356,
        B => S8365,
        Y => S1379
    );
NOT_167: ENTITY WORK.NOT
    PORT MAP (
        A => S1379,
        Y => controller_1115_S_0
    );
NAND_743: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_databusin_15,
        B => controller_1115_S_0,
        Y => S1380
    );
NAND_744: ENTITY WORK.NAND
    PORT MAP (
        A => controller_opcode_7,
        B => S1379,
        Y => S1381
    );
NAND_745: ENTITY WORK.NAND
    PORT MAP (
        A => S1380,
        B => S1381,
        Y => S2
    );
NOR_304: ENTITY WORK.NOR
    PORT MAP (
        A => controller_opcode_3,
        B => S369,
        Y => S1382
    );
NAND_746: ENTITY WORK.NAND
    PORT MAP (
        A => S8309,
        B => S368,
        Y => S1383
    );
NAND_747: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_adr_outreg_15,
        B => S1383,
        Y => S1384
    );
NAND_748: ENTITY WORK.NAND
    PORT MAP (
        A => S1306,
        B => S1382,
        Y => S1385
    );
NAND_749: ENTITY WORK.NAND
    PORT MAP (
        A => S1384,
        B => S1385,
        Y => S3
    );
NOR_305: ENTITY WORK.NOR
    PORT MAP (
        A => S8385,
        B => S383,
        Y => S1386
    );
NAND_750: ENTITY WORK.NAND
    PORT MAP (
        A => S8375,
        B => S382,
        Y => S1387
    );
NOR_306: ENTITY WORK.NOR
    PORT MAP (
        A => S8557,
        B => S1387,
        Y => S1388
    );
NAND_751: ENTITY WORK.NAND
    PORT MAP (
        A => S8375,
        B => S384,
        Y => S1389
    );
NOR_307: ENTITY WORK.NOR
    PORT MAP (
        A => S1220,
        B => S1389,
        Y => S1390
    );
NOR_308: ENTITY WORK.NOR
    PORT MAP (
        A => S8319,
        B => controller_opcode_5,
        Y => S1391
    );
NOT_168: ENTITY WORK.NOT
    PORT MAP (
        A => S1391,
        Y => S1392
    );
NAND_752: ENTITY WORK.NAND
    PORT MAP (
        A => S382,
        B => S1391,
        Y => S1393
    );
NAND_753: ENTITY WORK.NAND
    PORT MAP (
        A => S410,
        B => S1393,
        Y => S1394
    );
NOR_309: ENTITY WORK.NOR
    PORT MAP (
        A => S389,
        B => S1394,
        Y => S1395
    );
NOR_310: ENTITY WORK.NOR
    PORT MAP (
        A => S8385,
        B => S1395,
        Y => S1396
    );
NOT_169: ENTITY WORK.NOT
    PORT MAP (
        A => S1396,
        Y => S1397
    );
NAND_754: ENTITY WORK.NAND
    PORT MAP (
        A => S8375,
        B => S8416,
        Y => S1398
    );
NAND_755: ENTITY WORK.NAND
    PORT MAP (
        A => S8416,
        B => S1386,
        Y => S1399
    );
NOT_170: ENTITY WORK.NOT
    PORT MAP (
        A => S1399,
        Y => S1400
    );
NAND_756: ENTITY WORK.NAND
    PORT MAP (
        A => S1397,
        B => S1399,
        Y => S1401
    );
NOR_311: ENTITY WORK.NOR
    PORT MAP (
        A => controller_opcode_2,
        B => controller_opcode_3,
        Y => S1402
    );
NAND_757: ENTITY WORK.NAND
    PORT MAP (
        A => S8299,
        B => S8309,
        Y => S1403
    );
NOR_312: ENTITY WORK.NOR
    PORT MAP (
        A => S380,
        B => S1403,
        Y => S1404
    );
NAND_758: ENTITY WORK.NAND
    PORT MAP (
        A => S379,
        B => S1402,
        Y => S1405
    );
NOR_313: ENTITY WORK.NOR
    PORT MAP (
        A => S8278,
        B => S1405,
        Y => S1406
    );
NOT_171: ENTITY WORK.NOT
    PORT MAP (
        A => S1406,
        Y => S1407
    );
NOR_314: ENTITY WORK.NOR
    PORT MAP (
        A => S1401,
        B => S1406,
        Y => S1408
    );
NAND_759: ENTITY WORK.NAND
    PORT MAP (
        A => S371,
        B => S1408,
        Y => S1409
    );
NAND_760: ENTITY WORK.NAND
    PORT MAP (
        A => controller_fib_0,
        B => S1409,
        Y => S1410
    );
NOT_172: ENTITY WORK.NOT
    PORT MAP (
        A => S1410,
        Y => S1411
    );
NOR_315: ENTITY WORK.NOR
    PORT MAP (
        A => S1390,
        B => S1411,
        Y => S1412
    );
NOT_173: ENTITY WORK.NOT
    PORT MAP (
        A => S1412,
        Y => S1413
    );
NAND_761: ENTITY WORK.NAND
    PORT MAP (
        A => S8375,
        B => S392,
        Y => S1414
    );
NOT_174: ENTITY WORK.NOT
    PORT MAP (
        A => S1414,
        Y => S1415
    );
NOR_316: ENTITY WORK.NOR
    PORT MAP (
        A => S1406,
        B => S1415,
        Y => S1416
    );
NAND_762: ENTITY WORK.NAND
    PORT MAP (
        A => S1407,
        B => S1414,
        Y => S1417
    );
NAND_763: ENTITY WORK.NAND
    PORT MAP (
        A => S1413,
        B => S1417,
        Y => S1418
    );
NOR_317: ENTITY WORK.NOR
    PORT MAP (
        A => S401,
        B => S1403,
        Y => S1419
    );
NAND_764: ENTITY WORK.NAND
    PORT MAP (
        A => S400,
        B => S1402,
        Y => S1420
    );
NAND_765: ENTITY WORK.NAND
    PORT MAP (
        A => S8457,
        B => S8478,
        Y => S1421
    );
NOR_318: ENTITY WORK.NOR
    PORT MAP (
        A => S8557,
        B => S387,
        Y => S1422
    );
NOT_175: ENTITY WORK.NOT
    PORT MAP (
        A => S1422,
        Y => S1423
    );
NOR_319: ENTITY WORK.NOR
    PORT MAP (
        A => S8565,
        B => S387,
        Y => S1424
    );
NAND_766: ENTITY WORK.NAND
    PORT MAP (
        A => S1420,
        B => S1421,
        Y => S1425
    );
NOR_320: ENTITY WORK.NOR
    PORT MAP (
        A => S1419,
        B => S1424,
        Y => S1426
    );
NOR_321: ENTITY WORK.NOR
    PORT MAP (
        A => S1424,
        B => S1425,
        Y => S1427
    );
NAND_767: ENTITY WORK.NAND
    PORT MAP (
        A => S1421,
        B => S1426,
        Y => S1428
    );
NOR_322: ENTITY WORK.NOR
    PORT MAP (
        A => S8385,
        B => S1427,
        Y => S1429
    );
NAND_768: ENTITY WORK.NAND
    PORT MAP (
        A => S8375,
        B => S1428,
        Y => S1430
    );
NOR_323: ENTITY WORK.NOR
    PORT MAP (
        A => S8385,
        B => S1420,
        Y => S1431
    );
NAND_769: ENTITY WORK.NAND
    PORT MAP (
        A => S8375,
        B => S1419,
        Y => S1432
    );
NOR_324: ENTITY WORK.NOR
    PORT MAP (
        A => S8193,
        B => S1432,
        Y => S1433
    );
NAND_770: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_instruction_2,
        B => S1431,
        Y => S1434
    );
NOR_325: ENTITY WORK.NOR
    PORT MAP (
        A => S8299,
        B => S415,
        Y => S1435
    );
NAND_771: ENTITY WORK.NAND
    PORT MAP (
        A => controller_opcode_2,
        B => S414,
        Y => S1436
    );
NOR_326: ENTITY WORK.NOR
    PORT MAP (
        A => S1433,
        B => S1435,
        Y => S1437
    );
NAND_772: ENTITY WORK.NAND
    PORT MAP (
        A => S1434,
        B => S1436,
        Y => S1438
    );
NAND_773: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_instruction_1,
        B => S1431,
        Y => S1439
    );
NOT_176: ENTITY WORK.NOT
    PORT MAP (
        A => S1439,
        Y => S1440
    );
NAND_774: ENTITY WORK.NAND
    PORT MAP (
        A => controller_216_B_0,
        B => S414,
        Y => S1441
    );
NOT_177: ENTITY WORK.NOT
    PORT MAP (
        A => S1441,
        Y => S1442
    );
NOR_327: ENTITY WORK.NOR
    PORT MAP (
        A => S1440,
        B => S1442,
        Y => S1443
    );
NAND_775: ENTITY WORK.NAND
    PORT MAP (
        A => S1439,
        B => S1441,
        Y => S1444
    );
NAND_776: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_instruction_3,
        B => S1431,
        Y => S1445
    );
NOT_178: ENTITY WORK.NOT
    PORT MAP (
        A => S1445,
        Y => S1446
    );
NAND_777: ENTITY WORK.NAND
    PORT MAP (
        A => controller_opcode_3,
        B => S414,
        Y => S1447
    );
NOT_179: ENTITY WORK.NOT
    PORT MAP (
        A => S1447,
        Y => S1448
    );
NOR_328: ENTITY WORK.NOR
    PORT MAP (
        A => S1446,
        B => S1448,
        Y => S1449
    );
NAND_778: ENTITY WORK.NAND
    PORT MAP (
        A => S1445,
        B => S1447,
        Y => S1450
    );
NOR_329: ENTITY WORK.NOR
    PORT MAP (
        A => S1443,
        B => S1449,
        Y => S1451
    );
NAND_779: ENTITY WORK.NAND
    PORT MAP (
        A => S1444,
        B => S1450,
        Y => S1452
    );
NAND_780: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_instruction_0,
        B => S1431,
        Y => S1453
    );
NOT_180: ENTITY WORK.NOT
    PORT MAP (
        A => S1453,
        Y => S1454
    );
NAND_781: ENTITY WORK.NAND
    PORT MAP (
        A => controller_fib_4,
        B => S414,
        Y => S1455
    );
NOT_181: ENTITY WORK.NOT
    PORT MAP (
        A => S1455,
        Y => S1456
    );
NOR_330: ENTITY WORK.NOR
    PORT MAP (
        A => S1454,
        B => S1456,
        Y => S1457
    );
NAND_782: ENTITY WORK.NAND
    PORT MAP (
        A => S1453,
        B => S1455,
        Y => S1458
    );
NOR_331: ENTITY WORK.NOR
    PORT MAP (
        A => S1452,
        B => S1457,
        Y => S1459
    );
NAND_783: ENTITY WORK.NAND
    PORT MAP (
        A => S1451,
        B => S1458,
        Y => S1460
    );
NOR_332: ENTITY WORK.NOR
    PORT MAP (
        A => S1437,
        B => S1460,
        Y => S1461
    );
NAND_784: ENTITY WORK.NAND
    PORT MAP (
        A => S1438,
        B => S1459,
        Y => S1462
    );
NOR_333: ENTITY WORK.NOR
    PORT MAP (
        A => controller_outflag_0,
        B => S1462,
        Y => S1463
    );
NOT_182: ENTITY WORK.NOT
    PORT MAP (
        A => S1463,
        Y => S1464
    );
NAND_785: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_240,
        B => S1437,
        Y => S1465
    );
NAND_786: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_176,
        B => S1438,
        Y => S1466
    );
NAND_787: ENTITY WORK.NAND
    PORT MAP (
        A => S1465,
        B => S1466,
        Y => S1467
    );
NAND_788: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S1467,
        Y => S1468
    );
NAND_789: ENTITY WORK.NAND
    PORT MAP (
        A => S7783,
        B => S1437,
        Y => S1469
    );
NOR_334: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_160,
        B => S1437,
        Y => S1470
    );
NAND_790: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S1469,
        Y => S1471
    );
NOR_335: ENTITY WORK.NOR
    PORT MAP (
        A => S1470,
        B => S1471,
        Y => S1472
    );
NAND_791: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_208,
        B => S1437,
        Y => S1473
    );
NAND_792: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_144,
        B => S1438,
        Y => S1474
    );
NAND_793: ENTITY WORK.NAND
    PORT MAP (
        A => S1473,
        B => S1474,
        Y => S1475
    );
NAND_794: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S1475,
        Y => S1476
    );
NOR_336: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_128,
        B => S1437,
        Y => S1477
    );
NOR_337: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_192,
        B => S1438,
        Y => S1478
    );
NOR_338: ENTITY WORK.NOR
    PORT MAP (
        A => S1477,
        B => S1478,
        Y => S1479
    );
NAND_795: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S1479,
        Y => S1480
    );
NAND_796: ENTITY WORK.NAND
    PORT MAP (
        A => S1476,
        B => S1480,
        Y => S1481
    );
NOR_339: ENTITY WORK.NOR
    PORT MAP (
        A => S1443,
        B => S1481,
        Y => S1482
    );
NOR_340: ENTITY WORK.NOR
    PORT MAP (
        A => S1444,
        B => S1472,
        Y => S1483
    );
NAND_797: ENTITY WORK.NAND
    PORT MAP (
        A => S1468,
        B => S1483,
        Y => S1484
    );
NAND_798: ENTITY WORK.NAND
    PORT MAP (
        A => S1449,
        B => S1484,
        Y => S1485
    );
NOR_341: ENTITY WORK.NOR
    PORT MAP (
        A => S1482,
        B => S1485,
        Y => S1486
    );
NOR_342: ENTITY WORK.NOR
    PORT MAP (
        A => S1444,
        B => S1449,
        Y => S1487
    );
NAND_799: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_48,
        B => S1438,
        Y => S1488
    );
NAND_800: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_112,
        B => S1437,
        Y => S1489
    );
NAND_801: ENTITY WORK.NAND
    PORT MAP (
        A => S1488,
        B => S1489,
        Y => S1490
    );
NAND_802: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S1490,
        Y => S1491
    );
NAND_803: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_96,
        B => S1437,
        Y => S1492
    );
NAND_804: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_32,
        B => S1438,
        Y => S1493
    );
NAND_805: ENTITY WORK.NAND
    PORT MAP (
        A => S1492,
        B => S1493,
        Y => S1494
    );
NAND_806: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S1494,
        Y => S1495
    );
NAND_807: ENTITY WORK.NAND
    PORT MAP (
        A => S1491,
        B => S1495,
        Y => S1496
    );
NAND_808: ENTITY WORK.NAND
    PORT MAP (
        A => S1487,
        B => S1496,
        Y => S1497
    );
NOR_343: ENTITY WORK.NOR
    PORT MAP (
        A => S1438,
        B => S1458,
        Y => S1498
    );
NAND_809: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_80,
        B => S1498,
        Y => S1499
    );
NAND_810: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_16,
        B => S1438,
        Y => S1500
    );
NAND_811: ENTITY WORK.NAND
    PORT MAP (
        A => S1499,
        B => S1500,
        Y => S1501
    );
NOT_183: ENTITY WORK.NOT
    PORT MAP (
        A => S1501,
        Y => S1502
    );
NOR_344: ENTITY WORK.NOR
    PORT MAP (
        A => S1452,
        B => S1502,
        Y => S1503
    );
NAND_812: ENTITY WORK.NAND
    PORT MAP (
        A => S1451,
        B => S1501,
        Y => S1504
    );
NOR_345: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_64,
        B => S1438,
        Y => S1505
    );
NOT_184: ENTITY WORK.NOT
    PORT MAP (
        A => S1505,
        Y => S1506
    );
NOR_346: ENTITY WORK.NOR
    PORT MAP (
        A => S1460,
        B => S1505,
        Y => S1507
    );
NAND_813: ENTITY WORK.NAND
    PORT MAP (
        A => S1459,
        B => S1506,
        Y => S1508
    );
NOR_347: ENTITY WORK.NOR
    PORT MAP (
        A => S1503,
        B => S1507,
        Y => S1509
    );
NAND_814: ENTITY WORK.NAND
    PORT MAP (
        A => S1504,
        B => S1508,
        Y => S1510
    );
NAND_815: ENTITY WORK.NAND
    PORT MAP (
        A => S1497,
        B => S1509,
        Y => S1511
    );
NOR_348: ENTITY WORK.NOR
    PORT MAP (
        A => S1486,
        B => S1510,
        Y => S1512
    );
NOR_349: ENTITY WORK.NOR
    PORT MAP (
        A => S1486,
        B => S1511,
        Y => S1513
    );
NAND_816: ENTITY WORK.NAND
    PORT MAP (
        A => S1497,
        B => S1512,
        Y => S1514
    );
NOR_350: ENTITY WORK.NOR
    PORT MAP (
        A => S1463,
        B => S1513,
        Y => S1515
    );
NAND_817: ENTITY WORK.NAND
    PORT MAP (
        A => S1464,
        B => S1514,
        Y => S1516
    );
NAND_818: ENTITY WORK.NAND
    PORT MAP (
        A => S1429,
        B => S1515,
        Y => S1517
    );
NAND_819: ENTITY WORK.NAND
    PORT MAP (
        A => S1418,
        B => S1517,
        Y => S1518
    );
NOT_185: ENTITY WORK.NOT
    PORT MAP (
        A => S1518,
        Y => S1519
    );
NOR_351: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_0,
        B => S1519,
        Y => S1520
    );
NOR_352: ENTITY WORK.NOR
    PORT MAP (
        A => S1220,
        B => S1518,
        Y => S1521
    );
NOR_353: ENTITY WORK.NOR
    PORT MAP (
        A => S1520,
        B => S1521,
        Y => S1522
    );
NOR_354: ENTITY WORK.NOR
    PORT MAP (
        A => S409,
        B => S1422,
        Y => S1523
    );
NAND_820: ENTITY WORK.NAND
    PORT MAP (
        A => S410,
        B => S1423,
        Y => S1524
    );
NOR_355: ENTITY WORK.NOR
    PORT MAP (
        A => S8385,
        B => S1523,
        Y => S1525
    );
NAND_821: ENTITY WORK.NAND
    PORT MAP (
        A => S8375,
        B => S1524,
        Y => S1526
    );
NOR_356: ENTITY WORK.NOR
    PORT MAP (
        A => S378,
        B => S387,
        Y => S1527
    );
NAND_822: ENTITY WORK.NAND
    PORT MAP (
        A => S8375,
        B => S388,
        Y => S1528
    );
NOR_357: ENTITY WORK.NOR
    PORT MAP (
        A => S1525,
        B => S1527,
        Y => S1529
    );
NOR_358: ENTITY WORK.NOR
    PORT MAP (
        A => S1522,
        B => S1529,
        Y => S1530
    );
NAND_823: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_0,
        B => S1518,
        Y => S1531
    );
NOR_359: ENTITY WORK.NOR
    PORT MAP (
        A => S8385,
        B => S1421,
        Y => S1532
    );
NOR_360: ENTITY WORK.NOR
    PORT MAP (
        A => S1400,
        B => S1532,
        Y => S1533
    );
NOT_186: ENTITY WORK.NOT
    PORT MAP (
        A => S1533,
        Y => S1534
    );
NOR_361: ENTITY WORK.NOR
    PORT MAP (
        A => S1531,
        B => S1533,
        Y => S1535
    );
NOT_187: ENTITY WORK.NOT
    PORT MAP (
        A => S1535,
        Y => S1536
    );
NAND_824: ENTITY WORK.NAND
    PORT MAP (
        A => controller_opcode_3,
        B => S379,
        Y => S1537
    );
NOR_362: ENTITY WORK.NOR
    PORT MAP (
        A => S366,
        B => S380,
        Y => S1538
    );
NAND_825: ENTITY WORK.NAND
    PORT MAP (
        A => S367,
        B => S379,
        Y => S1539
    );
NOR_363: ENTITY WORK.NOR
    PORT MAP (
        A => S8267,
        B => S1539,
        Y => S1540
    );
NAND_826: ENTITY WORK.NAND
    PORT MAP (
        A => S1220,
        B => S1540,
        Y => S1541
    );
NOT_188: ENTITY WORK.NOT
    PORT MAP (
        A => S1541,
        Y => S1542
    );
NOR_364: ENTITY WORK.NOR
    PORT MAP (
        A => S1220,
        B => S1540,
        Y => S1543
    );
NOR_365: ENTITY WORK.NOR
    PORT MAP (
        A => S1539,
        B => S1543,
        Y => S1544
    );
NAND_827: ENTITY WORK.NAND
    PORT MAP (
        A => S1541,
        B => S1544,
        Y => S1545
    );
NOR_366: ENTITY WORK.NOR
    PORT MAP (
        A => S8565,
        B => S1387,
        Y => S1546
    );
NAND_828: ENTITY WORK.NAND
    PORT MAP (
        A => S8564,
        B => S1386,
        Y => S1547
    );
NOR_367: ENTITY WORK.NOR
    PORT MAP (
        A => S1412,
        B => S1547,
        Y => S1548
    );
NOR_368: ENTITY WORK.NOR
    PORT MAP (
        A => controller_389_B_0,
        B => S1462,
        Y => S1549
    );
NOT_189: ENTITY WORK.NOT
    PORT MAP (
        A => S1549,
        Y => S1550
    );
NAND_829: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_244,
        B => S1437,
        Y => S1551
    );
NAND_830: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_180,
        B => S1438,
        Y => S1552
    );
NAND_831: ENTITY WORK.NAND
    PORT MAP (
        A => S1551,
        B => S1552,
        Y => S1553
    );
NAND_832: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S1553,
        Y => S1554
    );
NAND_833: ENTITY WORK.NAND
    PORT MAP (
        A => S7816,
        B => S1437,
        Y => S1555
    );
NOR_369: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_164,
        B => S1437,
        Y => S1556
    );
NAND_834: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S1555,
        Y => S1557
    );
NOR_370: ENTITY WORK.NOR
    PORT MAP (
        A => S1556,
        B => S1557,
        Y => S1558
    );
NAND_835: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_148,
        B => S1438,
        Y => S1559
    );
NAND_836: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_212,
        B => S1437,
        Y => S1560
    );
NAND_837: ENTITY WORK.NAND
    PORT MAP (
        A => S1559,
        B => S1560,
        Y => S1561
    );
NAND_838: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S1561,
        Y => S1562
    );
NOR_371: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_132,
        B => S1437,
        Y => S1563
    );
NOR_372: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_196,
        B => S1438,
        Y => S1564
    );
NOR_373: ENTITY WORK.NOR
    PORT MAP (
        A => S1563,
        B => S1564,
        Y => S1565
    );
NAND_839: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S1565,
        Y => S1566
    );
NAND_840: ENTITY WORK.NAND
    PORT MAP (
        A => S1562,
        B => S1566,
        Y => S1567
    );
NOR_374: ENTITY WORK.NOR
    PORT MAP (
        A => S1443,
        B => S1567,
        Y => S1568
    );
NOR_375: ENTITY WORK.NOR
    PORT MAP (
        A => S1444,
        B => S1558,
        Y => S1569
    );
NAND_841: ENTITY WORK.NAND
    PORT MAP (
        A => S1554,
        B => S1569,
        Y => S1570
    );
NAND_842: ENTITY WORK.NAND
    PORT MAP (
        A => S1449,
        B => S1570,
        Y => S1571
    );
NOR_376: ENTITY WORK.NOR
    PORT MAP (
        A => S1568,
        B => S1571,
        Y => S1572
    );
NAND_843: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_100,
        B => S1458,
        Y => S1573
    );
NAND_844: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_116,
        B => S1457,
        Y => S1574
    );
NAND_845: ENTITY WORK.NAND
    PORT MAP (
        A => S1573,
        B => S1574,
        Y => S1575
    );
NAND_846: ENTITY WORK.NAND
    PORT MAP (
        A => S1437,
        B => S1575,
        Y => S1576
    );
NAND_847: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_36,
        B => S1458,
        Y => S1577
    );
NAND_848: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_52,
        B => S1457,
        Y => S1578
    );
NAND_849: ENTITY WORK.NAND
    PORT MAP (
        A => S1577,
        B => S1578,
        Y => S1579
    );
NAND_850: ENTITY WORK.NAND
    PORT MAP (
        A => S1438,
        B => S1579,
        Y => S1580
    );
NAND_851: ENTITY WORK.NAND
    PORT MAP (
        A => S1576,
        B => S1580,
        Y => S1581
    );
NAND_852: ENTITY WORK.NAND
    PORT MAP (
        A => S1487,
        B => S1581,
        Y => S1582
    );
NAND_853: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_84,
        B => S1498,
        Y => S1583
    );
NOR_377: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_68,
        B => S1438,
        Y => S1584
    );
NOT_190: ENTITY WORK.NOT
    PORT MAP (
        A => S1584,
        Y => S1585
    );
NAND_854: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_20,
        B => S1438,
        Y => S1586
    );
NAND_855: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S1586,
        Y => S1587
    );
NAND_856: ENTITY WORK.NAND
    PORT MAP (
        A => S1585,
        B => S1587,
        Y => S1588
    );
NAND_857: ENTITY WORK.NAND
    PORT MAP (
        A => S1583,
        B => S1588,
        Y => S1589
    );
NOT_191: ENTITY WORK.NOT
    PORT MAP (
        A => S1589,
        Y => S1590
    );
NOR_378: ENTITY WORK.NOR
    PORT MAP (
        A => S1452,
        B => S1590,
        Y => S1591
    );
NAND_858: ENTITY WORK.NAND
    PORT MAP (
        A => S1451,
        B => S1589,
        Y => S1592
    );
NAND_859: ENTITY WORK.NAND
    PORT MAP (
        A => S1582,
        B => S1592,
        Y => S1593
    );
NOR_379: ENTITY WORK.NOR
    PORT MAP (
        A => S1572,
        B => S1591,
        Y => S1594
    );
NOR_380: ENTITY WORK.NOR
    PORT MAP (
        A => S1572,
        B => S1593,
        Y => S1595
    );
NAND_860: ENTITY WORK.NAND
    PORT MAP (
        A => S1582,
        B => S1594,
        Y => S1596
    );
NOR_381: ENTITY WORK.NOR
    PORT MAP (
        A => S1549,
        B => S1595,
        Y => S1597
    );
NAND_861: ENTITY WORK.NAND
    PORT MAP (
        A => S1550,
        B => S1596,
        Y => S1598
    );
NOR_382: ENTITY WORK.NOR
    PORT MAP (
        A => S8468,
        B => S1387,
        Y => S1599
    );
NAND_862: ENTITY WORK.NAND
    PORT MAP (
        A => S8457,
        B => S1386,
        Y => S1600
    );
NOR_383: ENTITY WORK.NOR
    PORT MAP (
        A => S8426,
        B => S387,
        Y => S1601
    );
NOR_384: ENTITY WORK.NOR
    PORT MAP (
        A => S387,
        B => S1398,
        Y => S1602
    );
NAND_863: ENTITY WORK.NAND
    PORT MAP (
        A => S8375,
        B => S1601,
        Y => S1603
    );
NOR_385: ENTITY WORK.NOR
    PORT MAP (
        A => S1599,
        B => S1602,
        Y => S1604
    );
NAND_864: ENTITY WORK.NAND
    PORT MAP (
        A => S1600,
        B => S1603,
        Y => S1605
    );
NAND_865: ENTITY WORK.NAND
    PORT MAP (
        A => S1597,
        B => S1605,
        Y => S1606
    );
NOR_386: ENTITY WORK.NOR
    PORT MAP (
        A => S8385,
        B => S8545,
        Y => S1607
    );
NAND_866: ENTITY WORK.NAND
    PORT MAP (
        A => controller_fib_4,
        B => S1607,
        Y => S1608
    );
NAND_867: ENTITY WORK.NAND
    PORT MAP (
        A => S1606,
        B => S1608,
        Y => S1609
    );
NAND_868: ENTITY WORK.NAND
    PORT MAP (
        A => controller_216_B_0,
        B => S1607,
        Y => S1610
    );
NAND_869: ENTITY WORK.NAND
    PORT MAP (
        A => S1603,
        B => S1610,
        Y => S1611
    );
NOT_192: ENTITY WORK.NOT
    PORT MAP (
        A => S1611,
        Y => S1612
    );
NOR_387: ENTITY WORK.NOR
    PORT MAP (
        A => S1605,
        B => S1607,
        Y => S1613
    );
NOR_388: ENTITY WORK.NOR
    PORT MAP (
        A => S1609,
        B => S1613,
        Y => S1614
    );
NAND_870: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_shiftunit_2135_A,
        B => S1614,
        Y => S1615
    );
NAND_871: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_shiftunit_2439_A,
        B => S1609,
        Y => S1616
    );
NAND_872: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu2_0,
        B => S8570,
        Y => S1617
    );
NOR_389: ENTITY WORK.NOR
    PORT MAP (
        A => controller_216_B_0,
        B => controller_opcode_2,
        Y => S1618
    );
NOT_193: ENTITY WORK.NOT
    PORT MAP (
        A => S1618,
        Y => S1619
    );
NOR_390: ENTITY WORK.NOR
    PORT MAP (
        A => S8309,
        B => S1618,
        Y => S1620
    );
NAND_873: ENTITY WORK.NAND
    PORT MAP (
        A => controller_opcode_3,
        B => S1619,
        Y => S1621
    );
NOR_391: ENTITY WORK.NOR
    PORT MAP (
        A => S369,
        B => S1621,
        Y => S1622
    );
NAND_874: ENTITY WORK.NAND
    PORT MAP (
        A => S368,
        B => S1620,
        Y => S1623
    );
NAND_875: ENTITY WORK.NAND
    PORT MAP (
        A => S7884,
        B => S1622,
        Y => S1624
    );
NAND_876: ENTITY WORK.NAND
    PORT MAP (
        A => S1617,
        B => S1624,
        Y => S1625
    );
NAND_877: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu1_0,
        B => S1377,
        Y => S1626
    );
NOR_392: ENTITY WORK.NOR
    PORT MAP (
        A => controller_opcode_2,
        B => S8577,
        Y => S1627
    );
NAND_878: ENTITY WORK.NAND
    PORT MAP (
        A => S8299,
        B => S8576,
        Y => S1628
    );
NAND_879: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_databusin_0,
        B => S1627,
        Y => S1629
    );
NAND_880: ENTITY WORK.NAND
    PORT MAP (
        A => S1626,
        B => S1629,
        Y => S1630
    );
NOR_393: ENTITY WORK.NOR
    PORT MAP (
        A => S1625,
        B => S1630,
        Y => S1631
    );
NAND_881: ENTITY WORK.NAND
    PORT MAP (
        A => S1616,
        B => S1631,
        Y => S1632
    );
NOT_194: ENTITY WORK.NOT
    PORT MAP (
        A => S1632,
        Y => S1633
    );
NAND_882: ENTITY WORK.NAND
    PORT MAP (
        A => S1615,
        B => S1633,
        Y => S1634
    );
NOR_394: ENTITY WORK.NOR
    PORT MAP (
        A => S1548,
        B => S1634,
        Y => S1635
    );
NAND_883: ENTITY WORK.NAND
    PORT MAP (
        A => S1536,
        B => S1635,
        Y => S1636
    );
NOR_395: ENTITY WORK.NOR
    PORT MAP (
        A => S1530,
        B => S1636,
        Y => S1637
    );
NAND_884: ENTITY WORK.NAND
    PORT MAP (
        A => S1545,
        B => S1637,
        Y => datapath_indatatrf_0
    );
NAND_885: ENTITY WORK.NAND
    PORT MAP (
        A => S8375,
        B => S8520,
        Y => S1638
    );
NAND_886: ENTITY WORK.NAND
    PORT MAP (
        A => S1537,
        B => S1638,
        Y => S1639
    );
NOR_396: ENTITY WORK.NOR
    PORT MAP (
        A => S1622,
        B => S1639,
        Y => S1640
    );
NOR_397: ENTITY WORK.NOR
    PORT MAP (
        A => S1377,
        B => S1627,
        Y => S1641
    );
NAND_887: ENTITY WORK.NAND
    PORT MAP (
        A => S1640,
        B => S1641,
        Y => S1642
    );
NOT_195: ENTITY WORK.NOT
    PORT MAP (
        A => S1642,
        Y => S1643
    );
NAND_888: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_instruction_0,
        B => datapath_instruction_1,
        Y => S1644
    );
NOT_196: ENTITY WORK.NOT
    PORT MAP (
        A => S1644,
        Y => S1645
    );
NAND_889: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_instruction_2,
        B => S1645,
        Y => S1646
    );
NAND_890: ENTITY WORK.NAND
    PORT MAP (
        A => S8570,
        B => S1646,
        Y => S1647
    );
NOT_197: ENTITY WORK.NOT
    PORT MAP (
        A => S1647,
        Y => S1648
    );
NOR_398: ENTITY WORK.NOR
    PORT MAP (
        A => S1642,
        B => S1648,
        Y => S1649
    );
NAND_891: ENTITY WORK.NAND
    PORT MAP (
        A => S1643,
        B => S1647,
        Y => S1650
    );
NOR_399: ENTITY WORK.NOR
    PORT MAP (
        A => S8571,
        B => S1644,
        Y => S1651
    );
NOR_400: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_instruction_2,
        B => S1651,
        Y => S1652
    );
NOT_198: ENTITY WORK.NOT
    PORT MAP (
        A => S1652,
        Y => S1653
    );
NOR_401: ENTITY WORK.NOR
    PORT MAP (
        A => S1649,
        B => S1652,
        Y => S1654
    );
NAND_892: ENTITY WORK.NAND
    PORT MAP (
        A => S1650,
        B => S1653,
        Y => S1655
    );
NOR_402: ENTITY WORK.NOR
    PORT MAP (
        A => S8571,
        B => S1646,
        Y => S1656
    );
NOR_403: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_instruction_3,
        B => S1656,
        Y => S1657
    );
NOT_199: ENTITY WORK.NOT
    PORT MAP (
        A => S1657,
        Y => S1658
    );
NOR_404: ENTITY WORK.NOR
    PORT MAP (
        A => S8204,
        B => S1650,
        Y => S1659
    );
NAND_893: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_instruction_3,
        B => S1649,
        Y => S1660
    );
NOR_405: ENTITY WORK.NOR
    PORT MAP (
        A => S1657,
        B => S1659,
        Y => S1661
    );
NAND_894: ENTITY WORK.NAND
    PORT MAP (
        A => S1658,
        B => S1660,
        Y => S1662
    );
NOR_406: ENTITY WORK.NOR
    PORT MAP (
        A => S1654,
        B => S1662,
        Y => S1663
    );
NAND_895: ENTITY WORK.NAND
    PORT MAP (
        A => S1655,
        B => S1661,
        Y => S1664
    );
NOR_407: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_instruction_0,
        B => datapath_instruction_1,
        Y => S1665
    );
NOT_200: ENTITY WORK.NOT
    PORT MAP (
        A => S1665,
        Y => S1666
    );
NAND_896: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_instruction_1,
        B => S1642,
        Y => S1667
    );
NAND_897: ENTITY WORK.NAND
    PORT MAP (
        A => S8570,
        B => S1644,
        Y => S1668
    );
NAND_898: ENTITY WORK.NAND
    PORT MAP (
        A => S1667,
        B => S1668,
        Y => S1669
    );
NOT_201: ENTITY WORK.NOT
    PORT MAP (
        A => S1669,
        Y => S1670
    );
NOR_408: ENTITY WORK.NOR
    PORT MAP (
        A => S1665,
        B => S1670,
        Y => S1671
    );
NAND_899: ENTITY WORK.NAND
    PORT MAP (
        A => S1666,
        B => S1669,
        Y => S1672
    );
NOR_409: ENTITY WORK.NOR
    PORT MAP (
        A => S1664,
        B => S1672,
        Y => S1673
    );
NAND_900: ENTITY WORK.NAND
    PORT MAP (
        A => S1663,
        B => S1671,
        Y => S1674
    );
NOR_410: ENTITY WORK.NOR
    PORT MAP (
        A => S8572,
        B => S1628,
        Y => S1675
    );
NOR_411: ENTITY WORK.NOR
    PORT MAP (
        A => S8568,
        B => S1675,
        Y => S1676
    );
NAND_901: ENTITY WORK.NAND
    PORT MAP (
        A => S8569,
        B => S1640,
        Y => S1677
    );
NOR_412: ENTITY WORK.NOR
    PORT MAP (
        A => S1675,
        B => S1677,
        Y => S1678
    );
NAND_902: ENTITY WORK.NAND
    PORT MAP (
        A => S1640,
        B => S1676,
        Y => S1679
    );
NAND_903: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_instruction_0,
        B => S1642,
        Y => S1680
    );
NOT_202: ENTITY WORK.NOT
    PORT MAP (
        A => S1680,
        Y => S1681
    );
NOR_413: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_instruction_0,
        B => S8571,
        Y => S1682
    );
NOT_203: ENTITY WORK.NOT
    PORT MAP (
        A => S1682,
        Y => S1683
    );
NOR_414: ENTITY WORK.NOR
    PORT MAP (
        A => S1681,
        B => S1682,
        Y => S1684
    );
NAND_904: ENTITY WORK.NAND
    PORT MAP (
        A => S1680,
        B => S1683,
        Y => S1685
    );
NOR_415: ENTITY WORK.NOR
    PORT MAP (
        A => S1678,
        B => S1684,
        Y => S1686
    );
NAND_905: ENTITY WORK.NAND
    PORT MAP (
        A => S1679,
        B => S1685,
        Y => S1687
    );
NOR_416: ENTITY WORK.NOR
    PORT MAP (
        A => S1674,
        B => S1687,
        Y => S1688
    );
NAND_906: ENTITY WORK.NAND
    PORT MAP (
        A => S1673,
        B => S1686,
        Y => S1689
    );
NAND_907: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_0,
        B => S1688,
        Y => S1690
    );
NAND_908: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_64,
        B => S1689,
        Y => S1691
    );
NAND_909: ENTITY WORK.NAND
    PORT MAP (
        A => S1690,
        B => S1691,
        Y => S4
    );
NOR_417: ENTITY WORK.NOR
    PORT MAP (
        A => S1168,
        B => S1389,
        Y => S1692
    );
NAND_910: ENTITY WORK.NAND
    PORT MAP (
        A => controller_fib_1,
        B => S1409,
        Y => S1693
    );
NOT_204: ENTITY WORK.NOT
    PORT MAP (
        A => S1693,
        Y => S1694
    );
NOR_418: ENTITY WORK.NOR
    PORT MAP (
        A => S1692,
        B => S1694,
        Y => S1695
    );
NOR_419: ENTITY WORK.NOR
    PORT MAP (
        A => S1416,
        B => S1695,
        Y => S1696
    );
NOR_420: ENTITY WORK.NOR
    PORT MAP (
        A => controller_outflag_1,
        B => S1462,
        Y => S1697
    );
NOT_205: ENTITY WORK.NOT
    PORT MAP (
        A => S1697,
        Y => S1698
    );
NAND_911: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_241,
        B => S1437,
        Y => S1699
    );
NAND_912: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_177,
        B => S1438,
        Y => S1700
    );
NAND_913: ENTITY WORK.NAND
    PORT MAP (
        A => S1699,
        B => S1700,
        Y => S1701
    );
NAND_914: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S1701,
        Y => S1702
    );
NAND_915: ENTITY WORK.NAND
    PORT MAP (
        A => S7794,
        B => S1437,
        Y => S1703
    );
NOR_421: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_161,
        B => S1437,
        Y => S1704
    );
NAND_916: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S1703,
        Y => S1705
    );
NOR_422: ENTITY WORK.NOR
    PORT MAP (
        A => S1704,
        B => S1705,
        Y => S1706
    );
NAND_917: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_145,
        B => S1438,
        Y => S1707
    );
NAND_918: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_209,
        B => S1437,
        Y => S1708
    );
NAND_919: ENTITY WORK.NAND
    PORT MAP (
        A => S1707,
        B => S1708,
        Y => S1709
    );
NAND_920: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S1709,
        Y => S1710
    );
NOR_423: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_129,
        B => S1437,
        Y => S1711
    );
NOR_424: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_193,
        B => S1438,
        Y => S1712
    );
NOR_425: ENTITY WORK.NOR
    PORT MAP (
        A => S1711,
        B => S1712,
        Y => S1713
    );
NAND_921: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S1713,
        Y => S1714
    );
NAND_922: ENTITY WORK.NAND
    PORT MAP (
        A => S1710,
        B => S1714,
        Y => S1715
    );
NOR_426: ENTITY WORK.NOR
    PORT MAP (
        A => S1443,
        B => S1715,
        Y => S1716
    );
NOR_427: ENTITY WORK.NOR
    PORT MAP (
        A => S1444,
        B => S1706,
        Y => S1717
    );
NAND_923: ENTITY WORK.NAND
    PORT MAP (
        A => S1702,
        B => S1717,
        Y => S1718
    );
NAND_924: ENTITY WORK.NAND
    PORT MAP (
        A => S1449,
        B => S1718,
        Y => S1719
    );
NOR_428: ENTITY WORK.NOR
    PORT MAP (
        A => S1716,
        B => S1719,
        Y => S1720
    );
NAND_925: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_97,
        B => S1458,
        Y => S1721
    );
NAND_926: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_113,
        B => S1457,
        Y => S1722
    );
NAND_927: ENTITY WORK.NAND
    PORT MAP (
        A => S1721,
        B => S1722,
        Y => S1723
    );
NAND_928: ENTITY WORK.NAND
    PORT MAP (
        A => S1437,
        B => S1723,
        Y => S1724
    );
NAND_929: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_33,
        B => S1458,
        Y => S1725
    );
NAND_930: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_49,
        B => S1457,
        Y => S1726
    );
NAND_931: ENTITY WORK.NAND
    PORT MAP (
        A => S1725,
        B => S1726,
        Y => S1727
    );
NAND_932: ENTITY WORK.NAND
    PORT MAP (
        A => S1438,
        B => S1727,
        Y => S1728
    );
NAND_933: ENTITY WORK.NAND
    PORT MAP (
        A => S1724,
        B => S1728,
        Y => S1729
    );
NAND_934: ENTITY WORK.NAND
    PORT MAP (
        A => S1487,
        B => S1729,
        Y => S1730
    );
NAND_935: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_81,
        B => S1498,
        Y => S1731
    );
NOR_429: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_65,
        B => S1438,
        Y => S1732
    );
NOT_206: ENTITY WORK.NOT
    PORT MAP (
        A => S1732,
        Y => S1733
    );
NAND_936: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_17,
        B => S1438,
        Y => S1734
    );
NAND_937: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S1734,
        Y => S1735
    );
NAND_938: ENTITY WORK.NAND
    PORT MAP (
        A => S1733,
        B => S1735,
        Y => S1736
    );
NAND_939: ENTITY WORK.NAND
    PORT MAP (
        A => S1731,
        B => S1736,
        Y => S1737
    );
NOT_207: ENTITY WORK.NOT
    PORT MAP (
        A => S1737,
        Y => S1738
    );
NOR_430: ENTITY WORK.NOR
    PORT MAP (
        A => S1452,
        B => S1738,
        Y => S1739
    );
NAND_940: ENTITY WORK.NAND
    PORT MAP (
        A => S1451,
        B => S1737,
        Y => S1740
    );
NAND_941: ENTITY WORK.NAND
    PORT MAP (
        A => S1730,
        B => S1740,
        Y => S1741
    );
NOR_431: ENTITY WORK.NOR
    PORT MAP (
        A => S1720,
        B => S1739,
        Y => S1742
    );
NOR_432: ENTITY WORK.NOR
    PORT MAP (
        A => S1720,
        B => S1741,
        Y => S1743
    );
NAND_942: ENTITY WORK.NAND
    PORT MAP (
        A => S1730,
        B => S1742,
        Y => S1744
    );
NOR_433: ENTITY WORK.NOR
    PORT MAP (
        A => S1697,
        B => S1743,
        Y => S1745
    );
NAND_943: ENTITY WORK.NAND
    PORT MAP (
        A => S1698,
        B => S1744,
        Y => S1746
    );
NOR_434: ENTITY WORK.NOR
    PORT MAP (
        A => S1430,
        B => S1746,
        Y => S1747
    );
NOR_435: ENTITY WORK.NOR
    PORT MAP (
        A => S1696,
        B => S1747,
        Y => S1748
    );
NOT_208: ENTITY WORK.NOT
    PORT MAP (
        A => S1748,
        Y => S1749
    );
NOR_436: ENTITY WORK.NOR
    PORT MAP (
        A => S1168,
        B => S1749,
        Y => S1750
    );
NAND_944: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_1,
        B => S1748,
        Y => S1751
    );
NAND_945: ENTITY WORK.NAND
    PORT MAP (
        A => S1168,
        B => S1749,
        Y => S1752
    );
NOT_209: ENTITY WORK.NOT
    PORT MAP (
        A => S1752,
        Y => S1753
    );
NOR_437: ENTITY WORK.NOR
    PORT MAP (
        A => S1750,
        B => S1753,
        Y => S1754
    );
NOT_210: ENTITY WORK.NOT
    PORT MAP (
        A => S1754,
        Y => S1755
    );
NAND_946: ENTITY WORK.NAND
    PORT MAP (
        A => S1520,
        B => S1755,
        Y => S1756
    );
NOR_438: ENTITY WORK.NOR
    PORT MAP (
        A => S1520,
        B => S1755,
        Y => S1757
    );
NOR_439: ENTITY WORK.NOR
    PORT MAP (
        A => S1526,
        B => S1757,
        Y => S1758
    );
NAND_947: ENTITY WORK.NAND
    PORT MAP (
        A => S1756,
        B => S1758,
        Y => S1759
    );
NOR_440: ENTITY WORK.NOR
    PORT MAP (
        A => S1531,
        B => S1754,
        Y => S1760
    );
NOT_211: ENTITY WORK.NOT
    PORT MAP (
        A => S1760,
        Y => S1761
    );
NAND_948: ENTITY WORK.NAND
    PORT MAP (
        A => S1531,
        B => S1754,
        Y => S1762
    );
NAND_949: ENTITY WORK.NAND
    PORT MAP (
        A => S1527,
        B => S1762,
        Y => S1763
    );
NOR_441: ENTITY WORK.NOR
    PORT MAP (
        A => S1760,
        B => S1763,
        Y => S1764
    );
NOR_442: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_1,
        B => S1541,
        Y => S1765
    );
NOT_212: ENTITY WORK.NOT
    PORT MAP (
        A => S1765,
        Y => S1766
    );
NOR_443: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_1,
        B => S1539,
        Y => S1767
    );
NOR_444: ENTITY WORK.NOR
    PORT MAP (
        A => S1542,
        B => S1767,
        Y => S1768
    );
NOR_445: ENTITY WORK.NOR
    PORT MAP (
        A => S1765,
        B => S1768,
        Y => S1769
    );
NOR_446: ENTITY WORK.NOR
    PORT MAP (
        A => S1547,
        B => S1695,
        Y => S1770
    );
NAND_950: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_shiftunit_2153_A,
        B => S1614,
        Y => S1771
    );
NOR_447: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_muxmem_in2_0,
        B => datapath_muxmem_in2_1,
        Y => S1772
    );
NOR_448: ENTITY WORK.NOR
    PORT MAP (
        A => S1335,
        B => S1772,
        Y => S1773
    );
NOT_213: ENTITY WORK.NOT
    PORT MAP (
        A => S1773,
        Y => S1774
    );
NAND_951: ENTITY WORK.NAND
    PORT MAP (
        A => S1622,
        B => S1773,
        Y => S1775
    );
NAND_952: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu2_1,
        B => S8570,
        Y => S1776
    );
NAND_953: ENTITY WORK.NAND
    PORT MAP (
        A => S1775,
        B => S1776,
        Y => S1777
    );
NAND_954: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu1_1,
        B => S1377,
        Y => S1778
    );
NAND_955: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_databusin_1,
        B => S1627,
        Y => S1779
    );
NAND_956: ENTITY WORK.NAND
    PORT MAP (
        A => S1778,
        B => S1779,
        Y => S1780
    );
NOR_449: ENTITY WORK.NOR
    PORT MAP (
        A => S1777,
        B => S1780,
        Y => S1781
    );
NAND_957: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_shiftunit_2457_A,
        B => S1609,
        Y => S1782
    );
NAND_958: ENTITY WORK.NAND
    PORT MAP (
        A => S1771,
        B => S1781,
        Y => S1783
    );
NOR_450: ENTITY WORK.NOR
    PORT MAP (
        A => S1770,
        B => S1783,
        Y => S1784
    );
NAND_959: ENTITY WORK.NAND
    PORT MAP (
        A => S1782,
        B => S1784,
        Y => S1785
    );
NOR_451: ENTITY WORK.NOR
    PORT MAP (
        A => S1769,
        B => S1785,
        Y => S1786
    );
NOR_452: ENTITY WORK.NOR
    PORT MAP (
        A => S1168,
        B => S1748,
        Y => S1787
    );
NOT_214: ENTITY WORK.NOT
    PORT MAP (
        A => S1787,
        Y => S1788
    );
NAND_960: ENTITY WORK.NAND
    PORT MAP (
        A => S1534,
        B => S1787,
        Y => S1789
    );
NAND_961: ENTITY WORK.NAND
    PORT MAP (
        A => S1786,
        B => S1789,
        Y => S1790
    );
NOR_453: ENTITY WORK.NOR
    PORT MAP (
        A => S1764,
        B => S1790,
        Y => S1791
    );
NAND_962: ENTITY WORK.NAND
    PORT MAP (
        A => S1759,
        B => S1791,
        Y => datapath_indatatrf_1
    );
NAND_963: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_1,
        B => S1688,
        Y => S1792
    );
NAND_964: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_65,
        B => S1689,
        Y => S1793
    );
NAND_965: ENTITY WORK.NAND
    PORT MAP (
        A => S1792,
        B => S1793,
        Y => S5
    );
NOR_454: ENTITY WORK.NOR
    PORT MAP (
        A => S1116,
        B => S1389,
        Y => S1794
    );
NAND_966: ENTITY WORK.NAND
    PORT MAP (
        A => controller_fib_2,
        B => S1409,
        Y => S1795
    );
NOT_215: ENTITY WORK.NOT
    PORT MAP (
        A => S1795,
        Y => S1796
    );
NOR_455: ENTITY WORK.NOR
    PORT MAP (
        A => S1794,
        B => S1796,
        Y => S1797
    );
NOT_216: ENTITY WORK.NOT
    PORT MAP (
        A => S1797,
        Y => S1798
    );
NAND_967: ENTITY WORK.NAND
    PORT MAP (
        A => S1417,
        B => S1798,
        Y => S1799
    );
NOR_456: ENTITY WORK.NOR
    PORT MAP (
        A => controller_outflag_2,
        B => S1462,
        Y => S1800
    );
NOT_217: ENTITY WORK.NOT
    PORT MAP (
        A => S1800,
        Y => S1801
    );
NAND_968: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_242,
        B => S1437,
        Y => S1802
    );
NAND_969: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_178,
        B => S1438,
        Y => S1803
    );
NAND_970: ENTITY WORK.NAND
    PORT MAP (
        A => S1802,
        B => S1803,
        Y => S1804
    );
NAND_971: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S1804,
        Y => S1805
    );
NAND_972: ENTITY WORK.NAND
    PORT MAP (
        A => S7805,
        B => S1437,
        Y => S1806
    );
NOR_457: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_162,
        B => S1437,
        Y => S1807
    );
NAND_973: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S1806,
        Y => S1808
    );
NOR_458: ENTITY WORK.NOR
    PORT MAP (
        A => S1807,
        B => S1808,
        Y => S1809
    );
NAND_974: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_146,
        B => S1438,
        Y => S1810
    );
NAND_975: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_210,
        B => S1437,
        Y => S1811
    );
NAND_976: ENTITY WORK.NAND
    PORT MAP (
        A => S1810,
        B => S1811,
        Y => S1812
    );
NAND_977: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S1812,
        Y => S1813
    );
NOR_459: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_130,
        B => S1437,
        Y => S1814
    );
NOR_460: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_194,
        B => S1438,
        Y => S1815
    );
NOR_461: ENTITY WORK.NOR
    PORT MAP (
        A => S1814,
        B => S1815,
        Y => S1816
    );
NAND_978: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S1816,
        Y => S1817
    );
NAND_979: ENTITY WORK.NAND
    PORT MAP (
        A => S1813,
        B => S1817,
        Y => S1818
    );
NOR_462: ENTITY WORK.NOR
    PORT MAP (
        A => S1443,
        B => S1818,
        Y => S1819
    );
NOR_463: ENTITY WORK.NOR
    PORT MAP (
        A => S1444,
        B => S1809,
        Y => S1820
    );
NAND_980: ENTITY WORK.NAND
    PORT MAP (
        A => S1805,
        B => S1820,
        Y => S1821
    );
NAND_981: ENTITY WORK.NAND
    PORT MAP (
        A => S1449,
        B => S1821,
        Y => S1822
    );
NOR_464: ENTITY WORK.NOR
    PORT MAP (
        A => S1819,
        B => S1822,
        Y => S1823
    );
NAND_982: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_98,
        B => S1458,
        Y => S1824
    );
NAND_983: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_114,
        B => S1457,
        Y => S1825
    );
NAND_984: ENTITY WORK.NAND
    PORT MAP (
        A => S1824,
        B => S1825,
        Y => S1826
    );
NAND_985: ENTITY WORK.NAND
    PORT MAP (
        A => S1437,
        B => S1826,
        Y => S1827
    );
NAND_986: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_34,
        B => S1458,
        Y => S1828
    );
NAND_987: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_50,
        B => S1457,
        Y => S1829
    );
NAND_988: ENTITY WORK.NAND
    PORT MAP (
        A => S1828,
        B => S1829,
        Y => S1830
    );
NAND_989: ENTITY WORK.NAND
    PORT MAP (
        A => S1438,
        B => S1830,
        Y => S1831
    );
NAND_990: ENTITY WORK.NAND
    PORT MAP (
        A => S1827,
        B => S1831,
        Y => S1832
    );
NAND_991: ENTITY WORK.NAND
    PORT MAP (
        A => S1487,
        B => S1832,
        Y => S1833
    );
NAND_992: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_82,
        B => S1498,
        Y => S1834
    );
NOR_465: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_66,
        B => S1438,
        Y => S1835
    );
NOT_218: ENTITY WORK.NOT
    PORT MAP (
        A => S1835,
        Y => S1836
    );
NAND_993: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_18,
        B => S1438,
        Y => S1837
    );
NAND_994: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S1837,
        Y => S1838
    );
NAND_995: ENTITY WORK.NAND
    PORT MAP (
        A => S1836,
        B => S1838,
        Y => S1839
    );
NAND_996: ENTITY WORK.NAND
    PORT MAP (
        A => S1834,
        B => S1839,
        Y => S1840
    );
NOT_219: ENTITY WORK.NOT
    PORT MAP (
        A => S1840,
        Y => S1841
    );
NOR_466: ENTITY WORK.NOR
    PORT MAP (
        A => S1452,
        B => S1841,
        Y => S1842
    );
NAND_997: ENTITY WORK.NAND
    PORT MAP (
        A => S1451,
        B => S1840,
        Y => S1843
    );
NAND_998: ENTITY WORK.NAND
    PORT MAP (
        A => S1833,
        B => S1843,
        Y => S1844
    );
NOR_467: ENTITY WORK.NOR
    PORT MAP (
        A => S1823,
        B => S1842,
        Y => S1845
    );
NOR_468: ENTITY WORK.NOR
    PORT MAP (
        A => S1823,
        B => S1844,
        Y => S1846
    );
NAND_999: ENTITY WORK.NAND
    PORT MAP (
        A => S1833,
        B => S1845,
        Y => S1847
    );
NOR_469: ENTITY WORK.NOR
    PORT MAP (
        A => S1800,
        B => S1846,
        Y => S1848
    );
NAND_1000: ENTITY WORK.NAND
    PORT MAP (
        A => S1801,
        B => S1847,
        Y => S1849
    );
NAND_1001: ENTITY WORK.NAND
    PORT MAP (
        A => S1429,
        B => S1848,
        Y => S1850
    );
NAND_1002: ENTITY WORK.NAND
    PORT MAP (
        A => S1799,
        B => S1850,
        Y => S1851
    );
NOT_220: ENTITY WORK.NOT
    PORT MAP (
        A => S1851,
        Y => S1852
    );
NOR_470: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_2,
        B => S1852,
        Y => S1853
    );
NOT_221: ENTITY WORK.NOT
    PORT MAP (
        A => S1853,
        Y => S1854
    );
NOR_471: ENTITY WORK.NOR
    PORT MAP (
        A => S1116,
        B => S1851,
        Y => S1855
    );
NOT_222: ENTITY WORK.NOT
    PORT MAP (
        A => S1855,
        Y => S1856
    );
NAND_1003: ENTITY WORK.NAND
    PORT MAP (
        A => S1854,
        B => S1856,
        Y => S1857
    );
NOR_472: ENTITY WORK.NOR
    PORT MAP (
        A => S1750,
        B => S1757,
        Y => S1858
    );
NOR_473: ENTITY WORK.NOR
    PORT MAP (
        A => S1857,
        B => S1858,
        Y => S1859
    );
NAND_1004: ENTITY WORK.NAND
    PORT MAP (
        A => S1857,
        B => S1858,
        Y => S1860
    );
NOT_223: ENTITY WORK.NOT
    PORT MAP (
        A => S1860,
        Y => S1861
    );
NOR_474: ENTITY WORK.NOR
    PORT MAP (
        A => S1859,
        B => S1861,
        Y => S1862
    );
NAND_1005: ENTITY WORK.NAND
    PORT MAP (
        A => S1525,
        B => S1862,
        Y => S1863
    );
NAND_1006: ENTITY WORK.NAND
    PORT MAP (
        A => S1761,
        B => S1788,
        Y => S1864
    );
NOR_475: ENTITY WORK.NOR
    PORT MAP (
        A => S1857,
        B => S1864,
        Y => S1865
    );
NAND_1007: ENTITY WORK.NAND
    PORT MAP (
        A => S1857,
        B => S1864,
        Y => S1866
    );
NAND_1008: ENTITY WORK.NAND
    PORT MAP (
        A => S1527,
        B => S1866,
        Y => S1867
    );
NOR_476: ENTITY WORK.NOR
    PORT MAP (
        A => S1865,
        B => S1867,
        Y => S1868
    );
NAND_1009: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_2,
        B => S1851,
        Y => S1869
    );
NOR_477: ENTITY WORK.NOR
    PORT MAP (
        A => S1533,
        B => S1869,
        Y => S1870
    );
NOR_478: ENTITY WORK.NOR
    PORT MAP (
        A => S1547,
        B => S1797,
        Y => S1871
    );
NAND_1010: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_shiftunit_2171_A,
        B => S1614,
        Y => S1872
    );
NAND_1011: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_shiftunit_2475_A,
        B => S1609,
        Y => S1873
    );
NAND_1012: ENTITY WORK.NAND
    PORT MAP (
        A => S7897,
        B => S1336,
        Y => S1874
    );
NAND_1013: ENTITY WORK.NAND
    PORT MAP (
        A => S1338,
        B => S1874,
        Y => S1875
    );
NOR_479: ENTITY WORK.NOR
    PORT MAP (
        A => S1623,
        B => S1875,
        Y => S1876
    );
NOR_480: ENTITY WORK.NOR
    PORT MAP (
        A => S8054,
        B => S8571,
        Y => S1877
    );
NOR_481: ENTITY WORK.NOR
    PORT MAP (
        A => S8011,
        B => S1378,
        Y => S1878
    );
NAND_1014: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_databusin_2,
        B => S1627,
        Y => S1879
    );
NOR_482: ENTITY WORK.NOR
    PORT MAP (
        A => S1876,
        B => S1878,
        Y => S1880
    );
NAND_1015: ENTITY WORK.NAND
    PORT MAP (
        A => S1879,
        B => S1880,
        Y => S1881
    );
NOR_483: ENTITY WORK.NOR
    PORT MAP (
        A => S1877,
        B => S1881,
        Y => S1882
    );
NAND_1016: ENTITY WORK.NAND
    PORT MAP (
        A => S1873,
        B => S1882,
        Y => S1883
    );
NOR_484: ENTITY WORK.NOR
    PORT MAP (
        A => S1871,
        B => S1883,
        Y => S1884
    );
NAND_1017: ENTITY WORK.NAND
    PORT MAP (
        A => S1872,
        B => S1884,
        Y => S1885
    );
NOR_485: ENTITY WORK.NOR
    PORT MAP (
        A => S1116,
        B => S1765,
        Y => S1886
    );
NOR_486: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_2,
        B => S1766,
        Y => S1887
    );
NOR_487: ENTITY WORK.NOR
    PORT MAP (
        A => S1886,
        B => S1887,
        Y => S1888
    );
NAND_1018: ENTITY WORK.NAND
    PORT MAP (
        A => S1538,
        B => S1888,
        Y => S1889
    );
NOR_488: ENTITY WORK.NOR
    PORT MAP (
        A => S1870,
        B => S1885,
        Y => S1890
    );
NAND_1019: ENTITY WORK.NAND
    PORT MAP (
        A => S1889,
        B => S1890,
        Y => S1891
    );
NOR_489: ENTITY WORK.NOR
    PORT MAP (
        A => S1868,
        B => S1891,
        Y => S1892
    );
NAND_1020: ENTITY WORK.NAND
    PORT MAP (
        A => S1863,
        B => S1892,
        Y => datapath_indatatrf_2
    );
NAND_1021: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_2,
        B => S1688,
        Y => S1893
    );
NAND_1022: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_66,
        B => S1689,
        Y => S1894
    );
NAND_1023: ENTITY WORK.NAND
    PORT MAP (
        A => S1893,
        B => S1894,
        Y => S6
    );
NAND_1024: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_3,
        B => S1388,
        Y => S1895
    );
NAND_1025: ENTITY WORK.NAND
    PORT MAP (
        A => controller_fib_3,
        B => S1409,
        Y => S1896
    );
NAND_1026: ENTITY WORK.NAND
    PORT MAP (
        A => S1895,
        B => S1896,
        Y => S1897
    );
NOT_224: ENTITY WORK.NOT
    PORT MAP (
        A => S1897,
        Y => S1898
    );
NAND_1027: ENTITY WORK.NAND
    PORT MAP (
        A => S1417,
        B => S1897,
        Y => S1899
    );
NOR_490: ENTITY WORK.NOR
    PORT MAP (
        A => controller_outflag_3,
        B => S1462,
        Y => S1900
    );
NOT_225: ENTITY WORK.NOT
    PORT MAP (
        A => S1900,
        Y => S1901
    );
NAND_1028: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_243,
        B => S1437,
        Y => S1902
    );
NAND_1029: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_179,
        B => S1438,
        Y => S1903
    );
NAND_1030: ENTITY WORK.NAND
    PORT MAP (
        A => S1902,
        B => S1903,
        Y => S1904
    );
NAND_1031: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S1904,
        Y => S1905
    );
NAND_1032: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_163,
        B => S1438,
        Y => S1906
    );
NAND_1033: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_227,
        B => S1437,
        Y => S1907
    );
NAND_1034: ENTITY WORK.NAND
    PORT MAP (
        A => S1906,
        B => S1907,
        Y => S1908
    );
NAND_1035: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S1908,
        Y => S1909
    );
NAND_1036: ENTITY WORK.NAND
    PORT MAP (
        A => S1905,
        B => S1909,
        Y => S1910
    );
NAND_1037: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_147,
        B => S1438,
        Y => S1911
    );
NAND_1038: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_211,
        B => S1437,
        Y => S1912
    );
NAND_1039: ENTITY WORK.NAND
    PORT MAP (
        A => S1911,
        B => S1912,
        Y => S1913
    );
NAND_1040: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S1913,
        Y => S1914
    );
NOR_491: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_131,
        B => S1437,
        Y => S1915
    );
NAND_1041: ENTITY WORK.NAND
    PORT MAP (
        A => S7695,
        B => S1437,
        Y => S1916
    );
NAND_1042: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S1916,
        Y => S1917
    );
NOR_492: ENTITY WORK.NOR
    PORT MAP (
        A => S1915,
        B => S1917,
        Y => S1918
    );
NOR_493: ENTITY WORK.NOR
    PORT MAP (
        A => S1444,
        B => S1910,
        Y => S1919
    );
NOR_494: ENTITY WORK.NOR
    PORT MAP (
        A => S1443,
        B => S1918,
        Y => S1920
    );
NAND_1043: ENTITY WORK.NAND
    PORT MAP (
        A => S1914,
        B => S1920,
        Y => S1921
    );
NAND_1044: ENTITY WORK.NAND
    PORT MAP (
        A => S1449,
        B => S1921,
        Y => S1922
    );
NOR_495: ENTITY WORK.NOR
    PORT MAP (
        A => S1919,
        B => S1922,
        Y => S1923
    );
NAND_1045: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_67,
        B => S1459,
        Y => S1924
    );
NOT_226: ENTITY WORK.NOT
    PORT MAP (
        A => S1924,
        Y => S1925
    );
NOR_496: ENTITY WORK.NOR
    PORT MAP (
        A => S1452,
        B => S1458,
        Y => S1926
    );
NAND_1046: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_19,
        B => S1438,
        Y => S1927
    );
NAND_1047: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_83,
        B => S1437,
        Y => S1928
    );
NAND_1048: ENTITY WORK.NAND
    PORT MAP (
        A => S1927,
        B => S1928,
        Y => S1929
    );
NAND_1049: ENTITY WORK.NAND
    PORT MAP (
        A => S1926,
        B => S1929,
        Y => S1930
    );
NAND_1050: ENTITY WORK.NAND
    PORT MAP (
        A => S1462,
        B => S1930,
        Y => S1931
    );
NOR_497: ENTITY WORK.NOR
    PORT MAP (
        A => S1925,
        B => S1931,
        Y => S1932
    );
NAND_1051: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_115,
        B => S1437,
        Y => S1933
    );
NAND_1052: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_51,
        B => S1438,
        Y => S1934
    );
NAND_1053: ENTITY WORK.NAND
    PORT MAP (
        A => S1933,
        B => S1934,
        Y => S1935
    );
NAND_1054: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S1935,
        Y => S1936
    );
NAND_1055: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_99,
        B => S1437,
        Y => S1937
    );
NAND_1056: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_35,
        B => S1438,
        Y => S1938
    );
NAND_1057: ENTITY WORK.NAND
    PORT MAP (
        A => S1937,
        B => S1938,
        Y => S1939
    );
NOT_227: ENTITY WORK.NOT
    PORT MAP (
        A => S1939,
        Y => S1940
    );
NAND_1058: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S1939,
        Y => S1941
    );
NAND_1059: ENTITY WORK.NAND
    PORT MAP (
        A => S1936,
        B => S1941,
        Y => S1942
    );
NOR_498: ENTITY WORK.NOR
    PORT MAP (
        A => S1458,
        B => S1935,
        Y => S1943
    );
NAND_1060: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S1940,
        Y => S1944
    );
NAND_1061: ENTITY WORK.NAND
    PORT MAP (
        A => S1487,
        B => S1944,
        Y => S1945
    );
NOR_499: ENTITY WORK.NOR
    PORT MAP (
        A => S1943,
        B => S1945,
        Y => S1946
    );
NAND_1062: ENTITY WORK.NAND
    PORT MAP (
        A => S1487,
        B => S1942,
        Y => S1947
    );
NAND_1063: ENTITY WORK.NAND
    PORT MAP (
        A => S1932,
        B => S1947,
        Y => S1948
    );
NOR_500: ENTITY WORK.NOR
    PORT MAP (
        A => S1923,
        B => S1946,
        Y => S1949
    );
NOR_501: ENTITY WORK.NOR
    PORT MAP (
        A => S1923,
        B => S1948,
        Y => S1950
    );
NAND_1064: ENTITY WORK.NAND
    PORT MAP (
        A => S1932,
        B => S1949,
        Y => S1951
    );
NOR_502: ENTITY WORK.NOR
    PORT MAP (
        A => S1900,
        B => S1950,
        Y => S1952
    );
NAND_1065: ENTITY WORK.NAND
    PORT MAP (
        A => S1901,
        B => S1951,
        Y => S1953
    );
NAND_1066: ENTITY WORK.NAND
    PORT MAP (
        A => S1429,
        B => S1952,
        Y => S1954
    );
NAND_1067: ENTITY WORK.NAND
    PORT MAP (
        A => S1899,
        B => S1954,
        Y => S1955
    );
NOT_228: ENTITY WORK.NOT
    PORT MAP (
        A => S1955,
        Y => S1956
    );
NOR_503: ENTITY WORK.NOR
    PORT MAP (
        A => S1065,
        B => S1955,
        Y => S1957
    );
NOR_504: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_3,
        B => S1956,
        Y => S1958
    );
NOR_505: ENTITY WORK.NOR
    PORT MAP (
        A => S1065,
        B => S1956,
        Y => S1959
    );
NOT_229: ENTITY WORK.NOT
    PORT MAP (
        A => S1959,
        Y => S1960
    );
NOR_506: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_3,
        B => S1955,
        Y => S1961
    );
NOR_507: ENTITY WORK.NOR
    PORT MAP (
        A => S1959,
        B => S1961,
        Y => S1962
    );
NAND_1068: ENTITY WORK.NAND
    PORT MAP (
        A => S1866,
        B => S1869,
        Y => S1963
    );
NOR_508: ENTITY WORK.NOR
    PORT MAP (
        A => S1962,
        B => S1963,
        Y => S1964
    );
NAND_1069: ENTITY WORK.NAND
    PORT MAP (
        A => S1962,
        B => S1963,
        Y => S1965
    );
NOR_509: ENTITY WORK.NOR
    PORT MAP (
        A => S1528,
        B => S1964,
        Y => S1966
    );
NAND_1070: ENTITY WORK.NAND
    PORT MAP (
        A => S1965,
        B => S1966,
        Y => S1967
    );
NOR_510: ENTITY WORK.NOR
    PORT MAP (
        A => S1855,
        B => S1859,
        Y => S1968
    );
NOR_511: ENTITY WORK.NOR
    PORT MAP (
        A => S1962,
        B => S1968,
        Y => S1969
    );
NAND_1071: ENTITY WORK.NAND
    PORT MAP (
        A => S1962,
        B => S1968,
        Y => S1970
    );
NAND_1072: ENTITY WORK.NAND
    PORT MAP (
        A => S1525,
        B => S1970,
        Y => S1971
    );
NOR_512: ENTITY WORK.NOR
    PORT MAP (
        A => S1969,
        B => S1971,
        Y => S1972
    );
NOR_513: ENTITY WORK.NOR
    PORT MAP (
        A => S1533,
        B => S1960,
        Y => S1973
    );
NAND_1073: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_shiftunit_2189_A,
        B => S1614,
        Y => S1974
    );
NAND_1074: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_shiftunit_2493_A,
        B => S1609,
        Y => S1975
    );
NOR_514: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_muxmem_in2_3,
        B => S1337,
        Y => S1976
    );
NOR_515: ENTITY WORK.NOR
    PORT MAP (
        A => S1339,
        B => S1976,
        Y => S1977
    );
NOT_230: ENTITY WORK.NOT
    PORT MAP (
        A => S1977,
        Y => S1978
    );
NAND_1075: ENTITY WORK.NAND
    PORT MAP (
        A => S1622,
        B => S1977,
        Y => S1979
    );
NAND_1076: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu2_3,
        B => S8570,
        Y => S1980
    );
NAND_1077: ENTITY WORK.NAND
    PORT MAP (
        A => S1979,
        B => S1980,
        Y => S1981
    );
NAND_1078: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu1_3,
        B => S1377,
        Y => S1982
    );
NAND_1079: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_databusin_3,
        B => S1627,
        Y => S1983
    );
NAND_1080: ENTITY WORK.NAND
    PORT MAP (
        A => S1982,
        B => S1983,
        Y => S1984
    );
NOR_516: ENTITY WORK.NOR
    PORT MAP (
        A => S1981,
        B => S1984,
        Y => S1985
    );
NAND_1081: ENTITY WORK.NAND
    PORT MAP (
        A => S1975,
        B => S1985,
        Y => S1986
    );
NOR_517: ENTITY WORK.NOR
    PORT MAP (
        A => S1547,
        B => S1898,
        Y => S1987
    );
NOR_518: ENTITY WORK.NOR
    PORT MAP (
        A => S1986,
        B => S1987,
        Y => S1988
    );
NAND_1082: ENTITY WORK.NAND
    PORT MAP (
        A => S1974,
        B => S1988,
        Y => S1989
    );
NOR_519: ENTITY WORK.NOR
    PORT MAP (
        A => S1973,
        B => S1989,
        Y => S1990
    );
NOR_520: ENTITY WORK.NOR
    PORT MAP (
        A => S1065,
        B => S1887,
        Y => S1991
    );
NAND_1083: ENTITY WORK.NAND
    PORT MAP (
        A => S1065,
        B => S1887,
        Y => S1992
    );
NOR_521: ENTITY WORK.NOR
    PORT MAP (
        A => S1539,
        B => S1991,
        Y => S1993
    );
NAND_1084: ENTITY WORK.NAND
    PORT MAP (
        A => S1992,
        B => S1993,
        Y => S1994
    );
NAND_1085: ENTITY WORK.NAND
    PORT MAP (
        A => S1990,
        B => S1994,
        Y => S1995
    );
NOR_522: ENTITY WORK.NOR
    PORT MAP (
        A => S1972,
        B => S1995,
        Y => S1996
    );
NAND_1086: ENTITY WORK.NAND
    PORT MAP (
        A => S1967,
        B => S1996,
        Y => datapath_indatatrf_3
    );
NAND_1087: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_3,
        B => S1688,
        Y => S1997
    );
NAND_1088: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_67,
        B => S1689,
        Y => S1998
    );
NAND_1089: ENTITY WORK.NAND
    PORT MAP (
        A => S1997,
        B => S1998,
        Y => S7
    );
NAND_1090: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_4,
        B => S1388,
        Y => S1999
    );
NAND_1091: ENTITY WORK.NAND
    PORT MAP (
        A => controller_fib_4,
        B => S1409,
        Y => S2000
    );
NAND_1092: ENTITY WORK.NAND
    PORT MAP (
        A => S1999,
        B => S2000,
        Y => S2001
    );
NOT_231: ENTITY WORK.NOT
    PORT MAP (
        A => S2001,
        Y => S2002
    );
NAND_1093: ENTITY WORK.NAND
    PORT MAP (
        A => S1417,
        B => S2001,
        Y => S2003
    );
NAND_1094: ENTITY WORK.NAND
    PORT MAP (
        A => S1429,
        B => S1597,
        Y => S2004
    );
NAND_1095: ENTITY WORK.NAND
    PORT MAP (
        A => S2003,
        B => S2004,
        Y => S2005
    );
NOT_232: ENTITY WORK.NOT
    PORT MAP (
        A => S2005,
        Y => S2006
    );
NOR_523: ENTITY WORK.NOR
    PORT MAP (
        A => S1013,
        B => S2005,
        Y => S2007
    );
NOT_233: ENTITY WORK.NOT
    PORT MAP (
        A => S2007,
        Y => S2008
    );
NOR_524: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_4,
        B => S2006,
        Y => S2009
    );
NOT_234: ENTITY WORK.NOT
    PORT MAP (
        A => S2009,
        Y => S2010
    );
NAND_1096: ENTITY WORK.NAND
    PORT MAP (
        A => S2008,
        B => S2010,
        Y => S2011
    );
NOR_525: ENTITY WORK.NOR
    PORT MAP (
        A => S1957,
        B => S1969,
        Y => S2012
    );
NAND_1097: ENTITY WORK.NAND
    PORT MAP (
        A => S2011,
        B => S2012,
        Y => S2013
    );
NOR_526: ENTITY WORK.NOR
    PORT MAP (
        A => S2011,
        B => S2012,
        Y => S2014
    );
NAND_1098: ENTITY WORK.NAND
    PORT MAP (
        A => S1525,
        B => S2013,
        Y => S2015
    );
NOR_527: ENTITY WORK.NOR
    PORT MAP (
        A => S2014,
        B => S2015,
        Y => S2016
    );
NOR_528: ENTITY WORK.NOR
    PORT MAP (
        A => S1959,
        B => S1963,
        Y => S2017
    );
NOR_529: ENTITY WORK.NOR
    PORT MAP (
        A => S1961,
        B => S2017,
        Y => S2018
    );
NAND_1099: ENTITY WORK.NAND
    PORT MAP (
        A => S2011,
        B => S2018,
        Y => S2019
    );
NOR_530: ENTITY WORK.NOR
    PORT MAP (
        A => S2011,
        B => S2018,
        Y => S2020
    );
NOR_531: ENTITY WORK.NOR
    PORT MAP (
        A => S1528,
        B => S2020,
        Y => S2021
    );
NAND_1100: ENTITY WORK.NAND
    PORT MAP (
        A => S2019,
        B => S2021,
        Y => S2022
    );
NAND_1101: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_4,
        B => S2005,
        Y => S2023
    );
NOR_532: ENTITY WORK.NOR
    PORT MAP (
        A => S1533,
        B => S2023,
        Y => S2024
    );
NOR_533: ENTITY WORK.NOR
    PORT MAP (
        A => S1547,
        B => S2002,
        Y => S2025
    );
NAND_1102: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_shiftunit_2207_A,
        B => S1614,
        Y => S2026
    );
NAND_1103: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_shiftunit_2511_A,
        B => S1609,
        Y => S2027
    );
NAND_1104: ENTITY WORK.NAND
    PORT MAP (
        A => S7913,
        B => S1340,
        Y => S2028
    );
NAND_1105: ENTITY WORK.NAND
    PORT MAP (
        A => S1341,
        B => S2028,
        Y => S2029
    );
NOR_534: ENTITY WORK.NOR
    PORT MAP (
        A => S1623,
        B => S2029,
        Y => S2030
    );
NAND_1106: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_databusin_4,
        B => S1627,
        Y => S2031
    );
NAND_1107: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu2_4,
        B => S8570,
        Y => S2032
    );
NAND_1108: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu1_4,
        B => S1377,
        Y => S2033
    );
NAND_1109: ENTITY WORK.NAND
    PORT MAP (
        A => S2032,
        B => S2033,
        Y => S2034
    );
NAND_1110: ENTITY WORK.NAND
    PORT MAP (
        A => S2026,
        B => S2027,
        Y => S2035
    );
NOR_535: ENTITY WORK.NOR
    PORT MAP (
        A => S2025,
        B => S2035,
        Y => S2036
    );
NOR_536: ENTITY WORK.NOR
    PORT MAP (
        A => S2030,
        B => S2034,
        Y => S2037
    );
NAND_1111: ENTITY WORK.NAND
    PORT MAP (
        A => S2036,
        B => S2037,
        Y => S2038
    );
NOT_235: ENTITY WORK.NOT
    PORT MAP (
        A => S2038,
        Y => S2039
    );
NAND_1112: ENTITY WORK.NAND
    PORT MAP (
        A => S2031,
        B => S2039,
        Y => S2040
    );
NOR_537: ENTITY WORK.NOR
    PORT MAP (
        A => S2024,
        B => S2040,
        Y => S2041
    );
NAND_1113: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_4,
        B => S1992,
        Y => S2042
    );
NOR_538: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_4,
        B => S1992,
        Y => S2043
    );
NOR_539: ENTITY WORK.NOR
    PORT MAP (
        A => S1539,
        B => S2043,
        Y => S2044
    );
NAND_1114: ENTITY WORK.NAND
    PORT MAP (
        A => S2042,
        B => S2044,
        Y => S2045
    );
NAND_1115: ENTITY WORK.NAND
    PORT MAP (
        A => S2041,
        B => S2045,
        Y => S2046
    );
NOR_540: ENTITY WORK.NOR
    PORT MAP (
        A => S2016,
        B => S2046,
        Y => S2047
    );
NAND_1116: ENTITY WORK.NAND
    PORT MAP (
        A => S2022,
        B => S2047,
        Y => datapath_indatatrf_4
    );
NAND_1117: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_4,
        B => S1688,
        Y => S2048
    );
NAND_1118: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_68,
        B => S1689,
        Y => S2049
    );
NAND_1119: ENTITY WORK.NAND
    PORT MAP (
        A => S2048,
        B => S2049,
        Y => S8
    );
NOR_541: ENTITY WORK.NOR
    PORT MAP (
        A => S963,
        B => S1389,
        Y => S2050
    );
NAND_1120: ENTITY WORK.NAND
    PORT MAP (
        A => controller_216_B_0,
        B => S1401,
        Y => S2051
    );
NAND_1121: ENTITY WORK.NAND
    PORT MAP (
        A => controller_fib_4,
        B => S1406,
        Y => S2052
    );
NAND_1122: ENTITY WORK.NAND
    PORT MAP (
        A => S372,
        B => S2052,
        Y => S2053
    );
NOT_236: ENTITY WORK.NOT
    PORT MAP (
        A => S2053,
        Y => S2054
    );
NOR_542: ENTITY WORK.NOR
    PORT MAP (
        A => S2050,
        B => S2053,
        Y => S2055
    );
NAND_1123: ENTITY WORK.NAND
    PORT MAP (
        A => S2051,
        B => S2055,
        Y => S2056
    );
NAND_1124: ENTITY WORK.NAND
    PORT MAP (
        A => S1417,
        B => S2056,
        Y => S2057
    );
NOR_543: ENTITY WORK.NOR
    PORT MAP (
        A => controller_389_B_2,
        B => S1462,
        Y => S2058
    );
NOT_237: ENTITY WORK.NOT
    PORT MAP (
        A => S2058,
        Y => S2059
    );
NAND_1125: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_245,
        B => S1437,
        Y => S2060
    );
NAND_1126: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_181,
        B => S1438,
        Y => S2061
    );
NAND_1127: ENTITY WORK.NAND
    PORT MAP (
        A => S2060,
        B => S2061,
        Y => S2062
    );
NAND_1128: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S2062,
        Y => S2063
    );
NAND_1129: ENTITY WORK.NAND
    PORT MAP (
        A => S7822,
        B => S1437,
        Y => S2064
    );
NOR_544: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_165,
        B => S1437,
        Y => S2065
    );
NAND_1130: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S2064,
        Y => S2066
    );
NOR_545: ENTITY WORK.NOR
    PORT MAP (
        A => S2065,
        B => S2066,
        Y => S2067
    );
NAND_1131: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_149,
        B => S1438,
        Y => S2068
    );
NAND_1132: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_213,
        B => S1437,
        Y => S2069
    );
NAND_1133: ENTITY WORK.NAND
    PORT MAP (
        A => S2068,
        B => S2069,
        Y => S2070
    );
NAND_1134: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S2070,
        Y => S2071
    );
NOR_546: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_133,
        B => S1437,
        Y => S2072
    );
NOR_547: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_197,
        B => S1438,
        Y => S2073
    );
NOR_548: ENTITY WORK.NOR
    PORT MAP (
        A => S2072,
        B => S2073,
        Y => S2074
    );
NAND_1135: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S2074,
        Y => S2075
    );
NAND_1136: ENTITY WORK.NAND
    PORT MAP (
        A => S2071,
        B => S2075,
        Y => S2076
    );
NOR_549: ENTITY WORK.NOR
    PORT MAP (
        A => S1443,
        B => S2076,
        Y => S2077
    );
NOR_550: ENTITY WORK.NOR
    PORT MAP (
        A => S1444,
        B => S2067,
        Y => S2078
    );
NAND_1137: ENTITY WORK.NAND
    PORT MAP (
        A => S2063,
        B => S2078,
        Y => S2079
    );
NAND_1138: ENTITY WORK.NAND
    PORT MAP (
        A => S1449,
        B => S2079,
        Y => S2080
    );
NOR_551: ENTITY WORK.NOR
    PORT MAP (
        A => S2077,
        B => S2080,
        Y => S2081
    );
NAND_1139: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_101,
        B => S1458,
        Y => S2082
    );
NAND_1140: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_117,
        B => S1457,
        Y => S2083
    );
NAND_1141: ENTITY WORK.NAND
    PORT MAP (
        A => S2082,
        B => S2083,
        Y => S2084
    );
NAND_1142: ENTITY WORK.NAND
    PORT MAP (
        A => S1437,
        B => S2084,
        Y => S2085
    );
NAND_1143: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_37,
        B => S1458,
        Y => S2086
    );
NAND_1144: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_53,
        B => S1457,
        Y => S2087
    );
NAND_1145: ENTITY WORK.NAND
    PORT MAP (
        A => S2086,
        B => S2087,
        Y => S2088
    );
NAND_1146: ENTITY WORK.NAND
    PORT MAP (
        A => S1438,
        B => S2088,
        Y => S2089
    );
NAND_1147: ENTITY WORK.NAND
    PORT MAP (
        A => S2085,
        B => S2089,
        Y => S2090
    );
NAND_1148: ENTITY WORK.NAND
    PORT MAP (
        A => S1487,
        B => S2090,
        Y => S2091
    );
NAND_1149: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_85,
        B => S1498,
        Y => S2092
    );
NOR_552: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_69,
        B => S1438,
        Y => S2093
    );
NOT_238: ENTITY WORK.NOT
    PORT MAP (
        A => S2093,
        Y => S2094
    );
NAND_1150: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_21,
        B => S1438,
        Y => S2095
    );
NAND_1151: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S2095,
        Y => S2096
    );
NAND_1152: ENTITY WORK.NAND
    PORT MAP (
        A => S2094,
        B => S2096,
        Y => S2097
    );
NAND_1153: ENTITY WORK.NAND
    PORT MAP (
        A => S2092,
        B => S2097,
        Y => S2098
    );
NOT_239: ENTITY WORK.NOT
    PORT MAP (
        A => S2098,
        Y => S2099
    );
NOR_553: ENTITY WORK.NOR
    PORT MAP (
        A => S1452,
        B => S2099,
        Y => S2100
    );
NAND_1154: ENTITY WORK.NAND
    PORT MAP (
        A => S1451,
        B => S2098,
        Y => S2101
    );
NAND_1155: ENTITY WORK.NAND
    PORT MAP (
        A => S2091,
        B => S2101,
        Y => S2102
    );
NOR_554: ENTITY WORK.NOR
    PORT MAP (
        A => S2081,
        B => S2100,
        Y => S2103
    );
NOR_555: ENTITY WORK.NOR
    PORT MAP (
        A => S2081,
        B => S2102,
        Y => S2104
    );
NAND_1156: ENTITY WORK.NAND
    PORT MAP (
        A => S2091,
        B => S2103,
        Y => S2105
    );
NOR_556: ENTITY WORK.NOR
    PORT MAP (
        A => S2058,
        B => S2104,
        Y => S2106
    );
NAND_1157: ENTITY WORK.NAND
    PORT MAP (
        A => S2059,
        B => S2105,
        Y => S2107
    );
NAND_1158: ENTITY WORK.NAND
    PORT MAP (
        A => S1429,
        B => S2106,
        Y => S2108
    );
NAND_1159: ENTITY WORK.NAND
    PORT MAP (
        A => S2057,
        B => S2108,
        Y => S2109
    );
NOR_557: ENTITY WORK.NOR
    PORT MAP (
        A => S963,
        B => S2109,
        Y => S2110
    );
NOT_240: ENTITY WORK.NOT
    PORT MAP (
        A => S2110,
        Y => S2111
    );
NAND_1160: ENTITY WORK.NAND
    PORT MAP (
        A => S963,
        B => S2109,
        Y => S2112
    );
NAND_1161: ENTITY WORK.NAND
    PORT MAP (
        A => S2111,
        B => S2112,
        Y => S2113
    );
NOR_558: ENTITY WORK.NOR
    PORT MAP (
        A => S2007,
        B => S2014,
        Y => S2114
    );
NAND_1162: ENTITY WORK.NAND
    PORT MAP (
        A => S2113,
        B => S2114,
        Y => S2115
    );
NOR_559: ENTITY WORK.NOR
    PORT MAP (
        A => S2113,
        B => S2114,
        Y => S2116
    );
NAND_1163: ENTITY WORK.NAND
    PORT MAP (
        A => S1525,
        B => S2115,
        Y => S2117
    );
NOR_560: ENTITY WORK.NOR
    PORT MAP (
        A => S2116,
        B => S2117,
        Y => S2118
    );
NAND_1164: ENTITY WORK.NAND
    PORT MAP (
        A => S2019,
        B => S2023,
        Y => S2119
    );
NAND_1165: ENTITY WORK.NAND
    PORT MAP (
        A => S2113,
        B => S2119,
        Y => S2120
    );
NOR_561: ENTITY WORK.NOR
    PORT MAP (
        A => S2113,
        B => S2119,
        Y => S2121
    );
NOR_562: ENTITY WORK.NOR
    PORT MAP (
        A => S1528,
        B => S2121,
        Y => S2122
    );
NAND_1166: ENTITY WORK.NAND
    PORT MAP (
        A => S2120,
        B => S2122,
        Y => S2123
    );
NOR_563: ENTITY WORK.NOR
    PORT MAP (
        A => S963,
        B => S2043,
        Y => S2124
    );
NAND_1167: ENTITY WORK.NAND
    PORT MAP (
        A => S963,
        B => S2043,
        Y => S2125
    );
NOT_241: ENTITY WORK.NOT
    PORT MAP (
        A => S2125,
        Y => S2126
    );
NOR_564: ENTITY WORK.NOR
    PORT MAP (
        A => S2124,
        B => S2126,
        Y => S2127
    );
NAND_1168: ENTITY WORK.NAND
    PORT MAP (
        A => S1538,
        B => S2127,
        Y => S2128
    );
NAND_1169: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_5,
        B => S2109,
        Y => S2129
    );
NOR_565: ENTITY WORK.NOR
    PORT MAP (
        A => S1533,
        B => S2129,
        Y => S2130
    );
NAND_1170: ENTITY WORK.NAND
    PORT MAP (
        A => S1546,
        B => S2056,
        Y => S2131
    );
NAND_1171: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_shiftunit_2225_A,
        B => S1614,
        Y => S2132
    );
NOT_242: ENTITY WORK.NOT
    PORT MAP (
        A => S2132,
        Y => S2133
    );
NAND_1172: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_shiftunit_2529_A,
        B => S1609,
        Y => S2134
    );
NAND_1173: ENTITY WORK.NAND
    PORT MAP (
        A => S7920,
        B => S1341,
        Y => S2135
    );
NAND_1174: ENTITY WORK.NAND
    PORT MAP (
        A => S1344,
        B => S2135,
        Y => S2136
    );
NOR_566: ENTITY WORK.NOR
    PORT MAP (
        A => S1623,
        B => S2136,
        Y => S2137
    );
NOR_567: ENTITY WORK.NOR
    PORT MAP (
        A => S8236,
        B => S1628,
        Y => S2138
    );
NAND_1175: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu1_5,
        B => S1377,
        Y => S2139
    );
NOR_568: ENTITY WORK.NOR
    PORT MAP (
        A => S8087,
        B => S8571,
        Y => S2140
    );
NOR_569: ENTITY WORK.NOR
    PORT MAP (
        A => S2138,
        B => S2140,
        Y => S2141
    );
NAND_1176: ENTITY WORK.NAND
    PORT MAP (
        A => S2139,
        B => S2141,
        Y => S2142
    );
NOR_570: ENTITY WORK.NOR
    PORT MAP (
        A => S2137,
        B => S2142,
        Y => S2143
    );
NAND_1177: ENTITY WORK.NAND
    PORT MAP (
        A => S2134,
        B => S2143,
        Y => S2144
    );
NOR_571: ENTITY WORK.NOR
    PORT MAP (
        A => S2133,
        B => S2144,
        Y => S2145
    );
NAND_1178: ENTITY WORK.NAND
    PORT MAP (
        A => S2131,
        B => S2145,
        Y => S2146
    );
NOR_572: ENTITY WORK.NOR
    PORT MAP (
        A => S2130,
        B => S2146,
        Y => S2147
    );
NAND_1179: ENTITY WORK.NAND
    PORT MAP (
        A => S2128,
        B => S2147,
        Y => S2148
    );
NOR_573: ENTITY WORK.NOR
    PORT MAP (
        A => S2118,
        B => S2148,
        Y => S2149
    );
NAND_1180: ENTITY WORK.NAND
    PORT MAP (
        A => S2123,
        B => S2149,
        Y => datapath_indatatrf_5
    );
NAND_1181: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_5,
        B => S1688,
        Y => S2150
    );
NAND_1182: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_69,
        B => S1689,
        Y => S2151
    );
NAND_1183: ENTITY WORK.NAND
    PORT MAP (
        A => S2150,
        B => S2151,
        Y => S9
    );
NOR_574: ENTITY WORK.NOR
    PORT MAP (
        A => S910,
        B => S1389,
        Y => S2152
    );
NAND_1184: ENTITY WORK.NAND
    PORT MAP (
        A => controller_opcode_2,
        B => S1401,
        Y => S2153
    );
NAND_1185: ENTITY WORK.NAND
    PORT MAP (
        A => S2054,
        B => S2153,
        Y => S2154
    );
NOR_575: ENTITY WORK.NOR
    PORT MAP (
        A => S2152,
        B => S2154,
        Y => S2155
    );
NOR_576: ENTITY WORK.NOR
    PORT MAP (
        A => S1416,
        B => S2155,
        Y => S2156
    );
NOR_577: ENTITY WORK.NOR
    PORT MAP (
        A => controller_outflag_6,
        B => S1462,
        Y => S2157
    );
NOT_243: ENTITY WORK.NOT
    PORT MAP (
        A => S2157,
        Y => S2158
    );
NAND_1186: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_246,
        B => S1437,
        Y => S2159
    );
NAND_1187: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_182,
        B => S1438,
        Y => S2160
    );
NAND_1188: ENTITY WORK.NAND
    PORT MAP (
        A => S2159,
        B => S2160,
        Y => S2161
    );
NAND_1189: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S2161,
        Y => S2162
    );
NAND_1190: ENTITY WORK.NAND
    PORT MAP (
        A => S7823,
        B => S1437,
        Y => S2163
    );
NOR_578: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_166,
        B => S1437,
        Y => S2164
    );
NAND_1191: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S2163,
        Y => S2165
    );
NOR_579: ENTITY WORK.NOR
    PORT MAP (
        A => S2164,
        B => S2165,
        Y => S2166
    );
NAND_1192: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_150,
        B => S1438,
        Y => S2167
    );
NAND_1193: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_214,
        B => S1437,
        Y => S2168
    );
NAND_1194: ENTITY WORK.NAND
    PORT MAP (
        A => S2167,
        B => S2168,
        Y => S2169
    );
NAND_1195: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S2169,
        Y => S2170
    );
NOR_580: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_134,
        B => S1437,
        Y => S2171
    );
NOR_581: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_198,
        B => S1438,
        Y => S2172
    );
NOR_582: ENTITY WORK.NOR
    PORT MAP (
        A => S2171,
        B => S2172,
        Y => S2173
    );
NAND_1196: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S2173,
        Y => S2174
    );
NAND_1197: ENTITY WORK.NAND
    PORT MAP (
        A => S2170,
        B => S2174,
        Y => S2175
    );
NOR_583: ENTITY WORK.NOR
    PORT MAP (
        A => S1443,
        B => S2175,
        Y => S2176
    );
NOR_584: ENTITY WORK.NOR
    PORT MAP (
        A => S1444,
        B => S2166,
        Y => S2177
    );
NAND_1198: ENTITY WORK.NAND
    PORT MAP (
        A => S2162,
        B => S2177,
        Y => S2178
    );
NAND_1199: ENTITY WORK.NAND
    PORT MAP (
        A => S1449,
        B => S2178,
        Y => S2179
    );
NOR_585: ENTITY WORK.NOR
    PORT MAP (
        A => S2176,
        B => S2179,
        Y => S2180
    );
NAND_1200: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_102,
        B => S1458,
        Y => S2181
    );
NAND_1201: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_118,
        B => S1457,
        Y => S2182
    );
NAND_1202: ENTITY WORK.NAND
    PORT MAP (
        A => S2181,
        B => S2182,
        Y => S2183
    );
NAND_1203: ENTITY WORK.NAND
    PORT MAP (
        A => S1437,
        B => S2183,
        Y => S2184
    );
NAND_1204: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_38,
        B => S1458,
        Y => S2185
    );
NAND_1205: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_54,
        B => S1457,
        Y => S2186
    );
NAND_1206: ENTITY WORK.NAND
    PORT MAP (
        A => S2185,
        B => S2186,
        Y => S2187
    );
NAND_1207: ENTITY WORK.NAND
    PORT MAP (
        A => S1438,
        B => S2187,
        Y => S2188
    );
NAND_1208: ENTITY WORK.NAND
    PORT MAP (
        A => S2184,
        B => S2188,
        Y => S2189
    );
NAND_1209: ENTITY WORK.NAND
    PORT MAP (
        A => S1487,
        B => S2189,
        Y => S2190
    );
NAND_1210: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_86,
        B => S1498,
        Y => S2191
    );
NOR_586: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_70,
        B => S1438,
        Y => S2192
    );
NOT_244: ENTITY WORK.NOT
    PORT MAP (
        A => S2192,
        Y => S2193
    );
NAND_1211: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_22,
        B => S1438,
        Y => S2194
    );
NAND_1212: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S2194,
        Y => S2195
    );
NAND_1213: ENTITY WORK.NAND
    PORT MAP (
        A => S2193,
        B => S2195,
        Y => S2196
    );
NAND_1214: ENTITY WORK.NAND
    PORT MAP (
        A => S2191,
        B => S2196,
        Y => S2197
    );
NOT_245: ENTITY WORK.NOT
    PORT MAP (
        A => S2197,
        Y => S2198
    );
NOR_587: ENTITY WORK.NOR
    PORT MAP (
        A => S1452,
        B => S2198,
        Y => S2199
    );
NAND_1215: ENTITY WORK.NAND
    PORT MAP (
        A => S1451,
        B => S2197,
        Y => S2200
    );
NAND_1216: ENTITY WORK.NAND
    PORT MAP (
        A => S2190,
        B => S2200,
        Y => S2201
    );
NOR_588: ENTITY WORK.NOR
    PORT MAP (
        A => S2180,
        B => S2199,
        Y => S2202
    );
NOR_589: ENTITY WORK.NOR
    PORT MAP (
        A => S2180,
        B => S2201,
        Y => S2203
    );
NAND_1217: ENTITY WORK.NAND
    PORT MAP (
        A => S2190,
        B => S2202,
        Y => S2204
    );
NOR_590: ENTITY WORK.NOR
    PORT MAP (
        A => S2157,
        B => S2203,
        Y => S2205
    );
NAND_1218: ENTITY WORK.NAND
    PORT MAP (
        A => S2158,
        B => S2204,
        Y => S2206
    );
NOR_591: ENTITY WORK.NOR
    PORT MAP (
        A => S1430,
        B => S2206,
        Y => S2207
    );
NOR_592: ENTITY WORK.NOR
    PORT MAP (
        A => S2156,
        B => S2207,
        Y => S2208
    );
NOT_246: ENTITY WORK.NOT
    PORT MAP (
        A => S2208,
        Y => S2209
    );
NOR_593: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_6,
        B => S2208,
        Y => S2210
    );
NOT_247: ENTITY WORK.NOT
    PORT MAP (
        A => S2210,
        Y => S2211
    );
NOR_594: ENTITY WORK.NOR
    PORT MAP (
        A => S910,
        B => S2209,
        Y => S2212
    );
NOR_595: ENTITY WORK.NOR
    PORT MAP (
        A => S2210,
        B => S2212,
        Y => S2213
    );
NAND_1219: ENTITY WORK.NAND
    PORT MAP (
        A => S2111,
        B => S2114,
        Y => S2214
    );
NAND_1220: ENTITY WORK.NAND
    PORT MAP (
        A => S2112,
        B => S2214,
        Y => S2215
    );
NOT_248: ENTITY WORK.NOT
    PORT MAP (
        A => S2215,
        Y => S2216
    );
NOR_596: ENTITY WORK.NOR
    PORT MAP (
        A => S2213,
        B => S2216,
        Y => S2217
    );
NAND_1221: ENTITY WORK.NAND
    PORT MAP (
        A => S2213,
        B => S2216,
        Y => S2218
    );
NOT_249: ENTITY WORK.NOT
    PORT MAP (
        A => S2218,
        Y => S2219
    );
NAND_1222: ENTITY WORK.NAND
    PORT MAP (
        A => S1525,
        B => S2218,
        Y => S2220
    );
NOR_597: ENTITY WORK.NOR
    PORT MAP (
        A => S2217,
        B => S2220,
        Y => S2221
    );
NAND_1223: ENTITY WORK.NAND
    PORT MAP (
        A => S2120,
        B => S2129,
        Y => S2222
    );
NOT_250: ENTITY WORK.NOT
    PORT MAP (
        A => S2222,
        Y => S2223
    );
NAND_1224: ENTITY WORK.NAND
    PORT MAP (
        A => S2213,
        B => S2223,
        Y => S2224
    );
NOR_598: ENTITY WORK.NOR
    PORT MAP (
        A => S2213,
        B => S2223,
        Y => S2225
    );
NOR_599: ENTITY WORK.NOR
    PORT MAP (
        A => S1528,
        B => S2225,
        Y => S2226
    );
NAND_1225: ENTITY WORK.NAND
    PORT MAP (
        A => S2224,
        B => S2226,
        Y => S2227
    );
NOR_600: ENTITY WORK.NOR
    PORT MAP (
        A => S910,
        B => S2208,
        Y => S2228
    );
NOT_251: ENTITY WORK.NOT
    PORT MAP (
        A => S2228,
        Y => S2229
    );
NOR_601: ENTITY WORK.NOR
    PORT MAP (
        A => S1533,
        B => S2229,
        Y => S2230
    );
NOR_602: ENTITY WORK.NOR
    PORT MAP (
        A => S1547,
        B => S2155,
        Y => S2231
    );
NAND_1226: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_shiftunit_2243_A,
        B => S1614,
        Y => S2232
    );
NAND_1227: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_shiftunit_2547_A,
        B => S1609,
        Y => S2233
    );
NAND_1228: ENTITY WORK.NAND
    PORT MAP (
        A => S7928,
        B => S1344,
        Y => S2234
    );
NAND_1229: ENTITY WORK.NAND
    PORT MAP (
        A => S1346,
        B => S2234,
        Y => S2235
    );
NOR_603: ENTITY WORK.NOR
    PORT MAP (
        A => S1623,
        B => S2235,
        Y => S2236
    );
NAND_1230: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu2_6,
        B => S8570,
        Y => S2237
    );
NOR_604: ENTITY WORK.NOR
    PORT MAP (
        A => S8022,
        B => S1378,
        Y => S2238
    );
NOR_605: ENTITY WORK.NOR
    PORT MAP (
        A => S8257,
        B => S1628,
        Y => S2239
    );
NOR_606: ENTITY WORK.NOR
    PORT MAP (
        A => S2238,
        B => S2239,
        Y => S2240
    );
NAND_1231: ENTITY WORK.NAND
    PORT MAP (
        A => S2237,
        B => S2240,
        Y => S2241
    );
NOR_607: ENTITY WORK.NOR
    PORT MAP (
        A => S2236,
        B => S2241,
        Y => S2242
    );
NAND_1232: ENTITY WORK.NAND
    PORT MAP (
        A => S2232,
        B => S2233,
        Y => S2243
    );
NOR_608: ENTITY WORK.NOR
    PORT MAP (
        A => S2231,
        B => S2243,
        Y => S2244
    );
NAND_1233: ENTITY WORK.NAND
    PORT MAP (
        A => S2242,
        B => S2244,
        Y => S2245
    );
NOR_609: ENTITY WORK.NOR
    PORT MAP (
        A => S2230,
        B => S2245,
        Y => S2246
    );
NAND_1234: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_6,
        B => S2125,
        Y => S2247
    );
NOR_610: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_6,
        B => S2125,
        Y => S2248
    );
NOR_611: ENTITY WORK.NOR
    PORT MAP (
        A => S1539,
        B => S2248,
        Y => S2249
    );
NAND_1235: ENTITY WORK.NAND
    PORT MAP (
        A => S2247,
        B => S2249,
        Y => S2250
    );
NAND_1236: ENTITY WORK.NAND
    PORT MAP (
        A => S2246,
        B => S2250,
        Y => S2251
    );
NOR_612: ENTITY WORK.NOR
    PORT MAP (
        A => S2221,
        B => S2251,
        Y => S2252
    );
NAND_1237: ENTITY WORK.NAND
    PORT MAP (
        A => S2227,
        B => S2252,
        Y => datapath_indatatrf_6
    );
NAND_1238: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_6,
        B => S1688,
        Y => S2253
    );
NAND_1239: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_70,
        B => S1689,
        Y => S2254
    );
NAND_1240: ENTITY WORK.NAND
    PORT MAP (
        A => S2253,
        B => S2254,
        Y => S10
    );
NOR_613: ENTITY WORK.NOR
    PORT MAP (
        A => S858,
        B => S1389,
        Y => S2255
    );
NAND_1241: ENTITY WORK.NAND
    PORT MAP (
        A => controller_opcode_3,
        B => S1401,
        Y => S2256
    );
NOR_614: ENTITY WORK.NOR
    PORT MAP (
        A => S2053,
        B => S2255,
        Y => S2257
    );
NAND_1242: ENTITY WORK.NAND
    PORT MAP (
        A => S2256,
        B => S2257,
        Y => S2258
    );
NAND_1243: ENTITY WORK.NAND
    PORT MAP (
        A => S1417,
        B => S2258,
        Y => S2259
    );
NOR_615: ENTITY WORK.NOR
    PORT MAP (
        A => controller_outflag_7,
        B => S1462,
        Y => S2260
    );
NOT_252: ENTITY WORK.NOT
    PORT MAP (
        A => S2260,
        Y => S2261
    );
NAND_1244: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_247,
        B => S1437,
        Y => S2262
    );
NAND_1245: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_183,
        B => S1438,
        Y => S2263
    );
NAND_1246: ENTITY WORK.NAND
    PORT MAP (
        A => S2262,
        B => S2263,
        Y => S2264
    );
NAND_1247: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S2264,
        Y => S2265
    );
NAND_1248: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_167,
        B => S1438,
        Y => S2266
    );
NAND_1249: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_231,
        B => S1437,
        Y => S2267
    );
NAND_1250: ENTITY WORK.NAND
    PORT MAP (
        A => S2266,
        B => S2267,
        Y => S2268
    );
NAND_1251: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S2268,
        Y => S2269
    );
NAND_1252: ENTITY WORK.NAND
    PORT MAP (
        A => S2265,
        B => S2269,
        Y => S2270
    );
NAND_1253: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_151,
        B => S1438,
        Y => S2271
    );
NAND_1254: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_215,
        B => S1437,
        Y => S2272
    );
NAND_1255: ENTITY WORK.NAND
    PORT MAP (
        A => S2271,
        B => S2272,
        Y => S2273
    );
NAND_1256: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S2273,
        Y => S2274
    );
NOR_616: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_135,
        B => S1437,
        Y => S2275
    );
NAND_1257: ENTITY WORK.NAND
    PORT MAP (
        A => S7728,
        B => S1437,
        Y => S2276
    );
NAND_1258: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S2276,
        Y => S2277
    );
NOR_617: ENTITY WORK.NOR
    PORT MAP (
        A => S2275,
        B => S2277,
        Y => S2278
    );
NOR_618: ENTITY WORK.NOR
    PORT MAP (
        A => S1444,
        B => S2270,
        Y => S2279
    );
NOR_619: ENTITY WORK.NOR
    PORT MAP (
        A => S1443,
        B => S2278,
        Y => S2280
    );
NAND_1259: ENTITY WORK.NAND
    PORT MAP (
        A => S2274,
        B => S2280,
        Y => S2281
    );
NAND_1260: ENTITY WORK.NAND
    PORT MAP (
        A => S1449,
        B => S2281,
        Y => S2282
    );
NOR_620: ENTITY WORK.NOR
    PORT MAP (
        A => S2279,
        B => S2282,
        Y => S2283
    );
NAND_1261: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_71,
        B => S1459,
        Y => S2284
    );
NOT_253: ENTITY WORK.NOT
    PORT MAP (
        A => S2284,
        Y => S2285
    );
NAND_1262: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_23,
        B => S1438,
        Y => S2286
    );
NAND_1263: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_87,
        B => S1437,
        Y => S2287
    );
NAND_1264: ENTITY WORK.NAND
    PORT MAP (
        A => S2286,
        B => S2287,
        Y => S2288
    );
NAND_1265: ENTITY WORK.NAND
    PORT MAP (
        A => S1926,
        B => S2288,
        Y => S2289
    );
NAND_1266: ENTITY WORK.NAND
    PORT MAP (
        A => S1462,
        B => S2289,
        Y => S2290
    );
NOR_621: ENTITY WORK.NOR
    PORT MAP (
        A => S2285,
        B => S2290,
        Y => S2291
    );
NAND_1267: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_119,
        B => S1437,
        Y => S2292
    );
NAND_1268: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_55,
        B => S1438,
        Y => S2293
    );
NAND_1269: ENTITY WORK.NAND
    PORT MAP (
        A => S2292,
        B => S2293,
        Y => S2294
    );
NAND_1270: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S2294,
        Y => S2295
    );
NAND_1271: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_103,
        B => S1437,
        Y => S2296
    );
NAND_1272: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_39,
        B => S1438,
        Y => S2297
    );
NAND_1273: ENTITY WORK.NAND
    PORT MAP (
        A => S2296,
        B => S2297,
        Y => S2298
    );
NOT_254: ENTITY WORK.NOT
    PORT MAP (
        A => S2298,
        Y => S2299
    );
NAND_1274: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S2298,
        Y => S2300
    );
NAND_1275: ENTITY WORK.NAND
    PORT MAP (
        A => S2295,
        B => S2300,
        Y => S2301
    );
NOR_622: ENTITY WORK.NOR
    PORT MAP (
        A => S1458,
        B => S2294,
        Y => S2302
    );
NAND_1276: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S2299,
        Y => S2303
    );
NAND_1277: ENTITY WORK.NAND
    PORT MAP (
        A => S1487,
        B => S2303,
        Y => S2304
    );
NOR_623: ENTITY WORK.NOR
    PORT MAP (
        A => S2302,
        B => S2304,
        Y => S2305
    );
NAND_1278: ENTITY WORK.NAND
    PORT MAP (
        A => S1487,
        B => S2301,
        Y => S2306
    );
NAND_1279: ENTITY WORK.NAND
    PORT MAP (
        A => S2291,
        B => S2306,
        Y => S2307
    );
NOR_624: ENTITY WORK.NOR
    PORT MAP (
        A => S2283,
        B => S2305,
        Y => S2308
    );
NOR_625: ENTITY WORK.NOR
    PORT MAP (
        A => S2283,
        B => S2307,
        Y => S2309
    );
NAND_1280: ENTITY WORK.NAND
    PORT MAP (
        A => S2291,
        B => S2308,
        Y => S2310
    );
NOR_626: ENTITY WORK.NOR
    PORT MAP (
        A => S2260,
        B => S2309,
        Y => S2311
    );
NAND_1281: ENTITY WORK.NAND
    PORT MAP (
        A => S2261,
        B => S2310,
        Y => S2312
    );
NAND_1282: ENTITY WORK.NAND
    PORT MAP (
        A => S1429,
        B => S2311,
        Y => S2313
    );
NAND_1283: ENTITY WORK.NAND
    PORT MAP (
        A => S2259,
        B => S2313,
        Y => S2314
    );
NOT_255: ENTITY WORK.NOT
    PORT MAP (
        A => S2314,
        Y => S2315
    );
NOR_627: ENTITY WORK.NOR
    PORT MAP (
        A => S858,
        B => S2314,
        Y => S2316
    );
NAND_1284: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_7,
        B => S2315,
        Y => S2317
    );
NOR_628: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_7,
        B => S2315,
        Y => S2318
    );
NAND_1285: ENTITY WORK.NAND
    PORT MAP (
        A => S858,
        B => S2314,
        Y => S2319
    );
NAND_1286: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_7,
        B => S2314,
        Y => S2320
    );
NOR_629: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_7,
        B => S2314,
        Y => S2321
    );
NOR_630: ENTITY WORK.NOR
    PORT MAP (
        A => S2316,
        B => S2318,
        Y => S2322
    );
NOR_631: ENTITY WORK.NOR
    PORT MAP (
        A => S2225,
        B => S2228,
        Y => S2323
    );
NOR_632: ENTITY WORK.NOR
    PORT MAP (
        A => S2212,
        B => S2219,
        Y => S2324
    );
NOR_633: ENTITY WORK.NOR
    PORT MAP (
        A => S1533,
        B => S2320,
        Y => S2325
    );
NAND_1287: ENTITY WORK.NAND
    PORT MAP (
        A => S1546,
        B => S2258,
        Y => S2326
    );
NAND_1288: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_shiftunit_2261_A,
        B => S1614,
        Y => S2327
    );
NAND_1289: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_shiftunit_2565_A,
        B => S1609,
        Y => S2328
    );
NOT_256: ENTITY WORK.NOT
    PORT MAP (
        A => S2328,
        Y => S2329
    );
NAND_1290: ENTITY WORK.NAND
    PORT MAP (
        A => S7936,
        B => S1346,
        Y => S2330
    );
NAND_1291: ENTITY WORK.NAND
    PORT MAP (
        A => S1347,
        B => S2330,
        Y => S2331
    );
NOR_634: ENTITY WORK.NOR
    PORT MAP (
        A => S1623,
        B => S2331,
        Y => S2332
    );
NAND_1292: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu1_7,
        B => S1377,
        Y => S2333
    );
NAND_1293: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu2_7,
        B => S8570,
        Y => S2334
    );
NAND_1294: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_databusin_7,
        B => S1627,
        Y => S2335
    );
NAND_1295: ENTITY WORK.NAND
    PORT MAP (
        A => S2333,
        B => S2335,
        Y => S2336
    );
NOR_635: ENTITY WORK.NOR
    PORT MAP (
        A => S2332,
        B => S2336,
        Y => S2337
    );
NAND_1296: ENTITY WORK.NAND
    PORT MAP (
        A => S2334,
        B => S2337,
        Y => S2338
    );
NOR_636: ENTITY WORK.NOR
    PORT MAP (
        A => S2329,
        B => S2338,
        Y => S2339
    );
NOR_637: ENTITY WORK.NOR
    PORT MAP (
        A => S858,
        B => S2248,
        Y => S2340
    );
NAND_1297: ENTITY WORK.NAND
    PORT MAP (
        A => S858,
        B => S2248,
        Y => S2341
    );
NAND_1298: ENTITY WORK.NAND
    PORT MAP (
        A => S2326,
        B => S2339,
        Y => S2342
    );
NOR_638: ENTITY WORK.NOR
    PORT MAP (
        A => S2325,
        B => S2342,
        Y => S2343
    );
NOR_639: ENTITY WORK.NOR
    PORT MAP (
        A => S1539,
        B => S2340,
        Y => S2344
    );
NAND_1299: ENTITY WORK.NAND
    PORT MAP (
        A => S2341,
        B => S2344,
        Y => S2345
    );
NAND_1300: ENTITY WORK.NAND
    PORT MAP (
        A => S2327,
        B => S2345,
        Y => S2346
    );
NOT_257: ENTITY WORK.NOT
    PORT MAP (
        A => S2346,
        Y => S2347
    );
NAND_1301: ENTITY WORK.NAND
    PORT MAP (
        A => S2343,
        B => S2347,
        Y => S2348
    );
NOR_640: ENTITY WORK.NOR
    PORT MAP (
        A => S2322,
        B => S2324,
        Y => S2349
    );
NOT_258: ENTITY WORK.NOT
    PORT MAP (
        A => S2349,
        Y => S2350
    );
NAND_1302: ENTITY WORK.NAND
    PORT MAP (
        A => S2322,
        B => S2324,
        Y => S2351
    );
NAND_1303: ENTITY WORK.NAND
    PORT MAP (
        A => S2350,
        B => S2351,
        Y => S2352
    );
NAND_1304: ENTITY WORK.NAND
    PORT MAP (
        A => S1525,
        B => S2352,
        Y => S2353
    );
NOR_641: ENTITY WORK.NOR
    PORT MAP (
        A => S2322,
        B => S2323,
        Y => S2354
    );
NAND_1305: ENTITY WORK.NAND
    PORT MAP (
        A => S2322,
        B => S2323,
        Y => S2355
    );
NAND_1306: ENTITY WORK.NAND
    PORT MAP (
        A => S1527,
        B => S2355,
        Y => S2356
    );
NOR_642: ENTITY WORK.NOR
    PORT MAP (
        A => S2354,
        B => S2356,
        Y => S2357
    );
NOR_643: ENTITY WORK.NOR
    PORT MAP (
        A => S2348,
        B => S2357,
        Y => S2358
    );
NAND_1307: ENTITY WORK.NAND
    PORT MAP (
        A => S2353,
        B => S2358,
        Y => datapath_indatatrf_7
    );
NAND_1308: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_7,
        B => S1688,
        Y => S2359
    );
NAND_1309: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_71,
        B => S1689,
        Y => S2360
    );
NAND_1310: ENTITY WORK.NAND
    PORT MAP (
        A => S2359,
        B => S2360,
        Y => S11
    );
NOR_644: ENTITY WORK.NOR
    PORT MAP (
        A => controller_fib_0,
        B => S1396,
        Y => S2361
    );
NOR_645: ENTITY WORK.NOR
    PORT MAP (
        A => S1388,
        B => S1396,
        Y => S2362
    );
NOR_646: ENTITY WORK.NOR
    PORT MAP (
        A => S8309,
        B => S2362,
        Y => S2363
    );
NOR_647: ENTITY WORK.NOR
    PORT MAP (
        A => S1388,
        B => S2363,
        Y => S2364
    );
NOR_648: ENTITY WORK.NOR
    PORT MAP (
        A => S2361,
        B => S2364,
        Y => S2365
    );
NOR_649: ENTITY WORK.NOR
    PORT MAP (
        A => S2053,
        B => S2365,
        Y => S2366
    );
NOT_259: ENTITY WORK.NOT
    PORT MAP (
        A => S2366,
        Y => S2367
    );
NOR_650: ENTITY WORK.NOR
    PORT MAP (
        A => S1416,
        B => S2366,
        Y => S2368
    );
NAND_1311: ENTITY WORK.NAND
    PORT MAP (
        A => S1417,
        B => S2367,
        Y => S2369
    );
NAND_1312: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_248,
        B => S1437,
        Y => S2370
    );
NAND_1313: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_184,
        B => S1438,
        Y => S2371
    );
NAND_1314: ENTITY WORK.NAND
    PORT MAP (
        A => S2370,
        B => S2371,
        Y => S2372
    );
NAND_1315: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S2372,
        Y => S2373
    );
NAND_1316: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_168,
        B => S1438,
        Y => S2374
    );
NAND_1317: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_232,
        B => S1437,
        Y => S2375
    );
NAND_1318: ENTITY WORK.NAND
    PORT MAP (
        A => S2374,
        B => S2375,
        Y => S2376
    );
NAND_1319: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S2376,
        Y => S2377
    );
NAND_1320: ENTITY WORK.NAND
    PORT MAP (
        A => S2373,
        B => S2377,
        Y => S2378
    );
NAND_1321: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_152,
        B => S1438,
        Y => S2379
    );
NAND_1322: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_216,
        B => S1437,
        Y => S2380
    );
NAND_1323: ENTITY WORK.NAND
    PORT MAP (
        A => S2379,
        B => S2380,
        Y => S2381
    );
NAND_1324: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S2381,
        Y => S2382
    );
NOR_651: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_136,
        B => S1437,
        Y => S2383
    );
NAND_1325: ENTITY WORK.NAND
    PORT MAP (
        A => S7739,
        B => S1437,
        Y => S2384
    );
NAND_1326: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S2384,
        Y => S2385
    );
NOR_652: ENTITY WORK.NOR
    PORT MAP (
        A => S2383,
        B => S2385,
        Y => S2386
    );
NOR_653: ENTITY WORK.NOR
    PORT MAP (
        A => S1444,
        B => S2378,
        Y => S2387
    );
NOR_654: ENTITY WORK.NOR
    PORT MAP (
        A => S1443,
        B => S2386,
        Y => S2388
    );
NAND_1327: ENTITY WORK.NAND
    PORT MAP (
        A => S2382,
        B => S2388,
        Y => S2389
    );
NAND_1328: ENTITY WORK.NAND
    PORT MAP (
        A => S1449,
        B => S2389,
        Y => S2390
    );
NOR_655: ENTITY WORK.NOR
    PORT MAP (
        A => S2387,
        B => S2390,
        Y => S2391
    );
NAND_1329: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_104,
        B => S1458,
        Y => S2392
    );
NAND_1330: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_120,
        B => S1457,
        Y => S2393
    );
NAND_1331: ENTITY WORK.NAND
    PORT MAP (
        A => S2392,
        B => S2393,
        Y => S2394
    );
NAND_1332: ENTITY WORK.NAND
    PORT MAP (
        A => S1437,
        B => S2394,
        Y => S2395
    );
NAND_1333: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_40,
        B => S1458,
        Y => S2396
    );
NAND_1334: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_56,
        B => S1457,
        Y => S2397
    );
NAND_1335: ENTITY WORK.NAND
    PORT MAP (
        A => S2396,
        B => S2397,
        Y => S2398
    );
NAND_1336: ENTITY WORK.NAND
    PORT MAP (
        A => S1438,
        B => S2398,
        Y => S2399
    );
NAND_1337: ENTITY WORK.NAND
    PORT MAP (
        A => S2395,
        B => S2399,
        Y => S2400
    );
NAND_1338: ENTITY WORK.NAND
    PORT MAP (
        A => S1487,
        B => S2400,
        Y => S2401
    );
NOR_656: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_72,
        B => S1438,
        Y => S2402
    );
NOR_657: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_8,
        B => S1437,
        Y => S2403
    );
NOR_658: ENTITY WORK.NOR
    PORT MAP (
        A => S2402,
        B => S2403,
        Y => S2404
    );
NAND_1339: ENTITY WORK.NAND
    PORT MAP (
        A => S1459,
        B => S2404,
        Y => S2405
    );
NAND_1340: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_24,
        B => S1438,
        Y => S2406
    );
NAND_1341: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_88,
        B => S1437,
        Y => S2407
    );
NAND_1342: ENTITY WORK.NAND
    PORT MAP (
        A => S2406,
        B => S2407,
        Y => S2408
    );
NAND_1343: ENTITY WORK.NAND
    PORT MAP (
        A => S1926,
        B => S2408,
        Y => S2409
    );
NAND_1344: ENTITY WORK.NAND
    PORT MAP (
        A => S2405,
        B => S2409,
        Y => S2410
    );
NOT_260: ENTITY WORK.NOT
    PORT MAP (
        A => S2410,
        Y => S2411
    );
NAND_1345: ENTITY WORK.NAND
    PORT MAP (
        A => S2401,
        B => S2411,
        Y => S2412
    );
NAND_1346: ENTITY WORK.NAND
    PORT MAP (
        A => S2401,
        B => S2409,
        Y => S2413
    );
NOR_659: ENTITY WORK.NOR
    PORT MAP (
        A => S2391,
        B => S2413,
        Y => S2414
    );
NOR_660: ENTITY WORK.NOR
    PORT MAP (
        A => S2391,
        B => S2412,
        Y => S2415
    );
NAND_1347: ENTITY WORK.NAND
    PORT MAP (
        A => S2405,
        B => S2414,
        Y => S2416
    );
NOR_661: ENTITY WORK.NOR
    PORT MAP (
        A => S1461,
        B => S2415,
        Y => S2417
    );
NAND_1348: ENTITY WORK.NAND
    PORT MAP (
        A => S1462,
        B => S2416,
        Y => S2418
    );
NOR_662: ENTITY WORK.NOR
    PORT MAP (
        A => S1430,
        B => S2418,
        Y => S2419
    );
NOR_663: ENTITY WORK.NOR
    PORT MAP (
        A => S2368,
        B => S2419,
        Y => S2420
    );
NAND_1349: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_8,
        B => S2420,
        Y => S2421
    );
NOR_664: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_8,
        B => S2420,
        Y => S2422
    );
NOT_261: ENTITY WORK.NOT
    PORT MAP (
        A => S2422,
        Y => S2423
    );
NAND_1350: ENTITY WORK.NAND
    PORT MAP (
        A => S2421,
        B => S2423,
        Y => S2424
    );
NOT_262: ENTITY WORK.NOT
    PORT MAP (
        A => S2424,
        Y => S2425
    );
NOR_665: ENTITY WORK.NOR
    PORT MAP (
        A => S2321,
        B => S2323,
        Y => S2426
    );
NOT_263: ENTITY WORK.NOT
    PORT MAP (
        A => S2426,
        Y => S2427
    );
NAND_1351: ENTITY WORK.NAND
    PORT MAP (
        A => S2320,
        B => S2427,
        Y => S2428
    );
NOT_264: ENTITY WORK.NOT
    PORT MAP (
        A => S2428,
        Y => S2429
    );
NOR_666: ENTITY WORK.NOR
    PORT MAP (
        A => S2424,
        B => S2428,
        Y => S2430
    );
NOR_667: ENTITY WORK.NOR
    PORT MAP (
        A => S2425,
        B => S2429,
        Y => S2431
    );
NOR_668: ENTITY WORK.NOR
    PORT MAP (
        A => S2430,
        B => S2431,
        Y => S2432
    );
NAND_1352: ENTITY WORK.NAND
    PORT MAP (
        A => S1527,
        B => S2432,
        Y => S2433
    );
NOR_669: ENTITY WORK.NOR
    PORT MAP (
        A => S2318,
        B => S2324,
        Y => S2434
    );
NAND_1353: ENTITY WORK.NAND
    PORT MAP (
        A => S2213,
        B => S2322,
        Y => S2435
    );
NOR_670: ENTITY WORK.NOR
    PORT MAP (
        A => S2316,
        B => S2434,
        Y => S2436
    );
NOR_671: ENTITY WORK.NOR
    PORT MAP (
        A => S2424,
        B => S2436,
        Y => S2437
    );
NOT_265: ENTITY WORK.NOT
    PORT MAP (
        A => S2437,
        Y => S2438
    );
NAND_1354: ENTITY WORK.NAND
    PORT MAP (
        A => S2424,
        B => S2436,
        Y => S2439
    );
NAND_1355: ENTITY WORK.NAND
    PORT MAP (
        A => S1525,
        B => S2439,
        Y => S2440
    );
NOR_672: ENTITY WORK.NOR
    PORT MAP (
        A => S2437,
        B => S2440,
        Y => S2441
    );
NOR_673: ENTITY WORK.NOR
    PORT MAP (
        A => S805,
        B => S2420,
        Y => S2442
    );
NOT_266: ENTITY WORK.NOT
    PORT MAP (
        A => S2442,
        Y => S2443
    );
NOR_674: ENTITY WORK.NOR
    PORT MAP (
        A => S1533,
        B => S2443,
        Y => S2444
    );
NAND_1356: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_shiftunit_2279_A,
        B => S1614,
        Y => S2445
    );
NAND_1357: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_shiftunit_2583_A,
        B => S1609,
        Y => S2446
    );
NOR_675: ENTITY WORK.NOR
    PORT MAP (
        A => S1547,
        B => S2366,
        Y => S2447
    );
NAND_1358: ENTITY WORK.NAND
    PORT MAP (
        A => S7946,
        B => S1347,
        Y => S2448
    );
NAND_1359: ENTITY WORK.NAND
    PORT MAP (
        A => S1350,
        B => S2448,
        Y => S2449
    );
NOR_676: ENTITY WORK.NOR
    PORT MAP (
        A => S1623,
        B => S2449,
        Y => S2450
    );
NAND_1360: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_databusin_8,
        B => S1627,
        Y => S2451
    );
NAND_1361: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu1_8,
        B => S1377,
        Y => S2452
    );
NAND_1362: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu2_8,
        B => S8570,
        Y => S2453
    );
NAND_1363: ENTITY WORK.NAND
    PORT MAP (
        A => S2451,
        B => S2452,
        Y => S2454
    );
NOR_677: ENTITY WORK.NOR
    PORT MAP (
        A => S2447,
        B => S2454,
        Y => S2455
    );
NAND_1364: ENTITY WORK.NAND
    PORT MAP (
        A => S2453,
        B => S2455,
        Y => S2456
    );
NOR_678: ENTITY WORK.NOR
    PORT MAP (
        A => S2450,
        B => S2456,
        Y => S2457
    );
NAND_1365: ENTITY WORK.NAND
    PORT MAP (
        A => S2445,
        B => S2457,
        Y => S2458
    );
NOT_267: ENTITY WORK.NOT
    PORT MAP (
        A => S2458,
        Y => S2459
    );
NAND_1366: ENTITY WORK.NAND
    PORT MAP (
        A => S2446,
        B => S2459,
        Y => S2460
    );
NOR_679: ENTITY WORK.NOR
    PORT MAP (
        A => S2444,
        B => S2460,
        Y => S2461
    );
NAND_1367: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_8,
        B => S2341,
        Y => S2462
    );
NOR_680: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_8,
        B => S2341,
        Y => S2463
    );
NOT_268: ENTITY WORK.NOT
    PORT MAP (
        A => S2463,
        Y => S2464
    );
NOR_681: ENTITY WORK.NOR
    PORT MAP (
        A => S1539,
        B => S2463,
        Y => S2465
    );
NAND_1368: ENTITY WORK.NAND
    PORT MAP (
        A => S2462,
        B => S2465,
        Y => S2466
    );
NAND_1369: ENTITY WORK.NAND
    PORT MAP (
        A => S2461,
        B => S2466,
        Y => S2467
    );
NOR_682: ENTITY WORK.NOR
    PORT MAP (
        A => S2441,
        B => S2467,
        Y => S2468
    );
NAND_1370: ENTITY WORK.NAND
    PORT MAP (
        A => S2433,
        B => S2468,
        Y => datapath_indatatrf_8
    );
NAND_1371: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_8,
        B => S1688,
        Y => S2469
    );
NAND_1372: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_72,
        B => S1689,
        Y => S2470
    );
NAND_1373: ENTITY WORK.NAND
    PORT MAP (
        A => S2469,
        B => S2470,
        Y => S12
    );
NAND_1374: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_249,
        B => S1437,
        Y => S2471
    );
NAND_1375: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_185,
        B => S1438,
        Y => S2472
    );
NAND_1376: ENTITY WORK.NAND
    PORT MAP (
        A => S2471,
        B => S2472,
        Y => S2473
    );
NAND_1377: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S2473,
        Y => S2474
    );
NAND_1378: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_169,
        B => S1438,
        Y => S2475
    );
NAND_1379: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_233,
        B => S1437,
        Y => S2476
    );
NAND_1380: ENTITY WORK.NAND
    PORT MAP (
        A => S2475,
        B => S2476,
        Y => S2477
    );
NAND_1381: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S2477,
        Y => S2478
    );
NAND_1382: ENTITY WORK.NAND
    PORT MAP (
        A => S2474,
        B => S2478,
        Y => S2479
    );
NAND_1383: ENTITY WORK.NAND
    PORT MAP (
        A => S1443,
        B => S2479,
        Y => S2480
    );
NAND_1384: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_153,
        B => S1438,
        Y => S2481
    );
NAND_1385: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_217,
        B => S1437,
        Y => S2482
    );
NAND_1386: ENTITY WORK.NAND
    PORT MAP (
        A => S2481,
        B => S2482,
        Y => S2483
    );
NAND_1387: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S2483,
        Y => S2484
    );
NOR_683: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_137,
        B => S1437,
        Y => S2485
    );
NOR_684: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_201,
        B => S1438,
        Y => S2486
    );
NOR_685: ENTITY WORK.NOR
    PORT MAP (
        A => S2485,
        B => S2486,
        Y => S2487
    );
NAND_1388: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S2487,
        Y => S2488
    );
NAND_1389: ENTITY WORK.NAND
    PORT MAP (
        A => S2484,
        B => S2488,
        Y => S2489
    );
NAND_1390: ENTITY WORK.NAND
    PORT MAP (
        A => S1444,
        B => S2489,
        Y => S2490
    );
NAND_1391: ENTITY WORK.NAND
    PORT MAP (
        A => S2480,
        B => S2490,
        Y => S2491
    );
NAND_1392: ENTITY WORK.NAND
    PORT MAP (
        A => S1449,
        B => S2491,
        Y => S2492
    );
NAND_1393: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_25,
        B => S1438,
        Y => S2493
    );
NAND_1394: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_89,
        B => S1437,
        Y => S2494
    );
NAND_1395: ENTITY WORK.NAND
    PORT MAP (
        A => S2493,
        B => S2494,
        Y => S2495
    );
NAND_1396: ENTITY WORK.NAND
    PORT MAP (
        A => S1926,
        B => S2495,
        Y => S2496
    );
NAND_1397: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_9,
        B => S1438,
        Y => S2497
    );
NAND_1398: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_73,
        B => S1437,
        Y => S2498
    );
NAND_1399: ENTITY WORK.NAND
    PORT MAP (
        A => S2497,
        B => S2498,
        Y => S2499
    );
NAND_1400: ENTITY WORK.NAND
    PORT MAP (
        A => S1459,
        B => S2499,
        Y => S2500
    );
NAND_1401: ENTITY WORK.NAND
    PORT MAP (
        A => S2496,
        B => S2500,
        Y => S2501
    );
NAND_1402: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_57,
        B => S1438,
        Y => S2502
    );
NAND_1403: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_121,
        B => S1437,
        Y => S2503
    );
NAND_1404: ENTITY WORK.NAND
    PORT MAP (
        A => S2502,
        B => S2503,
        Y => S2504
    );
NOR_686: ENTITY WORK.NOR
    PORT MAP (
        A => S1458,
        B => S2504,
        Y => S2505
    );
NOR_687: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_41,
        B => S1437,
        Y => S2506
    );
NOR_688: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_105,
        B => S1438,
        Y => S2507
    );
NOR_689: ENTITY WORK.NOR
    PORT MAP (
        A => S2506,
        B => S2507,
        Y => S2508
    );
NOR_690: ENTITY WORK.NOR
    PORT MAP (
        A => S1457,
        B => S2508,
        Y => S2509
    );
NOR_691: ENTITY WORK.NOR
    PORT MAP (
        A => S2505,
        B => S2509,
        Y => S2510
    );
NAND_1405: ENTITY WORK.NAND
    PORT MAP (
        A => S1487,
        B => S2510,
        Y => S2511
    );
NOT_269: ENTITY WORK.NOT
    PORT MAP (
        A => S2511,
        Y => S2512
    );
NOR_692: ENTITY WORK.NOR
    PORT MAP (
        A => S2501,
        B => S2512,
        Y => S2513
    );
NAND_1406: ENTITY WORK.NAND
    PORT MAP (
        A => S2492,
        B => S2511,
        Y => S2514
    );
NOR_693: ENTITY WORK.NOR
    PORT MAP (
        A => S2501,
        B => S2514,
        Y => S2515
    );
NAND_1407: ENTITY WORK.NAND
    PORT MAP (
        A => S2492,
        B => S2513,
        Y => S2516
    );
NOR_694: ENTITY WORK.NOR
    PORT MAP (
        A => S1461,
        B => S2515,
        Y => S2517
    );
NAND_1408: ENTITY WORK.NAND
    PORT MAP (
        A => S1462,
        B => S2516,
        Y => S2518
    );
NOR_695: ENTITY WORK.NOR
    PORT MAP (
        A => S1430,
        B => S2518,
        Y => S2519
    );
NAND_1409: ENTITY WORK.NAND
    PORT MAP (
        A => S1429,
        B => S2517,
        Y => S2520
    );
NOR_696: ENTITY WORK.NOR
    PORT MAP (
        A => S2368,
        B => S2519,
        Y => S2521
    );
NAND_1410: ENTITY WORK.NAND
    PORT MAP (
        A => S2369,
        B => S2520,
        Y => S2522
    );
NOR_697: ENTITY WORK.NOR
    PORT MAP (
        A => S754,
        B => S2522,
        Y => S2523
    );
NOR_698: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_9,
        B => S2521,
        Y => S2524
    );
NOR_699: ENTITY WORK.NOR
    PORT MAP (
        A => S2523,
        B => S2524,
        Y => S2525
    );
NOT_270: ENTITY WORK.NOT
    PORT MAP (
        A => S2525,
        Y => S2526
    );
NAND_1411: ENTITY WORK.NAND
    PORT MAP (
        A => S2421,
        B => S2438,
        Y => S2527
    );
NOR_700: ENTITY WORK.NOR
    PORT MAP (
        A => S2525,
        B => S2527,
        Y => S2528
    );
NAND_1412: ENTITY WORK.NAND
    PORT MAP (
        A => S2525,
        B => S2527,
        Y => S2529
    );
NOR_701: ENTITY WORK.NOR
    PORT MAP (
        A => S1526,
        B => S2528,
        Y => S2530
    );
NAND_1413: ENTITY WORK.NAND
    PORT MAP (
        A => S2529,
        B => S2530,
        Y => S2531
    );
NAND_1414: ENTITY WORK.NAND
    PORT MAP (
        A => S2431,
        B => S2526,
        Y => S2532
    );
NOR_702: ENTITY WORK.NOR
    PORT MAP (
        A => S2431,
        B => S2442,
        Y => S2533
    );
NAND_1415: ENTITY WORK.NAND
    PORT MAP (
        A => S2525,
        B => S2533,
        Y => S2534
    );
NOR_703: ENTITY WORK.NOR
    PORT MAP (
        A => S2443,
        B => S2525,
        Y => S2535
    );
NOR_704: ENTITY WORK.NOR
    PORT MAP (
        A => S2525,
        B => S2533,
        Y => S2536
    );
NOR_705: ENTITY WORK.NOR
    PORT MAP (
        A => S1528,
        B => S2536,
        Y => S2537
    );
NAND_1416: ENTITY WORK.NAND
    PORT MAP (
        A => S2534,
        B => S2537,
        Y => S2538
    );
NAND_1417: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_9,
        B => S2464,
        Y => S2539
    );
NAND_1418: ENTITY WORK.NAND
    PORT MAP (
        A => S754,
        B => S2463,
        Y => S2540
    );
NOT_271: ENTITY WORK.NOT
    PORT MAP (
        A => S2540,
        Y => S2541
    );
NAND_1419: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_shiftunit_2297_A,
        B => S1614,
        Y => S2542
    );
NAND_1420: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_shiftunit_2601_A,
        B => S1609,
        Y => S2543
    );
NOT_272: ENTITY WORK.NOT
    PORT MAP (
        A => S2543,
        Y => S2544
    );
NOR_706: ENTITY WORK.NOR
    PORT MAP (
        A => controller_fib_1,
        B => S1396,
        Y => S2545
    );
NOR_707: ENTITY WORK.NOR
    PORT MAP (
        A => S2364,
        B => S2545,
        Y => S2546
    );
NOR_708: ENTITY WORK.NOR
    PORT MAP (
        A => S2053,
        B => S2546,
        Y => S2547
    );
NOR_709: ENTITY WORK.NOR
    PORT MAP (
        A => S1547,
        B => S2547,
        Y => S2548
    );
NOT_273: ENTITY WORK.NOT
    PORT MAP (
        A => S2548,
        Y => S2549
    );
NAND_1421: ENTITY WORK.NAND
    PORT MAP (
        A => S7957,
        B => S1350,
        Y => S2550
    );
NAND_1422: ENTITY WORK.NAND
    PORT MAP (
        A => S1352,
        B => S2550,
        Y => S2551
    );
NOR_710: ENTITY WORK.NOR
    PORT MAP (
        A => S1623,
        B => S2551,
        Y => S2552
    );
NOR_711: ENTITY WORK.NOR
    PORT MAP (
        A => S8129,
        B => S8571,
        Y => S2553
    );
NAND_1423: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu1_9,
        B => S1377,
        Y => S2554
    );
NOR_712: ENTITY WORK.NOR
    PORT MAP (
        A => S8288,
        B => S1628,
        Y => S2555
    );
NOR_713: ENTITY WORK.NOR
    PORT MAP (
        A => S2553,
        B => S2555,
        Y => S2556
    );
NAND_1424: ENTITY WORK.NAND
    PORT MAP (
        A => S2549,
        B => S2556,
        Y => S2557
    );
NOR_714: ENTITY WORK.NOR
    PORT MAP (
        A => S2552,
        B => S2557,
        Y => S2558
    );
NAND_1425: ENTITY WORK.NAND
    PORT MAP (
        A => S2554,
        B => S2558,
        Y => S2559
    );
NOR_715: ENTITY WORK.NOR
    PORT MAP (
        A => S2544,
        B => S2559,
        Y => S2560
    );
NAND_1426: ENTITY WORK.NAND
    PORT MAP (
        A => S2542,
        B => S2560,
        Y => S2561
    );
NAND_1427: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_9,
        B => S2522,
        Y => S2562
    );
NOR_716: ENTITY WORK.NOR
    PORT MAP (
        A => S1533,
        B => S2562,
        Y => S2563
    );
NAND_1428: ENTITY WORK.NAND
    PORT MAP (
        A => S2539,
        B => S2540,
        Y => S2564
    );
NOR_717: ENTITY WORK.NOR
    PORT MAP (
        A => S1539,
        B => S2564,
        Y => S2565
    );
NOR_718: ENTITY WORK.NOR
    PORT MAP (
        A => S2563,
        B => S2565,
        Y => S2566
    );
NAND_1429: ENTITY WORK.NAND
    PORT MAP (
        A => S2531,
        B => S2566,
        Y => S2567
    );
NOR_719: ENTITY WORK.NOR
    PORT MAP (
        A => S2561,
        B => S2567,
        Y => S2568
    );
NAND_1430: ENTITY WORK.NAND
    PORT MAP (
        A => S2538,
        B => S2568,
        Y => datapath_indatatrf_9
    );
NAND_1431: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_9,
        B => S1688,
        Y => S2569
    );
NAND_1432: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_73,
        B => S1689,
        Y => S2570
    );
NAND_1433: ENTITY WORK.NAND
    PORT MAP (
        A => S2569,
        B => S2570,
        Y => S13
    );
NAND_1434: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_250,
        B => S1443,
        Y => S2571
    );
NAND_1435: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_218,
        B => S1444,
        Y => S2572
    );
NAND_1436: ENTITY WORK.NAND
    PORT MAP (
        A => S2571,
        B => S2572,
        Y => S2573
    );
NAND_1437: ENTITY WORK.NAND
    PORT MAP (
        A => S1437,
        B => S2573,
        Y => S2574
    );
NAND_1438: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_186,
        B => S1443,
        Y => S2575
    );
NAND_1439: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_154,
        B => S1444,
        Y => S2576
    );
NAND_1440: ENTITY WORK.NAND
    PORT MAP (
        A => S2575,
        B => S2576,
        Y => S2577
    );
NAND_1441: ENTITY WORK.NAND
    PORT MAP (
        A => S1438,
        B => S2577,
        Y => S2578
    );
NAND_1442: ENTITY WORK.NAND
    PORT MAP (
        A => S2574,
        B => S2578,
        Y => S2579
    );
NAND_1443: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S2579,
        Y => S2580
    );
NAND_1444: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_234,
        B => S1443,
        Y => S2581
    );
NAND_1445: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_202,
        B => S1444,
        Y => S2582
    );
NAND_1446: ENTITY WORK.NAND
    PORT MAP (
        A => S2581,
        B => S2582,
        Y => S2583
    );
NAND_1447: ENTITY WORK.NAND
    PORT MAP (
        A => S1437,
        B => S2583,
        Y => S2584
    );
NAND_1448: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_170,
        B => S1443,
        Y => S2585
    );
NAND_1449: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_138,
        B => S1444,
        Y => S2586
    );
NAND_1450: ENTITY WORK.NAND
    PORT MAP (
        A => S2585,
        B => S2586,
        Y => S2587
    );
NAND_1451: ENTITY WORK.NAND
    PORT MAP (
        A => S1438,
        B => S2587,
        Y => S2588
    );
NAND_1452: ENTITY WORK.NAND
    PORT MAP (
        A => S2584,
        B => S2588,
        Y => S2589
    );
NAND_1453: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S2589,
        Y => S2590
    );
NAND_1454: ENTITY WORK.NAND
    PORT MAP (
        A => S2580,
        B => S2590,
        Y => S2591
    );
NAND_1455: ENTITY WORK.NAND
    PORT MAP (
        A => S1449,
        B => S2591,
        Y => S2592
    );
NOR_720: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_74,
        B => S1438,
        Y => S2593
    );
NOR_721: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_10,
        B => S1437,
        Y => S2594
    );
NOR_722: ENTITY WORK.NOR
    PORT MAP (
        A => S2593,
        B => S2594,
        Y => S2595
    );
NAND_1456: ENTITY WORK.NAND
    PORT MAP (
        A => S1459,
        B => S2595,
        Y => S2596
    );
NAND_1457: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_26,
        B => S1438,
        Y => S2597
    );
NAND_1458: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_90,
        B => S1437,
        Y => S2598
    );
NAND_1459: ENTITY WORK.NAND
    PORT MAP (
        A => S2597,
        B => S2598,
        Y => S2599
    );
NAND_1460: ENTITY WORK.NAND
    PORT MAP (
        A => S1926,
        B => S2599,
        Y => S2600
    );
NAND_1461: ENTITY WORK.NAND
    PORT MAP (
        A => S2596,
        B => S2600,
        Y => S2601
    );
NAND_1462: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_58,
        B => S1438,
        Y => S2602
    );
NAND_1463: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_122,
        B => S1437,
        Y => S2603
    );
NAND_1464: ENTITY WORK.NAND
    PORT MAP (
        A => S2602,
        B => S2603,
        Y => S2604
    );
NOR_723: ENTITY WORK.NOR
    PORT MAP (
        A => S1458,
        B => S2604,
        Y => S2605
    );
NOR_724: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_42,
        B => S1437,
        Y => S2606
    );
NOR_725: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_106,
        B => S1438,
        Y => S2607
    );
NOR_726: ENTITY WORK.NOR
    PORT MAP (
        A => S2606,
        B => S2607,
        Y => S2608
    );
NOR_727: ENTITY WORK.NOR
    PORT MAP (
        A => S1457,
        B => S2608,
        Y => S2609
    );
NOR_728: ENTITY WORK.NOR
    PORT MAP (
        A => S2605,
        B => S2609,
        Y => S2610
    );
NAND_1465: ENTITY WORK.NAND
    PORT MAP (
        A => S1487,
        B => S2610,
        Y => S2611
    );
NOT_274: ENTITY WORK.NOT
    PORT MAP (
        A => S2611,
        Y => S2612
    );
NOR_729: ENTITY WORK.NOR
    PORT MAP (
        A => S2601,
        B => S2612,
        Y => S2613
    );
NAND_1466: ENTITY WORK.NAND
    PORT MAP (
        A => S2592,
        B => S2611,
        Y => S2614
    );
NOR_730: ENTITY WORK.NOR
    PORT MAP (
        A => S2601,
        B => S2614,
        Y => S2615
    );
NAND_1467: ENTITY WORK.NAND
    PORT MAP (
        A => S2592,
        B => S2613,
        Y => S2616
    );
NOR_731: ENTITY WORK.NOR
    PORT MAP (
        A => S1461,
        B => S2615,
        Y => S2617
    );
NAND_1468: ENTITY WORK.NAND
    PORT MAP (
        A => S1462,
        B => S2616,
        Y => S2618
    );
NAND_1469: ENTITY WORK.NAND
    PORT MAP (
        A => S1429,
        B => S2617,
        Y => S2619
    );
NAND_1470: ENTITY WORK.NAND
    PORT MAP (
        A => S2369,
        B => S2619,
        Y => S2620
    );
NOT_275: ENTITY WORK.NOT
    PORT MAP (
        A => S2620,
        Y => S2621
    );
NAND_1471: ENTITY WORK.NAND
    PORT MAP (
        A => S702,
        B => S2620,
        Y => S2622
    );
NOT_276: ENTITY WORK.NOT
    PORT MAP (
        A => S2622,
        Y => S2623
    );
NAND_1472: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_10,
        B => S2621,
        Y => S2624
    );
NOT_277: ENTITY WORK.NOT
    PORT MAP (
        A => S2624,
        Y => S2625
    );
NOR_732: ENTITY WORK.NOR
    PORT MAP (
        A => S2623,
        B => S2625,
        Y => S2626
    );
NOR_733: ENTITY WORK.NOR
    PORT MAP (
        A => S2523,
        B => S2527,
        Y => S2627
    );
NOR_734: ENTITY WORK.NOR
    PORT MAP (
        A => S2524,
        B => S2627,
        Y => S2628
    );
NOR_735: ENTITY WORK.NOR
    PORT MAP (
        A => S2626,
        B => S2628,
        Y => S2629
    );
NAND_1473: ENTITY WORK.NAND
    PORT MAP (
        A => S2626,
        B => S2628,
        Y => S2630
    );
NOR_736: ENTITY WORK.NOR
    PORT MAP (
        A => S1526,
        B => S2629,
        Y => S2631
    );
NAND_1474: ENTITY WORK.NAND
    PORT MAP (
        A => S2630,
        B => S2631,
        Y => S2632
    );
NAND_1475: ENTITY WORK.NAND
    PORT MAP (
        A => S2532,
        B => S2562,
        Y => S2633
    );
NOR_737: ENTITY WORK.NOR
    PORT MAP (
        A => S2535,
        B => S2633,
        Y => S2634
    );
NOR_738: ENTITY WORK.NOR
    PORT MAP (
        A => S2626,
        B => S2634,
        Y => S2635
    );
NAND_1476: ENTITY WORK.NAND
    PORT MAP (
        A => S2626,
        B => S2634,
        Y => S2636
    );
NAND_1477: ENTITY WORK.NAND
    PORT MAP (
        A => S1527,
        B => S2636,
        Y => S2637
    );
NOR_739: ENTITY WORK.NOR
    PORT MAP (
        A => S2635,
        B => S2637,
        Y => S2638
    );
NAND_1478: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_10,
        B => S2620,
        Y => S2639
    );
NOT_278: ENTITY WORK.NOT
    PORT MAP (
        A => S2639,
        Y => S2640
    );
NOR_740: ENTITY WORK.NOR
    PORT MAP (
        A => S1533,
        B => S2639,
        Y => S2641
    );
NAND_1479: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_shiftunit_2315_A,
        B => S1614,
        Y => S2642
    );
NAND_1480: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_shiftunit_2619_A,
        B => S1609,
        Y => S2643
    );
NOT_279: ENTITY WORK.NOT
    PORT MAP (
        A => S2643,
        Y => S2644
    );
NAND_1481: ENTITY WORK.NAND
    PORT MAP (
        A => S7968,
        B => S1352,
        Y => S2645
    );
NAND_1482: ENTITY WORK.NAND
    PORT MAP (
        A => S1354,
        B => S2645,
        Y => S2646
    );
NOR_741: ENTITY WORK.NOR
    PORT MAP (
        A => S1623,
        B => S2646,
        Y => S2647
    );
NOR_742: ENTITY WORK.NOR
    PORT MAP (
        A => controller_fib_2,
        B => S1396,
        Y => S2648
    );
NOR_743: ENTITY WORK.NOR
    PORT MAP (
        A => S2364,
        B => S2648,
        Y => S2649
    );
NOR_744: ENTITY WORK.NOR
    PORT MAP (
        A => S2053,
        B => S2649,
        Y => S2650
    );
NOR_745: ENTITY WORK.NOR
    PORT MAP (
        A => S1547,
        B => S2650,
        Y => S2651
    );
NAND_1483: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu1_10,
        B => S1377,
        Y => S2652
    );
NAND_1484: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_databusin_10,
        B => S1627,
        Y => S2653
    );
NAND_1485: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu2_10,
        B => S8570,
        Y => S2654
    );
NOT_280: ENTITY WORK.NOT
    PORT MAP (
        A => S2654,
        Y => S2655
    );
NAND_1486: ENTITY WORK.NAND
    PORT MAP (
        A => S2652,
        B => S2653,
        Y => S2656
    );
NOR_746: ENTITY WORK.NOR
    PORT MAP (
        A => S2651,
        B => S2656,
        Y => S2657
    );
NOR_747: ENTITY WORK.NOR
    PORT MAP (
        A => S2647,
        B => S2655,
        Y => S2658
    );
NAND_1487: ENTITY WORK.NAND
    PORT MAP (
        A => S2657,
        B => S2658,
        Y => S2659
    );
NOR_748: ENTITY WORK.NOR
    PORT MAP (
        A => S2644,
        B => S2659,
        Y => S2660
    );
NAND_1488: ENTITY WORK.NAND
    PORT MAP (
        A => S2642,
        B => S2660,
        Y => S2661
    );
NOR_749: ENTITY WORK.NOR
    PORT MAP (
        A => S2641,
        B => S2661,
        Y => S2662
    );
NOR_750: ENTITY WORK.NOR
    PORT MAP (
        A => S702,
        B => S2541,
        Y => S2663
    );
NAND_1489: ENTITY WORK.NAND
    PORT MAP (
        A => S702,
        B => S2541,
        Y => S2664
    );
NOR_751: ENTITY WORK.NOR
    PORT MAP (
        A => S1539,
        B => S2663,
        Y => S2665
    );
NAND_1490: ENTITY WORK.NAND
    PORT MAP (
        A => S2664,
        B => S2665,
        Y => S2666
    );
NAND_1491: ENTITY WORK.NAND
    PORT MAP (
        A => S2662,
        B => S2666,
        Y => S2667
    );
NOR_752: ENTITY WORK.NOR
    PORT MAP (
        A => S2638,
        B => S2667,
        Y => S2668
    );
NAND_1492: ENTITY WORK.NAND
    PORT MAP (
        A => S2632,
        B => S2668,
        Y => datapath_indatatrf_10
    );
NAND_1493: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_10,
        B => S1688,
        Y => S2669
    );
NAND_1494: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_74,
        B => S1689,
        Y => S2670
    );
NAND_1495: ENTITY WORK.NAND
    PORT MAP (
        A => S2669,
        B => S2670,
        Y => S14
    );
NAND_1496: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_251,
        B => S1437,
        Y => S2671
    );
NAND_1497: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_187,
        B => S1438,
        Y => S2672
    );
NAND_1498: ENTITY WORK.NAND
    PORT MAP (
        A => S2671,
        B => S2672,
        Y => S2673
    );
NAND_1499: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S2673,
        Y => S2674
    );
NAND_1500: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_171,
        B => S1438,
        Y => S2675
    );
NAND_1501: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_235,
        B => S1437,
        Y => S2676
    );
NAND_1502: ENTITY WORK.NAND
    PORT MAP (
        A => S2675,
        B => S2676,
        Y => S2677
    );
NAND_1503: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S2677,
        Y => S2678
    );
NAND_1504: ENTITY WORK.NAND
    PORT MAP (
        A => S2674,
        B => S2678,
        Y => S2679
    );
NAND_1505: ENTITY WORK.NAND
    PORT MAP (
        A => S1443,
        B => S2679,
        Y => S2680
    );
NAND_1506: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_155,
        B => S1438,
        Y => S2681
    );
NAND_1507: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_219,
        B => S1437,
        Y => S2682
    );
NAND_1508: ENTITY WORK.NAND
    PORT MAP (
        A => S2681,
        B => S2682,
        Y => S2683
    );
NAND_1509: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S2683,
        Y => S2684
    );
NOR_753: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_139,
        B => S1437,
        Y => S2685
    );
NOR_754: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_203,
        B => S1438,
        Y => S2686
    );
NOR_755: ENTITY WORK.NOR
    PORT MAP (
        A => S2685,
        B => S2686,
        Y => S2687
    );
NAND_1510: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S2687,
        Y => S2688
    );
NAND_1511: ENTITY WORK.NAND
    PORT MAP (
        A => S2684,
        B => S2688,
        Y => S2689
    );
NAND_1512: ENTITY WORK.NAND
    PORT MAP (
        A => S1444,
        B => S2689,
        Y => S2690
    );
NAND_1513: ENTITY WORK.NAND
    PORT MAP (
        A => S2680,
        B => S2690,
        Y => S2691
    );
NAND_1514: ENTITY WORK.NAND
    PORT MAP (
        A => S1449,
        B => S2691,
        Y => S2692
    );
NAND_1515: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_27,
        B => S1438,
        Y => S2693
    );
NAND_1516: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_91,
        B => S1437,
        Y => S2694
    );
NAND_1517: ENTITY WORK.NAND
    PORT MAP (
        A => S2693,
        B => S2694,
        Y => S2695
    );
NAND_1518: ENTITY WORK.NAND
    PORT MAP (
        A => S1926,
        B => S2695,
        Y => S2696
    );
NAND_1519: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_11,
        B => S1438,
        Y => S2697
    );
NAND_1520: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_75,
        B => S1437,
        Y => S2698
    );
NAND_1521: ENTITY WORK.NAND
    PORT MAP (
        A => S2697,
        B => S2698,
        Y => S2699
    );
NAND_1522: ENTITY WORK.NAND
    PORT MAP (
        A => S1459,
        B => S2699,
        Y => S2700
    );
NAND_1523: ENTITY WORK.NAND
    PORT MAP (
        A => S2696,
        B => S2700,
        Y => S2701
    );
NAND_1524: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_123,
        B => S1437,
        Y => S2702
    );
NAND_1525: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_59,
        B => S1438,
        Y => S2703
    );
NAND_1526: ENTITY WORK.NAND
    PORT MAP (
        A => S2702,
        B => S2703,
        Y => S2704
    );
NAND_1527: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S2704,
        Y => S2705
    );
NAND_1528: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_107,
        B => S1437,
        Y => S2706
    );
NAND_1529: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_43,
        B => S1438,
        Y => S2707
    );
NAND_1530: ENTITY WORK.NAND
    PORT MAP (
        A => S2706,
        B => S2707,
        Y => S2708
    );
NAND_1531: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S2708,
        Y => S2709
    );
NAND_1532: ENTITY WORK.NAND
    PORT MAP (
        A => S2705,
        B => S2709,
        Y => S2710
    );
NAND_1533: ENTITY WORK.NAND
    PORT MAP (
        A => S1487,
        B => S2710,
        Y => S2711
    );
NOT_281: ENTITY WORK.NOT
    PORT MAP (
        A => S2711,
        Y => S2712
    );
NOR_756: ENTITY WORK.NOR
    PORT MAP (
        A => S2701,
        B => S2712,
        Y => S2713
    );
NAND_1534: ENTITY WORK.NAND
    PORT MAP (
        A => S2692,
        B => S2711,
        Y => S2714
    );
NOR_757: ENTITY WORK.NOR
    PORT MAP (
        A => S2701,
        B => S2714,
        Y => S2715
    );
NAND_1535: ENTITY WORK.NAND
    PORT MAP (
        A => S2692,
        B => S2713,
        Y => S2716
    );
NOR_758: ENTITY WORK.NOR
    PORT MAP (
        A => S1461,
        B => S2715,
        Y => S2717
    );
NAND_1536: ENTITY WORK.NAND
    PORT MAP (
        A => S1462,
        B => S2716,
        Y => S2718
    );
NAND_1537: ENTITY WORK.NAND
    PORT MAP (
        A => S1429,
        B => S2717,
        Y => S2719
    );
NAND_1538: ENTITY WORK.NAND
    PORT MAP (
        A => S2369,
        B => S2719,
        Y => S2720
    );
NOT_282: ENTITY WORK.NOT
    PORT MAP (
        A => S2720,
        Y => S2721
    );
NOR_759: ENTITY WORK.NOR
    PORT MAP (
        A => S651,
        B => S2720,
        Y => S2722
    );
NOR_760: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_11,
        B => S2721,
        Y => S2723
    );
NOR_761: ENTITY WORK.NOR
    PORT MAP (
        A => S2722,
        B => S2723,
        Y => S2724
    );
NOT_283: ENTITY WORK.NOT
    PORT MAP (
        A => S2724,
        Y => S2725
    );
NAND_1539: ENTITY WORK.NAND
    PORT MAP (
        A => S2624,
        B => S2630,
        Y => S2726
    );
NOR_762: ENTITY WORK.NOR
    PORT MAP (
        A => S2724,
        B => S2726,
        Y => S2727
    );
NAND_1540: ENTITY WORK.NAND
    PORT MAP (
        A => S2724,
        B => S2726,
        Y => S2728
    );
NAND_1541: ENTITY WORK.NAND
    PORT MAP (
        A => S1525,
        B => S2728,
        Y => S2729
    );
NOR_763: ENTITY WORK.NOR
    PORT MAP (
        A => S2727,
        B => S2729,
        Y => S2730
    );
NOR_764: ENTITY WORK.NOR
    PORT MAP (
        A => S2635,
        B => S2640,
        Y => S2731
    );
NAND_1542: ENTITY WORK.NAND
    PORT MAP (
        A => S2724,
        B => S2731,
        Y => S2732
    );
NOR_765: ENTITY WORK.NOR
    PORT MAP (
        A => S2724,
        B => S2731,
        Y => S2733
    );
NOR_766: ENTITY WORK.NOR
    PORT MAP (
        A => S1528,
        B => S2733,
        Y => S2734
    );
NAND_1543: ENTITY WORK.NAND
    PORT MAP (
        A => S2732,
        B => S2734,
        Y => S2735
    );
NAND_1544: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_11,
        B => S2664,
        Y => S2736
    );
NOR_767: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_11,
        B => S2664,
        Y => S2737
    );
NOR_768: ENTITY WORK.NOR
    PORT MAP (
        A => S1539,
        B => S2737,
        Y => S2738
    );
NAND_1545: ENTITY WORK.NAND
    PORT MAP (
        A => S2736,
        B => S2738,
        Y => S2739
    );
NAND_1546: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_11,
        B => S2720,
        Y => S2740
    );
NOR_769: ENTITY WORK.NOR
    PORT MAP (
        A => S1533,
        B => S2740,
        Y => S2741
    );
NAND_1547: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_shiftunit_2333_A,
        B => S1614,
        Y => S2742
    );
NAND_1548: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_shiftunit_2637_A,
        B => S1609,
        Y => S2743
    );
NOT_284: ENTITY WORK.NOT
    PORT MAP (
        A => S2743,
        Y => S2744
    );
NOR_770: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_muxmem_in2_11,
        B => S1353,
        Y => S2745
    );
NAND_1549: ENTITY WORK.NAND
    PORT MAP (
        A => S7978,
        B => S1354,
        Y => S2746
    );
NOR_771: ENTITY WORK.NOR
    PORT MAP (
        A => S1355,
        B => S2745,
        Y => S2747
    );
NAND_1550: ENTITY WORK.NAND
    PORT MAP (
        A => S1356,
        B => S2746,
        Y => S2748
    );
NAND_1551: ENTITY WORK.NAND
    PORT MAP (
        A => S1622,
        B => S2747,
        Y => S2749
    );
NOR_772: ENTITY WORK.NOR
    PORT MAP (
        A => controller_fib_3,
        B => S1396,
        Y => S2750
    );
NOR_773: ENTITY WORK.NOR
    PORT MAP (
        A => S2364,
        B => S2750,
        Y => S2751
    );
NOR_774: ENTITY WORK.NOR
    PORT MAP (
        A => S2053,
        B => S2751,
        Y => S2752
    );
NOR_775: ENTITY WORK.NOR
    PORT MAP (
        A => S1547,
        B => S2752,
        Y => S2753
    );
NAND_1552: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_databusin_11,
        B => S1627,
        Y => S2754
    );
NAND_1553: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu1_11,
        B => S1377,
        Y => S2755
    );
NAND_1554: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu2_11,
        B => S8570,
        Y => S2756
    );
NAND_1555: ENTITY WORK.NAND
    PORT MAP (
        A => S2755,
        B => S2756,
        Y => S2757
    );
NOT_285: ENTITY WORK.NOT
    PORT MAP (
        A => S2757,
        Y => S2758
    );
NAND_1556: ENTITY WORK.NAND
    PORT MAP (
        A => S2754,
        B => S2758,
        Y => S2759
    );
NOR_776: ENTITY WORK.NOR
    PORT MAP (
        A => S2753,
        B => S2759,
        Y => S2760
    );
NAND_1557: ENTITY WORK.NAND
    PORT MAP (
        A => S2749,
        B => S2760,
        Y => S2761
    );
NOR_777: ENTITY WORK.NOR
    PORT MAP (
        A => S2744,
        B => S2761,
        Y => S2762
    );
NAND_1558: ENTITY WORK.NAND
    PORT MAP (
        A => S2742,
        B => S2762,
        Y => S2763
    );
NOR_778: ENTITY WORK.NOR
    PORT MAP (
        A => S2741,
        B => S2763,
        Y => S2764
    );
NAND_1559: ENTITY WORK.NAND
    PORT MAP (
        A => S2739,
        B => S2764,
        Y => S2765
    );
NOR_779: ENTITY WORK.NOR
    PORT MAP (
        A => S2730,
        B => S2765,
        Y => S2766
    );
NAND_1560: ENTITY WORK.NAND
    PORT MAP (
        A => S2735,
        B => S2766,
        Y => datapath_indatatrf_11
    );
NAND_1561: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_11,
        B => S1688,
        Y => S2767
    );
NAND_1562: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_75,
        B => S1689,
        Y => S2768
    );
NAND_1563: ENTITY WORK.NAND
    PORT MAP (
        A => S2767,
        B => S2768,
        Y => S15
    );
NAND_1564: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_252,
        B => S1437,
        Y => S2769
    );
NAND_1565: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_188,
        B => S1438,
        Y => S2770
    );
NAND_1566: ENTITY WORK.NAND
    PORT MAP (
        A => S2769,
        B => S2770,
        Y => S2771
    );
NAND_1567: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S2771,
        Y => S2772
    );
NAND_1568: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_172,
        B => S1438,
        Y => S2773
    );
NAND_1569: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_236,
        B => S1437,
        Y => S2774
    );
NAND_1570: ENTITY WORK.NAND
    PORT MAP (
        A => S2773,
        B => S2774,
        Y => S2775
    );
NAND_1571: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S2775,
        Y => S2776
    );
NAND_1572: ENTITY WORK.NAND
    PORT MAP (
        A => S2772,
        B => S2776,
        Y => S2777
    );
NAND_1573: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_156,
        B => S1438,
        Y => S2778
    );
NAND_1574: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_220,
        B => S1437,
        Y => S2779
    );
NAND_1575: ENTITY WORK.NAND
    PORT MAP (
        A => S2778,
        B => S2779,
        Y => S2780
    );
NAND_1576: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S2780,
        Y => S2781
    );
NOR_780: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_140,
        B => S1437,
        Y => S2782
    );
NAND_1577: ENTITY WORK.NAND
    PORT MAP (
        A => S7750,
        B => S1437,
        Y => S2783
    );
NAND_1578: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S2783,
        Y => S2784
    );
NOR_781: ENTITY WORK.NOR
    PORT MAP (
        A => S2782,
        B => S2784,
        Y => S2785
    );
NOR_782: ENTITY WORK.NOR
    PORT MAP (
        A => S1444,
        B => S2777,
        Y => S2786
    );
NOR_783: ENTITY WORK.NOR
    PORT MAP (
        A => S1443,
        B => S2785,
        Y => S2787
    );
NAND_1579: ENTITY WORK.NAND
    PORT MAP (
        A => S2781,
        B => S2787,
        Y => S2788
    );
NAND_1580: ENTITY WORK.NAND
    PORT MAP (
        A => S1449,
        B => S2788,
        Y => S2789
    );
NOR_784: ENTITY WORK.NOR
    PORT MAP (
        A => S2786,
        B => S2789,
        Y => S2790
    );
NAND_1581: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_108,
        B => S1458,
        Y => S2791
    );
NAND_1582: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_124,
        B => S1457,
        Y => S2792
    );
NAND_1583: ENTITY WORK.NAND
    PORT MAP (
        A => S2791,
        B => S2792,
        Y => S2793
    );
NAND_1584: ENTITY WORK.NAND
    PORT MAP (
        A => S1437,
        B => S2793,
        Y => S2794
    );
NAND_1585: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_44,
        B => S1458,
        Y => S2795
    );
NAND_1586: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_60,
        B => S1457,
        Y => S2796
    );
NAND_1587: ENTITY WORK.NAND
    PORT MAP (
        A => S2795,
        B => S2796,
        Y => S2797
    );
NAND_1588: ENTITY WORK.NAND
    PORT MAP (
        A => S1438,
        B => S2797,
        Y => S2798
    );
NAND_1589: ENTITY WORK.NAND
    PORT MAP (
        A => S2794,
        B => S2798,
        Y => S2799
    );
NAND_1590: ENTITY WORK.NAND
    PORT MAP (
        A => S1487,
        B => S2799,
        Y => S2800
    );
NOR_785: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_76,
        B => S1438,
        Y => S2801
    );
NOR_786: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_12,
        B => S1437,
        Y => S2802
    );
NOR_787: ENTITY WORK.NOR
    PORT MAP (
        A => S2801,
        B => S2802,
        Y => S2803
    );
NAND_1591: ENTITY WORK.NAND
    PORT MAP (
        A => S1459,
        B => S2803,
        Y => S2804
    );
NAND_1592: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_28,
        B => S1438,
        Y => S2805
    );
NAND_1593: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_92,
        B => S1437,
        Y => S2806
    );
NAND_1594: ENTITY WORK.NAND
    PORT MAP (
        A => S2805,
        B => S2806,
        Y => S2807
    );
NAND_1595: ENTITY WORK.NAND
    PORT MAP (
        A => S1926,
        B => S2807,
        Y => S2808
    );
NAND_1596: ENTITY WORK.NAND
    PORT MAP (
        A => S2804,
        B => S2808,
        Y => S2809
    );
NOT_286: ENTITY WORK.NOT
    PORT MAP (
        A => S2809,
        Y => S2810
    );
NAND_1597: ENTITY WORK.NAND
    PORT MAP (
        A => S2800,
        B => S2810,
        Y => S2811
    );
NAND_1598: ENTITY WORK.NAND
    PORT MAP (
        A => S2800,
        B => S2808,
        Y => S2812
    );
NOR_788: ENTITY WORK.NOR
    PORT MAP (
        A => S2790,
        B => S2812,
        Y => S2813
    );
NOR_789: ENTITY WORK.NOR
    PORT MAP (
        A => S2790,
        B => S2811,
        Y => S2814
    );
NAND_1599: ENTITY WORK.NAND
    PORT MAP (
        A => S2804,
        B => S2813,
        Y => S2815
    );
NOR_790: ENTITY WORK.NOR
    PORT MAP (
        A => S1461,
        B => S2814,
        Y => S2816
    );
NAND_1600: ENTITY WORK.NAND
    PORT MAP (
        A => S1462,
        B => S2815,
        Y => S2817
    );
NAND_1601: ENTITY WORK.NAND
    PORT MAP (
        A => S1429,
        B => S2816,
        Y => S2818
    );
NAND_1602: ENTITY WORK.NAND
    PORT MAP (
        A => S2369,
        B => S2818,
        Y => S2819
    );
NOT_287: ENTITY WORK.NOT
    PORT MAP (
        A => S2819,
        Y => S2820
    );
NOR_791: ENTITY WORK.NOR
    PORT MAP (
        A => S599,
        B => S2819,
        Y => S2821
    );
NOT_288: ENTITY WORK.NOT
    PORT MAP (
        A => S2821,
        Y => S2822
    );
NOR_792: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_12,
        B => S2820,
        Y => S2823
    );
NOR_793: ENTITY WORK.NOR
    PORT MAP (
        A => S2821,
        B => S2823,
        Y => S2824
    );
NOR_794: ENTITY WORK.NOR
    PORT MAP (
        A => S2722,
        B => S2726,
        Y => S2825
    );
NOR_795: ENTITY WORK.NOR
    PORT MAP (
        A => S2723,
        B => S2825,
        Y => S2826
    );
NOR_796: ENTITY WORK.NOR
    PORT MAP (
        A => S2824,
        B => S2826,
        Y => S2827
    );
NAND_1603: ENTITY WORK.NAND
    PORT MAP (
        A => S2824,
        B => S2826,
        Y => S2828
    );
NAND_1604: ENTITY WORK.NAND
    PORT MAP (
        A => S1525,
        B => S2828,
        Y => S2829
    );
NOR_797: ENTITY WORK.NOR
    PORT MAP (
        A => S2827,
        B => S2829,
        Y => S2830
    );
NAND_1605: ENTITY WORK.NAND
    PORT MAP (
        A => S2635,
        B => S2725,
        Y => S2831
    );
NOR_798: ENTITY WORK.NOR
    PORT MAP (
        A => S2639,
        B => S2724,
        Y => S2832
    );
NAND_1606: ENTITY WORK.NAND
    PORT MAP (
        A => S2740,
        B => S2831,
        Y => S2833
    );
NOR_799: ENTITY WORK.NOR
    PORT MAP (
        A => S2832,
        B => S2833,
        Y => S2834
    );
NAND_1607: ENTITY WORK.NAND
    PORT MAP (
        A => S2824,
        B => S2834,
        Y => S2835
    );
NOR_800: ENTITY WORK.NOR
    PORT MAP (
        A => S2824,
        B => S2834,
        Y => S2836
    );
NOR_801: ENTITY WORK.NOR
    PORT MAP (
        A => S1528,
        B => S2836,
        Y => S2837
    );
NAND_1608: ENTITY WORK.NAND
    PORT MAP (
        A => S2835,
        B => S2837,
        Y => S2838
    );
NAND_1609: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_12,
        B => S2819,
        Y => S2839
    );
NOR_802: ENTITY WORK.NOR
    PORT MAP (
        A => S1533,
        B => S2839,
        Y => S2840
    );
NAND_1610: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_shiftunit_2351_A,
        B => S1614,
        Y => S2841
    );
NAND_1611: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_shiftunit_2655_A,
        B => S1609,
        Y => S2842
    );
NOT_289: ENTITY WORK.NOT
    PORT MAP (
        A => S2842,
        Y => S2843
    );
NOR_803: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_muxmem_in2_12,
        B => S1355,
        Y => S2844
    );
NAND_1612: ENTITY WORK.NAND
    PORT MAP (
        A => S7989,
        B => S1356,
        Y => S2845
    );
NOR_804: ENTITY WORK.NOR
    PORT MAP (
        A => S1357,
        B => S2844,
        Y => S2846
    );
NAND_1613: ENTITY WORK.NAND
    PORT MAP (
        A => S1358,
        B => S2845,
        Y => S2847
    );
NAND_1614: ENTITY WORK.NAND
    PORT MAP (
        A => S1622,
        B => S2846,
        Y => S2848
    );
NOR_805: ENTITY WORK.NOR
    PORT MAP (
        A => controller_fib_4,
        B => S1396,
        Y => S2849
    );
NOR_806: ENTITY WORK.NOR
    PORT MAP (
        A => S2364,
        B => S2849,
        Y => S2850
    );
NOR_807: ENTITY WORK.NOR
    PORT MAP (
        A => S2053,
        B => S2850,
        Y => S2851
    );
NOR_808: ENTITY WORK.NOR
    PORT MAP (
        A => S1547,
        B => S2851,
        Y => S2852
    );
NAND_1615: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_databusin_12,
        B => S1627,
        Y => S2853
    );
NAND_1616: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu1_12,
        B => S1377,
        Y => S2854
    );
NAND_1617: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu2_12,
        B => S8570,
        Y => S2855
    );
NAND_1618: ENTITY WORK.NAND
    PORT MAP (
        A => S2854,
        B => S2855,
        Y => S2856
    );
NOT_290: ENTITY WORK.NOT
    PORT MAP (
        A => S2856,
        Y => S2857
    );
NAND_1619: ENTITY WORK.NAND
    PORT MAP (
        A => S2853,
        B => S2857,
        Y => S2858
    );
NOR_809: ENTITY WORK.NOR
    PORT MAP (
        A => S2852,
        B => S2858,
        Y => S2859
    );
NAND_1620: ENTITY WORK.NAND
    PORT MAP (
        A => S2848,
        B => S2859,
        Y => S2860
    );
NOR_810: ENTITY WORK.NOR
    PORT MAP (
        A => S2843,
        B => S2860,
        Y => S2861
    );
NAND_1621: ENTITY WORK.NAND
    PORT MAP (
        A => S2841,
        B => S2861,
        Y => S2862
    );
NOR_811: ENTITY WORK.NOR
    PORT MAP (
        A => S2840,
        B => S2862,
        Y => S2863
    );
NAND_1622: ENTITY WORK.NAND
    PORT MAP (
        A => S599,
        B => S2737,
        Y => S2864
    );
NOR_812: ENTITY WORK.NOR
    PORT MAP (
        A => S599,
        B => S2737,
        Y => S2865
    );
NOR_813: ENTITY WORK.NOR
    PORT MAP (
        A => S1539,
        B => S2865,
        Y => S2866
    );
NAND_1623: ENTITY WORK.NAND
    PORT MAP (
        A => S2864,
        B => S2866,
        Y => S2867
    );
NAND_1624: ENTITY WORK.NAND
    PORT MAP (
        A => S2863,
        B => S2867,
        Y => S2868
    );
NOR_814: ENTITY WORK.NOR
    PORT MAP (
        A => S2830,
        B => S2868,
        Y => S2869
    );
NAND_1625: ENTITY WORK.NAND
    PORT MAP (
        A => S2838,
        B => S2869,
        Y => datapath_indatatrf_12
    );
NAND_1626: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_12,
        B => S1688,
        Y => S2870
    );
NAND_1627: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_76,
        B => S1689,
        Y => S2871
    );
NAND_1628: ENTITY WORK.NAND
    PORT MAP (
        A => S2870,
        B => S2871,
        Y => S16
    );
NAND_1629: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_253,
        B => S1437,
        Y => S2872
    );
NAND_1630: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_189,
        B => S1438,
        Y => S2873
    );
NAND_1631: ENTITY WORK.NAND
    PORT MAP (
        A => S2872,
        B => S2873,
        Y => S2874
    );
NAND_1632: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S2874,
        Y => S2875
    );
NAND_1633: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_173,
        B => S1438,
        Y => S2876
    );
NAND_1634: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_237,
        B => S1437,
        Y => S2877
    );
NAND_1635: ENTITY WORK.NAND
    PORT MAP (
        A => S2876,
        B => S2877,
        Y => S2878
    );
NAND_1636: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S2878,
        Y => S2879
    );
NAND_1637: ENTITY WORK.NAND
    PORT MAP (
        A => S2875,
        B => S2879,
        Y => S2880
    );
NAND_1638: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_157,
        B => S1438,
        Y => S2881
    );
NAND_1639: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_221,
        B => S1437,
        Y => S2882
    );
NAND_1640: ENTITY WORK.NAND
    PORT MAP (
        A => S2881,
        B => S2882,
        Y => S2883
    );
NAND_1641: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S2883,
        Y => S2884
    );
NOR_815: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_141,
        B => S1437,
        Y => S2885
    );
NAND_1642: ENTITY WORK.NAND
    PORT MAP (
        A => S7761,
        B => S1437,
        Y => S2886
    );
NAND_1643: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S2886,
        Y => S2887
    );
NOR_816: ENTITY WORK.NOR
    PORT MAP (
        A => S2885,
        B => S2887,
        Y => S2888
    );
NOR_817: ENTITY WORK.NOR
    PORT MAP (
        A => S1444,
        B => S2880,
        Y => S2889
    );
NOR_818: ENTITY WORK.NOR
    PORT MAP (
        A => S1443,
        B => S2888,
        Y => S2890
    );
NAND_1644: ENTITY WORK.NAND
    PORT MAP (
        A => S2884,
        B => S2890,
        Y => S2891
    );
NAND_1645: ENTITY WORK.NAND
    PORT MAP (
        A => S1449,
        B => S2891,
        Y => S2892
    );
NOR_819: ENTITY WORK.NOR
    PORT MAP (
        A => S2889,
        B => S2892,
        Y => S2893
    );
NAND_1646: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_109,
        B => S1458,
        Y => S2894
    );
NAND_1647: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_125,
        B => S1457,
        Y => S2895
    );
NAND_1648: ENTITY WORK.NAND
    PORT MAP (
        A => S2894,
        B => S2895,
        Y => S2896
    );
NAND_1649: ENTITY WORK.NAND
    PORT MAP (
        A => S1437,
        B => S2896,
        Y => S2897
    );
NAND_1650: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_45,
        B => S1458,
        Y => S2898
    );
NAND_1651: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_61,
        B => S1457,
        Y => S2899
    );
NAND_1652: ENTITY WORK.NAND
    PORT MAP (
        A => S2898,
        B => S2899,
        Y => S2900
    );
NAND_1653: ENTITY WORK.NAND
    PORT MAP (
        A => S1438,
        B => S2900,
        Y => S2901
    );
NAND_1654: ENTITY WORK.NAND
    PORT MAP (
        A => S2897,
        B => S2901,
        Y => S2902
    );
NAND_1655: ENTITY WORK.NAND
    PORT MAP (
        A => S1487,
        B => S2902,
        Y => S2903
    );
NOR_820: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_77,
        B => S1438,
        Y => S2904
    );
NOR_821: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_13,
        B => S1437,
        Y => S2905
    );
NOR_822: ENTITY WORK.NOR
    PORT MAP (
        A => S2904,
        B => S2905,
        Y => S2906
    );
NAND_1656: ENTITY WORK.NAND
    PORT MAP (
        A => S1459,
        B => S2906,
        Y => S2907
    );
NAND_1657: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_29,
        B => S1438,
        Y => S2908
    );
NAND_1658: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_93,
        B => S1437,
        Y => S2909
    );
NAND_1659: ENTITY WORK.NAND
    PORT MAP (
        A => S2908,
        B => S2909,
        Y => S2910
    );
NAND_1660: ENTITY WORK.NAND
    PORT MAP (
        A => S1926,
        B => S2910,
        Y => S2911
    );
NAND_1661: ENTITY WORK.NAND
    PORT MAP (
        A => S2907,
        B => S2911,
        Y => S2912
    );
NOT_291: ENTITY WORK.NOT
    PORT MAP (
        A => S2912,
        Y => S2913
    );
NAND_1662: ENTITY WORK.NAND
    PORT MAP (
        A => S2903,
        B => S2913,
        Y => S2914
    );
NAND_1663: ENTITY WORK.NAND
    PORT MAP (
        A => S2903,
        B => S2911,
        Y => S2915
    );
NOR_823: ENTITY WORK.NOR
    PORT MAP (
        A => S2893,
        B => S2915,
        Y => S2916
    );
NOR_824: ENTITY WORK.NOR
    PORT MAP (
        A => S2893,
        B => S2914,
        Y => S2917
    );
NAND_1664: ENTITY WORK.NAND
    PORT MAP (
        A => S2907,
        B => S2916,
        Y => S2918
    );
NOR_825: ENTITY WORK.NOR
    PORT MAP (
        A => S1461,
        B => S2917,
        Y => S2919
    );
NAND_1665: ENTITY WORK.NAND
    PORT MAP (
        A => S1462,
        B => S2918,
        Y => S2920
    );
NOR_826: ENTITY WORK.NOR
    PORT MAP (
        A => S1430,
        B => S2920,
        Y => S2921
    );
NOT_292: ENTITY WORK.NOT
    PORT MAP (
        A => S2921,
        Y => S2922
    );
NAND_1666: ENTITY WORK.NAND
    PORT MAP (
        A => S2369,
        B => S2922,
        Y => S2923
    );
NOT_293: ENTITY WORK.NOT
    PORT MAP (
        A => S2923,
        Y => S2924
    );
NOR_827: ENTITY WORK.NOR
    PORT MAP (
        A => S548,
        B => S2923,
        Y => S2925
    );
NOT_294: ENTITY WORK.NOT
    PORT MAP (
        A => S2925,
        Y => S2926
    );
NOR_828: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_13,
        B => S2924,
        Y => S2927
    );
NOT_295: ENTITY WORK.NOT
    PORT MAP (
        A => S2927,
        Y => S2928
    );
NAND_1667: ENTITY WORK.NAND
    PORT MAP (
        A => S2926,
        B => S2928,
        Y => S2929
    );
NOT_296: ENTITY WORK.NOT
    PORT MAP (
        A => S2929,
        Y => S2930
    );
NAND_1668: ENTITY WORK.NAND
    PORT MAP (
        A => S2822,
        B => S2828,
        Y => S2931
    );
NAND_1669: ENTITY WORK.NAND
    PORT MAP (
        A => S2929,
        B => S2931,
        Y => S2932
    );
NOR_829: ENTITY WORK.NOR
    PORT MAP (
        A => S2929,
        B => S2931,
        Y => S2933
    );
NOT_297: ENTITY WORK.NOT
    PORT MAP (
        A => S2933,
        Y => S2934
    );
NAND_1670: ENTITY WORK.NAND
    PORT MAP (
        A => S2932,
        B => S2934,
        Y => S2935
    );
NAND_1671: ENTITY WORK.NAND
    PORT MAP (
        A => S1525,
        B => S2935,
        Y => S2936
    );
NAND_1672: ENTITY WORK.NAND
    PORT MAP (
        A => S2839,
        B => S2930,
        Y => S2937
    );
NOR_830: ENTITY WORK.NOR
    PORT MAP (
        A => S2836,
        B => S2937,
        Y => S2938
    );
NAND_1673: ENTITY WORK.NAND
    PORT MAP (
        A => S2836,
        B => S2929,
        Y => S2939
    );
NOR_831: ENTITY WORK.NOR
    PORT MAP (
        A => S2839,
        B => S2930,
        Y => S2940
    );
NOR_832: ENTITY WORK.NOR
    PORT MAP (
        A => S1528,
        B => S2940,
        Y => S2941
    );
NAND_1674: ENTITY WORK.NAND
    PORT MAP (
        A => S2939,
        B => S2941,
        Y => S2942
    );
NOR_833: ENTITY WORK.NOR
    PORT MAP (
        A => S2938,
        B => S2942,
        Y => S2943
    );
NAND_1675: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_13,
        B => S2864,
        Y => S2944
    );
NOR_834: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_13,
        B => S2864,
        Y => S2945
    );
NOT_298: ENTITY WORK.NOT
    PORT MAP (
        A => S2945,
        Y => S2946
    );
NOR_835: ENTITY WORK.NOR
    PORT MAP (
        A => S1539,
        B => S2945,
        Y => S2947
    );
NAND_1676: ENTITY WORK.NAND
    PORT MAP (
        A => S2944,
        B => S2947,
        Y => S2948
    );
NAND_1677: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_13,
        B => S2923,
        Y => S2949
    );
NOR_836: ENTITY WORK.NOR
    PORT MAP (
        A => S1533,
        B => S2949,
        Y => S2950
    );
NAND_1678: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_shiftunit_2369_A,
        B => S1614,
        Y => S2951
    );
NAND_1679: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_shiftunit_2673_A,
        B => S1609,
        Y => S2952
    );
NOT_299: ENTITY WORK.NOT
    PORT MAP (
        A => S2952,
        Y => S2953
    );
NOR_837: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_muxmem_in2_13,
        B => S1357,
        Y => S2954
    );
NOR_838: ENTITY WORK.NOR
    PORT MAP (
        A => S1359,
        B => S2954,
        Y => S2955
    );
NOT_300: ENTITY WORK.NOT
    PORT MAP (
        A => S2955,
        Y => S2956
    );
NAND_1680: ENTITY WORK.NAND
    PORT MAP (
        A => S1622,
        B => S2955,
        Y => S2957
    );
NOR_839: ENTITY WORK.NOR
    PORT MAP (
        A => controller_216_B_0,
        B => S1396,
        Y => S2958
    );
NOR_840: ENTITY WORK.NOR
    PORT MAP (
        A => S2364,
        B => S2958,
        Y => S2959
    );
NOR_841: ENTITY WORK.NOR
    PORT MAP (
        A => S2053,
        B => S2959,
        Y => S2960
    );
NOR_842: ENTITY WORK.NOR
    PORT MAP (
        A => S1547,
        B => S2960,
        Y => S2961
    );
NAND_1681: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu1_13,
        B => S1377,
        Y => S2962
    );
NAND_1682: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu2_13,
        B => S8570,
        Y => S2963
    );
NAND_1683: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_databusin_13,
        B => S1627,
        Y => S2964
    );
NAND_1684: ENTITY WORK.NAND
    PORT MAP (
        A => S2963,
        B => S2964,
        Y => S2965
    );
NOT_301: ENTITY WORK.NOT
    PORT MAP (
        A => S2965,
        Y => S2966
    );
NAND_1685: ENTITY WORK.NAND
    PORT MAP (
        A => S2962,
        B => S2966,
        Y => S2967
    );
NOR_843: ENTITY WORK.NOR
    PORT MAP (
        A => S2961,
        B => S2967,
        Y => S2968
    );
NAND_1686: ENTITY WORK.NAND
    PORT MAP (
        A => S2957,
        B => S2968,
        Y => S2969
    );
NOR_844: ENTITY WORK.NOR
    PORT MAP (
        A => S2953,
        B => S2969,
        Y => S2970
    );
NAND_1687: ENTITY WORK.NAND
    PORT MAP (
        A => S2951,
        B => S2970,
        Y => S2971
    );
NOR_845: ENTITY WORK.NOR
    PORT MAP (
        A => S2950,
        B => S2971,
        Y => S2972
    );
NAND_1688: ENTITY WORK.NAND
    PORT MAP (
        A => S2948,
        B => S2972,
        Y => S2973
    );
NOR_846: ENTITY WORK.NOR
    PORT MAP (
        A => S2943,
        B => S2973,
        Y => S2974
    );
NAND_1689: ENTITY WORK.NAND
    PORT MAP (
        A => S2936,
        B => S2974,
        Y => datapath_indatatrf_13
    );
NAND_1690: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_13,
        B => S1688,
        Y => S2975
    );
NAND_1691: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_77,
        B => S1689,
        Y => S2976
    );
NAND_1692: ENTITY WORK.NAND
    PORT MAP (
        A => S2975,
        B => S2976,
        Y => S17
    );
NAND_1693: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_254,
        B => S1437,
        Y => S2977
    );
NAND_1694: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_190,
        B => S1438,
        Y => S2978
    );
NAND_1695: ENTITY WORK.NAND
    PORT MAP (
        A => S2977,
        B => S2978,
        Y => S2979
    );
NAND_1696: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S2979,
        Y => S2980
    );
NAND_1697: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_174,
        B => S1438,
        Y => S2981
    );
NAND_1698: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_238,
        B => S1437,
        Y => S2982
    );
NAND_1699: ENTITY WORK.NAND
    PORT MAP (
        A => S2981,
        B => S2982,
        Y => S2983
    );
NAND_1700: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S2983,
        Y => S2984
    );
NAND_1701: ENTITY WORK.NAND
    PORT MAP (
        A => S2980,
        B => S2984,
        Y => S2985
    );
NAND_1702: ENTITY WORK.NAND
    PORT MAP (
        A => S1443,
        B => S2985,
        Y => S2986
    );
NAND_1703: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_158,
        B => S1438,
        Y => S2987
    );
NAND_1704: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_222,
        B => S1437,
        Y => S2988
    );
NAND_1705: ENTITY WORK.NAND
    PORT MAP (
        A => S2987,
        B => S2988,
        Y => S2989
    );
NAND_1706: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S2989,
        Y => S2990
    );
NOR_847: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_142,
        B => S1437,
        Y => S2991
    );
NOR_848: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_206,
        B => S1438,
        Y => S2992
    );
NAND_1707: ENTITY WORK.NAND
    PORT MAP (
        A => S7772,
        B => S1437,
        Y => S2993
    );
NOR_849: ENTITY WORK.NOR
    PORT MAP (
        A => S2991,
        B => S2992,
        Y => S2994
    );
NAND_1708: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S2993,
        Y => S2995
    );
NOR_850: ENTITY WORK.NOR
    PORT MAP (
        A => S2991,
        B => S2995,
        Y => S2996
    );
NAND_1709: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S2994,
        Y => S2997
    );
NAND_1710: ENTITY WORK.NAND
    PORT MAP (
        A => S2990,
        B => S2997,
        Y => S2998
    );
NAND_1711: ENTITY WORK.NAND
    PORT MAP (
        A => S1444,
        B => S2998,
        Y => S2999
    );
NAND_1712: ENTITY WORK.NAND
    PORT MAP (
        A => S2986,
        B => S2999,
        Y => S3000
    );
NOR_851: ENTITY WORK.NOR
    PORT MAP (
        A => S1444,
        B => S2985,
        Y => S3001
    );
NOR_852: ENTITY WORK.NOR
    PORT MAP (
        A => S1443,
        B => S2996,
        Y => S3002
    );
NAND_1713: ENTITY WORK.NAND
    PORT MAP (
        A => S2990,
        B => S3002,
        Y => S3003
    );
NAND_1714: ENTITY WORK.NAND
    PORT MAP (
        A => S1449,
        B => S3003,
        Y => S3004
    );
NOR_853: ENTITY WORK.NOR
    PORT MAP (
        A => S3001,
        B => S3004,
        Y => S3005
    );
NAND_1715: ENTITY WORK.NAND
    PORT MAP (
        A => S1449,
        B => S3000,
        Y => S3006
    );
NOR_854: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_78,
        B => S1438,
        Y => S3007
    );
NAND_1716: ENTITY WORK.NAND
    PORT MAP (
        A => S7498,
        B => S1437,
        Y => S3008
    );
NOR_855: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_14,
        B => S1437,
        Y => S3009
    );
NAND_1717: ENTITY WORK.NAND
    PORT MAP (
        A => S7542,
        B => S1438,
        Y => S3010
    );
NOR_856: ENTITY WORK.NOR
    PORT MAP (
        A => S3007,
        B => S3009,
        Y => S3011
    );
NAND_1718: ENTITY WORK.NAND
    PORT MAP (
        A => S3008,
        B => S3010,
        Y => S3012
    );
NOR_857: ENTITY WORK.NOR
    PORT MAP (
        A => S1460,
        B => S3012,
        Y => S3013
    );
NAND_1719: ENTITY WORK.NAND
    PORT MAP (
        A => S1459,
        B => S3011,
        Y => S3014
    );
NAND_1720: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_30,
        B => S1438,
        Y => S3015
    );
NAND_1721: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_94,
        B => S1437,
        Y => S3016
    );
NAND_1722: ENTITY WORK.NAND
    PORT MAP (
        A => S3015,
        B => S3016,
        Y => S3017
    );
NAND_1723: ENTITY WORK.NAND
    PORT MAP (
        A => S1926,
        B => S3017,
        Y => S3018
    );
NAND_1724: ENTITY WORK.NAND
    PORT MAP (
        A => S3014,
        B => S3018,
        Y => S3019
    );
NOT_302: ENTITY WORK.NOT
    PORT MAP (
        A => S3019,
        Y => S3020
    );
NAND_1725: ENTITY WORK.NAND
    PORT MAP (
        A => S7509,
        B => S1438,
        Y => S3021
    );
NOR_858: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_126,
        B => S1438,
        Y => S3022
    );
NOR_859: ENTITY WORK.NOR
    PORT MAP (
        A => S1458,
        B => S3022,
        Y => S3023
    );
NAND_1726: ENTITY WORK.NAND
    PORT MAP (
        A => S3021,
        B => S3023,
        Y => S3024
    );
NOR_860: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_46,
        B => S1437,
        Y => S3025
    );
NOR_861: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_110,
        B => S1438,
        Y => S3026
    );
NOR_862: ENTITY WORK.NOR
    PORT MAP (
        A => S3025,
        B => S3026,
        Y => S3027
    );
NAND_1727: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S3027,
        Y => S3028
    );
NAND_1728: ENTITY WORK.NAND
    PORT MAP (
        A => S3024,
        B => S3028,
        Y => S3029
    );
NAND_1729: ENTITY WORK.NAND
    PORT MAP (
        A => S1487,
        B => S3029,
        Y => S3030
    );
NAND_1730: ENTITY WORK.NAND
    PORT MAP (
        A => S3018,
        B => S3030,
        Y => S3031
    );
NOR_863: ENTITY WORK.NOR
    PORT MAP (
        A => S3013,
        B => S3031,
        Y => S3032
    );
NAND_1731: ENTITY WORK.NAND
    PORT MAP (
        A => S3020,
        B => S3030,
        Y => S3033
    );
NOR_864: ENTITY WORK.NOR
    PORT MAP (
        A => S3005,
        B => S3033,
        Y => S3034
    );
NAND_1732: ENTITY WORK.NAND
    PORT MAP (
        A => S3006,
        B => S3032,
        Y => S3035
    );
NOR_865: ENTITY WORK.NOR
    PORT MAP (
        A => S1461,
        B => S3034,
        Y => S3036
    );
NAND_1733: ENTITY WORK.NAND
    PORT MAP (
        A => S1462,
        B => S3035,
        Y => S3037
    );
NAND_1734: ENTITY WORK.NAND
    PORT MAP (
        A => S1429,
        B => S3036,
        Y => S3038
    );
NAND_1735: ENTITY WORK.NAND
    PORT MAP (
        A => S2369,
        B => S3038,
        Y => S3039
    );
NOT_303: ENTITY WORK.NOT
    PORT MAP (
        A => S3039,
        Y => S3040
    );
NAND_1736: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_14,
        B => S3040,
        Y => S3041
    );
NOT_304: ENTITY WORK.NOT
    PORT MAP (
        A => S3041,
        Y => S3042
    );
NAND_1737: ENTITY WORK.NAND
    PORT MAP (
        A => S492,
        B => S3039,
        Y => S3043
    );
NOT_305: ENTITY WORK.NOT
    PORT MAP (
        A => S3043,
        Y => S3044
    );
NOR_866: ENTITY WORK.NOR
    PORT MAP (
        A => S3042,
        B => S3044,
        Y => S3045
    );
NOT_306: ENTITY WORK.NOT
    PORT MAP (
        A => S3045,
        Y => S3046
    );
NOR_867: ENTITY WORK.NOR
    PORT MAP (
        A => S2925,
        B => S2931,
        Y => S3047
    );
NOR_868: ENTITY WORK.NOR
    PORT MAP (
        A => S2927,
        B => S3047,
        Y => S3048
    );
NAND_1738: ENTITY WORK.NAND
    PORT MAP (
        A => S3045,
        B => S3048,
        Y => S3049
    );
NOR_869: ENTITY WORK.NOR
    PORT MAP (
        A => S3045,
        B => S3048,
        Y => S3050
    );
NOR_870: ENTITY WORK.NOR
    PORT MAP (
        A => S1526,
        B => S3050,
        Y => S3051
    );
NAND_1739: ENTITY WORK.NAND
    PORT MAP (
        A => S3049,
        B => S3051,
        Y => S3052
    );
NAND_1740: ENTITY WORK.NAND
    PORT MAP (
        A => S2939,
        B => S2949,
        Y => S3053
    );
NOR_871: ENTITY WORK.NOR
    PORT MAP (
        A => S2940,
        B => S3053,
        Y => S3054
    );
NOR_872: ENTITY WORK.NOR
    PORT MAP (
        A => S3045,
        B => S3054,
        Y => S3055
    );
NOT_307: ENTITY WORK.NOT
    PORT MAP (
        A => S3055,
        Y => S3056
    );
NAND_1741: ENTITY WORK.NAND
    PORT MAP (
        A => S3045,
        B => S3054,
        Y => S3057
    );
NAND_1742: ENTITY WORK.NAND
    PORT MAP (
        A => S1527,
        B => S3057,
        Y => S3058
    );
NOR_873: ENTITY WORK.NOR
    PORT MAP (
        A => S3055,
        B => S3058,
        Y => S3059
    );
NAND_1743: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_14,
        B => S3039,
        Y => S3060
    );
NOR_874: ENTITY WORK.NOR
    PORT MAP (
        A => S1533,
        B => S3060,
        Y => S3061
    );
NAND_1744: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_shiftunit_2387_A,
        B => S1614,
        Y => S3062
    );
NAND_1745: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_shiftunit_2691_A,
        B => S1609,
        Y => S3063
    );
NOR_875: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_muxmem_in2_14,
        B => S1359,
        Y => S3064
    );
NOT_308: ENTITY WORK.NOT
    PORT MAP (
        A => S3064,
        Y => S3065
    );
NAND_1746: ENTITY WORK.NAND
    PORT MAP (
        A => S1360,
        B => S3065,
        Y => S3066
    );
NOR_876: ENTITY WORK.NOR
    PORT MAP (
        A => S1623,
        B => S3066,
        Y => S3067
    );
NOR_877: ENTITY WORK.NOR
    PORT MAP (
        A => controller_opcode_2,
        B => S1396,
        Y => S3068
    );
NOR_878: ENTITY WORK.NOR
    PORT MAP (
        A => S2364,
        B => S3068,
        Y => S3069
    );
NOR_879: ENTITY WORK.NOR
    PORT MAP (
        A => S2053,
        B => S3069,
        Y => S3070
    );
NOR_880: ENTITY WORK.NOR
    PORT MAP (
        A => S1547,
        B => S3070,
        Y => S3071
    );
NAND_1747: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu2_14,
        B => S8570,
        Y => S3072
    );
NAND_1748: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_databusin_14,
        B => S1627,
        Y => S3073
    );
NAND_1749: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu1_14,
        B => S1377,
        Y => S3074
    );
NAND_1750: ENTITY WORK.NAND
    PORT MAP (
        A => S3072,
        B => S3073,
        Y => S3075
    );
NOR_881: ENTITY WORK.NOR
    PORT MAP (
        A => S3071,
        B => S3075,
        Y => S3076
    );
NAND_1751: ENTITY WORK.NAND
    PORT MAP (
        A => S3074,
        B => S3076,
        Y => S3077
    );
NOR_882: ENTITY WORK.NOR
    PORT MAP (
        A => S3067,
        B => S3077,
        Y => S3078
    );
NAND_1752: ENTITY WORK.NAND
    PORT MAP (
        A => S3063,
        B => S3078,
        Y => S3079
    );
NOT_309: ENTITY WORK.NOT
    PORT MAP (
        A => S3079,
        Y => S3080
    );
NAND_1753: ENTITY WORK.NAND
    PORT MAP (
        A => S3062,
        B => S3080,
        Y => S3081
    );
NOR_883: ENTITY WORK.NOR
    PORT MAP (
        A => S3061,
        B => S3081,
        Y => S3082
    );
NOR_884: ENTITY WORK.NOR
    PORT MAP (
        A => S492,
        B => S2945,
        Y => S3083
    );
NOR_885: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_14,
        B => S2946,
        Y => S3084
    );
NOR_886: ENTITY WORK.NOR
    PORT MAP (
        A => S3083,
        B => S3084,
        Y => S3085
    );
NAND_1754: ENTITY WORK.NAND
    PORT MAP (
        A => S1538,
        B => S3085,
        Y => S3086
    );
NAND_1755: ENTITY WORK.NAND
    PORT MAP (
        A => S3082,
        B => S3086,
        Y => S3087
    );
NOR_887: ENTITY WORK.NOR
    PORT MAP (
        A => S3059,
        B => S3087,
        Y => S3088
    );
NAND_1756: ENTITY WORK.NAND
    PORT MAP (
        A => S3052,
        B => S3088,
        Y => datapath_indatatrf_14
    );
NAND_1757: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_14,
        B => S1688,
        Y => S3089
    );
NAND_1758: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_78,
        B => S1689,
        Y => S3090
    );
NAND_1759: ENTITY WORK.NAND
    PORT MAP (
        A => S3089,
        B => S3090,
        Y => S18
    );
NAND_1760: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_159,
        B => S1438,
        Y => S3091
    );
NAND_1761: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_223,
        B => S1437,
        Y => S3092
    );
NAND_1762: ENTITY WORK.NAND
    PORT MAP (
        A => S3091,
        B => S3092,
        Y => S3093
    );
NAND_1763: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S3093,
        Y => S3094
    );
NOR_888: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_143,
        B => S1437,
        Y => S3095
    );
NOR_889: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_207,
        B => S1438,
        Y => S3096
    );
NOR_890: ENTITY WORK.NOR
    PORT MAP (
        A => S3095,
        B => S3096,
        Y => S3097
    );
NAND_1764: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S3097,
        Y => S3098
    );
NAND_1765: ENTITY WORK.NAND
    PORT MAP (
        A => S3094,
        B => S3098,
        Y => S3099
    );
NOR_891: ENTITY WORK.NOR
    PORT MAP (
        A => S1443,
        B => S3099,
        Y => S3100
    );
NOR_892: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_255,
        B => S1438,
        Y => S3101
    );
NAND_1766: ENTITY WORK.NAND
    PORT MAP (
        A => S7662,
        B => S1438,
        Y => S3102
    );
NAND_1767: ENTITY WORK.NAND
    PORT MAP (
        A => S1457,
        B => S3102,
        Y => S3103
    );
NOR_893: ENTITY WORK.NOR
    PORT MAP (
        A => S3101,
        B => S3103,
        Y => S3104
    );
NOR_894: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_239,
        B => S1438,
        Y => S3105
    );
NAND_1768: ENTITY WORK.NAND
    PORT MAP (
        A => S7574,
        B => S1438,
        Y => S3106
    );
NAND_1769: ENTITY WORK.NAND
    PORT MAP (
        A => S1458,
        B => S3106,
        Y => S3107
    );
NOR_895: ENTITY WORK.NOR
    PORT MAP (
        A => S3105,
        B => S3107,
        Y => S3108
    );
NOR_896: ENTITY WORK.NOR
    PORT MAP (
        A => S3104,
        B => S3108,
        Y => S3109
    );
NAND_1770: ENTITY WORK.NAND
    PORT MAP (
        A => S1443,
        B => S3109,
        Y => S3110
    );
NAND_1771: ENTITY WORK.NAND
    PORT MAP (
        A => S1449,
        B => S3110,
        Y => S3111
    );
NOR_897: ENTITY WORK.NOR
    PORT MAP (
        A => S1450,
        B => S3100,
        Y => S3112
    );
NOR_898: ENTITY WORK.NOR
    PORT MAP (
        A => S3100,
        B => S3111,
        Y => S3113
    );
NAND_1772: ENTITY WORK.NAND
    PORT MAP (
        A => S3110,
        B => S3112,
        Y => S3114
    );
NAND_1773: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_63,
        B => S1438,
        Y => S3115
    );
NAND_1774: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_127,
        B => S1437,
        Y => S3116
    );
NAND_1775: ENTITY WORK.NAND
    PORT MAP (
        A => S3115,
        B => S3116,
        Y => S3117
    );
NOR_899: ENTITY WORK.NOR
    PORT MAP (
        A => S1458,
        B => S3117,
        Y => S3118
    );
NOR_900: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_47,
        B => S1437,
        Y => S3119
    );
NOR_901: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_theregisterfile_memtrf_111,
        B => S1438,
        Y => S3120
    );
NOR_902: ENTITY WORK.NOR
    PORT MAP (
        A => S3119,
        B => S3120,
        Y => S3121
    );
NOR_903: ENTITY WORK.NOR
    PORT MAP (
        A => S1457,
        B => S3121,
        Y => S3122
    );
NOR_904: ENTITY WORK.NOR
    PORT MAP (
        A => S3118,
        B => S3122,
        Y => S3123
    );
NAND_1776: ENTITY WORK.NAND
    PORT MAP (
        A => S1487,
        B => S3123,
        Y => S3124
    );
NAND_1777: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_15,
        B => S1438,
        Y => S3125
    );
NAND_1778: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_79,
        B => S1437,
        Y => S3126
    );
NAND_1779: ENTITY WORK.NAND
    PORT MAP (
        A => S3125,
        B => S3126,
        Y => S3127
    );
NOT_310: ENTITY WORK.NOT
    PORT MAP (
        A => S3127,
        Y => S3128
    );
NOR_905: ENTITY WORK.NOR
    PORT MAP (
        A => S1460,
        B => S3128,
        Y => S3129
    );
NAND_1780: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_31,
        B => S1438,
        Y => S3130
    );
NAND_1781: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_95,
        B => S1437,
        Y => S3131
    );
NAND_1782: ENTITY WORK.NAND
    PORT MAP (
        A => S3130,
        B => S3131,
        Y => S3132
    );
NAND_1783: ENTITY WORK.NAND
    PORT MAP (
        A => S1926,
        B => S3132,
        Y => S3133
    );
NOT_311: ENTITY WORK.NOT
    PORT MAP (
        A => S3133,
        Y => S3134
    );
NOR_906: ENTITY WORK.NOR
    PORT MAP (
        A => S3129,
        B => S3134,
        Y => S3135
    );
NAND_1784: ENTITY WORK.NAND
    PORT MAP (
        A => S3124,
        B => S3133,
        Y => S3136
    );
NOR_907: ENTITY WORK.NOR
    PORT MAP (
        A => S3129,
        B => S3136,
        Y => S3137
    );
NAND_1785: ENTITY WORK.NAND
    PORT MAP (
        A => S3124,
        B => S3135,
        Y => S3138
    );
NOR_908: ENTITY WORK.NOR
    PORT MAP (
        A => S3113,
        B => S3138,
        Y => S3139
    );
NAND_1786: ENTITY WORK.NAND
    PORT MAP (
        A => S3114,
        B => S3137,
        Y => S3140
    );
NOR_909: ENTITY WORK.NOR
    PORT MAP (
        A => S1461,
        B => S3139,
        Y => S3141
    );
NAND_1787: ENTITY WORK.NAND
    PORT MAP (
        A => S1462,
        B => S3140,
        Y => S3142
    );
NOR_910: ENTITY WORK.NOR
    PORT MAP (
        A => S1430,
        B => S3142,
        Y => S3143
    );
NOR_911: ENTITY WORK.NOR
    PORT MAP (
        A => S2368,
        B => S3143,
        Y => S3144
    );
NOT_312: ENTITY WORK.NOT
    PORT MAP (
        A => S3144,
        Y => S3145
    );
NOR_912: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_15,
        B => S3144,
        Y => S3146
    );
NOT_313: ENTITY WORK.NOT
    PORT MAP (
        A => S3146,
        Y => S3147
    );
NOR_913: ENTITY WORK.NOR
    PORT MAP (
        A => S1304,
        B => S3145,
        Y => S3148
    );
NOT_314: ENTITY WORK.NOT
    PORT MAP (
        A => S3148,
        Y => S3149
    );
NAND_1788: ENTITY WORK.NAND
    PORT MAP (
        A => S3147,
        B => S3149,
        Y => S3150
    );
NAND_1789: ENTITY WORK.NAND
    PORT MAP (
        A => S3041,
        B => S3049,
        Y => S3151
    );
NOR_914: ENTITY WORK.NOR
    PORT MAP (
        A => S3150,
        B => S3151,
        Y => S3152
    );
NOT_315: ENTITY WORK.NOT
    PORT MAP (
        A => S3152,
        Y => S3153
    );
NAND_1790: ENTITY WORK.NAND
    PORT MAP (
        A => S3150,
        B => S3151,
        Y => S3154
    );
NAND_1791: ENTITY WORK.NAND
    PORT MAP (
        A => S3153,
        B => S3154,
        Y => S3155
    );
NAND_1792: ENTITY WORK.NAND
    PORT MAP (
        A => S1525,
        B => S3155,
        Y => S3156
    );
NAND_1793: ENTITY WORK.NAND
    PORT MAP (
        A => S3056,
        B => S3060,
        Y => S3157
    );
NAND_1794: ENTITY WORK.NAND
    PORT MAP (
        A => S3150,
        B => S3157,
        Y => S3158
    );
NOR_915: ENTITY WORK.NOR
    PORT MAP (
        A => S3150,
        B => S3157,
        Y => S3159
    );
NAND_1795: ENTITY WORK.NAND
    PORT MAP (
        A => S1527,
        B => S3158,
        Y => S3160
    );
NOR_916: ENTITY WORK.NOR
    PORT MAP (
        A => S3159,
        B => S3160,
        Y => S3161
    );
NAND_1796: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_shiftunit_2405_A,
        B => S1614,
        Y => S3162
    );
NOT_316: ENTITY WORK.NOT
    PORT MAP (
        A => S3162,
        Y => S3163
    );
NAND_1797: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_shiftunit_2708_A,
        B => S1609,
        Y => S3164
    );
NAND_1798: ENTITY WORK.NAND
    PORT MAP (
        A => S1364,
        B => S1622,
        Y => S3165
    );
NOR_917: ENTITY WORK.NOR
    PORT MAP (
        A => S2053,
        B => S2363,
        Y => S3166
    );
NOR_918: ENTITY WORK.NOR
    PORT MAP (
        A => S1547,
        B => S3166,
        Y => S3167
    );
NAND_1799: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_databusin_15,
        B => S1627,
        Y => S3168
    );
NAND_1800: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu2_15,
        B => S8570,
        Y => S3169
    );
NAND_1801: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu1_15,
        B => S1377,
        Y => S3170
    );
NAND_1802: ENTITY WORK.NAND
    PORT MAP (
        A => S3169,
        B => S3170,
        Y => S3171
    );
NOT_317: ENTITY WORK.NOT
    PORT MAP (
        A => S3171,
        Y => S3172
    );
NAND_1803: ENTITY WORK.NAND
    PORT MAP (
        A => S3168,
        B => S3172,
        Y => S3173
    );
NOR_919: ENTITY WORK.NOR
    PORT MAP (
        A => S3167,
        B => S3173,
        Y => S3174
    );
NAND_1804: ENTITY WORK.NAND
    PORT MAP (
        A => S3165,
        B => S3174,
        Y => S3175
    );
NOR_920: ENTITY WORK.NOR
    PORT MAP (
        A => S3163,
        B => S3175,
        Y => S3176
    );
NAND_1805: ENTITY WORK.NAND
    PORT MAP (
        A => S3164,
        B => S3176,
        Y => S3177
    );
NAND_1806: ENTITY WORK.NAND
    PORT MAP (
        A => S1534,
        B => S3145,
        Y => S3178
    );
NOR_921: ENTITY WORK.NOR
    PORT MAP (
        A => S1304,
        B => S3178,
        Y => S3179
    );
NOR_922: ENTITY WORK.NOR
    PORT MAP (
        A => S3177,
        B => S3179,
        Y => S3180
    );
NAND_1807: ENTITY WORK.NAND
    PORT MAP (
        A => S1304,
        B => S3084,
        Y => S3181
    );
NOR_923: ENTITY WORK.NOR
    PORT MAP (
        A => S1304,
        B => S3084,
        Y => S3182
    );
NOR_924: ENTITY WORK.NOR
    PORT MAP (
        A => S1539,
        B => S3182,
        Y => S3183
    );
NAND_1808: ENTITY WORK.NAND
    PORT MAP (
        A => S3181,
        B => S3183,
        Y => S3184
    );
NAND_1809: ENTITY WORK.NAND
    PORT MAP (
        A => S3180,
        B => S3184,
        Y => S3185
    );
NOR_925: ENTITY WORK.NOR
    PORT MAP (
        A => S3161,
        B => S3185,
        Y => S3186
    );
NAND_1810: ENTITY WORK.NAND
    PORT MAP (
        A => S3156,
        B => S3186,
        Y => datapath_indatatrf_15
    );
NAND_1811: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_15,
        B => S1688,
        Y => S3187
    );
NAND_1812: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_79,
        B => S1689,
        Y => S3188
    );
NAND_1813: ENTITY WORK.NAND
    PORT MAP (
        A => S3187,
        B => S3188,
        Y => S19
    );
NOR_926: ENTITY WORK.NOR
    PORT MAP (
        A => S1655,
        B => S1662,
        Y => S3189
    );
NAND_1814: ENTITY WORK.NAND
    PORT MAP (
        A => S1654,
        B => S1661,
        Y => S3190
    );
NOR_927: ENTITY WORK.NOR
    PORT MAP (
        A => S1671,
        B => S1687,
        Y => S3191
    );
NAND_1815: ENTITY WORK.NAND
    PORT MAP (
        A => S1672,
        B => S1686,
        Y => S3192
    );
NOR_928: ENTITY WORK.NOR
    PORT MAP (
        A => S3190,
        B => S3192,
        Y => S3193
    );
NAND_1816: ENTITY WORK.NAND
    PORT MAP (
        A => S3189,
        B => S3191,
        Y => S3194
    );
NAND_1817: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_0,
        B => S3193,
        Y => S3195
    );
NAND_1818: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_32,
        B => S3194,
        Y => S3196
    );
NAND_1819: ENTITY WORK.NAND
    PORT MAP (
        A => S3195,
        B => S3196,
        Y => S20
    );
NAND_1820: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_1,
        B => S3193,
        Y => S3197
    );
NAND_1821: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_33,
        B => S3194,
        Y => S3198
    );
NAND_1822: ENTITY WORK.NAND
    PORT MAP (
        A => S3197,
        B => S3198,
        Y => S21
    );
NAND_1823: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_2,
        B => S3193,
        Y => S3199
    );
NAND_1824: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_34,
        B => S3194,
        Y => S3200
    );
NAND_1825: ENTITY WORK.NAND
    PORT MAP (
        A => S3199,
        B => S3200,
        Y => S22
    );
NAND_1826: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_3,
        B => S3193,
        Y => S3201
    );
NAND_1827: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_35,
        B => S3194,
        Y => S3202
    );
NAND_1828: ENTITY WORK.NAND
    PORT MAP (
        A => S3201,
        B => S3202,
        Y => S23
    );
NAND_1829: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_4,
        B => S3193,
        Y => S3203
    );
NAND_1830: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_36,
        B => S3194,
        Y => S3204
    );
NAND_1831: ENTITY WORK.NAND
    PORT MAP (
        A => S3203,
        B => S3204,
        Y => S24
    );
NAND_1832: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_5,
        B => S3193,
        Y => S3205
    );
NAND_1833: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_37,
        B => S3194,
        Y => S3206
    );
NAND_1834: ENTITY WORK.NAND
    PORT MAP (
        A => S3205,
        B => S3206,
        Y => S25
    );
NAND_1835: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_6,
        B => S3193,
        Y => S3207
    );
NAND_1836: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_38,
        B => S3194,
        Y => S3208
    );
NAND_1837: ENTITY WORK.NAND
    PORT MAP (
        A => S3207,
        B => S3208,
        Y => S26
    );
NAND_1838: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_7,
        B => S3193,
        Y => S3209
    );
NAND_1839: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_39,
        B => S3194,
        Y => S3210
    );
NAND_1840: ENTITY WORK.NAND
    PORT MAP (
        A => S3209,
        B => S3210,
        Y => S27
    );
NAND_1841: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_8,
        B => S3193,
        Y => S3211
    );
NAND_1842: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_40,
        B => S3194,
        Y => S3212
    );
NAND_1843: ENTITY WORK.NAND
    PORT MAP (
        A => S3211,
        B => S3212,
        Y => S28
    );
NAND_1844: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_9,
        B => S3193,
        Y => S3213
    );
NAND_1845: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_41,
        B => S3194,
        Y => S3214
    );
NAND_1846: ENTITY WORK.NAND
    PORT MAP (
        A => S3213,
        B => S3214,
        Y => S29
    );
NAND_1847: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_10,
        B => S3193,
        Y => S3215
    );
NAND_1848: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_42,
        B => S3194,
        Y => S3216
    );
NAND_1849: ENTITY WORK.NAND
    PORT MAP (
        A => S3215,
        B => S3216,
        Y => S30
    );
NAND_1850: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_11,
        B => S3193,
        Y => S3217
    );
NAND_1851: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_43,
        B => S3194,
        Y => S3218
    );
NAND_1852: ENTITY WORK.NAND
    PORT MAP (
        A => S3217,
        B => S3218,
        Y => S31
    );
NAND_1853: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_12,
        B => S3193,
        Y => S3219
    );
NAND_1854: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_44,
        B => S3194,
        Y => S3220
    );
NAND_1855: ENTITY WORK.NAND
    PORT MAP (
        A => S3219,
        B => S3220,
        Y => S32
    );
NAND_1856: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_13,
        B => S3193,
        Y => S3221
    );
NAND_1857: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_45,
        B => S3194,
        Y => S3222
    );
NAND_1858: ENTITY WORK.NAND
    PORT MAP (
        A => S3221,
        B => S3222,
        Y => S33
    );
NAND_1859: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_14,
        B => S3193,
        Y => S3223
    );
NAND_1860: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_46,
        B => S3194,
        Y => S3224
    );
NAND_1861: ENTITY WORK.NAND
    PORT MAP (
        A => S3223,
        B => S3224,
        Y => S34
    );
NAND_1862: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_15,
        B => S3193,
        Y => S3225
    );
NAND_1863: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_47,
        B => S3194,
        Y => S3226
    );
NAND_1864: ENTITY WORK.NAND
    PORT MAP (
        A => S3225,
        B => S3226,
        Y => S35
    );
NOR_929: ENTITY WORK.NOR
    PORT MAP (
        A => S1678,
        B => S1685,
        Y => S3227
    );
NAND_1865: ENTITY WORK.NAND
    PORT MAP (
        A => S1679,
        B => S1684,
        Y => S3228
    );
NOR_930: ENTITY WORK.NOR
    PORT MAP (
        A => S1671,
        B => S3228,
        Y => S3229
    );
NAND_1866: ENTITY WORK.NAND
    PORT MAP (
        A => S1672,
        B => S3227,
        Y => S3230
    );
NOR_931: ENTITY WORK.NOR
    PORT MAP (
        A => S3190,
        B => S3230,
        Y => S3231
    );
NAND_1867: ENTITY WORK.NAND
    PORT MAP (
        A => S3189,
        B => S3229,
        Y => S3232
    );
NAND_1868: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_0,
        B => S3231,
        Y => S3233
    );
NAND_1869: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_48,
        B => S3232,
        Y => S3234
    );
NAND_1870: ENTITY WORK.NAND
    PORT MAP (
        A => S3233,
        B => S3234,
        Y => S36
    );
NAND_1871: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_1,
        B => S3231,
        Y => S3235
    );
NAND_1872: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_49,
        B => S3232,
        Y => S3236
    );
NAND_1873: ENTITY WORK.NAND
    PORT MAP (
        A => S3235,
        B => S3236,
        Y => S37
    );
NAND_1874: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_2,
        B => S3231,
        Y => S3237
    );
NAND_1875: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_50,
        B => S3232,
        Y => S3238
    );
NAND_1876: ENTITY WORK.NAND
    PORT MAP (
        A => S3237,
        B => S3238,
        Y => S38
    );
NAND_1877: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_3,
        B => S3231,
        Y => S3239
    );
NAND_1878: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_51,
        B => S3232,
        Y => S3240
    );
NAND_1879: ENTITY WORK.NAND
    PORT MAP (
        A => S3239,
        B => S3240,
        Y => S39
    );
NAND_1880: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_4,
        B => S3231,
        Y => S3241
    );
NAND_1881: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_52,
        B => S3232,
        Y => S3242
    );
NAND_1882: ENTITY WORK.NAND
    PORT MAP (
        A => S3241,
        B => S3242,
        Y => S40
    );
NAND_1883: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_5,
        B => S3231,
        Y => S3243
    );
NAND_1884: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_53,
        B => S3232,
        Y => S3244
    );
NAND_1885: ENTITY WORK.NAND
    PORT MAP (
        A => S3243,
        B => S3244,
        Y => S41
    );
NAND_1886: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_6,
        B => S3231,
        Y => S3245
    );
NAND_1887: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_54,
        B => S3232,
        Y => S3246
    );
NAND_1888: ENTITY WORK.NAND
    PORT MAP (
        A => S3245,
        B => S3246,
        Y => S42
    );
NAND_1889: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_7,
        B => S3231,
        Y => S3247
    );
NAND_1890: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_55,
        B => S3232,
        Y => S3248
    );
NAND_1891: ENTITY WORK.NAND
    PORT MAP (
        A => S3247,
        B => S3248,
        Y => S43
    );
NAND_1892: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_8,
        B => S3231,
        Y => S3249
    );
NAND_1893: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_56,
        B => S3232,
        Y => S3250
    );
NAND_1894: ENTITY WORK.NAND
    PORT MAP (
        A => S3249,
        B => S3250,
        Y => S44
    );
NAND_1895: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_9,
        B => S3231,
        Y => S3251
    );
NAND_1896: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_57,
        B => S3232,
        Y => S3252
    );
NAND_1897: ENTITY WORK.NAND
    PORT MAP (
        A => S3251,
        B => S3252,
        Y => S45
    );
NAND_1898: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_10,
        B => S3231,
        Y => S3253
    );
NAND_1899: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_58,
        B => S3232,
        Y => S3254
    );
NAND_1900: ENTITY WORK.NAND
    PORT MAP (
        A => S3253,
        B => S3254,
        Y => S46
    );
NAND_1901: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_11,
        B => S3231,
        Y => S3255
    );
NAND_1902: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_59,
        B => S3232,
        Y => S3256
    );
NAND_1903: ENTITY WORK.NAND
    PORT MAP (
        A => S3255,
        B => S3256,
        Y => S47
    );
NAND_1904: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_12,
        B => S3231,
        Y => S3257
    );
NAND_1905: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_60,
        B => S3232,
        Y => S3258
    );
NAND_1906: ENTITY WORK.NAND
    PORT MAP (
        A => S3257,
        B => S3258,
        Y => S48
    );
NAND_1907: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_13,
        B => S3231,
        Y => S3259
    );
NAND_1908: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_61,
        B => S3232,
        Y => S3260
    );
NAND_1909: ENTITY WORK.NAND
    PORT MAP (
        A => S3259,
        B => S3260,
        Y => S49
    );
NAND_1910: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_14,
        B => S3231,
        Y => S3261
    );
NAND_1911: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_62,
        B => S3232,
        Y => S3262
    );
NAND_1912: ENTITY WORK.NAND
    PORT MAP (
        A => S3261,
        B => S3262,
        Y => S50
    );
NAND_1913: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_15,
        B => S3231,
        Y => S3263
    );
NAND_1914: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_63,
        B => S3232,
        Y => S3264
    );
NAND_1915: ENTITY WORK.NAND
    PORT MAP (
        A => S3263,
        B => S3264,
        Y => S51
    );
NOR_932: ENTITY WORK.NOR
    PORT MAP (
        A => S1655,
        B => S1661,
        Y => S3265
    );
NAND_1916: ENTITY WORK.NAND
    PORT MAP (
        A => S1654,
        B => S1662,
        Y => S3266
    );
NOR_933: ENTITY WORK.NOR
    PORT MAP (
        A => S1672,
        B => S3266,
        Y => S3267
    );
NAND_1917: ENTITY WORK.NAND
    PORT MAP (
        A => S1671,
        B => S3265,
        Y => S3268
    );
NOR_934: ENTITY WORK.NOR
    PORT MAP (
        A => S1687,
        B => S3268,
        Y => S3269
    );
NAND_1918: ENTITY WORK.NAND
    PORT MAP (
        A => S1686,
        B => S3267,
        Y => S3270
    );
NAND_1919: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_0,
        B => S3269,
        Y => S3271
    );
NAND_1920: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_128,
        B => S3270,
        Y => S3272
    );
NAND_1921: ENTITY WORK.NAND
    PORT MAP (
        A => S3271,
        B => S3272,
        Y => S52
    );
NAND_1922: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_1,
        B => S3269,
        Y => S3273
    );
NAND_1923: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_129,
        B => S3270,
        Y => S3274
    );
NAND_1924: ENTITY WORK.NAND
    PORT MAP (
        A => S3273,
        B => S3274,
        Y => S53
    );
NAND_1925: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_2,
        B => S3269,
        Y => S3275
    );
NAND_1926: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_130,
        B => S3270,
        Y => S3276
    );
NAND_1927: ENTITY WORK.NAND
    PORT MAP (
        A => S3275,
        B => S3276,
        Y => S54
    );
NAND_1928: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_3,
        B => S3269,
        Y => S3277
    );
NAND_1929: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_131,
        B => S3270,
        Y => S3278
    );
NAND_1930: ENTITY WORK.NAND
    PORT MAP (
        A => S3277,
        B => S3278,
        Y => S55
    );
NAND_1931: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_4,
        B => S3269,
        Y => S3279
    );
NAND_1932: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_132,
        B => S3270,
        Y => S3280
    );
NAND_1933: ENTITY WORK.NAND
    PORT MAP (
        A => S3279,
        B => S3280,
        Y => S56
    );
NAND_1934: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_5,
        B => S3269,
        Y => S3281
    );
NAND_1935: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_133,
        B => S3270,
        Y => S3282
    );
NAND_1936: ENTITY WORK.NAND
    PORT MAP (
        A => S3281,
        B => S3282,
        Y => S57
    );
NAND_1937: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_6,
        B => S3269,
        Y => S3283
    );
NAND_1938: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_134,
        B => S3270,
        Y => S3284
    );
NAND_1939: ENTITY WORK.NAND
    PORT MAP (
        A => S3283,
        B => S3284,
        Y => S58
    );
NAND_1940: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_7,
        B => S3269,
        Y => S3285
    );
NAND_1941: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_135,
        B => S3270,
        Y => S3286
    );
NAND_1942: ENTITY WORK.NAND
    PORT MAP (
        A => S3285,
        B => S3286,
        Y => S59
    );
NAND_1943: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_8,
        B => S3269,
        Y => S3287
    );
NAND_1944: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_136,
        B => S3270,
        Y => S3288
    );
NAND_1945: ENTITY WORK.NAND
    PORT MAP (
        A => S3287,
        B => S3288,
        Y => S60
    );
NAND_1946: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_9,
        B => S3269,
        Y => S3289
    );
NAND_1947: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_137,
        B => S3270,
        Y => S3290
    );
NAND_1948: ENTITY WORK.NAND
    PORT MAP (
        A => S3289,
        B => S3290,
        Y => S61
    );
NAND_1949: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_10,
        B => S3269,
        Y => S3291
    );
NAND_1950: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_138,
        B => S3270,
        Y => S3292
    );
NAND_1951: ENTITY WORK.NAND
    PORT MAP (
        A => S3291,
        B => S3292,
        Y => S62
    );
NAND_1952: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_11,
        B => S3269,
        Y => S3293
    );
NAND_1953: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_139,
        B => S3270,
        Y => S3294
    );
NAND_1954: ENTITY WORK.NAND
    PORT MAP (
        A => S3293,
        B => S3294,
        Y => S63
    );
NAND_1955: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_12,
        B => S3269,
        Y => S3295
    );
NAND_1956: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_140,
        B => S3270,
        Y => S3296
    );
NAND_1957: ENTITY WORK.NAND
    PORT MAP (
        A => S3295,
        B => S3296,
        Y => S64
    );
NAND_1958: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_13,
        B => S3269,
        Y => S3297
    );
NAND_1959: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_141,
        B => S3270,
        Y => S3298
    );
NAND_1960: ENTITY WORK.NAND
    PORT MAP (
        A => S3297,
        B => S3298,
        Y => S65
    );
NAND_1961: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_14,
        B => S3269,
        Y => S3299
    );
NAND_1962: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_142,
        B => S3270,
        Y => S3300
    );
NAND_1963: ENTITY WORK.NAND
    PORT MAP (
        A => S3299,
        B => S3300,
        Y => S66
    );
NAND_1964: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_15,
        B => S3269,
        Y => S3301
    );
NAND_1965: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_143,
        B => S3270,
        Y => S3302
    );
NAND_1966: ENTITY WORK.NAND
    PORT MAP (
        A => S3301,
        B => S3302,
        Y => S67
    );
NOR_935: ENTITY WORK.NOR
    PORT MAP (
        A => S1672,
        B => S3190,
        Y => S3303
    );
NAND_1967: ENTITY WORK.NAND
    PORT MAP (
        A => S1671,
        B => S3189,
        Y => S3304
    );
NOR_936: ENTITY WORK.NOR
    PORT MAP (
        A => S3228,
        B => S3304,
        Y => S3305
    );
NAND_1968: ENTITY WORK.NAND
    PORT MAP (
        A => S3227,
        B => S3303,
        Y => S3306
    );
NAND_1969: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_0,
        B => S3305,
        Y => S3307
    );
NAND_1970: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_16,
        B => S3306,
        Y => S3308
    );
NAND_1971: ENTITY WORK.NAND
    PORT MAP (
        A => S3307,
        B => S3308,
        Y => S68
    );
NAND_1972: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_1,
        B => S3305,
        Y => S3309
    );
NAND_1973: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_17,
        B => S3306,
        Y => S3310
    );
NAND_1974: ENTITY WORK.NAND
    PORT MAP (
        A => S3309,
        B => S3310,
        Y => S69
    );
NAND_1975: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_2,
        B => S3305,
        Y => S3311
    );
NAND_1976: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_18,
        B => S3306,
        Y => S3312
    );
NAND_1977: ENTITY WORK.NAND
    PORT MAP (
        A => S3311,
        B => S3312,
        Y => S70
    );
NAND_1978: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_3,
        B => S3305,
        Y => S3313
    );
NAND_1979: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_19,
        B => S3306,
        Y => S3314
    );
NAND_1980: ENTITY WORK.NAND
    PORT MAP (
        A => S3313,
        B => S3314,
        Y => S71
    );
NAND_1981: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_4,
        B => S3305,
        Y => S3315
    );
NAND_1982: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_20,
        B => S3306,
        Y => S3316
    );
NAND_1983: ENTITY WORK.NAND
    PORT MAP (
        A => S3315,
        B => S3316,
        Y => S72
    );
NAND_1984: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_5,
        B => S3305,
        Y => S3317
    );
NAND_1985: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_21,
        B => S3306,
        Y => S3318
    );
NAND_1986: ENTITY WORK.NAND
    PORT MAP (
        A => S3317,
        B => S3318,
        Y => S73
    );
NAND_1987: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_6,
        B => S3305,
        Y => S3319
    );
NAND_1988: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_22,
        B => S3306,
        Y => S3320
    );
NAND_1989: ENTITY WORK.NAND
    PORT MAP (
        A => S3319,
        B => S3320,
        Y => S74
    );
NAND_1990: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_7,
        B => S3305,
        Y => S3321
    );
NAND_1991: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_23,
        B => S3306,
        Y => S3322
    );
NAND_1992: ENTITY WORK.NAND
    PORT MAP (
        A => S3321,
        B => S3322,
        Y => S75
    );
NAND_1993: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_8,
        B => S3305,
        Y => S3323
    );
NAND_1994: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_24,
        B => S3306,
        Y => S3324
    );
NAND_1995: ENTITY WORK.NAND
    PORT MAP (
        A => S3323,
        B => S3324,
        Y => S76
    );
NAND_1996: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_9,
        B => S3305,
        Y => S3325
    );
NAND_1997: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_25,
        B => S3306,
        Y => S3326
    );
NAND_1998: ENTITY WORK.NAND
    PORT MAP (
        A => S3325,
        B => S3326,
        Y => S77
    );
NAND_1999: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_10,
        B => S3305,
        Y => S3327
    );
NAND_2000: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_26,
        B => S3306,
        Y => S3328
    );
NAND_2001: ENTITY WORK.NAND
    PORT MAP (
        A => S3327,
        B => S3328,
        Y => S78
    );
NAND_2002: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_11,
        B => S3305,
        Y => S3329
    );
NAND_2003: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_27,
        B => S3306,
        Y => S3330
    );
NAND_2004: ENTITY WORK.NAND
    PORT MAP (
        A => S3329,
        B => S3330,
        Y => S79
    );
NAND_2005: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_12,
        B => S3305,
        Y => S3331
    );
NAND_2006: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_28,
        B => S3306,
        Y => S3332
    );
NAND_2007: ENTITY WORK.NAND
    PORT MAP (
        A => S3331,
        B => S3332,
        Y => S80
    );
NAND_2008: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_13,
        B => S3305,
        Y => S3333
    );
NAND_2009: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_29,
        B => S3306,
        Y => S3334
    );
NAND_2010: ENTITY WORK.NAND
    PORT MAP (
        A => S3333,
        B => S3334,
        Y => S81
    );
NAND_2011: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_14,
        B => S3305,
        Y => S3335
    );
NAND_2012: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_30,
        B => S3306,
        Y => S3336
    );
NAND_2013: ENTITY WORK.NAND
    PORT MAP (
        A => S3335,
        B => S3336,
        Y => S82
    );
NAND_2014: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_15,
        B => S3305,
        Y => S3337
    );
NAND_2015: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_31,
        B => S3306,
        Y => S3338
    );
NAND_2016: ENTITY WORK.NAND
    PORT MAP (
        A => S3337,
        B => S3338,
        Y => S83
    );
NOR_937: ENTITY WORK.NOR
    PORT MAP (
        A => S1674,
        B => S3228,
        Y => S3339
    );
NAND_2017: ENTITY WORK.NAND
    PORT MAP (
        A => S1673,
        B => S3227,
        Y => S3340
    );
NAND_2018: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_0,
        B => S3339,
        Y => S3341
    );
NAND_2019: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_80,
        B => S3340,
        Y => S3342
    );
NAND_2020: ENTITY WORK.NAND
    PORT MAP (
        A => S3341,
        B => S3342,
        Y => S84
    );
NAND_2021: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_1,
        B => S3339,
        Y => S3343
    );
NAND_2022: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_81,
        B => S3340,
        Y => S3344
    );
NAND_2023: ENTITY WORK.NAND
    PORT MAP (
        A => S3343,
        B => S3344,
        Y => S85
    );
NAND_2024: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_2,
        B => S3339,
        Y => S3345
    );
NAND_2025: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_82,
        B => S3340,
        Y => S3346
    );
NAND_2026: ENTITY WORK.NAND
    PORT MAP (
        A => S3345,
        B => S3346,
        Y => S86
    );
NAND_2027: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_3,
        B => S3339,
        Y => S3347
    );
NAND_2028: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_83,
        B => S3340,
        Y => S3348
    );
NAND_2029: ENTITY WORK.NAND
    PORT MAP (
        A => S3347,
        B => S3348,
        Y => S87
    );
NAND_2030: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_4,
        B => S3339,
        Y => S3349
    );
NAND_2031: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_84,
        B => S3340,
        Y => S3350
    );
NAND_2032: ENTITY WORK.NAND
    PORT MAP (
        A => S3349,
        B => S3350,
        Y => S88
    );
NAND_2033: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_5,
        B => S3339,
        Y => S3351
    );
NAND_2034: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_85,
        B => S3340,
        Y => S3352
    );
NAND_2035: ENTITY WORK.NAND
    PORT MAP (
        A => S3351,
        B => S3352,
        Y => S89
    );
NAND_2036: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_6,
        B => S3339,
        Y => S3353
    );
NAND_2037: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_86,
        B => S3340,
        Y => S3354
    );
NAND_2038: ENTITY WORK.NAND
    PORT MAP (
        A => S3353,
        B => S3354,
        Y => S90
    );
NAND_2039: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_7,
        B => S3339,
        Y => S3355
    );
NAND_2040: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_87,
        B => S3340,
        Y => S3356
    );
NAND_2041: ENTITY WORK.NAND
    PORT MAP (
        A => S3355,
        B => S3356,
        Y => S91
    );
NAND_2042: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_8,
        B => S3339,
        Y => S3357
    );
NAND_2043: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_88,
        B => S3340,
        Y => S3358
    );
NAND_2044: ENTITY WORK.NAND
    PORT MAP (
        A => S3357,
        B => S3358,
        Y => S92
    );
NAND_2045: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_9,
        B => S3339,
        Y => S3359
    );
NAND_2046: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_89,
        B => S3340,
        Y => S3360
    );
NAND_2047: ENTITY WORK.NAND
    PORT MAP (
        A => S3359,
        B => S3360,
        Y => S93
    );
NAND_2048: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_10,
        B => S3339,
        Y => S3361
    );
NAND_2049: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_90,
        B => S3340,
        Y => S3362
    );
NAND_2050: ENTITY WORK.NAND
    PORT MAP (
        A => S3361,
        B => S3362,
        Y => S94
    );
NAND_2051: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_11,
        B => S3339,
        Y => S3363
    );
NAND_2052: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_91,
        B => S3340,
        Y => S3364
    );
NAND_2053: ENTITY WORK.NAND
    PORT MAP (
        A => S3363,
        B => S3364,
        Y => S95
    );
NAND_2054: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_12,
        B => S3339,
        Y => S3365
    );
NAND_2055: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_92,
        B => S3340,
        Y => S3366
    );
NAND_2056: ENTITY WORK.NAND
    PORT MAP (
        A => S3365,
        B => S3366,
        Y => S96
    );
NAND_2057: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_13,
        B => S3339,
        Y => S3367
    );
NAND_2058: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_93,
        B => S3340,
        Y => S3368
    );
NAND_2059: ENTITY WORK.NAND
    PORT MAP (
        A => S3367,
        B => S3368,
        Y => S97
    );
NAND_2060: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_14,
        B => S3339,
        Y => S3369
    );
NAND_2061: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_94,
        B => S3340,
        Y => S3370
    );
NAND_2062: ENTITY WORK.NAND
    PORT MAP (
        A => S3369,
        B => S3370,
        Y => S98
    );
NAND_2063: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_15,
        B => S3339,
        Y => S3371
    );
NAND_2064: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_95,
        B => S3340,
        Y => S3372
    );
NAND_2065: ENTITY WORK.NAND
    PORT MAP (
        A => S3371,
        B => S3372,
        Y => S99
    );
NOR_938: ENTITY WORK.NOR
    PORT MAP (
        A => S1664,
        B => S3192,
        Y => S3373
    );
NAND_2066: ENTITY WORK.NAND
    PORT MAP (
        A => S1663,
        B => S3191,
        Y => S3374
    );
NAND_2067: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_0,
        B => S3373,
        Y => S3375
    );
NAND_2068: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_96,
        B => S3374,
        Y => S3376
    );
NAND_2069: ENTITY WORK.NAND
    PORT MAP (
        A => S3375,
        B => S3376,
        Y => S100
    );
NAND_2070: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_1,
        B => S3373,
        Y => S3377
    );
NAND_2071: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_97,
        B => S3374,
        Y => S3378
    );
NAND_2072: ENTITY WORK.NAND
    PORT MAP (
        A => S3377,
        B => S3378,
        Y => S101
    );
NAND_2073: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_2,
        B => S3373,
        Y => S3379
    );
NAND_2074: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_98,
        B => S3374,
        Y => S3380
    );
NAND_2075: ENTITY WORK.NAND
    PORT MAP (
        A => S3379,
        B => S3380,
        Y => S102
    );
NAND_2076: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_3,
        B => S3373,
        Y => S3381
    );
NAND_2077: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_99,
        B => S3374,
        Y => S3382
    );
NAND_2078: ENTITY WORK.NAND
    PORT MAP (
        A => S3381,
        B => S3382,
        Y => S103
    );
NAND_2079: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_4,
        B => S3373,
        Y => S3383
    );
NAND_2080: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_100,
        B => S3374,
        Y => S3384
    );
NAND_2081: ENTITY WORK.NAND
    PORT MAP (
        A => S3383,
        B => S3384,
        Y => S104
    );
NAND_2082: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_5,
        B => S3373,
        Y => S3385
    );
NAND_2083: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_101,
        B => S3374,
        Y => S3386
    );
NAND_2084: ENTITY WORK.NAND
    PORT MAP (
        A => S3385,
        B => S3386,
        Y => S105
    );
NAND_2085: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_6,
        B => S3373,
        Y => S3387
    );
NAND_2086: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_102,
        B => S3374,
        Y => S3388
    );
NAND_2087: ENTITY WORK.NAND
    PORT MAP (
        A => S3387,
        B => S3388,
        Y => S106
    );
NAND_2088: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_7,
        B => S3373,
        Y => S3389
    );
NAND_2089: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_103,
        B => S3374,
        Y => S3390
    );
NAND_2090: ENTITY WORK.NAND
    PORT MAP (
        A => S3389,
        B => S3390,
        Y => S107
    );
NAND_2091: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_8,
        B => S3373,
        Y => S3391
    );
NAND_2092: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_104,
        B => S3374,
        Y => S3392
    );
NAND_2093: ENTITY WORK.NAND
    PORT MAP (
        A => S3391,
        B => S3392,
        Y => S108
    );
NAND_2094: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_9,
        B => S3373,
        Y => S3393
    );
NAND_2095: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_105,
        B => S3374,
        Y => S3394
    );
NAND_2096: ENTITY WORK.NAND
    PORT MAP (
        A => S3393,
        B => S3394,
        Y => S109
    );
NAND_2097: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_10,
        B => S3373,
        Y => S3395
    );
NAND_2098: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_106,
        B => S3374,
        Y => S3396
    );
NAND_2099: ENTITY WORK.NAND
    PORT MAP (
        A => S3395,
        B => S3396,
        Y => S110
    );
NAND_2100: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_11,
        B => S3373,
        Y => S3397
    );
NAND_2101: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_107,
        B => S3374,
        Y => S3398
    );
NAND_2102: ENTITY WORK.NAND
    PORT MAP (
        A => S3397,
        B => S3398,
        Y => S111
    );
NAND_2103: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_12,
        B => S3373,
        Y => S3399
    );
NAND_2104: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_108,
        B => S3374,
        Y => S3400
    );
NAND_2105: ENTITY WORK.NAND
    PORT MAP (
        A => S3399,
        B => S3400,
        Y => S112
    );
NAND_2106: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_13,
        B => S3373,
        Y => S3401
    );
NAND_2107: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_109,
        B => S3374,
        Y => S3402
    );
NAND_2108: ENTITY WORK.NAND
    PORT MAP (
        A => S3401,
        B => S3402,
        Y => S113
    );
NAND_2109: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_14,
        B => S3373,
        Y => S3403
    );
NAND_2110: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_110,
        B => S3374,
        Y => S3404
    );
NAND_2111: ENTITY WORK.NAND
    PORT MAP (
        A => S3403,
        B => S3404,
        Y => S114
    );
NAND_2112: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_15,
        B => S3373,
        Y => S3405
    );
NAND_2113: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_111,
        B => S3374,
        Y => S3406
    );
NAND_2114: ENTITY WORK.NAND
    PORT MAP (
        A => S3405,
        B => S3406,
        Y => S115
    );
NOR_939: ENTITY WORK.NOR
    PORT MAP (
        A => S1664,
        B => S3230,
        Y => S3407
    );
NAND_2115: ENTITY WORK.NAND
    PORT MAP (
        A => S1663,
        B => S3229,
        Y => S3408
    );
NAND_2116: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_0,
        B => S3407,
        Y => S3409
    );
NAND_2117: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_112,
        B => S3408,
        Y => S3410
    );
NAND_2118: ENTITY WORK.NAND
    PORT MAP (
        A => S3409,
        B => S3410,
        Y => S116
    );
NAND_2119: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_1,
        B => S3407,
        Y => S3411
    );
NAND_2120: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_113,
        B => S3408,
        Y => S3412
    );
NAND_2121: ENTITY WORK.NAND
    PORT MAP (
        A => S3411,
        B => S3412,
        Y => S117
    );
NAND_2122: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_2,
        B => S3407,
        Y => S3413
    );
NAND_2123: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_114,
        B => S3408,
        Y => S3414
    );
NAND_2124: ENTITY WORK.NAND
    PORT MAP (
        A => S3413,
        B => S3414,
        Y => S118
    );
NAND_2125: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_3,
        B => S3407,
        Y => S3415
    );
NAND_2126: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_115,
        B => S3408,
        Y => S3416
    );
NAND_2127: ENTITY WORK.NAND
    PORT MAP (
        A => S3415,
        B => S3416,
        Y => S119
    );
NAND_2128: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_4,
        B => S3407,
        Y => S3417
    );
NAND_2129: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_116,
        B => S3408,
        Y => S3418
    );
NAND_2130: ENTITY WORK.NAND
    PORT MAP (
        A => S3417,
        B => S3418,
        Y => S120
    );
NAND_2131: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_5,
        B => S3407,
        Y => S3419
    );
NAND_2132: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_117,
        B => S3408,
        Y => S3420
    );
NAND_2133: ENTITY WORK.NAND
    PORT MAP (
        A => S3419,
        B => S3420,
        Y => S121
    );
NAND_2134: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_6,
        B => S3407,
        Y => S3421
    );
NAND_2135: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_118,
        B => S3408,
        Y => S3422
    );
NAND_2136: ENTITY WORK.NAND
    PORT MAP (
        A => S3421,
        B => S3422,
        Y => S122
    );
NAND_2137: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_7,
        B => S3407,
        Y => S3423
    );
NAND_2138: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_119,
        B => S3408,
        Y => S3424
    );
NAND_2139: ENTITY WORK.NAND
    PORT MAP (
        A => S3423,
        B => S3424,
        Y => S123
    );
NAND_2140: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_8,
        B => S3407,
        Y => S3425
    );
NAND_2141: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_120,
        B => S3408,
        Y => S3426
    );
NAND_2142: ENTITY WORK.NAND
    PORT MAP (
        A => S3425,
        B => S3426,
        Y => S124
    );
NAND_2143: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_9,
        B => S3407,
        Y => S3427
    );
NAND_2144: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_121,
        B => S3408,
        Y => S3428
    );
NAND_2145: ENTITY WORK.NAND
    PORT MAP (
        A => S3427,
        B => S3428,
        Y => S125
    );
NAND_2146: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_10,
        B => S3407,
        Y => S3429
    );
NAND_2147: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_122,
        B => S3408,
        Y => S3430
    );
NAND_2148: ENTITY WORK.NAND
    PORT MAP (
        A => S3429,
        B => S3430,
        Y => S126
    );
NAND_2149: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_11,
        B => S3407,
        Y => S3431
    );
NAND_2150: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_123,
        B => S3408,
        Y => S3432
    );
NAND_2151: ENTITY WORK.NAND
    PORT MAP (
        A => S3431,
        B => S3432,
        Y => S127
    );
NAND_2152: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_12,
        B => S3407,
        Y => S3433
    );
NAND_2153: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_124,
        B => S3408,
        Y => S3434
    );
NAND_2154: ENTITY WORK.NAND
    PORT MAP (
        A => S3433,
        B => S3434,
        Y => S128
    );
NAND_2155: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_13,
        B => S3407,
        Y => S3435
    );
NAND_2156: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_125,
        B => S3408,
        Y => S3436
    );
NAND_2157: ENTITY WORK.NAND
    PORT MAP (
        A => S3435,
        B => S3436,
        Y => S129
    );
NAND_2158: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_14,
        B => S3407,
        Y => S3437
    );
NAND_2159: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_126,
        B => S3408,
        Y => S3438
    );
NAND_2160: ENTITY WORK.NAND
    PORT MAP (
        A => S3437,
        B => S3438,
        Y => S130
    );
NAND_2161: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_15,
        B => S3407,
        Y => S3439
    );
NAND_2162: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_127,
        B => S3408,
        Y => S3440
    );
NAND_2163: ENTITY WORK.NAND
    PORT MAP (
        A => S3439,
        B => S3440,
        Y => S131
    );
NOR_940: ENTITY WORK.NOR
    PORT MAP (
        A => S1687,
        B => S3304,
        Y => S3441
    );
NAND_2164: ENTITY WORK.NAND
    PORT MAP (
        A => S1686,
        B => S3303,
        Y => S3442
    );
NAND_2165: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_0,
        B => S3441,
        Y => S3443
    );
NAND_2166: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_0,
        B => S3442,
        Y => S3444
    );
NAND_2167: ENTITY WORK.NAND
    PORT MAP (
        A => S3443,
        B => S3444,
        Y => S132
    );
NAND_2168: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_1,
        B => S3441,
        Y => S3445
    );
NAND_2169: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_1,
        B => S3442,
        Y => S3446
    );
NAND_2170: ENTITY WORK.NAND
    PORT MAP (
        A => S3445,
        B => S3446,
        Y => S133
    );
NAND_2171: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_2,
        B => S3441,
        Y => S3447
    );
NAND_2172: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_2,
        B => S3442,
        Y => S3448
    );
NAND_2173: ENTITY WORK.NAND
    PORT MAP (
        A => S3447,
        B => S3448,
        Y => S134
    );
NAND_2174: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_3,
        B => S3441,
        Y => S3449
    );
NAND_2175: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_3,
        B => S3442,
        Y => S3450
    );
NAND_2176: ENTITY WORK.NAND
    PORT MAP (
        A => S3449,
        B => S3450,
        Y => S135
    );
NAND_2177: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_4,
        B => S3441,
        Y => S3451
    );
NAND_2178: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_4,
        B => S3442,
        Y => S3452
    );
NAND_2179: ENTITY WORK.NAND
    PORT MAP (
        A => S3451,
        B => S3452,
        Y => S136
    );
NAND_2180: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_5,
        B => S3441,
        Y => S3453
    );
NAND_2181: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_5,
        B => S3442,
        Y => S3454
    );
NAND_2182: ENTITY WORK.NAND
    PORT MAP (
        A => S3453,
        B => S3454,
        Y => S137
    );
NAND_2183: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_6,
        B => S3441,
        Y => S3455
    );
NAND_2184: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_6,
        B => S3442,
        Y => S3456
    );
NAND_2185: ENTITY WORK.NAND
    PORT MAP (
        A => S3455,
        B => S3456,
        Y => S138
    );
NAND_2186: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_7,
        B => S3441,
        Y => S3457
    );
NAND_2187: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_7,
        B => S3442,
        Y => S3458
    );
NAND_2188: ENTITY WORK.NAND
    PORT MAP (
        A => S3457,
        B => S3458,
        Y => S139
    );
NAND_2189: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_8,
        B => S3441,
        Y => S3459
    );
NAND_2190: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_8,
        B => S3442,
        Y => S3460
    );
NAND_2191: ENTITY WORK.NAND
    PORT MAP (
        A => S3459,
        B => S3460,
        Y => S140
    );
NAND_2192: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_9,
        B => S3441,
        Y => S3461
    );
NAND_2193: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_9,
        B => S3442,
        Y => S3462
    );
NAND_2194: ENTITY WORK.NAND
    PORT MAP (
        A => S3461,
        B => S3462,
        Y => S141
    );
NAND_2195: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_10,
        B => S3441,
        Y => S3463
    );
NAND_2196: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_10,
        B => S3442,
        Y => S3464
    );
NAND_2197: ENTITY WORK.NAND
    PORT MAP (
        A => S3463,
        B => S3464,
        Y => S142
    );
NAND_2198: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_11,
        B => S3441,
        Y => S3465
    );
NAND_2199: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_11,
        B => S3442,
        Y => S3466
    );
NAND_2200: ENTITY WORK.NAND
    PORT MAP (
        A => S3465,
        B => S3466,
        Y => S143
    );
NAND_2201: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_12,
        B => S3441,
        Y => S3467
    );
NAND_2202: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_12,
        B => S3442,
        Y => S3468
    );
NAND_2203: ENTITY WORK.NAND
    PORT MAP (
        A => S3467,
        B => S3468,
        Y => S144
    );
NAND_2204: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_13,
        B => S3441,
        Y => S3469
    );
NAND_2205: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_13,
        B => S3442,
        Y => S3470
    );
NAND_2206: ENTITY WORK.NAND
    PORT MAP (
        A => S3469,
        B => S3470,
        Y => S145
    );
NAND_2207: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_14,
        B => S3441,
        Y => S3471
    );
NAND_2208: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_14,
        B => S3442,
        Y => S3472
    );
NAND_2209: ENTITY WORK.NAND
    PORT MAP (
        A => S3471,
        B => S3472,
        Y => S146
    );
NAND_2210: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_15,
        B => S3441,
        Y => S3473
    );
NAND_2211: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_15,
        B => S3442,
        Y => S3474
    );
NAND_2212: ENTITY WORK.NAND
    PORT MAP (
        A => S3473,
        B => S3474,
        Y => S147
    );
NOR_941: ENTITY WORK.NOR
    PORT MAP (
        A => S3228,
        B => S3268,
        Y => S3475
    );
NAND_2213: ENTITY WORK.NAND
    PORT MAP (
        A => S3227,
        B => S3267,
        Y => S3476
    );
NAND_2214: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_0,
        B => S3475,
        Y => S3477
    );
NAND_2215: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_144,
        B => S3476,
        Y => S3478
    );
NAND_2216: ENTITY WORK.NAND
    PORT MAP (
        A => S3477,
        B => S3478,
        Y => S148
    );
NAND_2217: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_1,
        B => S3475,
        Y => S3479
    );
NAND_2218: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_145,
        B => S3476,
        Y => S3480
    );
NAND_2219: ENTITY WORK.NAND
    PORT MAP (
        A => S3479,
        B => S3480,
        Y => S149
    );
NAND_2220: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_2,
        B => S3475,
        Y => S3481
    );
NAND_2221: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_146,
        B => S3476,
        Y => S3482
    );
NAND_2222: ENTITY WORK.NAND
    PORT MAP (
        A => S3481,
        B => S3482,
        Y => S150
    );
NAND_2223: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_3,
        B => S3475,
        Y => S3483
    );
NAND_2224: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_147,
        B => S3476,
        Y => S3484
    );
NAND_2225: ENTITY WORK.NAND
    PORT MAP (
        A => S3483,
        B => S3484,
        Y => S151
    );
NAND_2226: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_4,
        B => S3475,
        Y => S3485
    );
NAND_2227: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_148,
        B => S3476,
        Y => S3486
    );
NAND_2228: ENTITY WORK.NAND
    PORT MAP (
        A => S3485,
        B => S3486,
        Y => S152
    );
NAND_2229: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_5,
        B => S3475,
        Y => S3487
    );
NAND_2230: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_149,
        B => S3476,
        Y => S3488
    );
NAND_2231: ENTITY WORK.NAND
    PORT MAP (
        A => S3487,
        B => S3488,
        Y => S153
    );
NAND_2232: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_6,
        B => S3475,
        Y => S3489
    );
NAND_2233: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_150,
        B => S3476,
        Y => S3490
    );
NAND_2234: ENTITY WORK.NAND
    PORT MAP (
        A => S3489,
        B => S3490,
        Y => S154
    );
NAND_2235: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_7,
        B => S3475,
        Y => S3491
    );
NAND_2236: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_151,
        B => S3476,
        Y => S3492
    );
NAND_2237: ENTITY WORK.NAND
    PORT MAP (
        A => S3491,
        B => S3492,
        Y => S155
    );
NAND_2238: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_8,
        B => S3475,
        Y => S3493
    );
NAND_2239: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_152,
        B => S3476,
        Y => S3494
    );
NAND_2240: ENTITY WORK.NAND
    PORT MAP (
        A => S3493,
        B => S3494,
        Y => S156
    );
NAND_2241: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_9,
        B => S3475,
        Y => S3495
    );
NAND_2242: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_153,
        B => S3476,
        Y => S3496
    );
NAND_2243: ENTITY WORK.NAND
    PORT MAP (
        A => S3495,
        B => S3496,
        Y => S157
    );
NAND_2244: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_10,
        B => S3475,
        Y => S3497
    );
NAND_2245: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_154,
        B => S3476,
        Y => S3498
    );
NAND_2246: ENTITY WORK.NAND
    PORT MAP (
        A => S3497,
        B => S3498,
        Y => S158
    );
NAND_2247: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_11,
        B => S3475,
        Y => S3499
    );
NAND_2248: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_155,
        B => S3476,
        Y => S3500
    );
NAND_2249: ENTITY WORK.NAND
    PORT MAP (
        A => S3499,
        B => S3500,
        Y => S159
    );
NAND_2250: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_12,
        B => S3475,
        Y => S3501
    );
NAND_2251: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_156,
        B => S3476,
        Y => S3502
    );
NAND_2252: ENTITY WORK.NAND
    PORT MAP (
        A => S3501,
        B => S3502,
        Y => S160
    );
NAND_2253: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_13,
        B => S3475,
        Y => S3503
    );
NAND_2254: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_157,
        B => S3476,
        Y => S3504
    );
NAND_2255: ENTITY WORK.NAND
    PORT MAP (
        A => S3503,
        B => S3504,
        Y => S161
    );
NAND_2256: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_14,
        B => S3475,
        Y => S3505
    );
NAND_2257: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_158,
        B => S3476,
        Y => S3506
    );
NAND_2258: ENTITY WORK.NAND
    PORT MAP (
        A => S3505,
        B => S3506,
        Y => S162
    );
NAND_2259: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_15,
        B => S3475,
        Y => S3507
    );
NAND_2260: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_159,
        B => S3476,
        Y => S3508
    );
NAND_2261: ENTITY WORK.NAND
    PORT MAP (
        A => S3507,
        B => S3508,
        Y => S163
    );
NOR_942: ENTITY WORK.NOR
    PORT MAP (
        A => S3192,
        B => S3266,
        Y => S3509
    );
NAND_2262: ENTITY WORK.NAND
    PORT MAP (
        A => S3191,
        B => S3265,
        Y => S3510
    );
NAND_2263: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_0,
        B => S3509,
        Y => S3511
    );
NAND_2264: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_160,
        B => S3510,
        Y => S3512
    );
NAND_2265: ENTITY WORK.NAND
    PORT MAP (
        A => S3511,
        B => S3512,
        Y => S164
    );
NAND_2266: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_1,
        B => S3509,
        Y => S3513
    );
NAND_2267: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_161,
        B => S3510,
        Y => S3514
    );
NAND_2268: ENTITY WORK.NAND
    PORT MAP (
        A => S3513,
        B => S3514,
        Y => S165
    );
NAND_2269: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_2,
        B => S3509,
        Y => S3515
    );
NAND_2270: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_162,
        B => S3510,
        Y => S3516
    );
NAND_2271: ENTITY WORK.NAND
    PORT MAP (
        A => S3515,
        B => S3516,
        Y => S166
    );
NAND_2272: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_3,
        B => S3509,
        Y => S3517
    );
NAND_2273: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_163,
        B => S3510,
        Y => S3518
    );
NAND_2274: ENTITY WORK.NAND
    PORT MAP (
        A => S3517,
        B => S3518,
        Y => S167
    );
NAND_2275: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_4,
        B => S3509,
        Y => S3519
    );
NAND_2276: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_164,
        B => S3510,
        Y => S3520
    );
NAND_2277: ENTITY WORK.NAND
    PORT MAP (
        A => S3519,
        B => S3520,
        Y => S168
    );
NAND_2278: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_5,
        B => S3509,
        Y => S3521
    );
NAND_2279: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_165,
        B => S3510,
        Y => S3522
    );
NAND_2280: ENTITY WORK.NAND
    PORT MAP (
        A => S3521,
        B => S3522,
        Y => S169
    );
NAND_2281: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_6,
        B => S3509,
        Y => S3523
    );
NAND_2282: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_166,
        B => S3510,
        Y => S3524
    );
NAND_2283: ENTITY WORK.NAND
    PORT MAP (
        A => S3523,
        B => S3524,
        Y => S170
    );
NAND_2284: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_7,
        B => S3509,
        Y => S3525
    );
NAND_2285: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_167,
        B => S3510,
        Y => S3526
    );
NAND_2286: ENTITY WORK.NAND
    PORT MAP (
        A => S3525,
        B => S3526,
        Y => S171
    );
NAND_2287: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_8,
        B => S3509,
        Y => S3527
    );
NAND_2288: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_168,
        B => S3510,
        Y => S3528
    );
NAND_2289: ENTITY WORK.NAND
    PORT MAP (
        A => S3527,
        B => S3528,
        Y => S172
    );
NAND_2290: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_9,
        B => S3509,
        Y => S3529
    );
NAND_2291: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_169,
        B => S3510,
        Y => S3530
    );
NAND_2292: ENTITY WORK.NAND
    PORT MAP (
        A => S3529,
        B => S3530,
        Y => S173
    );
NAND_2293: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_10,
        B => S3509,
        Y => S3531
    );
NAND_2294: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_170,
        B => S3510,
        Y => S3532
    );
NAND_2295: ENTITY WORK.NAND
    PORT MAP (
        A => S3531,
        B => S3532,
        Y => S174
    );
NAND_2296: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_11,
        B => S3509,
        Y => S3533
    );
NAND_2297: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_171,
        B => S3510,
        Y => S3534
    );
NAND_2298: ENTITY WORK.NAND
    PORT MAP (
        A => S3533,
        B => S3534,
        Y => S175
    );
NAND_2299: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_12,
        B => S3509,
        Y => S3535
    );
NAND_2300: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_172,
        B => S3510,
        Y => S3536
    );
NAND_2301: ENTITY WORK.NAND
    PORT MAP (
        A => S3535,
        B => S3536,
        Y => S176
    );
NAND_2302: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_13,
        B => S3509,
        Y => S3537
    );
NAND_2303: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_173,
        B => S3510,
        Y => S3538
    );
NAND_2304: ENTITY WORK.NAND
    PORT MAP (
        A => S3537,
        B => S3538,
        Y => S177
    );
NAND_2305: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_14,
        B => S3509,
        Y => S3539
    );
NAND_2306: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_174,
        B => S3510,
        Y => S3540
    );
NAND_2307: ENTITY WORK.NAND
    PORT MAP (
        A => S3539,
        B => S3540,
        Y => S178
    );
NAND_2308: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_15,
        B => S3509,
        Y => S3541
    );
NAND_2309: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_175,
        B => S3510,
        Y => S3542
    );
NAND_2310: ENTITY WORK.NAND
    PORT MAP (
        A => S3541,
        B => S3542,
        Y => S179
    );
NOR_943: ENTITY WORK.NOR
    PORT MAP (
        A => S3230,
        B => S3266,
        Y => S3543
    );
NAND_2311: ENTITY WORK.NAND
    PORT MAP (
        A => S3229,
        B => S3265,
        Y => S3544
    );
NAND_2312: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_0,
        B => S3543,
        Y => S3545
    );
NAND_2313: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_176,
        B => S3544,
        Y => S3546
    );
NAND_2314: ENTITY WORK.NAND
    PORT MAP (
        A => S3545,
        B => S3546,
        Y => S180
    );
NAND_2315: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_1,
        B => S3543,
        Y => S3547
    );
NAND_2316: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_177,
        B => S3544,
        Y => S3548
    );
NAND_2317: ENTITY WORK.NAND
    PORT MAP (
        A => S3547,
        B => S3548,
        Y => S181
    );
NAND_2318: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_2,
        B => S3543,
        Y => S3549
    );
NAND_2319: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_178,
        B => S3544,
        Y => S3550
    );
NAND_2320: ENTITY WORK.NAND
    PORT MAP (
        A => S3549,
        B => S3550,
        Y => S182
    );
NAND_2321: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_3,
        B => S3543,
        Y => S3551
    );
NAND_2322: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_179,
        B => S3544,
        Y => S3552
    );
NAND_2323: ENTITY WORK.NAND
    PORT MAP (
        A => S3551,
        B => S3552,
        Y => S183
    );
NAND_2324: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_4,
        B => S3543,
        Y => S3553
    );
NAND_2325: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_180,
        B => S3544,
        Y => S3554
    );
NAND_2326: ENTITY WORK.NAND
    PORT MAP (
        A => S3553,
        B => S3554,
        Y => S184
    );
NAND_2327: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_5,
        B => S3543,
        Y => S3555
    );
NAND_2328: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_181,
        B => S3544,
        Y => S3556
    );
NAND_2329: ENTITY WORK.NAND
    PORT MAP (
        A => S3555,
        B => S3556,
        Y => S185
    );
NAND_2330: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_6,
        B => S3543,
        Y => S3557
    );
NAND_2331: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_182,
        B => S3544,
        Y => S3558
    );
NAND_2332: ENTITY WORK.NAND
    PORT MAP (
        A => S3557,
        B => S3558,
        Y => S186
    );
NAND_2333: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_7,
        B => S3543,
        Y => S3559
    );
NAND_2334: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_183,
        B => S3544,
        Y => S3560
    );
NAND_2335: ENTITY WORK.NAND
    PORT MAP (
        A => S3559,
        B => S3560,
        Y => S187
    );
NAND_2336: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_8,
        B => S3543,
        Y => S3561
    );
NAND_2337: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_184,
        B => S3544,
        Y => S3562
    );
NAND_2338: ENTITY WORK.NAND
    PORT MAP (
        A => S3561,
        B => S3562,
        Y => S188
    );
NAND_2339: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_9,
        B => S3543,
        Y => S3563
    );
NAND_2340: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_185,
        B => S3544,
        Y => S3564
    );
NAND_2341: ENTITY WORK.NAND
    PORT MAP (
        A => S3563,
        B => S3564,
        Y => S189
    );
NAND_2342: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_10,
        B => S3543,
        Y => S3565
    );
NAND_2343: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_186,
        B => S3544,
        Y => S3566
    );
NAND_2344: ENTITY WORK.NAND
    PORT MAP (
        A => S3565,
        B => S3566,
        Y => S190
    );
NAND_2345: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_11,
        B => S3543,
        Y => S3567
    );
NAND_2346: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_187,
        B => S3544,
        Y => S3568
    );
NAND_2347: ENTITY WORK.NAND
    PORT MAP (
        A => S3567,
        B => S3568,
        Y => S191
    );
NAND_2348: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_12,
        B => S3543,
        Y => S3569
    );
NAND_2349: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_188,
        B => S3544,
        Y => S3570
    );
NAND_2350: ENTITY WORK.NAND
    PORT MAP (
        A => S3569,
        B => S3570,
        Y => S192
    );
NAND_2351: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_13,
        B => S3543,
        Y => S3571
    );
NAND_2352: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_189,
        B => S3544,
        Y => S3572
    );
NAND_2353: ENTITY WORK.NAND
    PORT MAP (
        A => S3571,
        B => S3572,
        Y => S193
    );
NAND_2354: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_14,
        B => S3543,
        Y => S3573
    );
NAND_2355: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_190,
        B => S3544,
        Y => S3574
    );
NAND_2356: ENTITY WORK.NAND
    PORT MAP (
        A => S3573,
        B => S3574,
        Y => S194
    );
NAND_2357: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_15,
        B => S3543,
        Y => S3575
    );
NAND_2358: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_191,
        B => S3544,
        Y => S3576
    );
NAND_2359: ENTITY WORK.NAND
    PORT MAP (
        A => S3575,
        B => S3576,
        Y => S195
    );
NOR_944: ENTITY WORK.NOR
    PORT MAP (
        A => S1654,
        B => S1661,
        Y => S3577
    );
NAND_2360: ENTITY WORK.NAND
    PORT MAP (
        A => S1655,
        B => S1662,
        Y => S3578
    );
NOR_945: ENTITY WORK.NOR
    PORT MAP (
        A => S1672,
        B => S3578,
        Y => S3579
    );
NAND_2361: ENTITY WORK.NAND
    PORT MAP (
        A => S1671,
        B => S3577,
        Y => S3580
    );
NOR_946: ENTITY WORK.NOR
    PORT MAP (
        A => S1687,
        B => S3580,
        Y => S3581
    );
NAND_2362: ENTITY WORK.NAND
    PORT MAP (
        A => S1686,
        B => S3579,
        Y => S3582
    );
NAND_2363: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_0,
        B => S3581,
        Y => S3583
    );
NAND_2364: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_192,
        B => S3582,
        Y => S3584
    );
NAND_2365: ENTITY WORK.NAND
    PORT MAP (
        A => S3583,
        B => S3584,
        Y => S196
    );
NAND_2366: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_1,
        B => S3581,
        Y => S3585
    );
NAND_2367: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_193,
        B => S3582,
        Y => S3586
    );
NAND_2368: ENTITY WORK.NAND
    PORT MAP (
        A => S3585,
        B => S3586,
        Y => S197
    );
NAND_2369: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_2,
        B => S3581,
        Y => S3587
    );
NAND_2370: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_194,
        B => S3582,
        Y => S3588
    );
NAND_2371: ENTITY WORK.NAND
    PORT MAP (
        A => S3587,
        B => S3588,
        Y => S198
    );
NAND_2372: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_3,
        B => S3581,
        Y => S3589
    );
NAND_2373: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_195,
        B => S3582,
        Y => S3590
    );
NAND_2374: ENTITY WORK.NAND
    PORT MAP (
        A => S3589,
        B => S3590,
        Y => S199
    );
NAND_2375: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_4,
        B => S3581,
        Y => S3591
    );
NAND_2376: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_196,
        B => S3582,
        Y => S3592
    );
NAND_2377: ENTITY WORK.NAND
    PORT MAP (
        A => S3591,
        B => S3592,
        Y => S200
    );
NAND_2378: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_5,
        B => S3581,
        Y => S3593
    );
NAND_2379: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_197,
        B => S3582,
        Y => S3594
    );
NAND_2380: ENTITY WORK.NAND
    PORT MAP (
        A => S3593,
        B => S3594,
        Y => S201
    );
NAND_2381: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_6,
        B => S3581,
        Y => S3595
    );
NAND_2382: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_198,
        B => S3582,
        Y => S3596
    );
NAND_2383: ENTITY WORK.NAND
    PORT MAP (
        A => S3595,
        B => S3596,
        Y => S202
    );
NAND_2384: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_7,
        B => S3581,
        Y => S3597
    );
NAND_2385: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_199,
        B => S3582,
        Y => S3598
    );
NAND_2386: ENTITY WORK.NAND
    PORT MAP (
        A => S3597,
        B => S3598,
        Y => S203
    );
NAND_2387: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_8,
        B => S3581,
        Y => S3599
    );
NAND_2388: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_200,
        B => S3582,
        Y => S3600
    );
NAND_2389: ENTITY WORK.NAND
    PORT MAP (
        A => S3599,
        B => S3600,
        Y => S204
    );
NAND_2390: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_9,
        B => S3581,
        Y => S3601
    );
NAND_2391: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_201,
        B => S3582,
        Y => S3602
    );
NAND_2392: ENTITY WORK.NAND
    PORT MAP (
        A => S3601,
        B => S3602,
        Y => S205
    );
NAND_2393: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_10,
        B => S3581,
        Y => S3603
    );
NAND_2394: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_202,
        B => S3582,
        Y => S3604
    );
NAND_2395: ENTITY WORK.NAND
    PORT MAP (
        A => S3603,
        B => S3604,
        Y => S206
    );
NAND_2396: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_11,
        B => S3581,
        Y => S3605
    );
NAND_2397: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_203,
        B => S3582,
        Y => S3606
    );
NAND_2398: ENTITY WORK.NAND
    PORT MAP (
        A => S3605,
        B => S3606,
        Y => S207
    );
NAND_2399: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_12,
        B => S3581,
        Y => S3607
    );
NAND_2400: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_204,
        B => S3582,
        Y => S3608
    );
NAND_2401: ENTITY WORK.NAND
    PORT MAP (
        A => S3607,
        B => S3608,
        Y => S208
    );
NAND_2402: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_13,
        B => S3581,
        Y => S3609
    );
NAND_2403: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_205,
        B => S3582,
        Y => S3610
    );
NAND_2404: ENTITY WORK.NAND
    PORT MAP (
        A => S3609,
        B => S3610,
        Y => S209
    );
NAND_2405: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_14,
        B => S3581,
        Y => S3611
    );
NAND_2406: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_206,
        B => S3582,
        Y => S3612
    );
NAND_2407: ENTITY WORK.NAND
    PORT MAP (
        A => S3611,
        B => S3612,
        Y => S210
    );
NAND_2408: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_15,
        B => S3581,
        Y => S3613
    );
NAND_2409: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_207,
        B => S3582,
        Y => S3614
    );
NAND_2410: ENTITY WORK.NAND
    PORT MAP (
        A => S3613,
        B => S3614,
        Y => S211
    );
NOR_947: ENTITY WORK.NOR
    PORT MAP (
        A => S3228,
        B => S3580,
        Y => S3615
    );
NAND_2411: ENTITY WORK.NAND
    PORT MAP (
        A => S3227,
        B => S3579,
        Y => S3616
    );
NAND_2412: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_0,
        B => S3615,
        Y => S3617
    );
NAND_2413: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_208,
        B => S3616,
        Y => S3618
    );
NAND_2414: ENTITY WORK.NAND
    PORT MAP (
        A => S3617,
        B => S3618,
        Y => S212
    );
NAND_2415: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_1,
        B => S3615,
        Y => S3619
    );
NAND_2416: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_209,
        B => S3616,
        Y => S3620
    );
NAND_2417: ENTITY WORK.NAND
    PORT MAP (
        A => S3619,
        B => S3620,
        Y => S213
    );
NAND_2418: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_2,
        B => S3615,
        Y => S3621
    );
NAND_2419: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_210,
        B => S3616,
        Y => S3622
    );
NAND_2420: ENTITY WORK.NAND
    PORT MAP (
        A => S3621,
        B => S3622,
        Y => S214
    );
NAND_2421: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_3,
        B => S3615,
        Y => S3623
    );
NAND_2422: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_211,
        B => S3616,
        Y => S3624
    );
NAND_2423: ENTITY WORK.NAND
    PORT MAP (
        A => S3623,
        B => S3624,
        Y => S215
    );
NAND_2424: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_4,
        B => S3615,
        Y => S3625
    );
NAND_2425: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_212,
        B => S3616,
        Y => S3626
    );
NAND_2426: ENTITY WORK.NAND
    PORT MAP (
        A => S3625,
        B => S3626,
        Y => S216
    );
NAND_2427: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_5,
        B => S3615,
        Y => S3627
    );
NAND_2428: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_213,
        B => S3616,
        Y => S3628
    );
NAND_2429: ENTITY WORK.NAND
    PORT MAP (
        A => S3627,
        B => S3628,
        Y => S217
    );
NAND_2430: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_6,
        B => S3615,
        Y => S3629
    );
NAND_2431: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_214,
        B => S3616,
        Y => S3630
    );
NAND_2432: ENTITY WORK.NAND
    PORT MAP (
        A => S3629,
        B => S3630,
        Y => S218
    );
NAND_2433: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_7,
        B => S3615,
        Y => S3631
    );
NAND_2434: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_215,
        B => S3616,
        Y => S3632
    );
NAND_2435: ENTITY WORK.NAND
    PORT MAP (
        A => S3631,
        B => S3632,
        Y => S219
    );
NAND_2436: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_8,
        B => S3615,
        Y => S3633
    );
NAND_2437: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_216,
        B => S3616,
        Y => S3634
    );
NAND_2438: ENTITY WORK.NAND
    PORT MAP (
        A => S3633,
        B => S3634,
        Y => S220
    );
NAND_2439: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_9,
        B => S3615,
        Y => S3635
    );
NAND_2440: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_217,
        B => S3616,
        Y => S3636
    );
NAND_2441: ENTITY WORK.NAND
    PORT MAP (
        A => S3635,
        B => S3636,
        Y => S221
    );
NAND_2442: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_10,
        B => S3615,
        Y => S3637
    );
NAND_2443: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_218,
        B => S3616,
        Y => S3638
    );
NAND_2444: ENTITY WORK.NAND
    PORT MAP (
        A => S3637,
        B => S3638,
        Y => S222
    );
NAND_2445: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_11,
        B => S3615,
        Y => S3639
    );
NAND_2446: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_219,
        B => S3616,
        Y => S3640
    );
NAND_2447: ENTITY WORK.NAND
    PORT MAP (
        A => S3639,
        B => S3640,
        Y => S223
    );
NAND_2448: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_12,
        B => S3615,
        Y => S3641
    );
NAND_2449: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_220,
        B => S3616,
        Y => S3642
    );
NAND_2450: ENTITY WORK.NAND
    PORT MAP (
        A => S3641,
        B => S3642,
        Y => S224
    );
NAND_2451: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_13,
        B => S3615,
        Y => S3643
    );
NAND_2452: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_221,
        B => S3616,
        Y => S3644
    );
NAND_2453: ENTITY WORK.NAND
    PORT MAP (
        A => S3643,
        B => S3644,
        Y => S225
    );
NAND_2454: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_14,
        B => S3615,
        Y => S3645
    );
NAND_2455: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_222,
        B => S3616,
        Y => S3646
    );
NAND_2456: ENTITY WORK.NAND
    PORT MAP (
        A => S3645,
        B => S3646,
        Y => S226
    );
NAND_2457: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_15,
        B => S3615,
        Y => S3647
    );
NAND_2458: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_223,
        B => S3616,
        Y => S3648
    );
NAND_2459: ENTITY WORK.NAND
    PORT MAP (
        A => S3647,
        B => S3648,
        Y => S227
    );
NOR_948: ENTITY WORK.NOR
    PORT MAP (
        A => S3192,
        B => S3578,
        Y => S3649
    );
NAND_2460: ENTITY WORK.NAND
    PORT MAP (
        A => S3191,
        B => S3577,
        Y => S3650
    );
NAND_2461: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_0,
        B => S3649,
        Y => S3651
    );
NAND_2462: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_224,
        B => S3650,
        Y => S3652
    );
NAND_2463: ENTITY WORK.NAND
    PORT MAP (
        A => S3651,
        B => S3652,
        Y => S228
    );
NAND_2464: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_1,
        B => S3649,
        Y => S3653
    );
NAND_2465: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_225,
        B => S3650,
        Y => S3654
    );
NAND_2466: ENTITY WORK.NAND
    PORT MAP (
        A => S3653,
        B => S3654,
        Y => S229
    );
NAND_2467: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_2,
        B => S3649,
        Y => S3655
    );
NAND_2468: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_226,
        B => S3650,
        Y => S3656
    );
NAND_2469: ENTITY WORK.NAND
    PORT MAP (
        A => S3655,
        B => S3656,
        Y => S230
    );
NAND_2470: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_3,
        B => S3649,
        Y => S3657
    );
NAND_2471: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_227,
        B => S3650,
        Y => S3658
    );
NAND_2472: ENTITY WORK.NAND
    PORT MAP (
        A => S3657,
        B => S3658,
        Y => S231
    );
NAND_2473: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_4,
        B => S3649,
        Y => S3659
    );
NAND_2474: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_228,
        B => S3650,
        Y => S3660
    );
NAND_2475: ENTITY WORK.NAND
    PORT MAP (
        A => S3659,
        B => S3660,
        Y => S232
    );
NAND_2476: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_5,
        B => S3649,
        Y => S3661
    );
NAND_2477: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_229,
        B => S3650,
        Y => S3662
    );
NAND_2478: ENTITY WORK.NAND
    PORT MAP (
        A => S3661,
        B => S3662,
        Y => S233
    );
NAND_2479: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_6,
        B => S3649,
        Y => S3663
    );
NAND_2480: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_230,
        B => S3650,
        Y => S3664
    );
NAND_2481: ENTITY WORK.NAND
    PORT MAP (
        A => S3663,
        B => S3664,
        Y => S234
    );
NAND_2482: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_7,
        B => S3649,
        Y => S3665
    );
NAND_2483: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_231,
        B => S3650,
        Y => S3666
    );
NAND_2484: ENTITY WORK.NAND
    PORT MAP (
        A => S3665,
        B => S3666,
        Y => S235
    );
NAND_2485: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_8,
        B => S3649,
        Y => S3667
    );
NAND_2486: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_232,
        B => S3650,
        Y => S3668
    );
NAND_2487: ENTITY WORK.NAND
    PORT MAP (
        A => S3667,
        B => S3668,
        Y => S236
    );
NAND_2488: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_9,
        B => S3649,
        Y => S3669
    );
NAND_2489: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_233,
        B => S3650,
        Y => S3670
    );
NAND_2490: ENTITY WORK.NAND
    PORT MAP (
        A => S3669,
        B => S3670,
        Y => S237
    );
NAND_2491: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_10,
        B => S3649,
        Y => S3671
    );
NAND_2492: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_234,
        B => S3650,
        Y => S3672
    );
NAND_2493: ENTITY WORK.NAND
    PORT MAP (
        A => S3671,
        B => S3672,
        Y => S238
    );
NAND_2494: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_11,
        B => S3649,
        Y => S3673
    );
NAND_2495: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_235,
        B => S3650,
        Y => S3674
    );
NAND_2496: ENTITY WORK.NAND
    PORT MAP (
        A => S3673,
        B => S3674,
        Y => S239
    );
NAND_2497: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_12,
        B => S3649,
        Y => S3675
    );
NAND_2498: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_236,
        B => S3650,
        Y => S3676
    );
NAND_2499: ENTITY WORK.NAND
    PORT MAP (
        A => S3675,
        B => S3676,
        Y => S240
    );
NAND_2500: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_13,
        B => S3649,
        Y => S3677
    );
NAND_2501: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_237,
        B => S3650,
        Y => S3678
    );
NAND_2502: ENTITY WORK.NAND
    PORT MAP (
        A => S3677,
        B => S3678,
        Y => S241
    );
NAND_2503: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_14,
        B => S3649,
        Y => S3679
    );
NAND_2504: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_238,
        B => S3650,
        Y => S3680
    );
NAND_2505: ENTITY WORK.NAND
    PORT MAP (
        A => S3679,
        B => S3680,
        Y => S242
    );
NAND_2506: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_indatatrf_15,
        B => S3649,
        Y => S3681
    );
NAND_2507: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_theregisterfile_memtrf_239,
        B => S3650,
        Y => S3682
    );
NAND_2508: ENTITY WORK.NAND
    PORT MAP (
        A => S3681,
        B => S3682,
        Y => S243
    );
NOR_949: ENTITY WORK.NOR
    PORT MAP (
        A => S1857,
        B => S1962,
        Y => S3683
    );
NOT_318: ENTITY WORK.NOT
    PORT MAP (
        A => S3683,
        Y => S3684
    );
NOR_950: ENTITY WORK.NOR
    PORT MAP (
        A => S3046,
        B => S3150,
        Y => S3685
    );
NAND_2509: ENTITY WORK.NAND
    PORT MAP (
        A => S2824,
        B => S3685,
        Y => S3686
    );
NOR_951: ENTITY WORK.NOR
    PORT MAP (
        A => S2929,
        B => S3686,
        Y => S3687
    );
NAND_2510: ENTITY WORK.NAND
    PORT MAP (
        A => S2626,
        B => S2724,
        Y => S3688
    );
NOT_319: ENTITY WORK.NOT
    PORT MAP (
        A => S3688,
        Y => S3689
    );
NOR_952: ENTITY WORK.NOR
    PORT MAP (
        A => S2424,
        B => S3688,
        Y => S3690
    );
NOT_320: ENTITY WORK.NOT
    PORT MAP (
        A => S3690,
        Y => S3691
    );
NAND_2511: ENTITY WORK.NAND
    PORT MAP (
        A => S2525,
        B => S3687,
        Y => S3692
    );
NOR_953: ENTITY WORK.NOR
    PORT MAP (
        A => S3691,
        B => S3692,
        Y => S3693
    );
NOR_954: ENTITY WORK.NOR
    PORT MAP (
        A => S2011,
        B => S2113,
        Y => S3694
    );
NAND_2512: ENTITY WORK.NAND
    PORT MAP (
        A => S1754,
        B => S3694,
        Y => S3695
    );
NAND_2513: ENTITY WORK.NAND
    PORT MAP (
        A => S1522,
        B => S3683,
        Y => S3696
    );
NOR_955: ENTITY WORK.NOR
    PORT MAP (
        A => S3695,
        B => S3696,
        Y => S3697
    );
NAND_2514: ENTITY WORK.NAND
    PORT MAP (
        A => S3693,
        B => S3697,
        Y => S3698
    );
NOR_956: ENTITY WORK.NOR
    PORT MAP (
        A => S2435,
        B => S3698,
        Y => S3699
    );
NOR_957: ENTITY WORK.NOR
    PORT MAP (
        A => S1405,
        B => S3699,
        Y => S3700
    );
NOR_958: ENTITY WORK.NOR
    PORT MAP (
        A => controller_389_B_0,
        B => S1404,
        Y => S3701
    );
NOR_959: ENTITY WORK.NOR
    PORT MAP (
        A => S3700,
        B => S3701,
        Y => S264
    );
NAND_2515: ENTITY WORK.NAND
    PORT MAP (
        A => controller_389_B_2,
        B => S1405,
        Y => S3702
    );
NAND_2516: ENTITY WORK.NAND
    PORT MAP (
        A => S2211,
        B => S2319,
        Y => S3703
    );
NOR_960: ENTITY WORK.NOR
    PORT MAP (
        A => S1853,
        B => S1958,
        Y => S3704
    );
NOR_961: ENTITY WORK.NOR
    PORT MAP (
        A => S1957,
        B => S3704,
        Y => S3705
    );
NAND_2517: ENTITY WORK.NAND
    PORT MAP (
        A => S1521,
        B => S1752,
        Y => S3706
    );
NAND_2518: ENTITY WORK.NAND
    PORT MAP (
        A => S1751,
        B => S3706,
        Y => S3707
    );
NOR_962: ENTITY WORK.NOR
    PORT MAP (
        A => S3684,
        B => S3707,
        Y => S3708
    );
NOR_963: ENTITY WORK.NOR
    PORT MAP (
        A => S3705,
        B => S3708,
        Y => S3709
    );
NOR_964: ENTITY WORK.NOR
    PORT MAP (
        A => S2007,
        B => S3709,
        Y => S3710
    );
NAND_2519: ENTITY WORK.NAND
    PORT MAP (
        A => S2010,
        B => S2112,
        Y => S3711
    );
NOR_965: ENTITY WORK.NOR
    PORT MAP (
        A => S3710,
        B => S3711,
        Y => S3712
    );
NOR_966: ENTITY WORK.NOR
    PORT MAP (
        A => S2435,
        B => S3712,
        Y => S3713
    );
NAND_2520: ENTITY WORK.NAND
    PORT MAP (
        A => S2111,
        B => S3713,
        Y => S3714
    );
NAND_2521: ENTITY WORK.NAND
    PORT MAP (
        A => S2317,
        B => S3703,
        Y => S3715
    );
NAND_2522: ENTITY WORK.NAND
    PORT MAP (
        A => S3714,
        B => S3715,
        Y => S3716
    );
NAND_2523: ENTITY WORK.NAND
    PORT MAP (
        A => S3693,
        B => S3716,
        Y => S3717
    );
NOT_321: ENTITY WORK.NOT
    PORT MAP (
        A => S3717,
        Y => S3718
    );
NOR_967: ENTITY WORK.NOR
    PORT MAP (
        A => S2422,
        B => S2524,
        Y => S3719
    );
NOR_968: ENTITY WORK.NOR
    PORT MAP (
        A => S2523,
        B => S3719,
        Y => S3720
    );
NAND_2524: ENTITY WORK.NAND
    PORT MAP (
        A => S3689,
        B => S3720,
        Y => S3721
    );
NOR_969: ENTITY WORK.NOR
    PORT MAP (
        A => S2622,
        B => S2722,
        Y => S3722
    );
NOR_970: ENTITY WORK.NOR
    PORT MAP (
        A => S2723,
        B => S3722,
        Y => S3723
    );
NAND_2525: ENTITY WORK.NAND
    PORT MAP (
        A => S3721,
        B => S3723,
        Y => S3724
    );
NAND_2526: ENTITY WORK.NAND
    PORT MAP (
        A => S3687,
        B => S3724,
        Y => S3725
    );
NOR_971: ENTITY WORK.NOR
    PORT MAP (
        A => S2823,
        B => S2927,
        Y => S3726
    );
NOR_972: ENTITY WORK.NOR
    PORT MAP (
        A => S2925,
        B => S3726,
        Y => S3727
    );
NAND_2527: ENTITY WORK.NAND
    PORT MAP (
        A => S3685,
        B => S3727,
        Y => S3728
    );
NOR_973: ENTITY WORK.NOR
    PORT MAP (
        A => S3043,
        B => S3148,
        Y => S3729
    );
NOR_974: ENTITY WORK.NOR
    PORT MAP (
        A => S3146,
        B => S3729,
        Y => S3730
    );
NAND_2528: ENTITY WORK.NAND
    PORT MAP (
        A => S3728,
        B => S3730,
        Y => S3731
    );
NOR_975: ENTITY WORK.NOR
    PORT MAP (
        A => S3718,
        B => S3731,
        Y => S3732
    );
NAND_2529: ENTITY WORK.NAND
    PORT MAP (
        A => S3725,
        B => S3732,
        Y => S3733
    );
NAND_2530: ENTITY WORK.NAND
    PORT MAP (
        A => S3700,
        B => S3733,
        Y => S3734
    );
NAND_2531: ENTITY WORK.NAND
    PORT MAP (
        A => S3702,
        B => S3734,
        Y => S265
    );
NAND_2532: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_0,
        B => S8580,
        Y => S3735
    );
NOR_976: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_muxmem_in2_0,
        B => S1222,
        Y => S3736
    );
NOR_977: ENTITY WORK.NOR
    PORT MAP (
        A => S364,
        B => S3736,
        Y => S3737
    );
NAND_2533: ENTITY WORK.NAND
    PORT MAP (
        A => S1223,
        B => S3737,
        Y => S3738
    );
NOR_978: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_muxmem_in2_0,
        B => S1334,
        Y => S3739
    );
NOR_979: ENTITY WORK.NOR
    PORT MAP (
        A => S1370,
        B => S3739,
        Y => S3740
    );
NAND_2534: ENTITY WORK.NAND
    PORT MAP (
        A => S3738,
        B => S3740,
        Y => S3741
    );
NOR_980: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_0,
        B => S1371,
        Y => S3742
    );
NOR_981: ENTITY WORK.NOR
    PORT MAP (
        A => S8580,
        B => S3742,
        Y => S3743
    );
NAND_2535: ENTITY WORK.NAND
    PORT MAP (
        A => S3741,
        B => S3743,
        Y => S3744
    );
NAND_2536: ENTITY WORK.NAND
    PORT MAP (
        A => S3735,
        B => S3744,
        Y => S267
    );
NAND_2537: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_1,
        B => S8580,
        Y => S3745
    );
NOR_982: ENTITY WORK.NOR
    PORT MAP (
        A => S1224,
        B => S1226,
        Y => S3746
    );
NOR_983: ENTITY WORK.NOR
    PORT MAP (
        A => S1228,
        B => S3746,
        Y => S3747
    );
NAND_2538: ENTITY WORK.NAND
    PORT MAP (
        A => S365,
        B => S3747,
        Y => S3748
    );
NOR_984: ENTITY WORK.NOR
    PORT MAP (
        A => S1334,
        B => S1774,
        Y => S3749
    );
NOR_985: ENTITY WORK.NOR
    PORT MAP (
        A => S1370,
        B => S3749,
        Y => S3750
    );
NAND_2539: ENTITY WORK.NAND
    PORT MAP (
        A => S3748,
        B => S3750,
        Y => S3751
    );
NOR_986: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_1,
        B => S1371,
        Y => S3752
    );
NOR_987: ENTITY WORK.NOR
    PORT MAP (
        A => S8580,
        B => S3752,
        Y => S3753
    );
NAND_2540: ENTITY WORK.NAND
    PORT MAP (
        A => S3751,
        B => S3753,
        Y => S3754
    );
NAND_2541: ENTITY WORK.NAND
    PORT MAP (
        A => S3745,
        B => S3754,
        Y => S268
    );
NAND_2542: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_2,
        B => S8580,
        Y => S3755
    );
NOR_988: ENTITY WORK.NOR
    PORT MAP (
        A => S1229,
        B => S1231,
        Y => S3756
    );
NOR_989: ENTITY WORK.NOR
    PORT MAP (
        A => S364,
        B => S3756,
        Y => S3757
    );
NAND_2543: ENTITY WORK.NAND
    PORT MAP (
        A => S1232,
        B => S3757,
        Y => S3758
    );
NOR_990: ENTITY WORK.NOR
    PORT MAP (
        A => S1334,
        B => S1875,
        Y => S3759
    );
NOR_991: ENTITY WORK.NOR
    PORT MAP (
        A => S1370,
        B => S3759,
        Y => S3760
    );
NAND_2544: ENTITY WORK.NAND
    PORT MAP (
        A => S3758,
        B => S3760,
        Y => S3761
    );
NOR_992: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_2,
        B => S1371,
        Y => S3762
    );
NOR_993: ENTITY WORK.NOR
    PORT MAP (
        A => S8580,
        B => S3762,
        Y => S3763
    );
NAND_2545: ENTITY WORK.NAND
    PORT MAP (
        A => S3761,
        B => S3763,
        Y => S3764
    );
NAND_2546: ENTITY WORK.NAND
    PORT MAP (
        A => S3755,
        B => S3764,
        Y => S269
    );
NAND_2547: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_3,
        B => S8580,
        Y => S3765
    );
NOR_994: ENTITY WORK.NOR
    PORT MAP (
        A => S1069,
        B => S1070,
        Y => S3766
    );
NAND_2548: ENTITY WORK.NAND
    PORT MAP (
        A => S1233,
        B => S3766,
        Y => S3767
    );
NOR_995: ENTITY WORK.NOR
    PORT MAP (
        A => S1233,
        B => S3766,
        Y => S3768
    );
NOR_996: ENTITY WORK.NOR
    PORT MAP (
        A => S364,
        B => S3768,
        Y => S3769
    );
NAND_2549: ENTITY WORK.NAND
    PORT MAP (
        A => S3767,
        B => S3769,
        Y => S3770
    );
NOR_997: ENTITY WORK.NOR
    PORT MAP (
        A => S1334,
        B => S1978,
        Y => S3771
    );
NOR_998: ENTITY WORK.NOR
    PORT MAP (
        A => S1370,
        B => S3771,
        Y => S3772
    );
NAND_2550: ENTITY WORK.NAND
    PORT MAP (
        A => S3770,
        B => S3772,
        Y => S3773
    );
NOR_999: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_3,
        B => S1371,
        Y => S3774
    );
NOR_1000: ENTITY WORK.NOR
    PORT MAP (
        A => S8580,
        B => S3774,
        Y => S3775
    );
NAND_2551: ENTITY WORK.NAND
    PORT MAP (
        A => S3773,
        B => S3775,
        Y => S3776
    );
NAND_2552: ENTITY WORK.NAND
    PORT MAP (
        A => S3765,
        B => S3776,
        Y => S270
    );
NAND_2553: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_4,
        B => S8580,
        Y => S3777
    );
NOR_1001: ENTITY WORK.NOR
    PORT MAP (
        A => S1019,
        B => S1235,
        Y => S3778
    );
NOR_1002: ENTITY WORK.NOR
    PORT MAP (
        A => S1334,
        B => S2029,
        Y => S3779
    );
NOR_1003: ENTITY WORK.NOR
    PORT MAP (
        A => S364,
        B => S3778,
        Y => S3780
    );
NAND_2554: ENTITY WORK.NAND
    PORT MAP (
        A => S1236,
        B => S3780,
        Y => S3781
    );
NOT_322: ENTITY WORK.NOT
    PORT MAP (
        A => S3781,
        Y => S3782
    );
NOR_1004: ENTITY WORK.NOR
    PORT MAP (
        A => S3779,
        B => S3782,
        Y => S3783
    );
NAND_2555: ENTITY WORK.NAND
    PORT MAP (
        A => S1371,
        B => S3783,
        Y => S3784
    );
NOR_1005: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_4,
        B => S1371,
        Y => S3785
    );
NOR_1006: ENTITY WORK.NOR
    PORT MAP (
        A => S8580,
        B => S3785,
        Y => S3786
    );
NAND_2556: ENTITY WORK.NAND
    PORT MAP (
        A => S3784,
        B => S3786,
        Y => S3787
    );
NAND_2557: ENTITY WORK.NAND
    PORT MAP (
        A => S3777,
        B => S3787,
        Y => S271
    );
NAND_2558: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_5,
        B => S8580,
        Y => S3788
    );
NOR_1007: ENTITY WORK.NOR
    PORT MAP (
        A => S967,
        B => S968,
        Y => S3789
    );
NAND_2559: ENTITY WORK.NAND
    PORT MAP (
        A => S1237,
        B => S3789,
        Y => S3790
    );
NOR_1008: ENTITY WORK.NOR
    PORT MAP (
        A => S1237,
        B => S3789,
        Y => S3791
    );
NOR_1009: ENTITY WORK.NOR
    PORT MAP (
        A => S364,
        B => S3791,
        Y => S3792
    );
NAND_2560: ENTITY WORK.NAND
    PORT MAP (
        A => S3790,
        B => S3792,
        Y => S3793
    );
NOR_1010: ENTITY WORK.NOR
    PORT MAP (
        A => S1334,
        B => S2136,
        Y => S3794
    );
NOR_1011: ENTITY WORK.NOR
    PORT MAP (
        A => S1370,
        B => S3794,
        Y => S3795
    );
NAND_2561: ENTITY WORK.NAND
    PORT MAP (
        A => S3793,
        B => S3795,
        Y => S3796
    );
NOR_1012: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_5,
        B => S1371,
        Y => S3797
    );
NOR_1013: ENTITY WORK.NOR
    PORT MAP (
        A => S8580,
        B => S3797,
        Y => S3798
    );
NAND_2562: ENTITY WORK.NAND
    PORT MAP (
        A => S3796,
        B => S3798,
        Y => S3799
    );
NAND_2563: ENTITY WORK.NAND
    PORT MAP (
        A => S3788,
        B => S3799,
        Y => S272
    );
NAND_2564: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_6,
        B => S8580,
        Y => S3800
    );
NOR_1014: ENTITY WORK.NOR
    PORT MAP (
        A => S916,
        B => S1239,
        Y => S3801
    );
NOR_1015: ENTITY WORK.NOR
    PORT MAP (
        A => S364,
        B => S3801,
        Y => S3802
    );
NAND_2565: ENTITY WORK.NAND
    PORT MAP (
        A => S1240,
        B => S3802,
        Y => S3803
    );
NOR_1016: ENTITY WORK.NOR
    PORT MAP (
        A => S1334,
        B => S2235,
        Y => S3804
    );
NOR_1017: ENTITY WORK.NOR
    PORT MAP (
        A => S1370,
        B => S3804,
        Y => S3805
    );
NAND_2566: ENTITY WORK.NAND
    PORT MAP (
        A => S3803,
        B => S3805,
        Y => S3806
    );
NOR_1018: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_6,
        B => S1371,
        Y => S3807
    );
NOR_1019: ENTITY WORK.NOR
    PORT MAP (
        A => S8580,
        B => S3807,
        Y => S3808
    );
NAND_2567: ENTITY WORK.NAND
    PORT MAP (
        A => S3806,
        B => S3808,
        Y => S3809
    );
NAND_2568: ENTITY WORK.NAND
    PORT MAP (
        A => S3800,
        B => S3809,
        Y => S273
    );
NAND_2569: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_7,
        B => S8580,
        Y => S3810
    );
NOR_1020: ENTITY WORK.NOR
    PORT MAP (
        A => S862,
        B => S863,
        Y => S3811
    );
NAND_2570: ENTITY WORK.NAND
    PORT MAP (
        A => S1241,
        B => S3811,
        Y => S3812
    );
NOR_1021: ENTITY WORK.NOR
    PORT MAP (
        A => S1241,
        B => S3811,
        Y => S3813
    );
NOR_1022: ENTITY WORK.NOR
    PORT MAP (
        A => S364,
        B => S3813,
        Y => S3814
    );
NAND_2571: ENTITY WORK.NAND
    PORT MAP (
        A => S3812,
        B => S3814,
        Y => S3815
    );
NOR_1023: ENTITY WORK.NOR
    PORT MAP (
        A => S1334,
        B => S2331,
        Y => S3816
    );
NOR_1024: ENTITY WORK.NOR
    PORT MAP (
        A => S1370,
        B => S3816,
        Y => S3817
    );
NAND_2572: ENTITY WORK.NAND
    PORT MAP (
        A => S3815,
        B => S3817,
        Y => S3818
    );
NOR_1025: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_7,
        B => S1371,
        Y => S3819
    );
NOR_1026: ENTITY WORK.NOR
    PORT MAP (
        A => S8580,
        B => S3819,
        Y => S3820
    );
NAND_2573: ENTITY WORK.NAND
    PORT MAP (
        A => S3818,
        B => S3820,
        Y => S3821
    );
NAND_2574: ENTITY WORK.NAND
    PORT MAP (
        A => S3810,
        B => S3821,
        Y => S274
    );
NAND_2575: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_8,
        B => S8580,
        Y => S3822
    );
NOR_1027: ENTITY WORK.NOR
    PORT MAP (
        A => S811,
        B => S1243,
        Y => S3823
    );
NOR_1028: ENTITY WORK.NOR
    PORT MAP (
        A => S364,
        B => S3823,
        Y => S3824
    );
NAND_2576: ENTITY WORK.NAND
    PORT MAP (
        A => S1244,
        B => S3824,
        Y => S3825
    );
NOR_1029: ENTITY WORK.NOR
    PORT MAP (
        A => S1334,
        B => S2449,
        Y => S3826
    );
NOR_1030: ENTITY WORK.NOR
    PORT MAP (
        A => S1370,
        B => S3826,
        Y => S3827
    );
NAND_2577: ENTITY WORK.NAND
    PORT MAP (
        A => S3825,
        B => S3827,
        Y => S3828
    );
NOR_1031: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_8,
        B => S1371,
        Y => S3829
    );
NOR_1032: ENTITY WORK.NOR
    PORT MAP (
        A => S8580,
        B => S3829,
        Y => S3830
    );
NAND_2578: ENTITY WORK.NAND
    PORT MAP (
        A => S3828,
        B => S3830,
        Y => S3831
    );
NAND_2579: ENTITY WORK.NAND
    PORT MAP (
        A => S3822,
        B => S3831,
        Y => S275
    );
NAND_2580: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_9,
        B => S8580,
        Y => S3832
    );
NOR_1033: ENTITY WORK.NOR
    PORT MAP (
        A => S758,
        B => S759,
        Y => S3833
    );
NAND_2581: ENTITY WORK.NAND
    PORT MAP (
        A => S1245,
        B => S3833,
        Y => S3834
    );
NOR_1034: ENTITY WORK.NOR
    PORT MAP (
        A => S1245,
        B => S3833,
        Y => S3835
    );
NOR_1035: ENTITY WORK.NOR
    PORT MAP (
        A => S364,
        B => S3835,
        Y => S3836
    );
NAND_2582: ENTITY WORK.NAND
    PORT MAP (
        A => S3834,
        B => S3836,
        Y => S3837
    );
NOR_1036: ENTITY WORK.NOR
    PORT MAP (
        A => S1334,
        B => S2551,
        Y => S3838
    );
NOR_1037: ENTITY WORK.NOR
    PORT MAP (
        A => S1370,
        B => S3838,
        Y => S3839
    );
NAND_2583: ENTITY WORK.NAND
    PORT MAP (
        A => S3837,
        B => S3839,
        Y => S3840
    );
NOR_1038: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_9,
        B => S1371,
        Y => S3841
    );
NOR_1039: ENTITY WORK.NOR
    PORT MAP (
        A => S8580,
        B => S3841,
        Y => S3842
    );
NAND_2584: ENTITY WORK.NAND
    PORT MAP (
        A => S3840,
        B => S3842,
        Y => S3843
    );
NAND_2585: ENTITY WORK.NAND
    PORT MAP (
        A => S3832,
        B => S3843,
        Y => S276
    );
NAND_2586: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_10,
        B => S8580,
        Y => S3844
    );
NOR_1040: ENTITY WORK.NOR
    PORT MAP (
        A => S708,
        B => S1247,
        Y => S3845
    );
NOR_1041: ENTITY WORK.NOR
    PORT MAP (
        A => S364,
        B => S3845,
        Y => S3846
    );
NAND_2587: ENTITY WORK.NAND
    PORT MAP (
        A => S1248,
        B => S3846,
        Y => S3847
    );
NOR_1042: ENTITY WORK.NOR
    PORT MAP (
        A => S1334,
        B => S2646,
        Y => S3848
    );
NOR_1043: ENTITY WORK.NOR
    PORT MAP (
        A => S1370,
        B => S3848,
        Y => S3849
    );
NAND_2588: ENTITY WORK.NAND
    PORT MAP (
        A => S3847,
        B => S3849,
        Y => S3850
    );
NOR_1044: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_10,
        B => S1371,
        Y => S3851
    );
NOR_1045: ENTITY WORK.NOR
    PORT MAP (
        A => S8580,
        B => S3851,
        Y => S3852
    );
NAND_2589: ENTITY WORK.NAND
    PORT MAP (
        A => S3850,
        B => S3852,
        Y => S3853
    );
NAND_2590: ENTITY WORK.NAND
    PORT MAP (
        A => S3844,
        B => S3853,
        Y => S277
    );
NAND_2591: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_11,
        B => S8580,
        Y => S3854
    );
NOR_1046: ENTITY WORK.NOR
    PORT MAP (
        A => S655,
        B => S656,
        Y => S3855
    );
NAND_2592: ENTITY WORK.NAND
    PORT MAP (
        A => S1249,
        B => S3855,
        Y => S3856
    );
NOR_1047: ENTITY WORK.NOR
    PORT MAP (
        A => S1249,
        B => S3855,
        Y => S3857
    );
NOR_1048: ENTITY WORK.NOR
    PORT MAP (
        A => S364,
        B => S3857,
        Y => S3858
    );
NAND_2593: ENTITY WORK.NAND
    PORT MAP (
        A => S3856,
        B => S3858,
        Y => S3859
    );
NOR_1049: ENTITY WORK.NOR
    PORT MAP (
        A => S1334,
        B => S2748,
        Y => S3860
    );
NOR_1050: ENTITY WORK.NOR
    PORT MAP (
        A => S1370,
        B => S3860,
        Y => S3861
    );
NAND_2594: ENTITY WORK.NAND
    PORT MAP (
        A => S3859,
        B => S3861,
        Y => S3862
    );
NOR_1051: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_11,
        B => S1371,
        Y => S3863
    );
NOR_1052: ENTITY WORK.NOR
    PORT MAP (
        A => S8580,
        B => S3863,
        Y => S3864
    );
NAND_2595: ENTITY WORK.NAND
    PORT MAP (
        A => S3862,
        B => S3864,
        Y => S3865
    );
NAND_2596: ENTITY WORK.NAND
    PORT MAP (
        A => S3854,
        B => S3865,
        Y => S278
    );
NAND_2597: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_12,
        B => S8580,
        Y => S3866
    );
NOR_1053: ENTITY WORK.NOR
    PORT MAP (
        A => S605,
        B => S1251,
        Y => S3867
    );
NOR_1054: ENTITY WORK.NOR
    PORT MAP (
        A => S364,
        B => S3867,
        Y => S3868
    );
NAND_2598: ENTITY WORK.NAND
    PORT MAP (
        A => S1252,
        B => S3868,
        Y => S3869
    );
NOR_1055: ENTITY WORK.NOR
    PORT MAP (
        A => S1334,
        B => S2847,
        Y => S3870
    );
NOR_1056: ENTITY WORK.NOR
    PORT MAP (
        A => S1370,
        B => S3870,
        Y => S3871
    );
NAND_2599: ENTITY WORK.NAND
    PORT MAP (
        A => S3869,
        B => S3871,
        Y => S3872
    );
NOR_1057: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_12,
        B => S1371,
        Y => S3873
    );
NOR_1058: ENTITY WORK.NOR
    PORT MAP (
        A => S8580,
        B => S3873,
        Y => S3874
    );
NAND_2600: ENTITY WORK.NAND
    PORT MAP (
        A => S3872,
        B => S3874,
        Y => S3875
    );
NAND_2601: ENTITY WORK.NAND
    PORT MAP (
        A => S3866,
        B => S3875,
        Y => S279
    );
NAND_2602: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_13,
        B => S8580,
        Y => S3876
    );
NOR_1059: ENTITY WORK.NOR
    PORT MAP (
        A => S552,
        B => S553,
        Y => S3877
    );
NAND_2603: ENTITY WORK.NAND
    PORT MAP (
        A => S1253,
        B => S3877,
        Y => S3878
    );
NOR_1060: ENTITY WORK.NOR
    PORT MAP (
        A => S1253,
        B => S3877,
        Y => S3879
    );
NOR_1061: ENTITY WORK.NOR
    PORT MAP (
        A => S364,
        B => S3879,
        Y => S3880
    );
NAND_2604: ENTITY WORK.NAND
    PORT MAP (
        A => S3878,
        B => S3880,
        Y => S3881
    );
NOR_1062: ENTITY WORK.NOR
    PORT MAP (
        A => S1334,
        B => S2956,
        Y => S3882
    );
NOR_1063: ENTITY WORK.NOR
    PORT MAP (
        A => S1370,
        B => S3882,
        Y => S3883
    );
NAND_2605: ENTITY WORK.NAND
    PORT MAP (
        A => S3881,
        B => S3883,
        Y => S3884
    );
NOR_1064: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_13,
        B => S1371,
        Y => S3885
    );
NOR_1065: ENTITY WORK.NOR
    PORT MAP (
        A => S8580,
        B => S3885,
        Y => S3886
    );
NAND_2606: ENTITY WORK.NAND
    PORT MAP (
        A => S3884,
        B => S3886,
        Y => S3887
    );
NAND_2607: ENTITY WORK.NAND
    PORT MAP (
        A => S3876,
        B => S3887,
        Y => S280
    );
NAND_2608: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_14,
        B => S8580,
        Y => S3888
    );
NOR_1066: ENTITY WORK.NOR
    PORT MAP (
        A => S502,
        B => S1255,
        Y => S3889
    );
NOR_1067: ENTITY WORK.NOR
    PORT MAP (
        A => S364,
        B => S3889,
        Y => S3890
    );
NAND_2609: ENTITY WORK.NAND
    PORT MAP (
        A => S1256,
        B => S3890,
        Y => S3891
    );
NOR_1068: ENTITY WORK.NOR
    PORT MAP (
        A => S1334,
        B => S3066,
        Y => S3892
    );
NOR_1069: ENTITY WORK.NOR
    PORT MAP (
        A => S1370,
        B => S3892,
        Y => S3893
    );
NAND_2610: ENTITY WORK.NAND
    PORT MAP (
        A => S3891,
        B => S3893,
        Y => S3894
    );
NOR_1070: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_14,
        B => S1371,
        Y => S3895
    );
NOR_1071: ENTITY WORK.NOR
    PORT MAP (
        A => S8580,
        B => S3895,
        Y => S3896
    );
NAND_2611: ENTITY WORK.NAND
    PORT MAP (
        A => S3894,
        B => S3896,
        Y => S3897
    );
NAND_2612: ENTITY WORK.NAND
    PORT MAP (
        A => S3888,
        B => S3897,
        Y => S281
    );
NOR_1072: ENTITY WORK.NOR
    PORT MAP (
        A => S8557,
        B => S377,
        Y => S3898
    );
NAND_2613: ENTITY WORK.NAND
    PORT MAP (
        A => S8556,
        B => S376,
        Y => S3899
    );
NOR_1073: ENTITY WORK.NOR
    PORT MAP (
        A => S3036,
        B => S3141,
        Y => S3900
    );
NAND_2614: ENTITY WORK.NAND
    PORT MAP (
        A => S3037,
        B => S3142,
        Y => S3901
    );
NOR_1074: ENTITY WORK.NOR
    PORT MAP (
        A => S2919,
        B => S3901,
        Y => S3902
    );
NAND_2615: ENTITY WORK.NAND
    PORT MAP (
        A => S2920,
        B => S3900,
        Y => S3903
    );
NOR_1075: ENTITY WORK.NOR
    PORT MAP (
        A => S2816,
        B => S3903,
        Y => S3904
    );
NAND_2616: ENTITY WORK.NAND
    PORT MAP (
        A => S2817,
        B => S3902,
        Y => S3905
    );
NOR_1076: ENTITY WORK.NOR
    PORT MAP (
        A => S2717,
        B => S3905,
        Y => S3906
    );
NAND_2617: ENTITY WORK.NAND
    PORT MAP (
        A => S2718,
        B => S3904,
        Y => S3907
    );
NOR_1077: ENTITY WORK.NOR
    PORT MAP (
        A => S2617,
        B => S3907,
        Y => S3908
    );
NAND_2618: ENTITY WORK.NAND
    PORT MAP (
        A => S2618,
        B => S3906,
        Y => S3909
    );
NOR_1078: ENTITY WORK.NOR
    PORT MAP (
        A => S2517,
        B => S3909,
        Y => S3910
    );
NAND_2619: ENTITY WORK.NAND
    PORT MAP (
        A => S2518,
        B => S3908,
        Y => S3911
    );
NOR_1079: ENTITY WORK.NOR
    PORT MAP (
        A => S2417,
        B => S3911,
        Y => S3912
    );
NAND_2620: ENTITY WORK.NAND
    PORT MAP (
        A => S2418,
        B => S3910,
        Y => S3913
    );
NOR_1080: ENTITY WORK.NOR
    PORT MAP (
        A => S2311,
        B => S3913,
        Y => S3914
    );
NAND_2621: ENTITY WORK.NAND
    PORT MAP (
        A => S2312,
        B => S3912,
        Y => S3915
    );
NOR_1081: ENTITY WORK.NOR
    PORT MAP (
        A => S2205,
        B => S3915,
        Y => S3916
    );
NAND_2622: ENTITY WORK.NAND
    PORT MAP (
        A => S2206,
        B => S3914,
        Y => S3917
    );
NOR_1082: ENTITY WORK.NOR
    PORT MAP (
        A => S2106,
        B => S3917,
        Y => S3918
    );
NAND_2623: ENTITY WORK.NAND
    PORT MAP (
        A => S2107,
        B => S3916,
        Y => S3919
    );
NOR_1083: ENTITY WORK.NOR
    PORT MAP (
        A => S1597,
        B => S3919,
        Y => S3920
    );
NAND_2624: ENTITY WORK.NAND
    PORT MAP (
        A => S1598,
        B => S3918,
        Y => S3921
    );
NOR_1084: ENTITY WORK.NOR
    PORT MAP (
        A => S1952,
        B => S3921,
        Y => S3922
    );
NAND_2625: ENTITY WORK.NAND
    PORT MAP (
        A => S1953,
        B => S3920,
        Y => S3923
    );
NOR_1085: ENTITY WORK.NOR
    PORT MAP (
        A => S1848,
        B => S3923,
        Y => S3924
    );
NAND_2626: ENTITY WORK.NAND
    PORT MAP (
        A => S1849,
        B => S3922,
        Y => S3925
    );
NOR_1086: ENTITY WORK.NOR
    PORT MAP (
        A => S1745,
        B => S3925,
        Y => S3926
    );
NAND_2627: ENTITY WORK.NAND
    PORT MAP (
        A => S1746,
        B => S3924,
        Y => S3927
    );
NOR_1087: ENTITY WORK.NOR
    PORT MAP (
        A => S1516,
        B => S3927,
        Y => S3928
    );
NAND_2628: ENTITY WORK.NAND
    PORT MAP (
        A => S1515,
        B => S3926,
        Y => S3929
    );
NOR_1088: ENTITY WORK.NOR
    PORT MAP (
        A => S1304,
        B => S3928,
        Y => S3930
    );
NAND_2629: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_15,
        B => S3929,
        Y => S3931
    );
NOR_1089: ENTITY WORK.NOR
    PORT MAP (
        A => S1745,
        B => S3931,
        Y => S3932
    );
NAND_2630: ENTITY WORK.NAND
    PORT MAP (
        A => S1746,
        B => S3930,
        Y => S3933
    );
NOR_1090: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_15,
        B => S1746,
        Y => S3934
    );
NAND_2631: ENTITY WORK.NAND
    PORT MAP (
        A => S1304,
        B => S1745,
        Y => S3935
    );
NOR_1091: ENTITY WORK.NOR
    PORT MAP (
        A => S3932,
        B => S3934,
        Y => S3936
    );
NAND_2632: ENTITY WORK.NAND
    PORT MAP (
        A => S3933,
        B => S3935,
        Y => S3937
    );
NOR_1092: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_14,
        B => S1516,
        Y => S3938
    );
NOT_323: ENTITY WORK.NOT
    PORT MAP (
        A => S3938,
        Y => S3939
    );
NOR_1093: ENTITY WORK.NOR
    PORT MAP (
        A => S3937,
        B => S3938,
        Y => S3940
    );
NAND_2633: ENTITY WORK.NAND
    PORT MAP (
        A => S3936,
        B => S3939,
        Y => S3941
    );
NOR_1094: ENTITY WORK.NOR
    PORT MAP (
        A => S3932,
        B => S3940,
        Y => S3942
    );
NAND_2634: ENTITY WORK.NAND
    PORT MAP (
        A => S3933,
        B => S3941,
        Y => S3943
    );
NOR_1095: ENTITY WORK.NOR
    PORT MAP (
        A => S3925,
        B => S3942,
        Y => S3944
    );
NAND_2635: ENTITY WORK.NAND
    PORT MAP (
        A => S3924,
        B => S3943,
        Y => S3945
    );
NAND_2636: ENTITY WORK.NAND
    PORT MAP (
        A => S3937,
        B => S3938,
        Y => S3946
    );
NAND_2637: ENTITY WORK.NAND
    PORT MAP (
        A => S3941,
        B => S3946,
        Y => S3947
    );
NAND_2638: ENTITY WORK.NAND
    PORT MAP (
        A => S3930,
        B => S3945,
        Y => S3948
    );
NOT_324: ENTITY WORK.NOT
    PORT MAP (
        A => S3948,
        Y => S3949
    );
NOR_1096: ENTITY WORK.NOR
    PORT MAP (
        A => S3945,
        B => S3947,
        Y => S3950
    );
NOT_325: ENTITY WORK.NOT
    PORT MAP (
        A => S3950,
        Y => S3951
    );
NAND_2639: ENTITY WORK.NAND
    PORT MAP (
        A => S3948,
        B => S3951,
        Y => S3952
    );
NOR_1097: ENTITY WORK.NOR
    PORT MAP (
        A => S3949,
        B => S3950,
        Y => S3953
    );
NOR_1098: ENTITY WORK.NOR
    PORT MAP (
        A => S1516,
        B => S3945,
        Y => S3954
    );
NAND_2640: ENTITY WORK.NAND
    PORT MAP (
        A => S1515,
        B => S3944,
        Y => S3955
    );
NOR_1099: ENTITY WORK.NOR
    PORT MAP (
        A => S492,
        B => S3954,
        Y => S3956
    );
NAND_2641: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_14,
        B => S3955,
        Y => S3957
    );
NOR_1100: ENTITY WORK.NOR
    PORT MAP (
        A => S1745,
        B => S3957,
        Y => S3958
    );
NAND_2642: ENTITY WORK.NAND
    PORT MAP (
        A => S1746,
        B => S3956,
        Y => S3959
    );
NOR_1101: ENTITY WORK.NOR
    PORT MAP (
        A => S1746,
        B => S3956,
        Y => S3960
    );
NAND_2643: ENTITY WORK.NAND
    PORT MAP (
        A => S1745,
        B => S3957,
        Y => S3961
    );
NOR_1102: ENTITY WORK.NOR
    PORT MAP (
        A => S3958,
        B => S3960,
        Y => S3962
    );
NAND_2644: ENTITY WORK.NAND
    PORT MAP (
        A => S3959,
        B => S3961,
        Y => S3963
    );
NOR_1103: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_13,
        B => S1516,
        Y => S3964
    );
NAND_2645: ENTITY WORK.NAND
    PORT MAP (
        A => S548,
        B => S1515,
        Y => S3965
    );
NOR_1104: ENTITY WORK.NOR
    PORT MAP (
        A => S3963,
        B => S3964,
        Y => S3966
    );
NAND_2646: ENTITY WORK.NAND
    PORT MAP (
        A => S3962,
        B => S3965,
        Y => S3967
    );
NOR_1105: ENTITY WORK.NOR
    PORT MAP (
        A => S3958,
        B => S3966,
        Y => S3968
    );
NAND_2647: ENTITY WORK.NAND
    PORT MAP (
        A => S3959,
        B => S3967,
        Y => S3969
    );
NOR_1106: ENTITY WORK.NOR
    PORT MAP (
        A => S1849,
        B => S3923,
        Y => S3970
    );
NAND_2648: ENTITY WORK.NAND
    PORT MAP (
        A => S3969,
        B => S3970,
        Y => S3971
    );
NOR_1107: ENTITY WORK.NOR
    PORT MAP (
        A => S3925,
        B => S3969,
        Y => S3972
    );
NAND_2649: ENTITY WORK.NAND
    PORT MAP (
        A => S3952,
        B => S3971,
        Y => S3973
    );
NOR_1108: ENTITY WORK.NOR
    PORT MAP (
        A => S3972,
        B => S3973,
        Y => S3974
    );
NOT_326: ENTITY WORK.NOT
    PORT MAP (
        A => S3974,
        Y => S3975
    );
NOR_1109: ENTITY WORK.NOR
    PORT MAP (
        A => S1848,
        B => S3953,
        Y => S3976
    );
NAND_2650: ENTITY WORK.NAND
    PORT MAP (
        A => S1849,
        B => S3952,
        Y => S3977
    );
NOR_1110: ENTITY WORK.NOR
    PORT MAP (
        A => S3969,
        B => S3976,
        Y => S3978
    );
NAND_2651: ENTITY WORK.NAND
    PORT MAP (
        A => S3968,
        B => S3977,
        Y => S3979
    );
NOR_1111: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_15,
        B => S1849,
        Y => S3980
    );
NAND_2652: ENTITY WORK.NAND
    PORT MAP (
        A => S1304,
        B => S1848,
        Y => S3981
    );
NOR_1112: ENTITY WORK.NOR
    PORT MAP (
        A => S3923,
        B => S3980,
        Y => S3982
    );
NAND_2653: ENTITY WORK.NAND
    PORT MAP (
        A => S3922,
        B => S3981,
        Y => S3983
    );
NOR_1113: ENTITY WORK.NOR
    PORT MAP (
        A => S3978,
        B => S3983,
        Y => S3984
    );
NAND_2654: ENTITY WORK.NAND
    PORT MAP (
        A => S3979,
        B => S3982,
        Y => S3985
    );
NOR_1114: ENTITY WORK.NOR
    PORT MAP (
        A => S3962,
        B => S3965,
        Y => S3986
    );
NOR_1115: ENTITY WORK.NOR
    PORT MAP (
        A => S3966,
        B => S3986,
        Y => S3987
    );
NOR_1116: ENTITY WORK.NOR
    PORT MAP (
        A => S3985,
        B => S3987,
        Y => S3988
    );
NOT_327: ENTITY WORK.NOT
    PORT MAP (
        A => S3988,
        Y => S3989
    );
NOR_1117: ENTITY WORK.NOR
    PORT MAP (
        A => S3956,
        B => S3984,
        Y => S3990
    );
NAND_2655: ENTITY WORK.NAND
    PORT MAP (
        A => S3957,
        B => S3985,
        Y => S3991
    );
NOR_1118: ENTITY WORK.NOR
    PORT MAP (
        A => S3988,
        B => S3990,
        Y => S3992
    );
NAND_2656: ENTITY WORK.NAND
    PORT MAP (
        A => S3989,
        B => S3991,
        Y => S3993
    );
NOR_1119: ENTITY WORK.NOR
    PORT MAP (
        A => S1848,
        B => S3993,
        Y => S3994
    );
NAND_2657: ENTITY WORK.NAND
    PORT MAP (
        A => S1849,
        B => S3992,
        Y => S3995
    );
NOR_1120: ENTITY WORK.NOR
    PORT MAP (
        A => S1849,
        B => S3992,
        Y => S3996
    );
NAND_2658: ENTITY WORK.NAND
    PORT MAP (
        A => S1848,
        B => S3993,
        Y => S3997
    );
NOR_1121: ENTITY WORK.NOR
    PORT MAP (
        A => S3994,
        B => S3996,
        Y => S3998
    );
NAND_2659: ENTITY WORK.NAND
    PORT MAP (
        A => S3995,
        B => S3997,
        Y => S3999
    );
NOR_1122: ENTITY WORK.NOR
    PORT MAP (
        A => S1516,
        B => S3985,
        Y => S4000
    );
NAND_2660: ENTITY WORK.NAND
    PORT MAP (
        A => S1515,
        B => S3984,
        Y => S4001
    );
NOR_1123: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_13,
        B => S4000,
        Y => S4002
    );
NAND_2661: ENTITY WORK.NAND
    PORT MAP (
        A => S548,
        B => S4001,
        Y => S4003
    );
NOR_1124: ENTITY WORK.NOR
    PORT MAP (
        A => S548,
        B => S4001,
        Y => S4004
    );
NAND_2662: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_13,
        B => S4000,
        Y => S4005
    );
NOR_1125: ENTITY WORK.NOR
    PORT MAP (
        A => S4002,
        B => S4004,
        Y => S4006
    );
NAND_2663: ENTITY WORK.NAND
    PORT MAP (
        A => S4003,
        B => S4005,
        Y => S4007
    );
NOR_1126: ENTITY WORK.NOR
    PORT MAP (
        A => S1745,
        B => S4007,
        Y => S4008
    );
NAND_2664: ENTITY WORK.NAND
    PORT MAP (
        A => S1746,
        B => S4006,
        Y => S4009
    );
NOR_1127: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_12,
        B => S1516,
        Y => S4010
    );
NAND_2665: ENTITY WORK.NAND
    PORT MAP (
        A => S599,
        B => S1515,
        Y => S4011
    );
NOR_1128: ENTITY WORK.NOR
    PORT MAP (
        A => S1746,
        B => S4006,
        Y => S4012
    );
NAND_2666: ENTITY WORK.NAND
    PORT MAP (
        A => S1745,
        B => S4007,
        Y => S4013
    );
NOR_1129: ENTITY WORK.NOR
    PORT MAP (
        A => S4008,
        B => S4012,
        Y => S4014
    );
NAND_2667: ENTITY WORK.NAND
    PORT MAP (
        A => S4009,
        B => S4013,
        Y => S4015
    );
NOR_1130: ENTITY WORK.NOR
    PORT MAP (
        A => S4010,
        B => S4015,
        Y => S4016
    );
NAND_2668: ENTITY WORK.NAND
    PORT MAP (
        A => S4011,
        B => S4014,
        Y => S4017
    );
NOR_1131: ENTITY WORK.NOR
    PORT MAP (
        A => S4008,
        B => S4016,
        Y => S4018
    );
NAND_2669: ENTITY WORK.NAND
    PORT MAP (
        A => S4009,
        B => S4017,
        Y => S4019
    );
NOR_1132: ENTITY WORK.NOR
    PORT MAP (
        A => S3999,
        B => S4018,
        Y => S4020
    );
NAND_2670: ENTITY WORK.NAND
    PORT MAP (
        A => S3998,
        B => S4019,
        Y => S4021
    );
NOR_1133: ENTITY WORK.NOR
    PORT MAP (
        A => S3994,
        B => S4020,
        Y => S4022
    );
NAND_2671: ENTITY WORK.NAND
    PORT MAP (
        A => S3995,
        B => S4021,
        Y => S4023
    );
NOR_1134: ENTITY WORK.NOR
    PORT MAP (
        A => S1952,
        B => S4022,
        Y => S4024
    );
NAND_2672: ENTITY WORK.NAND
    PORT MAP (
        A => S1953,
        B => S4023,
        Y => S4025
    );
NOR_1135: ENTITY WORK.NOR
    PORT MAP (
        A => S1953,
        B => S4023,
        Y => S4026
    );
NAND_2673: ENTITY WORK.NAND
    PORT MAP (
        A => S1952,
        B => S4022,
        Y => S4027
    );
NOR_1136: ENTITY WORK.NOR
    PORT MAP (
        A => S3921,
        B => S4026,
        Y => S4028
    );
NAND_2674: ENTITY WORK.NAND
    PORT MAP (
        A => S3920,
        B => S4027,
        Y => S4029
    );
NAND_2675: ENTITY WORK.NAND
    PORT MAP (
        A => S4025,
        B => S4028,
        Y => S4030
    );
NAND_2676: ENTITY WORK.NAND
    PORT MAP (
        A => S3974,
        B => S4030,
        Y => S4031
    );
NOR_1137: ENTITY WORK.NOR
    PORT MAP (
        A => S3974,
        B => S4024,
        Y => S4032
    );
NAND_2677: ENTITY WORK.NAND
    PORT MAP (
        A => S3975,
        B => S4025,
        Y => S4033
    );
NOR_1138: ENTITY WORK.NOR
    PORT MAP (
        A => S4029,
        B => S4032,
        Y => S4034
    );
NAND_2678: ENTITY WORK.NAND
    PORT MAP (
        A => S4028,
        B => S4033,
        Y => S4035
    );
NOR_1139: ENTITY WORK.NOR
    PORT MAP (
        A => S3998,
        B => S4019,
        Y => S4036
    );
NOR_1140: ENTITY WORK.NOR
    PORT MAP (
        A => S4020,
        B => S4036,
        Y => S4037
    );
NOR_1141: ENTITY WORK.NOR
    PORT MAP (
        A => S4035,
        B => S4037,
        Y => S4038
    );
NOT_328: ENTITY WORK.NOT
    PORT MAP (
        A => S4038,
        Y => S4039
    );
NOR_1142: ENTITY WORK.NOR
    PORT MAP (
        A => S3992,
        B => S4034,
        Y => S4040
    );
NAND_2679: ENTITY WORK.NAND
    PORT MAP (
        A => S3993,
        B => S4035,
        Y => S4041
    );
NOR_1143: ENTITY WORK.NOR
    PORT MAP (
        A => S4038,
        B => S4040,
        Y => S4042
    );
NAND_2680: ENTITY WORK.NAND
    PORT MAP (
        A => S4039,
        B => S4041,
        Y => S4043
    );
NOR_1144: ENTITY WORK.NOR
    PORT MAP (
        A => S1952,
        B => S4043,
        Y => S4044
    );
NAND_2681: ENTITY WORK.NAND
    PORT MAP (
        A => S1953,
        B => S4042,
        Y => S4045
    );
NOR_1145: ENTITY WORK.NOR
    PORT MAP (
        A => S1953,
        B => S4042,
        Y => S4046
    );
NAND_2682: ENTITY WORK.NAND
    PORT MAP (
        A => S1952,
        B => S4043,
        Y => S4047
    );
NOR_1146: ENTITY WORK.NOR
    PORT MAP (
        A => S4044,
        B => S4046,
        Y => S4048
    );
NAND_2683: ENTITY WORK.NAND
    PORT MAP (
        A => S4045,
        B => S4047,
        Y => S4049
    );
NOR_1147: ENTITY WORK.NOR
    PORT MAP (
        A => S4011,
        B => S4014,
        Y => S4050
    );
NOR_1148: ENTITY WORK.NOR
    PORT MAP (
        A => S4016,
        B => S4050,
        Y => S4051
    );
NOR_1149: ENTITY WORK.NOR
    PORT MAP (
        A => S4035,
        B => S4051,
        Y => S4052
    );
NOT_329: ENTITY WORK.NOT
    PORT MAP (
        A => S4052,
        Y => S4053
    );
NAND_2684: ENTITY WORK.NAND
    PORT MAP (
        A => S4007,
        B => S4035,
        Y => S4054
    );
NOT_330: ENTITY WORK.NOT
    PORT MAP (
        A => S4054,
        Y => S4055
    );
NOR_1150: ENTITY WORK.NOR
    PORT MAP (
        A => S4052,
        B => S4055,
        Y => S4056
    );
NAND_2685: ENTITY WORK.NAND
    PORT MAP (
        A => S4053,
        B => S4054,
        Y => S4057
    );
NOR_1151: ENTITY WORK.NOR
    PORT MAP (
        A => S1848,
        B => S4057,
        Y => S4058
    );
NAND_2686: ENTITY WORK.NAND
    PORT MAP (
        A => S1849,
        B => S4056,
        Y => S4059
    );
NOR_1152: ENTITY WORK.NOR
    PORT MAP (
        A => S1849,
        B => S4056,
        Y => S4060
    );
NAND_2687: ENTITY WORK.NAND
    PORT MAP (
        A => S1848,
        B => S4057,
        Y => S4061
    );
NOR_1153: ENTITY WORK.NOR
    PORT MAP (
        A => S4058,
        B => S4060,
        Y => S4062
    );
NAND_2688: ENTITY WORK.NAND
    PORT MAP (
        A => S4059,
        B => S4061,
        Y => S4063
    );
NOR_1154: ENTITY WORK.NOR
    PORT MAP (
        A => S1516,
        B => S4035,
        Y => S4064
    );
NAND_2689: ENTITY WORK.NAND
    PORT MAP (
        A => S1515,
        B => S4034,
        Y => S4065
    );
NOR_1155: ENTITY WORK.NOR
    PORT MAP (
        A => S599,
        B => S4064,
        Y => S4066
    );
NAND_2690: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_12,
        B => S4065,
        Y => S4067
    );
NOR_1156: ENTITY WORK.NOR
    PORT MAP (
        A => S4011,
        B => S4035,
        Y => S4068
    );
NOT_331: ENTITY WORK.NOT
    PORT MAP (
        A => S4068,
        Y => S4069
    );
NOR_1157: ENTITY WORK.NOR
    PORT MAP (
        A => S4066,
        B => S4068,
        Y => S4070
    );
NAND_2691: ENTITY WORK.NAND
    PORT MAP (
        A => S4067,
        B => S4069,
        Y => S4071
    );
NOR_1158: ENTITY WORK.NOR
    PORT MAP (
        A => S1745,
        B => S4070,
        Y => S4072
    );
NAND_2692: ENTITY WORK.NAND
    PORT MAP (
        A => S1746,
        B => S4071,
        Y => S4073
    );
NOR_1159: ENTITY WORK.NOR
    PORT MAP (
        A => S1746,
        B => S4071,
        Y => S4074
    );
NAND_2693: ENTITY WORK.NAND
    PORT MAP (
        A => S1745,
        B => S4070,
        Y => S4075
    );
NOR_1160: ENTITY WORK.NOR
    PORT MAP (
        A => S4072,
        B => S4074,
        Y => S4076
    );
NAND_2694: ENTITY WORK.NAND
    PORT MAP (
        A => S4073,
        B => S4075,
        Y => S4077
    );
NOR_1161: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_11,
        B => S1516,
        Y => S4078
    );
NAND_2695: ENTITY WORK.NAND
    PORT MAP (
        A => S651,
        B => S1515,
        Y => S4079
    );
NOR_1162: ENTITY WORK.NOR
    PORT MAP (
        A => S4077,
        B => S4078,
        Y => S4080
    );
NAND_2696: ENTITY WORK.NAND
    PORT MAP (
        A => S4076,
        B => S4079,
        Y => S4081
    );
NOR_1163: ENTITY WORK.NOR
    PORT MAP (
        A => S4072,
        B => S4080,
        Y => S4082
    );
NAND_2697: ENTITY WORK.NAND
    PORT MAP (
        A => S4073,
        B => S4081,
        Y => S4083
    );
NOR_1164: ENTITY WORK.NOR
    PORT MAP (
        A => S4063,
        B => S4082,
        Y => S4084
    );
NAND_2698: ENTITY WORK.NAND
    PORT MAP (
        A => S4062,
        B => S4083,
        Y => S4085
    );
NOR_1165: ENTITY WORK.NOR
    PORT MAP (
        A => S4058,
        B => S4084,
        Y => S4086
    );
NAND_2699: ENTITY WORK.NAND
    PORT MAP (
        A => S4059,
        B => S4085,
        Y => S4087
    );
NOR_1166: ENTITY WORK.NOR
    PORT MAP (
        A => S4049,
        B => S4086,
        Y => S4088
    );
NAND_2700: ENTITY WORK.NAND
    PORT MAP (
        A => S4048,
        B => S4087,
        Y => S4089
    );
NOR_1167: ENTITY WORK.NOR
    PORT MAP (
        A => S4044,
        B => S4088,
        Y => S4090
    );
NAND_2701: ENTITY WORK.NAND
    PORT MAP (
        A => S4045,
        B => S4089,
        Y => S4091
    );
NAND_2702: ENTITY WORK.NAND
    PORT MAP (
        A => S1597,
        B => S3918,
        Y => S4092
    );
NAND_2703: ENTITY WORK.NAND
    PORT MAP (
        A => S3920,
        B => S4090,
        Y => S4093
    );
NOR_1168: ENTITY WORK.NOR
    PORT MAP (
        A => S4090,
        B => S4092,
        Y => S4094
    );
NOT_332: ENTITY WORK.NOT
    PORT MAP (
        A => S4094,
        Y => S4095
    );
NOR_1169: ENTITY WORK.NOR
    PORT MAP (
        A => S4031,
        B => S4094,
        Y => S4096
    );
NAND_2704: ENTITY WORK.NAND
    PORT MAP (
        A => S4093,
        B => S4095,
        Y => S4097
    );
NOR_1170: ENTITY WORK.NOR
    PORT MAP (
        A => S4031,
        B => S4097,
        Y => S4098
    );
NAND_2705: ENTITY WORK.NAND
    PORT MAP (
        A => S4093,
        B => S4096,
        Y => S4099
    );
NOR_1171: ENTITY WORK.NOR
    PORT MAP (
        A => S1597,
        B => S4031,
        Y => S4100
    );
NOT_333: ENTITY WORK.NOT
    PORT MAP (
        A => S4100,
        Y => S4101
    );
NOR_1172: ENTITY WORK.NOR
    PORT MAP (
        A => S4091,
        B => S4100,
        Y => S4102
    );
NAND_2706: ENTITY WORK.NAND
    PORT MAP (
        A => S4090,
        B => S4101,
        Y => S4103
    );
NAND_2707: ENTITY WORK.NAND
    PORT MAP (
        A => S1597,
        B => S3975,
        Y => S4104
    );
NAND_2708: ENTITY WORK.NAND
    PORT MAP (
        A => S3918,
        B => S4104,
        Y => S4105
    );
NOT_334: ENTITY WORK.NOT
    PORT MAP (
        A => S4105,
        Y => S4106
    );
NOR_1173: ENTITY WORK.NOR
    PORT MAP (
        A => S4102,
        B => S4105,
        Y => S4107
    );
NAND_2709: ENTITY WORK.NAND
    PORT MAP (
        A => S4103,
        B => S4106,
        Y => S4108
    );
NOR_1174: ENTITY WORK.NOR
    PORT MAP (
        A => S4048,
        B => S4087,
        Y => S4109
    );
NOR_1175: ENTITY WORK.NOR
    PORT MAP (
        A => S4088,
        B => S4109,
        Y => S4110
    );
NOR_1176: ENTITY WORK.NOR
    PORT MAP (
        A => S4108,
        B => S4110,
        Y => S4111
    );
NOT_335: ENTITY WORK.NOT
    PORT MAP (
        A => S4111,
        Y => S4112
    );
NOR_1177: ENTITY WORK.NOR
    PORT MAP (
        A => S4042,
        B => S4107,
        Y => S4113
    );
NAND_2710: ENTITY WORK.NAND
    PORT MAP (
        A => S4043,
        B => S4108,
        Y => S4114
    );
NOR_1178: ENTITY WORK.NOR
    PORT MAP (
        A => S4111,
        B => S4113,
        Y => S4115
    );
NAND_2711: ENTITY WORK.NAND
    PORT MAP (
        A => S4112,
        B => S4114,
        Y => S4116
    );
NOR_1179: ENTITY WORK.NOR
    PORT MAP (
        A => S1597,
        B => S4116,
        Y => S4117
    );
NAND_2712: ENTITY WORK.NAND
    PORT MAP (
        A => S1598,
        B => S4115,
        Y => S4118
    );
NOR_1180: ENTITY WORK.NOR
    PORT MAP (
        A => S1598,
        B => S4115,
        Y => S4119
    );
NAND_2713: ENTITY WORK.NAND
    PORT MAP (
        A => S1597,
        B => S4116,
        Y => S4120
    );
NOR_1181: ENTITY WORK.NOR
    PORT MAP (
        A => S4117,
        B => S4119,
        Y => S4121
    );
NAND_2714: ENTITY WORK.NAND
    PORT MAP (
        A => S4118,
        B => S4120,
        Y => S4122
    );
NOR_1182: ENTITY WORK.NOR
    PORT MAP (
        A => S4062,
        B => S4083,
        Y => S4123
    );
NOR_1183: ENTITY WORK.NOR
    PORT MAP (
        A => S4084,
        B => S4123,
        Y => S4124
    );
NOR_1184: ENTITY WORK.NOR
    PORT MAP (
        A => S4108,
        B => S4124,
        Y => S4125
    );
NOT_336: ENTITY WORK.NOT
    PORT MAP (
        A => S4125,
        Y => S4126
    );
NOR_1185: ENTITY WORK.NOR
    PORT MAP (
        A => S4056,
        B => S4107,
        Y => S4127
    );
NAND_2715: ENTITY WORK.NAND
    PORT MAP (
        A => S4057,
        B => S4108,
        Y => S4128
    );
NOR_1186: ENTITY WORK.NOR
    PORT MAP (
        A => S4125,
        B => S4127,
        Y => S4129
    );
NAND_2716: ENTITY WORK.NAND
    PORT MAP (
        A => S4126,
        B => S4128,
        Y => S4130
    );
NOR_1187: ENTITY WORK.NOR
    PORT MAP (
        A => S1952,
        B => S4130,
        Y => S4131
    );
NAND_2717: ENTITY WORK.NAND
    PORT MAP (
        A => S1953,
        B => S4129,
        Y => S4132
    );
NOR_1188: ENTITY WORK.NOR
    PORT MAP (
        A => S1953,
        B => S4129,
        Y => S4133
    );
NAND_2718: ENTITY WORK.NAND
    PORT MAP (
        A => S1952,
        B => S4130,
        Y => S4134
    );
NOR_1189: ENTITY WORK.NOR
    PORT MAP (
        A => S4131,
        B => S4133,
        Y => S4135
    );
NAND_2719: ENTITY WORK.NAND
    PORT MAP (
        A => S4132,
        B => S4134,
        Y => S4136
    );
NOR_1190: ENTITY WORK.NOR
    PORT MAP (
        A => S4076,
        B => S4079,
        Y => S4137
    );
NOR_1191: ENTITY WORK.NOR
    PORT MAP (
        A => S4080,
        B => S4137,
        Y => S4138
    );
NOR_1192: ENTITY WORK.NOR
    PORT MAP (
        A => S4108,
        B => S4138,
        Y => S4139
    );
NOT_337: ENTITY WORK.NOT
    PORT MAP (
        A => S4139,
        Y => S4140
    );
NAND_2720: ENTITY WORK.NAND
    PORT MAP (
        A => S4070,
        B => S4108,
        Y => S4141
    );
NOT_338: ENTITY WORK.NOT
    PORT MAP (
        A => S4141,
        Y => S4142
    );
NOR_1193: ENTITY WORK.NOR
    PORT MAP (
        A => S4139,
        B => S4142,
        Y => S4143
    );
NAND_2721: ENTITY WORK.NAND
    PORT MAP (
        A => S4140,
        B => S4141,
        Y => S4144
    );
NOR_1194: ENTITY WORK.NOR
    PORT MAP (
        A => S1848,
        B => S4144,
        Y => S4145
    );
NAND_2722: ENTITY WORK.NAND
    PORT MAP (
        A => S1849,
        B => S4143,
        Y => S4146
    );
NOR_1195: ENTITY WORK.NOR
    PORT MAP (
        A => S1849,
        B => S4143,
        Y => S4147
    );
NAND_2723: ENTITY WORK.NAND
    PORT MAP (
        A => S1848,
        B => S4144,
        Y => S4148
    );
NOR_1196: ENTITY WORK.NOR
    PORT MAP (
        A => S4145,
        B => S4147,
        Y => S4149
    );
NAND_2724: ENTITY WORK.NAND
    PORT MAP (
        A => S4146,
        B => S4148,
        Y => S4150
    );
NOR_1197: ENTITY WORK.NOR
    PORT MAP (
        A => S1516,
        B => S4108,
        Y => S4151
    );
NAND_2725: ENTITY WORK.NAND
    PORT MAP (
        A => S1515,
        B => S4107,
        Y => S4152
    );
NOR_1198: ENTITY WORK.NOR
    PORT MAP (
        A => S651,
        B => S4152,
        Y => S4153
    );
NAND_2726: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_11,
        B => S4151,
        Y => S4154
    );
NOR_1199: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_11,
        B => S4151,
        Y => S4155
    );
NAND_2727: ENTITY WORK.NAND
    PORT MAP (
        A => S651,
        B => S4152,
        Y => S4156
    );
NAND_2728: ENTITY WORK.NAND
    PORT MAP (
        A => S4154,
        B => S4156,
        Y => S4157
    );
NOR_1200: ENTITY WORK.NOR
    PORT MAP (
        A => S4153,
        B => S4155,
        Y => S4158
    );
NOR_1201: ENTITY WORK.NOR
    PORT MAP (
        A => S1745,
        B => S4157,
        Y => S4159
    );
NAND_2729: ENTITY WORK.NAND
    PORT MAP (
        A => S1746,
        B => S4158,
        Y => S4160
    );
NOR_1202: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_10,
        B => S1516,
        Y => S4161
    );
NAND_2730: ENTITY WORK.NAND
    PORT MAP (
        A => S702,
        B => S1515,
        Y => S4162
    );
NOR_1203: ENTITY WORK.NOR
    PORT MAP (
        A => S1746,
        B => S4158,
        Y => S4163
    );
NAND_2731: ENTITY WORK.NAND
    PORT MAP (
        A => S1745,
        B => S4157,
        Y => S4164
    );
NOR_1204: ENTITY WORK.NOR
    PORT MAP (
        A => S4159,
        B => S4163,
        Y => S4165
    );
NAND_2732: ENTITY WORK.NAND
    PORT MAP (
        A => S4160,
        B => S4164,
        Y => S4166
    );
NOR_1205: ENTITY WORK.NOR
    PORT MAP (
        A => S4161,
        B => S4166,
        Y => S4167
    );
NAND_2733: ENTITY WORK.NAND
    PORT MAP (
        A => S4162,
        B => S4165,
        Y => S4168
    );
NOR_1206: ENTITY WORK.NOR
    PORT MAP (
        A => S4159,
        B => S4167,
        Y => S4169
    );
NAND_2734: ENTITY WORK.NAND
    PORT MAP (
        A => S4160,
        B => S4168,
        Y => S4170
    );
NOR_1207: ENTITY WORK.NOR
    PORT MAP (
        A => S4150,
        B => S4169,
        Y => S4171
    );
NAND_2735: ENTITY WORK.NAND
    PORT MAP (
        A => S4149,
        B => S4170,
        Y => S4172
    );
NOR_1208: ENTITY WORK.NOR
    PORT MAP (
        A => S4145,
        B => S4171,
        Y => S4173
    );
NAND_2736: ENTITY WORK.NAND
    PORT MAP (
        A => S4146,
        B => S4172,
        Y => S4174
    );
NOR_1209: ENTITY WORK.NOR
    PORT MAP (
        A => S4136,
        B => S4173,
        Y => S4175
    );
NAND_2737: ENTITY WORK.NAND
    PORT MAP (
        A => S4135,
        B => S4174,
        Y => S4176
    );
NOR_1210: ENTITY WORK.NOR
    PORT MAP (
        A => S4131,
        B => S4175,
        Y => S4177
    );
NAND_2738: ENTITY WORK.NAND
    PORT MAP (
        A => S4132,
        B => S4176,
        Y => S4178
    );
NOR_1211: ENTITY WORK.NOR
    PORT MAP (
        A => S4122,
        B => S4177,
        Y => S4179
    );
NAND_2739: ENTITY WORK.NAND
    PORT MAP (
        A => S4121,
        B => S4178,
        Y => S4180
    );
NOR_1212: ENTITY WORK.NOR
    PORT MAP (
        A => S4117,
        B => S4179,
        Y => S4181
    );
NAND_2740: ENTITY WORK.NAND
    PORT MAP (
        A => S4118,
        B => S4180,
        Y => S4182
    );
NOR_1213: ENTITY WORK.NOR
    PORT MAP (
        A => S2106,
        B => S4181,
        Y => S4183
    );
NAND_2741: ENTITY WORK.NAND
    PORT MAP (
        A => S2107,
        B => S4182,
        Y => S4184
    );
NOR_1214: ENTITY WORK.NOR
    PORT MAP (
        A => S2107,
        B => S4182,
        Y => S4185
    );
NAND_2742: ENTITY WORK.NAND
    PORT MAP (
        A => S2106,
        B => S4181,
        Y => S4186
    );
NOR_1215: ENTITY WORK.NOR
    PORT MAP (
        A => S3917,
        B => S4185,
        Y => S4187
    );
NAND_2743: ENTITY WORK.NAND
    PORT MAP (
        A => S3916,
        B => S4186,
        Y => S4188
    );
NOR_1216: ENTITY WORK.NOR
    PORT MAP (
        A => S4183,
        B => S4188,
        Y => S4189
    );
NOR_1217: ENTITY WORK.NOR
    PORT MAP (
        A => S4099,
        B => S4189,
        Y => S4190
    );
NOT_339: ENTITY WORK.NOT
    PORT MAP (
        A => S4190,
        Y => S4191
    );
NOR_1218: ENTITY WORK.NOR
    PORT MAP (
        A => S4098,
        B => S4183,
        Y => S4192
    );
NAND_2744: ENTITY WORK.NAND
    PORT MAP (
        A => S4099,
        B => S4184,
        Y => S4193
    );
NOR_1219: ENTITY WORK.NOR
    PORT MAP (
        A => S4188,
        B => S4192,
        Y => S4194
    );
NAND_2745: ENTITY WORK.NAND
    PORT MAP (
        A => S4187,
        B => S4193,
        Y => S4195
    );
NOR_1220: ENTITY WORK.NOR
    PORT MAP (
        A => S4121,
        B => S4178,
        Y => S4196
    );
NAND_2746: ENTITY WORK.NAND
    PORT MAP (
        A => S4122,
        B => S4177,
        Y => S4197
    );
NOR_1221: ENTITY WORK.NOR
    PORT MAP (
        A => S4179,
        B => S4196,
        Y => S4198
    );
NAND_2747: ENTITY WORK.NAND
    PORT MAP (
        A => S4180,
        B => S4197,
        Y => S4199
    );
NOR_1222: ENTITY WORK.NOR
    PORT MAP (
        A => S4195,
        B => S4198,
        Y => S4200
    );
NAND_2748: ENTITY WORK.NAND
    PORT MAP (
        A => S4194,
        B => S4199,
        Y => S4201
    );
NOR_1223: ENTITY WORK.NOR
    PORT MAP (
        A => S4115,
        B => S4194,
        Y => S4202
    );
NAND_2749: ENTITY WORK.NAND
    PORT MAP (
        A => S4116,
        B => S4195,
        Y => S4203
    );
NOR_1224: ENTITY WORK.NOR
    PORT MAP (
        A => S4200,
        B => S4202,
        Y => S4204
    );
NAND_2750: ENTITY WORK.NAND
    PORT MAP (
        A => S4201,
        B => S4203,
        Y => S4205
    );
NOR_1225: ENTITY WORK.NOR
    PORT MAP (
        A => S2106,
        B => S4205,
        Y => S4206
    );
NAND_2751: ENTITY WORK.NAND
    PORT MAP (
        A => S2107,
        B => S4204,
        Y => S4207
    );
NOR_1226: ENTITY WORK.NOR
    PORT MAP (
        A => S2107,
        B => S4204,
        Y => S4208
    );
NAND_2752: ENTITY WORK.NAND
    PORT MAP (
        A => S2106,
        B => S4205,
        Y => S4209
    );
NOR_1227: ENTITY WORK.NOR
    PORT MAP (
        A => S4206,
        B => S4208,
        Y => S4210
    );
NAND_2753: ENTITY WORK.NAND
    PORT MAP (
        A => S4207,
        B => S4209,
        Y => S4211
    );
NOR_1228: ENTITY WORK.NOR
    PORT MAP (
        A => S4135,
        B => S4174,
        Y => S4212
    );
NAND_2754: ENTITY WORK.NAND
    PORT MAP (
        A => S4136,
        B => S4173,
        Y => S4213
    );
NOR_1229: ENTITY WORK.NOR
    PORT MAP (
        A => S4175,
        B => S4212,
        Y => S4214
    );
NAND_2755: ENTITY WORK.NAND
    PORT MAP (
        A => S4176,
        B => S4213,
        Y => S4215
    );
NOR_1230: ENTITY WORK.NOR
    PORT MAP (
        A => S4195,
        B => S4214,
        Y => S4216
    );
NAND_2756: ENTITY WORK.NAND
    PORT MAP (
        A => S4194,
        B => S4215,
        Y => S4217
    );
NOR_1231: ENTITY WORK.NOR
    PORT MAP (
        A => S4129,
        B => S4194,
        Y => S4218
    );
NAND_2757: ENTITY WORK.NAND
    PORT MAP (
        A => S4130,
        B => S4195,
        Y => S4219
    );
NOR_1232: ENTITY WORK.NOR
    PORT MAP (
        A => S4216,
        B => S4218,
        Y => S4220
    );
NAND_2758: ENTITY WORK.NAND
    PORT MAP (
        A => S4217,
        B => S4219,
        Y => S4221
    );
NOR_1233: ENTITY WORK.NOR
    PORT MAP (
        A => S1597,
        B => S4221,
        Y => S4222
    );
NAND_2759: ENTITY WORK.NAND
    PORT MAP (
        A => S1598,
        B => S4220,
        Y => S4223
    );
NOR_1234: ENTITY WORK.NOR
    PORT MAP (
        A => S1598,
        B => S4220,
        Y => S4224
    );
NAND_2760: ENTITY WORK.NAND
    PORT MAP (
        A => S1597,
        B => S4221,
        Y => S4225
    );
NOR_1235: ENTITY WORK.NOR
    PORT MAP (
        A => S4222,
        B => S4224,
        Y => S4226
    );
NAND_2761: ENTITY WORK.NAND
    PORT MAP (
        A => S4223,
        B => S4225,
        Y => S4227
    );
NOR_1236: ENTITY WORK.NOR
    PORT MAP (
        A => S4149,
        B => S4170,
        Y => S4228
    );
NAND_2762: ENTITY WORK.NAND
    PORT MAP (
        A => S4150,
        B => S4169,
        Y => S4229
    );
NOR_1237: ENTITY WORK.NOR
    PORT MAP (
        A => S4171,
        B => S4228,
        Y => S4230
    );
NAND_2763: ENTITY WORK.NAND
    PORT MAP (
        A => S4172,
        B => S4229,
        Y => S4231
    );
NOR_1238: ENTITY WORK.NOR
    PORT MAP (
        A => S4195,
        B => S4230,
        Y => S4232
    );
NAND_2764: ENTITY WORK.NAND
    PORT MAP (
        A => S4194,
        B => S4231,
        Y => S4233
    );
NOR_1239: ENTITY WORK.NOR
    PORT MAP (
        A => S4143,
        B => S4194,
        Y => S4234
    );
NAND_2765: ENTITY WORK.NAND
    PORT MAP (
        A => S4144,
        B => S4195,
        Y => S4235
    );
NOR_1240: ENTITY WORK.NOR
    PORT MAP (
        A => S4232,
        B => S4234,
        Y => S4236
    );
NAND_2766: ENTITY WORK.NAND
    PORT MAP (
        A => S4233,
        B => S4235,
        Y => S4237
    );
NOR_1241: ENTITY WORK.NOR
    PORT MAP (
        A => S1952,
        B => S4237,
        Y => S4238
    );
NAND_2767: ENTITY WORK.NAND
    PORT MAP (
        A => S1953,
        B => S4236,
        Y => S4239
    );
NOR_1242: ENTITY WORK.NOR
    PORT MAP (
        A => S1953,
        B => S4236,
        Y => S4240
    );
NAND_2768: ENTITY WORK.NAND
    PORT MAP (
        A => S1952,
        B => S4237,
        Y => S4241
    );
NOR_1243: ENTITY WORK.NOR
    PORT MAP (
        A => S4238,
        B => S4240,
        Y => S4242
    );
NAND_2769: ENTITY WORK.NAND
    PORT MAP (
        A => S4239,
        B => S4241,
        Y => S4243
    );
NOR_1244: ENTITY WORK.NOR
    PORT MAP (
        A => S4158,
        B => S4194,
        Y => S4244
    );
NAND_2770: ENTITY WORK.NAND
    PORT MAP (
        A => S4157,
        B => S4195,
        Y => S4245
    );
NOR_1245: ENTITY WORK.NOR
    PORT MAP (
        A => S4162,
        B => S4165,
        Y => S4246
    );
NAND_2771: ENTITY WORK.NAND
    PORT MAP (
        A => S4161,
        B => S4166,
        Y => S4247
    );
NOR_1246: ENTITY WORK.NOR
    PORT MAP (
        A => S4167,
        B => S4246,
        Y => S4248
    );
NAND_2772: ENTITY WORK.NAND
    PORT MAP (
        A => S4168,
        B => S4247,
        Y => S4249
    );
NOR_1247: ENTITY WORK.NOR
    PORT MAP (
        A => S4195,
        B => S4248,
        Y => S4250
    );
NAND_2773: ENTITY WORK.NAND
    PORT MAP (
        A => S4194,
        B => S4249,
        Y => S4251
    );
NOR_1248: ENTITY WORK.NOR
    PORT MAP (
        A => S4244,
        B => S4250,
        Y => S4252
    );
NAND_2774: ENTITY WORK.NAND
    PORT MAP (
        A => S4245,
        B => S4251,
        Y => S4253
    );
NOR_1249: ENTITY WORK.NOR
    PORT MAP (
        A => S1848,
        B => S4253,
        Y => S4254
    );
NAND_2775: ENTITY WORK.NAND
    PORT MAP (
        A => S1849,
        B => S4252,
        Y => S4255
    );
NOR_1250: ENTITY WORK.NOR
    PORT MAP (
        A => S1849,
        B => S4252,
        Y => S4256
    );
NAND_2776: ENTITY WORK.NAND
    PORT MAP (
        A => S1848,
        B => S4253,
        Y => S4257
    );
NOR_1251: ENTITY WORK.NOR
    PORT MAP (
        A => S4254,
        B => S4256,
        Y => S4258
    );
NAND_2777: ENTITY WORK.NAND
    PORT MAP (
        A => S4255,
        B => S4257,
        Y => S4259
    );
NOR_1252: ENTITY WORK.NOR
    PORT MAP (
        A => S1516,
        B => S4195,
        Y => S4260
    );
NAND_2778: ENTITY WORK.NAND
    PORT MAP (
        A => S1515,
        B => S4194,
        Y => S4261
    );
NOR_1253: ENTITY WORK.NOR
    PORT MAP (
        A => S702,
        B => S4261,
        Y => S4262
    );
NAND_2779: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_10,
        B => S4260,
        Y => S4263
    );
NOR_1254: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_10,
        B => S4260,
        Y => S4264
    );
NAND_2780: ENTITY WORK.NAND
    PORT MAP (
        A => S702,
        B => S4261,
        Y => S4265
    );
NOR_1255: ENTITY WORK.NOR
    PORT MAP (
        A => S4262,
        B => S4264,
        Y => S4266
    );
NAND_2781: ENTITY WORK.NAND
    PORT MAP (
        A => S4263,
        B => S4265,
        Y => S4267
    );
NOR_1256: ENTITY WORK.NOR
    PORT MAP (
        A => S1745,
        B => S4267,
        Y => S4268
    );
NAND_2782: ENTITY WORK.NAND
    PORT MAP (
        A => S1746,
        B => S4266,
        Y => S4269
    );
NOR_1257: ENTITY WORK.NOR
    PORT MAP (
        A => S1746,
        B => S4266,
        Y => S4270
    );
NAND_2783: ENTITY WORK.NAND
    PORT MAP (
        A => S1745,
        B => S4267,
        Y => S4271
    );
NOR_1258: ENTITY WORK.NOR
    PORT MAP (
        A => S4268,
        B => S4270,
        Y => S4272
    );
NAND_2784: ENTITY WORK.NAND
    PORT MAP (
        A => S4269,
        B => S4271,
        Y => S4273
    );
NOR_1259: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_9,
        B => S1516,
        Y => S4274
    );
NAND_2785: ENTITY WORK.NAND
    PORT MAP (
        A => S754,
        B => S1515,
        Y => S4275
    );
NOR_1260: ENTITY WORK.NOR
    PORT MAP (
        A => S4273,
        B => S4274,
        Y => S4276
    );
NAND_2786: ENTITY WORK.NAND
    PORT MAP (
        A => S4272,
        B => S4275,
        Y => S4277
    );
NOR_1261: ENTITY WORK.NOR
    PORT MAP (
        A => S4268,
        B => S4276,
        Y => S4278
    );
NAND_2787: ENTITY WORK.NAND
    PORT MAP (
        A => S4269,
        B => S4277,
        Y => S4279
    );
NOR_1262: ENTITY WORK.NOR
    PORT MAP (
        A => S4259,
        B => S4278,
        Y => S4280
    );
NAND_2788: ENTITY WORK.NAND
    PORT MAP (
        A => S4258,
        B => S4279,
        Y => S4281
    );
NOR_1263: ENTITY WORK.NOR
    PORT MAP (
        A => S4254,
        B => S4280,
        Y => S4282
    );
NAND_2789: ENTITY WORK.NAND
    PORT MAP (
        A => S4255,
        B => S4281,
        Y => S4283
    );
NOR_1264: ENTITY WORK.NOR
    PORT MAP (
        A => S4243,
        B => S4282,
        Y => S4284
    );
NAND_2790: ENTITY WORK.NAND
    PORT MAP (
        A => S4242,
        B => S4283,
        Y => S4285
    );
NOR_1265: ENTITY WORK.NOR
    PORT MAP (
        A => S4238,
        B => S4284,
        Y => S4286
    );
NAND_2791: ENTITY WORK.NAND
    PORT MAP (
        A => S4239,
        B => S4285,
        Y => S4287
    );
NOR_1266: ENTITY WORK.NOR
    PORT MAP (
        A => S4227,
        B => S4286,
        Y => S4288
    );
NAND_2792: ENTITY WORK.NAND
    PORT MAP (
        A => S4226,
        B => S4287,
        Y => S4289
    );
NOR_1267: ENTITY WORK.NOR
    PORT MAP (
        A => S4222,
        B => S4288,
        Y => S4290
    );
NAND_2793: ENTITY WORK.NAND
    PORT MAP (
        A => S4223,
        B => S4289,
        Y => S4291
    );
NOR_1268: ENTITY WORK.NOR
    PORT MAP (
        A => S4211,
        B => S4290,
        Y => S4292
    );
NAND_2794: ENTITY WORK.NAND
    PORT MAP (
        A => S4210,
        B => S4291,
        Y => S4293
    );
NOR_1269: ENTITY WORK.NOR
    PORT MAP (
        A => S4206,
        B => S4292,
        Y => S4294
    );
NAND_2795: ENTITY WORK.NAND
    PORT MAP (
        A => S4207,
        B => S4293,
        Y => S4295
    );
NAND_2796: ENTITY WORK.NAND
    PORT MAP (
        A => S2206,
        B => S4295,
        Y => S4296
    );
NAND_2797: ENTITY WORK.NAND
    PORT MAP (
        A => S3914,
        B => S4295,
        Y => S4297
    );
NAND_2798: ENTITY WORK.NAND
    PORT MAP (
        A => S3917,
        B => S4297,
        Y => S4298
    );
NAND_2799: ENTITY WORK.NAND
    PORT MAP (
        A => S4296,
        B => S4298,
        Y => S4299
    );
NAND_2800: ENTITY WORK.NAND
    PORT MAP (
        A => S4190,
        B => S4299,
        Y => S4300
    );
NOT_340: ENTITY WORK.NOT
    PORT MAP (
        A => S4300,
        Y => S4301
    );
NOR_1270: ENTITY WORK.NOR
    PORT MAP (
        A => S2311,
        B => S4300,
        Y => S4302
    );
NAND_2801: ENTITY WORK.NAND
    PORT MAP (
        A => S2312,
        B => S4301,
        Y => S4303
    );
NOR_1271: ENTITY WORK.NOR
    PORT MAP (
        A => S2312,
        B => S4190,
        Y => S4304
    );
NOR_1272: ENTITY WORK.NOR
    PORT MAP (
        A => S4302,
        B => S4304,
        Y => S4305
    );
NOT_341: ENTITY WORK.NOT
    PORT MAP (
        A => S4305,
        Y => S4306
    );
NOR_1273: ENTITY WORK.NOR
    PORT MAP (
        A => S3917,
        B => S4191,
        Y => S4307
    );
NAND_2802: ENTITY WORK.NAND
    PORT MAP (
        A => S3916,
        B => S4190,
        Y => S4308
    );
NOR_1274: ENTITY WORK.NOR
    PORT MAP (
        A => S2206,
        B => S4098,
        Y => S4309
    );
NOR_1275: ENTITY WORK.NOR
    PORT MAP (
        A => S4294,
        B => S4309,
        Y => S4310
    );
NOR_1276: ENTITY WORK.NOR
    PORT MAP (
        A => S4297,
        B => S4309,
        Y => S4311
    );
NAND_2803: ENTITY WORK.NAND
    PORT MAP (
        A => S3914,
        B => S4310,
        Y => S4312
    );
NOR_1277: ENTITY WORK.NOR
    PORT MAP (
        A => S4307,
        B => S4311,
        Y => S4313
    );
NAND_2804: ENTITY WORK.NAND
    PORT MAP (
        A => S4308,
        B => S4312,
        Y => S4314
    );
NOR_1278: ENTITY WORK.NOR
    PORT MAP (
        A => S4210,
        B => S4291,
        Y => S4315
    );
NOR_1279: ENTITY WORK.NOR
    PORT MAP (
        A => S4292,
        B => S4315,
        Y => S4316
    );
NOR_1280: ENTITY WORK.NOR
    PORT MAP (
        A => S4313,
        B => S4316,
        Y => S4317
    );
NOT_342: ENTITY WORK.NOT
    PORT MAP (
        A => S4317,
        Y => S4318
    );
NOR_1281: ENTITY WORK.NOR
    PORT MAP (
        A => S4204,
        B => S4314,
        Y => S4319
    );
NAND_2805: ENTITY WORK.NAND
    PORT MAP (
        A => S4205,
        B => S4313,
        Y => S4320
    );
NOR_1282: ENTITY WORK.NOR
    PORT MAP (
        A => S4317,
        B => S4319,
        Y => S4321
    );
NAND_2806: ENTITY WORK.NAND
    PORT MAP (
        A => S4318,
        B => S4320,
        Y => S4322
    );
NOR_1283: ENTITY WORK.NOR
    PORT MAP (
        A => S2205,
        B => S4322,
        Y => S4323
    );
NAND_2807: ENTITY WORK.NAND
    PORT MAP (
        A => S2206,
        B => S4321,
        Y => S4324
    );
NOR_1284: ENTITY WORK.NOR
    PORT MAP (
        A => S2206,
        B => S4321,
        Y => S4325
    );
NAND_2808: ENTITY WORK.NAND
    PORT MAP (
        A => S2205,
        B => S4322,
        Y => S4326
    );
NOR_1285: ENTITY WORK.NOR
    PORT MAP (
        A => S4323,
        B => S4325,
        Y => S4327
    );
NAND_2809: ENTITY WORK.NAND
    PORT MAP (
        A => S4324,
        B => S4326,
        Y => S4328
    );
NOR_1286: ENTITY WORK.NOR
    PORT MAP (
        A => S4226,
        B => S4287,
        Y => S4329
    );
NOR_1287: ENTITY WORK.NOR
    PORT MAP (
        A => S4288,
        B => S4329,
        Y => S4330
    );
NOR_1288: ENTITY WORK.NOR
    PORT MAP (
        A => S4313,
        B => S4330,
        Y => S4331
    );
NOT_343: ENTITY WORK.NOT
    PORT MAP (
        A => S4331,
        Y => S4332
    );
NOR_1289: ENTITY WORK.NOR
    PORT MAP (
        A => S4220,
        B => S4314,
        Y => S4333
    );
NAND_2810: ENTITY WORK.NAND
    PORT MAP (
        A => S4221,
        B => S4313,
        Y => S4334
    );
NOR_1290: ENTITY WORK.NOR
    PORT MAP (
        A => S4331,
        B => S4333,
        Y => S4335
    );
NAND_2811: ENTITY WORK.NAND
    PORT MAP (
        A => S4332,
        B => S4334,
        Y => S4336
    );
NOR_1291: ENTITY WORK.NOR
    PORT MAP (
        A => S2106,
        B => S4336,
        Y => S4337
    );
NAND_2812: ENTITY WORK.NAND
    PORT MAP (
        A => S2107,
        B => S4335,
        Y => S4338
    );
NOR_1292: ENTITY WORK.NOR
    PORT MAP (
        A => S2107,
        B => S4335,
        Y => S4339
    );
NAND_2813: ENTITY WORK.NAND
    PORT MAP (
        A => S2106,
        B => S4336,
        Y => S4340
    );
NOR_1293: ENTITY WORK.NOR
    PORT MAP (
        A => S4337,
        B => S4339,
        Y => S4341
    );
NAND_2814: ENTITY WORK.NAND
    PORT MAP (
        A => S4338,
        B => S4340,
        Y => S4342
    );
NOR_1294: ENTITY WORK.NOR
    PORT MAP (
        A => S4242,
        B => S4283,
        Y => S4343
    );
NOR_1295: ENTITY WORK.NOR
    PORT MAP (
        A => S4284,
        B => S4343,
        Y => S4344
    );
NOR_1296: ENTITY WORK.NOR
    PORT MAP (
        A => S4313,
        B => S4344,
        Y => S4345
    );
NOT_344: ENTITY WORK.NOT
    PORT MAP (
        A => S4345,
        Y => S4346
    );
NOR_1297: ENTITY WORK.NOR
    PORT MAP (
        A => S4236,
        B => S4314,
        Y => S4347
    );
NAND_2815: ENTITY WORK.NAND
    PORT MAP (
        A => S4237,
        B => S4313,
        Y => S4348
    );
NOR_1298: ENTITY WORK.NOR
    PORT MAP (
        A => S4345,
        B => S4347,
        Y => S4349
    );
NAND_2816: ENTITY WORK.NAND
    PORT MAP (
        A => S4346,
        B => S4348,
        Y => S4350
    );
NOR_1299: ENTITY WORK.NOR
    PORT MAP (
        A => S1597,
        B => S4350,
        Y => S4351
    );
NAND_2817: ENTITY WORK.NAND
    PORT MAP (
        A => S1598,
        B => S4349,
        Y => S4352
    );
NOR_1300: ENTITY WORK.NOR
    PORT MAP (
        A => S1598,
        B => S4349,
        Y => S4353
    );
NAND_2818: ENTITY WORK.NAND
    PORT MAP (
        A => S1597,
        B => S4350,
        Y => S4354
    );
NOR_1301: ENTITY WORK.NOR
    PORT MAP (
        A => S4351,
        B => S4353,
        Y => S4355
    );
NAND_2819: ENTITY WORK.NAND
    PORT MAP (
        A => S4352,
        B => S4354,
        Y => S4356
    );
NOR_1302: ENTITY WORK.NOR
    PORT MAP (
        A => S4258,
        B => S4279,
        Y => S4357
    );
NOR_1303: ENTITY WORK.NOR
    PORT MAP (
        A => S4280,
        B => S4357,
        Y => S4358
    );
NOR_1304: ENTITY WORK.NOR
    PORT MAP (
        A => S4313,
        B => S4358,
        Y => S4359
    );
NOT_345: ENTITY WORK.NOT
    PORT MAP (
        A => S4359,
        Y => S4360
    );
NAND_2820: ENTITY WORK.NAND
    PORT MAP (
        A => S4253,
        B => S4313,
        Y => S4361
    );
NOT_346: ENTITY WORK.NOT
    PORT MAP (
        A => S4361,
        Y => S4362
    );
NOR_1305: ENTITY WORK.NOR
    PORT MAP (
        A => S4359,
        B => S4362,
        Y => S4363
    );
NAND_2821: ENTITY WORK.NAND
    PORT MAP (
        A => S4360,
        B => S4361,
        Y => S4364
    );
NOR_1306: ENTITY WORK.NOR
    PORT MAP (
        A => S1952,
        B => S4364,
        Y => S4365
    );
NAND_2822: ENTITY WORK.NAND
    PORT MAP (
        A => S1953,
        B => S4363,
        Y => S4366
    );
NOR_1307: ENTITY WORK.NOR
    PORT MAP (
        A => S1953,
        B => S4363,
        Y => S4367
    );
NAND_2823: ENTITY WORK.NAND
    PORT MAP (
        A => S1952,
        B => S4364,
        Y => S4368
    );
NOR_1308: ENTITY WORK.NOR
    PORT MAP (
        A => S4365,
        B => S4367,
        Y => S4369
    );
NAND_2824: ENTITY WORK.NAND
    PORT MAP (
        A => S4366,
        B => S4368,
        Y => S4370
    );
NOR_1309: ENTITY WORK.NOR
    PORT MAP (
        A => S4272,
        B => S4275,
        Y => S4371
    );
NOR_1310: ENTITY WORK.NOR
    PORT MAP (
        A => S4276,
        B => S4371,
        Y => S4372
    );
NOR_1311: ENTITY WORK.NOR
    PORT MAP (
        A => S4313,
        B => S4372,
        Y => S4373
    );
NOT_347: ENTITY WORK.NOT
    PORT MAP (
        A => S4373,
        Y => S4374
    );
NOR_1312: ENTITY WORK.NOR
    PORT MAP (
        A => S4266,
        B => S4314,
        Y => S4375
    );
NAND_2825: ENTITY WORK.NAND
    PORT MAP (
        A => S4267,
        B => S4313,
        Y => S4376
    );
NOR_1313: ENTITY WORK.NOR
    PORT MAP (
        A => S4373,
        B => S4375,
        Y => S4377
    );
NAND_2826: ENTITY WORK.NAND
    PORT MAP (
        A => S4374,
        B => S4376,
        Y => S4378
    );
NOR_1314: ENTITY WORK.NOR
    PORT MAP (
        A => S1848,
        B => S4378,
        Y => S4379
    );
NAND_2827: ENTITY WORK.NAND
    PORT MAP (
        A => S1849,
        B => S4377,
        Y => S4380
    );
NOR_1315: ENTITY WORK.NOR
    PORT MAP (
        A => S1849,
        B => S4377,
        Y => S4381
    );
NAND_2828: ENTITY WORK.NAND
    PORT MAP (
        A => S1848,
        B => S4378,
        Y => S4382
    );
NOR_1316: ENTITY WORK.NOR
    PORT MAP (
        A => S4379,
        B => S4381,
        Y => S4383
    );
NAND_2829: ENTITY WORK.NAND
    PORT MAP (
        A => S4380,
        B => S4382,
        Y => S4384
    );
NOR_1317: ENTITY WORK.NOR
    PORT MAP (
        A => S1516,
        B => S4313,
        Y => S4385
    );
NAND_2830: ENTITY WORK.NAND
    PORT MAP (
        A => S1515,
        B => S4314,
        Y => S4386
    );
NOR_1318: ENTITY WORK.NOR
    PORT MAP (
        A => S754,
        B => S4386,
        Y => S4387
    );
NAND_2831: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_9,
        B => S4385,
        Y => S4388
    );
NOR_1319: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_9,
        B => S4385,
        Y => S4389
    );
NAND_2832: ENTITY WORK.NAND
    PORT MAP (
        A => S754,
        B => S4386,
        Y => S4390
    );
NOR_1320: ENTITY WORK.NOR
    PORT MAP (
        A => S4387,
        B => S4389,
        Y => S4391
    );
NAND_2833: ENTITY WORK.NAND
    PORT MAP (
        A => S4388,
        B => S4390,
        Y => S4392
    );
NOR_1321: ENTITY WORK.NOR
    PORT MAP (
        A => S1745,
        B => S4392,
        Y => S4393
    );
NAND_2834: ENTITY WORK.NAND
    PORT MAP (
        A => S1746,
        B => S4391,
        Y => S4394
    );
NOR_1322: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_8,
        B => S1516,
        Y => S4395
    );
NAND_2835: ENTITY WORK.NAND
    PORT MAP (
        A => S805,
        B => S1515,
        Y => S4396
    );
NOR_1323: ENTITY WORK.NOR
    PORT MAP (
        A => S1746,
        B => S4391,
        Y => S4397
    );
NAND_2836: ENTITY WORK.NAND
    PORT MAP (
        A => S1745,
        B => S4392,
        Y => S4398
    );
NOR_1324: ENTITY WORK.NOR
    PORT MAP (
        A => S4393,
        B => S4397,
        Y => S4399
    );
NAND_2837: ENTITY WORK.NAND
    PORT MAP (
        A => S4394,
        B => S4398,
        Y => S4400
    );
NOR_1325: ENTITY WORK.NOR
    PORT MAP (
        A => S4395,
        B => S4400,
        Y => S4401
    );
NAND_2838: ENTITY WORK.NAND
    PORT MAP (
        A => S4396,
        B => S4399,
        Y => S4402
    );
NOR_1326: ENTITY WORK.NOR
    PORT MAP (
        A => S4393,
        B => S4401,
        Y => S4403
    );
NAND_2839: ENTITY WORK.NAND
    PORT MAP (
        A => S4394,
        B => S4402,
        Y => S4404
    );
NOR_1327: ENTITY WORK.NOR
    PORT MAP (
        A => S4384,
        B => S4403,
        Y => S4405
    );
NAND_2840: ENTITY WORK.NAND
    PORT MAP (
        A => S4383,
        B => S4404,
        Y => S4406
    );
NOR_1328: ENTITY WORK.NOR
    PORT MAP (
        A => S4379,
        B => S4405,
        Y => S4407
    );
NAND_2841: ENTITY WORK.NAND
    PORT MAP (
        A => S4380,
        B => S4406,
        Y => S4408
    );
NOR_1329: ENTITY WORK.NOR
    PORT MAP (
        A => S4370,
        B => S4407,
        Y => S4409
    );
NAND_2842: ENTITY WORK.NAND
    PORT MAP (
        A => S4369,
        B => S4408,
        Y => S4410
    );
NOR_1330: ENTITY WORK.NOR
    PORT MAP (
        A => S4365,
        B => S4409,
        Y => S4411
    );
NAND_2843: ENTITY WORK.NAND
    PORT MAP (
        A => S4366,
        B => S4410,
        Y => S4412
    );
NOR_1331: ENTITY WORK.NOR
    PORT MAP (
        A => S4356,
        B => S4411,
        Y => S4413
    );
NAND_2844: ENTITY WORK.NAND
    PORT MAP (
        A => S4355,
        B => S4412,
        Y => S4414
    );
NOR_1332: ENTITY WORK.NOR
    PORT MAP (
        A => S4351,
        B => S4413,
        Y => S4415
    );
NAND_2845: ENTITY WORK.NAND
    PORT MAP (
        A => S4352,
        B => S4414,
        Y => S4416
    );
NOR_1333: ENTITY WORK.NOR
    PORT MAP (
        A => S4342,
        B => S4415,
        Y => S4417
    );
NAND_2846: ENTITY WORK.NAND
    PORT MAP (
        A => S4341,
        B => S4416,
        Y => S4418
    );
NOR_1334: ENTITY WORK.NOR
    PORT MAP (
        A => S4337,
        B => S4417,
        Y => S4419
    );
NAND_2847: ENTITY WORK.NAND
    PORT MAP (
        A => S4338,
        B => S4418,
        Y => S4420
    );
NOR_1335: ENTITY WORK.NOR
    PORT MAP (
        A => S4328,
        B => S4419,
        Y => S4421
    );
NAND_2848: ENTITY WORK.NAND
    PORT MAP (
        A => S4327,
        B => S4420,
        Y => S4422
    );
NOR_1336: ENTITY WORK.NOR
    PORT MAP (
        A => S4323,
        B => S4421,
        Y => S4423
    );
NAND_2849: ENTITY WORK.NAND
    PORT MAP (
        A => S4324,
        B => S4422,
        Y => S4424
    );
NOR_1337: ENTITY WORK.NOR
    PORT MAP (
        A => S4306,
        B => S4423,
        Y => S4425
    );
NAND_2850: ENTITY WORK.NAND
    PORT MAP (
        A => S4305,
        B => S4424,
        Y => S4426
    );
NOR_1338: ENTITY WORK.NOR
    PORT MAP (
        A => S4302,
        B => S4425,
        Y => S4427
    );
NAND_2851: ENTITY WORK.NAND
    PORT MAP (
        A => S4303,
        B => S4426,
        Y => S4428
    );
NOR_1339: ENTITY WORK.NOR
    PORT MAP (
        A => S3913,
        B => S4427,
        Y => S4429
    );
NAND_2852: ENTITY WORK.NAND
    PORT MAP (
        A => S3912,
        B => S4428,
        Y => S4430
    );
NOR_1340: ENTITY WORK.NOR
    PORT MAP (
        A => S4327,
        B => S4420,
        Y => S4431
    );
NAND_2853: ENTITY WORK.NAND
    PORT MAP (
        A => S4328,
        B => S4419,
        Y => S4432
    );
NOR_1341: ENTITY WORK.NOR
    PORT MAP (
        A => S4421,
        B => S4431,
        Y => S4433
    );
NAND_2854: ENTITY WORK.NAND
    PORT MAP (
        A => S4422,
        B => S4432,
        Y => S4434
    );
NOR_1342: ENTITY WORK.NOR
    PORT MAP (
        A => S4430,
        B => S4433,
        Y => S4435
    );
NAND_2855: ENTITY WORK.NAND
    PORT MAP (
        A => S4429,
        B => S4434,
        Y => S4436
    );
NOR_1343: ENTITY WORK.NOR
    PORT MAP (
        A => S4321,
        B => S4429,
        Y => S4437
    );
NAND_2856: ENTITY WORK.NAND
    PORT MAP (
        A => S4322,
        B => S4430,
        Y => S4438
    );
NOR_1344: ENTITY WORK.NOR
    PORT MAP (
        A => S4435,
        B => S4437,
        Y => S4439
    );
NAND_2857: ENTITY WORK.NAND
    PORT MAP (
        A => S4436,
        B => S4438,
        Y => S4440
    );
NOR_1345: ENTITY WORK.NOR
    PORT MAP (
        A => S2311,
        B => S4440,
        Y => S4441
    );
NAND_2858: ENTITY WORK.NAND
    PORT MAP (
        A => S2312,
        B => S4439,
        Y => S4442
    );
NOR_1346: ENTITY WORK.NOR
    PORT MAP (
        A => S2312,
        B => S4439,
        Y => S4443
    );
NAND_2859: ENTITY WORK.NAND
    PORT MAP (
        A => S2311,
        B => S4440,
        Y => S4444
    );
NOR_1347: ENTITY WORK.NOR
    PORT MAP (
        A => S4441,
        B => S4443,
        Y => S4445
    );
NAND_2860: ENTITY WORK.NAND
    PORT MAP (
        A => S4442,
        B => S4444,
        Y => S4446
    );
NAND_2861: ENTITY WORK.NAND
    PORT MAP (
        A => S4342,
        B => S4415,
        Y => S4447
    );
NAND_2862: ENTITY WORK.NAND
    PORT MAP (
        A => S4418,
        B => S4447,
        Y => S4448
    );
NAND_2863: ENTITY WORK.NAND
    PORT MAP (
        A => S4429,
        B => S4448,
        Y => S4449
    );
NAND_2864: ENTITY WORK.NAND
    PORT MAP (
        A => S4336,
        B => S4430,
        Y => S4450
    );
NAND_2865: ENTITY WORK.NAND
    PORT MAP (
        A => S4449,
        B => S4450,
        Y => S4451
    );
NOT_348: ENTITY WORK.NOT
    PORT MAP (
        A => S4451,
        Y => S4452
    );
NAND_2866: ENTITY WORK.NAND
    PORT MAP (
        A => S2206,
        B => S4452,
        Y => S4453
    );
NAND_2867: ENTITY WORK.NAND
    PORT MAP (
        A => S2205,
        B => S4451,
        Y => S4454
    );
NAND_2868: ENTITY WORK.NAND
    PORT MAP (
        A => S4356,
        B => S4411,
        Y => S4455
    );
NAND_2869: ENTITY WORK.NAND
    PORT MAP (
        A => S4414,
        B => S4455,
        Y => S4456
    );
NAND_2870: ENTITY WORK.NAND
    PORT MAP (
        A => S4429,
        B => S4456,
        Y => S4457
    );
NAND_2871: ENTITY WORK.NAND
    PORT MAP (
        A => S4350,
        B => S4430,
        Y => S4458
    );
NAND_2872: ENTITY WORK.NAND
    PORT MAP (
        A => S4457,
        B => S4458,
        Y => S4459
    );
NOT_349: ENTITY WORK.NOT
    PORT MAP (
        A => S4459,
        Y => S4460
    );
NOR_1348: ENTITY WORK.NOR
    PORT MAP (
        A => S2106,
        B => S4459,
        Y => S4461
    );
NAND_2873: ENTITY WORK.NAND
    PORT MAP (
        A => S2107,
        B => S4460,
        Y => S4462
    );
NAND_2874: ENTITY WORK.NAND
    PORT MAP (
        A => S2106,
        B => S4459,
        Y => S4463
    );
NOT_350: ENTITY WORK.NOT
    PORT MAP (
        A => S4463,
        Y => S4464
    );
NOR_1349: ENTITY WORK.NOR
    PORT MAP (
        A => S4461,
        B => S4464,
        Y => S4465
    );
NOT_351: ENTITY WORK.NOT
    PORT MAP (
        A => S4465,
        Y => S4466
    );
NOR_1350: ENTITY WORK.NOR
    PORT MAP (
        A => S4363,
        B => S4429,
        Y => S4467
    );
NAND_2875: ENTITY WORK.NAND
    PORT MAP (
        A => S4364,
        B => S4430,
        Y => S4468
    );
NOR_1351: ENTITY WORK.NOR
    PORT MAP (
        A => S4369,
        B => S4408,
        Y => S4469
    );
NAND_2876: ENTITY WORK.NAND
    PORT MAP (
        A => S4370,
        B => S4407,
        Y => S4470
    );
NOR_1352: ENTITY WORK.NOR
    PORT MAP (
        A => S4409,
        B => S4469,
        Y => S4471
    );
NAND_2877: ENTITY WORK.NAND
    PORT MAP (
        A => S4410,
        B => S4470,
        Y => S4472
    );
NOR_1353: ENTITY WORK.NOR
    PORT MAP (
        A => S4430,
        B => S4471,
        Y => S4473
    );
NAND_2878: ENTITY WORK.NAND
    PORT MAP (
        A => S4429,
        B => S4472,
        Y => S4474
    );
NOR_1354: ENTITY WORK.NOR
    PORT MAP (
        A => S4467,
        B => S4473,
        Y => S4475
    );
NAND_2879: ENTITY WORK.NAND
    PORT MAP (
        A => S4468,
        B => S4474,
        Y => S4476
    );
NOR_1355: ENTITY WORK.NOR
    PORT MAP (
        A => S1597,
        B => S4476,
        Y => S4477
    );
NAND_2880: ENTITY WORK.NAND
    PORT MAP (
        A => S1598,
        B => S4475,
        Y => S4478
    );
NOR_1356: ENTITY WORK.NOR
    PORT MAP (
        A => S1598,
        B => S4475,
        Y => S4479
    );
NAND_2881: ENTITY WORK.NAND
    PORT MAP (
        A => S1597,
        B => S4476,
        Y => S4480
    );
NOR_1357: ENTITY WORK.NOR
    PORT MAP (
        A => S4477,
        B => S4479,
        Y => S4481
    );
NAND_2882: ENTITY WORK.NAND
    PORT MAP (
        A => S4478,
        B => S4480,
        Y => S4482
    );
NOR_1358: ENTITY WORK.NOR
    PORT MAP (
        A => S4383,
        B => S4404,
        Y => S4483
    );
NAND_2883: ENTITY WORK.NAND
    PORT MAP (
        A => S4384,
        B => S4403,
        Y => S4484
    );
NOR_1359: ENTITY WORK.NOR
    PORT MAP (
        A => S4405,
        B => S4483,
        Y => S4485
    );
NAND_2884: ENTITY WORK.NAND
    PORT MAP (
        A => S4406,
        B => S4484,
        Y => S4486
    );
NOR_1360: ENTITY WORK.NOR
    PORT MAP (
        A => S4430,
        B => S4485,
        Y => S4487
    );
NAND_2885: ENTITY WORK.NAND
    PORT MAP (
        A => S4429,
        B => S4486,
        Y => S4488
    );
NOR_1361: ENTITY WORK.NOR
    PORT MAP (
        A => S4377,
        B => S4429,
        Y => S4489
    );
NAND_2886: ENTITY WORK.NAND
    PORT MAP (
        A => S4378,
        B => S4430,
        Y => S4490
    );
NOR_1362: ENTITY WORK.NOR
    PORT MAP (
        A => S4487,
        B => S4489,
        Y => S4491
    );
NAND_2887: ENTITY WORK.NAND
    PORT MAP (
        A => S4488,
        B => S4490,
        Y => S4492
    );
NOR_1363: ENTITY WORK.NOR
    PORT MAP (
        A => S1952,
        B => S4492,
        Y => S4493
    );
NAND_2888: ENTITY WORK.NAND
    PORT MAP (
        A => S1953,
        B => S4491,
        Y => S4494
    );
NOR_1364: ENTITY WORK.NOR
    PORT MAP (
        A => S1953,
        B => S4491,
        Y => S4495
    );
NAND_2889: ENTITY WORK.NAND
    PORT MAP (
        A => S1952,
        B => S4492,
        Y => S4496
    );
NOR_1365: ENTITY WORK.NOR
    PORT MAP (
        A => S4493,
        B => S4495,
        Y => S4497
    );
NAND_2890: ENTITY WORK.NAND
    PORT MAP (
        A => S4494,
        B => S4496,
        Y => S4498
    );
NOR_1366: ENTITY WORK.NOR
    PORT MAP (
        A => S4396,
        B => S4399,
        Y => S4499
    );
NAND_2891: ENTITY WORK.NAND
    PORT MAP (
        A => S4395,
        B => S4400,
        Y => S4500
    );
NOR_1367: ENTITY WORK.NOR
    PORT MAP (
        A => S4401,
        B => S4499,
        Y => S4501
    );
NAND_2892: ENTITY WORK.NAND
    PORT MAP (
        A => S4402,
        B => S4500,
        Y => S4502
    );
NOR_1368: ENTITY WORK.NOR
    PORT MAP (
        A => S4430,
        B => S4501,
        Y => S4503
    );
NAND_2893: ENTITY WORK.NAND
    PORT MAP (
        A => S4429,
        B => S4502,
        Y => S4504
    );
NOR_1369: ENTITY WORK.NOR
    PORT MAP (
        A => S4391,
        B => S4429,
        Y => S4505
    );
NAND_2894: ENTITY WORK.NAND
    PORT MAP (
        A => S4392,
        B => S4430,
        Y => S4506
    );
NOR_1370: ENTITY WORK.NOR
    PORT MAP (
        A => S4503,
        B => S4505,
        Y => S4507
    );
NAND_2895: ENTITY WORK.NAND
    PORT MAP (
        A => S4504,
        B => S4506,
        Y => S4508
    );
NOR_1371: ENTITY WORK.NOR
    PORT MAP (
        A => S1848,
        B => S4508,
        Y => S4509
    );
NAND_2896: ENTITY WORK.NAND
    PORT MAP (
        A => S1849,
        B => S4507,
        Y => S4510
    );
NOR_1372: ENTITY WORK.NOR
    PORT MAP (
        A => S1849,
        B => S4507,
        Y => S4511
    );
NAND_2897: ENTITY WORK.NAND
    PORT MAP (
        A => S1848,
        B => S4508,
        Y => S4512
    );
NOR_1373: ENTITY WORK.NOR
    PORT MAP (
        A => S4509,
        B => S4511,
        Y => S4513
    );
NAND_2898: ENTITY WORK.NAND
    PORT MAP (
        A => S4510,
        B => S4512,
        Y => S4514
    );
NOR_1374: ENTITY WORK.NOR
    PORT MAP (
        A => S1516,
        B => S4430,
        Y => S4515
    );
NAND_2899: ENTITY WORK.NAND
    PORT MAP (
        A => S1515,
        B => S4429,
        Y => S4516
    );
NOR_1375: ENTITY WORK.NOR
    PORT MAP (
        A => S805,
        B => S4515,
        Y => S4517
    );
NAND_2900: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_8,
        B => S4516,
        Y => S4518
    );
NOR_1376: ENTITY WORK.NOR
    PORT MAP (
        A => S4396,
        B => S4430,
        Y => S4519
    );
NAND_2901: ENTITY WORK.NAND
    PORT MAP (
        A => S4395,
        B => S4429,
        Y => S4520
    );
NOR_1377: ENTITY WORK.NOR
    PORT MAP (
        A => S4517,
        B => S4519,
        Y => S4521
    );
NAND_2902: ENTITY WORK.NAND
    PORT MAP (
        A => S4518,
        B => S4520,
        Y => S4522
    );
NOR_1378: ENTITY WORK.NOR
    PORT MAP (
        A => S1745,
        B => S4521,
        Y => S4523
    );
NAND_2903: ENTITY WORK.NAND
    PORT MAP (
        A => S1746,
        B => S4522,
        Y => S4524
    );
NAND_2904: ENTITY WORK.NAND
    PORT MAP (
        A => S858,
        B => S1515,
        Y => S4525
    );
NOT_352: ENTITY WORK.NOT
    PORT MAP (
        A => S4525,
        Y => S4526
    );
NOR_1379: ENTITY WORK.NOR
    PORT MAP (
        A => S1746,
        B => S4522,
        Y => S4527
    );
NAND_2905: ENTITY WORK.NAND
    PORT MAP (
        A => S1745,
        B => S4521,
        Y => S4528
    );
NOR_1380: ENTITY WORK.NOR
    PORT MAP (
        A => S4523,
        B => S4527,
        Y => S4529
    );
NAND_2906: ENTITY WORK.NAND
    PORT MAP (
        A => S4524,
        B => S4528,
        Y => S4530
    );
NOR_1381: ENTITY WORK.NOR
    PORT MAP (
        A => S4526,
        B => S4530,
        Y => S4531
    );
NAND_2907: ENTITY WORK.NAND
    PORT MAP (
        A => S4525,
        B => S4529,
        Y => S4532
    );
NOR_1382: ENTITY WORK.NOR
    PORT MAP (
        A => S4523,
        B => S4531,
        Y => S4533
    );
NAND_2908: ENTITY WORK.NAND
    PORT MAP (
        A => S4524,
        B => S4532,
        Y => S4534
    );
NOR_1383: ENTITY WORK.NOR
    PORT MAP (
        A => S4514,
        B => S4533,
        Y => S4535
    );
NAND_2909: ENTITY WORK.NAND
    PORT MAP (
        A => S4513,
        B => S4534,
        Y => S4536
    );
NOR_1384: ENTITY WORK.NOR
    PORT MAP (
        A => S4509,
        B => S4535,
        Y => S4537
    );
NAND_2910: ENTITY WORK.NAND
    PORT MAP (
        A => S4510,
        B => S4536,
        Y => S4538
    );
NOR_1385: ENTITY WORK.NOR
    PORT MAP (
        A => S4498,
        B => S4537,
        Y => S4539
    );
NAND_2911: ENTITY WORK.NAND
    PORT MAP (
        A => S4497,
        B => S4538,
        Y => S4540
    );
NOR_1386: ENTITY WORK.NOR
    PORT MAP (
        A => S4493,
        B => S4539,
        Y => S4541
    );
NAND_2912: ENTITY WORK.NAND
    PORT MAP (
        A => S4494,
        B => S4540,
        Y => S4542
    );
NOR_1387: ENTITY WORK.NOR
    PORT MAP (
        A => S4482,
        B => S4541,
        Y => S4543
    );
NAND_2913: ENTITY WORK.NAND
    PORT MAP (
        A => S4481,
        B => S4542,
        Y => S4544
    );
NOR_1388: ENTITY WORK.NOR
    PORT MAP (
        A => S4477,
        B => S4543,
        Y => S4545
    );
NAND_2914: ENTITY WORK.NAND
    PORT MAP (
        A => S4478,
        B => S4544,
        Y => S4546
    );
NOR_1389: ENTITY WORK.NOR
    PORT MAP (
        A => S4466,
        B => S4545,
        Y => S4547
    );
NAND_2915: ENTITY WORK.NAND
    PORT MAP (
        A => S4465,
        B => S4546,
        Y => S4548
    );
NOR_1390: ENTITY WORK.NOR
    PORT MAP (
        A => S4461,
        B => S4547,
        Y => S4549
    );
NAND_2916: ENTITY WORK.NAND
    PORT MAP (
        A => S4462,
        B => S4548,
        Y => S4550
    );
NAND_2917: ENTITY WORK.NAND
    PORT MAP (
        A => S4454,
        B => S4550,
        Y => S4551
    );
NAND_2918: ENTITY WORK.NAND
    PORT MAP (
        A => S4453,
        B => S4549,
        Y => S4552
    );
NAND_2919: ENTITY WORK.NAND
    PORT MAP (
        A => S4454,
        B => S4552,
        Y => S4553
    );
NAND_2920: ENTITY WORK.NAND
    PORT MAP (
        A => S4453,
        B => S4551,
        Y => S4554
    );
NOR_1391: ENTITY WORK.NOR
    PORT MAP (
        A => S4446,
        B => S4553,
        Y => S4555
    );
NAND_2921: ENTITY WORK.NAND
    PORT MAP (
        A => S4445,
        B => S4554,
        Y => S4556
    );
NOR_1392: ENTITY WORK.NOR
    PORT MAP (
        A => S4441,
        B => S4555,
        Y => S4557
    );
NAND_2922: ENTITY WORK.NAND
    PORT MAP (
        A => S4442,
        B => S4556,
        Y => S4558
    );
NOR_1393: ENTITY WORK.NOR
    PORT MAP (
        A => S4300,
        B => S4429,
        Y => S4559
    );
NOR_1394: ENTITY WORK.NOR
    PORT MAP (
        A => S3950,
        B => S4559,
        Y => S4560
    );
NOT_353: ENTITY WORK.NOT
    PORT MAP (
        A => S4560,
        Y => S4561
    );
NOR_1395: ENTITY WORK.NOR
    PORT MAP (
        A => S2417,
        B => S4560,
        Y => S4562
    );
NAND_2923: ENTITY WORK.NAND
    PORT MAP (
        A => S2418,
        B => S4561,
        Y => S4563
    );
NOR_1396: ENTITY WORK.NOR
    PORT MAP (
        A => S4558,
        B => S4562,
        Y => S4564
    );
NAND_2924: ENTITY WORK.NAND
    PORT MAP (
        A => S4557,
        B => S4563,
        Y => S4565
    );
NOR_1397: ENTITY WORK.NOR
    PORT MAP (
        A => S2418,
        B => S4561,
        Y => S4566
    );
NAND_2925: ENTITY WORK.NAND
    PORT MAP (
        A => S2417,
        B => S4560,
        Y => S4567
    );
NOR_1398: ENTITY WORK.NOR
    PORT MAP (
        A => S3911,
        B => S4566,
        Y => S4568
    );
NAND_2926: ENTITY WORK.NAND
    PORT MAP (
        A => S3910,
        B => S4567,
        Y => S4569
    );
NOR_1399: ENTITY WORK.NOR
    PORT MAP (
        A => S4564,
        B => S4569,
        Y => S4570
    );
NAND_2927: ENTITY WORK.NAND
    PORT MAP (
        A => S4565,
        B => S4568,
        Y => S4571
    );
NOR_1400: ENTITY WORK.NOR
    PORT MAP (
        A => S4445,
        B => S4554,
        Y => S4572
    );
NOR_1401: ENTITY WORK.NOR
    PORT MAP (
        A => S4555,
        B => S4572,
        Y => S4573
    );
NOR_1402: ENTITY WORK.NOR
    PORT MAP (
        A => S4571,
        B => S4573,
        Y => S4574
    );
NOR_1403: ENTITY WORK.NOR
    PORT MAP (
        A => S4439,
        B => S4570,
        Y => S4575
    );
NOR_1404: ENTITY WORK.NOR
    PORT MAP (
        A => S4574,
        B => S4575,
        Y => S4576
    );
NOT_354: ENTITY WORK.NOT
    PORT MAP (
        A => S4576,
        Y => S4577
    );
NOR_1405: ENTITY WORK.NOR
    PORT MAP (
        A => S2417,
        B => S4577,
        Y => S4578
    );
NAND_2928: ENTITY WORK.NAND
    PORT MAP (
        A => S2418,
        B => S4576,
        Y => S4579
    );
NOR_1406: ENTITY WORK.NOR
    PORT MAP (
        A => S2418,
        B => S4576,
        Y => S4580
    );
NOT_355: ENTITY WORK.NOT
    PORT MAP (
        A => S4580,
        Y => S4581
    );
NAND_2929: ENTITY WORK.NAND
    PORT MAP (
        A => S4579,
        B => S4581,
        Y => S4582
    );
NOT_356: ENTITY WORK.NOT
    PORT MAP (
        A => S4582,
        Y => S4583
    );
NAND_2930: ENTITY WORK.NAND
    PORT MAP (
        A => S4453,
        B => S4454,
        Y => S4584
    );
NAND_2931: ENTITY WORK.NAND
    PORT MAP (
        A => S4549,
        B => S4584,
        Y => S4585
    );
NOT_357: ENTITY WORK.NOT
    PORT MAP (
        A => S4585,
        Y => S4586
    );
NOR_1407: ENTITY WORK.NOR
    PORT MAP (
        A => S4549,
        B => S4584,
        Y => S4587
    );
NOR_1408: ENTITY WORK.NOR
    PORT MAP (
        A => S4586,
        B => S4587,
        Y => S4588
    );
NOR_1409: ENTITY WORK.NOR
    PORT MAP (
        A => S4571,
        B => S4588,
        Y => S4589
    );
NOR_1410: ENTITY WORK.NOR
    PORT MAP (
        A => S4452,
        B => S4570,
        Y => S4590
    );
NOR_1411: ENTITY WORK.NOR
    PORT MAP (
        A => S4589,
        B => S4590,
        Y => S4591
    );
NOT_358: ENTITY WORK.NOT
    PORT MAP (
        A => S4591,
        Y => S4592
    );
NOR_1412: ENTITY WORK.NOR
    PORT MAP (
        A => S2311,
        B => S4592,
        Y => S4593
    );
NOR_1413: ENTITY WORK.NOR
    PORT MAP (
        A => S2312,
        B => S4591,
        Y => S4594
    );
NOR_1414: ENTITY WORK.NOR
    PORT MAP (
        A => S4465,
        B => S4546,
        Y => S4595
    );
NOR_1415: ENTITY WORK.NOR
    PORT MAP (
        A => S4547,
        B => S4595,
        Y => S4596
    );
NOR_1416: ENTITY WORK.NOR
    PORT MAP (
        A => S4571,
        B => S4596,
        Y => S4597
    );
NOR_1417: ENTITY WORK.NOR
    PORT MAP (
        A => S4460,
        B => S4570,
        Y => S4598
    );
NOR_1418: ENTITY WORK.NOR
    PORT MAP (
        A => S4597,
        B => S4598,
        Y => S4599
    );
NOT_359: ENTITY WORK.NOT
    PORT MAP (
        A => S4599,
        Y => S4600
    );
NOR_1419: ENTITY WORK.NOR
    PORT MAP (
        A => S2205,
        B => S4600,
        Y => S4601
    );
NAND_2932: ENTITY WORK.NAND
    PORT MAP (
        A => S2206,
        B => S4599,
        Y => S4602
    );
NAND_2933: ENTITY WORK.NAND
    PORT MAP (
        A => S2205,
        B => S4600,
        Y => S4603
    );
NAND_2934: ENTITY WORK.NAND
    PORT MAP (
        A => S4602,
        B => S4603,
        Y => S4604
    );
NOT_360: ENTITY WORK.NOT
    PORT MAP (
        A => S4604,
        Y => S4605
    );
NOR_1420: ENTITY WORK.NOR
    PORT MAP (
        A => S4481,
        B => S4542,
        Y => S4606
    );
NOR_1421: ENTITY WORK.NOR
    PORT MAP (
        A => S4543,
        B => S4606,
        Y => S4607
    );
NOR_1422: ENTITY WORK.NOR
    PORT MAP (
        A => S4571,
        B => S4607,
        Y => S4608
    );
NOR_1423: ENTITY WORK.NOR
    PORT MAP (
        A => S4475,
        B => S4570,
        Y => S4609
    );
NOR_1424: ENTITY WORK.NOR
    PORT MAP (
        A => S4608,
        B => S4609,
        Y => S4610
    );
NOT_361: ENTITY WORK.NOT
    PORT MAP (
        A => S4610,
        Y => S4611
    );
NOR_1425: ENTITY WORK.NOR
    PORT MAP (
        A => S2106,
        B => S4611,
        Y => S4612
    );
NAND_2935: ENTITY WORK.NAND
    PORT MAP (
        A => S2107,
        B => S4610,
        Y => S4613
    );
NAND_2936: ENTITY WORK.NAND
    PORT MAP (
        A => S2106,
        B => S4611,
        Y => S4614
    );
NAND_2937: ENTITY WORK.NAND
    PORT MAP (
        A => S4613,
        B => S4614,
        Y => S4615
    );
NOT_362: ENTITY WORK.NOT
    PORT MAP (
        A => S4615,
        Y => S4616
    );
NOR_1426: ENTITY WORK.NOR
    PORT MAP (
        A => S4491,
        B => S4570,
        Y => S4617
    );
NOR_1427: ENTITY WORK.NOR
    PORT MAP (
        A => S4497,
        B => S4538,
        Y => S4618
    );
NOR_1428: ENTITY WORK.NOR
    PORT MAP (
        A => S4539,
        B => S4618,
        Y => S4619
    );
NOR_1429: ENTITY WORK.NOR
    PORT MAP (
        A => S4571,
        B => S4619,
        Y => S4620
    );
NOR_1430: ENTITY WORK.NOR
    PORT MAP (
        A => S4617,
        B => S4620,
        Y => S4621
    );
NOT_363: ENTITY WORK.NOT
    PORT MAP (
        A => S4621,
        Y => S4622
    );
NOR_1431: ENTITY WORK.NOR
    PORT MAP (
        A => S1597,
        B => S4622,
        Y => S4623
    );
NAND_2938: ENTITY WORK.NAND
    PORT MAP (
        A => S1598,
        B => S4621,
        Y => S4624
    );
NAND_2939: ENTITY WORK.NAND
    PORT MAP (
        A => S1597,
        B => S4622,
        Y => S4625
    );
NAND_2940: ENTITY WORK.NAND
    PORT MAP (
        A => S4624,
        B => S4625,
        Y => S4626
    );
NOT_364: ENTITY WORK.NOT
    PORT MAP (
        A => S4626,
        Y => S4627
    );
NOR_1432: ENTITY WORK.NOR
    PORT MAP (
        A => S4513,
        B => S4534,
        Y => S4628
    );
NOR_1433: ENTITY WORK.NOR
    PORT MAP (
        A => S4535,
        B => S4628,
        Y => S4629
    );
NOR_1434: ENTITY WORK.NOR
    PORT MAP (
        A => S4571,
        B => S4629,
        Y => S4630
    );
NOR_1435: ENTITY WORK.NOR
    PORT MAP (
        A => S4507,
        B => S4570,
        Y => S4631
    );
NOR_1436: ENTITY WORK.NOR
    PORT MAP (
        A => S4630,
        B => S4631,
        Y => S4632
    );
NOT_365: ENTITY WORK.NOT
    PORT MAP (
        A => S4632,
        Y => S4633
    );
NAND_2941: ENTITY WORK.NAND
    PORT MAP (
        A => S1953,
        B => S4632,
        Y => S4634
    );
NAND_2942: ENTITY WORK.NAND
    PORT MAP (
        A => S1952,
        B => S4633,
        Y => S4635
    );
NOR_1437: ENTITY WORK.NOR
    PORT MAP (
        A => S4525,
        B => S4529,
        Y => S4636
    );
NOR_1438: ENTITY WORK.NOR
    PORT MAP (
        A => S4531,
        B => S4636,
        Y => S4637
    );
NOR_1439: ENTITY WORK.NOR
    PORT MAP (
        A => S4571,
        B => S4637,
        Y => S4638
    );
NOR_1440: ENTITY WORK.NOR
    PORT MAP (
        A => S4522,
        B => S4570,
        Y => S4639
    );
NOR_1441: ENTITY WORK.NOR
    PORT MAP (
        A => S4638,
        B => S4639,
        Y => S4640
    );
NOT_366: ENTITY WORK.NOT
    PORT MAP (
        A => S4640,
        Y => S4641
    );
NOR_1442: ENTITY WORK.NOR
    PORT MAP (
        A => S1848,
        B => S4641,
        Y => S4642
    );
NAND_2943: ENTITY WORK.NAND
    PORT MAP (
        A => S1849,
        B => S4640,
        Y => S4643
    );
NOR_1443: ENTITY WORK.NOR
    PORT MAP (
        A => S1516,
        B => S4571,
        Y => S4644
    );
NAND_2944: ENTITY WORK.NAND
    PORT MAP (
        A => S1515,
        B => S4570,
        Y => S4645
    );
NOR_1444: ENTITY WORK.NOR
    PORT MAP (
        A => S858,
        B => S4644,
        Y => S4646
    );
NAND_2945: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_7,
        B => S4645,
        Y => S4647
    );
NOR_1445: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_7,
        B => S4645,
        Y => S4648
    );
NAND_2946: ENTITY WORK.NAND
    PORT MAP (
        A => S858,
        B => S4644,
        Y => S4649
    );
NOR_1446: ENTITY WORK.NOR
    PORT MAP (
        A => S4646,
        B => S4648,
        Y => S4650
    );
NAND_2947: ENTITY WORK.NAND
    PORT MAP (
        A => S4647,
        B => S4649,
        Y => S4651
    );
NOR_1447: ENTITY WORK.NOR
    PORT MAP (
        A => S1745,
        B => S4650,
        Y => S4652
    );
NAND_2948: ENTITY WORK.NAND
    PORT MAP (
        A => S1746,
        B => S4651,
        Y => S4653
    );
NAND_2949: ENTITY WORK.NAND
    PORT MAP (
        A => S910,
        B => S1515,
        Y => S4654
    );
NOT_367: ENTITY WORK.NOT
    PORT MAP (
        A => S4654,
        Y => S4655
    );
NOR_1448: ENTITY WORK.NOR
    PORT MAP (
        A => S1746,
        B => S4651,
        Y => S4656
    );
NAND_2950: ENTITY WORK.NAND
    PORT MAP (
        A => S1745,
        B => S4650,
        Y => S4657
    );
NOR_1449: ENTITY WORK.NOR
    PORT MAP (
        A => S4652,
        B => S4656,
        Y => S4658
    );
NAND_2951: ENTITY WORK.NAND
    PORT MAP (
        A => S4653,
        B => S4657,
        Y => S4659
    );
NOR_1450: ENTITY WORK.NOR
    PORT MAP (
        A => S4655,
        B => S4659,
        Y => S4660
    );
NAND_2952: ENTITY WORK.NAND
    PORT MAP (
        A => S4654,
        B => S4658,
        Y => S4661
    );
NOR_1451: ENTITY WORK.NOR
    PORT MAP (
        A => S4652,
        B => S4660,
        Y => S4662
    );
NAND_2953: ENTITY WORK.NAND
    PORT MAP (
        A => S4653,
        B => S4661,
        Y => S4663
    );
NAND_2954: ENTITY WORK.NAND
    PORT MAP (
        A => S1848,
        B => S4641,
        Y => S4664
    );
NAND_2955: ENTITY WORK.NAND
    PORT MAP (
        A => S4643,
        B => S4664,
        Y => S4665
    );
NOT_368: ENTITY WORK.NOT
    PORT MAP (
        A => S4665,
        Y => S4666
    );
NOR_1452: ENTITY WORK.NOR
    PORT MAP (
        A => S4662,
        B => S4665,
        Y => S4667
    );
NAND_2956: ENTITY WORK.NAND
    PORT MAP (
        A => S4663,
        B => S4666,
        Y => S4668
    );
NOR_1453: ENTITY WORK.NOR
    PORT MAP (
        A => S4642,
        B => S4667,
        Y => S4669
    );
NAND_2957: ENTITY WORK.NAND
    PORT MAP (
        A => S4643,
        B => S4668,
        Y => S4670
    );
NAND_2958: ENTITY WORK.NAND
    PORT MAP (
        A => S4635,
        B => S4670,
        Y => S4671
    );
NAND_2959: ENTITY WORK.NAND
    PORT MAP (
        A => S4634,
        B => S4669,
        Y => S4672
    );
NAND_2960: ENTITY WORK.NAND
    PORT MAP (
        A => S4635,
        B => S4672,
        Y => S4673
    );
NAND_2961: ENTITY WORK.NAND
    PORT MAP (
        A => S4634,
        B => S4671,
        Y => S4674
    );
NOR_1454: ENTITY WORK.NOR
    PORT MAP (
        A => S4626,
        B => S4673,
        Y => S4675
    );
NAND_2962: ENTITY WORK.NAND
    PORT MAP (
        A => S4627,
        B => S4674,
        Y => S4676
    );
NOR_1455: ENTITY WORK.NOR
    PORT MAP (
        A => S4623,
        B => S4675,
        Y => S4677
    );
NAND_2963: ENTITY WORK.NAND
    PORT MAP (
        A => S4624,
        B => S4676,
        Y => S4678
    );
NOR_1456: ENTITY WORK.NOR
    PORT MAP (
        A => S4615,
        B => S4677,
        Y => S4679
    );
NAND_2964: ENTITY WORK.NAND
    PORT MAP (
        A => S4616,
        B => S4678,
        Y => S4680
    );
NOR_1457: ENTITY WORK.NOR
    PORT MAP (
        A => S4612,
        B => S4679,
        Y => S4681
    );
NAND_2965: ENTITY WORK.NAND
    PORT MAP (
        A => S4613,
        B => S4680,
        Y => S4682
    );
NOR_1458: ENTITY WORK.NOR
    PORT MAP (
        A => S4604,
        B => S4681,
        Y => S4683
    );
NAND_2966: ENTITY WORK.NAND
    PORT MAP (
        A => S4605,
        B => S4682,
        Y => S4684
    );
NOR_1459: ENTITY WORK.NOR
    PORT MAP (
        A => S4601,
        B => S4683,
        Y => S4685
    );
NAND_2967: ENTITY WORK.NAND
    PORT MAP (
        A => S4602,
        B => S4684,
        Y => S4686
    );
NOR_1460: ENTITY WORK.NOR
    PORT MAP (
        A => S4594,
        B => S4685,
        Y => S4687
    );
NOR_1461: ENTITY WORK.NOR
    PORT MAP (
        A => S4593,
        B => S4686,
        Y => S4688
    );
NOR_1462: ENTITY WORK.NOR
    PORT MAP (
        A => S4593,
        B => S4687,
        Y => S4689
    );
NOR_1463: ENTITY WORK.NOR
    PORT MAP (
        A => S4594,
        B => S4688,
        Y => S4690
    );
NOR_1464: ENTITY WORK.NOR
    PORT MAP (
        A => S4582,
        B => S4689,
        Y => S4691
    );
NAND_2968: ENTITY WORK.NAND
    PORT MAP (
        A => S4583,
        B => S4690,
        Y => S4692
    );
NOR_1465: ENTITY WORK.NOR
    PORT MAP (
        A => S4578,
        B => S4691,
        Y => S4693
    );
NAND_2969: ENTITY WORK.NAND
    PORT MAP (
        A => S4579,
        B => S4692,
        Y => S4694
    );
NOR_1466: ENTITY WORK.NOR
    PORT MAP (
        A => S2418,
        B => S3911,
        Y => S4695
    );
NOR_1467: ENTITY WORK.NOR
    PORT MAP (
        A => S4557,
        B => S4695,
        Y => S4696
    );
NOR_1468: ENTITY WORK.NOR
    PORT MAP (
        A => S3912,
        B => S4558,
        Y => S4697
    );
NOR_1469: ENTITY WORK.NOR
    PORT MAP (
        A => S4696,
        B => S4697,
        Y => S4698
    );
NOR_1470: ENTITY WORK.NOR
    PORT MAP (
        A => S4560,
        B => S4698,
        Y => S4699
    );
NOT_369: ENTITY WORK.NOT
    PORT MAP (
        A => S4699,
        Y => S4700
    );
NOR_1471: ENTITY WORK.NOR
    PORT MAP (
        A => S2517,
        B => S4700,
        Y => S4701
    );
NAND_2970: ENTITY WORK.NAND
    PORT MAP (
        A => S2518,
        B => S4699,
        Y => S4702
    );
NOR_1472: ENTITY WORK.NOR
    PORT MAP (
        A => S4694,
        B => S4701,
        Y => S4703
    );
NAND_2971: ENTITY WORK.NAND
    PORT MAP (
        A => S4693,
        B => S4702,
        Y => S4704
    );
NAND_2972: ENTITY WORK.NAND
    PORT MAP (
        A => S2517,
        B => S4560,
        Y => S4705
    );
NAND_2973: ENTITY WORK.NAND
    PORT MAP (
        A => S3908,
        B => S4705,
        Y => S4706
    );
NOT_370: ENTITY WORK.NOT
    PORT MAP (
        A => S4706,
        Y => S4707
    );
NOR_1473: ENTITY WORK.NOR
    PORT MAP (
        A => S4703,
        B => S4706,
        Y => S4708
    );
NAND_2974: ENTITY WORK.NAND
    PORT MAP (
        A => S4704,
        B => S4707,
        Y => S4709
    );
NAND_2975: ENTITY WORK.NAND
    PORT MAP (
        A => S4582,
        B => S4689,
        Y => S4710
    );
NAND_2976: ENTITY WORK.NAND
    PORT MAP (
        A => S4692,
        B => S4710,
        Y => S4711
    );
NAND_2977: ENTITY WORK.NAND
    PORT MAP (
        A => S4708,
        B => S4711,
        Y => S4712
    );
NOT_371: ENTITY WORK.NOT
    PORT MAP (
        A => S4712,
        Y => S4713
    );
NOR_1474: ENTITY WORK.NOR
    PORT MAP (
        A => S4576,
        B => S4708,
        Y => S4714
    );
NOT_372: ENTITY WORK.NOT
    PORT MAP (
        A => S4714,
        Y => S4715
    );
NOR_1475: ENTITY WORK.NOR
    PORT MAP (
        A => S4713,
        B => S4714,
        Y => S4716
    );
NAND_2978: ENTITY WORK.NAND
    PORT MAP (
        A => S4712,
        B => S4715,
        Y => S4717
    );
NOR_1476: ENTITY WORK.NOR
    PORT MAP (
        A => S2517,
        B => S4717,
        Y => S4718
    );
NAND_2979: ENTITY WORK.NAND
    PORT MAP (
        A => S2518,
        B => S4716,
        Y => S4719
    );
NOR_1477: ENTITY WORK.NOR
    PORT MAP (
        A => S2518,
        B => S4716,
        Y => S4720
    );
NAND_2980: ENTITY WORK.NAND
    PORT MAP (
        A => S2517,
        B => S4717,
        Y => S4721
    );
NOR_1478: ENTITY WORK.NOR
    PORT MAP (
        A => S4718,
        B => S4720,
        Y => S4722
    );
NAND_2981: ENTITY WORK.NAND
    PORT MAP (
        A => S4719,
        B => S4721,
        Y => S4723
    );
NOR_1479: ENTITY WORK.NOR
    PORT MAP (
        A => S4593,
        B => S4594,
        Y => S4724
    );
NOR_1480: ENTITY WORK.NOR
    PORT MAP (
        A => S4686,
        B => S4724,
        Y => S4725
    );
NOT_373: ENTITY WORK.NOT
    PORT MAP (
        A => S4725,
        Y => S4726
    );
NAND_2982: ENTITY WORK.NAND
    PORT MAP (
        A => S4686,
        B => S4724,
        Y => S4727
    );
NAND_2983: ENTITY WORK.NAND
    PORT MAP (
        A => S4726,
        B => S4727,
        Y => S4728
    );
NAND_2984: ENTITY WORK.NAND
    PORT MAP (
        A => S4708,
        B => S4728,
        Y => S4729
    );
NOT_374: ENTITY WORK.NOT
    PORT MAP (
        A => S4729,
        Y => S4730
    );
NOR_1481: ENTITY WORK.NOR
    PORT MAP (
        A => S4591,
        B => S4708,
        Y => S4731
    );
NOT_375: ENTITY WORK.NOT
    PORT MAP (
        A => S4731,
        Y => S4732
    );
NOR_1482: ENTITY WORK.NOR
    PORT MAP (
        A => S4730,
        B => S4731,
        Y => S4733
    );
NAND_2985: ENTITY WORK.NAND
    PORT MAP (
        A => S4729,
        B => S4732,
        Y => S4734
    );
NOR_1483: ENTITY WORK.NOR
    PORT MAP (
        A => S2417,
        B => S4734,
        Y => S4735
    );
NAND_2986: ENTITY WORK.NAND
    PORT MAP (
        A => S2418,
        B => S4733,
        Y => S4736
    );
NOR_1484: ENTITY WORK.NOR
    PORT MAP (
        A => S2418,
        B => S4733,
        Y => S4737
    );
NAND_2987: ENTITY WORK.NAND
    PORT MAP (
        A => S2417,
        B => S4734,
        Y => S4738
    );
NAND_2988: ENTITY WORK.NAND
    PORT MAP (
        A => S4604,
        B => S4681,
        Y => S4739
    );
NAND_2989: ENTITY WORK.NAND
    PORT MAP (
        A => S4684,
        B => S4739,
        Y => S4740
    );
NAND_2990: ENTITY WORK.NAND
    PORT MAP (
        A => S4708,
        B => S4740,
        Y => S4741
    );
NOT_376: ENTITY WORK.NOT
    PORT MAP (
        A => S4741,
        Y => S4742
    );
NOR_1485: ENTITY WORK.NOR
    PORT MAP (
        A => S4599,
        B => S4708,
        Y => S4743
    );
NOT_377: ENTITY WORK.NOT
    PORT MAP (
        A => S4743,
        Y => S4744
    );
NOR_1486: ENTITY WORK.NOR
    PORT MAP (
        A => S4742,
        B => S4743,
        Y => S4745
    );
NAND_2991: ENTITY WORK.NAND
    PORT MAP (
        A => S4741,
        B => S4744,
        Y => S4746
    );
NOR_1487: ENTITY WORK.NOR
    PORT MAP (
        A => S2311,
        B => S4746,
        Y => S4747
    );
NAND_2992: ENTITY WORK.NAND
    PORT MAP (
        A => S2312,
        B => S4745,
        Y => S4748
    );
NOR_1488: ENTITY WORK.NOR
    PORT MAP (
        A => S2312,
        B => S4745,
        Y => S4749
    );
NAND_2993: ENTITY WORK.NAND
    PORT MAP (
        A => S2311,
        B => S4746,
        Y => S4750
    );
NOR_1489: ENTITY WORK.NOR
    PORT MAP (
        A => S4747,
        B => S4749,
        Y => S4751
    );
NAND_2994: ENTITY WORK.NAND
    PORT MAP (
        A => S4748,
        B => S4750,
        Y => S4752
    );
NAND_2995: ENTITY WORK.NAND
    PORT MAP (
        A => S4615,
        B => S4677,
        Y => S4753
    );
NAND_2996: ENTITY WORK.NAND
    PORT MAP (
        A => S4680,
        B => S4753,
        Y => S4754
    );
NAND_2997: ENTITY WORK.NAND
    PORT MAP (
        A => S4708,
        B => S4754,
        Y => S4755
    );
NOT_378: ENTITY WORK.NOT
    PORT MAP (
        A => S4755,
        Y => S4756
    );
NOR_1490: ENTITY WORK.NOR
    PORT MAP (
        A => S4610,
        B => S4708,
        Y => S4757
    );
NOT_379: ENTITY WORK.NOT
    PORT MAP (
        A => S4757,
        Y => S4758
    );
NOR_1491: ENTITY WORK.NOR
    PORT MAP (
        A => S4756,
        B => S4757,
        Y => S4759
    );
NAND_2998: ENTITY WORK.NAND
    PORT MAP (
        A => S4755,
        B => S4758,
        Y => S4760
    );
NOR_1492: ENTITY WORK.NOR
    PORT MAP (
        A => S2205,
        B => S4760,
        Y => S4761
    );
NAND_2999: ENTITY WORK.NAND
    PORT MAP (
        A => S2206,
        B => S4759,
        Y => S4762
    );
NOR_1493: ENTITY WORK.NOR
    PORT MAP (
        A => S2206,
        B => S4759,
        Y => S4763
    );
NAND_3000: ENTITY WORK.NAND
    PORT MAP (
        A => S2205,
        B => S4760,
        Y => S4764
    );
NOR_1494: ENTITY WORK.NOR
    PORT MAP (
        A => S4761,
        B => S4763,
        Y => S4765
    );
NAND_3001: ENTITY WORK.NAND
    PORT MAP (
        A => S4762,
        B => S4764,
        Y => S4766
    );
NAND_3002: ENTITY WORK.NAND
    PORT MAP (
        A => S4626,
        B => S4673,
        Y => S4767
    );
NAND_3003: ENTITY WORK.NAND
    PORT MAP (
        A => S4676,
        B => S4767,
        Y => S4768
    );
NAND_3004: ENTITY WORK.NAND
    PORT MAP (
        A => S4708,
        B => S4768,
        Y => S4769
    );
NOT_380: ENTITY WORK.NOT
    PORT MAP (
        A => S4769,
        Y => S4770
    );
NOR_1495: ENTITY WORK.NOR
    PORT MAP (
        A => S4621,
        B => S4708,
        Y => S4771
    );
NOT_381: ENTITY WORK.NOT
    PORT MAP (
        A => S4771,
        Y => S4772
    );
NOR_1496: ENTITY WORK.NOR
    PORT MAP (
        A => S4770,
        B => S4771,
        Y => S4773
    );
NAND_3005: ENTITY WORK.NAND
    PORT MAP (
        A => S4769,
        B => S4772,
        Y => S4774
    );
NOR_1497: ENTITY WORK.NOR
    PORT MAP (
        A => S2106,
        B => S4774,
        Y => S4775
    );
NAND_3006: ENTITY WORK.NAND
    PORT MAP (
        A => S2107,
        B => S4773,
        Y => S4776
    );
NOR_1498: ENTITY WORK.NOR
    PORT MAP (
        A => S2107,
        B => S4773,
        Y => S4777
    );
NAND_3007: ENTITY WORK.NAND
    PORT MAP (
        A => S2106,
        B => S4774,
        Y => S4778
    );
NOR_1499: ENTITY WORK.NOR
    PORT MAP (
        A => S4775,
        B => S4777,
        Y => S4779
    );
NAND_3008: ENTITY WORK.NAND
    PORT MAP (
        A => S4776,
        B => S4778,
        Y => S4780
    );
NAND_3009: ENTITY WORK.NAND
    PORT MAP (
        A => S4634,
        B => S4635,
        Y => S4781
    );
NOR_1500: ENTITY WORK.NOR
    PORT MAP (
        A => S4670,
        B => S4781,
        Y => S4782
    );
NAND_3010: ENTITY WORK.NAND
    PORT MAP (
        A => S4670,
        B => S4781,
        Y => S4783
    );
NOT_382: ENTITY WORK.NOT
    PORT MAP (
        A => S4783,
        Y => S4784
    );
NOR_1501: ENTITY WORK.NOR
    PORT MAP (
        A => S4782,
        B => S4784,
        Y => S4785
    );
NAND_3011: ENTITY WORK.NAND
    PORT MAP (
        A => S4708,
        B => S4785,
        Y => S4786
    );
NOT_383: ENTITY WORK.NOT
    PORT MAP (
        A => S4786,
        Y => S4787
    );
NOR_1502: ENTITY WORK.NOR
    PORT MAP (
        A => S4632,
        B => S4708,
        Y => S4788
    );
NOT_384: ENTITY WORK.NOT
    PORT MAP (
        A => S4788,
        Y => S4789
    );
NOR_1503: ENTITY WORK.NOR
    PORT MAP (
        A => S4787,
        B => S4788,
        Y => S4790
    );
NAND_3012: ENTITY WORK.NAND
    PORT MAP (
        A => S4786,
        B => S4789,
        Y => S4791
    );
NOR_1504: ENTITY WORK.NOR
    PORT MAP (
        A => S1597,
        B => S4791,
        Y => S4792
    );
NAND_3013: ENTITY WORK.NAND
    PORT MAP (
        A => S1598,
        B => S4790,
        Y => S4793
    );
NOR_1505: ENTITY WORK.NOR
    PORT MAP (
        A => S1598,
        B => S4790,
        Y => S4794
    );
NAND_3014: ENTITY WORK.NAND
    PORT MAP (
        A => S1597,
        B => S4791,
        Y => S4795
    );
NOR_1506: ENTITY WORK.NOR
    PORT MAP (
        A => S4792,
        B => S4794,
        Y => S4796
    );
NAND_3015: ENTITY WORK.NAND
    PORT MAP (
        A => S4793,
        B => S4795,
        Y => S4797
    );
NOR_1507: ENTITY WORK.NOR
    PORT MAP (
        A => S4640,
        B => S4708,
        Y => S4798
    );
NOT_385: ENTITY WORK.NOT
    PORT MAP (
        A => S4798,
        Y => S4799
    );
NAND_3016: ENTITY WORK.NAND
    PORT MAP (
        A => S4662,
        B => S4665,
        Y => S4800
    );
NAND_3017: ENTITY WORK.NAND
    PORT MAP (
        A => S4668,
        B => S4800,
        Y => S4801
    );
NAND_3018: ENTITY WORK.NAND
    PORT MAP (
        A => S4708,
        B => S4801,
        Y => S4802
    );
NOT_386: ENTITY WORK.NOT
    PORT MAP (
        A => S4802,
        Y => S4803
    );
NOR_1508: ENTITY WORK.NOR
    PORT MAP (
        A => S4798,
        B => S4803,
        Y => S4804
    );
NAND_3019: ENTITY WORK.NAND
    PORT MAP (
        A => S4799,
        B => S4802,
        Y => S4805
    );
NOR_1509: ENTITY WORK.NOR
    PORT MAP (
        A => S1952,
        B => S4805,
        Y => S4806
    );
NAND_3020: ENTITY WORK.NAND
    PORT MAP (
        A => S1953,
        B => S4804,
        Y => S4807
    );
NOR_1510: ENTITY WORK.NOR
    PORT MAP (
        A => S4654,
        B => S4658,
        Y => S4808
    );
NOR_1511: ENTITY WORK.NOR
    PORT MAP (
        A => S4660,
        B => S4808,
        Y => S4809
    );
NAND_3021: ENTITY WORK.NAND
    PORT MAP (
        A => S4708,
        B => S4809,
        Y => S4810
    );
NOT_387: ENTITY WORK.NOT
    PORT MAP (
        A => S4810,
        Y => S4811
    );
NOR_1512: ENTITY WORK.NOR
    PORT MAP (
        A => S4650,
        B => S4708,
        Y => S4812
    );
NOT_388: ENTITY WORK.NOT
    PORT MAP (
        A => S4812,
        Y => S4813
    );
NOR_1513: ENTITY WORK.NOR
    PORT MAP (
        A => S4811,
        B => S4812,
        Y => S4814
    );
NAND_3022: ENTITY WORK.NAND
    PORT MAP (
        A => S4810,
        B => S4813,
        Y => S4815
    );
NOR_1514: ENTITY WORK.NOR
    PORT MAP (
        A => S1848,
        B => S4814,
        Y => S4816
    );
NAND_3023: ENTITY WORK.NAND
    PORT MAP (
        A => S1849,
        B => S4815,
        Y => S4817
    );
NOR_1515: ENTITY WORK.NOR
    PORT MAP (
        A => S1849,
        B => S4815,
        Y => S4818
    );
NAND_3024: ENTITY WORK.NAND
    PORT MAP (
        A => S1848,
        B => S4814,
        Y => S4819
    );
NOR_1516: ENTITY WORK.NOR
    PORT MAP (
        A => S4816,
        B => S4818,
        Y => S4820
    );
NAND_3025: ENTITY WORK.NAND
    PORT MAP (
        A => S4817,
        B => S4819,
        Y => S4821
    );
NOR_1517: ENTITY WORK.NOR
    PORT MAP (
        A => S1516,
        B => S4709,
        Y => S4822
    );
NAND_3026: ENTITY WORK.NAND
    PORT MAP (
        A => S1515,
        B => S4708,
        Y => S4823
    );
NOR_1518: ENTITY WORK.NOR
    PORT MAP (
        A => S910,
        B => S4822,
        Y => S4824
    );
NAND_3027: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_6,
        B => S4823,
        Y => S4825
    );
NOR_1519: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_6,
        B => S4823,
        Y => S4826
    );
NAND_3028: ENTITY WORK.NAND
    PORT MAP (
        A => S910,
        B => S4822,
        Y => S4827
    );
NOR_1520: ENTITY WORK.NOR
    PORT MAP (
        A => S4824,
        B => S4826,
        Y => S4828
    );
NAND_3029: ENTITY WORK.NAND
    PORT MAP (
        A => S4825,
        B => S4827,
        Y => S4829
    );
NOR_1521: ENTITY WORK.NOR
    PORT MAP (
        A => S1745,
        B => S4828,
        Y => S4830
    );
NAND_3030: ENTITY WORK.NAND
    PORT MAP (
        A => S1746,
        B => S4829,
        Y => S4831
    );
NOR_1522: ENTITY WORK.NOR
    PORT MAP (
        A => S1746,
        B => S4829,
        Y => S4832
    );
NAND_3031: ENTITY WORK.NAND
    PORT MAP (
        A => S1745,
        B => S4828,
        Y => S4833
    );
NOR_1523: ENTITY WORK.NOR
    PORT MAP (
        A => S4830,
        B => S4832,
        Y => S4834
    );
NAND_3032: ENTITY WORK.NAND
    PORT MAP (
        A => S4831,
        B => S4833,
        Y => S4835
    );
NOR_1524: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_5,
        B => S1516,
        Y => S4836
    );
NAND_3033: ENTITY WORK.NAND
    PORT MAP (
        A => S963,
        B => S1515,
        Y => S4837
    );
NOR_1525: ENTITY WORK.NOR
    PORT MAP (
        A => S4835,
        B => S4836,
        Y => S4838
    );
NAND_3034: ENTITY WORK.NAND
    PORT MAP (
        A => S4834,
        B => S4837,
        Y => S4839
    );
NOR_1526: ENTITY WORK.NOR
    PORT MAP (
        A => S4830,
        B => S4838,
        Y => S4840
    );
NAND_3035: ENTITY WORK.NAND
    PORT MAP (
        A => S4831,
        B => S4839,
        Y => S4841
    );
NOR_1527: ENTITY WORK.NOR
    PORT MAP (
        A => S4821,
        B => S4840,
        Y => S4842
    );
NAND_3036: ENTITY WORK.NAND
    PORT MAP (
        A => S4820,
        B => S4841,
        Y => S4843
    );
NOR_1528: ENTITY WORK.NOR
    PORT MAP (
        A => S4816,
        B => S4842,
        Y => S4844
    );
NAND_3037: ENTITY WORK.NAND
    PORT MAP (
        A => S4817,
        B => S4843,
        Y => S4845
    );
NOR_1529: ENTITY WORK.NOR
    PORT MAP (
        A => S1953,
        B => S4804,
        Y => S4846
    );
NAND_3038: ENTITY WORK.NAND
    PORT MAP (
        A => S1952,
        B => S4805,
        Y => S4847
    );
NOR_1530: ENTITY WORK.NOR
    PORT MAP (
        A => S4806,
        B => S4846,
        Y => S4848
    );
NAND_3039: ENTITY WORK.NAND
    PORT MAP (
        A => S4807,
        B => S4847,
        Y => S4849
    );
NOR_1531: ENTITY WORK.NOR
    PORT MAP (
        A => S4844,
        B => S4849,
        Y => S4850
    );
NAND_3040: ENTITY WORK.NAND
    PORT MAP (
        A => S4845,
        B => S4848,
        Y => S4851
    );
NOR_1532: ENTITY WORK.NOR
    PORT MAP (
        A => S4806,
        B => S4850,
        Y => S4852
    );
NAND_3041: ENTITY WORK.NAND
    PORT MAP (
        A => S4807,
        B => S4851,
        Y => S4853
    );
NOR_1533: ENTITY WORK.NOR
    PORT MAP (
        A => S4797,
        B => S4852,
        Y => S4854
    );
NAND_3042: ENTITY WORK.NAND
    PORT MAP (
        A => S4796,
        B => S4853,
        Y => S4855
    );
NOR_1534: ENTITY WORK.NOR
    PORT MAP (
        A => S4792,
        B => S4854,
        Y => S4856
    );
NAND_3043: ENTITY WORK.NAND
    PORT MAP (
        A => S4793,
        B => S4855,
        Y => S4857
    );
NOR_1535: ENTITY WORK.NOR
    PORT MAP (
        A => S4780,
        B => S4856,
        Y => S4858
    );
NAND_3044: ENTITY WORK.NAND
    PORT MAP (
        A => S4779,
        B => S4857,
        Y => S4859
    );
NOR_1536: ENTITY WORK.NOR
    PORT MAP (
        A => S4775,
        B => S4858,
        Y => S4860
    );
NAND_3045: ENTITY WORK.NAND
    PORT MAP (
        A => S4776,
        B => S4859,
        Y => S4861
    );
NOR_1537: ENTITY WORK.NOR
    PORT MAP (
        A => S4766,
        B => S4860,
        Y => S4862
    );
NAND_3046: ENTITY WORK.NAND
    PORT MAP (
        A => S4765,
        B => S4861,
        Y => S4863
    );
NOR_1538: ENTITY WORK.NOR
    PORT MAP (
        A => S4761,
        B => S4862,
        Y => S4864
    );
NAND_3047: ENTITY WORK.NAND
    PORT MAP (
        A => S4762,
        B => S4863,
        Y => S4865
    );
NOR_1539: ENTITY WORK.NOR
    PORT MAP (
        A => S4752,
        B => S4864,
        Y => S4866
    );
NAND_3048: ENTITY WORK.NAND
    PORT MAP (
        A => S4751,
        B => S4865,
        Y => S4867
    );
NOR_1540: ENTITY WORK.NOR
    PORT MAP (
        A => S4747,
        B => S4866,
        Y => S4868
    );
NAND_3049: ENTITY WORK.NAND
    PORT MAP (
        A => S4748,
        B => S4867,
        Y => S4869
    );
NOR_1541: ENTITY WORK.NOR
    PORT MAP (
        A => S4737,
        B => S4868,
        Y => S4870
    );
NAND_3050: ENTITY WORK.NAND
    PORT MAP (
        A => S4738,
        B => S4869,
        Y => S4871
    );
NOR_1542: ENTITY WORK.NOR
    PORT MAP (
        A => S4735,
        B => S4870,
        Y => S4872
    );
NAND_3051: ENTITY WORK.NAND
    PORT MAP (
        A => S4736,
        B => S4871,
        Y => S4873
    );
NOR_1543: ENTITY WORK.NOR
    PORT MAP (
        A => S4723,
        B => S4872,
        Y => S4874
    );
NAND_3052: ENTITY WORK.NAND
    PORT MAP (
        A => S4722,
        B => S4873,
        Y => S4875
    );
NAND_3053: ENTITY WORK.NAND
    PORT MAP (
        A => S2517,
        B => S3908,
        Y => S4876
    );
NOT_389: ENTITY WORK.NOT
    PORT MAP (
        A => S4876,
        Y => S4877
    );
NOR_1544: ENTITY WORK.NOR
    PORT MAP (
        A => S4693,
        B => S4877,
        Y => S4878
    );
NOR_1545: ENTITY WORK.NOR
    PORT MAP (
        A => S3910,
        B => S4694,
        Y => S4879
    );
NOR_1546: ENTITY WORK.NOR
    PORT MAP (
        A => S4878,
        B => S4879,
        Y => S4880
    );
NOR_1547: ENTITY WORK.NOR
    PORT MAP (
        A => S4700,
        B => S4880,
        Y => S4881
    );
NOT_390: ENTITY WORK.NOT
    PORT MAP (
        A => S4881,
        Y => S4882
    );
NOR_1548: ENTITY WORK.NOR
    PORT MAP (
        A => S2617,
        B => S4882,
        Y => S4883
    );
NAND_3054: ENTITY WORK.NAND
    PORT MAP (
        A => S2618,
        B => S4881,
        Y => S4884
    );
NOR_1549: ENTITY WORK.NOR
    PORT MAP (
        A => S4718,
        B => S4883,
        Y => S4885
    );
NAND_3055: ENTITY WORK.NAND
    PORT MAP (
        A => S4719,
        B => S4884,
        Y => S4886
    );
NOR_1550: ENTITY WORK.NOR
    PORT MAP (
        A => S4874,
        B => S4886,
        Y => S4887
    );
NAND_3056: ENTITY WORK.NAND
    PORT MAP (
        A => S4875,
        B => S4885,
        Y => S4888
    );
NOR_1551: ENTITY WORK.NOR
    PORT MAP (
        A => S2618,
        B => S4699,
        Y => S4889
    );
NAND_3057: ENTITY WORK.NAND
    PORT MAP (
        A => S2617,
        B => S4700,
        Y => S4890
    );
NOR_1552: ENTITY WORK.NOR
    PORT MAP (
        A => S3907,
        B => S4889,
        Y => S4891
    );
NAND_3058: ENTITY WORK.NAND
    PORT MAP (
        A => S3906,
        B => S4890,
        Y => S4892
    );
NOR_1553: ENTITY WORK.NOR
    PORT MAP (
        A => S4883,
        B => S4889,
        Y => S4893
    );
NAND_3059: ENTITY WORK.NAND
    PORT MAP (
        A => S4884,
        B => S4890,
        Y => S4894
    );
NOR_1554: ENTITY WORK.NOR
    PORT MAP (
        A => S4887,
        B => S4892,
        Y => S4895
    );
NAND_3060: ENTITY WORK.NAND
    PORT MAP (
        A => S4888,
        B => S4891,
        Y => S4896
    );
NOR_1555: ENTITY WORK.NOR
    PORT MAP (
        A => S4722,
        B => S4873,
        Y => S4897
    );
NAND_3061: ENTITY WORK.NAND
    PORT MAP (
        A => S4723,
        B => S4872,
        Y => S4898
    );
NOR_1556: ENTITY WORK.NOR
    PORT MAP (
        A => S4874,
        B => S4897,
        Y => S4899
    );
NAND_3062: ENTITY WORK.NAND
    PORT MAP (
        A => S4875,
        B => S4898,
        Y => S4900
    );
NOR_1557: ENTITY WORK.NOR
    PORT MAP (
        A => S4896,
        B => S4899,
        Y => S4901
    );
NAND_3063: ENTITY WORK.NAND
    PORT MAP (
        A => S4895,
        B => S4900,
        Y => S4902
    );
NOR_1558: ENTITY WORK.NOR
    PORT MAP (
        A => S4716,
        B => S4895,
        Y => S4903
    );
NAND_3064: ENTITY WORK.NAND
    PORT MAP (
        A => S4717,
        B => S4896,
        Y => S4904
    );
NOR_1559: ENTITY WORK.NOR
    PORT MAP (
        A => S4901,
        B => S4903,
        Y => S4905
    );
NAND_3065: ENTITY WORK.NAND
    PORT MAP (
        A => S4902,
        B => S4904,
        Y => S4906
    );
NOR_1560: ENTITY WORK.NOR
    PORT MAP (
        A => S2617,
        B => S4906,
        Y => S4907
    );
NAND_3066: ENTITY WORK.NAND
    PORT MAP (
        A => S2618,
        B => S4905,
        Y => S4908
    );
NOR_1561: ENTITY WORK.NOR
    PORT MAP (
        A => S2618,
        B => S4905,
        Y => S4909
    );
NAND_3067: ENTITY WORK.NAND
    PORT MAP (
        A => S2617,
        B => S4906,
        Y => S4910
    );
NOR_1562: ENTITY WORK.NOR
    PORT MAP (
        A => S4907,
        B => S4909,
        Y => S4911
    );
NAND_3068: ENTITY WORK.NAND
    PORT MAP (
        A => S4908,
        B => S4910,
        Y => S4912
    );
NOR_1563: ENTITY WORK.NOR
    PORT MAP (
        A => S4735,
        B => S4737,
        Y => S4913
    );
NAND_3069: ENTITY WORK.NAND
    PORT MAP (
        A => S4736,
        B => S4738,
        Y => S4914
    );
NOR_1564: ENTITY WORK.NOR
    PORT MAP (
        A => S4869,
        B => S4913,
        Y => S4915
    );
NAND_3070: ENTITY WORK.NAND
    PORT MAP (
        A => S4868,
        B => S4914,
        Y => S4916
    );
NOR_1565: ENTITY WORK.NOR
    PORT MAP (
        A => S4868,
        B => S4914,
        Y => S4917
    );
NAND_3071: ENTITY WORK.NAND
    PORT MAP (
        A => S4869,
        B => S4913,
        Y => S4918
    );
NOR_1566: ENTITY WORK.NOR
    PORT MAP (
        A => S4915,
        B => S4917,
        Y => S4919
    );
NAND_3072: ENTITY WORK.NAND
    PORT MAP (
        A => S4916,
        B => S4918,
        Y => S4920
    );
NOR_1567: ENTITY WORK.NOR
    PORT MAP (
        A => S4896,
        B => S4919,
        Y => S4921
    );
NAND_3073: ENTITY WORK.NAND
    PORT MAP (
        A => S4895,
        B => S4920,
        Y => S4922
    );
NOR_1568: ENTITY WORK.NOR
    PORT MAP (
        A => S4733,
        B => S4895,
        Y => S4923
    );
NAND_3074: ENTITY WORK.NAND
    PORT MAP (
        A => S4734,
        B => S4896,
        Y => S4924
    );
NOR_1569: ENTITY WORK.NOR
    PORT MAP (
        A => S4921,
        B => S4923,
        Y => S4925
    );
NAND_3075: ENTITY WORK.NAND
    PORT MAP (
        A => S4922,
        B => S4924,
        Y => S4926
    );
NOR_1570: ENTITY WORK.NOR
    PORT MAP (
        A => S2518,
        B => S4925,
        Y => S4927
    );
NAND_3076: ENTITY WORK.NAND
    PORT MAP (
        A => S2517,
        B => S4926,
        Y => S4928
    );
NOR_1571: ENTITY WORK.NOR
    PORT MAP (
        A => S2517,
        B => S4926,
        Y => S4929
    );
NAND_3077: ENTITY WORK.NAND
    PORT MAP (
        A => S2518,
        B => S4925,
        Y => S4930
    );
NOR_1572: ENTITY WORK.NOR
    PORT MAP (
        A => S4751,
        B => S4865,
        Y => S4931
    );
NAND_3078: ENTITY WORK.NAND
    PORT MAP (
        A => S4752,
        B => S4864,
        Y => S4932
    );
NOR_1573: ENTITY WORK.NOR
    PORT MAP (
        A => S4866,
        B => S4931,
        Y => S4933
    );
NAND_3079: ENTITY WORK.NAND
    PORT MAP (
        A => S4867,
        B => S4932,
        Y => S4934
    );
NOR_1574: ENTITY WORK.NOR
    PORT MAP (
        A => S4896,
        B => S4933,
        Y => S4935
    );
NAND_3080: ENTITY WORK.NAND
    PORT MAP (
        A => S4895,
        B => S4934,
        Y => S4936
    );
NOR_1575: ENTITY WORK.NOR
    PORT MAP (
        A => S4745,
        B => S4895,
        Y => S4937
    );
NAND_3081: ENTITY WORK.NAND
    PORT MAP (
        A => S4746,
        B => S4896,
        Y => S4938
    );
NOR_1576: ENTITY WORK.NOR
    PORT MAP (
        A => S4935,
        B => S4937,
        Y => S4939
    );
NAND_3082: ENTITY WORK.NAND
    PORT MAP (
        A => S4936,
        B => S4938,
        Y => S4940
    );
NOR_1577: ENTITY WORK.NOR
    PORT MAP (
        A => S2417,
        B => S4940,
        Y => S4941
    );
NAND_3083: ENTITY WORK.NAND
    PORT MAP (
        A => S2418,
        B => S4939,
        Y => S4942
    );
NOR_1578: ENTITY WORK.NOR
    PORT MAP (
        A => S2418,
        B => S4939,
        Y => S4943
    );
NAND_3084: ENTITY WORK.NAND
    PORT MAP (
        A => S2417,
        B => S4940,
        Y => S4944
    );
NOR_1579: ENTITY WORK.NOR
    PORT MAP (
        A => S4941,
        B => S4943,
        Y => S4945
    );
NAND_3085: ENTITY WORK.NAND
    PORT MAP (
        A => S4942,
        B => S4944,
        Y => S4946
    );
NOR_1580: ENTITY WORK.NOR
    PORT MAP (
        A => S4765,
        B => S4861,
        Y => S4947
    );
NAND_3086: ENTITY WORK.NAND
    PORT MAP (
        A => S4766,
        B => S4860,
        Y => S4948
    );
NOR_1581: ENTITY WORK.NOR
    PORT MAP (
        A => S4862,
        B => S4947,
        Y => S4949
    );
NAND_3087: ENTITY WORK.NAND
    PORT MAP (
        A => S4863,
        B => S4948,
        Y => S4950
    );
NOR_1582: ENTITY WORK.NOR
    PORT MAP (
        A => S4896,
        B => S4949,
        Y => S4951
    );
NAND_3088: ENTITY WORK.NAND
    PORT MAP (
        A => S4895,
        B => S4950,
        Y => S4952
    );
NOR_1583: ENTITY WORK.NOR
    PORT MAP (
        A => S4759,
        B => S4895,
        Y => S4953
    );
NAND_3089: ENTITY WORK.NAND
    PORT MAP (
        A => S4760,
        B => S4896,
        Y => S4954
    );
NOR_1584: ENTITY WORK.NOR
    PORT MAP (
        A => S4951,
        B => S4953,
        Y => S4955
    );
NAND_3090: ENTITY WORK.NAND
    PORT MAP (
        A => S4952,
        B => S4954,
        Y => S4956
    );
NOR_1585: ENTITY WORK.NOR
    PORT MAP (
        A => S2311,
        B => S4956,
        Y => S4957
    );
NAND_3091: ENTITY WORK.NAND
    PORT MAP (
        A => S2312,
        B => S4955,
        Y => S4958
    );
NOR_1586: ENTITY WORK.NOR
    PORT MAP (
        A => S2312,
        B => S4955,
        Y => S4959
    );
NAND_3092: ENTITY WORK.NAND
    PORT MAP (
        A => S2311,
        B => S4956,
        Y => S4960
    );
NOR_1587: ENTITY WORK.NOR
    PORT MAP (
        A => S4773,
        B => S4895,
        Y => S4961
    );
NAND_3093: ENTITY WORK.NAND
    PORT MAP (
        A => S4774,
        B => S4896,
        Y => S4962
    );
NOR_1588: ENTITY WORK.NOR
    PORT MAP (
        A => S4779,
        B => S4857,
        Y => S4963
    );
NAND_3094: ENTITY WORK.NAND
    PORT MAP (
        A => S4780,
        B => S4856,
        Y => S4964
    );
NOR_1589: ENTITY WORK.NOR
    PORT MAP (
        A => S4858,
        B => S4963,
        Y => S4965
    );
NAND_3095: ENTITY WORK.NAND
    PORT MAP (
        A => S4859,
        B => S4964,
        Y => S4966
    );
NOR_1590: ENTITY WORK.NOR
    PORT MAP (
        A => S4896,
        B => S4965,
        Y => S4967
    );
NAND_3096: ENTITY WORK.NAND
    PORT MAP (
        A => S4895,
        B => S4966,
        Y => S4968
    );
NOR_1591: ENTITY WORK.NOR
    PORT MAP (
        A => S4961,
        B => S4967,
        Y => S4969
    );
NAND_3097: ENTITY WORK.NAND
    PORT MAP (
        A => S4962,
        B => S4968,
        Y => S4970
    );
NOR_1592: ENTITY WORK.NOR
    PORT MAP (
        A => S2205,
        B => S4970,
        Y => S4971
    );
NAND_3098: ENTITY WORK.NAND
    PORT MAP (
        A => S2206,
        B => S4969,
        Y => S4972
    );
NOR_1593: ENTITY WORK.NOR
    PORT MAP (
        A => S2206,
        B => S4969,
        Y => S4973
    );
NAND_3099: ENTITY WORK.NAND
    PORT MAP (
        A => S2205,
        B => S4970,
        Y => S4974
    );
NOR_1594: ENTITY WORK.NOR
    PORT MAP (
        A => S4971,
        B => S4973,
        Y => S4975
    );
NAND_3100: ENTITY WORK.NAND
    PORT MAP (
        A => S4972,
        B => S4974,
        Y => S4976
    );
NOR_1595: ENTITY WORK.NOR
    PORT MAP (
        A => S4796,
        B => S4853,
        Y => S4977
    );
NAND_3101: ENTITY WORK.NAND
    PORT MAP (
        A => S4797,
        B => S4852,
        Y => S4978
    );
NOR_1596: ENTITY WORK.NOR
    PORT MAP (
        A => S4854,
        B => S4977,
        Y => S4979
    );
NAND_3102: ENTITY WORK.NAND
    PORT MAP (
        A => S4855,
        B => S4978,
        Y => S4980
    );
NOR_1597: ENTITY WORK.NOR
    PORT MAP (
        A => S4896,
        B => S4979,
        Y => S4981
    );
NAND_3103: ENTITY WORK.NAND
    PORT MAP (
        A => S4895,
        B => S4980,
        Y => S4982
    );
NOR_1598: ENTITY WORK.NOR
    PORT MAP (
        A => S4790,
        B => S4895,
        Y => S4983
    );
NAND_3104: ENTITY WORK.NAND
    PORT MAP (
        A => S4791,
        B => S4896,
        Y => S4984
    );
NOR_1599: ENTITY WORK.NOR
    PORT MAP (
        A => S4981,
        B => S4983,
        Y => S4985
    );
NAND_3105: ENTITY WORK.NAND
    PORT MAP (
        A => S4982,
        B => S4984,
        Y => S4986
    );
NOR_1600: ENTITY WORK.NOR
    PORT MAP (
        A => S2106,
        B => S4986,
        Y => S4987
    );
NAND_3106: ENTITY WORK.NAND
    PORT MAP (
        A => S2107,
        B => S4985,
        Y => S4988
    );
NOR_1601: ENTITY WORK.NOR
    PORT MAP (
        A => S2107,
        B => S4985,
        Y => S4989
    );
NAND_3107: ENTITY WORK.NAND
    PORT MAP (
        A => S2106,
        B => S4986,
        Y => S4990
    );
NOR_1602: ENTITY WORK.NOR
    PORT MAP (
        A => S4804,
        B => S4895,
        Y => S4991
    );
NAND_3108: ENTITY WORK.NAND
    PORT MAP (
        A => S4805,
        B => S4896,
        Y => S4992
    );
NOR_1603: ENTITY WORK.NOR
    PORT MAP (
        A => S4845,
        B => S4848,
        Y => S4993
    );
NAND_3109: ENTITY WORK.NAND
    PORT MAP (
        A => S4844,
        B => S4849,
        Y => S4994
    );
NOR_1604: ENTITY WORK.NOR
    PORT MAP (
        A => S4850,
        B => S4993,
        Y => S4995
    );
NAND_3110: ENTITY WORK.NAND
    PORT MAP (
        A => S4851,
        B => S4994,
        Y => S4996
    );
NOR_1605: ENTITY WORK.NOR
    PORT MAP (
        A => S4896,
        B => S4995,
        Y => S4997
    );
NAND_3111: ENTITY WORK.NAND
    PORT MAP (
        A => S4895,
        B => S4996,
        Y => S4998
    );
NOR_1606: ENTITY WORK.NOR
    PORT MAP (
        A => S4991,
        B => S4997,
        Y => S4999
    );
NAND_3112: ENTITY WORK.NAND
    PORT MAP (
        A => S4992,
        B => S4998,
        Y => S5000
    );
NOR_1607: ENTITY WORK.NOR
    PORT MAP (
        A => S1597,
        B => S5000,
        Y => S5001
    );
NAND_3113: ENTITY WORK.NAND
    PORT MAP (
        A => S1598,
        B => S4999,
        Y => S5002
    );
NOR_1608: ENTITY WORK.NOR
    PORT MAP (
        A => S4815,
        B => S4895,
        Y => S5003
    );
NAND_3114: ENTITY WORK.NAND
    PORT MAP (
        A => S4814,
        B => S4896,
        Y => S5004
    );
NOR_1609: ENTITY WORK.NOR
    PORT MAP (
        A => S4820,
        B => S4841,
        Y => S5005
    );
NAND_3115: ENTITY WORK.NAND
    PORT MAP (
        A => S4821,
        B => S4840,
        Y => S5006
    );
NOR_1610: ENTITY WORK.NOR
    PORT MAP (
        A => S4842,
        B => S5005,
        Y => S5007
    );
NAND_3116: ENTITY WORK.NAND
    PORT MAP (
        A => S4843,
        B => S5006,
        Y => S5008
    );
NOR_1611: ENTITY WORK.NOR
    PORT MAP (
        A => S4896,
        B => S5007,
        Y => S5009
    );
NAND_3117: ENTITY WORK.NAND
    PORT MAP (
        A => S4895,
        B => S5008,
        Y => S5010
    );
NOR_1612: ENTITY WORK.NOR
    PORT MAP (
        A => S5003,
        B => S5009,
        Y => S5011
    );
NAND_3118: ENTITY WORK.NAND
    PORT MAP (
        A => S5004,
        B => S5010,
        Y => S5012
    );
NOR_1613: ENTITY WORK.NOR
    PORT MAP (
        A => S1952,
        B => S5012,
        Y => S5013
    );
NAND_3119: ENTITY WORK.NAND
    PORT MAP (
        A => S1953,
        B => S5011,
        Y => S5014
    );
NOR_1614: ENTITY WORK.NOR
    PORT MAP (
        A => S1953,
        B => S5011,
        Y => S5015
    );
NAND_3120: ENTITY WORK.NAND
    PORT MAP (
        A => S1952,
        B => S5012,
        Y => S5016
    );
NOR_1615: ENTITY WORK.NOR
    PORT MAP (
        A => S5013,
        B => S5015,
        Y => S5017
    );
NAND_3121: ENTITY WORK.NAND
    PORT MAP (
        A => S5014,
        B => S5016,
        Y => S5018
    );
NOR_1616: ENTITY WORK.NOR
    PORT MAP (
        A => S4834,
        B => S4837,
        Y => S5019
    );
NAND_3122: ENTITY WORK.NAND
    PORT MAP (
        A => S4835,
        B => S4836,
        Y => S5020
    );
NOR_1617: ENTITY WORK.NOR
    PORT MAP (
        A => S4838,
        B => S5019,
        Y => S5021
    );
NAND_3123: ENTITY WORK.NAND
    PORT MAP (
        A => S4839,
        B => S5020,
        Y => S5022
    );
NOR_1618: ENTITY WORK.NOR
    PORT MAP (
        A => S4896,
        B => S5021,
        Y => S5023
    );
NAND_3124: ENTITY WORK.NAND
    PORT MAP (
        A => S4895,
        B => S5022,
        Y => S5024
    );
NOR_1619: ENTITY WORK.NOR
    PORT MAP (
        A => S4829,
        B => S4895,
        Y => S5025
    );
NAND_3125: ENTITY WORK.NAND
    PORT MAP (
        A => S4828,
        B => S4896,
        Y => S5026
    );
NOR_1620: ENTITY WORK.NOR
    PORT MAP (
        A => S5023,
        B => S5025,
        Y => S5027
    );
NAND_3126: ENTITY WORK.NAND
    PORT MAP (
        A => S5024,
        B => S5026,
        Y => S5028
    );
NOR_1621: ENTITY WORK.NOR
    PORT MAP (
        A => S1848,
        B => S5028,
        Y => S5029
    );
NAND_3127: ENTITY WORK.NAND
    PORT MAP (
        A => S1849,
        B => S5027,
        Y => S5030
    );
NOR_1622: ENTITY WORK.NOR
    PORT MAP (
        A => S1849,
        B => S5027,
        Y => S5031
    );
NAND_3128: ENTITY WORK.NAND
    PORT MAP (
        A => S1848,
        B => S5028,
        Y => S5032
    );
NOR_1623: ENTITY WORK.NOR
    PORT MAP (
        A => S5029,
        B => S5031,
        Y => S5033
    );
NAND_3129: ENTITY WORK.NAND
    PORT MAP (
        A => S5030,
        B => S5032,
        Y => S5034
    );
NOR_1624: ENTITY WORK.NOR
    PORT MAP (
        A => S1516,
        B => S4896,
        Y => S5035
    );
NAND_3130: ENTITY WORK.NAND
    PORT MAP (
        A => S1515,
        B => S4895,
        Y => S5036
    );
NOR_1625: ENTITY WORK.NOR
    PORT MAP (
        A => S963,
        B => S5035,
        Y => S5037
    );
NAND_3131: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_5,
        B => S5036,
        Y => S5038
    );
NOR_1626: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_5,
        B => S5036,
        Y => S5039
    );
NAND_3132: ENTITY WORK.NAND
    PORT MAP (
        A => S963,
        B => S5035,
        Y => S5040
    );
NOR_1627: ENTITY WORK.NOR
    PORT MAP (
        A => S5037,
        B => S5039,
        Y => S5041
    );
NAND_3133: ENTITY WORK.NAND
    PORT MAP (
        A => S5038,
        B => S5040,
        Y => S5042
    );
NOR_1628: ENTITY WORK.NOR
    PORT MAP (
        A => S1745,
        B => S5041,
        Y => S5043
    );
NAND_3134: ENTITY WORK.NAND
    PORT MAP (
        A => S1746,
        B => S5042,
        Y => S5044
    );
NOR_1629: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_4,
        B => S1516,
        Y => S5045
    );
NAND_3135: ENTITY WORK.NAND
    PORT MAP (
        A => S1013,
        B => S1515,
        Y => S5046
    );
NOR_1630: ENTITY WORK.NOR
    PORT MAP (
        A => S1746,
        B => S5042,
        Y => S5047
    );
NAND_3136: ENTITY WORK.NAND
    PORT MAP (
        A => S1745,
        B => S5041,
        Y => S5048
    );
NOR_1631: ENTITY WORK.NOR
    PORT MAP (
        A => S5043,
        B => S5047,
        Y => S5049
    );
NAND_3137: ENTITY WORK.NAND
    PORT MAP (
        A => S5044,
        B => S5048,
        Y => S5050
    );
NOR_1632: ENTITY WORK.NOR
    PORT MAP (
        A => S5045,
        B => S5050,
        Y => S5051
    );
NAND_3138: ENTITY WORK.NAND
    PORT MAP (
        A => S5046,
        B => S5049,
        Y => S5052
    );
NOR_1633: ENTITY WORK.NOR
    PORT MAP (
        A => S5043,
        B => S5051,
        Y => S5053
    );
NAND_3139: ENTITY WORK.NAND
    PORT MAP (
        A => S5044,
        B => S5052,
        Y => S5054
    );
NOR_1634: ENTITY WORK.NOR
    PORT MAP (
        A => S5034,
        B => S5053,
        Y => S5055
    );
NAND_3140: ENTITY WORK.NAND
    PORT MAP (
        A => S5033,
        B => S5054,
        Y => S5056
    );
NOR_1635: ENTITY WORK.NOR
    PORT MAP (
        A => S5029,
        B => S5055,
        Y => S5057
    );
NAND_3141: ENTITY WORK.NAND
    PORT MAP (
        A => S5030,
        B => S5056,
        Y => S5058
    );
NOR_1636: ENTITY WORK.NOR
    PORT MAP (
        A => S5018,
        B => S5057,
        Y => S5059
    );
NAND_3142: ENTITY WORK.NAND
    PORT MAP (
        A => S5017,
        B => S5058,
        Y => S5060
    );
NOR_1637: ENTITY WORK.NOR
    PORT MAP (
        A => S5013,
        B => S5059,
        Y => S5061
    );
NAND_3143: ENTITY WORK.NAND
    PORT MAP (
        A => S5014,
        B => S5060,
        Y => S5062
    );
NOR_1638: ENTITY WORK.NOR
    PORT MAP (
        A => S1598,
        B => S4999,
        Y => S5063
    );
NAND_3144: ENTITY WORK.NAND
    PORT MAP (
        A => S1597,
        B => S5000,
        Y => S5064
    );
NOR_1639: ENTITY WORK.NOR
    PORT MAP (
        A => S5001,
        B => S5063,
        Y => S5065
    );
NAND_3145: ENTITY WORK.NAND
    PORT MAP (
        A => S5002,
        B => S5064,
        Y => S5066
    );
NOR_1640: ENTITY WORK.NOR
    PORT MAP (
        A => S5061,
        B => S5066,
        Y => S5067
    );
NAND_3146: ENTITY WORK.NAND
    PORT MAP (
        A => S5062,
        B => S5065,
        Y => S5068
    );
NOR_1641: ENTITY WORK.NOR
    PORT MAP (
        A => S5001,
        B => S5067,
        Y => S5069
    );
NAND_3147: ENTITY WORK.NAND
    PORT MAP (
        A => S5002,
        B => S5068,
        Y => S5070
    );
NOR_1642: ENTITY WORK.NOR
    PORT MAP (
        A => S4989,
        B => S5069,
        Y => S5071
    );
NAND_3148: ENTITY WORK.NAND
    PORT MAP (
        A => S4990,
        B => S5070,
        Y => S5072
    );
NOR_1643: ENTITY WORK.NOR
    PORT MAP (
        A => S4987,
        B => S5071,
        Y => S5073
    );
NAND_3149: ENTITY WORK.NAND
    PORT MAP (
        A => S4988,
        B => S5072,
        Y => S5074
    );
NOR_1644: ENTITY WORK.NOR
    PORT MAP (
        A => S4976,
        B => S5073,
        Y => S5075
    );
NAND_3150: ENTITY WORK.NAND
    PORT MAP (
        A => S4975,
        B => S5074,
        Y => S5076
    );
NOR_1645: ENTITY WORK.NOR
    PORT MAP (
        A => S4971,
        B => S5075,
        Y => S5077
    );
NAND_3151: ENTITY WORK.NAND
    PORT MAP (
        A => S4972,
        B => S5076,
        Y => S5078
    );
NOR_1646: ENTITY WORK.NOR
    PORT MAP (
        A => S4959,
        B => S5077,
        Y => S5079
    );
NAND_3152: ENTITY WORK.NAND
    PORT MAP (
        A => S4960,
        B => S5078,
        Y => S5080
    );
NOR_1647: ENTITY WORK.NOR
    PORT MAP (
        A => S4957,
        B => S5079,
        Y => S5081
    );
NAND_3153: ENTITY WORK.NAND
    PORT MAP (
        A => S4958,
        B => S5080,
        Y => S5082
    );
NOR_1648: ENTITY WORK.NOR
    PORT MAP (
        A => S4946,
        B => S5081,
        Y => S5083
    );
NAND_3154: ENTITY WORK.NAND
    PORT MAP (
        A => S4945,
        B => S5082,
        Y => S5084
    );
NOR_1649: ENTITY WORK.NOR
    PORT MAP (
        A => S4941,
        B => S5083,
        Y => S5085
    );
NAND_3155: ENTITY WORK.NAND
    PORT MAP (
        A => S4942,
        B => S5084,
        Y => S5086
    );
NOR_1650: ENTITY WORK.NOR
    PORT MAP (
        A => S4929,
        B => S5086,
        Y => S5087
    );
NAND_3156: ENTITY WORK.NAND
    PORT MAP (
        A => S4930,
        B => S5085,
        Y => S5088
    );
NOR_1651: ENTITY WORK.NOR
    PORT MAP (
        A => S4927,
        B => S5087,
        Y => S5089
    );
NAND_3157: ENTITY WORK.NAND
    PORT MAP (
        A => S4928,
        B => S5088,
        Y => S5090
    );
NOR_1652: ENTITY WORK.NOR
    PORT MAP (
        A => S4912,
        B => S5090,
        Y => S5091
    );
NAND_3158: ENTITY WORK.NAND
    PORT MAP (
        A => S4911,
        B => S5089,
        Y => S5092
    );
NOR_1653: ENTITY WORK.NOR
    PORT MAP (
        A => S4881,
        B => S4895,
        Y => S5093
    );
NOR_1654: ENTITY WORK.NOR
    PORT MAP (
        A => S4718,
        B => S4874,
        Y => S5094
    );
NAND_3159: ENTITY WORK.NAND
    PORT MAP (
        A => S4719,
        B => S4875,
        Y => S5095
    );
NOR_1655: ENTITY WORK.NOR
    PORT MAP (
        A => S4894,
        B => S5094,
        Y => S5096
    );
NOR_1656: ENTITY WORK.NOR
    PORT MAP (
        A => S4893,
        B => S5095,
        Y => S5097
    );
NOR_1657: ENTITY WORK.NOR
    PORT MAP (
        A => S5096,
        B => S5097,
        Y => S5098
    );
NOR_1658: ENTITY WORK.NOR
    PORT MAP (
        A => S4896,
        B => S5098,
        Y => S5099
    );
NOR_1659: ENTITY WORK.NOR
    PORT MAP (
        A => S5093,
        B => S5099,
        Y => S5100
    );
NOT_391: ENTITY WORK.NOT
    PORT MAP (
        A => S5100,
        Y => S5101
    );
NOR_1660: ENTITY WORK.NOR
    PORT MAP (
        A => S2717,
        B => S5101,
        Y => S5102
    );
NAND_3160: ENTITY WORK.NAND
    PORT MAP (
        A => S2718,
        B => S5100,
        Y => S5103
    );
NOR_1661: ENTITY WORK.NOR
    PORT MAP (
        A => S4907,
        B => S5102,
        Y => S5104
    );
NAND_3161: ENTITY WORK.NAND
    PORT MAP (
        A => S4908,
        B => S5103,
        Y => S5105
    );
NOR_1662: ENTITY WORK.NOR
    PORT MAP (
        A => S5091,
        B => S5105,
        Y => S5106
    );
NAND_3162: ENTITY WORK.NAND
    PORT MAP (
        A => S5092,
        B => S5104,
        Y => S5107
    );
NOR_1663: ENTITY WORK.NOR
    PORT MAP (
        A => S2718,
        B => S5100,
        Y => S5108
    );
NAND_3163: ENTITY WORK.NAND
    PORT MAP (
        A => S2717,
        B => S5101,
        Y => S5109
    );
NOR_1664: ENTITY WORK.NOR
    PORT MAP (
        A => S3905,
        B => S5108,
        Y => S5110
    );
NAND_3164: ENTITY WORK.NAND
    PORT MAP (
        A => S3904,
        B => S5109,
        Y => S5111
    );
NOR_1665: ENTITY WORK.NOR
    PORT MAP (
        A => S5106,
        B => S5111,
        Y => S5112
    );
NAND_3165: ENTITY WORK.NAND
    PORT MAP (
        A => S5107,
        B => S5110,
        Y => S5113
    );
NOR_1666: ENTITY WORK.NOR
    PORT MAP (
        A => S5102,
        B => S5108,
        Y => S5114
    );
NAND_3166: ENTITY WORK.NAND
    PORT MAP (
        A => S5103,
        B => S5109,
        Y => S5115
    );
NOR_1667: ENTITY WORK.NOR
    PORT MAP (
        A => S4907,
        B => S5091,
        Y => S5116
    );
NAND_3167: ENTITY WORK.NAND
    PORT MAP (
        A => S4908,
        B => S5092,
        Y => S5117
    );
NOR_1668: ENTITY WORK.NOR
    PORT MAP (
        A => S5114,
        B => S5117,
        Y => S5118
    );
NOR_1669: ENTITY WORK.NOR
    PORT MAP (
        A => S5115,
        B => S5116,
        Y => S5119
    );
NOR_1670: ENTITY WORK.NOR
    PORT MAP (
        A => S5118,
        B => S5119,
        Y => S5120
    );
NAND_3168: ENTITY WORK.NAND
    PORT MAP (
        A => S5112,
        B => S5120,
        Y => S5121
    );
NAND_3169: ENTITY WORK.NAND
    PORT MAP (
        A => S5100,
        B => S5113,
        Y => S5122
    );
NAND_3170: ENTITY WORK.NAND
    PORT MAP (
        A => S5121,
        B => S5122,
        Y => S5123
    );
NOR_1671: ENTITY WORK.NOR
    PORT MAP (
        A => S4911,
        B => S5089,
        Y => S5124
    );
NAND_3171: ENTITY WORK.NAND
    PORT MAP (
        A => S4912,
        B => S5090,
        Y => S5125
    );
NOR_1672: ENTITY WORK.NOR
    PORT MAP (
        A => S5091,
        B => S5124,
        Y => S5126
    );
NAND_3172: ENTITY WORK.NAND
    PORT MAP (
        A => S5092,
        B => S5125,
        Y => S5127
    );
NOR_1673: ENTITY WORK.NOR
    PORT MAP (
        A => S5113,
        B => S5126,
        Y => S5128
    );
NAND_3173: ENTITY WORK.NAND
    PORT MAP (
        A => S5112,
        B => S5127,
        Y => S5129
    );
NOR_1674: ENTITY WORK.NOR
    PORT MAP (
        A => S4905,
        B => S5112,
        Y => S5130
    );
NAND_3174: ENTITY WORK.NAND
    PORT MAP (
        A => S4906,
        B => S5113,
        Y => S5131
    );
NOR_1675: ENTITY WORK.NOR
    PORT MAP (
        A => S5128,
        B => S5130,
        Y => S5132
    );
NAND_3175: ENTITY WORK.NAND
    PORT MAP (
        A => S5129,
        B => S5131,
        Y => S5133
    );
NOR_1676: ENTITY WORK.NOR
    PORT MAP (
        A => S2717,
        B => S5133,
        Y => S5134
    );
NAND_3176: ENTITY WORK.NAND
    PORT MAP (
        A => S2718,
        B => S5132,
        Y => S5135
    );
NAND_3177: ENTITY WORK.NAND
    PORT MAP (
        A => S2717,
        B => S5133,
        Y => S5136
    );
NAND_3178: ENTITY WORK.NAND
    PORT MAP (
        A => S5135,
        B => S5136,
        Y => S5137
    );
NOT_392: ENTITY WORK.NOT
    PORT MAP (
        A => S5137,
        Y => S5138
    );
NOR_1677: ENTITY WORK.NOR
    PORT MAP (
        A => S4927,
        B => S4929,
        Y => S5139
    );
NAND_3179: ENTITY WORK.NAND
    PORT MAP (
        A => S4928,
        B => S4930,
        Y => S5140
    );
NOR_1678: ENTITY WORK.NOR
    PORT MAP (
        A => S5086,
        B => S5139,
        Y => S5141
    );
NOR_1679: ENTITY WORK.NOR
    PORT MAP (
        A => S5085,
        B => S5140,
        Y => S5142
    );
NOR_1680: ENTITY WORK.NOR
    PORT MAP (
        A => S5141,
        B => S5142,
        Y => S5143
    );
NOR_1681: ENTITY WORK.NOR
    PORT MAP (
        A => S5113,
        B => S5143,
        Y => S5144
    );
NOR_1682: ENTITY WORK.NOR
    PORT MAP (
        A => S4925,
        B => S5112,
        Y => S5145
    );
NOR_1683: ENTITY WORK.NOR
    PORT MAP (
        A => S5144,
        B => S5145,
        Y => S5146
    );
NOT_393: ENTITY WORK.NOT
    PORT MAP (
        A => S5146,
        Y => S5147
    );
NAND_3180: ENTITY WORK.NAND
    PORT MAP (
        A => S2617,
        B => S5147,
        Y => S5148
    );
NAND_3181: ENTITY WORK.NAND
    PORT MAP (
        A => S2618,
        B => S5146,
        Y => S5149
    );
NOR_1684: ENTITY WORK.NOR
    PORT MAP (
        A => S4945,
        B => S5082,
        Y => S5150
    );
NOR_1685: ENTITY WORK.NOR
    PORT MAP (
        A => S5083,
        B => S5150,
        Y => S5151
    );
NOR_1686: ENTITY WORK.NOR
    PORT MAP (
        A => S5113,
        B => S5151,
        Y => S5152
    );
NOR_1687: ENTITY WORK.NOR
    PORT MAP (
        A => S4939,
        B => S5112,
        Y => S5153
    );
NOR_1688: ENTITY WORK.NOR
    PORT MAP (
        A => S5152,
        B => S5153,
        Y => S5154
    );
NOT_394: ENTITY WORK.NOT
    PORT MAP (
        A => S5154,
        Y => S5155
    );
NOR_1689: ENTITY WORK.NOR
    PORT MAP (
        A => S2517,
        B => S5155,
        Y => S5156
    );
NAND_3182: ENTITY WORK.NAND
    PORT MAP (
        A => S2518,
        B => S5154,
        Y => S5157
    );
NOR_1690: ENTITY WORK.NOR
    PORT MAP (
        A => S2518,
        B => S5154,
        Y => S5158
    );
NOR_1691: ENTITY WORK.NOR
    PORT MAP (
        A => S5156,
        B => S5158,
        Y => S5159
    );
NOT_395: ENTITY WORK.NOT
    PORT MAP (
        A => S5159,
        Y => S5160
    );
NOR_1692: ENTITY WORK.NOR
    PORT MAP (
        A => S4957,
        B => S4959,
        Y => S5161
    );
NAND_3183: ENTITY WORK.NAND
    PORT MAP (
        A => S4958,
        B => S4960,
        Y => S5162
    );
NOR_1693: ENTITY WORK.NOR
    PORT MAP (
        A => S5077,
        B => S5161,
        Y => S5163
    );
NAND_3184: ENTITY WORK.NAND
    PORT MAP (
        A => S5078,
        B => S5162,
        Y => S5164
    );
NOR_1694: ENTITY WORK.NOR
    PORT MAP (
        A => S5078,
        B => S5162,
        Y => S5165
    );
NAND_3185: ENTITY WORK.NAND
    PORT MAP (
        A => S5077,
        B => S5161,
        Y => S5166
    );
NOR_1695: ENTITY WORK.NOR
    PORT MAP (
        A => S5163,
        B => S5165,
        Y => S5167
    );
NAND_3186: ENTITY WORK.NAND
    PORT MAP (
        A => S5164,
        B => S5166,
        Y => S5168
    );
NOR_1696: ENTITY WORK.NOR
    PORT MAP (
        A => S5113,
        B => S5168,
        Y => S5169
    );
NAND_3187: ENTITY WORK.NAND
    PORT MAP (
        A => S5112,
        B => S5167,
        Y => S5170
    );
NOR_1697: ENTITY WORK.NOR
    PORT MAP (
        A => S4955,
        B => S5112,
        Y => S5171
    );
NAND_3188: ENTITY WORK.NAND
    PORT MAP (
        A => S4956,
        B => S5113,
        Y => S5172
    );
NOR_1698: ENTITY WORK.NOR
    PORT MAP (
        A => S5169,
        B => S5171,
        Y => S5173
    );
NAND_3189: ENTITY WORK.NAND
    PORT MAP (
        A => S5170,
        B => S5172,
        Y => S5174
    );
NOR_1699: ENTITY WORK.NOR
    PORT MAP (
        A => S2417,
        B => S5174,
        Y => S5175
    );
NAND_3190: ENTITY WORK.NAND
    PORT MAP (
        A => S2418,
        B => S5173,
        Y => S5176
    );
NOR_1700: ENTITY WORK.NOR
    PORT MAP (
        A => S2418,
        B => S5173,
        Y => S5177
    );
NAND_3191: ENTITY WORK.NAND
    PORT MAP (
        A => S2417,
        B => S5174,
        Y => S5178
    );
NOR_1701: ENTITY WORK.NOR
    PORT MAP (
        A => S4975,
        B => S5074,
        Y => S5179
    );
NAND_3192: ENTITY WORK.NAND
    PORT MAP (
        A => S4976,
        B => S5073,
        Y => S5180
    );
NOR_1702: ENTITY WORK.NOR
    PORT MAP (
        A => S5075,
        B => S5179,
        Y => S5181
    );
NAND_3193: ENTITY WORK.NAND
    PORT MAP (
        A => S5076,
        B => S5180,
        Y => S5182
    );
NOR_1703: ENTITY WORK.NOR
    PORT MAP (
        A => S5113,
        B => S5181,
        Y => S5183
    );
NAND_3194: ENTITY WORK.NAND
    PORT MAP (
        A => S5112,
        B => S5182,
        Y => S5184
    );
NOR_1704: ENTITY WORK.NOR
    PORT MAP (
        A => S4969,
        B => S5112,
        Y => S5185
    );
NAND_3195: ENTITY WORK.NAND
    PORT MAP (
        A => S4970,
        B => S5113,
        Y => S5186
    );
NOR_1705: ENTITY WORK.NOR
    PORT MAP (
        A => S5183,
        B => S5185,
        Y => S5187
    );
NAND_3196: ENTITY WORK.NAND
    PORT MAP (
        A => S5184,
        B => S5186,
        Y => S5188
    );
NOR_1706: ENTITY WORK.NOR
    PORT MAP (
        A => S2311,
        B => S5188,
        Y => S5189
    );
NAND_3197: ENTITY WORK.NAND
    PORT MAP (
        A => S2312,
        B => S5187,
        Y => S5190
    );
NOR_1707: ENTITY WORK.NOR
    PORT MAP (
        A => S2312,
        B => S5187,
        Y => S5191
    );
NAND_3198: ENTITY WORK.NAND
    PORT MAP (
        A => S2311,
        B => S5188,
        Y => S5192
    );
NOR_1708: ENTITY WORK.NOR
    PORT MAP (
        A => S5189,
        B => S5191,
        Y => S5193
    );
NAND_3199: ENTITY WORK.NAND
    PORT MAP (
        A => S5190,
        B => S5192,
        Y => S5194
    );
NOR_1709: ENTITY WORK.NOR
    PORT MAP (
        A => S4987,
        B => S4989,
        Y => S5195
    );
NAND_3200: ENTITY WORK.NAND
    PORT MAP (
        A => S4988,
        B => S4990,
        Y => S5196
    );
NOR_1710: ENTITY WORK.NOR
    PORT MAP (
        A => S5070,
        B => S5195,
        Y => S5197
    );
NAND_3201: ENTITY WORK.NAND
    PORT MAP (
        A => S5069,
        B => S5196,
        Y => S5198
    );
NOR_1711: ENTITY WORK.NOR
    PORT MAP (
        A => S5069,
        B => S5196,
        Y => S5199
    );
NAND_3202: ENTITY WORK.NAND
    PORT MAP (
        A => S5070,
        B => S5195,
        Y => S5200
    );
NOR_1712: ENTITY WORK.NOR
    PORT MAP (
        A => S5197,
        B => S5199,
        Y => S5201
    );
NAND_3203: ENTITY WORK.NAND
    PORT MAP (
        A => S5198,
        B => S5200,
        Y => S5202
    );
NOR_1713: ENTITY WORK.NOR
    PORT MAP (
        A => S5113,
        B => S5201,
        Y => S5203
    );
NAND_3204: ENTITY WORK.NAND
    PORT MAP (
        A => S5112,
        B => S5202,
        Y => S5204
    );
NOR_1714: ENTITY WORK.NOR
    PORT MAP (
        A => S4985,
        B => S5112,
        Y => S5205
    );
NAND_3205: ENTITY WORK.NAND
    PORT MAP (
        A => S4986,
        B => S5113,
        Y => S5206
    );
NOR_1715: ENTITY WORK.NOR
    PORT MAP (
        A => S5203,
        B => S5205,
        Y => S5207
    );
NAND_3206: ENTITY WORK.NAND
    PORT MAP (
        A => S5204,
        B => S5206,
        Y => S5208
    );
NOR_1716: ENTITY WORK.NOR
    PORT MAP (
        A => S2205,
        B => S5208,
        Y => S5209
    );
NAND_3207: ENTITY WORK.NAND
    PORT MAP (
        A => S2206,
        B => S5207,
        Y => S5210
    );
NOR_1717: ENTITY WORK.NOR
    PORT MAP (
        A => S2206,
        B => S5207,
        Y => S5211
    );
NAND_3208: ENTITY WORK.NAND
    PORT MAP (
        A => S2205,
        B => S5208,
        Y => S5212
    );
NOR_1718: ENTITY WORK.NOR
    PORT MAP (
        A => S5062,
        B => S5065,
        Y => S5213
    );
NAND_3209: ENTITY WORK.NAND
    PORT MAP (
        A => S5061,
        B => S5066,
        Y => S5214
    );
NOR_1719: ENTITY WORK.NOR
    PORT MAP (
        A => S5067,
        B => S5213,
        Y => S5215
    );
NAND_3210: ENTITY WORK.NAND
    PORT MAP (
        A => S5068,
        B => S5214,
        Y => S5216
    );
NOR_1720: ENTITY WORK.NOR
    PORT MAP (
        A => S5113,
        B => S5215,
        Y => S5217
    );
NAND_3211: ENTITY WORK.NAND
    PORT MAP (
        A => S5112,
        B => S5216,
        Y => S5218
    );
NOR_1721: ENTITY WORK.NOR
    PORT MAP (
        A => S4999,
        B => S5112,
        Y => S5219
    );
NAND_3212: ENTITY WORK.NAND
    PORT MAP (
        A => S5000,
        B => S5113,
        Y => S5220
    );
NOR_1722: ENTITY WORK.NOR
    PORT MAP (
        A => S5217,
        B => S5219,
        Y => S5221
    );
NAND_3213: ENTITY WORK.NAND
    PORT MAP (
        A => S5218,
        B => S5220,
        Y => S5222
    );
NOR_1723: ENTITY WORK.NOR
    PORT MAP (
        A => S2106,
        B => S5222,
        Y => S5223
    );
NAND_3214: ENTITY WORK.NAND
    PORT MAP (
        A => S2107,
        B => S5221,
        Y => S5224
    );
NAND_3215: ENTITY WORK.NAND
    PORT MAP (
        A => S5012,
        B => S5113,
        Y => S5225
    );
NAND_3216: ENTITY WORK.NAND
    PORT MAP (
        A => S5018,
        B => S5057,
        Y => S5226
    );
NAND_3217: ENTITY WORK.NAND
    PORT MAP (
        A => S5060,
        B => S5226,
        Y => S5227
    );
NAND_3218: ENTITY WORK.NAND
    PORT MAP (
        A => S5112,
        B => S5227,
        Y => S5228
    );
NAND_3219: ENTITY WORK.NAND
    PORT MAP (
        A => S5225,
        B => S5228,
        Y => S5229
    );
NOT_396: ENTITY WORK.NOT
    PORT MAP (
        A => S5229,
        Y => S5230
    );
NOR_1724: ENTITY WORK.NOR
    PORT MAP (
        A => S1597,
        B => S5229,
        Y => S5231
    );
NAND_3220: ENTITY WORK.NAND
    PORT MAP (
        A => S1598,
        B => S5230,
        Y => S5232
    );
NAND_3221: ENTITY WORK.NAND
    PORT MAP (
        A => S1597,
        B => S5229,
        Y => S5233
    );
NAND_3222: ENTITY WORK.NAND
    PORT MAP (
        A => S5232,
        B => S5233,
        Y => S5234
    );
NOT_397: ENTITY WORK.NOT
    PORT MAP (
        A => S5234,
        Y => S5235
    );
NAND_3223: ENTITY WORK.NAND
    PORT MAP (
        A => S5034,
        B => S5053,
        Y => S5236
    );
NAND_3224: ENTITY WORK.NAND
    PORT MAP (
        A => S5056,
        B => S5236,
        Y => S5237
    );
NAND_3225: ENTITY WORK.NAND
    PORT MAP (
        A => S5112,
        B => S5237,
        Y => S5238
    );
NAND_3226: ENTITY WORK.NAND
    PORT MAP (
        A => S5028,
        B => S5113,
        Y => S5239
    );
NAND_3227: ENTITY WORK.NAND
    PORT MAP (
        A => S5238,
        B => S5239,
        Y => S5240
    );
NOT_398: ENTITY WORK.NOT
    PORT MAP (
        A => S5240,
        Y => S5241
    );
NOR_1725: ENTITY WORK.NOR
    PORT MAP (
        A => S1952,
        B => S5240,
        Y => S5242
    );
NAND_3228: ENTITY WORK.NAND
    PORT MAP (
        A => S1953,
        B => S5241,
        Y => S5243
    );
NAND_3229: ENTITY WORK.NAND
    PORT MAP (
        A => S1952,
        B => S5240,
        Y => S5244
    );
NAND_3230: ENTITY WORK.NAND
    PORT MAP (
        A => S5243,
        B => S5244,
        Y => S5245
    );
NOT_399: ENTITY WORK.NOT
    PORT MAP (
        A => S5245,
        Y => S5246
    );
NOR_1726: ENTITY WORK.NOR
    PORT MAP (
        A => S5046,
        B => S5049,
        Y => S5247
    );
NOR_1727: ENTITY WORK.NOR
    PORT MAP (
        A => S5051,
        B => S5247,
        Y => S5248
    );
NOR_1728: ENTITY WORK.NOR
    PORT MAP (
        A => S5113,
        B => S5248,
        Y => S5249
    );
NOR_1729: ENTITY WORK.NOR
    PORT MAP (
        A => S5042,
        B => S5112,
        Y => S5250
    );
NOR_1730: ENTITY WORK.NOR
    PORT MAP (
        A => S5249,
        B => S5250,
        Y => S5251
    );
NOT_400: ENTITY WORK.NOT
    PORT MAP (
        A => S5251,
        Y => S5252
    );
NOR_1731: ENTITY WORK.NOR
    PORT MAP (
        A => S1848,
        B => S5252,
        Y => S5253
    );
NAND_3231: ENTITY WORK.NAND
    PORT MAP (
        A => S1849,
        B => S5251,
        Y => S5254
    );
NOR_1732: ENTITY WORK.NOR
    PORT MAP (
        A => S1849,
        B => S5251,
        Y => S5255
    );
NAND_3232: ENTITY WORK.NAND
    PORT MAP (
        A => S1848,
        B => S5252,
        Y => S5256
    );
NOR_1733: ENTITY WORK.NOR
    PORT MAP (
        A => S1516,
        B => S5113,
        Y => S5257
    );
NAND_3233: ENTITY WORK.NAND
    PORT MAP (
        A => S1515,
        B => S5112,
        Y => S5258
    );
NOR_1734: ENTITY WORK.NOR
    PORT MAP (
        A => S1013,
        B => S5257,
        Y => S5259
    );
NAND_3234: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_4,
        B => S5258,
        Y => S5260
    );
NOR_1735: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_4,
        B => S5258,
        Y => S5261
    );
NAND_3235: ENTITY WORK.NAND
    PORT MAP (
        A => S1013,
        B => S5257,
        Y => S5262
    );
NOR_1736: ENTITY WORK.NOR
    PORT MAP (
        A => S5259,
        B => S5261,
        Y => S5263
    );
NAND_3236: ENTITY WORK.NAND
    PORT MAP (
        A => S5260,
        B => S5262,
        Y => S5264
    );
NOR_1737: ENTITY WORK.NOR
    PORT MAP (
        A => S1745,
        B => S5263,
        Y => S5265
    );
NAND_3237: ENTITY WORK.NAND
    PORT MAP (
        A => S1746,
        B => S5264,
        Y => S5266
    );
NOR_1738: ENTITY WORK.NOR
    PORT MAP (
        A => S1746,
        B => S5264,
        Y => S5267
    );
NAND_3238: ENTITY WORK.NAND
    PORT MAP (
        A => S1745,
        B => S5263,
        Y => S5268
    );
NOR_1739: ENTITY WORK.NOR
    PORT MAP (
        A => S5265,
        B => S5267,
        Y => S5269
    );
NAND_3239: ENTITY WORK.NAND
    PORT MAP (
        A => S5266,
        B => S5268,
        Y => S5270
    );
NOR_1740: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_3,
        B => S1516,
        Y => S5271
    );
NAND_3240: ENTITY WORK.NAND
    PORT MAP (
        A => S1065,
        B => S1515,
        Y => S5272
    );
NOR_1741: ENTITY WORK.NOR
    PORT MAP (
        A => S5270,
        B => S5271,
        Y => S5273
    );
NAND_3241: ENTITY WORK.NAND
    PORT MAP (
        A => S5269,
        B => S5272,
        Y => S5274
    );
NOR_1742: ENTITY WORK.NOR
    PORT MAP (
        A => S5265,
        B => S5273,
        Y => S5275
    );
NAND_3242: ENTITY WORK.NAND
    PORT MAP (
        A => S5266,
        B => S5274,
        Y => S5276
    );
NOR_1743: ENTITY WORK.NOR
    PORT MAP (
        A => S5255,
        B => S5275,
        Y => S5277
    );
NAND_3243: ENTITY WORK.NAND
    PORT MAP (
        A => S5256,
        B => S5276,
        Y => S5278
    );
NOR_1744: ENTITY WORK.NOR
    PORT MAP (
        A => S5253,
        B => S5277,
        Y => S5279
    );
NAND_3244: ENTITY WORK.NAND
    PORT MAP (
        A => S5254,
        B => S5278,
        Y => S5280
    );
NOR_1745: ENTITY WORK.NOR
    PORT MAP (
        A => S5245,
        B => S5279,
        Y => S5281
    );
NAND_3245: ENTITY WORK.NAND
    PORT MAP (
        A => S5246,
        B => S5280,
        Y => S5282
    );
NOR_1746: ENTITY WORK.NOR
    PORT MAP (
        A => S5242,
        B => S5281,
        Y => S5283
    );
NAND_3246: ENTITY WORK.NAND
    PORT MAP (
        A => S5243,
        B => S5282,
        Y => S5284
    );
NOR_1747: ENTITY WORK.NOR
    PORT MAP (
        A => S5234,
        B => S5283,
        Y => S5285
    );
NAND_3247: ENTITY WORK.NAND
    PORT MAP (
        A => S5235,
        B => S5284,
        Y => S5286
    );
NOR_1748: ENTITY WORK.NOR
    PORT MAP (
        A => S5231,
        B => S5285,
        Y => S5287
    );
NAND_3248: ENTITY WORK.NAND
    PORT MAP (
        A => S5232,
        B => S5286,
        Y => S5288
    );
NOR_1749: ENTITY WORK.NOR
    PORT MAP (
        A => S2107,
        B => S5221,
        Y => S5289
    );
NAND_3249: ENTITY WORK.NAND
    PORT MAP (
        A => S2106,
        B => S5222,
        Y => S5290
    );
NOR_1750: ENTITY WORK.NOR
    PORT MAP (
        A => S5223,
        B => S5289,
        Y => S5291
    );
NAND_3250: ENTITY WORK.NAND
    PORT MAP (
        A => S5224,
        B => S5290,
        Y => S5292
    );
NOR_1751: ENTITY WORK.NOR
    PORT MAP (
        A => S5287,
        B => S5292,
        Y => S5293
    );
NAND_3251: ENTITY WORK.NAND
    PORT MAP (
        A => S5288,
        B => S5291,
        Y => S5294
    );
NOR_1752: ENTITY WORK.NOR
    PORT MAP (
        A => S5223,
        B => S5293,
        Y => S5295
    );
NAND_3252: ENTITY WORK.NAND
    PORT MAP (
        A => S5224,
        B => S5294,
        Y => S5296
    );
NOR_1753: ENTITY WORK.NOR
    PORT MAP (
        A => S5211,
        B => S5295,
        Y => S5297
    );
NAND_3253: ENTITY WORK.NAND
    PORT MAP (
        A => S5212,
        B => S5296,
        Y => S5298
    );
NOR_1754: ENTITY WORK.NOR
    PORT MAP (
        A => S5209,
        B => S5297,
        Y => S5299
    );
NAND_3254: ENTITY WORK.NAND
    PORT MAP (
        A => S5210,
        B => S5298,
        Y => S5300
    );
NOR_1755: ENTITY WORK.NOR
    PORT MAP (
        A => S5194,
        B => S5299,
        Y => S5301
    );
NAND_3255: ENTITY WORK.NAND
    PORT MAP (
        A => S5193,
        B => S5300,
        Y => S5302
    );
NOR_1756: ENTITY WORK.NOR
    PORT MAP (
        A => S5189,
        B => S5301,
        Y => S5303
    );
NAND_3256: ENTITY WORK.NAND
    PORT MAP (
        A => S5190,
        B => S5302,
        Y => S5304
    );
NOR_1757: ENTITY WORK.NOR
    PORT MAP (
        A => S5177,
        B => S5303,
        Y => S5305
    );
NAND_3257: ENTITY WORK.NAND
    PORT MAP (
        A => S5178,
        B => S5304,
        Y => S5306
    );
NOR_1758: ENTITY WORK.NOR
    PORT MAP (
        A => S5175,
        B => S5305,
        Y => S5307
    );
NAND_3258: ENTITY WORK.NAND
    PORT MAP (
        A => S5176,
        B => S5306,
        Y => S5308
    );
NOR_1759: ENTITY WORK.NOR
    PORT MAP (
        A => S5160,
        B => S5307,
        Y => S5309
    );
NAND_3259: ENTITY WORK.NAND
    PORT MAP (
        A => S5159,
        B => S5308,
        Y => S5310
    );
NOR_1760: ENTITY WORK.NOR
    PORT MAP (
        A => S5156,
        B => S5309,
        Y => S5311
    );
NAND_3260: ENTITY WORK.NAND
    PORT MAP (
        A => S5157,
        B => S5310,
        Y => S5312
    );
NAND_3261: ENTITY WORK.NAND
    PORT MAP (
        A => S5149,
        B => S5311,
        Y => S5313
    );
NAND_3262: ENTITY WORK.NAND
    PORT MAP (
        A => S5148,
        B => S5312,
        Y => S5314
    );
NAND_3263: ENTITY WORK.NAND
    PORT MAP (
        A => S5149,
        B => S5314,
        Y => S5315
    );
NAND_3264: ENTITY WORK.NAND
    PORT MAP (
        A => S5148,
        B => S5313,
        Y => S5316
    );
NOR_1761: ENTITY WORK.NOR
    PORT MAP (
        A => S5137,
        B => S5316,
        Y => S5317
    );
NAND_3265: ENTITY WORK.NAND
    PORT MAP (
        A => S5138,
        B => S5315,
        Y => S5318
    );
NOR_1762: ENTITY WORK.NOR
    PORT MAP (
        A => S5134,
        B => S5317,
        Y => S5319
    );
NAND_3266: ENTITY WORK.NAND
    PORT MAP (
        A => S5135,
        B => S5318,
        Y => S5320
    );
NOR_1763: ENTITY WORK.NOR
    PORT MAP (
        A => S2817,
        B => S3903,
        Y => S5321
    );
NOR_1764: ENTITY WORK.NOR
    PORT MAP (
        A => S3905,
        B => S5320,
        Y => S5322
    );
NAND_3267: ENTITY WORK.NAND
    PORT MAP (
        A => S5320,
        B => S5321,
        Y => S5323
    );
NAND_3268: ENTITY WORK.NAND
    PORT MAP (
        A => S5123,
        B => S5323,
        Y => S5324
    );
NAND_3269: ENTITY WORK.NAND
    PORT MAP (
        A => S2817,
        B => S5123,
        Y => S5325
    );
NOT_401: ENTITY WORK.NOT
    PORT MAP (
        A => S5325,
        Y => S5326
    );
NOR_1765: ENTITY WORK.NOR
    PORT MAP (
        A => S5320,
        B => S5326,
        Y => S5327
    );
NAND_3270: ENTITY WORK.NAND
    PORT MAP (
        A => S5319,
        B => S5325,
        Y => S5328
    );
NOR_1766: ENTITY WORK.NOR
    PORT MAP (
        A => S2817,
        B => S5123,
        Y => S5329
    );
NOR_1767: ENTITY WORK.NOR
    PORT MAP (
        A => S3903,
        B => S5329,
        Y => S5330
    );
NOT_402: ENTITY WORK.NOT
    PORT MAP (
        A => S5330,
        Y => S5331
    );
NOR_1768: ENTITY WORK.NOR
    PORT MAP (
        A => S5327,
        B => S5331,
        Y => S5332
    );
NAND_3271: ENTITY WORK.NAND
    PORT MAP (
        A => S5328,
        B => S5330,
        Y => S5333
    );
NOR_1769: ENTITY WORK.NOR
    PORT MAP (
        A => S5322,
        B => S5324,
        Y => S5334
    );
NAND_3272: ENTITY WORK.NAND
    PORT MAP (
        A => S2920,
        B => S5334,
        Y => S5335
    );
NOT_403: ENTITY WORK.NOT
    PORT MAP (
        A => S5335,
        Y => S5336
    );
NAND_3273: ENTITY WORK.NAND
    PORT MAP (
        A => S5137,
        B => S5316,
        Y => S5337
    );
NAND_3274: ENTITY WORK.NAND
    PORT MAP (
        A => S5318,
        B => S5337,
        Y => S5338
    );
NAND_3275: ENTITY WORK.NAND
    PORT MAP (
        A => S5332,
        B => S5338,
        Y => S5339
    );
NAND_3276: ENTITY WORK.NAND
    PORT MAP (
        A => S5133,
        B => S5333,
        Y => S5340
    );
NAND_3277: ENTITY WORK.NAND
    PORT MAP (
        A => S5339,
        B => S5340,
        Y => S5341
    );
NOT_404: ENTITY WORK.NOT
    PORT MAP (
        A => S5341,
        Y => S5342
    );
NOR_1770: ENTITY WORK.NOR
    PORT MAP (
        A => S2816,
        B => S5341,
        Y => S5343
    );
NAND_3278: ENTITY WORK.NAND
    PORT MAP (
        A => S2817,
        B => S5342,
        Y => S5344
    );
NAND_3279: ENTITY WORK.NAND
    PORT MAP (
        A => S2816,
        B => S5341,
        Y => S5345
    );
NAND_3280: ENTITY WORK.NAND
    PORT MAP (
        A => S5344,
        B => S5345,
        Y => S5346
    );
NOT_405: ENTITY WORK.NOT
    PORT MAP (
        A => S5346,
        Y => S5347
    );
NAND_3281: ENTITY WORK.NAND
    PORT MAP (
        A => S5148,
        B => S5149,
        Y => S5348
    );
NAND_3282: ENTITY WORK.NAND
    PORT MAP (
        A => S5311,
        B => S5348,
        Y => S5349
    );
NOR_1771: ENTITY WORK.NOR
    PORT MAP (
        A => S5311,
        B => S5348,
        Y => S5350
    );
NOT_406: ENTITY WORK.NOT
    PORT MAP (
        A => S5350,
        Y => S5351
    );
NAND_3283: ENTITY WORK.NAND
    PORT MAP (
        A => S5349,
        B => S5351,
        Y => S5352
    );
NAND_3284: ENTITY WORK.NAND
    PORT MAP (
        A => S5332,
        B => S5352,
        Y => S5353
    );
NOT_407: ENTITY WORK.NOT
    PORT MAP (
        A => S5353,
        Y => S5354
    );
NOR_1772: ENTITY WORK.NOR
    PORT MAP (
        A => S5146,
        B => S5332,
        Y => S5355
    );
NOR_1773: ENTITY WORK.NOR
    PORT MAP (
        A => S5354,
        B => S5355,
        Y => S5356
    );
NOT_408: ENTITY WORK.NOT
    PORT MAP (
        A => S5356,
        Y => S5357
    );
NAND_3285: ENTITY WORK.NAND
    PORT MAP (
        A => S2717,
        B => S5357,
        Y => S5358
    );
NAND_3286: ENTITY WORK.NAND
    PORT MAP (
        A => S2718,
        B => S5356,
        Y => S5359
    );
NOR_1774: ENTITY WORK.NOR
    PORT MAP (
        A => S5159,
        B => S5308,
        Y => S5360
    );
NOR_1775: ENTITY WORK.NOR
    PORT MAP (
        A => S5309,
        B => S5360,
        Y => S5361
    );
NOR_1776: ENTITY WORK.NOR
    PORT MAP (
        A => S5333,
        B => S5361,
        Y => S5362
    );
NOR_1777: ENTITY WORK.NOR
    PORT MAP (
        A => S5154,
        B => S5332,
        Y => S5363
    );
NOR_1778: ENTITY WORK.NOR
    PORT MAP (
        A => S5362,
        B => S5363,
        Y => S5364
    );
NOT_409: ENTITY WORK.NOT
    PORT MAP (
        A => S5364,
        Y => S5365
    );
NOR_1779: ENTITY WORK.NOR
    PORT MAP (
        A => S2617,
        B => S5365,
        Y => S5366
    );
NOT_410: ENTITY WORK.NOT
    PORT MAP (
        A => S5366,
        Y => S5367
    );
NOR_1780: ENTITY WORK.NOR
    PORT MAP (
        A => S2618,
        B => S5364,
        Y => S5368
    );
NOR_1781: ENTITY WORK.NOR
    PORT MAP (
        A => S5366,
        B => S5368,
        Y => S5369
    );
NOT_411: ENTITY WORK.NOT
    PORT MAP (
        A => S5369,
        Y => S5370
    );
NOR_1782: ENTITY WORK.NOR
    PORT MAP (
        A => S5175,
        B => S5177,
        Y => S5371
    );
NAND_3287: ENTITY WORK.NAND
    PORT MAP (
        A => S5176,
        B => S5178,
        Y => S5372
    );
NOR_1783: ENTITY WORK.NOR
    PORT MAP (
        A => S5304,
        B => S5371,
        Y => S5373
    );
NOR_1784: ENTITY WORK.NOR
    PORT MAP (
        A => S5303,
        B => S5372,
        Y => S5374
    );
NOR_1785: ENTITY WORK.NOR
    PORT MAP (
        A => S5373,
        B => S5374,
        Y => S5375
    );
NOR_1786: ENTITY WORK.NOR
    PORT MAP (
        A => S5174,
        B => S5332,
        Y => S5376
    );
NAND_3288: ENTITY WORK.NAND
    PORT MAP (
        A => S5173,
        B => S5333,
        Y => S5377
    );
NAND_3289: ENTITY WORK.NAND
    PORT MAP (
        A => S5332,
        B => S5375,
        Y => S5378
    );
NOT_412: ENTITY WORK.NOT
    PORT MAP (
        A => S5378,
        Y => S5379
    );
NAND_3290: ENTITY WORK.NAND
    PORT MAP (
        A => S5377,
        B => S5378,
        Y => S5380
    );
NOR_1787: ENTITY WORK.NOR
    PORT MAP (
        A => S5376,
        B => S5379,
        Y => S5381
    );
NOR_1788: ENTITY WORK.NOR
    PORT MAP (
        A => S2518,
        B => S5380,
        Y => S5382
    );
NOR_1789: ENTITY WORK.NOR
    PORT MAP (
        A => S2517,
        B => S5381,
        Y => S5383
    );
NAND_3291: ENTITY WORK.NAND
    PORT MAP (
        A => S5194,
        B => S5299,
        Y => S5384
    );
NAND_3292: ENTITY WORK.NAND
    PORT MAP (
        A => S5302,
        B => S5384,
        Y => S5385
    );
NAND_3293: ENTITY WORK.NAND
    PORT MAP (
        A => S5332,
        B => S5385,
        Y => S5386
    );
NAND_3294: ENTITY WORK.NAND
    PORT MAP (
        A => S5188,
        B => S5333,
        Y => S5387
    );
NAND_3295: ENTITY WORK.NAND
    PORT MAP (
        A => S5386,
        B => S5387,
        Y => S5388
    );
NOT_413: ENTITY WORK.NOT
    PORT MAP (
        A => S5388,
        Y => S5389
    );
NOR_1790: ENTITY WORK.NOR
    PORT MAP (
        A => S2417,
        B => S5388,
        Y => S5390
    );
NAND_3296: ENTITY WORK.NAND
    PORT MAP (
        A => S2418,
        B => S5389,
        Y => S5391
    );
NAND_3297: ENTITY WORK.NAND
    PORT MAP (
        A => S2417,
        B => S5388,
        Y => S5392
    );
NAND_3298: ENTITY WORK.NAND
    PORT MAP (
        A => S5391,
        B => S5392,
        Y => S5393
    );
NOT_414: ENTITY WORK.NOT
    PORT MAP (
        A => S5393,
        Y => S5394
    );
NOR_1791: ENTITY WORK.NOR
    PORT MAP (
        A => S5209,
        B => S5211,
        Y => S5395
    );
NAND_3299: ENTITY WORK.NAND
    PORT MAP (
        A => S5210,
        B => S5212,
        Y => S5396
    );
NOR_1792: ENTITY WORK.NOR
    PORT MAP (
        A => S5296,
        B => S5395,
        Y => S5397
    );
NOR_1793: ENTITY WORK.NOR
    PORT MAP (
        A => S5295,
        B => S5396,
        Y => S5398
    );
NOR_1794: ENTITY WORK.NOR
    PORT MAP (
        A => S5397,
        B => S5398,
        Y => S5399
    );
NOR_1795: ENTITY WORK.NOR
    PORT MAP (
        A => S5333,
        B => S5399,
        Y => S5400
    );
NOR_1796: ENTITY WORK.NOR
    PORT MAP (
        A => S5207,
        B => S5332,
        Y => S5401
    );
NOR_1797: ENTITY WORK.NOR
    PORT MAP (
        A => S5400,
        B => S5401,
        Y => S5402
    );
NOT_415: ENTITY WORK.NOT
    PORT MAP (
        A => S5402,
        Y => S5403
    );
NOR_1798: ENTITY WORK.NOR
    PORT MAP (
        A => S2311,
        B => S5403,
        Y => S5404
    );
NOR_1799: ENTITY WORK.NOR
    PORT MAP (
        A => S2312,
        B => S5402,
        Y => S5405
    );
NOR_1800: ENTITY WORK.NOR
    PORT MAP (
        A => S5288,
        B => S5291,
        Y => S5406
    );
NOT_416: ENTITY WORK.NOT
    PORT MAP (
        A => S5406,
        Y => S5407
    );
NAND_3300: ENTITY WORK.NAND
    PORT MAP (
        A => S5294,
        B => S5407,
        Y => S5408
    );
NAND_3301: ENTITY WORK.NAND
    PORT MAP (
        A => S5332,
        B => S5408,
        Y => S5409
    );
NAND_3302: ENTITY WORK.NAND
    PORT MAP (
        A => S5222,
        B => S5333,
        Y => S5410
    );
NAND_3303: ENTITY WORK.NAND
    PORT MAP (
        A => S5409,
        B => S5410,
        Y => S5411
    );
NOT_417: ENTITY WORK.NOT
    PORT MAP (
        A => S5411,
        Y => S5412
    );
NOR_1801: ENTITY WORK.NOR
    PORT MAP (
        A => S2205,
        B => S5411,
        Y => S5413
    );
NAND_3304: ENTITY WORK.NAND
    PORT MAP (
        A => S2206,
        B => S5412,
        Y => S5414
    );
NAND_3305: ENTITY WORK.NAND
    PORT MAP (
        A => S5234,
        B => S5283,
        Y => S5415
    );
NAND_3306: ENTITY WORK.NAND
    PORT MAP (
        A => S5286,
        B => S5415,
        Y => S5416
    );
NAND_3307: ENTITY WORK.NAND
    PORT MAP (
        A => S5332,
        B => S5416,
        Y => S5417
    );
NAND_3308: ENTITY WORK.NAND
    PORT MAP (
        A => S5229,
        B => S5333,
        Y => S5418
    );
NAND_3309: ENTITY WORK.NAND
    PORT MAP (
        A => S5417,
        B => S5418,
        Y => S5419
    );
NOT_418: ENTITY WORK.NOT
    PORT MAP (
        A => S5419,
        Y => S5420
    );
NAND_3310: ENTITY WORK.NAND
    PORT MAP (
        A => S2107,
        B => S5420,
        Y => S5421
    );
NOT_419: ENTITY WORK.NOT
    PORT MAP (
        A => S5421,
        Y => S5422
    );
NAND_3311: ENTITY WORK.NAND
    PORT MAP (
        A => S2106,
        B => S5419,
        Y => S5423
    );
NAND_3312: ENTITY WORK.NAND
    PORT MAP (
        A => S5421,
        B => S5423,
        Y => S5424
    );
NOT_420: ENTITY WORK.NOT
    PORT MAP (
        A => S5424,
        Y => S5425
    );
NAND_3313: ENTITY WORK.NAND
    PORT MAP (
        A => S5245,
        B => S5279,
        Y => S5426
    );
NAND_3314: ENTITY WORK.NAND
    PORT MAP (
        A => S5282,
        B => S5426,
        Y => S5427
    );
NAND_3315: ENTITY WORK.NAND
    PORT MAP (
        A => S5332,
        B => S5427,
        Y => S5428
    );
NAND_3316: ENTITY WORK.NAND
    PORT MAP (
        A => S5240,
        B => S5333,
        Y => S5429
    );
NAND_3317: ENTITY WORK.NAND
    PORT MAP (
        A => S5428,
        B => S5429,
        Y => S5430
    );
NOT_421: ENTITY WORK.NOT
    PORT MAP (
        A => S5430,
        Y => S5431
    );
NAND_3318: ENTITY WORK.NAND
    PORT MAP (
        A => S1598,
        B => S5431,
        Y => S5432
    );
NOT_422: ENTITY WORK.NOT
    PORT MAP (
        A => S5432,
        Y => S5433
    );
NAND_3319: ENTITY WORK.NAND
    PORT MAP (
        A => S1597,
        B => S5430,
        Y => S5434
    );
NAND_3320: ENTITY WORK.NAND
    PORT MAP (
        A => S5432,
        B => S5434,
        Y => S5435
    );
NOT_423: ENTITY WORK.NOT
    PORT MAP (
        A => S5435,
        Y => S5436
    );
NOR_1802: ENTITY WORK.NOR
    PORT MAP (
        A => S5253,
        B => S5255,
        Y => S5437
    );
NAND_3321: ENTITY WORK.NAND
    PORT MAP (
        A => S5254,
        B => S5256,
        Y => S5438
    );
NAND_3322: ENTITY WORK.NAND
    PORT MAP (
        A => S5275,
        B => S5437,
        Y => S5439
    );
NAND_3323: ENTITY WORK.NAND
    PORT MAP (
        A => S5276,
        B => S5438,
        Y => S5440
    );
NAND_3324: ENTITY WORK.NAND
    PORT MAP (
        A => S5439,
        B => S5440,
        Y => S5441
    );
NAND_3325: ENTITY WORK.NAND
    PORT MAP (
        A => S5332,
        B => S5441,
        Y => S5442
    );
NAND_3326: ENTITY WORK.NAND
    PORT MAP (
        A => S5251,
        B => S5333,
        Y => S5443
    );
NAND_3327: ENTITY WORK.NAND
    PORT MAP (
        A => S5442,
        B => S5443,
        Y => S5444
    );
NOT_424: ENTITY WORK.NOT
    PORT MAP (
        A => S5444,
        Y => S5445
    );
NOR_1803: ENTITY WORK.NOR
    PORT MAP (
        A => S1952,
        B => S5445,
        Y => S5446
    );
NAND_3328: ENTITY WORK.NAND
    PORT MAP (
        A => S1953,
        B => S5444,
        Y => S5447
    );
NOR_1804: ENTITY WORK.NOR
    PORT MAP (
        A => S1953,
        B => S5444,
        Y => S5448
    );
NAND_3329: ENTITY WORK.NAND
    PORT MAP (
        A => S1952,
        B => S5445,
        Y => S5449
    );
NOR_1805: ENTITY WORK.NOR
    PORT MAP (
        A => S5269,
        B => S5272,
        Y => S5450
    );
NOR_1806: ENTITY WORK.NOR
    PORT MAP (
        A => S5273,
        B => S5450,
        Y => S5451
    );
NAND_3330: ENTITY WORK.NAND
    PORT MAP (
        A => S5332,
        B => S5451,
        Y => S5452
    );
NOT_425: ENTITY WORK.NOT
    PORT MAP (
        A => S5452,
        Y => S5453
    );
NOR_1807: ENTITY WORK.NOR
    PORT MAP (
        A => S5263,
        B => S5332,
        Y => S5454
    );
NOT_426: ENTITY WORK.NOT
    PORT MAP (
        A => S5454,
        Y => S5455
    );
NOR_1808: ENTITY WORK.NOR
    PORT MAP (
        A => S5453,
        B => S5454,
        Y => S5456
    );
NAND_3331: ENTITY WORK.NAND
    PORT MAP (
        A => S5452,
        B => S5455,
        Y => S5457
    );
NOR_1809: ENTITY WORK.NOR
    PORT MAP (
        A => S1848,
        B => S5456,
        Y => S5458
    );
NAND_3332: ENTITY WORK.NAND
    PORT MAP (
        A => S1849,
        B => S5457,
        Y => S5459
    );
NOR_1810: ENTITY WORK.NOR
    PORT MAP (
        A => S1849,
        B => S5457,
        Y => S5460
    );
NAND_3333: ENTITY WORK.NAND
    PORT MAP (
        A => S1848,
        B => S5456,
        Y => S5461
    );
NOR_1811: ENTITY WORK.NOR
    PORT MAP (
        A => S5458,
        B => S5460,
        Y => S5462
    );
NAND_3334: ENTITY WORK.NAND
    PORT MAP (
        A => S5459,
        B => S5461,
        Y => S5463
    );
NOR_1812: ENTITY WORK.NOR
    PORT MAP (
        A => S1516,
        B => S5333,
        Y => S5464
    );
NAND_3335: ENTITY WORK.NAND
    PORT MAP (
        A => S1515,
        B => S5332,
        Y => S5465
    );
NOR_1813: ENTITY WORK.NOR
    PORT MAP (
        A => S1065,
        B => S5464,
        Y => S5466
    );
NAND_3336: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_3,
        B => S5465,
        Y => S5467
    );
NAND_3337: ENTITY WORK.NAND
    PORT MAP (
        A => S5271,
        B => S5332,
        Y => S5468
    );
NOT_427: ENTITY WORK.NOT
    PORT MAP (
        A => S5468,
        Y => S5469
    );
NOR_1814: ENTITY WORK.NOR
    PORT MAP (
        A => S5466,
        B => S5469,
        Y => S5470
    );
NAND_3338: ENTITY WORK.NAND
    PORT MAP (
        A => S5467,
        B => S5468,
        Y => S5471
    );
NOR_1815: ENTITY WORK.NOR
    PORT MAP (
        A => S1745,
        B => S5470,
        Y => S5472
    );
NAND_3339: ENTITY WORK.NAND
    PORT MAP (
        A => S1746,
        B => S5471,
        Y => S5473
    );
NOR_1816: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_2,
        B => S1516,
        Y => S5474
    );
NAND_3340: ENTITY WORK.NAND
    PORT MAP (
        A => S1116,
        B => S1515,
        Y => S5475
    );
NOR_1817: ENTITY WORK.NOR
    PORT MAP (
        A => S1746,
        B => S5471,
        Y => S5476
    );
NAND_3341: ENTITY WORK.NAND
    PORT MAP (
        A => S1745,
        B => S5470,
        Y => S5477
    );
NOR_1818: ENTITY WORK.NOR
    PORT MAP (
        A => S5472,
        B => S5476,
        Y => S5478
    );
NAND_3342: ENTITY WORK.NAND
    PORT MAP (
        A => S5473,
        B => S5477,
        Y => S5479
    );
NOR_1819: ENTITY WORK.NOR
    PORT MAP (
        A => S5474,
        B => S5479,
        Y => S5480
    );
NAND_3343: ENTITY WORK.NAND
    PORT MAP (
        A => S5475,
        B => S5478,
        Y => S5481
    );
NOR_1820: ENTITY WORK.NOR
    PORT MAP (
        A => S5472,
        B => S5480,
        Y => S5482
    );
NAND_3344: ENTITY WORK.NAND
    PORT MAP (
        A => S5473,
        B => S5481,
        Y => S5483
    );
NOR_1821: ENTITY WORK.NOR
    PORT MAP (
        A => S5463,
        B => S5482,
        Y => S5484
    );
NAND_3345: ENTITY WORK.NAND
    PORT MAP (
        A => S5462,
        B => S5483,
        Y => S5485
    );
NOR_1822: ENTITY WORK.NOR
    PORT MAP (
        A => S5458,
        B => S5484,
        Y => S5486
    );
NAND_3346: ENTITY WORK.NAND
    PORT MAP (
        A => S5459,
        B => S5485,
        Y => S5487
    );
NOR_1823: ENTITY WORK.NOR
    PORT MAP (
        A => S5448,
        B => S5486,
        Y => S5488
    );
NAND_3347: ENTITY WORK.NAND
    PORT MAP (
        A => S5449,
        B => S5487,
        Y => S5489
    );
NOR_1824: ENTITY WORK.NOR
    PORT MAP (
        A => S5446,
        B => S5488,
        Y => S5490
    );
NAND_3348: ENTITY WORK.NAND
    PORT MAP (
        A => S5447,
        B => S5489,
        Y => S5491
    );
NOR_1825: ENTITY WORK.NOR
    PORT MAP (
        A => S5435,
        B => S5490,
        Y => S5492
    );
NAND_3349: ENTITY WORK.NAND
    PORT MAP (
        A => S5436,
        B => S5491,
        Y => S5493
    );
NOR_1826: ENTITY WORK.NOR
    PORT MAP (
        A => S5433,
        B => S5492,
        Y => S5494
    );
NAND_3350: ENTITY WORK.NAND
    PORT MAP (
        A => S5432,
        B => S5493,
        Y => S5495
    );
NOR_1827: ENTITY WORK.NOR
    PORT MAP (
        A => S5424,
        B => S5494,
        Y => S5496
    );
NAND_3351: ENTITY WORK.NAND
    PORT MAP (
        A => S5425,
        B => S5495,
        Y => S5497
    );
NOR_1828: ENTITY WORK.NOR
    PORT MAP (
        A => S5422,
        B => S5496,
        Y => S5498
    );
NAND_3352: ENTITY WORK.NAND
    PORT MAP (
        A => S5421,
        B => S5497,
        Y => S5499
    );
NAND_3353: ENTITY WORK.NAND
    PORT MAP (
        A => S2205,
        B => S5411,
        Y => S5500
    );
NOT_428: ENTITY WORK.NOT
    PORT MAP (
        A => S5500,
        Y => S5501
    );
NOR_1829: ENTITY WORK.NOR
    PORT MAP (
        A => S5413,
        B => S5501,
        Y => S5502
    );
NOT_429: ENTITY WORK.NOT
    PORT MAP (
        A => S5502,
        Y => S5503
    );
NOR_1830: ENTITY WORK.NOR
    PORT MAP (
        A => S5498,
        B => S5503,
        Y => S5504
    );
NAND_3354: ENTITY WORK.NAND
    PORT MAP (
        A => S5499,
        B => S5502,
        Y => S5505
    );
NOR_1831: ENTITY WORK.NOR
    PORT MAP (
        A => S5413,
        B => S5504,
        Y => S5506
    );
NAND_3355: ENTITY WORK.NAND
    PORT MAP (
        A => S5414,
        B => S5505,
        Y => S5507
    );
NOR_1832: ENTITY WORK.NOR
    PORT MAP (
        A => S5405,
        B => S5506,
        Y => S5508
    );
NOR_1833: ENTITY WORK.NOR
    PORT MAP (
        A => S5404,
        B => S5507,
        Y => S5509
    );
NOR_1834: ENTITY WORK.NOR
    PORT MAP (
        A => S5404,
        B => S5508,
        Y => S5510
    );
NOR_1835: ENTITY WORK.NOR
    PORT MAP (
        A => S5405,
        B => S5509,
        Y => S5511
    );
NOR_1836: ENTITY WORK.NOR
    PORT MAP (
        A => S5393,
        B => S5510,
        Y => S5512
    );
NAND_3356: ENTITY WORK.NAND
    PORT MAP (
        A => S5394,
        B => S5511,
        Y => S5513
    );
NOR_1837: ENTITY WORK.NOR
    PORT MAP (
        A => S5390,
        B => S5512,
        Y => S5514
    );
NAND_3357: ENTITY WORK.NAND
    PORT MAP (
        A => S5391,
        B => S5513,
        Y => S5515
    );
NOR_1838: ENTITY WORK.NOR
    PORT MAP (
        A => S5383,
        B => S5515,
        Y => S5516
    );
NOR_1839: ENTITY WORK.NOR
    PORT MAP (
        A => S5382,
        B => S5514,
        Y => S5517
    );
NOR_1840: ENTITY WORK.NOR
    PORT MAP (
        A => S5382,
        B => S5516,
        Y => S5518
    );
NOR_1841: ENTITY WORK.NOR
    PORT MAP (
        A => S5383,
        B => S5517,
        Y => S5519
    );
NOR_1842: ENTITY WORK.NOR
    PORT MAP (
        A => S5370,
        B => S5519,
        Y => S5520
    );
NAND_3358: ENTITY WORK.NAND
    PORT MAP (
        A => S5369,
        B => S5518,
        Y => S5521
    );
NOR_1843: ENTITY WORK.NOR
    PORT MAP (
        A => S5366,
        B => S5520,
        Y => S5522
    );
NAND_3359: ENTITY WORK.NAND
    PORT MAP (
        A => S5367,
        B => S5521,
        Y => S5523
    );
NAND_3360: ENTITY WORK.NAND
    PORT MAP (
        A => S5359,
        B => S5522,
        Y => S5524
    );
NAND_3361: ENTITY WORK.NAND
    PORT MAP (
        A => S5358,
        B => S5523,
        Y => S5525
    );
NAND_3362: ENTITY WORK.NAND
    PORT MAP (
        A => S5359,
        B => S5525,
        Y => S5526
    );
NAND_3363: ENTITY WORK.NAND
    PORT MAP (
        A => S5358,
        B => S5524,
        Y => S5527
    );
NOR_1844: ENTITY WORK.NOR
    PORT MAP (
        A => S5346,
        B => S5527,
        Y => S5528
    );
NAND_3364: ENTITY WORK.NAND
    PORT MAP (
        A => S5347,
        B => S5526,
        Y => S5529
    );
NOR_1845: ENTITY WORK.NOR
    PORT MAP (
        A => S5343,
        B => S5528,
        Y => S5530
    );
NAND_3365: ENTITY WORK.NAND
    PORT MAP (
        A => S5344,
        B => S5529,
        Y => S5531
    );
NOR_1846: ENTITY WORK.NOR
    PORT MAP (
        A => S5336,
        B => S5531,
        Y => S5532
    );
NAND_3366: ENTITY WORK.NAND
    PORT MAP (
        A => S5335,
        B => S5530,
        Y => S5533
    );
NOR_1847: ENTITY WORK.NOR
    PORT MAP (
        A => S2920,
        B => S5334,
        Y => S5534
    );
NOT_430: ENTITY WORK.NOT
    PORT MAP (
        A => S5534,
        Y => S5535
    );
NOR_1848: ENTITY WORK.NOR
    PORT MAP (
        A => S3901,
        B => S5534,
        Y => S5536
    );
NAND_3367: ENTITY WORK.NAND
    PORT MAP (
        A => S3900,
        B => S5535,
        Y => S5537
    );
NOR_1849: ENTITY WORK.NOR
    PORT MAP (
        A => S5532,
        B => S5537,
        Y => S5538
    );
NAND_3368: ENTITY WORK.NAND
    PORT MAP (
        A => S5533,
        B => S5536,
        Y => S5539
    );
NAND_3369: ENTITY WORK.NAND
    PORT MAP (
        A => S5346,
        B => S5527,
        Y => S5540
    );
NAND_3370: ENTITY WORK.NAND
    PORT MAP (
        A => S5529,
        B => S5540,
        Y => S5541
    );
NAND_3371: ENTITY WORK.NAND
    PORT MAP (
        A => S5538,
        B => S5541,
        Y => S5542
    );
NAND_3372: ENTITY WORK.NAND
    PORT MAP (
        A => S5341,
        B => S5539,
        Y => S5543
    );
NAND_3373: ENTITY WORK.NAND
    PORT MAP (
        A => S5542,
        B => S5543,
        Y => S5544
    );
NOT_431: ENTITY WORK.NOT
    PORT MAP (
        A => S5544,
        Y => S5545
    );
NAND_3374: ENTITY WORK.NAND
    PORT MAP (
        A => S2920,
        B => S5545,
        Y => S5546
    );
NOT_432: ENTITY WORK.NOT
    PORT MAP (
        A => S5546,
        Y => S5547
    );
NAND_3375: ENTITY WORK.NAND
    PORT MAP (
        A => S2919,
        B => S5544,
        Y => S5548
    );
NAND_3376: ENTITY WORK.NAND
    PORT MAP (
        A => S5546,
        B => S5548,
        Y => S5549
    );
NOT_433: ENTITY WORK.NOT
    PORT MAP (
        A => S5549,
        Y => S5550
    );
NAND_3377: ENTITY WORK.NAND
    PORT MAP (
        A => S5358,
        B => S5359,
        Y => S5551
    );
NAND_3378: ENTITY WORK.NAND
    PORT MAP (
        A => S5522,
        B => S5551,
        Y => S5552
    );
NOT_434: ENTITY WORK.NOT
    PORT MAP (
        A => S5552,
        Y => S5553
    );
NOR_1850: ENTITY WORK.NOR
    PORT MAP (
        A => S5522,
        B => S5551,
        Y => S5554
    );
NOR_1851: ENTITY WORK.NOR
    PORT MAP (
        A => S5553,
        B => S5554,
        Y => S5555
    );
NOR_1852: ENTITY WORK.NOR
    PORT MAP (
        A => S5539,
        B => S5555,
        Y => S5556
    );
NOR_1853: ENTITY WORK.NOR
    PORT MAP (
        A => S5356,
        B => S5538,
        Y => S5557
    );
NOR_1854: ENTITY WORK.NOR
    PORT MAP (
        A => S5556,
        B => S5557,
        Y => S5558
    );
NOT_435: ENTITY WORK.NOT
    PORT MAP (
        A => S5558,
        Y => S5559
    );
NAND_3379: ENTITY WORK.NAND
    PORT MAP (
        A => S2817,
        B => S5558,
        Y => S5560
    );
NAND_3380: ENTITY WORK.NAND
    PORT MAP (
        A => S2816,
        B => S5559,
        Y => S5561
    );
NOR_1855: ENTITY WORK.NOR
    PORT MAP (
        A => S5369,
        B => S5518,
        Y => S5562
    );
NOR_1856: ENTITY WORK.NOR
    PORT MAP (
        A => S5520,
        B => S5562,
        Y => S5563
    );
NOR_1857: ENTITY WORK.NOR
    PORT MAP (
        A => S5539,
        B => S5563,
        Y => S5564
    );
NOR_1858: ENTITY WORK.NOR
    PORT MAP (
        A => S5364,
        B => S5538,
        Y => S5565
    );
NOR_1859: ENTITY WORK.NOR
    PORT MAP (
        A => S5564,
        B => S5565,
        Y => S5566
    );
NOT_436: ENTITY WORK.NOT
    PORT MAP (
        A => S5566,
        Y => S5567
    );
NOR_1860: ENTITY WORK.NOR
    PORT MAP (
        A => S2717,
        B => S5567,
        Y => S5568
    );
NOT_437: ENTITY WORK.NOT
    PORT MAP (
        A => S5568,
        Y => S5569
    );
NOR_1861: ENTITY WORK.NOR
    PORT MAP (
        A => S2718,
        B => S5566,
        Y => S5570
    );
NOR_1862: ENTITY WORK.NOR
    PORT MAP (
        A => S5568,
        B => S5570,
        Y => S5571
    );
NOT_438: ENTITY WORK.NOT
    PORT MAP (
        A => S5571,
        Y => S5572
    );
NOR_1863: ENTITY WORK.NOR
    PORT MAP (
        A => S5382,
        B => S5383,
        Y => S5573
    );
NOR_1864: ENTITY WORK.NOR
    PORT MAP (
        A => S5515,
        B => S5573,
        Y => S5574
    );
NOT_439: ENTITY WORK.NOT
    PORT MAP (
        A => S5574,
        Y => S5575
    );
NAND_3381: ENTITY WORK.NAND
    PORT MAP (
        A => S5515,
        B => S5573,
        Y => S5576
    );
NOT_440: ENTITY WORK.NOT
    PORT MAP (
        A => S5576,
        Y => S5577
    );
NOR_1865: ENTITY WORK.NOR
    PORT MAP (
        A => S5574,
        B => S5577,
        Y => S5578
    );
NAND_3382: ENTITY WORK.NAND
    PORT MAP (
        A => S5575,
        B => S5576,
        Y => S5579
    );
NOR_1866: ENTITY WORK.NOR
    PORT MAP (
        A => S5539,
        B => S5578,
        Y => S5580
    );
NAND_3383: ENTITY WORK.NAND
    PORT MAP (
        A => S5538,
        B => S5579,
        Y => S5581
    );
NOR_1867: ENTITY WORK.NOR
    PORT MAP (
        A => S5380,
        B => S5538,
        Y => S5582
    );
NAND_3384: ENTITY WORK.NAND
    PORT MAP (
        A => S5381,
        B => S5539,
        Y => S5583
    );
NOR_1868: ENTITY WORK.NOR
    PORT MAP (
        A => S5580,
        B => S5582,
        Y => S5584
    );
NAND_3385: ENTITY WORK.NAND
    PORT MAP (
        A => S5581,
        B => S5583,
        Y => S5585
    );
NAND_3386: ENTITY WORK.NAND
    PORT MAP (
        A => S2618,
        B => S5584,
        Y => S5586
    );
NAND_3387: ENTITY WORK.NAND
    PORT MAP (
        A => S2617,
        B => S5585,
        Y => S5587
    );
NAND_3388: ENTITY WORK.NAND
    PORT MAP (
        A => S5393,
        B => S5510,
        Y => S5588
    );
NAND_3389: ENTITY WORK.NAND
    PORT MAP (
        A => S5513,
        B => S5588,
        Y => S5589
    );
NAND_3390: ENTITY WORK.NAND
    PORT MAP (
        A => S5538,
        B => S5589,
        Y => S5590
    );
NAND_3391: ENTITY WORK.NAND
    PORT MAP (
        A => S5388,
        B => S5539,
        Y => S5591
    );
NAND_3392: ENTITY WORK.NAND
    PORT MAP (
        A => S5590,
        B => S5591,
        Y => S5592
    );
NOT_441: ENTITY WORK.NOT
    PORT MAP (
        A => S5592,
        Y => S5593
    );
NAND_3393: ENTITY WORK.NAND
    PORT MAP (
        A => S2518,
        B => S5593,
        Y => S5594
    );
NOT_442: ENTITY WORK.NOT
    PORT MAP (
        A => S5594,
        Y => S5595
    );
NAND_3394: ENTITY WORK.NAND
    PORT MAP (
        A => S2517,
        B => S5592,
        Y => S5596
    );
NAND_3395: ENTITY WORK.NAND
    PORT MAP (
        A => S5594,
        B => S5596,
        Y => S5597
    );
NOT_443: ENTITY WORK.NOT
    PORT MAP (
        A => S5597,
        Y => S5598
    );
NOR_1869: ENTITY WORK.NOR
    PORT MAP (
        A => S5404,
        B => S5405,
        Y => S5599
    );
NOR_1870: ENTITY WORK.NOR
    PORT MAP (
        A => S5507,
        B => S5599,
        Y => S5600
    );
NAND_3396: ENTITY WORK.NAND
    PORT MAP (
        A => S5507,
        B => S5599,
        Y => S5601
    );
NOT_444: ENTITY WORK.NOT
    PORT MAP (
        A => S5601,
        Y => S5602
    );
NOR_1871: ENTITY WORK.NOR
    PORT MAP (
        A => S5600,
        B => S5602,
        Y => S5603
    );
NOR_1872: ENTITY WORK.NOR
    PORT MAP (
        A => S5539,
        B => S5603,
        Y => S5604
    );
NOR_1873: ENTITY WORK.NOR
    PORT MAP (
        A => S5402,
        B => S5538,
        Y => S5605
    );
NOR_1874: ENTITY WORK.NOR
    PORT MAP (
        A => S5604,
        B => S5605,
        Y => S5606
    );
NOT_445: ENTITY WORK.NOT
    PORT MAP (
        A => S5606,
        Y => S5607
    );
NOR_1875: ENTITY WORK.NOR
    PORT MAP (
        A => S2417,
        B => S5607,
        Y => S5608
    );
NOR_1876: ENTITY WORK.NOR
    PORT MAP (
        A => S2418,
        B => S5606,
        Y => S5609
    );
NOR_1877: ENTITY WORK.NOR
    PORT MAP (
        A => S5499,
        B => S5502,
        Y => S5610
    );
NOT_446: ENTITY WORK.NOT
    PORT MAP (
        A => S5610,
        Y => S5611
    );
NAND_3397: ENTITY WORK.NAND
    PORT MAP (
        A => S5505,
        B => S5611,
        Y => S5612
    );
NAND_3398: ENTITY WORK.NAND
    PORT MAP (
        A => S5538,
        B => S5612,
        Y => S5613
    );
NAND_3399: ENTITY WORK.NAND
    PORT MAP (
        A => S5411,
        B => S5539,
        Y => S5614
    );
NAND_3400: ENTITY WORK.NAND
    PORT MAP (
        A => S5613,
        B => S5614,
        Y => S5615
    );
NOT_447: ENTITY WORK.NOT
    PORT MAP (
        A => S5615,
        Y => S5616
    );
NAND_3401: ENTITY WORK.NAND
    PORT MAP (
        A => S2312,
        B => S5616,
        Y => S5617
    );
NOT_448: ENTITY WORK.NOT
    PORT MAP (
        A => S5617,
        Y => S5618
    );
NAND_3402: ENTITY WORK.NAND
    PORT MAP (
        A => S2311,
        B => S5615,
        Y => S5619
    );
NAND_3403: ENTITY WORK.NAND
    PORT MAP (
        A => S5617,
        B => S5619,
        Y => S5620
    );
NOT_449: ENTITY WORK.NOT
    PORT MAP (
        A => S5620,
        Y => S5621
    );
NAND_3404: ENTITY WORK.NAND
    PORT MAP (
        A => S5424,
        B => S5494,
        Y => S5622
    );
NAND_3405: ENTITY WORK.NAND
    PORT MAP (
        A => S5497,
        B => S5622,
        Y => S5623
    );
NAND_3406: ENTITY WORK.NAND
    PORT MAP (
        A => S5538,
        B => S5623,
        Y => S5624
    );
NAND_3407: ENTITY WORK.NAND
    PORT MAP (
        A => S5419,
        B => S5539,
        Y => S5625
    );
NAND_3408: ENTITY WORK.NAND
    PORT MAP (
        A => S5624,
        B => S5625,
        Y => S5626
    );
NOT_450: ENTITY WORK.NOT
    PORT MAP (
        A => S5626,
        Y => S5627
    );
NOR_1878: ENTITY WORK.NOR
    PORT MAP (
        A => S2205,
        B => S5626,
        Y => S5628
    );
NOR_1879: ENTITY WORK.NOR
    PORT MAP (
        A => S2206,
        B => S5627,
        Y => S5629
    );
NAND_3409: ENTITY WORK.NAND
    PORT MAP (
        A => S5435,
        B => S5490,
        Y => S5630
    );
NAND_3410: ENTITY WORK.NAND
    PORT MAP (
        A => S5493,
        B => S5630,
        Y => S5631
    );
NAND_3411: ENTITY WORK.NAND
    PORT MAP (
        A => S5538,
        B => S5631,
        Y => S5632
    );
NAND_3412: ENTITY WORK.NAND
    PORT MAP (
        A => S5430,
        B => S5539,
        Y => S5633
    );
NAND_3413: ENTITY WORK.NAND
    PORT MAP (
        A => S5632,
        B => S5633,
        Y => S5634
    );
NOT_451: ENTITY WORK.NOT
    PORT MAP (
        A => S5634,
        Y => S5635
    );
NAND_3414: ENTITY WORK.NAND
    PORT MAP (
        A => S2107,
        B => S5635,
        Y => S5636
    );
NOT_452: ENTITY WORK.NOT
    PORT MAP (
        A => S5636,
        Y => S5637
    );
NAND_3415: ENTITY WORK.NAND
    PORT MAP (
        A => S2106,
        B => S5634,
        Y => S5638
    );
NAND_3416: ENTITY WORK.NAND
    PORT MAP (
        A => S5636,
        B => S5638,
        Y => S5639
    );
NOT_453: ENTITY WORK.NOT
    PORT MAP (
        A => S5639,
        Y => S5640
    );
NOR_1880: ENTITY WORK.NOR
    PORT MAP (
        A => S5446,
        B => S5448,
        Y => S5641
    );
NAND_3417: ENTITY WORK.NAND
    PORT MAP (
        A => S5447,
        B => S5449,
        Y => S5642
    );
NOR_1881: ENTITY WORK.NOR
    PORT MAP (
        A => S5486,
        B => S5642,
        Y => S5643
    );
NOR_1882: ENTITY WORK.NOR
    PORT MAP (
        A => S5487,
        B => S5641,
        Y => S5644
    );
NOR_1883: ENTITY WORK.NOR
    PORT MAP (
        A => S5643,
        B => S5644,
        Y => S5645
    );
NAND_3418: ENTITY WORK.NAND
    PORT MAP (
        A => S5538,
        B => S5645,
        Y => S5646
    );
NAND_3419: ENTITY WORK.NAND
    PORT MAP (
        A => S5444,
        B => S5539,
        Y => S5647
    );
NAND_3420: ENTITY WORK.NAND
    PORT MAP (
        A => S5646,
        B => S5647,
        Y => S5648
    );
NOT_454: ENTITY WORK.NOT
    PORT MAP (
        A => S5648,
        Y => S5649
    );
NOR_1884: ENTITY WORK.NOR
    PORT MAP (
        A => S1597,
        B => S5649,
        Y => S5650
    );
NAND_3421: ENTITY WORK.NAND
    PORT MAP (
        A => S1598,
        B => S5648,
        Y => S5651
    );
NOR_1885: ENTITY WORK.NOR
    PORT MAP (
        A => S1598,
        B => S5648,
        Y => S5652
    );
NAND_3422: ENTITY WORK.NAND
    PORT MAP (
        A => S1597,
        B => S5649,
        Y => S5653
    );
NOR_1886: ENTITY WORK.NOR
    PORT MAP (
        A => S5462,
        B => S5483,
        Y => S5654
    );
NAND_3423: ENTITY WORK.NAND
    PORT MAP (
        A => S5463,
        B => S5482,
        Y => S5655
    );
NOR_1887: ENTITY WORK.NOR
    PORT MAP (
        A => S5484,
        B => S5654,
        Y => S5656
    );
NAND_3424: ENTITY WORK.NAND
    PORT MAP (
        A => S5485,
        B => S5655,
        Y => S5657
    );
NOR_1888: ENTITY WORK.NOR
    PORT MAP (
        A => S5539,
        B => S5656,
        Y => S5658
    );
NAND_3425: ENTITY WORK.NAND
    PORT MAP (
        A => S5538,
        B => S5657,
        Y => S5659
    );
NOR_1889: ENTITY WORK.NOR
    PORT MAP (
        A => S5457,
        B => S5538,
        Y => S5660
    );
NAND_3426: ENTITY WORK.NAND
    PORT MAP (
        A => S5456,
        B => S5539,
        Y => S5661
    );
NOR_1890: ENTITY WORK.NOR
    PORT MAP (
        A => S5658,
        B => S5660,
        Y => S5662
    );
NAND_3427: ENTITY WORK.NAND
    PORT MAP (
        A => S5659,
        B => S5661,
        Y => S5663
    );
NOR_1891: ENTITY WORK.NOR
    PORT MAP (
        A => S1952,
        B => S5663,
        Y => S5664
    );
NAND_3428: ENTITY WORK.NAND
    PORT MAP (
        A => S1953,
        B => S5662,
        Y => S5665
    );
NOR_1892: ENTITY WORK.NOR
    PORT MAP (
        A => S1953,
        B => S5662,
        Y => S5666
    );
NAND_3429: ENTITY WORK.NAND
    PORT MAP (
        A => S1952,
        B => S5663,
        Y => S5667
    );
NOR_1893: ENTITY WORK.NOR
    PORT MAP (
        A => S5664,
        B => S5666,
        Y => S5668
    );
NAND_3430: ENTITY WORK.NAND
    PORT MAP (
        A => S5665,
        B => S5667,
        Y => S5669
    );
NOR_1894: ENTITY WORK.NOR
    PORT MAP (
        A => S5475,
        B => S5478,
        Y => S5670
    );
NAND_3431: ENTITY WORK.NAND
    PORT MAP (
        A => S5474,
        B => S5479,
        Y => S5671
    );
NOR_1895: ENTITY WORK.NOR
    PORT MAP (
        A => S5480,
        B => S5670,
        Y => S5672
    );
NAND_3432: ENTITY WORK.NAND
    PORT MAP (
        A => S5481,
        B => S5671,
        Y => S5673
    );
NOR_1896: ENTITY WORK.NOR
    PORT MAP (
        A => S5539,
        B => S5672,
        Y => S5674
    );
NAND_3433: ENTITY WORK.NAND
    PORT MAP (
        A => S5538,
        B => S5673,
        Y => S5675
    );
NOR_1897: ENTITY WORK.NOR
    PORT MAP (
        A => S5471,
        B => S5538,
        Y => S5676
    );
NAND_3434: ENTITY WORK.NAND
    PORT MAP (
        A => S5470,
        B => S5539,
        Y => S5677
    );
NOR_1898: ENTITY WORK.NOR
    PORT MAP (
        A => S5674,
        B => S5676,
        Y => S5678
    );
NAND_3435: ENTITY WORK.NAND
    PORT MAP (
        A => S5675,
        B => S5677,
        Y => S5679
    );
NOR_1899: ENTITY WORK.NOR
    PORT MAP (
        A => S1848,
        B => S5679,
        Y => S5680
    );
NAND_3436: ENTITY WORK.NAND
    PORT MAP (
        A => S1849,
        B => S5678,
        Y => S5681
    );
NOR_1900: ENTITY WORK.NOR
    PORT MAP (
        A => S1849,
        B => S5678,
        Y => S5682
    );
NAND_3437: ENTITY WORK.NAND
    PORT MAP (
        A => S1848,
        B => S5679,
        Y => S5683
    );
NOR_1901: ENTITY WORK.NOR
    PORT MAP (
        A => S1516,
        B => S5539,
        Y => S5684
    );
NAND_3438: ENTITY WORK.NAND
    PORT MAP (
        A => S1515,
        B => S5538,
        Y => S5685
    );
NOR_1902: ENTITY WORK.NOR
    PORT MAP (
        A => S1116,
        B => S5684,
        Y => S5686
    );
NAND_3439: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_2,
        B => S5685,
        Y => S5687
    );
NOR_1903: ENTITY WORK.NOR
    PORT MAP (
        A => S5475,
        B => S5539,
        Y => S5688
    );
NAND_3440: ENTITY WORK.NAND
    PORT MAP (
        A => S5474,
        B => S5538,
        Y => S5689
    );
NOR_1904: ENTITY WORK.NOR
    PORT MAP (
        A => S5686,
        B => S5688,
        Y => S5690
    );
NAND_3441: ENTITY WORK.NAND
    PORT MAP (
        A => S5687,
        B => S5689,
        Y => S5691
    );
NOR_1905: ENTITY WORK.NOR
    PORT MAP (
        A => S1745,
        B => S5690,
        Y => S5692
    );
NAND_3442: ENTITY WORK.NAND
    PORT MAP (
        A => S1746,
        B => S5691,
        Y => S5693
    );
NOR_1906: ENTITY WORK.NOR
    PORT MAP (
        A => S1746,
        B => S5691,
        Y => S5694
    );
NAND_3443: ENTITY WORK.NAND
    PORT MAP (
        A => S1745,
        B => S5690,
        Y => S5695
    );
NOR_1907: ENTITY WORK.NOR
    PORT MAP (
        A => S5692,
        B => S5694,
        Y => S5696
    );
NAND_3444: ENTITY WORK.NAND
    PORT MAP (
        A => S5693,
        B => S5695,
        Y => S5697
    );
NAND_3445: ENTITY WORK.NAND
    PORT MAP (
        A => S1168,
        B => S1515,
        Y => S5698
    );
NOT_455: ENTITY WORK.NOT
    PORT MAP (
        A => S5698,
        Y => S5699
    );
NOR_1908: ENTITY WORK.NOR
    PORT MAP (
        A => S5697,
        B => S5699,
        Y => S5700
    );
NAND_3446: ENTITY WORK.NAND
    PORT MAP (
        A => S5696,
        B => S5698,
        Y => S5701
    );
NOR_1909: ENTITY WORK.NOR
    PORT MAP (
        A => S5692,
        B => S5700,
        Y => S5702
    );
NAND_3447: ENTITY WORK.NAND
    PORT MAP (
        A => S5693,
        B => S5701,
        Y => S5703
    );
NOR_1910: ENTITY WORK.NOR
    PORT MAP (
        A => S5682,
        B => S5702,
        Y => S5704
    );
NAND_3448: ENTITY WORK.NAND
    PORT MAP (
        A => S5683,
        B => S5703,
        Y => S5705
    );
NOR_1911: ENTITY WORK.NOR
    PORT MAP (
        A => S5680,
        B => S5704,
        Y => S5706
    );
NAND_3449: ENTITY WORK.NAND
    PORT MAP (
        A => S5681,
        B => S5705,
        Y => S5707
    );
NOR_1912: ENTITY WORK.NOR
    PORT MAP (
        A => S5669,
        B => S5706,
        Y => S5708
    );
NAND_3450: ENTITY WORK.NAND
    PORT MAP (
        A => S5668,
        B => S5707,
        Y => S5709
    );
NOR_1913: ENTITY WORK.NOR
    PORT MAP (
        A => S5664,
        B => S5708,
        Y => S5710
    );
NAND_3451: ENTITY WORK.NAND
    PORT MAP (
        A => S5665,
        B => S5709,
        Y => S5711
    );
NOR_1914: ENTITY WORK.NOR
    PORT MAP (
        A => S5652,
        B => S5710,
        Y => S5712
    );
NAND_3452: ENTITY WORK.NAND
    PORT MAP (
        A => S5653,
        B => S5711,
        Y => S5713
    );
NOR_1915: ENTITY WORK.NOR
    PORT MAP (
        A => S5650,
        B => S5712,
        Y => S5714
    );
NAND_3453: ENTITY WORK.NAND
    PORT MAP (
        A => S5651,
        B => S5713,
        Y => S5715
    );
NOR_1916: ENTITY WORK.NOR
    PORT MAP (
        A => S5639,
        B => S5714,
        Y => S5716
    );
NAND_3454: ENTITY WORK.NAND
    PORT MAP (
        A => S5640,
        B => S5715,
        Y => S5717
    );
NOR_1917: ENTITY WORK.NOR
    PORT MAP (
        A => S5637,
        B => S5716,
        Y => S5718
    );
NAND_3455: ENTITY WORK.NAND
    PORT MAP (
        A => S5636,
        B => S5717,
        Y => S5719
    );
NOR_1918: ENTITY WORK.NOR
    PORT MAP (
        A => S5629,
        B => S5718,
        Y => S5720
    );
NOR_1919: ENTITY WORK.NOR
    PORT MAP (
        A => S5628,
        B => S5719,
        Y => S5721
    );
NOR_1920: ENTITY WORK.NOR
    PORT MAP (
        A => S5628,
        B => S5720,
        Y => S5722
    );
NOR_1921: ENTITY WORK.NOR
    PORT MAP (
        A => S5629,
        B => S5721,
        Y => S5723
    );
NOR_1922: ENTITY WORK.NOR
    PORT MAP (
        A => S5620,
        B => S5722,
        Y => S5724
    );
NAND_3456: ENTITY WORK.NAND
    PORT MAP (
        A => S5621,
        B => S5723,
        Y => S5725
    );
NOR_1923: ENTITY WORK.NOR
    PORT MAP (
        A => S5618,
        B => S5724,
        Y => S5726
    );
NAND_3457: ENTITY WORK.NAND
    PORT MAP (
        A => S5617,
        B => S5725,
        Y => S5727
    );
NOR_1924: ENTITY WORK.NOR
    PORT MAP (
        A => S5609,
        B => S5726,
        Y => S5728
    );
NOR_1925: ENTITY WORK.NOR
    PORT MAP (
        A => S5608,
        B => S5727,
        Y => S5729
    );
NOR_1926: ENTITY WORK.NOR
    PORT MAP (
        A => S5608,
        B => S5728,
        Y => S5730
    );
NOR_1927: ENTITY WORK.NOR
    PORT MAP (
        A => S5609,
        B => S5729,
        Y => S5731
    );
NOR_1928: ENTITY WORK.NOR
    PORT MAP (
        A => S5597,
        B => S5730,
        Y => S5732
    );
NAND_3458: ENTITY WORK.NAND
    PORT MAP (
        A => S5598,
        B => S5731,
        Y => S5733
    );
NOR_1929: ENTITY WORK.NOR
    PORT MAP (
        A => S5595,
        B => S5732,
        Y => S5734
    );
NAND_3459: ENTITY WORK.NAND
    PORT MAP (
        A => S5594,
        B => S5733,
        Y => S5735
    );
NAND_3460: ENTITY WORK.NAND
    PORT MAP (
        A => S5587,
        B => S5735,
        Y => S5736
    );
NAND_3461: ENTITY WORK.NAND
    PORT MAP (
        A => S5586,
        B => S5734,
        Y => S5737
    );
NAND_3462: ENTITY WORK.NAND
    PORT MAP (
        A => S5587,
        B => S5737,
        Y => S5738
    );
NAND_3463: ENTITY WORK.NAND
    PORT MAP (
        A => S5586,
        B => S5736,
        Y => S5739
    );
NOR_1930: ENTITY WORK.NOR
    PORT MAP (
        A => S5572,
        B => S5738,
        Y => S5740
    );
NAND_3464: ENTITY WORK.NAND
    PORT MAP (
        A => S5571,
        B => S5739,
        Y => S5741
    );
NOR_1931: ENTITY WORK.NOR
    PORT MAP (
        A => S5568,
        B => S5740,
        Y => S5742
    );
NAND_3465: ENTITY WORK.NAND
    PORT MAP (
        A => S5569,
        B => S5741,
        Y => S5743
    );
NAND_3466: ENTITY WORK.NAND
    PORT MAP (
        A => S5561,
        B => S5743,
        Y => S5744
    );
NAND_3467: ENTITY WORK.NAND
    PORT MAP (
        A => S5560,
        B => S5742,
        Y => S5745
    );
NAND_3468: ENTITY WORK.NAND
    PORT MAP (
        A => S5561,
        B => S5745,
        Y => S5746
    );
NAND_3469: ENTITY WORK.NAND
    PORT MAP (
        A => S5560,
        B => S5744,
        Y => S5747
    );
NOR_1932: ENTITY WORK.NOR
    PORT MAP (
        A => S5549,
        B => S5746,
        Y => S5748
    );
NAND_3470: ENTITY WORK.NAND
    PORT MAP (
        A => S5550,
        B => S5747,
        Y => S5749
    );
NAND_3471: ENTITY WORK.NAND
    PORT MAP (
        A => S5334,
        B => S5539,
        Y => S5750
    );
NOT_456: ENTITY WORK.NOT
    PORT MAP (
        A => S5750,
        Y => S5751
    );
NOR_1933: ENTITY WORK.NOR
    PORT MAP (
        A => S3950,
        B => S5751,
        Y => S5752
    );
NOR_1934: ENTITY WORK.NOR
    PORT MAP (
        A => S3036,
        B => S5752,
        Y => S5753
    );
NOT_457: ENTITY WORK.NOT
    PORT MAP (
        A => S5753,
        Y => S5754
    );
NOR_1935: ENTITY WORK.NOR
    PORT MAP (
        A => S5547,
        B => S5753,
        Y => S5755
    );
NAND_3472: ENTITY WORK.NAND
    PORT MAP (
        A => S5546,
        B => S5754,
        Y => S5756
    );
NOR_1936: ENTITY WORK.NOR
    PORT MAP (
        A => S5748,
        B => S5756,
        Y => S5757
    );
NAND_3473: ENTITY WORK.NAND
    PORT MAP (
        A => S5749,
        B => S5755,
        Y => S5758
    );
NAND_3474: ENTITY WORK.NAND
    PORT MAP (
        A => S3036,
        B => S5752,
        Y => S5759
    );
NAND_3475: ENTITY WORK.NAND
    PORT MAP (
        A => S3142,
        B => S5759,
        Y => S5760
    );
NOT_458: ENTITY WORK.NOT
    PORT MAP (
        A => S5760,
        Y => S5761
    );
NOR_1937: ENTITY WORK.NOR
    PORT MAP (
        A => S5757,
        B => S5760,
        Y => S5762
    );
NAND_3476: ENTITY WORK.NAND
    PORT MAP (
        A => S5758,
        B => S5761,
        Y => S5763
    );
NAND_3477: ENTITY WORK.NAND
    PORT MAP (
        A => S5639,
        B => S5714,
        Y => S5764
    );
NAND_3478: ENTITY WORK.NAND
    PORT MAP (
        A => S5717,
        B => S5764,
        Y => S5765
    );
NAND_3479: ENTITY WORK.NAND
    PORT MAP (
        A => S5762,
        B => S5765,
        Y => S5766
    );
NAND_3480: ENTITY WORK.NAND
    PORT MAP (
        A => S5634,
        B => S5763,
        Y => S5767
    );
NAND_3481: ENTITY WORK.NAND
    PORT MAP (
        A => S5766,
        B => S5767,
        Y => S5768
    );
NAND_3482: ENTITY WORK.NAND
    PORT MAP (
        A => S2205,
        B => S5768,
        Y => S5769
    );
NOR_1938: ENTITY WORK.NOR
    PORT MAP (
        A => S5650,
        B => S5652,
        Y => S5770
    );
NAND_3483: ENTITY WORK.NAND
    PORT MAP (
        A => S5651,
        B => S5653,
        Y => S5771
    );
NOR_1939: ENTITY WORK.NOR
    PORT MAP (
        A => S5710,
        B => S5771,
        Y => S5772
    );
NOR_1940: ENTITY WORK.NOR
    PORT MAP (
        A => S5711,
        B => S5770,
        Y => S5773
    );
NOR_1941: ENTITY WORK.NOR
    PORT MAP (
        A => S5772,
        B => S5773,
        Y => S5774
    );
NAND_3484: ENTITY WORK.NAND
    PORT MAP (
        A => S5762,
        B => S5774,
        Y => S5775
    );
NAND_3485: ENTITY WORK.NAND
    PORT MAP (
        A => S5648,
        B => S5763,
        Y => S5776
    );
NAND_3486: ENTITY WORK.NAND
    PORT MAP (
        A => S5775,
        B => S5776,
        Y => S5777
    );
NAND_3487: ENTITY WORK.NAND
    PORT MAP (
        A => S2107,
        B => S5777,
        Y => S5778
    );
NOR_1942: ENTITY WORK.NOR
    PORT MAP (
        A => S5696,
        B => S5698,
        Y => S5779
    );
NOR_1943: ENTITY WORK.NOR
    PORT MAP (
        A => S5700,
        B => S5779,
        Y => S5780
    );
NOR_1944: ENTITY WORK.NOR
    PORT MAP (
        A => S5763,
        B => S5780,
        Y => S5781
    );
NOR_1945: ENTITY WORK.NOR
    PORT MAP (
        A => S5691,
        B => S5762,
        Y => S5782
    );
NOR_1946: ENTITY WORK.NOR
    PORT MAP (
        A => S5781,
        B => S5782,
        Y => S5783
    );
NAND_3488: ENTITY WORK.NAND
    PORT MAP (
        A => S1849,
        B => S5783,
        Y => S5784
    );
NAND_3489: ENTITY WORK.NAND
    PORT MAP (
        A => S1515,
        B => S5762,
        Y => S5785
    );
NAND_3490: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_1,
        B => S5785,
        Y => S5786
    );
NOR_1947: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_0,
        B => S1516,
        Y => S5787
    );
NOR_1948: ENTITY WORK.NOR
    PORT MAP (
        A => S1745,
        B => S5787,
        Y => S5788
    );
NOR_1949: ENTITY WORK.NOR
    PORT MAP (
        A => S5698,
        B => S5763,
        Y => S5789
    );
NOR_1950: ENTITY WORK.NOR
    PORT MAP (
        A => S5788,
        B => S5789,
        Y => S5790
    );
NAND_3491: ENTITY WORK.NAND
    PORT MAP (
        A => S5786,
        B => S5790,
        Y => S5791
    );
NAND_3492: ENTITY WORK.NAND
    PORT MAP (
        A => S1745,
        B => S5787,
        Y => S5792
    );
NAND_3493: ENTITY WORK.NAND
    PORT MAP (
        A => S5791,
        B => S5792,
        Y => S5793
    );
NAND_3494: ENTITY WORK.NAND
    PORT MAP (
        A => S5784,
        B => S5793,
        Y => S5794
    );
NOR_1951: ENTITY WORK.NOR
    PORT MAP (
        A => S5680,
        B => S5682,
        Y => S5795
    );
NAND_3495: ENTITY WORK.NAND
    PORT MAP (
        A => S5681,
        B => S5683,
        Y => S5796
    );
NAND_3496: ENTITY WORK.NAND
    PORT MAP (
        A => S5702,
        B => S5795,
        Y => S5797
    );
NAND_3497: ENTITY WORK.NAND
    PORT MAP (
        A => S5703,
        B => S5796,
        Y => S5798
    );
NAND_3498: ENTITY WORK.NAND
    PORT MAP (
        A => S5797,
        B => S5798,
        Y => S5799
    );
NAND_3499: ENTITY WORK.NAND
    PORT MAP (
        A => S5762,
        B => S5799,
        Y => S5800
    );
NOT_459: ENTITY WORK.NOT
    PORT MAP (
        A => S5800,
        Y => S5801
    );
NOR_1952: ENTITY WORK.NOR
    PORT MAP (
        A => S5679,
        B => S5762,
        Y => S5802
    );
NAND_3500: ENTITY WORK.NAND
    PORT MAP (
        A => S5678,
        B => S5763,
        Y => S5803
    );
NOR_1953: ENTITY WORK.NOR
    PORT MAP (
        A => S5801,
        B => S5802,
        Y => S5804
    );
NAND_3501: ENTITY WORK.NAND
    PORT MAP (
        A => S5800,
        B => S5803,
        Y => S5805
    );
NOR_1954: ENTITY WORK.NOR
    PORT MAP (
        A => S1953,
        B => S5805,
        Y => S5806
    );
NOR_1955: ENTITY WORK.NOR
    PORT MAP (
        A => S1849,
        B => S5783,
        Y => S5807
    );
NOR_1956: ENTITY WORK.NOR
    PORT MAP (
        A => S5806,
        B => S5807,
        Y => S5808
    );
NAND_3502: ENTITY WORK.NAND
    PORT MAP (
        A => S5794,
        B => S5808,
        Y => S5809
    );
NOR_1957: ENTITY WORK.NOR
    PORT MAP (
        A => S1952,
        B => S5804,
        Y => S5810
    );
NAND_3503: ENTITY WORK.NAND
    PORT MAP (
        A => S5669,
        B => S5706,
        Y => S5811
    );
NAND_3504: ENTITY WORK.NAND
    PORT MAP (
        A => S5709,
        B => S5811,
        Y => S5812
    );
NAND_3505: ENTITY WORK.NAND
    PORT MAP (
        A => S5762,
        B => S5812,
        Y => S5813
    );
NOT_460: ENTITY WORK.NOT
    PORT MAP (
        A => S5813,
        Y => S5814
    );
NOR_1958: ENTITY WORK.NOR
    PORT MAP (
        A => S5662,
        B => S5762,
        Y => S5815
    );
NOT_461: ENTITY WORK.NOT
    PORT MAP (
        A => S5815,
        Y => S5816
    );
NOR_1959: ENTITY WORK.NOR
    PORT MAP (
        A => S5814,
        B => S5815,
        Y => S5817
    );
NAND_3506: ENTITY WORK.NAND
    PORT MAP (
        A => S5813,
        B => S5816,
        Y => S5818
    );
NOR_1960: ENTITY WORK.NOR
    PORT MAP (
        A => S1597,
        B => S5818,
        Y => S5819
    );
NOR_1961: ENTITY WORK.NOR
    PORT MAP (
        A => S5810,
        B => S5819,
        Y => S5820
    );
NAND_3507: ENTITY WORK.NAND
    PORT MAP (
        A => S5809,
        B => S5820,
        Y => S5821
    );
NOR_1962: ENTITY WORK.NOR
    PORT MAP (
        A => S2107,
        B => S5777,
        Y => S5822
    );
NOR_1963: ENTITY WORK.NOR
    PORT MAP (
        A => S1598,
        B => S5817,
        Y => S5823
    );
NOR_1964: ENTITY WORK.NOR
    PORT MAP (
        A => S5822,
        B => S5823,
        Y => S5824
    );
NAND_3508: ENTITY WORK.NAND
    PORT MAP (
        A => S5821,
        B => S5824,
        Y => S5825
    );
NAND_3509: ENTITY WORK.NAND
    PORT MAP (
        A => S5778,
        B => S5825,
        Y => S5826
    );
NAND_3510: ENTITY WORK.NAND
    PORT MAP (
        A => S5769,
        B => S5826,
        Y => S5827
    );
NOR_1965: ENTITY WORK.NOR
    PORT MAP (
        A => S5628,
        B => S5629,
        Y => S5828
    );
NOR_1966: ENTITY WORK.NOR
    PORT MAP (
        A => S5719,
        B => S5828,
        Y => S5829
    );
NAND_3511: ENTITY WORK.NAND
    PORT MAP (
        A => S5719,
        B => S5828,
        Y => S5830
    );
NOT_462: ENTITY WORK.NOT
    PORT MAP (
        A => S5830,
        Y => S5831
    );
NOR_1967: ENTITY WORK.NOR
    PORT MAP (
        A => S5829,
        B => S5831,
        Y => S5832
    );
NOR_1968: ENTITY WORK.NOR
    PORT MAP (
        A => S5626,
        B => S5762,
        Y => S5833
    );
NAND_3512: ENTITY WORK.NAND
    PORT MAP (
        A => S5762,
        B => S5832,
        Y => S5834
    );
NOT_463: ENTITY WORK.NOT
    PORT MAP (
        A => S5834,
        Y => S5835
    );
NOR_1969: ENTITY WORK.NOR
    PORT MAP (
        A => S5833,
        B => S5835,
        Y => S5836
    );
NOR_1970: ENTITY WORK.NOR
    PORT MAP (
        A => S2311,
        B => S5836,
        Y => S5837
    );
NOR_1971: ENTITY WORK.NOR
    PORT MAP (
        A => S2205,
        B => S5768,
        Y => S5838
    );
NOR_1972: ENTITY WORK.NOR
    PORT MAP (
        A => S5837,
        B => S5838,
        Y => S5839
    );
NAND_3513: ENTITY WORK.NAND
    PORT MAP (
        A => S5827,
        B => S5839,
        Y => S5840
    );
NAND_3514: ENTITY WORK.NAND
    PORT MAP (
        A => S5597,
        B => S5730,
        Y => S5841
    );
NAND_3515: ENTITY WORK.NAND
    PORT MAP (
        A => S5733,
        B => S5841,
        Y => S5842
    );
NAND_3516: ENTITY WORK.NAND
    PORT MAP (
        A => S5762,
        B => S5842,
        Y => S5843
    );
NAND_3517: ENTITY WORK.NAND
    PORT MAP (
        A => S5592,
        B => S5763,
        Y => S5844
    );
NAND_3518: ENTITY WORK.NAND
    PORT MAP (
        A => S5843,
        B => S5844,
        Y => S5845
    );
NOR_1973: ENTITY WORK.NOR
    PORT MAP (
        A => S2617,
        B => S5845,
        Y => S5846
    );
NAND_3519: ENTITY WORK.NAND
    PORT MAP (
        A => S5586,
        B => S5587,
        Y => S5847
    );
NAND_3520: ENTITY WORK.NAND
    PORT MAP (
        A => S5735,
        B => S5847,
        Y => S5848
    );
NOT_464: ENTITY WORK.NOT
    PORT MAP (
        A => S5848,
        Y => S5849
    );
NOR_1974: ENTITY WORK.NOR
    PORT MAP (
        A => S5735,
        B => S5847,
        Y => S5850
    );
NOR_1975: ENTITY WORK.NOR
    PORT MAP (
        A => S5849,
        B => S5850,
        Y => S5851
    );
NAND_3521: ENTITY WORK.NAND
    PORT MAP (
        A => S5762,
        B => S5851,
        Y => S5852
    );
NOT_465: ENTITY WORK.NOT
    PORT MAP (
        A => S5852,
        Y => S5853
    );
NOR_1976: ENTITY WORK.NOR
    PORT MAP (
        A => S5584,
        B => S5762,
        Y => S5854
    );
NOT_466: ENTITY WORK.NOT
    PORT MAP (
        A => S5854,
        Y => S5855
    );
NOR_1977: ENTITY WORK.NOR
    PORT MAP (
        A => S5853,
        B => S5854,
        Y => S5856
    );
NAND_3522: ENTITY WORK.NAND
    PORT MAP (
        A => S5852,
        B => S5855,
        Y => S5857
    );
NOR_1978: ENTITY WORK.NOR
    PORT MAP (
        A => S2717,
        B => S5857,
        Y => S5858
    );
NOR_1979: ENTITY WORK.NOR
    PORT MAP (
        A => S5846,
        B => S5858,
        Y => S5859
    );
NOT_467: ENTITY WORK.NOT
    PORT MAP (
        A => S5859,
        Y => S5860
    );
NAND_3523: ENTITY WORK.NAND
    PORT MAP (
        A => S2617,
        B => S5845,
        Y => S5861
    );
NOR_1980: ENTITY WORK.NOR
    PORT MAP (
        A => S2718,
        B => S5856,
        Y => S5862
    );
NAND_3524: ENTITY WORK.NAND
    PORT MAP (
        A => S2717,
        B => S5857,
        Y => S5863
    );
NAND_3525: ENTITY WORK.NAND
    PORT MAP (
        A => S5861,
        B => S5863,
        Y => S5864
    );
NOR_1981: ENTITY WORK.NOR
    PORT MAP (
        A => S5860,
        B => S5864,
        Y => S5865
    );
NAND_3526: ENTITY WORK.NAND
    PORT MAP (
        A => S5620,
        B => S5722,
        Y => S5866
    );
NAND_3527: ENTITY WORK.NAND
    PORT MAP (
        A => S5725,
        B => S5866,
        Y => S5867
    );
NAND_3528: ENTITY WORK.NAND
    PORT MAP (
        A => S5762,
        B => S5867,
        Y => S5868
    );
NAND_3529: ENTITY WORK.NAND
    PORT MAP (
        A => S5615,
        B => S5763,
        Y => S5869
    );
NAND_3530: ENTITY WORK.NAND
    PORT MAP (
        A => S5868,
        B => S5869,
        Y => S5870
    );
NOT_468: ENTITY WORK.NOT
    PORT MAP (
        A => S5870,
        Y => S5871
    );
NOR_1982: ENTITY WORK.NOR
    PORT MAP (
        A => S2417,
        B => S5870,
        Y => S5872
    );
NAND_3531: ENTITY WORK.NAND
    PORT MAP (
        A => S2418,
        B => S5871,
        Y => S5873
    );
NAND_3532: ENTITY WORK.NAND
    PORT MAP (
        A => S2311,
        B => S5836,
        Y => S5874
    );
NOR_1983: ENTITY WORK.NOR
    PORT MAP (
        A => S5608,
        B => S5609,
        Y => S5875
    );
NOR_1984: ENTITY WORK.NOR
    PORT MAP (
        A => S5727,
        B => S5875,
        Y => S5876
    );
NOT_469: ENTITY WORK.NOT
    PORT MAP (
        A => S5876,
        Y => S5877
    );
NAND_3533: ENTITY WORK.NAND
    PORT MAP (
        A => S5727,
        B => S5875,
        Y => S5878
    );
NAND_3534: ENTITY WORK.NAND
    PORT MAP (
        A => S5877,
        B => S5878,
        Y => S5879
    );
NAND_3535: ENTITY WORK.NAND
    PORT MAP (
        A => S5762,
        B => S5879,
        Y => S5880
    );
NOT_470: ENTITY WORK.NOT
    PORT MAP (
        A => S5880,
        Y => S5881
    );
NOR_1985: ENTITY WORK.NOR
    PORT MAP (
        A => S5606,
        B => S5762,
        Y => S5882
    );
NOR_1986: ENTITY WORK.NOR
    PORT MAP (
        A => S5881,
        B => S5882,
        Y => S5883
    );
NOT_471: ENTITY WORK.NOT
    PORT MAP (
        A => S5883,
        Y => S5884
    );
NAND_3536: ENTITY WORK.NAND
    PORT MAP (
        A => S2518,
        B => S5883,
        Y => S5885
    );
NOR_1987: ENTITY WORK.NOR
    PORT MAP (
        A => S2518,
        B => S5883,
        Y => S5886
    );
NAND_3537: ENTITY WORK.NAND
    PORT MAP (
        A => S2517,
        B => S5884,
        Y => S5887
    );
NAND_3538: ENTITY WORK.NAND
    PORT MAP (
        A => S2417,
        B => S5870,
        Y => S5888
    );
NAND_3539: ENTITY WORK.NAND
    PORT MAP (
        A => S5874,
        B => S5887,
        Y => S5889
    );
NAND_3540: ENTITY WORK.NAND
    PORT MAP (
        A => S5885,
        B => S5888,
        Y => S5890
    );
NOR_1988: ENTITY WORK.NOR
    PORT MAP (
        A => S5889,
        B => S5890,
        Y => S5891
    );
NAND_3541: ENTITY WORK.NAND
    PORT MAP (
        A => S5865,
        B => S5891,
        Y => S5892
    );
NOR_1989: ENTITY WORK.NOR
    PORT MAP (
        A => S5872,
        B => S5892,
        Y => S5893
    );
NAND_3542: ENTITY WORK.NAND
    PORT MAP (
        A => S5840,
        B => S5893,
        Y => S5894
    );
NAND_3543: ENTITY WORK.NAND
    PORT MAP (
        A => S5873,
        B => S5885,
        Y => S5895
    );
NAND_3544: ENTITY WORK.NAND
    PORT MAP (
        A => S5865,
        B => S5895,
        Y => S5896
    );
NOR_1990: ENTITY WORK.NOR
    PORT MAP (
        A => S5886,
        B => S5896,
        Y => S5897
    );
NOR_1991: ENTITY WORK.NOR
    PORT MAP (
        A => S5859,
        B => S5862,
        Y => S5898
    );
NOR_1992: ENTITY WORK.NOR
    PORT MAP (
        A => S5897,
        B => S5898,
        Y => S5899
    );
NAND_3545: ENTITY WORK.NAND
    PORT MAP (
        A => S5894,
        B => S5899,
        Y => S5900
    );
NOR_1993: ENTITY WORK.NOR
    PORT MAP (
        A => S5752,
        B => S5762,
        Y => S5901
    );
NOT_472: ENTITY WORK.NOT
    PORT MAP (
        A => S5901,
        Y => S5902
    );
NAND_3546: ENTITY WORK.NAND
    PORT MAP (
        A => S5121,
        B => S5902,
        Y => S5903
    );
NAND_3547: ENTITY WORK.NAND
    PORT MAP (
        A => S3142,
        B => S5903,
        Y => S5904
    );
NAND_3548: ENTITY WORK.NAND
    PORT MAP (
        A => S5549,
        B => S5746,
        Y => S5905
    );
NAND_3549: ENTITY WORK.NAND
    PORT MAP (
        A => S5749,
        B => S5905,
        Y => S5906
    );
NAND_3550: ENTITY WORK.NAND
    PORT MAP (
        A => S5762,
        B => S5906,
        Y => S5907
    );
NAND_3551: ENTITY WORK.NAND
    PORT MAP (
        A => S5544,
        B => S5763,
        Y => S5908
    );
NAND_3552: ENTITY WORK.NAND
    PORT MAP (
        A => S5907,
        B => S5908,
        Y => S5909
    );
NOR_1994: ENTITY WORK.NOR
    PORT MAP (
        A => S3036,
        B => S5909,
        Y => S5910
    );
NOT_473: ENTITY WORK.NOT
    PORT MAP (
        A => S5910,
        Y => S5911
    );
NAND_3553: ENTITY WORK.NAND
    PORT MAP (
        A => S5904,
        B => S5911,
        Y => S5912
    );
NOR_1995: ENTITY WORK.NOR
    PORT MAP (
        A => S3142,
        B => S5903,
        Y => S5913
    );
NOT_474: ENTITY WORK.NOT
    PORT MAP (
        A => S5913,
        Y => S5914
    );
NAND_3554: ENTITY WORK.NAND
    PORT MAP (
        A => S3036,
        B => S5909,
        Y => S5915
    );
NAND_3555: ENTITY WORK.NAND
    PORT MAP (
        A => S5914,
        B => S5915,
        Y => S5916
    );
NOR_1996: ENTITY WORK.NOR
    PORT MAP (
        A => S5912,
        B => S5916,
        Y => S5917
    );
NOR_1997: ENTITY WORK.NOR
    PORT MAP (
        A => S5571,
        B => S5739,
        Y => S5918
    );
NOR_1998: ENTITY WORK.NOR
    PORT MAP (
        A => S5740,
        B => S5918,
        Y => S5919
    );
NOR_1999: ENTITY WORK.NOR
    PORT MAP (
        A => S5763,
        B => S5919,
        Y => S5920
    );
NOR_2000: ENTITY WORK.NOR
    PORT MAP (
        A => S5566,
        B => S5762,
        Y => S5921
    );
NOR_2001: ENTITY WORK.NOR
    PORT MAP (
        A => S5920,
        B => S5921,
        Y => S5922
    );
NAND_3556: ENTITY WORK.NAND
    PORT MAP (
        A => S2817,
        B => S5922,
        Y => S5923
    );
NAND_3557: ENTITY WORK.NAND
    PORT MAP (
        A => S5560,
        B => S5561,
        Y => S5924
    );
NAND_3558: ENTITY WORK.NAND
    PORT MAP (
        A => S5742,
        B => S5924,
        Y => S5925
    );
NOR_2002: ENTITY WORK.NOR
    PORT MAP (
        A => S5742,
        B => S5924,
        Y => S5926
    );
NOT_475: ENTITY WORK.NOT
    PORT MAP (
        A => S5926,
        Y => S5927
    );
NAND_3559: ENTITY WORK.NAND
    PORT MAP (
        A => S5925,
        B => S5927,
        Y => S5928
    );
NAND_3560: ENTITY WORK.NAND
    PORT MAP (
        A => S5762,
        B => S5928,
        Y => S5929
    );
NOT_476: ENTITY WORK.NOT
    PORT MAP (
        A => S5929,
        Y => S5930
    );
NOR_2003: ENTITY WORK.NOR
    PORT MAP (
        A => S5558,
        B => S5762,
        Y => S5931
    );
NOR_2004: ENTITY WORK.NOR
    PORT MAP (
        A => S5930,
        B => S5931,
        Y => S5932
    );
NAND_3561: ENTITY WORK.NAND
    PORT MAP (
        A => S2920,
        B => S5932,
        Y => S5933
    );
NAND_3562: ENTITY WORK.NAND
    PORT MAP (
        A => S5923,
        B => S5933,
        Y => S5934
    );
NOR_2005: ENTITY WORK.NOR
    PORT MAP (
        A => S2817,
        B => S5922,
        Y => S5935
    );
NOR_2006: ENTITY WORK.NOR
    PORT MAP (
        A => S2920,
        B => S5932,
        Y => S5936
    );
NOR_2007: ENTITY WORK.NOR
    PORT MAP (
        A => S5934,
        B => S5936,
        Y => S5937
    );
NAND_3563: ENTITY WORK.NAND
    PORT MAP (
        A => S5917,
        B => S5937,
        Y => S5938
    );
NOR_2008: ENTITY WORK.NOR
    PORT MAP (
        A => S5935,
        B => S5938,
        Y => S5939
    );
NAND_3564: ENTITY WORK.NAND
    PORT MAP (
        A => S5900,
        B => S5939,
        Y => S5940
    );
NAND_3565: ENTITY WORK.NAND
    PORT MAP (
        A => S5910,
        B => S5914,
        Y => S5941
    );
NAND_3566: ENTITY WORK.NAND
    PORT MAP (
        A => S5904,
        B => S5941,
        Y => S5942
    );
NAND_3567: ENTITY WORK.NAND
    PORT MAP (
        A => S5917,
        B => S5934,
        Y => S5943
    );
NOR_2009: ENTITY WORK.NOR
    PORT MAP (
        A => S5936,
        B => S5943,
        Y => S5944
    );
NOR_2010: ENTITY WORK.NOR
    PORT MAP (
        A => S5942,
        B => S5944,
        Y => S5945
    );
NAND_3568: ENTITY WORK.NAND
    PORT MAP (
        A => S5940,
        B => S5945,
        Y => S5946
    );
NAND_3569: ENTITY WORK.NAND
    PORT MAP (
        A => S3898,
        B => S5946,
        Y => S5947
    );
NOR_2011: ENTITY WORK.NOR
    PORT MAP (
        A => S377,
        B => S1392,
        Y => S5948
    );
NAND_3570: ENTITY WORK.NAND
    PORT MAP (
        A => S376,
        B => S1391,
        Y => S5949
    );
NAND_3571: ENTITY WORK.NAND
    PORT MAP (
        A => S8564,
        B => S376,
        Y => S5950
    );
NAND_3572: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu1_0,
        B => S5950,
        Y => S5951
    );
NOT_477: ENTITY WORK.NOT
    PORT MAP (
        A => S5951,
        Y => S5952
    );
NAND_3573: ENTITY WORK.NAND
    PORT MAP (
        A => S1515,
        B => S5948,
        Y => S5953
    );
NOR_2012: ENTITY WORK.NOR
    PORT MAP (
        A => S1220,
        B => S5953,
        Y => S5954
    );
NOR_2013: ENTITY WORK.NOR
    PORT MAP (
        A => S5952,
        B => S5954,
        Y => S5955
    );
NAND_3574: ENTITY WORK.NAND
    PORT MAP (
        A => S5947,
        B => S5955,
        Y => S282
    );
NAND_3575: ENTITY WORK.NAND
    PORT MAP (
        A => S3898,
        B => S5762,
        Y => S5956
    );
NOR_2014: ENTITY WORK.NOR
    PORT MAP (
        A => S1168,
        B => S1516,
        Y => S5957
    );
NAND_3576: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_0,
        B => S1745,
        Y => S5958
    );
NOT_478: ENTITY WORK.NOT
    PORT MAP (
        A => S5958,
        Y => S5959
    );
NAND_3577: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_1,
        B => S1745,
        Y => S5960
    );
NAND_3578: ENTITY WORK.NAND
    PORT MAP (
        A => S5957,
        B => S5959,
        Y => S5961
    );
NOR_2015: ENTITY WORK.NOR
    PORT MAP (
        A => S5957,
        B => S5959,
        Y => S5962
    );
NAND_3579: ENTITY WORK.NAND
    PORT MAP (
        A => S5948,
        B => S5961,
        Y => S5963
    );
NOR_2016: ENTITY WORK.NOR
    PORT MAP (
        A => S5962,
        B => S5963,
        Y => S5964
    );
NAND_3580: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu1_1,
        B => S5950,
        Y => S5965
    );
NOT_479: ENTITY WORK.NOT
    PORT MAP (
        A => S5965,
        Y => S5966
    );
NOR_2017: ENTITY WORK.NOR
    PORT MAP (
        A => S5964,
        B => S5966,
        Y => S5967
    );
NAND_3581: ENTITY WORK.NAND
    PORT MAP (
        A => S5956,
        B => S5967,
        Y => S283
    );
NOR_2018: ENTITY WORK.NOR
    PORT MAP (
        A => S3899,
        B => S5539,
        Y => S5968
    );
NAND_3582: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu1_2,
        B => S5950,
        Y => S5969
    );
NAND_3583: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_0,
        B => S1848,
        Y => S5970
    );
NOT_480: ENTITY WORK.NOT
    PORT MAP (
        A => S5970,
        Y => S5971
    );
NAND_3584: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_2,
        B => S1515,
        Y => S5972
    );
NAND_3585: ENTITY WORK.NAND
    PORT MAP (
        A => S5960,
        B => S5972,
        Y => S5973
    );
NOR_2019: ENTITY WORK.NOR
    PORT MAP (
        A => S1116,
        B => S1746,
        Y => S5974
    );
NAND_3586: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_2,
        B => S1745,
        Y => S5975
    );
NAND_3587: ENTITY WORK.NAND
    PORT MAP (
        A => S5957,
        B => S5974,
        Y => S5976
    );
NOT_481: ENTITY WORK.NOT
    PORT MAP (
        A => S5976,
        Y => S5977
    );
NAND_3588: ENTITY WORK.NAND
    PORT MAP (
        A => S5973,
        B => S5976,
        Y => S5978
    );
NOT_482: ENTITY WORK.NOT
    PORT MAP (
        A => S5978,
        Y => S5979
    );
NAND_3589: ENTITY WORK.NAND
    PORT MAP (
        A => S5971,
        B => S5979,
        Y => S5980
    );
NOT_483: ENTITY WORK.NOT
    PORT MAP (
        A => S5980,
        Y => S5981
    );
NAND_3590: ENTITY WORK.NAND
    PORT MAP (
        A => S5970,
        B => S5978,
        Y => S5982
    );
NAND_3591: ENTITY WORK.NAND
    PORT MAP (
        A => S5980,
        B => S5982,
        Y => S5983
    );
NOR_2020: ENTITY WORK.NOR
    PORT MAP (
        A => S5961,
        B => S5983,
        Y => S5984
    );
NAND_3592: ENTITY WORK.NAND
    PORT MAP (
        A => S5961,
        B => S5983,
        Y => S5985
    );
NAND_3593: ENTITY WORK.NAND
    PORT MAP (
        A => S5948,
        B => S5985,
        Y => S5986
    );
NOR_2021: ENTITY WORK.NOR
    PORT MAP (
        A => S5984,
        B => S5986,
        Y => S5987
    );
NOR_2022: ENTITY WORK.NOR
    PORT MAP (
        A => S5968,
        B => S5987,
        Y => S5988
    );
NAND_3594: ENTITY WORK.NAND
    PORT MAP (
        A => S5969,
        B => S5988,
        Y => S284
    );
NOR_2023: ENTITY WORK.NOR
    PORT MAP (
        A => S3899,
        B => S5333,
        Y => S5989
    );
NAND_3595: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu1_3,
        B => S5950,
        Y => S5990
    );
NOR_2024: ENTITY WORK.NOR
    PORT MAP (
        A => S1220,
        B => S1953,
        Y => S5991
    );
NAND_3596: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_0,
        B => S1952,
        Y => S5992
    );
NOR_2025: ENTITY WORK.NOR
    PORT MAP (
        A => S5977,
        B => S5981,
        Y => S5993
    );
NOR_2026: ENTITY WORK.NOR
    PORT MAP (
        A => S1168,
        B => S1849,
        Y => S5994
    );
NAND_3597: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_1,
        B => S1848,
        Y => S5995
    );
NOR_2027: ENTITY WORK.NOR
    PORT MAP (
        A => S1065,
        B => S1516,
        Y => S5996
    );
NAND_3598: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_3,
        B => S1515,
        Y => S5997
    );
NOR_2028: ENTITY WORK.NOR
    PORT MAP (
        A => S5974,
        B => S5996,
        Y => S5998
    );
NAND_3599: ENTITY WORK.NAND
    PORT MAP (
        A => S5975,
        B => S5997,
        Y => S5999
    );
NOR_2029: ENTITY WORK.NOR
    PORT MAP (
        A => S1065,
        B => S1746,
        Y => S6000
    );
NAND_3600: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_3,
        B => S1745,
        Y => S6001
    );
NOR_2030: ENTITY WORK.NOR
    PORT MAP (
        A => S5975,
        B => S5997,
        Y => S6002
    );
NAND_3601: ENTITY WORK.NAND
    PORT MAP (
        A => S5974,
        B => S5996,
        Y => S6003
    );
NOR_2031: ENTITY WORK.NOR
    PORT MAP (
        A => S5998,
        B => S6002,
        Y => S6004
    );
NAND_3602: ENTITY WORK.NAND
    PORT MAP (
        A => S5999,
        B => S6003,
        Y => S6005
    );
NOR_2032: ENTITY WORK.NOR
    PORT MAP (
        A => S5995,
        B => S6005,
        Y => S6006
    );
NAND_3603: ENTITY WORK.NAND
    PORT MAP (
        A => S5994,
        B => S6004,
        Y => S6007
    );
NAND_3604: ENTITY WORK.NAND
    PORT MAP (
        A => S5995,
        B => S6005,
        Y => S6008
    );
NAND_3605: ENTITY WORK.NAND
    PORT MAP (
        A => S6007,
        B => S6008,
        Y => S6009
    );
NOR_2033: ENTITY WORK.NOR
    PORT MAP (
        A => S5993,
        B => S6009,
        Y => S6010
    );
NOT_484: ENTITY WORK.NOT
    PORT MAP (
        A => S6010,
        Y => S6011
    );
NAND_3606: ENTITY WORK.NAND
    PORT MAP (
        A => S5993,
        B => S6009,
        Y => S6012
    );
NAND_3607: ENTITY WORK.NAND
    PORT MAP (
        A => S6011,
        B => S6012,
        Y => S6013
    );
NOT_485: ENTITY WORK.NOT
    PORT MAP (
        A => S6013,
        Y => S6014
    );
NAND_3608: ENTITY WORK.NAND
    PORT MAP (
        A => S5991,
        B => S6014,
        Y => S6015
    );
NOT_486: ENTITY WORK.NOT
    PORT MAP (
        A => S6015,
        Y => S6016
    );
NAND_3609: ENTITY WORK.NAND
    PORT MAP (
        A => S5992,
        B => S6013,
        Y => S6017
    );
NOT_487: ENTITY WORK.NOT
    PORT MAP (
        A => S6017,
        Y => S6018
    );
NOR_2034: ENTITY WORK.NOR
    PORT MAP (
        A => S6016,
        B => S6018,
        Y => S6019
    );
NAND_3610: ENTITY WORK.NAND
    PORT MAP (
        A => S5984,
        B => S6019,
        Y => S6020
    );
NOR_2035: ENTITY WORK.NOR
    PORT MAP (
        A => S5984,
        B => S6019,
        Y => S6021
    );
NAND_3611: ENTITY WORK.NAND
    PORT MAP (
        A => S5948,
        B => S6020,
        Y => S6022
    );
NOR_2036: ENTITY WORK.NOR
    PORT MAP (
        A => S6021,
        B => S6022,
        Y => S6023
    );
NOR_2037: ENTITY WORK.NOR
    PORT MAP (
        A => S5989,
        B => S6023,
        Y => S6024
    );
NAND_3612: ENTITY WORK.NAND
    PORT MAP (
        A => S5990,
        B => S6024,
        Y => S285
    );
NOR_2038: ENTITY WORK.NOR
    PORT MAP (
        A => S3899,
        B => S5113,
        Y => S6025
    );
NOR_2039: ENTITY WORK.NOR
    PORT MAP (
        A => S6010,
        B => S6016,
        Y => S6026
    );
NAND_3613: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_0,
        B => S1597,
        Y => S6027
    );
NAND_3614: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_1,
        B => S1952,
        Y => S6028
    );
NAND_3615: ENTITY WORK.NAND
    PORT MAP (
        A => S6027,
        B => S6028,
        Y => S6029
    );
NOR_2040: ENTITY WORK.NOR
    PORT MAP (
        A => S1168,
        B => S1598,
        Y => S6030
    );
NAND_3616: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_1,
        B => S1597,
        Y => S6031
    );
NOR_2041: ENTITY WORK.NOR
    PORT MAP (
        A => S5992,
        B => S6031,
        Y => S6032
    );
NAND_3617: ENTITY WORK.NAND
    PORT MAP (
        A => S5991,
        B => S6030,
        Y => S6033
    );
NAND_3618: ENTITY WORK.NAND
    PORT MAP (
        A => S6029,
        B => S6033,
        Y => S6034
    );
NOT_488: ENTITY WORK.NOT
    PORT MAP (
        A => S6034,
        Y => S6035
    );
NOR_2042: ENTITY WORK.NOR
    PORT MAP (
        A => S6002,
        B => S6006,
        Y => S6036
    );
NAND_3619: ENTITY WORK.NAND
    PORT MAP (
        A => S6003,
        B => S6007,
        Y => S6037
    );
NOR_2043: ENTITY WORK.NOR
    PORT MAP (
        A => S1116,
        B => S1849,
        Y => S6038
    );
NAND_3620: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_2,
        B => S1848,
        Y => S6039
    );
NOR_2044: ENTITY WORK.NOR
    PORT MAP (
        A => S1013,
        B => S1516,
        Y => S6040
    );
NAND_3621: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_4,
        B => S1515,
        Y => S6041
    );
NOR_2045: ENTITY WORK.NOR
    PORT MAP (
        A => S6000,
        B => S6040,
        Y => S6042
    );
NAND_3622: ENTITY WORK.NAND
    PORT MAP (
        A => S6001,
        B => S6041,
        Y => S6043
    );
NOR_2046: ENTITY WORK.NOR
    PORT MAP (
        A => S1013,
        B => S1746,
        Y => S6044
    );
NAND_3623: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_4,
        B => S1745,
        Y => S6045
    );
NOR_2047: ENTITY WORK.NOR
    PORT MAP (
        A => S6001,
        B => S6041,
        Y => S6046
    );
NAND_3624: ENTITY WORK.NAND
    PORT MAP (
        A => S6000,
        B => S6040,
        Y => S6047
    );
NOR_2048: ENTITY WORK.NOR
    PORT MAP (
        A => S6042,
        B => S6046,
        Y => S6048
    );
NAND_3625: ENTITY WORK.NAND
    PORT MAP (
        A => S6043,
        B => S6047,
        Y => S6049
    );
NOR_2049: ENTITY WORK.NOR
    PORT MAP (
        A => S6039,
        B => S6049,
        Y => S6050
    );
NAND_3626: ENTITY WORK.NAND
    PORT MAP (
        A => S6038,
        B => S6048,
        Y => S6051
    );
NOR_2050: ENTITY WORK.NOR
    PORT MAP (
        A => S6038,
        B => S6048,
        Y => S6052
    );
NAND_3627: ENTITY WORK.NAND
    PORT MAP (
        A => S6039,
        B => S6049,
        Y => S6053
    );
NOR_2051: ENTITY WORK.NOR
    PORT MAP (
        A => S6050,
        B => S6052,
        Y => S6054
    );
NAND_3628: ENTITY WORK.NAND
    PORT MAP (
        A => S6051,
        B => S6053,
        Y => S6055
    );
NOR_2052: ENTITY WORK.NOR
    PORT MAP (
        A => S6036,
        B => S6055,
        Y => S6056
    );
NAND_3629: ENTITY WORK.NAND
    PORT MAP (
        A => S6037,
        B => S6054,
        Y => S6057
    );
NAND_3630: ENTITY WORK.NAND
    PORT MAP (
        A => S6036,
        B => S6055,
        Y => S6058
    );
NAND_3631: ENTITY WORK.NAND
    PORT MAP (
        A => S6057,
        B => S6058,
        Y => S6059
    );
NOT_489: ENTITY WORK.NOT
    PORT MAP (
        A => S6059,
        Y => S6060
    );
NAND_3632: ENTITY WORK.NAND
    PORT MAP (
        A => S6035,
        B => S6060,
        Y => S6061
    );
NOT_490: ENTITY WORK.NOT
    PORT MAP (
        A => S6061,
        Y => S6062
    );
NAND_3633: ENTITY WORK.NAND
    PORT MAP (
        A => S6034,
        B => S6059,
        Y => S6063
    );
NAND_3634: ENTITY WORK.NAND
    PORT MAP (
        A => S6061,
        B => S6063,
        Y => S6064
    );
NAND_3635: ENTITY WORK.NAND
    PORT MAP (
        A => S6026,
        B => S6064,
        Y => S6065
    );
NOR_2053: ENTITY WORK.NOR
    PORT MAP (
        A => S6026,
        B => S6064,
        Y => S6066
    );
NOT_491: ENTITY WORK.NOT
    PORT MAP (
        A => S6066,
        Y => S6067
    );
NAND_3636: ENTITY WORK.NAND
    PORT MAP (
        A => S6065,
        B => S6067,
        Y => S6068
    );
NAND_3637: ENTITY WORK.NAND
    PORT MAP (
        A => S6020,
        B => S6068,
        Y => S6069
    );
NOR_2054: ENTITY WORK.NOR
    PORT MAP (
        A => S6020,
        B => S6068,
        Y => S6070
    );
NOR_2055: ENTITY WORK.NOR
    PORT MAP (
        A => S5949,
        B => S6070,
        Y => S6071
    );
NAND_3638: ENTITY WORK.NAND
    PORT MAP (
        A => S6069,
        B => S6071,
        Y => S6072
    );
NAND_3639: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu1_4,
        B => S5950,
        Y => S6073
    );
NOT_492: ENTITY WORK.NOT
    PORT MAP (
        A => S6073,
        Y => S6074
    );
NOR_2056: ENTITY WORK.NOR
    PORT MAP (
        A => S6025,
        B => S6074,
        Y => S6075
    );
NAND_3640: ENTITY WORK.NAND
    PORT MAP (
        A => S6072,
        B => S6075,
        Y => S286
    );
NOR_2057: ENTITY WORK.NOR
    PORT MAP (
        A => S3899,
        B => S4896,
        Y => S6076
    );
NAND_3641: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu1_5,
        B => S5950,
        Y => S6077
    );
NOR_2058: ENTITY WORK.NOR
    PORT MAP (
        A => S6056,
        B => S6062,
        Y => S6078
    );
NAND_3642: ENTITY WORK.NAND
    PORT MAP (
        A => S6057,
        B => S6061,
        Y => S6079
    );
NOR_2059: ENTITY WORK.NOR
    PORT MAP (
        A => S1220,
        B => S2107,
        Y => S6080
    );
NAND_3643: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_0,
        B => S2106,
        Y => S6081
    );
NOR_2060: ENTITY WORK.NOR
    PORT MAP (
        A => S1116,
        B => S1953,
        Y => S6082
    );
NAND_3644: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_2,
        B => S1952,
        Y => S6083
    );
NOR_2061: ENTITY WORK.NOR
    PORT MAP (
        A => S6030,
        B => S6082,
        Y => S6084
    );
NAND_3645: ENTITY WORK.NAND
    PORT MAP (
        A => S6031,
        B => S6083,
        Y => S6085
    );
NOR_2062: ENTITY WORK.NOR
    PORT MAP (
        A => S1116,
        B => S1598,
        Y => S6086
    );
NAND_3646: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_2,
        B => S1597,
        Y => S6087
    );
NOR_2063: ENTITY WORK.NOR
    PORT MAP (
        A => S6031,
        B => S6083,
        Y => S6088
    );
NAND_3647: ENTITY WORK.NAND
    PORT MAP (
        A => S6030,
        B => S6082,
        Y => S6089
    );
NOR_2064: ENTITY WORK.NOR
    PORT MAP (
        A => S6084,
        B => S6088,
        Y => S6090
    );
NAND_3648: ENTITY WORK.NAND
    PORT MAP (
        A => S6085,
        B => S6089,
        Y => S6091
    );
NOR_2065: ENTITY WORK.NOR
    PORT MAP (
        A => S6081,
        B => S6091,
        Y => S6092
    );
NAND_3649: ENTITY WORK.NAND
    PORT MAP (
        A => S6080,
        B => S6090,
        Y => S6093
    );
NOR_2066: ENTITY WORK.NOR
    PORT MAP (
        A => S6080,
        B => S6090,
        Y => S6094
    );
NAND_3650: ENTITY WORK.NAND
    PORT MAP (
        A => S6081,
        B => S6091,
        Y => S6095
    );
NOR_2067: ENTITY WORK.NOR
    PORT MAP (
        A => S6092,
        B => S6094,
        Y => S6096
    );
NAND_3651: ENTITY WORK.NAND
    PORT MAP (
        A => S6093,
        B => S6095,
        Y => S6097
    );
NOR_2068: ENTITY WORK.NOR
    PORT MAP (
        A => S6046,
        B => S6050,
        Y => S6098
    );
NAND_3652: ENTITY WORK.NAND
    PORT MAP (
        A => S6047,
        B => S6051,
        Y => S6099
    );
NOR_2069: ENTITY WORK.NOR
    PORT MAP (
        A => S1065,
        B => S1849,
        Y => S6100
    );
NAND_3653: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_3,
        B => S1848,
        Y => S6101
    );
NOR_2070: ENTITY WORK.NOR
    PORT MAP (
        A => S963,
        B => S1516,
        Y => S6102
    );
NAND_3654: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_5,
        B => S1515,
        Y => S6103
    );
NOR_2071: ENTITY WORK.NOR
    PORT MAP (
        A => S6044,
        B => S6102,
        Y => S6104
    );
NAND_3655: ENTITY WORK.NAND
    PORT MAP (
        A => S6045,
        B => S6103,
        Y => S6105
    );
NOR_2072: ENTITY WORK.NOR
    PORT MAP (
        A => S963,
        B => S1746,
        Y => S6106
    );
NAND_3656: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_5,
        B => S1745,
        Y => S6107
    );
NOR_2073: ENTITY WORK.NOR
    PORT MAP (
        A => S6045,
        B => S6103,
        Y => S6108
    );
NAND_3657: ENTITY WORK.NAND
    PORT MAP (
        A => S6044,
        B => S6102,
        Y => S6109
    );
NOR_2074: ENTITY WORK.NOR
    PORT MAP (
        A => S6104,
        B => S6108,
        Y => S6110
    );
NAND_3658: ENTITY WORK.NAND
    PORT MAP (
        A => S6105,
        B => S6109,
        Y => S6111
    );
NOR_2075: ENTITY WORK.NOR
    PORT MAP (
        A => S6101,
        B => S6111,
        Y => S6112
    );
NAND_3659: ENTITY WORK.NAND
    PORT MAP (
        A => S6100,
        B => S6110,
        Y => S6113
    );
NOR_2076: ENTITY WORK.NOR
    PORT MAP (
        A => S6100,
        B => S6110,
        Y => S6114
    );
NAND_3660: ENTITY WORK.NAND
    PORT MAP (
        A => S6101,
        B => S6111,
        Y => S6115
    );
NOR_2077: ENTITY WORK.NOR
    PORT MAP (
        A => S6112,
        B => S6114,
        Y => S6116
    );
NAND_3661: ENTITY WORK.NAND
    PORT MAP (
        A => S6113,
        B => S6115,
        Y => S6117
    );
NOR_2078: ENTITY WORK.NOR
    PORT MAP (
        A => S6098,
        B => S6117,
        Y => S6118
    );
NAND_3662: ENTITY WORK.NAND
    PORT MAP (
        A => S6099,
        B => S6116,
        Y => S6119
    );
NOR_2079: ENTITY WORK.NOR
    PORT MAP (
        A => S6099,
        B => S6116,
        Y => S6120
    );
NAND_3663: ENTITY WORK.NAND
    PORT MAP (
        A => S6098,
        B => S6117,
        Y => S6121
    );
NOR_2080: ENTITY WORK.NOR
    PORT MAP (
        A => S6118,
        B => S6120,
        Y => S6122
    );
NAND_3664: ENTITY WORK.NAND
    PORT MAP (
        A => S6119,
        B => S6121,
        Y => S6123
    );
NOR_2081: ENTITY WORK.NOR
    PORT MAP (
        A => S6097,
        B => S6123,
        Y => S6124
    );
NAND_3665: ENTITY WORK.NAND
    PORT MAP (
        A => S6096,
        B => S6122,
        Y => S6125
    );
NOR_2082: ENTITY WORK.NOR
    PORT MAP (
        A => S6096,
        B => S6122,
        Y => S6126
    );
NAND_3666: ENTITY WORK.NAND
    PORT MAP (
        A => S6097,
        B => S6123,
        Y => S6127
    );
NOR_2083: ENTITY WORK.NOR
    PORT MAP (
        A => S6124,
        B => S6126,
        Y => S6128
    );
NAND_3667: ENTITY WORK.NAND
    PORT MAP (
        A => S6125,
        B => S6127,
        Y => S6129
    );
NOR_2084: ENTITY WORK.NOR
    PORT MAP (
        A => S6078,
        B => S6129,
        Y => S6130
    );
NOR_2085: ENTITY WORK.NOR
    PORT MAP (
        A => S6079,
        B => S6128,
        Y => S6131
    );
NOR_2086: ENTITY WORK.NOR
    PORT MAP (
        A => S6130,
        B => S6131,
        Y => S6132
    );
NOT_493: ENTITY WORK.NOT
    PORT MAP (
        A => S6132,
        Y => S6133
    );
NOR_2087: ENTITY WORK.NOR
    PORT MAP (
        A => S6033,
        B => S6133,
        Y => S6134
    );
NOR_2088: ENTITY WORK.NOR
    PORT MAP (
        A => S6032,
        B => S6132,
        Y => S6135
    );
NOR_2089: ENTITY WORK.NOR
    PORT MAP (
        A => S6134,
        B => S6135,
        Y => S6136
    );
NAND_3668: ENTITY WORK.NAND
    PORT MAP (
        A => S6066,
        B => S6136,
        Y => S6137
    );
NOT_494: ENTITY WORK.NOT
    PORT MAP (
        A => S6137,
        Y => S6138
    );
NOR_2090: ENTITY WORK.NOR
    PORT MAP (
        A => S6066,
        B => S6136,
        Y => S6139
    );
NOR_2091: ENTITY WORK.NOR
    PORT MAP (
        A => S6138,
        B => S6139,
        Y => S6140
    );
NAND_3669: ENTITY WORK.NAND
    PORT MAP (
        A => S6070,
        B => S6140,
        Y => S6141
    );
NOR_2092: ENTITY WORK.NOR
    PORT MAP (
        A => S6070,
        B => S6140,
        Y => S6142
    );
NAND_3670: ENTITY WORK.NAND
    PORT MAP (
        A => S5948,
        B => S6141,
        Y => S6143
    );
NOR_2093: ENTITY WORK.NOR
    PORT MAP (
        A => S6142,
        B => S6143,
        Y => S6144
    );
NOR_2094: ENTITY WORK.NOR
    PORT MAP (
        A => S6076,
        B => S6144,
        Y => S6145
    );
NAND_3671: ENTITY WORK.NAND
    PORT MAP (
        A => S6077,
        B => S6145,
        Y => S287
    );
NOR_2095: ENTITY WORK.NOR
    PORT MAP (
        A => S3899,
        B => S4709,
        Y => S6146
    );
NAND_3672: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu1_6,
        B => S5950,
        Y => S6147
    );
NOR_2096: ENTITY WORK.NOR
    PORT MAP (
        A => S6130,
        B => S6134,
        Y => S6148
    );
NOT_495: ENTITY WORK.NOT
    PORT MAP (
        A => S6148,
        Y => S6149
    );
NOR_2097: ENTITY WORK.NOR
    PORT MAP (
        A => S1220,
        B => S2206,
        Y => S6150
    );
NAND_3673: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_0,
        B => S2205,
        Y => S6151
    );
NOR_2098: ENTITY WORK.NOR
    PORT MAP (
        A => S6088,
        B => S6092,
        Y => S6152
    );
NAND_3674: ENTITY WORK.NAND
    PORT MAP (
        A => S6089,
        B => S6093,
        Y => S6153
    );
NOR_2099: ENTITY WORK.NOR
    PORT MAP (
        A => S6151,
        B => S6152,
        Y => S6154
    );
NAND_3675: ENTITY WORK.NAND
    PORT MAP (
        A => S6150,
        B => S6153,
        Y => S6155
    );
NAND_3676: ENTITY WORK.NAND
    PORT MAP (
        A => S6151,
        B => S6152,
        Y => S6156
    );
NAND_3677: ENTITY WORK.NAND
    PORT MAP (
        A => S6155,
        B => S6156,
        Y => S6157
    );
NOT_496: ENTITY WORK.NOT
    PORT MAP (
        A => S6157,
        Y => S6158
    );
NOR_2100: ENTITY WORK.NOR
    PORT MAP (
        A => S6118,
        B => S6124,
        Y => S6159
    );
NAND_3678: ENTITY WORK.NAND
    PORT MAP (
        A => S6119,
        B => S6125,
        Y => S6160
    );
NOR_2101: ENTITY WORK.NOR
    PORT MAP (
        A => S1168,
        B => S2107,
        Y => S6161
    );
NAND_3679: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_1,
        B => S2106,
        Y => S6162
    );
NOR_2102: ENTITY WORK.NOR
    PORT MAP (
        A => S1065,
        B => S1953,
        Y => S6163
    );
NAND_3680: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_3,
        B => S1952,
        Y => S6164
    );
NOR_2103: ENTITY WORK.NOR
    PORT MAP (
        A => S6086,
        B => S6163,
        Y => S6165
    );
NAND_3681: ENTITY WORK.NAND
    PORT MAP (
        A => S6087,
        B => S6164,
        Y => S6166
    );
NOR_2104: ENTITY WORK.NOR
    PORT MAP (
        A => S1065,
        B => S1598,
        Y => S6167
    );
NAND_3682: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_3,
        B => S1597,
        Y => S6168
    );
NOR_2105: ENTITY WORK.NOR
    PORT MAP (
        A => S6087,
        B => S6164,
        Y => S6169
    );
NAND_3683: ENTITY WORK.NAND
    PORT MAP (
        A => S6086,
        B => S6163,
        Y => S6170
    );
NOR_2106: ENTITY WORK.NOR
    PORT MAP (
        A => S6165,
        B => S6169,
        Y => S6171
    );
NAND_3684: ENTITY WORK.NAND
    PORT MAP (
        A => S6166,
        B => S6170,
        Y => S6172
    );
NOR_2107: ENTITY WORK.NOR
    PORT MAP (
        A => S6162,
        B => S6172,
        Y => S6173
    );
NAND_3685: ENTITY WORK.NAND
    PORT MAP (
        A => S6161,
        B => S6171,
        Y => S6174
    );
NOR_2108: ENTITY WORK.NOR
    PORT MAP (
        A => S6161,
        B => S6171,
        Y => S6175
    );
NAND_3686: ENTITY WORK.NAND
    PORT MAP (
        A => S6162,
        B => S6172,
        Y => S6176
    );
NOR_2109: ENTITY WORK.NOR
    PORT MAP (
        A => S6173,
        B => S6175,
        Y => S6177
    );
NAND_3687: ENTITY WORK.NAND
    PORT MAP (
        A => S6174,
        B => S6176,
        Y => S6178
    );
NOR_2110: ENTITY WORK.NOR
    PORT MAP (
        A => S6108,
        B => S6112,
        Y => S6179
    );
NAND_3688: ENTITY WORK.NAND
    PORT MAP (
        A => S6109,
        B => S6113,
        Y => S6180
    );
NOR_2111: ENTITY WORK.NOR
    PORT MAP (
        A => S1013,
        B => S1849,
        Y => S6181
    );
NAND_3689: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_4,
        B => S1848,
        Y => S6182
    );
NOR_2112: ENTITY WORK.NOR
    PORT MAP (
        A => S910,
        B => S1516,
        Y => S6183
    );
NAND_3690: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_6,
        B => S1515,
        Y => S6184
    );
NOR_2113: ENTITY WORK.NOR
    PORT MAP (
        A => S6106,
        B => S6183,
        Y => S6185
    );
NAND_3691: ENTITY WORK.NAND
    PORT MAP (
        A => S6107,
        B => S6184,
        Y => S6186
    );
NOR_2114: ENTITY WORK.NOR
    PORT MAP (
        A => S910,
        B => S1746,
        Y => S6187
    );
NAND_3692: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_6,
        B => S1745,
        Y => S6188
    );
NOR_2115: ENTITY WORK.NOR
    PORT MAP (
        A => S6107,
        B => S6184,
        Y => S6189
    );
NAND_3693: ENTITY WORK.NAND
    PORT MAP (
        A => S6106,
        B => S6183,
        Y => S6190
    );
NOR_2116: ENTITY WORK.NOR
    PORT MAP (
        A => S6185,
        B => S6189,
        Y => S6191
    );
NAND_3694: ENTITY WORK.NAND
    PORT MAP (
        A => S6186,
        B => S6190,
        Y => S6192
    );
NOR_2117: ENTITY WORK.NOR
    PORT MAP (
        A => S6182,
        B => S6192,
        Y => S6193
    );
NAND_3695: ENTITY WORK.NAND
    PORT MAP (
        A => S6181,
        B => S6191,
        Y => S6194
    );
NOR_2118: ENTITY WORK.NOR
    PORT MAP (
        A => S6181,
        B => S6191,
        Y => S6195
    );
NAND_3696: ENTITY WORK.NAND
    PORT MAP (
        A => S6182,
        B => S6192,
        Y => S6196
    );
NOR_2119: ENTITY WORK.NOR
    PORT MAP (
        A => S6193,
        B => S6195,
        Y => S6197
    );
NAND_3697: ENTITY WORK.NAND
    PORT MAP (
        A => S6194,
        B => S6196,
        Y => S6198
    );
NOR_2120: ENTITY WORK.NOR
    PORT MAP (
        A => S6179,
        B => S6198,
        Y => S6199
    );
NAND_3698: ENTITY WORK.NAND
    PORT MAP (
        A => S6180,
        B => S6197,
        Y => S6200
    );
NOR_2121: ENTITY WORK.NOR
    PORT MAP (
        A => S6180,
        B => S6197,
        Y => S6201
    );
NAND_3699: ENTITY WORK.NAND
    PORT MAP (
        A => S6179,
        B => S6198,
        Y => S6202
    );
NOR_2122: ENTITY WORK.NOR
    PORT MAP (
        A => S6199,
        B => S6201,
        Y => S6203
    );
NAND_3700: ENTITY WORK.NAND
    PORT MAP (
        A => S6200,
        B => S6202,
        Y => S6204
    );
NOR_2123: ENTITY WORK.NOR
    PORT MAP (
        A => S6178,
        B => S6204,
        Y => S6205
    );
NAND_3701: ENTITY WORK.NAND
    PORT MAP (
        A => S6177,
        B => S6203,
        Y => S6206
    );
NOR_2124: ENTITY WORK.NOR
    PORT MAP (
        A => S6177,
        B => S6203,
        Y => S6207
    );
NAND_3702: ENTITY WORK.NAND
    PORT MAP (
        A => S6178,
        B => S6204,
        Y => S6208
    );
NOR_2125: ENTITY WORK.NOR
    PORT MAP (
        A => S6205,
        B => S6207,
        Y => S6209
    );
NAND_3703: ENTITY WORK.NAND
    PORT MAP (
        A => S6206,
        B => S6208,
        Y => S6210
    );
NOR_2126: ENTITY WORK.NOR
    PORT MAP (
        A => S6159,
        B => S6210,
        Y => S6211
    );
NAND_3704: ENTITY WORK.NAND
    PORT MAP (
        A => S6160,
        B => S6209,
        Y => S6212
    );
NAND_3705: ENTITY WORK.NAND
    PORT MAP (
        A => S6159,
        B => S6210,
        Y => S6213
    );
NAND_3706: ENTITY WORK.NAND
    PORT MAP (
        A => S6212,
        B => S6213,
        Y => S6214
    );
NOT_497: ENTITY WORK.NOT
    PORT MAP (
        A => S6214,
        Y => S6215
    );
NAND_3707: ENTITY WORK.NAND
    PORT MAP (
        A => S6158,
        B => S6215,
        Y => S6216
    );
NOT_498: ENTITY WORK.NOT
    PORT MAP (
        A => S6216,
        Y => S6217
    );
NAND_3708: ENTITY WORK.NAND
    PORT MAP (
        A => S6157,
        B => S6214,
        Y => S6218
    );
NAND_3709: ENTITY WORK.NAND
    PORT MAP (
        A => S6216,
        B => S6218,
        Y => S6219
    );
NOT_499: ENTITY WORK.NOT
    PORT MAP (
        A => S6219,
        Y => S6220
    );
NAND_3710: ENTITY WORK.NAND
    PORT MAP (
        A => S6148,
        B => S6219,
        Y => S6221
    );
NAND_3711: ENTITY WORK.NAND
    PORT MAP (
        A => S6149,
        B => S6220,
        Y => S6222
    );
NOT_500: ENTITY WORK.NOT
    PORT MAP (
        A => S6222,
        Y => S6223
    );
NAND_3712: ENTITY WORK.NAND
    PORT MAP (
        A => S6221,
        B => S6222,
        Y => S6224
    );
NOR_2127: ENTITY WORK.NOR
    PORT MAP (
        A => S6137,
        B => S6224,
        Y => S6225
    );
NOT_501: ENTITY WORK.NOT
    PORT MAP (
        A => S6225,
        Y => S6226
    );
NAND_3713: ENTITY WORK.NAND
    PORT MAP (
        A => S6137,
        B => S6224,
        Y => S6227
    );
NAND_3714: ENTITY WORK.NAND
    PORT MAP (
        A => S6226,
        B => S6227,
        Y => S6228
    );
NOR_2128: ENTITY WORK.NOR
    PORT MAP (
        A => S6141,
        B => S6228,
        Y => S6229
    );
NAND_3715: ENTITY WORK.NAND
    PORT MAP (
        A => S6141,
        B => S6228,
        Y => S6230
    );
NAND_3716: ENTITY WORK.NAND
    PORT MAP (
        A => S5948,
        B => S6230,
        Y => S6231
    );
NOR_2129: ENTITY WORK.NOR
    PORT MAP (
        A => S6229,
        B => S6231,
        Y => S6232
    );
NOR_2130: ENTITY WORK.NOR
    PORT MAP (
        A => S6146,
        B => S6232,
        Y => S6233
    );
NAND_3717: ENTITY WORK.NAND
    PORT MAP (
        A => S6147,
        B => S6233,
        Y => S288
    );
NOR_2131: ENTITY WORK.NOR
    PORT MAP (
        A => S3899,
        B => S4571,
        Y => S6234
    );
NAND_3718: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu1_7,
        B => S5950,
        Y => S6235
    );
NOR_2132: ENTITY WORK.NOR
    PORT MAP (
        A => S6211,
        B => S6217,
        Y => S6236
    );
NAND_3719: ENTITY WORK.NAND
    PORT MAP (
        A => S6212,
        B => S6216,
        Y => S6237
    );
NOR_2133: ENTITY WORK.NOR
    PORT MAP (
        A => S1220,
        B => S2312,
        Y => S6238
    );
NAND_3720: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_0,
        B => S2311,
        Y => S6239
    );
NOR_2134: ENTITY WORK.NOR
    PORT MAP (
        A => S1168,
        B => S2206,
        Y => S6240
    );
NAND_3721: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_1,
        B => S2205,
        Y => S6241
    );
NOR_2135: ENTITY WORK.NOR
    PORT MAP (
        A => S6238,
        B => S6240,
        Y => S6242
    );
NAND_3722: ENTITY WORK.NAND
    PORT MAP (
        A => S6239,
        B => S6241,
        Y => S6243
    );
NOR_2136: ENTITY WORK.NOR
    PORT MAP (
        A => S1168,
        B => S2312,
        Y => S6244
    );
NAND_3723: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_1,
        B => S2311,
        Y => S6245
    );
NOR_2137: ENTITY WORK.NOR
    PORT MAP (
        A => S6151,
        B => S6245,
        Y => S6246
    );
NAND_3724: ENTITY WORK.NAND
    PORT MAP (
        A => S6150,
        B => S6244,
        Y => S6247
    );
NOR_2138: ENTITY WORK.NOR
    PORT MAP (
        A => S6242,
        B => S6246,
        Y => S6248
    );
NAND_3725: ENTITY WORK.NAND
    PORT MAP (
        A => S6243,
        B => S6247,
        Y => S6249
    );
NOR_2139: ENTITY WORK.NOR
    PORT MAP (
        A => S6169,
        B => S6173,
        Y => S6250
    );
NAND_3726: ENTITY WORK.NAND
    PORT MAP (
        A => S6170,
        B => S6174,
        Y => S6251
    );
NOR_2140: ENTITY WORK.NOR
    PORT MAP (
        A => S6248,
        B => S6251,
        Y => S6252
    );
NAND_3727: ENTITY WORK.NAND
    PORT MAP (
        A => S6249,
        B => S6250,
        Y => S6253
    );
NOR_2141: ENTITY WORK.NOR
    PORT MAP (
        A => S6249,
        B => S6250,
        Y => S6254
    );
NAND_3728: ENTITY WORK.NAND
    PORT MAP (
        A => S6248,
        B => S6251,
        Y => S6255
    );
NOR_2142: ENTITY WORK.NOR
    PORT MAP (
        A => S6252,
        B => S6254,
        Y => S6256
    );
NAND_3729: ENTITY WORK.NAND
    PORT MAP (
        A => S6253,
        B => S6255,
        Y => S6257
    );
NOR_2143: ENTITY WORK.NOR
    PORT MAP (
        A => S6199,
        B => S6205,
        Y => S6258
    );
NAND_3730: ENTITY WORK.NAND
    PORT MAP (
        A => S6200,
        B => S6206,
        Y => S6259
    );
NOR_2144: ENTITY WORK.NOR
    PORT MAP (
        A => S1116,
        B => S2107,
        Y => S6260
    );
NAND_3731: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_2,
        B => S2106,
        Y => S6261
    );
NOR_2145: ENTITY WORK.NOR
    PORT MAP (
        A => S1013,
        B => S1953,
        Y => S6262
    );
NAND_3732: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_4,
        B => S1952,
        Y => S6263
    );
NOR_2146: ENTITY WORK.NOR
    PORT MAP (
        A => S6167,
        B => S6262,
        Y => S6264
    );
NAND_3733: ENTITY WORK.NAND
    PORT MAP (
        A => S6168,
        B => S6263,
        Y => S6265
    );
NOR_2147: ENTITY WORK.NOR
    PORT MAP (
        A => S1013,
        B => S1598,
        Y => S6266
    );
NAND_3734: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_4,
        B => S1597,
        Y => S6267
    );
NOR_2148: ENTITY WORK.NOR
    PORT MAP (
        A => S6168,
        B => S6263,
        Y => S6268
    );
NAND_3735: ENTITY WORK.NAND
    PORT MAP (
        A => S6167,
        B => S6262,
        Y => S6269
    );
NOR_2149: ENTITY WORK.NOR
    PORT MAP (
        A => S6264,
        B => S6268,
        Y => S6270
    );
NAND_3736: ENTITY WORK.NAND
    PORT MAP (
        A => S6265,
        B => S6269,
        Y => S6271
    );
NOR_2150: ENTITY WORK.NOR
    PORT MAP (
        A => S6261,
        B => S6271,
        Y => S6272
    );
NAND_3737: ENTITY WORK.NAND
    PORT MAP (
        A => S6260,
        B => S6270,
        Y => S6273
    );
NOR_2151: ENTITY WORK.NOR
    PORT MAP (
        A => S6260,
        B => S6270,
        Y => S6274
    );
NAND_3738: ENTITY WORK.NAND
    PORT MAP (
        A => S6261,
        B => S6271,
        Y => S6275
    );
NOR_2152: ENTITY WORK.NOR
    PORT MAP (
        A => S6272,
        B => S6274,
        Y => S6276
    );
NAND_3739: ENTITY WORK.NAND
    PORT MAP (
        A => S6273,
        B => S6275,
        Y => S6277
    );
NOR_2153: ENTITY WORK.NOR
    PORT MAP (
        A => S6189,
        B => S6193,
        Y => S6278
    );
NAND_3740: ENTITY WORK.NAND
    PORT MAP (
        A => S6190,
        B => S6194,
        Y => S6279
    );
NOR_2154: ENTITY WORK.NOR
    PORT MAP (
        A => S963,
        B => S1849,
        Y => S6280
    );
NAND_3741: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_5,
        B => S1848,
        Y => S6281
    );
NOR_2155: ENTITY WORK.NOR
    PORT MAP (
        A => S858,
        B => S1516,
        Y => S6282
    );
NAND_3742: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_7,
        B => S1515,
        Y => S6283
    );
NOR_2156: ENTITY WORK.NOR
    PORT MAP (
        A => S6187,
        B => S6282,
        Y => S6284
    );
NAND_3743: ENTITY WORK.NAND
    PORT MAP (
        A => S6188,
        B => S6283,
        Y => S6285
    );
NOR_2157: ENTITY WORK.NOR
    PORT MAP (
        A => S858,
        B => S1746,
        Y => S6286
    );
NAND_3744: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_7,
        B => S1745,
        Y => S6287
    );
NOR_2158: ENTITY WORK.NOR
    PORT MAP (
        A => S6188,
        B => S6283,
        Y => S6288
    );
NAND_3745: ENTITY WORK.NAND
    PORT MAP (
        A => S6187,
        B => S6282,
        Y => S6289
    );
NOR_2159: ENTITY WORK.NOR
    PORT MAP (
        A => S6284,
        B => S6288,
        Y => S6290
    );
NAND_3746: ENTITY WORK.NAND
    PORT MAP (
        A => S6285,
        B => S6289,
        Y => S6291
    );
NOR_2160: ENTITY WORK.NOR
    PORT MAP (
        A => S6281,
        B => S6291,
        Y => S6292
    );
NAND_3747: ENTITY WORK.NAND
    PORT MAP (
        A => S6280,
        B => S6290,
        Y => S6293
    );
NOR_2161: ENTITY WORK.NOR
    PORT MAP (
        A => S6280,
        B => S6290,
        Y => S6294
    );
NAND_3748: ENTITY WORK.NAND
    PORT MAP (
        A => S6281,
        B => S6291,
        Y => S6295
    );
NOR_2162: ENTITY WORK.NOR
    PORT MAP (
        A => S6292,
        B => S6294,
        Y => S6296
    );
NAND_3749: ENTITY WORK.NAND
    PORT MAP (
        A => S6293,
        B => S6295,
        Y => S6297
    );
NOR_2163: ENTITY WORK.NOR
    PORT MAP (
        A => S6278,
        B => S6297,
        Y => S6298
    );
NAND_3750: ENTITY WORK.NAND
    PORT MAP (
        A => S6279,
        B => S6296,
        Y => S6299
    );
NOR_2164: ENTITY WORK.NOR
    PORT MAP (
        A => S6279,
        B => S6296,
        Y => S6300
    );
NAND_3751: ENTITY WORK.NAND
    PORT MAP (
        A => S6278,
        B => S6297,
        Y => S6301
    );
NOR_2165: ENTITY WORK.NOR
    PORT MAP (
        A => S6298,
        B => S6300,
        Y => S6302
    );
NAND_3752: ENTITY WORK.NAND
    PORT MAP (
        A => S6299,
        B => S6301,
        Y => S6303
    );
NOR_2166: ENTITY WORK.NOR
    PORT MAP (
        A => S6277,
        B => S6303,
        Y => S6304
    );
NAND_3753: ENTITY WORK.NAND
    PORT MAP (
        A => S6276,
        B => S6302,
        Y => S6305
    );
NOR_2167: ENTITY WORK.NOR
    PORT MAP (
        A => S6276,
        B => S6302,
        Y => S6306
    );
NAND_3754: ENTITY WORK.NAND
    PORT MAP (
        A => S6277,
        B => S6303,
        Y => S6307
    );
NOR_2168: ENTITY WORK.NOR
    PORT MAP (
        A => S6304,
        B => S6306,
        Y => S6308
    );
NAND_3755: ENTITY WORK.NAND
    PORT MAP (
        A => S6305,
        B => S6307,
        Y => S6309
    );
NOR_2169: ENTITY WORK.NOR
    PORT MAP (
        A => S6258,
        B => S6309,
        Y => S6310
    );
NAND_3756: ENTITY WORK.NAND
    PORT MAP (
        A => S6259,
        B => S6308,
        Y => S6311
    );
NOR_2170: ENTITY WORK.NOR
    PORT MAP (
        A => S6259,
        B => S6308,
        Y => S6312
    );
NAND_3757: ENTITY WORK.NAND
    PORT MAP (
        A => S6258,
        B => S6309,
        Y => S6313
    );
NOR_2171: ENTITY WORK.NOR
    PORT MAP (
        A => S6310,
        B => S6312,
        Y => S6314
    );
NAND_3758: ENTITY WORK.NAND
    PORT MAP (
        A => S6311,
        B => S6313,
        Y => S6315
    );
NOR_2172: ENTITY WORK.NOR
    PORT MAP (
        A => S6257,
        B => S6315,
        Y => S6316
    );
NAND_3759: ENTITY WORK.NAND
    PORT MAP (
        A => S6256,
        B => S6314,
        Y => S6317
    );
NOR_2173: ENTITY WORK.NOR
    PORT MAP (
        A => S6256,
        B => S6314,
        Y => S6318
    );
NAND_3760: ENTITY WORK.NAND
    PORT MAP (
        A => S6257,
        B => S6315,
        Y => S6319
    );
NOR_2174: ENTITY WORK.NOR
    PORT MAP (
        A => S6316,
        B => S6318,
        Y => S6320
    );
NAND_3761: ENTITY WORK.NAND
    PORT MAP (
        A => S6317,
        B => S6319,
        Y => S6321
    );
NOR_2175: ENTITY WORK.NOR
    PORT MAP (
        A => S6236,
        B => S6321,
        Y => S6322
    );
NAND_3762: ENTITY WORK.NAND
    PORT MAP (
        A => S6237,
        B => S6320,
        Y => S6323
    );
NAND_3763: ENTITY WORK.NAND
    PORT MAP (
        A => S6236,
        B => S6321,
        Y => S6324
    );
NAND_3764: ENTITY WORK.NAND
    PORT MAP (
        A => S6323,
        B => S6324,
        Y => S6325
    );
NOT_502: ENTITY WORK.NOT
    PORT MAP (
        A => S6325,
        Y => S6326
    );
NAND_3765: ENTITY WORK.NAND
    PORT MAP (
        A => S6154,
        B => S6326,
        Y => S6327
    );
NOT_503: ENTITY WORK.NOT
    PORT MAP (
        A => S6327,
        Y => S6328
    );
NAND_3766: ENTITY WORK.NAND
    PORT MAP (
        A => S6155,
        B => S6325,
        Y => S6329
    );
NAND_3767: ENTITY WORK.NAND
    PORT MAP (
        A => S6327,
        B => S6329,
        Y => S6330
    );
NOT_504: ENTITY WORK.NOT
    PORT MAP (
        A => S6330,
        Y => S6331
    );
NAND_3768: ENTITY WORK.NAND
    PORT MAP (
        A => S6223,
        B => S6331,
        Y => S6332
    );
NOT_505: ENTITY WORK.NOT
    PORT MAP (
        A => S6332,
        Y => S6333
    );
NAND_3769: ENTITY WORK.NAND
    PORT MAP (
        A => S6222,
        B => S6330,
        Y => S6334
    );
NAND_3770: ENTITY WORK.NAND
    PORT MAP (
        A => S6332,
        B => S6334,
        Y => S6335
    );
NOT_506: ENTITY WORK.NOT
    PORT MAP (
        A => S6335,
        Y => S6336
    );
NAND_3771: ENTITY WORK.NAND
    PORT MAP (
        A => S6229,
        B => S6336,
        Y => S6337
    );
NAND_3772: ENTITY WORK.NAND
    PORT MAP (
        A => S5948,
        B => S6337,
        Y => S6338
    );
NOR_2176: ENTITY WORK.NOR
    PORT MAP (
        A => S6225,
        B => S6229,
        Y => S6339
    );
NAND_3773: ENTITY WORK.NAND
    PORT MAP (
        A => S6335,
        B => S6339,
        Y => S6340
    );
NAND_3774: ENTITY WORK.NAND
    PORT MAP (
        A => S6225,
        B => S6336,
        Y => S6341
    );
NAND_3775: ENTITY WORK.NAND
    PORT MAP (
        A => S6340,
        B => S6341,
        Y => S6342
    );
NOR_2177: ENTITY WORK.NOR
    PORT MAP (
        A => S6338,
        B => S6342,
        Y => S6343
    );
NOR_2178: ENTITY WORK.NOR
    PORT MAP (
        A => S6234,
        B => S6343,
        Y => S6344
    );
NAND_3776: ENTITY WORK.NAND
    PORT MAP (
        A => S6235,
        B => S6344,
        Y => S289
    );
NOR_2179: ENTITY WORK.NOR
    PORT MAP (
        A => S3899,
        B => S4430,
        Y => S6345
    );
NAND_3777: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu1_8,
        B => S5950,
        Y => S6346
    );
NOR_2180: ENTITY WORK.NOR
    PORT MAP (
        A => S6322,
        B => S6328,
        Y => S6347
    );
NAND_3778: ENTITY WORK.NAND
    PORT MAP (
        A => S6323,
        B => S6327,
        Y => S6348
    );
NOR_2181: ENTITY WORK.NOR
    PORT MAP (
        A => S6310,
        B => S6316,
        Y => S6349
    );
NAND_3779: ENTITY WORK.NAND
    PORT MAP (
        A => S6311,
        B => S6317,
        Y => S6350
    );
NOR_2182: ENTITY WORK.NOR
    PORT MAP (
        A => S1220,
        B => S2418,
        Y => S6351
    );
NAND_3780: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_0,
        B => S2417,
        Y => S6352
    );
NOR_2183: ENTITY WORK.NOR
    PORT MAP (
        A => S1116,
        B => S2206,
        Y => S6353
    );
NAND_3781: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_2,
        B => S2205,
        Y => S6354
    );
NOR_2184: ENTITY WORK.NOR
    PORT MAP (
        A => S6244,
        B => S6353,
        Y => S6355
    );
NAND_3782: ENTITY WORK.NAND
    PORT MAP (
        A => S6245,
        B => S6354,
        Y => S6356
    );
NOR_2185: ENTITY WORK.NOR
    PORT MAP (
        A => S1116,
        B => S2312,
        Y => S6357
    );
NAND_3783: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_2,
        B => S2311,
        Y => S6358
    );
NOR_2186: ENTITY WORK.NOR
    PORT MAP (
        A => S6245,
        B => S6354,
        Y => S6359
    );
NAND_3784: ENTITY WORK.NAND
    PORT MAP (
        A => S6244,
        B => S6353,
        Y => S6360
    );
NOR_2187: ENTITY WORK.NOR
    PORT MAP (
        A => S6355,
        B => S6359,
        Y => S6361
    );
NAND_3785: ENTITY WORK.NAND
    PORT MAP (
        A => S6356,
        B => S6360,
        Y => S6362
    );
NOR_2188: ENTITY WORK.NOR
    PORT MAP (
        A => S6352,
        B => S6362,
        Y => S6363
    );
NAND_3786: ENTITY WORK.NAND
    PORT MAP (
        A => S6351,
        B => S6361,
        Y => S6364
    );
NOR_2189: ENTITY WORK.NOR
    PORT MAP (
        A => S6351,
        B => S6361,
        Y => S6365
    );
NAND_3787: ENTITY WORK.NAND
    PORT MAP (
        A => S6352,
        B => S6362,
        Y => S6366
    );
NOR_2190: ENTITY WORK.NOR
    PORT MAP (
        A => S6363,
        B => S6365,
        Y => S6367
    );
NAND_3788: ENTITY WORK.NAND
    PORT MAP (
        A => S6364,
        B => S6366,
        Y => S6368
    );
NOR_2191: ENTITY WORK.NOR
    PORT MAP (
        A => S6268,
        B => S6272,
        Y => S6369
    );
NAND_3789: ENTITY WORK.NAND
    PORT MAP (
        A => S6269,
        B => S6273,
        Y => S6370
    );
NOR_2192: ENTITY WORK.NOR
    PORT MAP (
        A => S6368,
        B => S6369,
        Y => S6371
    );
NAND_3790: ENTITY WORK.NAND
    PORT MAP (
        A => S6367,
        B => S6370,
        Y => S6372
    );
NOR_2193: ENTITY WORK.NOR
    PORT MAP (
        A => S6367,
        B => S6370,
        Y => S6373
    );
NAND_3791: ENTITY WORK.NAND
    PORT MAP (
        A => S6368,
        B => S6369,
        Y => S6374
    );
NOR_2194: ENTITY WORK.NOR
    PORT MAP (
        A => S6371,
        B => S6373,
        Y => S6375
    );
NAND_3792: ENTITY WORK.NAND
    PORT MAP (
        A => S6372,
        B => S6374,
        Y => S6376
    );
NOR_2195: ENTITY WORK.NOR
    PORT MAP (
        A => S6247,
        B => S6376,
        Y => S6377
    );
NAND_3793: ENTITY WORK.NAND
    PORT MAP (
        A => S6246,
        B => S6375,
        Y => S6378
    );
NOR_2196: ENTITY WORK.NOR
    PORT MAP (
        A => S6246,
        B => S6375,
        Y => S6379
    );
NAND_3794: ENTITY WORK.NAND
    PORT MAP (
        A => S6247,
        B => S6376,
        Y => S6380
    );
NOR_2197: ENTITY WORK.NOR
    PORT MAP (
        A => S6377,
        B => S6379,
        Y => S6381
    );
NAND_3795: ENTITY WORK.NAND
    PORT MAP (
        A => S6378,
        B => S6380,
        Y => S6382
    );
NOR_2198: ENTITY WORK.NOR
    PORT MAP (
        A => S6298,
        B => S6304,
        Y => S6383
    );
NAND_3796: ENTITY WORK.NAND
    PORT MAP (
        A => S6299,
        B => S6305,
        Y => S6384
    );
NOR_2199: ENTITY WORK.NOR
    PORT MAP (
        A => S1065,
        B => S2107,
        Y => S6385
    );
NAND_3797: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_3,
        B => S2106,
        Y => S6386
    );
NOR_2200: ENTITY WORK.NOR
    PORT MAP (
        A => S963,
        B => S1953,
        Y => S6387
    );
NAND_3798: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_5,
        B => S1952,
        Y => S6388
    );
NOR_2201: ENTITY WORK.NOR
    PORT MAP (
        A => S6266,
        B => S6387,
        Y => S6389
    );
NAND_3799: ENTITY WORK.NAND
    PORT MAP (
        A => S6267,
        B => S6388,
        Y => S6390
    );
NOR_2202: ENTITY WORK.NOR
    PORT MAP (
        A => S963,
        B => S1598,
        Y => S6391
    );
NAND_3800: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_5,
        B => S1597,
        Y => S6392
    );
NOR_2203: ENTITY WORK.NOR
    PORT MAP (
        A => S6267,
        B => S6388,
        Y => S6393
    );
NAND_3801: ENTITY WORK.NAND
    PORT MAP (
        A => S6266,
        B => S6387,
        Y => S6394
    );
NOR_2204: ENTITY WORK.NOR
    PORT MAP (
        A => S6389,
        B => S6393,
        Y => S6395
    );
NAND_3802: ENTITY WORK.NAND
    PORT MAP (
        A => S6390,
        B => S6394,
        Y => S6396
    );
NOR_2205: ENTITY WORK.NOR
    PORT MAP (
        A => S6386,
        B => S6396,
        Y => S6397
    );
NAND_3803: ENTITY WORK.NAND
    PORT MAP (
        A => S6385,
        B => S6395,
        Y => S6398
    );
NOR_2206: ENTITY WORK.NOR
    PORT MAP (
        A => S6385,
        B => S6395,
        Y => S6399
    );
NAND_3804: ENTITY WORK.NAND
    PORT MAP (
        A => S6386,
        B => S6396,
        Y => S6400
    );
NOR_2207: ENTITY WORK.NOR
    PORT MAP (
        A => S6397,
        B => S6399,
        Y => S6401
    );
NAND_3805: ENTITY WORK.NAND
    PORT MAP (
        A => S6398,
        B => S6400,
        Y => S6402
    );
NOR_2208: ENTITY WORK.NOR
    PORT MAP (
        A => S6288,
        B => S6292,
        Y => S6403
    );
NAND_3806: ENTITY WORK.NAND
    PORT MAP (
        A => S6289,
        B => S6293,
        Y => S6404
    );
NOR_2209: ENTITY WORK.NOR
    PORT MAP (
        A => S910,
        B => S1849,
        Y => S6405
    );
NAND_3807: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_6,
        B => S1848,
        Y => S6406
    );
NOR_2210: ENTITY WORK.NOR
    PORT MAP (
        A => S805,
        B => S1516,
        Y => S6407
    );
NAND_3808: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_8,
        B => S1515,
        Y => S6408
    );
NOR_2211: ENTITY WORK.NOR
    PORT MAP (
        A => S6286,
        B => S6407,
        Y => S6409
    );
NAND_3809: ENTITY WORK.NAND
    PORT MAP (
        A => S6287,
        B => S6408,
        Y => S6410
    );
NOR_2212: ENTITY WORK.NOR
    PORT MAP (
        A => S805,
        B => S1746,
        Y => S6411
    );
NAND_3810: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_8,
        B => S1745,
        Y => S6412
    );
NOR_2213: ENTITY WORK.NOR
    PORT MAP (
        A => S6287,
        B => S6408,
        Y => S6413
    );
NAND_3811: ENTITY WORK.NAND
    PORT MAP (
        A => S6286,
        B => S6407,
        Y => S6414
    );
NOR_2214: ENTITY WORK.NOR
    PORT MAP (
        A => S6409,
        B => S6413,
        Y => S6415
    );
NAND_3812: ENTITY WORK.NAND
    PORT MAP (
        A => S6410,
        B => S6414,
        Y => S6416
    );
NOR_2215: ENTITY WORK.NOR
    PORT MAP (
        A => S6406,
        B => S6416,
        Y => S6417
    );
NAND_3813: ENTITY WORK.NAND
    PORT MAP (
        A => S6405,
        B => S6415,
        Y => S6418
    );
NOR_2216: ENTITY WORK.NOR
    PORT MAP (
        A => S6405,
        B => S6415,
        Y => S6419
    );
NAND_3814: ENTITY WORK.NAND
    PORT MAP (
        A => S6406,
        B => S6416,
        Y => S6420
    );
NOR_2217: ENTITY WORK.NOR
    PORT MAP (
        A => S6417,
        B => S6419,
        Y => S6421
    );
NAND_3815: ENTITY WORK.NAND
    PORT MAP (
        A => S6418,
        B => S6420,
        Y => S6422
    );
NOR_2218: ENTITY WORK.NOR
    PORT MAP (
        A => S6403,
        B => S6422,
        Y => S6423
    );
NAND_3816: ENTITY WORK.NAND
    PORT MAP (
        A => S6404,
        B => S6421,
        Y => S6424
    );
NOR_2219: ENTITY WORK.NOR
    PORT MAP (
        A => S6404,
        B => S6421,
        Y => S6425
    );
NAND_3817: ENTITY WORK.NAND
    PORT MAP (
        A => S6403,
        B => S6422,
        Y => S6426
    );
NOR_2220: ENTITY WORK.NOR
    PORT MAP (
        A => S6423,
        B => S6425,
        Y => S6427
    );
NAND_3818: ENTITY WORK.NAND
    PORT MAP (
        A => S6424,
        B => S6426,
        Y => S6428
    );
NOR_2221: ENTITY WORK.NOR
    PORT MAP (
        A => S6402,
        B => S6428,
        Y => S6429
    );
NAND_3819: ENTITY WORK.NAND
    PORT MAP (
        A => S6401,
        B => S6427,
        Y => S6430
    );
NOR_2222: ENTITY WORK.NOR
    PORT MAP (
        A => S6401,
        B => S6427,
        Y => S6431
    );
NAND_3820: ENTITY WORK.NAND
    PORT MAP (
        A => S6402,
        B => S6428,
        Y => S6432
    );
NOR_2223: ENTITY WORK.NOR
    PORT MAP (
        A => S6429,
        B => S6431,
        Y => S6433
    );
NAND_3821: ENTITY WORK.NAND
    PORT MAP (
        A => S6430,
        B => S6432,
        Y => S6434
    );
NOR_2224: ENTITY WORK.NOR
    PORT MAP (
        A => S6383,
        B => S6434,
        Y => S6435
    );
NAND_3822: ENTITY WORK.NAND
    PORT MAP (
        A => S6384,
        B => S6433,
        Y => S6436
    );
NOR_2225: ENTITY WORK.NOR
    PORT MAP (
        A => S6384,
        B => S6433,
        Y => S6437
    );
NAND_3823: ENTITY WORK.NAND
    PORT MAP (
        A => S6383,
        B => S6434,
        Y => S6438
    );
NOR_2226: ENTITY WORK.NOR
    PORT MAP (
        A => S6435,
        B => S6437,
        Y => S6439
    );
NAND_3824: ENTITY WORK.NAND
    PORT MAP (
        A => S6436,
        B => S6438,
        Y => S6440
    );
NOR_2227: ENTITY WORK.NOR
    PORT MAP (
        A => S6382,
        B => S6440,
        Y => S6441
    );
NAND_3825: ENTITY WORK.NAND
    PORT MAP (
        A => S6381,
        B => S6439,
        Y => S6442
    );
NOR_2228: ENTITY WORK.NOR
    PORT MAP (
        A => S6381,
        B => S6439,
        Y => S6443
    );
NAND_3826: ENTITY WORK.NAND
    PORT MAP (
        A => S6382,
        B => S6440,
        Y => S6444
    );
NOR_2229: ENTITY WORK.NOR
    PORT MAP (
        A => S6441,
        B => S6443,
        Y => S6445
    );
NAND_3827: ENTITY WORK.NAND
    PORT MAP (
        A => S6442,
        B => S6444,
        Y => S6446
    );
NOR_2230: ENTITY WORK.NOR
    PORT MAP (
        A => S6349,
        B => S6446,
        Y => S6447
    );
NAND_3828: ENTITY WORK.NAND
    PORT MAP (
        A => S6350,
        B => S6445,
        Y => S6448
    );
NOR_2231: ENTITY WORK.NOR
    PORT MAP (
        A => S6350,
        B => S6445,
        Y => S6449
    );
NAND_3829: ENTITY WORK.NAND
    PORT MAP (
        A => S6349,
        B => S6446,
        Y => S6450
    );
NOR_2232: ENTITY WORK.NOR
    PORT MAP (
        A => S6447,
        B => S6449,
        Y => S6451
    );
NAND_3830: ENTITY WORK.NAND
    PORT MAP (
        A => S6448,
        B => S6450,
        Y => S6452
    );
NOR_2233: ENTITY WORK.NOR
    PORT MAP (
        A => S6255,
        B => S6452,
        Y => S6453
    );
NAND_3831: ENTITY WORK.NAND
    PORT MAP (
        A => S6254,
        B => S6451,
        Y => S6454
    );
NOR_2234: ENTITY WORK.NOR
    PORT MAP (
        A => S6254,
        B => S6451,
        Y => S6455
    );
NAND_3832: ENTITY WORK.NAND
    PORT MAP (
        A => S6255,
        B => S6452,
        Y => S6456
    );
NOR_2235: ENTITY WORK.NOR
    PORT MAP (
        A => S6453,
        B => S6455,
        Y => S6457
    );
NAND_3833: ENTITY WORK.NAND
    PORT MAP (
        A => S6454,
        B => S6456,
        Y => S6458
    );
NAND_3834: ENTITY WORK.NAND
    PORT MAP (
        A => S6347,
        B => S6458,
        Y => S6459
    );
NOR_2236: ENTITY WORK.NOR
    PORT MAP (
        A => S6347,
        B => S6458,
        Y => S6460
    );
NAND_3835: ENTITY WORK.NAND
    PORT MAP (
        A => S6348,
        B => S6457,
        Y => S6461
    );
NAND_3836: ENTITY WORK.NAND
    PORT MAP (
        A => S6459,
        B => S6461,
        Y => S6462
    );
NOT_507: ENTITY WORK.NOT
    PORT MAP (
        A => S6462,
        Y => S6463
    );
NAND_3837: ENTITY WORK.NAND
    PORT MAP (
        A => S6333,
        B => S6463,
        Y => S6464
    );
NOT_508: ENTITY WORK.NOT
    PORT MAP (
        A => S6464,
        Y => S6465
    );
NAND_3838: ENTITY WORK.NAND
    PORT MAP (
        A => S6332,
        B => S6462,
        Y => S6466
    );
NAND_3839: ENTITY WORK.NAND
    PORT MAP (
        A => S6464,
        B => S6466,
        Y => S6467
    );
NOR_2237: ENTITY WORK.NOR
    PORT MAP (
        A => S6341,
        B => S6467,
        Y => S6468
    );
NOT_509: ENTITY WORK.NOT
    PORT MAP (
        A => S6468,
        Y => S6469
    );
NAND_3840: ENTITY WORK.NAND
    PORT MAP (
        A => S6341,
        B => S6467,
        Y => S6470
    );
NAND_3841: ENTITY WORK.NAND
    PORT MAP (
        A => S6469,
        B => S6470,
        Y => S6471
    );
NOR_2238: ENTITY WORK.NOR
    PORT MAP (
        A => S6337,
        B => S6471,
        Y => S6472
    );
NAND_3842: ENTITY WORK.NAND
    PORT MAP (
        A => S6337,
        B => S6471,
        Y => S6473
    );
NAND_3843: ENTITY WORK.NAND
    PORT MAP (
        A => S5948,
        B => S6473,
        Y => S6474
    );
NOR_2239: ENTITY WORK.NOR
    PORT MAP (
        A => S6472,
        B => S6474,
        Y => S6475
    );
NOR_2240: ENTITY WORK.NOR
    PORT MAP (
        A => S6345,
        B => S6475,
        Y => S6476
    );
NAND_3844: ENTITY WORK.NAND
    PORT MAP (
        A => S6346,
        B => S6476,
        Y => S290
    );
NOR_2241: ENTITY WORK.NOR
    PORT MAP (
        A => S3899,
        B => S4313,
        Y => S6477
    );
NAND_3845: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu1_9,
        B => S5950,
        Y => S6478
    );
NOR_2242: ENTITY WORK.NOR
    PORT MAP (
        A => S6468,
        B => S6472,
        Y => S6479
    );
NOR_2243: ENTITY WORK.NOR
    PORT MAP (
        A => S6447,
        B => S6453,
        Y => S6480
    );
NOR_2244: ENTITY WORK.NOR
    PORT MAP (
        A => S1220,
        B => S2518,
        Y => S6481
    );
NAND_3846: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_0,
        B => S2517,
        Y => S6482
    );
NOR_2245: ENTITY WORK.NOR
    PORT MAP (
        A => S6371,
        B => S6377,
        Y => S6483
    );
NAND_3847: ENTITY WORK.NAND
    PORT MAP (
        A => S6372,
        B => S6378,
        Y => S6484
    );
NOR_2246: ENTITY WORK.NOR
    PORT MAP (
        A => S6482,
        B => S6483,
        Y => S6485
    );
NOT_510: ENTITY WORK.NOT
    PORT MAP (
        A => S6485,
        Y => S6486
    );
NOR_2247: ENTITY WORK.NOR
    PORT MAP (
        A => S6481,
        B => S6484,
        Y => S6487
    );
NAND_3848: ENTITY WORK.NAND
    PORT MAP (
        A => S6482,
        B => S6483,
        Y => S6488
    );
NOR_2248: ENTITY WORK.NOR
    PORT MAP (
        A => S6485,
        B => S6487,
        Y => S6489
    );
NAND_3849: ENTITY WORK.NAND
    PORT MAP (
        A => S6486,
        B => S6488,
        Y => S6490
    );
NOR_2249: ENTITY WORK.NOR
    PORT MAP (
        A => S6435,
        B => S6441,
        Y => S6491
    );
NAND_3850: ENTITY WORK.NAND
    PORT MAP (
        A => S6436,
        B => S6442,
        Y => S6492
    );
NOR_2250: ENTITY WORK.NOR
    PORT MAP (
        A => S6359,
        B => S6363,
        Y => S6493
    );
NAND_3851: ENTITY WORK.NAND
    PORT MAP (
        A => S6360,
        B => S6364,
        Y => S6494
    );
NOR_2251: ENTITY WORK.NOR
    PORT MAP (
        A => S1168,
        B => S2418,
        Y => S6495
    );
NAND_3852: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_1,
        B => S2417,
        Y => S6496
    );
NOR_2252: ENTITY WORK.NOR
    PORT MAP (
        A => S1065,
        B => S2206,
        Y => S6497
    );
NAND_3853: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_3,
        B => S2205,
        Y => S6498
    );
NOR_2253: ENTITY WORK.NOR
    PORT MAP (
        A => S6357,
        B => S6497,
        Y => S6499
    );
NAND_3854: ENTITY WORK.NAND
    PORT MAP (
        A => S6358,
        B => S6498,
        Y => S6500
    );
NOR_2254: ENTITY WORK.NOR
    PORT MAP (
        A => S1065,
        B => S2312,
        Y => S6501
    );
NAND_3855: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_3,
        B => S2311,
        Y => S6502
    );
NOR_2255: ENTITY WORK.NOR
    PORT MAP (
        A => S6358,
        B => S6498,
        Y => S6503
    );
NAND_3856: ENTITY WORK.NAND
    PORT MAP (
        A => S6357,
        B => S6497,
        Y => S6504
    );
NOR_2256: ENTITY WORK.NOR
    PORT MAP (
        A => S6499,
        B => S6503,
        Y => S6505
    );
NAND_3857: ENTITY WORK.NAND
    PORT MAP (
        A => S6500,
        B => S6504,
        Y => S6506
    );
NOR_2257: ENTITY WORK.NOR
    PORT MAP (
        A => S6496,
        B => S6506,
        Y => S6507
    );
NAND_3858: ENTITY WORK.NAND
    PORT MAP (
        A => S6495,
        B => S6505,
        Y => S6508
    );
NOR_2258: ENTITY WORK.NOR
    PORT MAP (
        A => S6495,
        B => S6505,
        Y => S6509
    );
NAND_3859: ENTITY WORK.NAND
    PORT MAP (
        A => S6496,
        B => S6506,
        Y => S6510
    );
NOR_2259: ENTITY WORK.NOR
    PORT MAP (
        A => S6507,
        B => S6509,
        Y => S6511
    );
NAND_3860: ENTITY WORK.NAND
    PORT MAP (
        A => S6508,
        B => S6510,
        Y => S6512
    );
NOR_2260: ENTITY WORK.NOR
    PORT MAP (
        A => S6393,
        B => S6397,
        Y => S6513
    );
NAND_3861: ENTITY WORK.NAND
    PORT MAP (
        A => S6394,
        B => S6398,
        Y => S6514
    );
NOR_2261: ENTITY WORK.NOR
    PORT MAP (
        A => S6512,
        B => S6513,
        Y => S6515
    );
NAND_3862: ENTITY WORK.NAND
    PORT MAP (
        A => S6511,
        B => S6514,
        Y => S6516
    );
NOR_2262: ENTITY WORK.NOR
    PORT MAP (
        A => S6511,
        B => S6514,
        Y => S6517
    );
NAND_3863: ENTITY WORK.NAND
    PORT MAP (
        A => S6512,
        B => S6513,
        Y => S6518
    );
NOR_2263: ENTITY WORK.NOR
    PORT MAP (
        A => S6515,
        B => S6517,
        Y => S6519
    );
NAND_3864: ENTITY WORK.NAND
    PORT MAP (
        A => S6516,
        B => S6518,
        Y => S6520
    );
NOR_2264: ENTITY WORK.NOR
    PORT MAP (
        A => S6494,
        B => S6519,
        Y => S6521
    );
NAND_3865: ENTITY WORK.NAND
    PORT MAP (
        A => S6493,
        B => S6520,
        Y => S6522
    );
NOR_2265: ENTITY WORK.NOR
    PORT MAP (
        A => S6493,
        B => S6520,
        Y => S6523
    );
NAND_3866: ENTITY WORK.NAND
    PORT MAP (
        A => S6494,
        B => S6519,
        Y => S6524
    );
NOR_2266: ENTITY WORK.NOR
    PORT MAP (
        A => S6521,
        B => S6523,
        Y => S6525
    );
NAND_3867: ENTITY WORK.NAND
    PORT MAP (
        A => S6522,
        B => S6524,
        Y => S6526
    );
NOR_2267: ENTITY WORK.NOR
    PORT MAP (
        A => S6423,
        B => S6429,
        Y => S6527
    );
NAND_3868: ENTITY WORK.NAND
    PORT MAP (
        A => S6424,
        B => S6430,
        Y => S6528
    );
NOR_2268: ENTITY WORK.NOR
    PORT MAP (
        A => S1013,
        B => S2107,
        Y => S6529
    );
NAND_3869: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_4,
        B => S2106,
        Y => S6530
    );
NOR_2269: ENTITY WORK.NOR
    PORT MAP (
        A => S910,
        B => S1953,
        Y => S6531
    );
NAND_3870: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_6,
        B => S1952,
        Y => S6532
    );
NOR_2270: ENTITY WORK.NOR
    PORT MAP (
        A => S6391,
        B => S6531,
        Y => S6533
    );
NAND_3871: ENTITY WORK.NAND
    PORT MAP (
        A => S6392,
        B => S6532,
        Y => S6534
    );
NOR_2271: ENTITY WORK.NOR
    PORT MAP (
        A => S910,
        B => S1598,
        Y => S6535
    );
NAND_3872: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_6,
        B => S1597,
        Y => S6536
    );
NOR_2272: ENTITY WORK.NOR
    PORT MAP (
        A => S6392,
        B => S6532,
        Y => S6537
    );
NAND_3873: ENTITY WORK.NAND
    PORT MAP (
        A => S6391,
        B => S6531,
        Y => S6538
    );
NOR_2273: ENTITY WORK.NOR
    PORT MAP (
        A => S6533,
        B => S6537,
        Y => S6539
    );
NAND_3874: ENTITY WORK.NAND
    PORT MAP (
        A => S6534,
        B => S6538,
        Y => S6540
    );
NOR_2274: ENTITY WORK.NOR
    PORT MAP (
        A => S6530,
        B => S6540,
        Y => S6541
    );
NAND_3875: ENTITY WORK.NAND
    PORT MAP (
        A => S6529,
        B => S6539,
        Y => S6542
    );
NOR_2275: ENTITY WORK.NOR
    PORT MAP (
        A => S6529,
        B => S6539,
        Y => S6543
    );
NAND_3876: ENTITY WORK.NAND
    PORT MAP (
        A => S6530,
        B => S6540,
        Y => S6544
    );
NOR_2276: ENTITY WORK.NOR
    PORT MAP (
        A => S6541,
        B => S6543,
        Y => S6545
    );
NAND_3877: ENTITY WORK.NAND
    PORT MAP (
        A => S6542,
        B => S6544,
        Y => S6546
    );
NOR_2277: ENTITY WORK.NOR
    PORT MAP (
        A => S6413,
        B => S6417,
        Y => S6547
    );
NAND_3878: ENTITY WORK.NAND
    PORT MAP (
        A => S6414,
        B => S6418,
        Y => S6548
    );
NOR_2278: ENTITY WORK.NOR
    PORT MAP (
        A => S858,
        B => S1849,
        Y => S6549
    );
NAND_3879: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_7,
        B => S1848,
        Y => S6550
    );
NOR_2279: ENTITY WORK.NOR
    PORT MAP (
        A => S754,
        B => S1516,
        Y => S6551
    );
NAND_3880: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_9,
        B => S1515,
        Y => S6552
    );
NOR_2280: ENTITY WORK.NOR
    PORT MAP (
        A => S6411,
        B => S6551,
        Y => S6553
    );
NAND_3881: ENTITY WORK.NAND
    PORT MAP (
        A => S6412,
        B => S6552,
        Y => S6554
    );
NOR_2281: ENTITY WORK.NOR
    PORT MAP (
        A => S754,
        B => S1746,
        Y => S6555
    );
NAND_3882: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_9,
        B => S1745,
        Y => S6556
    );
NOR_2282: ENTITY WORK.NOR
    PORT MAP (
        A => S6412,
        B => S6552,
        Y => S6557
    );
NAND_3883: ENTITY WORK.NAND
    PORT MAP (
        A => S6411,
        B => S6551,
        Y => S6558
    );
NOR_2283: ENTITY WORK.NOR
    PORT MAP (
        A => S6553,
        B => S6557,
        Y => S6559
    );
NAND_3884: ENTITY WORK.NAND
    PORT MAP (
        A => S6554,
        B => S6558,
        Y => S6560
    );
NOR_2284: ENTITY WORK.NOR
    PORT MAP (
        A => S6550,
        B => S6560,
        Y => S6561
    );
NAND_3885: ENTITY WORK.NAND
    PORT MAP (
        A => S6549,
        B => S6559,
        Y => S6562
    );
NOR_2285: ENTITY WORK.NOR
    PORT MAP (
        A => S6549,
        B => S6559,
        Y => S6563
    );
NAND_3886: ENTITY WORK.NAND
    PORT MAP (
        A => S6550,
        B => S6560,
        Y => S6564
    );
NOR_2286: ENTITY WORK.NOR
    PORT MAP (
        A => S6561,
        B => S6563,
        Y => S6565
    );
NAND_3887: ENTITY WORK.NAND
    PORT MAP (
        A => S6562,
        B => S6564,
        Y => S6566
    );
NOR_2287: ENTITY WORK.NOR
    PORT MAP (
        A => S6547,
        B => S6566,
        Y => S6567
    );
NAND_3888: ENTITY WORK.NAND
    PORT MAP (
        A => S6548,
        B => S6565,
        Y => S6568
    );
NOR_2288: ENTITY WORK.NOR
    PORT MAP (
        A => S6548,
        B => S6565,
        Y => S6569
    );
NAND_3889: ENTITY WORK.NAND
    PORT MAP (
        A => S6547,
        B => S6566,
        Y => S6570
    );
NOR_2289: ENTITY WORK.NOR
    PORT MAP (
        A => S6567,
        B => S6569,
        Y => S6571
    );
NAND_3890: ENTITY WORK.NAND
    PORT MAP (
        A => S6568,
        B => S6570,
        Y => S6572
    );
NOR_2290: ENTITY WORK.NOR
    PORT MAP (
        A => S6546,
        B => S6572,
        Y => S6573
    );
NAND_3891: ENTITY WORK.NAND
    PORT MAP (
        A => S6545,
        B => S6571,
        Y => S6574
    );
NOR_2291: ENTITY WORK.NOR
    PORT MAP (
        A => S6545,
        B => S6571,
        Y => S6575
    );
NAND_3892: ENTITY WORK.NAND
    PORT MAP (
        A => S6546,
        B => S6572,
        Y => S6576
    );
NOR_2292: ENTITY WORK.NOR
    PORT MAP (
        A => S6573,
        B => S6575,
        Y => S6577
    );
NAND_3893: ENTITY WORK.NAND
    PORT MAP (
        A => S6574,
        B => S6576,
        Y => S6578
    );
NOR_2293: ENTITY WORK.NOR
    PORT MAP (
        A => S6527,
        B => S6578,
        Y => S6579
    );
NAND_3894: ENTITY WORK.NAND
    PORT MAP (
        A => S6528,
        B => S6577,
        Y => S6580
    );
NOR_2294: ENTITY WORK.NOR
    PORT MAP (
        A => S6528,
        B => S6577,
        Y => S6581
    );
NAND_3895: ENTITY WORK.NAND
    PORT MAP (
        A => S6527,
        B => S6578,
        Y => S6582
    );
NOR_2295: ENTITY WORK.NOR
    PORT MAP (
        A => S6579,
        B => S6581,
        Y => S6583
    );
NAND_3896: ENTITY WORK.NAND
    PORT MAP (
        A => S6580,
        B => S6582,
        Y => S6584
    );
NOR_2296: ENTITY WORK.NOR
    PORT MAP (
        A => S6526,
        B => S6584,
        Y => S6585
    );
NAND_3897: ENTITY WORK.NAND
    PORT MAP (
        A => S6525,
        B => S6583,
        Y => S6586
    );
NOR_2297: ENTITY WORK.NOR
    PORT MAP (
        A => S6525,
        B => S6583,
        Y => S6587
    );
NAND_3898: ENTITY WORK.NAND
    PORT MAP (
        A => S6526,
        B => S6584,
        Y => S6588
    );
NOR_2298: ENTITY WORK.NOR
    PORT MAP (
        A => S6585,
        B => S6587,
        Y => S6589
    );
NAND_3899: ENTITY WORK.NAND
    PORT MAP (
        A => S6586,
        B => S6588,
        Y => S6590
    );
NOR_2299: ENTITY WORK.NOR
    PORT MAP (
        A => S6491,
        B => S6590,
        Y => S6591
    );
NAND_3900: ENTITY WORK.NAND
    PORT MAP (
        A => S6492,
        B => S6589,
        Y => S6592
    );
NOR_2300: ENTITY WORK.NOR
    PORT MAP (
        A => S6492,
        B => S6589,
        Y => S6593
    );
NAND_3901: ENTITY WORK.NAND
    PORT MAP (
        A => S6491,
        B => S6590,
        Y => S6594
    );
NOR_2301: ENTITY WORK.NOR
    PORT MAP (
        A => S6591,
        B => S6593,
        Y => S6595
    );
NAND_3902: ENTITY WORK.NAND
    PORT MAP (
        A => S6592,
        B => S6594,
        Y => S6596
    );
NOR_2302: ENTITY WORK.NOR
    PORT MAP (
        A => S6490,
        B => S6596,
        Y => S6597
    );
NAND_3903: ENTITY WORK.NAND
    PORT MAP (
        A => S6489,
        B => S6595,
        Y => S6598
    );
NAND_3904: ENTITY WORK.NAND
    PORT MAP (
        A => S6490,
        B => S6596,
        Y => S6599
    );
NAND_3905: ENTITY WORK.NAND
    PORT MAP (
        A => S6598,
        B => S6599,
        Y => S6600
    );
NAND_3906: ENTITY WORK.NAND
    PORT MAP (
        A => S6480,
        B => S6600,
        Y => S6601
    );
NOT_511: ENTITY WORK.NOT
    PORT MAP (
        A => S6601,
        Y => S6602
    );
NOR_2303: ENTITY WORK.NOR
    PORT MAP (
        A => S6480,
        B => S6600,
        Y => S6603
    );
NOT_512: ENTITY WORK.NOT
    PORT MAP (
        A => S6603,
        Y => S6604
    );
NOR_2304: ENTITY WORK.NOR
    PORT MAP (
        A => S6602,
        B => S6603,
        Y => S6605
    );
NAND_3907: ENTITY WORK.NAND
    PORT MAP (
        A => S6601,
        B => S6604,
        Y => S6606
    );
NOR_2305: ENTITY WORK.NOR
    PORT MAP (
        A => S6461,
        B => S6606,
        Y => S6607
    );
NAND_3908: ENTITY WORK.NAND
    PORT MAP (
        A => S6460,
        B => S6605,
        Y => S6608
    );
NOR_2306: ENTITY WORK.NOR
    PORT MAP (
        A => S6460,
        B => S6605,
        Y => S6609
    );
NAND_3909: ENTITY WORK.NAND
    PORT MAP (
        A => S6461,
        B => S6606,
        Y => S6610
    );
NOR_2307: ENTITY WORK.NOR
    PORT MAP (
        A => S6607,
        B => S6609,
        Y => S6611
    );
NAND_3910: ENTITY WORK.NAND
    PORT MAP (
        A => S6608,
        B => S6610,
        Y => S6612
    );
NAND_3911: ENTITY WORK.NAND
    PORT MAP (
        A => S6465,
        B => S6611,
        Y => S6613
    );
NAND_3912: ENTITY WORK.NAND
    PORT MAP (
        A => S6464,
        B => S6612,
        Y => S6614
    );
NAND_3913: ENTITY WORK.NAND
    PORT MAP (
        A => S6613,
        B => S6614,
        Y => S6615
    );
NOR_2308: ENTITY WORK.NOR
    PORT MAP (
        A => S6479,
        B => S6615,
        Y => S6616
    );
NOT_513: ENTITY WORK.NOT
    PORT MAP (
        A => S6616,
        Y => S6617
    );
NAND_3914: ENTITY WORK.NAND
    PORT MAP (
        A => S6479,
        B => S6615,
        Y => S6618
    );
NAND_3915: ENTITY WORK.NAND
    PORT MAP (
        A => S5948,
        B => S6618,
        Y => S6619
    );
NOR_2309: ENTITY WORK.NOR
    PORT MAP (
        A => S6616,
        B => S6619,
        Y => S6620
    );
NOR_2310: ENTITY WORK.NOR
    PORT MAP (
        A => S6477,
        B => S6620,
        Y => S6621
    );
NAND_3916: ENTITY WORK.NAND
    PORT MAP (
        A => S6478,
        B => S6621,
        Y => S291
    );
NOR_2311: ENTITY WORK.NOR
    PORT MAP (
        A => S3899,
        B => S4195,
        Y => S6622
    );
NAND_3917: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu1_10,
        B => S5950,
        Y => S6623
    );
NAND_3918: ENTITY WORK.NAND
    PORT MAP (
        A => S6613,
        B => S6617,
        Y => S6624
    );
NOR_2312: ENTITY WORK.NOR
    PORT MAP (
        A => S6591,
        B => S6597,
        Y => S6625
    );
NAND_3919: ENTITY WORK.NAND
    PORT MAP (
        A => S6592,
        B => S6598,
        Y => S6626
    );
NOR_2313: ENTITY WORK.NOR
    PORT MAP (
        A => S1220,
        B => S2618,
        Y => S6627
    );
NAND_3920: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_0,
        B => S2617,
        Y => S6628
    );
NOR_2314: ENTITY WORK.NOR
    PORT MAP (
        A => S1168,
        B => S2518,
        Y => S6629
    );
NAND_3921: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_1,
        B => S2517,
        Y => S6630
    );
NOR_2315: ENTITY WORK.NOR
    PORT MAP (
        A => S6627,
        B => S6629,
        Y => S6631
    );
NAND_3922: ENTITY WORK.NAND
    PORT MAP (
        A => S6628,
        B => S6630,
        Y => S6632
    );
NOR_2316: ENTITY WORK.NOR
    PORT MAP (
        A => S1168,
        B => S2618,
        Y => S6633
    );
NAND_3923: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_1,
        B => S2617,
        Y => S6634
    );
NOR_2317: ENTITY WORK.NOR
    PORT MAP (
        A => S6482,
        B => S6634,
        Y => S6635
    );
NAND_3924: ENTITY WORK.NAND
    PORT MAP (
        A => S6481,
        B => S6633,
        Y => S6636
    );
NOR_2318: ENTITY WORK.NOR
    PORT MAP (
        A => S6631,
        B => S6635,
        Y => S6637
    );
NAND_3925: ENTITY WORK.NAND
    PORT MAP (
        A => S6632,
        B => S6636,
        Y => S6638
    );
NOR_2319: ENTITY WORK.NOR
    PORT MAP (
        A => S6515,
        B => S6523,
        Y => S6639
    );
NAND_3926: ENTITY WORK.NAND
    PORT MAP (
        A => S6516,
        B => S6524,
        Y => S6640
    );
NOR_2320: ENTITY WORK.NOR
    PORT MAP (
        A => S6637,
        B => S6640,
        Y => S6641
    );
NAND_3927: ENTITY WORK.NAND
    PORT MAP (
        A => S6638,
        B => S6639,
        Y => S6642
    );
NOR_2321: ENTITY WORK.NOR
    PORT MAP (
        A => S6638,
        B => S6639,
        Y => S6643
    );
NAND_3928: ENTITY WORK.NAND
    PORT MAP (
        A => S6637,
        B => S6640,
        Y => S6644
    );
NOR_2322: ENTITY WORK.NOR
    PORT MAP (
        A => S6641,
        B => S6643,
        Y => S6645
    );
NAND_3929: ENTITY WORK.NAND
    PORT MAP (
        A => S6642,
        B => S6644,
        Y => S6646
    );
NOR_2323: ENTITY WORK.NOR
    PORT MAP (
        A => S6579,
        B => S6585,
        Y => S6647
    );
NAND_3930: ENTITY WORK.NAND
    PORT MAP (
        A => S6580,
        B => S6586,
        Y => S6648
    );
NOR_2324: ENTITY WORK.NOR
    PORT MAP (
        A => S6503,
        B => S6507,
        Y => S6649
    );
NAND_3931: ENTITY WORK.NAND
    PORT MAP (
        A => S6504,
        B => S6508,
        Y => S6650
    );
NOR_2325: ENTITY WORK.NOR
    PORT MAP (
        A => S1116,
        B => S2418,
        Y => S6651
    );
NAND_3932: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_2,
        B => S2417,
        Y => S6652
    );
NOR_2326: ENTITY WORK.NOR
    PORT MAP (
        A => S1013,
        B => S2206,
        Y => S6653
    );
NAND_3933: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_4,
        B => S2205,
        Y => S6654
    );
NOR_2327: ENTITY WORK.NOR
    PORT MAP (
        A => S6501,
        B => S6653,
        Y => S6655
    );
NAND_3934: ENTITY WORK.NAND
    PORT MAP (
        A => S6502,
        B => S6654,
        Y => S6656
    );
NOR_2328: ENTITY WORK.NOR
    PORT MAP (
        A => S1013,
        B => S2312,
        Y => S6657
    );
NAND_3935: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_4,
        B => S2311,
        Y => S6658
    );
NOR_2329: ENTITY WORK.NOR
    PORT MAP (
        A => S6502,
        B => S6654,
        Y => S6659
    );
NAND_3936: ENTITY WORK.NAND
    PORT MAP (
        A => S6501,
        B => S6653,
        Y => S6660
    );
NOR_2330: ENTITY WORK.NOR
    PORT MAP (
        A => S6655,
        B => S6659,
        Y => S6661
    );
NAND_3937: ENTITY WORK.NAND
    PORT MAP (
        A => S6656,
        B => S6660,
        Y => S6662
    );
NOR_2331: ENTITY WORK.NOR
    PORT MAP (
        A => S6652,
        B => S6662,
        Y => S6663
    );
NAND_3938: ENTITY WORK.NAND
    PORT MAP (
        A => S6651,
        B => S6661,
        Y => S6664
    );
NOR_2332: ENTITY WORK.NOR
    PORT MAP (
        A => S6651,
        B => S6661,
        Y => S6665
    );
NAND_3939: ENTITY WORK.NAND
    PORT MAP (
        A => S6652,
        B => S6662,
        Y => S6666
    );
NOR_2333: ENTITY WORK.NOR
    PORT MAP (
        A => S6663,
        B => S6665,
        Y => S6667
    );
NAND_3940: ENTITY WORK.NAND
    PORT MAP (
        A => S6664,
        B => S6666,
        Y => S6668
    );
NOR_2334: ENTITY WORK.NOR
    PORT MAP (
        A => S6537,
        B => S6541,
        Y => S6669
    );
NAND_3941: ENTITY WORK.NAND
    PORT MAP (
        A => S6538,
        B => S6542,
        Y => S6670
    );
NOR_2335: ENTITY WORK.NOR
    PORT MAP (
        A => S6668,
        B => S6669,
        Y => S6671
    );
NAND_3942: ENTITY WORK.NAND
    PORT MAP (
        A => S6667,
        B => S6670,
        Y => S6672
    );
NOR_2336: ENTITY WORK.NOR
    PORT MAP (
        A => S6667,
        B => S6670,
        Y => S6673
    );
NAND_3943: ENTITY WORK.NAND
    PORT MAP (
        A => S6668,
        B => S6669,
        Y => S6674
    );
NOR_2337: ENTITY WORK.NOR
    PORT MAP (
        A => S6671,
        B => S6673,
        Y => S6675
    );
NAND_3944: ENTITY WORK.NAND
    PORT MAP (
        A => S6672,
        B => S6674,
        Y => S6676
    );
NOR_2338: ENTITY WORK.NOR
    PORT MAP (
        A => S6650,
        B => S6675,
        Y => S6677
    );
NAND_3945: ENTITY WORK.NAND
    PORT MAP (
        A => S6649,
        B => S6676,
        Y => S6678
    );
NOR_2339: ENTITY WORK.NOR
    PORT MAP (
        A => S6649,
        B => S6676,
        Y => S6679
    );
NAND_3946: ENTITY WORK.NAND
    PORT MAP (
        A => S6650,
        B => S6675,
        Y => S6680
    );
NOR_2340: ENTITY WORK.NOR
    PORT MAP (
        A => S6677,
        B => S6679,
        Y => S6681
    );
NAND_3947: ENTITY WORK.NAND
    PORT MAP (
        A => S6678,
        B => S6680,
        Y => S6682
    );
NOR_2341: ENTITY WORK.NOR
    PORT MAP (
        A => S6567,
        B => S6573,
        Y => S6683
    );
NAND_3948: ENTITY WORK.NAND
    PORT MAP (
        A => S6568,
        B => S6574,
        Y => S6684
    );
NOR_2342: ENTITY WORK.NOR
    PORT MAP (
        A => S963,
        B => S2107,
        Y => S6685
    );
NAND_3949: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_5,
        B => S2106,
        Y => S6686
    );
NOR_2343: ENTITY WORK.NOR
    PORT MAP (
        A => S858,
        B => S1953,
        Y => S6687
    );
NAND_3950: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_7,
        B => S1952,
        Y => S6688
    );
NOR_2344: ENTITY WORK.NOR
    PORT MAP (
        A => S6535,
        B => S6687,
        Y => S6689
    );
NAND_3951: ENTITY WORK.NAND
    PORT MAP (
        A => S6536,
        B => S6688,
        Y => S6690
    );
NOR_2345: ENTITY WORK.NOR
    PORT MAP (
        A => S858,
        B => S1598,
        Y => S6691
    );
NAND_3952: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_7,
        B => S1597,
        Y => S6692
    );
NOR_2346: ENTITY WORK.NOR
    PORT MAP (
        A => S6536,
        B => S6688,
        Y => S6693
    );
NAND_3953: ENTITY WORK.NAND
    PORT MAP (
        A => S6535,
        B => S6687,
        Y => S6694
    );
NOR_2347: ENTITY WORK.NOR
    PORT MAP (
        A => S6689,
        B => S6693,
        Y => S6695
    );
NAND_3954: ENTITY WORK.NAND
    PORT MAP (
        A => S6690,
        B => S6694,
        Y => S6696
    );
NOR_2348: ENTITY WORK.NOR
    PORT MAP (
        A => S6686,
        B => S6696,
        Y => S6697
    );
NAND_3955: ENTITY WORK.NAND
    PORT MAP (
        A => S6685,
        B => S6695,
        Y => S6698
    );
NOR_2349: ENTITY WORK.NOR
    PORT MAP (
        A => S6685,
        B => S6695,
        Y => S6699
    );
NAND_3956: ENTITY WORK.NAND
    PORT MAP (
        A => S6686,
        B => S6696,
        Y => S6700
    );
NOR_2350: ENTITY WORK.NOR
    PORT MAP (
        A => S6697,
        B => S6699,
        Y => S6701
    );
NAND_3957: ENTITY WORK.NAND
    PORT MAP (
        A => S6698,
        B => S6700,
        Y => S6702
    );
NOR_2351: ENTITY WORK.NOR
    PORT MAP (
        A => S6557,
        B => S6561,
        Y => S6703
    );
NAND_3958: ENTITY WORK.NAND
    PORT MAP (
        A => S6558,
        B => S6562,
        Y => S6704
    );
NOR_2352: ENTITY WORK.NOR
    PORT MAP (
        A => S805,
        B => S1849,
        Y => S6705
    );
NAND_3959: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_8,
        B => S1848,
        Y => S6706
    );
NOR_2353: ENTITY WORK.NOR
    PORT MAP (
        A => S702,
        B => S1516,
        Y => S6707
    );
NAND_3960: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_10,
        B => S1515,
        Y => S6708
    );
NOR_2354: ENTITY WORK.NOR
    PORT MAP (
        A => S6555,
        B => S6707,
        Y => S6709
    );
NAND_3961: ENTITY WORK.NAND
    PORT MAP (
        A => S6556,
        B => S6708,
        Y => S6710
    );
NOR_2355: ENTITY WORK.NOR
    PORT MAP (
        A => S702,
        B => S1746,
        Y => S6711
    );
NAND_3962: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_10,
        B => S1745,
        Y => S6712
    );
NOR_2356: ENTITY WORK.NOR
    PORT MAP (
        A => S6556,
        B => S6708,
        Y => S6713
    );
NAND_3963: ENTITY WORK.NAND
    PORT MAP (
        A => S6555,
        B => S6707,
        Y => S6714
    );
NOR_2357: ENTITY WORK.NOR
    PORT MAP (
        A => S6709,
        B => S6713,
        Y => S6715
    );
NAND_3964: ENTITY WORK.NAND
    PORT MAP (
        A => S6710,
        B => S6714,
        Y => S6716
    );
NOR_2358: ENTITY WORK.NOR
    PORT MAP (
        A => S6706,
        B => S6716,
        Y => S6717
    );
NAND_3965: ENTITY WORK.NAND
    PORT MAP (
        A => S6705,
        B => S6715,
        Y => S6718
    );
NOR_2359: ENTITY WORK.NOR
    PORT MAP (
        A => S6705,
        B => S6715,
        Y => S6719
    );
NAND_3966: ENTITY WORK.NAND
    PORT MAP (
        A => S6706,
        B => S6716,
        Y => S6720
    );
NOR_2360: ENTITY WORK.NOR
    PORT MAP (
        A => S6717,
        B => S6719,
        Y => S6721
    );
NAND_3967: ENTITY WORK.NAND
    PORT MAP (
        A => S6718,
        B => S6720,
        Y => S6722
    );
NOR_2361: ENTITY WORK.NOR
    PORT MAP (
        A => S6703,
        B => S6722,
        Y => S6723
    );
NAND_3968: ENTITY WORK.NAND
    PORT MAP (
        A => S6704,
        B => S6721,
        Y => S6724
    );
NOR_2362: ENTITY WORK.NOR
    PORT MAP (
        A => S6704,
        B => S6721,
        Y => S6725
    );
NAND_3969: ENTITY WORK.NAND
    PORT MAP (
        A => S6703,
        B => S6722,
        Y => S6726
    );
NOR_2363: ENTITY WORK.NOR
    PORT MAP (
        A => S6723,
        B => S6725,
        Y => S6727
    );
NAND_3970: ENTITY WORK.NAND
    PORT MAP (
        A => S6724,
        B => S6726,
        Y => S6728
    );
NOR_2364: ENTITY WORK.NOR
    PORT MAP (
        A => S6702,
        B => S6728,
        Y => S6729
    );
NAND_3971: ENTITY WORK.NAND
    PORT MAP (
        A => S6701,
        B => S6727,
        Y => S6730
    );
NOR_2365: ENTITY WORK.NOR
    PORT MAP (
        A => S6701,
        B => S6727,
        Y => S6731
    );
NAND_3972: ENTITY WORK.NAND
    PORT MAP (
        A => S6702,
        B => S6728,
        Y => S6732
    );
NOR_2366: ENTITY WORK.NOR
    PORT MAP (
        A => S6729,
        B => S6731,
        Y => S6733
    );
NAND_3973: ENTITY WORK.NAND
    PORT MAP (
        A => S6730,
        B => S6732,
        Y => S6734
    );
NOR_2367: ENTITY WORK.NOR
    PORT MAP (
        A => S6683,
        B => S6734,
        Y => S6735
    );
NAND_3974: ENTITY WORK.NAND
    PORT MAP (
        A => S6684,
        B => S6733,
        Y => S6736
    );
NOR_2368: ENTITY WORK.NOR
    PORT MAP (
        A => S6684,
        B => S6733,
        Y => S6737
    );
NAND_3975: ENTITY WORK.NAND
    PORT MAP (
        A => S6683,
        B => S6734,
        Y => S6738
    );
NOR_2369: ENTITY WORK.NOR
    PORT MAP (
        A => S6735,
        B => S6737,
        Y => S6739
    );
NAND_3976: ENTITY WORK.NAND
    PORT MAP (
        A => S6736,
        B => S6738,
        Y => S6740
    );
NOR_2370: ENTITY WORK.NOR
    PORT MAP (
        A => S6682,
        B => S6740,
        Y => S6741
    );
NAND_3977: ENTITY WORK.NAND
    PORT MAP (
        A => S6681,
        B => S6739,
        Y => S6742
    );
NOR_2371: ENTITY WORK.NOR
    PORT MAP (
        A => S6681,
        B => S6739,
        Y => S6743
    );
NAND_3978: ENTITY WORK.NAND
    PORT MAP (
        A => S6682,
        B => S6740,
        Y => S6744
    );
NOR_2372: ENTITY WORK.NOR
    PORT MAP (
        A => S6741,
        B => S6743,
        Y => S6745
    );
NAND_3979: ENTITY WORK.NAND
    PORT MAP (
        A => S6742,
        B => S6744,
        Y => S6746
    );
NOR_2373: ENTITY WORK.NOR
    PORT MAP (
        A => S6647,
        B => S6746,
        Y => S6747
    );
NAND_3980: ENTITY WORK.NAND
    PORT MAP (
        A => S6648,
        B => S6745,
        Y => S6748
    );
NOR_2374: ENTITY WORK.NOR
    PORT MAP (
        A => S6648,
        B => S6745,
        Y => S6749
    );
NAND_3981: ENTITY WORK.NAND
    PORT MAP (
        A => S6647,
        B => S6746,
        Y => S6750
    );
NOR_2375: ENTITY WORK.NOR
    PORT MAP (
        A => S6747,
        B => S6749,
        Y => S6751
    );
NAND_3982: ENTITY WORK.NAND
    PORT MAP (
        A => S6748,
        B => S6750,
        Y => S6752
    );
NOR_2376: ENTITY WORK.NOR
    PORT MAP (
        A => S6646,
        B => S6752,
        Y => S6753
    );
NAND_3983: ENTITY WORK.NAND
    PORT MAP (
        A => S6645,
        B => S6751,
        Y => S6754
    );
NOR_2377: ENTITY WORK.NOR
    PORT MAP (
        A => S6645,
        B => S6751,
        Y => S6755
    );
NAND_3984: ENTITY WORK.NAND
    PORT MAP (
        A => S6646,
        B => S6752,
        Y => S6756
    );
NOR_2378: ENTITY WORK.NOR
    PORT MAP (
        A => S6753,
        B => S6755,
        Y => S6757
    );
NAND_3985: ENTITY WORK.NAND
    PORT MAP (
        A => S6754,
        B => S6756,
        Y => S6758
    );
NOR_2379: ENTITY WORK.NOR
    PORT MAP (
        A => S6625,
        B => S6758,
        Y => S6759
    );
NAND_3986: ENTITY WORK.NAND
    PORT MAP (
        A => S6626,
        B => S6757,
        Y => S6760
    );
NOR_2380: ENTITY WORK.NOR
    PORT MAP (
        A => S6626,
        B => S6757,
        Y => S6761
    );
NOR_2381: ENTITY WORK.NOR
    PORT MAP (
        A => S6759,
        B => S6761,
        Y => S6762
    );
NOT_514: ENTITY WORK.NOT
    PORT MAP (
        A => S6762,
        Y => S6763
    );
NOR_2382: ENTITY WORK.NOR
    PORT MAP (
        A => S6486,
        B => S6763,
        Y => S6764
    );
NOT_515: ENTITY WORK.NOT
    PORT MAP (
        A => S6764,
        Y => S6765
    );
NOR_2383: ENTITY WORK.NOR
    PORT MAP (
        A => S6485,
        B => S6762,
        Y => S6766
    );
NOR_2384: ENTITY WORK.NOR
    PORT MAP (
        A => S6764,
        B => S6766,
        Y => S6767
    );
NAND_3987: ENTITY WORK.NAND
    PORT MAP (
        A => S6603,
        B => S6767,
        Y => S6768
    );
NOT_516: ENTITY WORK.NOT
    PORT MAP (
        A => S6768,
        Y => S6769
    );
NOR_2385: ENTITY WORK.NOR
    PORT MAP (
        A => S6603,
        B => S6767,
        Y => S6770
    );
NOT_517: ENTITY WORK.NOT
    PORT MAP (
        A => S6770,
        Y => S6771
    );
NOR_2386: ENTITY WORK.NOR
    PORT MAP (
        A => S6769,
        B => S6770,
        Y => S6772
    );
NAND_3988: ENTITY WORK.NAND
    PORT MAP (
        A => S6768,
        B => S6771,
        Y => S6773
    );
NOR_2387: ENTITY WORK.NOR
    PORT MAP (
        A => S6608,
        B => S6773,
        Y => S6774
    );
NOR_2388: ENTITY WORK.NOR
    PORT MAP (
        A => S6607,
        B => S6772,
        Y => S6775
    );
NOR_2389: ENTITY WORK.NOR
    PORT MAP (
        A => S6774,
        B => S6775,
        Y => S6776
    );
NAND_3989: ENTITY WORK.NAND
    PORT MAP (
        A => S6624,
        B => S6776,
        Y => S6777
    );
NOT_518: ENTITY WORK.NOT
    PORT MAP (
        A => S6777,
        Y => S6778
    );
NOR_2390: ENTITY WORK.NOR
    PORT MAP (
        A => S6624,
        B => S6776,
        Y => S6779
    );
NAND_3990: ENTITY WORK.NAND
    PORT MAP (
        A => S5948,
        B => S6777,
        Y => S6780
    );
NOR_2391: ENTITY WORK.NOR
    PORT MAP (
        A => S6779,
        B => S6780,
        Y => S6781
    );
NOR_2392: ENTITY WORK.NOR
    PORT MAP (
        A => S6622,
        B => S6781,
        Y => S6782
    );
NAND_3991: ENTITY WORK.NAND
    PORT MAP (
        A => S6623,
        B => S6782,
        Y => S292
    );
NOR_2393: ENTITY WORK.NOR
    PORT MAP (
        A => S3899,
        B => S4108,
        Y => S6783
    );
NAND_3992: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu1_11,
        B => S5950,
        Y => S6784
    );
NOR_2394: ENTITY WORK.NOR
    PORT MAP (
        A => S6774,
        B => S6778,
        Y => S6785
    );
NOR_2395: ENTITY WORK.NOR
    PORT MAP (
        A => S6759,
        B => S6764,
        Y => S6786
    );
NAND_3993: ENTITY WORK.NAND
    PORT MAP (
        A => S6760,
        B => S6765,
        Y => S6787
    );
NOR_2396: ENTITY WORK.NOR
    PORT MAP (
        A => S6747,
        B => S6753,
        Y => S6788
    );
NAND_3994: ENTITY WORK.NAND
    PORT MAP (
        A => S6748,
        B => S6754,
        Y => S6789
    );
NOR_2397: ENTITY WORK.NOR
    PORT MAP (
        A => S1220,
        B => S2718,
        Y => S6790
    );
NAND_3995: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_0,
        B => S2717,
        Y => S6791
    );
NOR_2398: ENTITY WORK.NOR
    PORT MAP (
        A => S1116,
        B => S2518,
        Y => S6792
    );
NAND_3996: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_2,
        B => S2517,
        Y => S6793
    );
NOR_2399: ENTITY WORK.NOR
    PORT MAP (
        A => S6633,
        B => S6792,
        Y => S6794
    );
NAND_3997: ENTITY WORK.NAND
    PORT MAP (
        A => S6634,
        B => S6793,
        Y => S6795
    );
NOR_2400: ENTITY WORK.NOR
    PORT MAP (
        A => S1116,
        B => S2618,
        Y => S6796
    );
NAND_3998: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_2,
        B => S2617,
        Y => S6797
    );
NOR_2401: ENTITY WORK.NOR
    PORT MAP (
        A => S6634,
        B => S6793,
        Y => S6798
    );
NAND_3999: ENTITY WORK.NAND
    PORT MAP (
        A => S6633,
        B => S6792,
        Y => S6799
    );
NOR_2402: ENTITY WORK.NOR
    PORT MAP (
        A => S6794,
        B => S6798,
        Y => S6800
    );
NAND_4000: ENTITY WORK.NAND
    PORT MAP (
        A => S6795,
        B => S6799,
        Y => S6801
    );
NOR_2403: ENTITY WORK.NOR
    PORT MAP (
        A => S6791,
        B => S6801,
        Y => S6802
    );
NAND_4001: ENTITY WORK.NAND
    PORT MAP (
        A => S6790,
        B => S6800,
        Y => S6803
    );
NOR_2404: ENTITY WORK.NOR
    PORT MAP (
        A => S6790,
        B => S6800,
        Y => S6804
    );
NAND_4002: ENTITY WORK.NAND
    PORT MAP (
        A => S6791,
        B => S6801,
        Y => S6805
    );
NOR_2405: ENTITY WORK.NOR
    PORT MAP (
        A => S6802,
        B => S6804,
        Y => S6806
    );
NAND_4003: ENTITY WORK.NAND
    PORT MAP (
        A => S6803,
        B => S6805,
        Y => S6807
    );
NOR_2406: ENTITY WORK.NOR
    PORT MAP (
        A => S6636,
        B => S6807,
        Y => S6808
    );
NAND_4004: ENTITY WORK.NAND
    PORT MAP (
        A => S6635,
        B => S6806,
        Y => S6809
    );
NOR_2407: ENTITY WORK.NOR
    PORT MAP (
        A => S6635,
        B => S6806,
        Y => S6810
    );
NAND_4005: ENTITY WORK.NAND
    PORT MAP (
        A => S6636,
        B => S6807,
        Y => S6811
    );
NOR_2408: ENTITY WORK.NOR
    PORT MAP (
        A => S6808,
        B => S6810,
        Y => S6812
    );
NAND_4006: ENTITY WORK.NAND
    PORT MAP (
        A => S6809,
        B => S6811,
        Y => S6813
    );
NOR_2409: ENTITY WORK.NOR
    PORT MAP (
        A => S6671,
        B => S6679,
        Y => S6814
    );
NAND_4007: ENTITY WORK.NAND
    PORT MAP (
        A => S6672,
        B => S6680,
        Y => S6815
    );
NOR_2410: ENTITY WORK.NOR
    PORT MAP (
        A => S6812,
        B => S6815,
        Y => S6816
    );
NAND_4008: ENTITY WORK.NAND
    PORT MAP (
        A => S6813,
        B => S6814,
        Y => S6817
    );
NOR_2411: ENTITY WORK.NOR
    PORT MAP (
        A => S6813,
        B => S6814,
        Y => S6818
    );
NAND_4009: ENTITY WORK.NAND
    PORT MAP (
        A => S6812,
        B => S6815,
        Y => S6819
    );
NOR_2412: ENTITY WORK.NOR
    PORT MAP (
        A => S6816,
        B => S6818,
        Y => S6820
    );
NAND_4010: ENTITY WORK.NAND
    PORT MAP (
        A => S6817,
        B => S6819,
        Y => S6821
    );
NOR_2413: ENTITY WORK.NOR
    PORT MAP (
        A => S6735,
        B => S6741,
        Y => S6822
    );
NAND_4011: ENTITY WORK.NAND
    PORT MAP (
        A => S6736,
        B => S6742,
        Y => S6823
    );
NOR_2414: ENTITY WORK.NOR
    PORT MAP (
        A => S6659,
        B => S6663,
        Y => S6824
    );
NAND_4012: ENTITY WORK.NAND
    PORT MAP (
        A => S6660,
        B => S6664,
        Y => S6825
    );
NOR_2415: ENTITY WORK.NOR
    PORT MAP (
        A => S1065,
        B => S2418,
        Y => S6826
    );
NAND_4013: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_3,
        B => S2417,
        Y => S6827
    );
NOR_2416: ENTITY WORK.NOR
    PORT MAP (
        A => S963,
        B => S2206,
        Y => S6828
    );
NAND_4014: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_5,
        B => S2205,
        Y => S6829
    );
NOR_2417: ENTITY WORK.NOR
    PORT MAP (
        A => S6657,
        B => S6828,
        Y => S6830
    );
NAND_4015: ENTITY WORK.NAND
    PORT MAP (
        A => S6658,
        B => S6829,
        Y => S6831
    );
NOR_2418: ENTITY WORK.NOR
    PORT MAP (
        A => S963,
        B => S2312,
        Y => S6832
    );
NAND_4016: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_5,
        B => S2311,
        Y => S6833
    );
NOR_2419: ENTITY WORK.NOR
    PORT MAP (
        A => S6658,
        B => S6829,
        Y => S6834
    );
NAND_4017: ENTITY WORK.NAND
    PORT MAP (
        A => S6657,
        B => S6828,
        Y => S6835
    );
NOR_2420: ENTITY WORK.NOR
    PORT MAP (
        A => S6830,
        B => S6834,
        Y => S6836
    );
NAND_4018: ENTITY WORK.NAND
    PORT MAP (
        A => S6831,
        B => S6835,
        Y => S6837
    );
NOR_2421: ENTITY WORK.NOR
    PORT MAP (
        A => S6827,
        B => S6837,
        Y => S6838
    );
NAND_4019: ENTITY WORK.NAND
    PORT MAP (
        A => S6826,
        B => S6836,
        Y => S6839
    );
NOR_2422: ENTITY WORK.NOR
    PORT MAP (
        A => S6826,
        B => S6836,
        Y => S6840
    );
NAND_4020: ENTITY WORK.NAND
    PORT MAP (
        A => S6827,
        B => S6837,
        Y => S6841
    );
NOR_2423: ENTITY WORK.NOR
    PORT MAP (
        A => S6838,
        B => S6840,
        Y => S6842
    );
NAND_4021: ENTITY WORK.NAND
    PORT MAP (
        A => S6839,
        B => S6841,
        Y => S6843
    );
NOR_2424: ENTITY WORK.NOR
    PORT MAP (
        A => S6693,
        B => S6697,
        Y => S6844
    );
NAND_4022: ENTITY WORK.NAND
    PORT MAP (
        A => S6694,
        B => S6698,
        Y => S6845
    );
NOR_2425: ENTITY WORK.NOR
    PORT MAP (
        A => S6843,
        B => S6844,
        Y => S6846
    );
NAND_4023: ENTITY WORK.NAND
    PORT MAP (
        A => S6842,
        B => S6845,
        Y => S6847
    );
NOR_2426: ENTITY WORK.NOR
    PORT MAP (
        A => S6842,
        B => S6845,
        Y => S6848
    );
NAND_4024: ENTITY WORK.NAND
    PORT MAP (
        A => S6843,
        B => S6844,
        Y => S6849
    );
NOR_2427: ENTITY WORK.NOR
    PORT MAP (
        A => S6846,
        B => S6848,
        Y => S6850
    );
NAND_4025: ENTITY WORK.NAND
    PORT MAP (
        A => S6847,
        B => S6849,
        Y => S6851
    );
NOR_2428: ENTITY WORK.NOR
    PORT MAP (
        A => S6825,
        B => S6850,
        Y => S6852
    );
NAND_4026: ENTITY WORK.NAND
    PORT MAP (
        A => S6824,
        B => S6851,
        Y => S6853
    );
NOR_2429: ENTITY WORK.NOR
    PORT MAP (
        A => S6824,
        B => S6851,
        Y => S6854
    );
NAND_4027: ENTITY WORK.NAND
    PORT MAP (
        A => S6825,
        B => S6850,
        Y => S6855
    );
NOR_2430: ENTITY WORK.NOR
    PORT MAP (
        A => S6852,
        B => S6854,
        Y => S6856
    );
NAND_4028: ENTITY WORK.NAND
    PORT MAP (
        A => S6853,
        B => S6855,
        Y => S6857
    );
NOR_2431: ENTITY WORK.NOR
    PORT MAP (
        A => S6723,
        B => S6729,
        Y => S6858
    );
NAND_4029: ENTITY WORK.NAND
    PORT MAP (
        A => S6724,
        B => S6730,
        Y => S6859
    );
NOR_2432: ENTITY WORK.NOR
    PORT MAP (
        A => S910,
        B => S2107,
        Y => S6860
    );
NAND_4030: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_6,
        B => S2106,
        Y => S6861
    );
NOR_2433: ENTITY WORK.NOR
    PORT MAP (
        A => S805,
        B => S1953,
        Y => S6862
    );
NAND_4031: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_8,
        B => S1952,
        Y => S6863
    );
NOR_2434: ENTITY WORK.NOR
    PORT MAP (
        A => S6691,
        B => S6862,
        Y => S6864
    );
NAND_4032: ENTITY WORK.NAND
    PORT MAP (
        A => S6692,
        B => S6863,
        Y => S6865
    );
NOR_2435: ENTITY WORK.NOR
    PORT MAP (
        A => S805,
        B => S1598,
        Y => S6866
    );
NAND_4033: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_8,
        B => S1597,
        Y => S6867
    );
NOR_2436: ENTITY WORK.NOR
    PORT MAP (
        A => S6692,
        B => S6863,
        Y => S6868
    );
NAND_4034: ENTITY WORK.NAND
    PORT MAP (
        A => S6691,
        B => S6862,
        Y => S6869
    );
NOR_2437: ENTITY WORK.NOR
    PORT MAP (
        A => S6864,
        B => S6868,
        Y => S6870
    );
NAND_4035: ENTITY WORK.NAND
    PORT MAP (
        A => S6865,
        B => S6869,
        Y => S6871
    );
NOR_2438: ENTITY WORK.NOR
    PORT MAP (
        A => S6861,
        B => S6871,
        Y => S6872
    );
NAND_4036: ENTITY WORK.NAND
    PORT MAP (
        A => S6860,
        B => S6870,
        Y => S6873
    );
NOR_2439: ENTITY WORK.NOR
    PORT MAP (
        A => S6860,
        B => S6870,
        Y => S6874
    );
NAND_4037: ENTITY WORK.NAND
    PORT MAP (
        A => S6861,
        B => S6871,
        Y => S6875
    );
NOR_2440: ENTITY WORK.NOR
    PORT MAP (
        A => S6872,
        B => S6874,
        Y => S6876
    );
NAND_4038: ENTITY WORK.NAND
    PORT MAP (
        A => S6873,
        B => S6875,
        Y => S6877
    );
NOR_2441: ENTITY WORK.NOR
    PORT MAP (
        A => S6713,
        B => S6717,
        Y => S6878
    );
NAND_4039: ENTITY WORK.NAND
    PORT MAP (
        A => S6714,
        B => S6718,
        Y => S6879
    );
NOR_2442: ENTITY WORK.NOR
    PORT MAP (
        A => S754,
        B => S1849,
        Y => S6880
    );
NAND_4040: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_9,
        B => S1848,
        Y => S6881
    );
NOR_2443: ENTITY WORK.NOR
    PORT MAP (
        A => S651,
        B => S1516,
        Y => S6882
    );
NAND_4041: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_11,
        B => S1515,
        Y => S6883
    );
NOR_2444: ENTITY WORK.NOR
    PORT MAP (
        A => S6711,
        B => S6882,
        Y => S6884
    );
NAND_4042: ENTITY WORK.NAND
    PORT MAP (
        A => S6712,
        B => S6883,
        Y => S6885
    );
NOR_2445: ENTITY WORK.NOR
    PORT MAP (
        A => S651,
        B => S1746,
        Y => S6886
    );
NAND_4043: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_11,
        B => S1745,
        Y => S6887
    );
NOR_2446: ENTITY WORK.NOR
    PORT MAP (
        A => S6712,
        B => S6883,
        Y => S6888
    );
NAND_4044: ENTITY WORK.NAND
    PORT MAP (
        A => S6711,
        B => S6882,
        Y => S6889
    );
NOR_2447: ENTITY WORK.NOR
    PORT MAP (
        A => S6884,
        B => S6888,
        Y => S6890
    );
NAND_4045: ENTITY WORK.NAND
    PORT MAP (
        A => S6885,
        B => S6889,
        Y => S6891
    );
NOR_2448: ENTITY WORK.NOR
    PORT MAP (
        A => S6881,
        B => S6891,
        Y => S6892
    );
NAND_4046: ENTITY WORK.NAND
    PORT MAP (
        A => S6880,
        B => S6890,
        Y => S6893
    );
NOR_2449: ENTITY WORK.NOR
    PORT MAP (
        A => S6880,
        B => S6890,
        Y => S6894
    );
NAND_4047: ENTITY WORK.NAND
    PORT MAP (
        A => S6881,
        B => S6891,
        Y => S6895
    );
NOR_2450: ENTITY WORK.NOR
    PORT MAP (
        A => S6892,
        B => S6894,
        Y => S6896
    );
NAND_4048: ENTITY WORK.NAND
    PORT MAP (
        A => S6893,
        B => S6895,
        Y => S6897
    );
NOR_2451: ENTITY WORK.NOR
    PORT MAP (
        A => S6878,
        B => S6897,
        Y => S6898
    );
NAND_4049: ENTITY WORK.NAND
    PORT MAP (
        A => S6879,
        B => S6896,
        Y => S6899
    );
NOR_2452: ENTITY WORK.NOR
    PORT MAP (
        A => S6879,
        B => S6896,
        Y => S6900
    );
NAND_4050: ENTITY WORK.NAND
    PORT MAP (
        A => S6878,
        B => S6897,
        Y => S6901
    );
NOR_2453: ENTITY WORK.NOR
    PORT MAP (
        A => S6898,
        B => S6900,
        Y => S6902
    );
NAND_4051: ENTITY WORK.NAND
    PORT MAP (
        A => S6899,
        B => S6901,
        Y => S6903
    );
NOR_2454: ENTITY WORK.NOR
    PORT MAP (
        A => S6877,
        B => S6903,
        Y => S6904
    );
NAND_4052: ENTITY WORK.NAND
    PORT MAP (
        A => S6876,
        B => S6902,
        Y => S6905
    );
NOR_2455: ENTITY WORK.NOR
    PORT MAP (
        A => S6876,
        B => S6902,
        Y => S6906
    );
NAND_4053: ENTITY WORK.NAND
    PORT MAP (
        A => S6877,
        B => S6903,
        Y => S6907
    );
NOR_2456: ENTITY WORK.NOR
    PORT MAP (
        A => S6904,
        B => S6906,
        Y => S6908
    );
NAND_4054: ENTITY WORK.NAND
    PORT MAP (
        A => S6905,
        B => S6907,
        Y => S6909
    );
NOR_2457: ENTITY WORK.NOR
    PORT MAP (
        A => S6858,
        B => S6909,
        Y => S6910
    );
NAND_4055: ENTITY WORK.NAND
    PORT MAP (
        A => S6859,
        B => S6908,
        Y => S6911
    );
NOR_2458: ENTITY WORK.NOR
    PORT MAP (
        A => S6859,
        B => S6908,
        Y => S6912
    );
NAND_4056: ENTITY WORK.NAND
    PORT MAP (
        A => S6858,
        B => S6909,
        Y => S6913
    );
NOR_2459: ENTITY WORK.NOR
    PORT MAP (
        A => S6910,
        B => S6912,
        Y => S6914
    );
NAND_4057: ENTITY WORK.NAND
    PORT MAP (
        A => S6911,
        B => S6913,
        Y => S6915
    );
NOR_2460: ENTITY WORK.NOR
    PORT MAP (
        A => S6857,
        B => S6915,
        Y => S6916
    );
NAND_4058: ENTITY WORK.NAND
    PORT MAP (
        A => S6856,
        B => S6914,
        Y => S6917
    );
NOR_2461: ENTITY WORK.NOR
    PORT MAP (
        A => S6856,
        B => S6914,
        Y => S6918
    );
NAND_4059: ENTITY WORK.NAND
    PORT MAP (
        A => S6857,
        B => S6915,
        Y => S6919
    );
NOR_2462: ENTITY WORK.NOR
    PORT MAP (
        A => S6916,
        B => S6918,
        Y => S6920
    );
NAND_4060: ENTITY WORK.NAND
    PORT MAP (
        A => S6917,
        B => S6919,
        Y => S6921
    );
NOR_2463: ENTITY WORK.NOR
    PORT MAP (
        A => S6822,
        B => S6921,
        Y => S6922
    );
NAND_4061: ENTITY WORK.NAND
    PORT MAP (
        A => S6823,
        B => S6920,
        Y => S6923
    );
NOR_2464: ENTITY WORK.NOR
    PORT MAP (
        A => S6823,
        B => S6920,
        Y => S6924
    );
NAND_4062: ENTITY WORK.NAND
    PORT MAP (
        A => S6822,
        B => S6921,
        Y => S6925
    );
NOR_2465: ENTITY WORK.NOR
    PORT MAP (
        A => S6922,
        B => S6924,
        Y => S6926
    );
NAND_4063: ENTITY WORK.NAND
    PORT MAP (
        A => S6923,
        B => S6925,
        Y => S6927
    );
NOR_2466: ENTITY WORK.NOR
    PORT MAP (
        A => S6821,
        B => S6927,
        Y => S6928
    );
NAND_4064: ENTITY WORK.NAND
    PORT MAP (
        A => S6820,
        B => S6926,
        Y => S6929
    );
NOR_2467: ENTITY WORK.NOR
    PORT MAP (
        A => S6820,
        B => S6926,
        Y => S6930
    );
NAND_4065: ENTITY WORK.NAND
    PORT MAP (
        A => S6821,
        B => S6927,
        Y => S6931
    );
NOR_2468: ENTITY WORK.NOR
    PORT MAP (
        A => S6928,
        B => S6930,
        Y => S6932
    );
NAND_4066: ENTITY WORK.NAND
    PORT MAP (
        A => S6929,
        B => S6931,
        Y => S6933
    );
NOR_2469: ENTITY WORK.NOR
    PORT MAP (
        A => S6788,
        B => S6933,
        Y => S6934
    );
NAND_4067: ENTITY WORK.NAND
    PORT MAP (
        A => S6789,
        B => S6932,
        Y => S6935
    );
NOR_2470: ENTITY WORK.NOR
    PORT MAP (
        A => S6789,
        B => S6932,
        Y => S6936
    );
NAND_4068: ENTITY WORK.NAND
    PORT MAP (
        A => S6788,
        B => S6933,
        Y => S6937
    );
NOR_2471: ENTITY WORK.NOR
    PORT MAP (
        A => S6934,
        B => S6936,
        Y => S6938
    );
NAND_4069: ENTITY WORK.NAND
    PORT MAP (
        A => S6935,
        B => S6937,
        Y => S6939
    );
NOR_2472: ENTITY WORK.NOR
    PORT MAP (
        A => S6644,
        B => S6939,
        Y => S6940
    );
NAND_4070: ENTITY WORK.NAND
    PORT MAP (
        A => S6643,
        B => S6938,
        Y => S6941
    );
NOR_2473: ENTITY WORK.NOR
    PORT MAP (
        A => S6643,
        B => S6938,
        Y => S6942
    );
NAND_4071: ENTITY WORK.NAND
    PORT MAP (
        A => S6644,
        B => S6939,
        Y => S6943
    );
NOR_2474: ENTITY WORK.NOR
    PORT MAP (
        A => S6940,
        B => S6942,
        Y => S6944
    );
NAND_4072: ENTITY WORK.NAND
    PORT MAP (
        A => S6941,
        B => S6943,
        Y => S6945
    );
NAND_4073: ENTITY WORK.NAND
    PORT MAP (
        A => S6786,
        B => S6945,
        Y => S6946
    );
NAND_4074: ENTITY WORK.NAND
    PORT MAP (
        A => S6787,
        B => S6944,
        Y => S6947
    );
NAND_4075: ENTITY WORK.NAND
    PORT MAP (
        A => S6946,
        B => S6947,
        Y => S6948
    );
NOR_2475: ENTITY WORK.NOR
    PORT MAP (
        A => S6768,
        B => S6948,
        Y => S6949
    );
NOT_519: ENTITY WORK.NOT
    PORT MAP (
        A => S6949,
        Y => S6950
    );
NAND_4076: ENTITY WORK.NAND
    PORT MAP (
        A => S6768,
        B => S6948,
        Y => S6951
    );
NAND_4077: ENTITY WORK.NAND
    PORT MAP (
        A => S6950,
        B => S6951,
        Y => S6952
    );
NOR_2476: ENTITY WORK.NOR
    PORT MAP (
        A => S6785,
        B => S6952,
        Y => S6953
    );
NAND_4078: ENTITY WORK.NAND
    PORT MAP (
        A => S6785,
        B => S6952,
        Y => S6954
    );
NAND_4079: ENTITY WORK.NAND
    PORT MAP (
        A => S5948,
        B => S6954,
        Y => S6955
    );
NOR_2477: ENTITY WORK.NOR
    PORT MAP (
        A => S6953,
        B => S6955,
        Y => S6956
    );
NOR_2478: ENTITY WORK.NOR
    PORT MAP (
        A => S6783,
        B => S6956,
        Y => S6957
    );
NAND_4080: ENTITY WORK.NAND
    PORT MAP (
        A => S6784,
        B => S6957,
        Y => S293
    );
NOR_2479: ENTITY WORK.NOR
    PORT MAP (
        A => S3899,
        B => S4035,
        Y => S6958
    );
NAND_4081: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu1_12,
        B => S5950,
        Y => S6959
    );
NOR_2480: ENTITY WORK.NOR
    PORT MAP (
        A => S6949,
        B => S6953,
        Y => S6960
    );
NOR_2481: ENTITY WORK.NOR
    PORT MAP (
        A => S6934,
        B => S6940,
        Y => S6961
    );
NAND_4082: ENTITY WORK.NAND
    PORT MAP (
        A => S6935,
        B => S6941,
        Y => S6962
    );
NOR_2482: ENTITY WORK.NOR
    PORT MAP (
        A => S6922,
        B => S6928,
        Y => S6963
    );
NAND_4083: ENTITY WORK.NAND
    PORT MAP (
        A => S6923,
        B => S6929,
        Y => S6964
    );
NOR_2483: ENTITY WORK.NOR
    PORT MAP (
        A => S1220,
        B => S2817,
        Y => S6965
    );
NAND_4084: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_0,
        B => S2816,
        Y => S6966
    );
NOR_2484: ENTITY WORK.NOR
    PORT MAP (
        A => S6798,
        B => S6802,
        Y => S6967
    );
NAND_4085: ENTITY WORK.NAND
    PORT MAP (
        A => S6799,
        B => S6803,
        Y => S6968
    );
NOR_2485: ENTITY WORK.NOR
    PORT MAP (
        A => S1168,
        B => S2718,
        Y => S6969
    );
NAND_4086: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_1,
        B => S2717,
        Y => S6970
    );
NOR_2486: ENTITY WORK.NOR
    PORT MAP (
        A => S1065,
        B => S2518,
        Y => S6971
    );
NAND_4087: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_3,
        B => S2517,
        Y => S6972
    );
NOR_2487: ENTITY WORK.NOR
    PORT MAP (
        A => S6796,
        B => S6971,
        Y => S6973
    );
NAND_4088: ENTITY WORK.NAND
    PORT MAP (
        A => S6797,
        B => S6972,
        Y => S6974
    );
NOR_2488: ENTITY WORK.NOR
    PORT MAP (
        A => S1065,
        B => S2618,
        Y => S6975
    );
NAND_4089: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_3,
        B => S2617,
        Y => S6976
    );
NOR_2489: ENTITY WORK.NOR
    PORT MAP (
        A => S6797,
        B => S6972,
        Y => S6977
    );
NAND_4090: ENTITY WORK.NAND
    PORT MAP (
        A => S6796,
        B => S6971,
        Y => S6978
    );
NOR_2490: ENTITY WORK.NOR
    PORT MAP (
        A => S6973,
        B => S6977,
        Y => S6979
    );
NAND_4091: ENTITY WORK.NAND
    PORT MAP (
        A => S6974,
        B => S6978,
        Y => S6980
    );
NOR_2491: ENTITY WORK.NOR
    PORT MAP (
        A => S6970,
        B => S6980,
        Y => S6981
    );
NAND_4092: ENTITY WORK.NAND
    PORT MAP (
        A => S6969,
        B => S6979,
        Y => S6982
    );
NOR_2492: ENTITY WORK.NOR
    PORT MAP (
        A => S6969,
        B => S6979,
        Y => S6983
    );
NAND_4093: ENTITY WORK.NAND
    PORT MAP (
        A => S6970,
        B => S6980,
        Y => S6984
    );
NOR_2493: ENTITY WORK.NOR
    PORT MAP (
        A => S6981,
        B => S6983,
        Y => S6985
    );
NAND_4094: ENTITY WORK.NAND
    PORT MAP (
        A => S6982,
        B => S6984,
        Y => S6986
    );
NOR_2494: ENTITY WORK.NOR
    PORT MAP (
        A => S6967,
        B => S6986,
        Y => S6987
    );
NAND_4095: ENTITY WORK.NAND
    PORT MAP (
        A => S6968,
        B => S6985,
        Y => S6988
    );
NOR_2495: ENTITY WORK.NOR
    PORT MAP (
        A => S6968,
        B => S6985,
        Y => S6989
    );
NAND_4096: ENTITY WORK.NAND
    PORT MAP (
        A => S6967,
        B => S6986,
        Y => S6990
    );
NOR_2496: ENTITY WORK.NOR
    PORT MAP (
        A => S6987,
        B => S6989,
        Y => S6991
    );
NAND_4097: ENTITY WORK.NAND
    PORT MAP (
        A => S6988,
        B => S6990,
        Y => S6992
    );
NOR_2497: ENTITY WORK.NOR
    PORT MAP (
        A => S6966,
        B => S6992,
        Y => S6993
    );
NAND_4098: ENTITY WORK.NAND
    PORT MAP (
        A => S6965,
        B => S6991,
        Y => S6994
    );
NOR_2498: ENTITY WORK.NOR
    PORT MAP (
        A => S6965,
        B => S6991,
        Y => S6995
    );
NAND_4099: ENTITY WORK.NAND
    PORT MAP (
        A => S6966,
        B => S6992,
        Y => S6996
    );
NOR_2499: ENTITY WORK.NOR
    PORT MAP (
        A => S6993,
        B => S6995,
        Y => S6997
    );
NAND_4100: ENTITY WORK.NAND
    PORT MAP (
        A => S6994,
        B => S6996,
        Y => S6998
    );
NOR_2500: ENTITY WORK.NOR
    PORT MAP (
        A => S6846,
        B => S6854,
        Y => S6999
    );
NAND_4101: ENTITY WORK.NAND
    PORT MAP (
        A => S6847,
        B => S6855,
        Y => S7000
    );
NOR_2501: ENTITY WORK.NOR
    PORT MAP (
        A => S6998,
        B => S6999,
        Y => S7001
    );
NAND_4102: ENTITY WORK.NAND
    PORT MAP (
        A => S6997,
        B => S7000,
        Y => S7002
    );
NOR_2502: ENTITY WORK.NOR
    PORT MAP (
        A => S6997,
        B => S7000,
        Y => S7003
    );
NAND_4103: ENTITY WORK.NAND
    PORT MAP (
        A => S6998,
        B => S6999,
        Y => S7004
    );
NOR_2503: ENTITY WORK.NOR
    PORT MAP (
        A => S7001,
        B => S7003,
        Y => S7005
    );
NAND_4104: ENTITY WORK.NAND
    PORT MAP (
        A => S7002,
        B => S7004,
        Y => S7006
    );
NOR_2504: ENTITY WORK.NOR
    PORT MAP (
        A => S6809,
        B => S7006,
        Y => S7007
    );
NAND_4105: ENTITY WORK.NAND
    PORT MAP (
        A => S6808,
        B => S7005,
        Y => S7008
    );
NOR_2505: ENTITY WORK.NOR
    PORT MAP (
        A => S6808,
        B => S7005,
        Y => S7009
    );
NAND_4106: ENTITY WORK.NAND
    PORT MAP (
        A => S6809,
        B => S7006,
        Y => S7010
    );
NOR_2506: ENTITY WORK.NOR
    PORT MAP (
        A => S7007,
        B => S7009,
        Y => S7011
    );
NAND_4107: ENTITY WORK.NAND
    PORT MAP (
        A => S7008,
        B => S7010,
        Y => S7012
    );
NOR_2507: ENTITY WORK.NOR
    PORT MAP (
        A => S6910,
        B => S6916,
        Y => S7013
    );
NAND_4108: ENTITY WORK.NAND
    PORT MAP (
        A => S6911,
        B => S6917,
        Y => S7014
    );
NOR_2508: ENTITY WORK.NOR
    PORT MAP (
        A => S6834,
        B => S6838,
        Y => S7015
    );
NAND_4109: ENTITY WORK.NAND
    PORT MAP (
        A => S6835,
        B => S6839,
        Y => S7016
    );
NOR_2509: ENTITY WORK.NOR
    PORT MAP (
        A => S1013,
        B => S2418,
        Y => S7017
    );
NAND_4110: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_4,
        B => S2417,
        Y => S7018
    );
NOR_2510: ENTITY WORK.NOR
    PORT MAP (
        A => S910,
        B => S2206,
        Y => S7019
    );
NAND_4111: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_6,
        B => S2205,
        Y => S7020
    );
NOR_2511: ENTITY WORK.NOR
    PORT MAP (
        A => S6832,
        B => S7019,
        Y => S7021
    );
NAND_4112: ENTITY WORK.NAND
    PORT MAP (
        A => S6833,
        B => S7020,
        Y => S7022
    );
NOR_2512: ENTITY WORK.NOR
    PORT MAP (
        A => S910,
        B => S2312,
        Y => S7023
    );
NAND_4113: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_6,
        B => S2311,
        Y => S7024
    );
NOR_2513: ENTITY WORK.NOR
    PORT MAP (
        A => S6833,
        B => S7020,
        Y => S7025
    );
NAND_4114: ENTITY WORK.NAND
    PORT MAP (
        A => S6832,
        B => S7019,
        Y => S7026
    );
NOR_2514: ENTITY WORK.NOR
    PORT MAP (
        A => S7021,
        B => S7025,
        Y => S7027
    );
NAND_4115: ENTITY WORK.NAND
    PORT MAP (
        A => S7022,
        B => S7026,
        Y => S7028
    );
NOR_2515: ENTITY WORK.NOR
    PORT MAP (
        A => S7018,
        B => S7028,
        Y => S7029
    );
NAND_4116: ENTITY WORK.NAND
    PORT MAP (
        A => S7017,
        B => S7027,
        Y => S7030
    );
NOR_2516: ENTITY WORK.NOR
    PORT MAP (
        A => S7017,
        B => S7027,
        Y => S7031
    );
NAND_4117: ENTITY WORK.NAND
    PORT MAP (
        A => S7018,
        B => S7028,
        Y => S7032
    );
NOR_2517: ENTITY WORK.NOR
    PORT MAP (
        A => S7029,
        B => S7031,
        Y => S7033
    );
NAND_4118: ENTITY WORK.NAND
    PORT MAP (
        A => S7030,
        B => S7032,
        Y => S7034
    );
NOR_2518: ENTITY WORK.NOR
    PORT MAP (
        A => S6868,
        B => S6872,
        Y => S7035
    );
NAND_4119: ENTITY WORK.NAND
    PORT MAP (
        A => S6869,
        B => S6873,
        Y => S7036
    );
NOR_2519: ENTITY WORK.NOR
    PORT MAP (
        A => S7034,
        B => S7035,
        Y => S7037
    );
NAND_4120: ENTITY WORK.NAND
    PORT MAP (
        A => S7033,
        B => S7036,
        Y => S7038
    );
NOR_2520: ENTITY WORK.NOR
    PORT MAP (
        A => S7033,
        B => S7036,
        Y => S7039
    );
NAND_4121: ENTITY WORK.NAND
    PORT MAP (
        A => S7034,
        B => S7035,
        Y => S7040
    );
NOR_2521: ENTITY WORK.NOR
    PORT MAP (
        A => S7037,
        B => S7039,
        Y => S7041
    );
NAND_4122: ENTITY WORK.NAND
    PORT MAP (
        A => S7038,
        B => S7040,
        Y => S7042
    );
NOR_2522: ENTITY WORK.NOR
    PORT MAP (
        A => S7016,
        B => S7041,
        Y => S7043
    );
NAND_4123: ENTITY WORK.NAND
    PORT MAP (
        A => S7015,
        B => S7042,
        Y => S7044
    );
NOR_2523: ENTITY WORK.NOR
    PORT MAP (
        A => S7015,
        B => S7042,
        Y => S7045
    );
NAND_4124: ENTITY WORK.NAND
    PORT MAP (
        A => S7016,
        B => S7041,
        Y => S7046
    );
NOR_2524: ENTITY WORK.NOR
    PORT MAP (
        A => S7043,
        B => S7045,
        Y => S7047
    );
NAND_4125: ENTITY WORK.NAND
    PORT MAP (
        A => S7044,
        B => S7046,
        Y => S7048
    );
NOR_2525: ENTITY WORK.NOR
    PORT MAP (
        A => S6898,
        B => S6904,
        Y => S7049
    );
NAND_4126: ENTITY WORK.NAND
    PORT MAP (
        A => S6899,
        B => S6905,
        Y => S7050
    );
NOR_2526: ENTITY WORK.NOR
    PORT MAP (
        A => S858,
        B => S2107,
        Y => S7051
    );
NAND_4127: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_7,
        B => S2106,
        Y => S7052
    );
NOR_2527: ENTITY WORK.NOR
    PORT MAP (
        A => S754,
        B => S1953,
        Y => S7053
    );
NAND_4128: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_9,
        B => S1952,
        Y => S7054
    );
NOR_2528: ENTITY WORK.NOR
    PORT MAP (
        A => S6866,
        B => S7053,
        Y => S7055
    );
NAND_4129: ENTITY WORK.NAND
    PORT MAP (
        A => S6867,
        B => S7054,
        Y => S7056
    );
NOR_2529: ENTITY WORK.NOR
    PORT MAP (
        A => S754,
        B => S1598,
        Y => S7057
    );
NAND_4130: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_9,
        B => S1597,
        Y => S7058
    );
NOR_2530: ENTITY WORK.NOR
    PORT MAP (
        A => S6867,
        B => S7054,
        Y => S7059
    );
NAND_4131: ENTITY WORK.NAND
    PORT MAP (
        A => S6866,
        B => S7053,
        Y => S7060
    );
NOR_2531: ENTITY WORK.NOR
    PORT MAP (
        A => S7055,
        B => S7059,
        Y => S7061
    );
NAND_4132: ENTITY WORK.NAND
    PORT MAP (
        A => S7056,
        B => S7060,
        Y => S7062
    );
NOR_2532: ENTITY WORK.NOR
    PORT MAP (
        A => S7052,
        B => S7062,
        Y => S7063
    );
NAND_4133: ENTITY WORK.NAND
    PORT MAP (
        A => S7051,
        B => S7061,
        Y => S7064
    );
NOR_2533: ENTITY WORK.NOR
    PORT MAP (
        A => S7051,
        B => S7061,
        Y => S7065
    );
NAND_4134: ENTITY WORK.NAND
    PORT MAP (
        A => S7052,
        B => S7062,
        Y => S7066
    );
NOR_2534: ENTITY WORK.NOR
    PORT MAP (
        A => S7063,
        B => S7065,
        Y => S7067
    );
NAND_4135: ENTITY WORK.NAND
    PORT MAP (
        A => S7064,
        B => S7066,
        Y => S7068
    );
NOR_2535: ENTITY WORK.NOR
    PORT MAP (
        A => S6888,
        B => S6892,
        Y => S7069
    );
NAND_4136: ENTITY WORK.NAND
    PORT MAP (
        A => S6889,
        B => S6893,
        Y => S7070
    );
NOR_2536: ENTITY WORK.NOR
    PORT MAP (
        A => S702,
        B => S1849,
        Y => S7071
    );
NAND_4137: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_10,
        B => S1848,
        Y => S7072
    );
NOR_2537: ENTITY WORK.NOR
    PORT MAP (
        A => S599,
        B => S1516,
        Y => S7073
    );
NAND_4138: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_12,
        B => S1515,
        Y => S7074
    );
NOR_2538: ENTITY WORK.NOR
    PORT MAP (
        A => S6886,
        B => S7073,
        Y => S7075
    );
NAND_4139: ENTITY WORK.NAND
    PORT MAP (
        A => S6887,
        B => S7074,
        Y => S7076
    );
NOR_2539: ENTITY WORK.NOR
    PORT MAP (
        A => S599,
        B => S1746,
        Y => S7077
    );
NAND_4140: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_12,
        B => S1745,
        Y => S7078
    );
NOR_2540: ENTITY WORK.NOR
    PORT MAP (
        A => S6887,
        B => S7074,
        Y => S7079
    );
NAND_4141: ENTITY WORK.NAND
    PORT MAP (
        A => S6886,
        B => S7073,
        Y => S7080
    );
NOR_2541: ENTITY WORK.NOR
    PORT MAP (
        A => S7075,
        B => S7079,
        Y => S7081
    );
NAND_4142: ENTITY WORK.NAND
    PORT MAP (
        A => S7076,
        B => S7080,
        Y => S7082
    );
NOR_2542: ENTITY WORK.NOR
    PORT MAP (
        A => S7072,
        B => S7082,
        Y => S7083
    );
NAND_4143: ENTITY WORK.NAND
    PORT MAP (
        A => S7071,
        B => S7081,
        Y => S7084
    );
NOR_2543: ENTITY WORK.NOR
    PORT MAP (
        A => S7071,
        B => S7081,
        Y => S7085
    );
NAND_4144: ENTITY WORK.NAND
    PORT MAP (
        A => S7072,
        B => S7082,
        Y => S7086
    );
NOR_2544: ENTITY WORK.NOR
    PORT MAP (
        A => S7083,
        B => S7085,
        Y => S7087
    );
NAND_4145: ENTITY WORK.NAND
    PORT MAP (
        A => S7084,
        B => S7086,
        Y => S7088
    );
NOR_2545: ENTITY WORK.NOR
    PORT MAP (
        A => S7069,
        B => S7088,
        Y => S7089
    );
NAND_4146: ENTITY WORK.NAND
    PORT MAP (
        A => S7070,
        B => S7087,
        Y => S7090
    );
NOR_2546: ENTITY WORK.NOR
    PORT MAP (
        A => S7070,
        B => S7087,
        Y => S7091
    );
NAND_4147: ENTITY WORK.NAND
    PORT MAP (
        A => S7069,
        B => S7088,
        Y => S7092
    );
NOR_2547: ENTITY WORK.NOR
    PORT MAP (
        A => S7089,
        B => S7091,
        Y => S7093
    );
NAND_4148: ENTITY WORK.NAND
    PORT MAP (
        A => S7090,
        B => S7092,
        Y => S7094
    );
NOR_2548: ENTITY WORK.NOR
    PORT MAP (
        A => S7068,
        B => S7094,
        Y => S7095
    );
NAND_4149: ENTITY WORK.NAND
    PORT MAP (
        A => S7067,
        B => S7093,
        Y => S7096
    );
NOR_2549: ENTITY WORK.NOR
    PORT MAP (
        A => S7067,
        B => S7093,
        Y => S7097
    );
NAND_4150: ENTITY WORK.NAND
    PORT MAP (
        A => S7068,
        B => S7094,
        Y => S7098
    );
NOR_2550: ENTITY WORK.NOR
    PORT MAP (
        A => S7095,
        B => S7097,
        Y => S7099
    );
NAND_4151: ENTITY WORK.NAND
    PORT MAP (
        A => S7096,
        B => S7098,
        Y => S7100
    );
NOR_2551: ENTITY WORK.NOR
    PORT MAP (
        A => S7049,
        B => S7100,
        Y => S7101
    );
NAND_4152: ENTITY WORK.NAND
    PORT MAP (
        A => S7050,
        B => S7099,
        Y => S7102
    );
NOR_2552: ENTITY WORK.NOR
    PORT MAP (
        A => S7050,
        B => S7099,
        Y => S7103
    );
NAND_4153: ENTITY WORK.NAND
    PORT MAP (
        A => S7049,
        B => S7100,
        Y => S7104
    );
NOR_2553: ENTITY WORK.NOR
    PORT MAP (
        A => S7101,
        B => S7103,
        Y => S7105
    );
NAND_4154: ENTITY WORK.NAND
    PORT MAP (
        A => S7102,
        B => S7104,
        Y => S7106
    );
NOR_2554: ENTITY WORK.NOR
    PORT MAP (
        A => S7048,
        B => S7106,
        Y => S7107
    );
NAND_4155: ENTITY WORK.NAND
    PORT MAP (
        A => S7047,
        B => S7105,
        Y => S7108
    );
NOR_2555: ENTITY WORK.NOR
    PORT MAP (
        A => S7047,
        B => S7105,
        Y => S7109
    );
NAND_4156: ENTITY WORK.NAND
    PORT MAP (
        A => S7048,
        B => S7106,
        Y => S7110
    );
NOR_2556: ENTITY WORK.NOR
    PORT MAP (
        A => S7107,
        B => S7109,
        Y => S7111
    );
NAND_4157: ENTITY WORK.NAND
    PORT MAP (
        A => S7108,
        B => S7110,
        Y => S7112
    );
NOR_2557: ENTITY WORK.NOR
    PORT MAP (
        A => S7013,
        B => S7112,
        Y => S7113
    );
NAND_4158: ENTITY WORK.NAND
    PORT MAP (
        A => S7014,
        B => S7111,
        Y => S7114
    );
NOR_2558: ENTITY WORK.NOR
    PORT MAP (
        A => S7014,
        B => S7111,
        Y => S7115
    );
NAND_4159: ENTITY WORK.NAND
    PORT MAP (
        A => S7013,
        B => S7112,
        Y => S7116
    );
NOR_2559: ENTITY WORK.NOR
    PORT MAP (
        A => S7113,
        B => S7115,
        Y => S7117
    );
NAND_4160: ENTITY WORK.NAND
    PORT MAP (
        A => S7114,
        B => S7116,
        Y => S7118
    );
NOR_2560: ENTITY WORK.NOR
    PORT MAP (
        A => S7012,
        B => S7118,
        Y => S7119
    );
NAND_4161: ENTITY WORK.NAND
    PORT MAP (
        A => S7011,
        B => S7117,
        Y => S7120
    );
NOR_2561: ENTITY WORK.NOR
    PORT MAP (
        A => S7011,
        B => S7117,
        Y => S7121
    );
NAND_4162: ENTITY WORK.NAND
    PORT MAP (
        A => S7012,
        B => S7118,
        Y => S7122
    );
NOR_2562: ENTITY WORK.NOR
    PORT MAP (
        A => S7119,
        B => S7121,
        Y => S7123
    );
NAND_4163: ENTITY WORK.NAND
    PORT MAP (
        A => S7120,
        B => S7122,
        Y => S7124
    );
NOR_2563: ENTITY WORK.NOR
    PORT MAP (
        A => S6963,
        B => S7124,
        Y => S7125
    );
NAND_4164: ENTITY WORK.NAND
    PORT MAP (
        A => S6964,
        B => S7123,
        Y => S7126
    );
NOR_2564: ENTITY WORK.NOR
    PORT MAP (
        A => S6964,
        B => S7123,
        Y => S7127
    );
NAND_4165: ENTITY WORK.NAND
    PORT MAP (
        A => S6963,
        B => S7124,
        Y => S7128
    );
NOR_2565: ENTITY WORK.NOR
    PORT MAP (
        A => S7125,
        B => S7127,
        Y => S7129
    );
NAND_4166: ENTITY WORK.NAND
    PORT MAP (
        A => S7126,
        B => S7128,
        Y => S7130
    );
NOR_2566: ENTITY WORK.NOR
    PORT MAP (
        A => S6819,
        B => S7130,
        Y => S7131
    );
NAND_4167: ENTITY WORK.NAND
    PORT MAP (
        A => S6818,
        B => S7129,
        Y => S7132
    );
NOR_2567: ENTITY WORK.NOR
    PORT MAP (
        A => S6818,
        B => S7129,
        Y => S7133
    );
NAND_4168: ENTITY WORK.NAND
    PORT MAP (
        A => S6819,
        B => S7130,
        Y => S7134
    );
NOR_2568: ENTITY WORK.NOR
    PORT MAP (
        A => S7131,
        B => S7133,
        Y => S7135
    );
NAND_4169: ENTITY WORK.NAND
    PORT MAP (
        A => S7132,
        B => S7134,
        Y => S7136
    );
NAND_4170: ENTITY WORK.NAND
    PORT MAP (
        A => S6961,
        B => S7136,
        Y => S7137
    );
NAND_4171: ENTITY WORK.NAND
    PORT MAP (
        A => S6962,
        B => S7135,
        Y => S7138
    );
NAND_4172: ENTITY WORK.NAND
    PORT MAP (
        A => S7137,
        B => S7138,
        Y => S7139
    );
NOR_2569: ENTITY WORK.NOR
    PORT MAP (
        A => S6947,
        B => S7139,
        Y => S7140
    );
NOT_520: ENTITY WORK.NOT
    PORT MAP (
        A => S7140,
        Y => S7141
    );
NAND_4173: ENTITY WORK.NAND
    PORT MAP (
        A => S6947,
        B => S7139,
        Y => S7142
    );
NAND_4174: ENTITY WORK.NAND
    PORT MAP (
        A => S7141,
        B => S7142,
        Y => S7143
    );
NOR_2570: ENTITY WORK.NOR
    PORT MAP (
        A => S6960,
        B => S7143,
        Y => S7144
    );
NAND_4175: ENTITY WORK.NAND
    PORT MAP (
        A => S6960,
        B => S7143,
        Y => S7145
    );
NAND_4176: ENTITY WORK.NAND
    PORT MAP (
        A => S5948,
        B => S7145,
        Y => S7146
    );
NOR_2571: ENTITY WORK.NOR
    PORT MAP (
        A => S7144,
        B => S7146,
        Y => S7147
    );
NOR_2572: ENTITY WORK.NOR
    PORT MAP (
        A => S6958,
        B => S7147,
        Y => S7148
    );
NAND_4177: ENTITY WORK.NAND
    PORT MAP (
        A => S6959,
        B => S7148,
        Y => S294
    );
NOR_2573: ENTITY WORK.NOR
    PORT MAP (
        A => S7140,
        B => S7144,
        Y => S7149
    );
NOR_2574: ENTITY WORK.NOR
    PORT MAP (
        A => S7125,
        B => S7131,
        Y => S7150
    );
NAND_4178: ENTITY WORK.NAND
    PORT MAP (
        A => S7126,
        B => S7132,
        Y => S7151
    );
NOR_2575: ENTITY WORK.NOR
    PORT MAP (
        A => S7001,
        B => S7007,
        Y => S7152
    );
NAND_4179: ENTITY WORK.NAND
    PORT MAP (
        A => S7002,
        B => S7008,
        Y => S7153
    );
NOR_2576: ENTITY WORK.NOR
    PORT MAP (
        A => S7113,
        B => S7119,
        Y => S7154
    );
NAND_4180: ENTITY WORK.NAND
    PORT MAP (
        A => S7114,
        B => S7120,
        Y => S7155
    );
NOR_2577: ENTITY WORK.NOR
    PORT MAP (
        A => S6987,
        B => S6993,
        Y => S7156
    );
NAND_4181: ENTITY WORK.NAND
    PORT MAP (
        A => S6988,
        B => S6994,
        Y => S7157
    );
NOR_2578: ENTITY WORK.NOR
    PORT MAP (
        A => S1220,
        B => S2920,
        Y => S7158
    );
NOR_2579: ENTITY WORK.NOR
    PORT MAP (
        A => S1168,
        B => S2817,
        Y => S7159
    );
NAND_4182: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_1,
        B => S2816,
        Y => S7160
    );
NOR_2580: ENTITY WORK.NOR
    PORT MAP (
        A => S7158,
        B => S7159,
        Y => S7161
    );
NOT_521: ENTITY WORK.NOT
    PORT MAP (
        A => S7161,
        Y => S7162
    );
NOR_2581: ENTITY WORK.NOR
    PORT MAP (
        A => S1168,
        B => S2920,
        Y => S7163
    );
NAND_4183: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_1,
        B => S2919,
        Y => S7164
    );
NOR_2582: ENTITY WORK.NOR
    PORT MAP (
        A => S6966,
        B => S7164,
        Y => S7165
    );
NAND_4184: ENTITY WORK.NAND
    PORT MAP (
        A => S6965,
        B => S7163,
        Y => S7166
    );
NOR_2583: ENTITY WORK.NOR
    PORT MAP (
        A => S7161,
        B => S7165,
        Y => S7167
    );
NAND_4185: ENTITY WORK.NAND
    PORT MAP (
        A => S7162,
        B => S7166,
        Y => S7168
    );
NOR_2584: ENTITY WORK.NOR
    PORT MAP (
        A => S6977,
        B => S6981,
        Y => S7169
    );
NAND_4186: ENTITY WORK.NAND
    PORT MAP (
        A => S6978,
        B => S6982,
        Y => S7170
    );
NOR_2585: ENTITY WORK.NOR
    PORT MAP (
        A => S1116,
        B => S2718,
        Y => S7171
    );
NAND_4187: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_2,
        B => S2717,
        Y => S7172
    );
NOR_2586: ENTITY WORK.NOR
    PORT MAP (
        A => S1013,
        B => S2518,
        Y => S7173
    );
NAND_4188: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_4,
        B => S2517,
        Y => S7174
    );
NOR_2587: ENTITY WORK.NOR
    PORT MAP (
        A => S6975,
        B => S7173,
        Y => S7175
    );
NAND_4189: ENTITY WORK.NAND
    PORT MAP (
        A => S6976,
        B => S7174,
        Y => S7176
    );
NOR_2588: ENTITY WORK.NOR
    PORT MAP (
        A => S1013,
        B => S2618,
        Y => S7177
    );
NAND_4190: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_4,
        B => S2617,
        Y => S7178
    );
NOR_2589: ENTITY WORK.NOR
    PORT MAP (
        A => S6976,
        B => S7174,
        Y => S7179
    );
NAND_4191: ENTITY WORK.NAND
    PORT MAP (
        A => S6975,
        B => S7173,
        Y => S7180
    );
NOR_2590: ENTITY WORK.NOR
    PORT MAP (
        A => S7175,
        B => S7179,
        Y => S7181
    );
NAND_4192: ENTITY WORK.NAND
    PORT MAP (
        A => S7176,
        B => S7180,
        Y => S7182
    );
NOR_2591: ENTITY WORK.NOR
    PORT MAP (
        A => S7172,
        B => S7182,
        Y => S7183
    );
NAND_4193: ENTITY WORK.NAND
    PORT MAP (
        A => S7171,
        B => S7181,
        Y => S7184
    );
NOR_2592: ENTITY WORK.NOR
    PORT MAP (
        A => S7171,
        B => S7181,
        Y => S7185
    );
NAND_4194: ENTITY WORK.NAND
    PORT MAP (
        A => S7172,
        B => S7182,
        Y => S7186
    );
NOR_2593: ENTITY WORK.NOR
    PORT MAP (
        A => S7183,
        B => S7185,
        Y => S7187
    );
NAND_4195: ENTITY WORK.NAND
    PORT MAP (
        A => S7184,
        B => S7186,
        Y => S7188
    );
NOR_2594: ENTITY WORK.NOR
    PORT MAP (
        A => S7169,
        B => S7188,
        Y => S7189
    );
NAND_4196: ENTITY WORK.NAND
    PORT MAP (
        A => S7170,
        B => S7187,
        Y => S7190
    );
NOR_2595: ENTITY WORK.NOR
    PORT MAP (
        A => S7170,
        B => S7187,
        Y => S7191
    );
NAND_4197: ENTITY WORK.NAND
    PORT MAP (
        A => S7169,
        B => S7188,
        Y => S7192
    );
NOR_2596: ENTITY WORK.NOR
    PORT MAP (
        A => S7189,
        B => S7191,
        Y => S7193
    );
NAND_4198: ENTITY WORK.NAND
    PORT MAP (
        A => S7190,
        B => S7192,
        Y => S7194
    );
NOR_2597: ENTITY WORK.NOR
    PORT MAP (
        A => S7167,
        B => S7193,
        Y => S7195
    );
NAND_4199: ENTITY WORK.NAND
    PORT MAP (
        A => S7168,
        B => S7194,
        Y => S7196
    );
NOR_2598: ENTITY WORK.NOR
    PORT MAP (
        A => S7168,
        B => S7194,
        Y => S7197
    );
NAND_4200: ENTITY WORK.NAND
    PORT MAP (
        A => S7167,
        B => S7193,
        Y => S7198
    );
NOR_2599: ENTITY WORK.NOR
    PORT MAP (
        A => S7195,
        B => S7197,
        Y => S7199
    );
NAND_4201: ENTITY WORK.NAND
    PORT MAP (
        A => S7196,
        B => S7198,
        Y => S7200
    );
NOR_2600: ENTITY WORK.NOR
    PORT MAP (
        A => S7037,
        B => S7045,
        Y => S7201
    );
NAND_4202: ENTITY WORK.NAND
    PORT MAP (
        A => S7038,
        B => S7046,
        Y => S7202
    );
NOR_2601: ENTITY WORK.NOR
    PORT MAP (
        A => S7200,
        B => S7201,
        Y => S7203
    );
NAND_4203: ENTITY WORK.NAND
    PORT MAP (
        A => S7199,
        B => S7202,
        Y => S7204
    );
NOR_2602: ENTITY WORK.NOR
    PORT MAP (
        A => S7199,
        B => S7202,
        Y => S7205
    );
NAND_4204: ENTITY WORK.NAND
    PORT MAP (
        A => S7200,
        B => S7201,
        Y => S7206
    );
NOR_2603: ENTITY WORK.NOR
    PORT MAP (
        A => S7203,
        B => S7205,
        Y => S7207
    );
NAND_4205: ENTITY WORK.NAND
    PORT MAP (
        A => S7204,
        B => S7206,
        Y => S7208
    );
NOR_2604: ENTITY WORK.NOR
    PORT MAP (
        A => S7157,
        B => S7207,
        Y => S7209
    );
NAND_4206: ENTITY WORK.NAND
    PORT MAP (
        A => S7156,
        B => S7208,
        Y => S7210
    );
NOR_2605: ENTITY WORK.NOR
    PORT MAP (
        A => S7156,
        B => S7208,
        Y => S7211
    );
NAND_4207: ENTITY WORK.NAND
    PORT MAP (
        A => S7157,
        B => S7207,
        Y => S7212
    );
NOR_2606: ENTITY WORK.NOR
    PORT MAP (
        A => S7209,
        B => S7211,
        Y => S7213
    );
NAND_4208: ENTITY WORK.NAND
    PORT MAP (
        A => S7210,
        B => S7212,
        Y => S7214
    );
NOR_2607: ENTITY WORK.NOR
    PORT MAP (
        A => S7101,
        B => S7107,
        Y => S7215
    );
NAND_4209: ENTITY WORK.NAND
    PORT MAP (
        A => S7102,
        B => S7108,
        Y => S7216
    );
NOR_2608: ENTITY WORK.NOR
    PORT MAP (
        A => S7025,
        B => S7029,
        Y => S7217
    );
NAND_4210: ENTITY WORK.NAND
    PORT MAP (
        A => S7026,
        B => S7030,
        Y => S7218
    );
NOR_2609: ENTITY WORK.NOR
    PORT MAP (
        A => S963,
        B => S2418,
        Y => S7219
    );
NAND_4211: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_5,
        B => S2417,
        Y => S7220
    );
NOR_2610: ENTITY WORK.NOR
    PORT MAP (
        A => S858,
        B => S2206,
        Y => S7221
    );
NAND_4212: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_7,
        B => S2205,
        Y => S7222
    );
NOR_2611: ENTITY WORK.NOR
    PORT MAP (
        A => S7023,
        B => S7221,
        Y => S7223
    );
NAND_4213: ENTITY WORK.NAND
    PORT MAP (
        A => S7024,
        B => S7222,
        Y => S7224
    );
NOR_2612: ENTITY WORK.NOR
    PORT MAP (
        A => S858,
        B => S2312,
        Y => S7225
    );
NAND_4214: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_7,
        B => S2311,
        Y => S7226
    );
NOR_2613: ENTITY WORK.NOR
    PORT MAP (
        A => S7024,
        B => S7222,
        Y => S7227
    );
NAND_4215: ENTITY WORK.NAND
    PORT MAP (
        A => S7023,
        B => S7221,
        Y => S7228
    );
NOR_2614: ENTITY WORK.NOR
    PORT MAP (
        A => S7223,
        B => S7227,
        Y => S7229
    );
NAND_4216: ENTITY WORK.NAND
    PORT MAP (
        A => S7224,
        B => S7228,
        Y => S7230
    );
NOR_2615: ENTITY WORK.NOR
    PORT MAP (
        A => S7220,
        B => S7230,
        Y => S7231
    );
NAND_4217: ENTITY WORK.NAND
    PORT MAP (
        A => S7219,
        B => S7229,
        Y => S7232
    );
NOR_2616: ENTITY WORK.NOR
    PORT MAP (
        A => S7219,
        B => S7229,
        Y => S7233
    );
NAND_4218: ENTITY WORK.NAND
    PORT MAP (
        A => S7220,
        B => S7230,
        Y => S7234
    );
NOR_2617: ENTITY WORK.NOR
    PORT MAP (
        A => S7231,
        B => S7233,
        Y => S7235
    );
NAND_4219: ENTITY WORK.NAND
    PORT MAP (
        A => S7232,
        B => S7234,
        Y => S7236
    );
NOR_2618: ENTITY WORK.NOR
    PORT MAP (
        A => S7059,
        B => S7063,
        Y => S7237
    );
NAND_4220: ENTITY WORK.NAND
    PORT MAP (
        A => S7060,
        B => S7064,
        Y => S7238
    );
NOR_2619: ENTITY WORK.NOR
    PORT MAP (
        A => S7236,
        B => S7237,
        Y => S7239
    );
NAND_4221: ENTITY WORK.NAND
    PORT MAP (
        A => S7235,
        B => S7238,
        Y => S7240
    );
NOR_2620: ENTITY WORK.NOR
    PORT MAP (
        A => S7235,
        B => S7238,
        Y => S7241
    );
NAND_4222: ENTITY WORK.NAND
    PORT MAP (
        A => S7236,
        B => S7237,
        Y => S7242
    );
NOR_2621: ENTITY WORK.NOR
    PORT MAP (
        A => S7239,
        B => S7241,
        Y => S7243
    );
NAND_4223: ENTITY WORK.NAND
    PORT MAP (
        A => S7240,
        B => S7242,
        Y => S7244
    );
NOR_2622: ENTITY WORK.NOR
    PORT MAP (
        A => S7218,
        B => S7243,
        Y => S7245
    );
NAND_4224: ENTITY WORK.NAND
    PORT MAP (
        A => S7217,
        B => S7244,
        Y => S7246
    );
NOR_2623: ENTITY WORK.NOR
    PORT MAP (
        A => S7217,
        B => S7244,
        Y => S7247
    );
NAND_4225: ENTITY WORK.NAND
    PORT MAP (
        A => S7218,
        B => S7243,
        Y => S7248
    );
NOR_2624: ENTITY WORK.NOR
    PORT MAP (
        A => S7245,
        B => S7247,
        Y => S7249
    );
NAND_4226: ENTITY WORK.NAND
    PORT MAP (
        A => S7246,
        B => S7248,
        Y => S7250
    );
NOR_2625: ENTITY WORK.NOR
    PORT MAP (
        A => S7089,
        B => S7095,
        Y => S7251
    );
NAND_4227: ENTITY WORK.NAND
    PORT MAP (
        A => S7090,
        B => S7096,
        Y => S7252
    );
NOR_2626: ENTITY WORK.NOR
    PORT MAP (
        A => S805,
        B => S2107,
        Y => S7253
    );
NAND_4228: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_8,
        B => S2106,
        Y => S7254
    );
NOR_2627: ENTITY WORK.NOR
    PORT MAP (
        A => S702,
        B => S1953,
        Y => S7255
    );
NAND_4229: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_10,
        B => S1952,
        Y => S7256
    );
NOR_2628: ENTITY WORK.NOR
    PORT MAP (
        A => S7057,
        B => S7255,
        Y => S7257
    );
NAND_4230: ENTITY WORK.NAND
    PORT MAP (
        A => S7058,
        B => S7256,
        Y => S7258
    );
NAND_4231: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_10,
        B => S1597,
        Y => S7259
    );
NOR_2629: ENTITY WORK.NOR
    PORT MAP (
        A => S7058,
        B => S7256,
        Y => S7260
    );
NAND_4232: ENTITY WORK.NAND
    PORT MAP (
        A => S7057,
        B => S7255,
        Y => S7261
    );
NOR_2630: ENTITY WORK.NOR
    PORT MAP (
        A => S7257,
        B => S7260,
        Y => S7262
    );
NAND_4233: ENTITY WORK.NAND
    PORT MAP (
        A => S7258,
        B => S7261,
        Y => S7263
    );
NOR_2631: ENTITY WORK.NOR
    PORT MAP (
        A => S7254,
        B => S7263,
        Y => S7264
    );
NAND_4234: ENTITY WORK.NAND
    PORT MAP (
        A => S7253,
        B => S7262,
        Y => S7265
    );
NOR_2632: ENTITY WORK.NOR
    PORT MAP (
        A => S7253,
        B => S7262,
        Y => S7266
    );
NAND_4235: ENTITY WORK.NAND
    PORT MAP (
        A => S7254,
        B => S7263,
        Y => S7267
    );
NOR_2633: ENTITY WORK.NOR
    PORT MAP (
        A => S7264,
        B => S7266,
        Y => S7268
    );
NAND_4236: ENTITY WORK.NAND
    PORT MAP (
        A => S7265,
        B => S7267,
        Y => S7269
    );
NOR_2634: ENTITY WORK.NOR
    PORT MAP (
        A => S7079,
        B => S7083,
        Y => S7270
    );
NAND_4237: ENTITY WORK.NAND
    PORT MAP (
        A => S7080,
        B => S7084,
        Y => S7271
    );
NOR_2635: ENTITY WORK.NOR
    PORT MAP (
        A => S651,
        B => S1849,
        Y => S7272
    );
NAND_4238: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_11,
        B => S1848,
        Y => S7273
    );
NOR_2636: ENTITY WORK.NOR
    PORT MAP (
        A => S548,
        B => S1516,
        Y => S7274
    );
NAND_4239: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_13,
        B => S1515,
        Y => S7275
    );
NOR_2637: ENTITY WORK.NOR
    PORT MAP (
        A => S7077,
        B => S7274,
        Y => S7276
    );
NAND_4240: ENTITY WORK.NAND
    PORT MAP (
        A => S7078,
        B => S7275,
        Y => S7277
    );
NAND_4241: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_13,
        B => S1745,
        Y => S7278
    );
NOR_2638: ENTITY WORK.NOR
    PORT MAP (
        A => S7078,
        B => S7275,
        Y => S7279
    );
NAND_4242: ENTITY WORK.NAND
    PORT MAP (
        A => S7077,
        B => S7274,
        Y => S7280
    );
NOR_2639: ENTITY WORK.NOR
    PORT MAP (
        A => S7276,
        B => S7279,
        Y => S7281
    );
NAND_4243: ENTITY WORK.NAND
    PORT MAP (
        A => S7277,
        B => S7280,
        Y => S7282
    );
NOR_2640: ENTITY WORK.NOR
    PORT MAP (
        A => S7273,
        B => S7282,
        Y => S7283
    );
NAND_4244: ENTITY WORK.NAND
    PORT MAP (
        A => S7272,
        B => S7281,
        Y => S7284
    );
NOR_2641: ENTITY WORK.NOR
    PORT MAP (
        A => S7272,
        B => S7281,
        Y => S7285
    );
NAND_4245: ENTITY WORK.NAND
    PORT MAP (
        A => S7273,
        B => S7282,
        Y => S7286
    );
NOR_2642: ENTITY WORK.NOR
    PORT MAP (
        A => S7283,
        B => S7285,
        Y => S7287
    );
NAND_4246: ENTITY WORK.NAND
    PORT MAP (
        A => S7284,
        B => S7286,
        Y => S7288
    );
NOR_2643: ENTITY WORK.NOR
    PORT MAP (
        A => S7270,
        B => S7288,
        Y => S7289
    );
NAND_4247: ENTITY WORK.NAND
    PORT MAP (
        A => S7271,
        B => S7287,
        Y => S7290
    );
NOR_2644: ENTITY WORK.NOR
    PORT MAP (
        A => S7271,
        B => S7287,
        Y => S7291
    );
NAND_4248: ENTITY WORK.NAND
    PORT MAP (
        A => S7270,
        B => S7288,
        Y => S7292
    );
NOR_2645: ENTITY WORK.NOR
    PORT MAP (
        A => S7289,
        B => S7291,
        Y => S7293
    );
NAND_4249: ENTITY WORK.NAND
    PORT MAP (
        A => S7290,
        B => S7292,
        Y => S7294
    );
NOR_2646: ENTITY WORK.NOR
    PORT MAP (
        A => S7269,
        B => S7294,
        Y => S7295
    );
NAND_4250: ENTITY WORK.NAND
    PORT MAP (
        A => S7268,
        B => S7293,
        Y => S7296
    );
NOR_2647: ENTITY WORK.NOR
    PORT MAP (
        A => S7268,
        B => S7293,
        Y => S7297
    );
NAND_4251: ENTITY WORK.NAND
    PORT MAP (
        A => S7269,
        B => S7294,
        Y => S7298
    );
NOR_2648: ENTITY WORK.NOR
    PORT MAP (
        A => S7295,
        B => S7297,
        Y => S7299
    );
NAND_4252: ENTITY WORK.NAND
    PORT MAP (
        A => S7296,
        B => S7298,
        Y => S7300
    );
NOR_2649: ENTITY WORK.NOR
    PORT MAP (
        A => S7251,
        B => S7300,
        Y => S7301
    );
NAND_4253: ENTITY WORK.NAND
    PORT MAP (
        A => S7252,
        B => S7299,
        Y => S7302
    );
NOR_2650: ENTITY WORK.NOR
    PORT MAP (
        A => S7252,
        B => S7299,
        Y => S7303
    );
NAND_4254: ENTITY WORK.NAND
    PORT MAP (
        A => S7251,
        B => S7300,
        Y => S7304
    );
NOR_2651: ENTITY WORK.NOR
    PORT MAP (
        A => S7301,
        B => S7303,
        Y => S7305
    );
NAND_4255: ENTITY WORK.NAND
    PORT MAP (
        A => S7302,
        B => S7304,
        Y => S7306
    );
NOR_2652: ENTITY WORK.NOR
    PORT MAP (
        A => S7250,
        B => S7306,
        Y => S7307
    );
NAND_4256: ENTITY WORK.NAND
    PORT MAP (
        A => S7249,
        B => S7305,
        Y => S7308
    );
NOR_2653: ENTITY WORK.NOR
    PORT MAP (
        A => S7249,
        B => S7305,
        Y => S7309
    );
NAND_4257: ENTITY WORK.NAND
    PORT MAP (
        A => S7250,
        B => S7306,
        Y => S7310
    );
NOR_2654: ENTITY WORK.NOR
    PORT MAP (
        A => S7307,
        B => S7309,
        Y => S7311
    );
NAND_4258: ENTITY WORK.NAND
    PORT MAP (
        A => S7308,
        B => S7310,
        Y => S7312
    );
NOR_2655: ENTITY WORK.NOR
    PORT MAP (
        A => S7215,
        B => S7312,
        Y => S7313
    );
NAND_4259: ENTITY WORK.NAND
    PORT MAP (
        A => S7216,
        B => S7311,
        Y => S7314
    );
NOR_2656: ENTITY WORK.NOR
    PORT MAP (
        A => S7216,
        B => S7311,
        Y => S7315
    );
NAND_4260: ENTITY WORK.NAND
    PORT MAP (
        A => S7215,
        B => S7312,
        Y => S7316
    );
NOR_2657: ENTITY WORK.NOR
    PORT MAP (
        A => S7313,
        B => S7315,
        Y => S7317
    );
NAND_4261: ENTITY WORK.NAND
    PORT MAP (
        A => S7314,
        B => S7316,
        Y => S7318
    );
NOR_2658: ENTITY WORK.NOR
    PORT MAP (
        A => S7214,
        B => S7318,
        Y => S7319
    );
NAND_4262: ENTITY WORK.NAND
    PORT MAP (
        A => S7213,
        B => S7317,
        Y => S7320
    );
NOR_2659: ENTITY WORK.NOR
    PORT MAP (
        A => S7213,
        B => S7317,
        Y => S7321
    );
NAND_4263: ENTITY WORK.NAND
    PORT MAP (
        A => S7214,
        B => S7318,
        Y => S7322
    );
NOR_2660: ENTITY WORK.NOR
    PORT MAP (
        A => S7319,
        B => S7321,
        Y => S7323
    );
NAND_4264: ENTITY WORK.NAND
    PORT MAP (
        A => S7320,
        B => S7322,
        Y => S7324
    );
NOR_2661: ENTITY WORK.NOR
    PORT MAP (
        A => S7154,
        B => S7324,
        Y => S7325
    );
NOT_522: ENTITY WORK.NOT
    PORT MAP (
        A => S7325,
        Y => S7326
    );
NOR_2662: ENTITY WORK.NOR
    PORT MAP (
        A => S7155,
        B => S7323,
        Y => S7327
    );
NAND_4265: ENTITY WORK.NAND
    PORT MAP (
        A => S7154,
        B => S7324,
        Y => S7328
    );
NOR_2663: ENTITY WORK.NOR
    PORT MAP (
        A => S7325,
        B => S7327,
        Y => S7329
    );
NAND_4266: ENTITY WORK.NAND
    PORT MAP (
        A => S7326,
        B => S7328,
        Y => S7330
    );
NOR_2664: ENTITY WORK.NOR
    PORT MAP (
        A => S7152,
        B => S7330,
        Y => S7331
    );
NOR_2665: ENTITY WORK.NOR
    PORT MAP (
        A => S7153,
        B => S7329,
        Y => S7332
    );
NOR_2666: ENTITY WORK.NOR
    PORT MAP (
        A => S7331,
        B => S7332,
        Y => S7333
    );
NOT_523: ENTITY WORK.NOT
    PORT MAP (
        A => S7333,
        Y => S7334
    );
NAND_4267: ENTITY WORK.NAND
    PORT MAP (
        A => S7150,
        B => S7334,
        Y => S7335
    );
NAND_4268: ENTITY WORK.NAND
    PORT MAP (
        A => S7151,
        B => S7333,
        Y => S7336
    );
NAND_4269: ENTITY WORK.NAND
    PORT MAP (
        A => S7335,
        B => S7336,
        Y => S7337
    );
NOR_2667: ENTITY WORK.NOR
    PORT MAP (
        A => S7138,
        B => S7337,
        Y => S7338
    );
NOT_524: ENTITY WORK.NOT
    PORT MAP (
        A => S7338,
        Y => S7339
    );
NAND_4270: ENTITY WORK.NAND
    PORT MAP (
        A => S7138,
        B => S7337,
        Y => S7340
    );
NAND_4271: ENTITY WORK.NAND
    PORT MAP (
        A => S7339,
        B => S7340,
        Y => S7341
    );
NOR_2668: ENTITY WORK.NOR
    PORT MAP (
        A => S7149,
        B => S7341,
        Y => S7342
    );
NAND_4272: ENTITY WORK.NAND
    PORT MAP (
        A => S7149,
        B => S7341,
        Y => S7343
    );
NOR_2669: ENTITY WORK.NOR
    PORT MAP (
        A => S5949,
        B => S7342,
        Y => S7344
    );
NAND_4273: ENTITY WORK.NAND
    PORT MAP (
        A => S7343,
        B => S7344,
        Y => S7345
    );
NAND_4274: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu1_13,
        B => S5950,
        Y => S7346
    );
NOT_525: ENTITY WORK.NOT
    PORT MAP (
        A => S7346,
        Y => S7347
    );
NOR_2670: ENTITY WORK.NOR
    PORT MAP (
        A => S3899,
        B => S3985,
        Y => S7348
    );
NOR_2671: ENTITY WORK.NOR
    PORT MAP (
        A => S7347,
        B => S7348,
        Y => S7349
    );
NAND_4275: ENTITY WORK.NAND
    PORT MAP (
        A => S7345,
        B => S7349,
        Y => S295
    );
NOR_2672: ENTITY WORK.NOR
    PORT MAP (
        A => S7325,
        B => S7331,
        Y => S7350
    );
NOT_526: ENTITY WORK.NOT
    PORT MAP (
        A => S7350,
        Y => S7351
    );
NOR_2673: ENTITY WORK.NOR
    PORT MAP (
        A => S7203,
        B => S7211,
        Y => S7352
    );
NOR_2674: ENTITY WORK.NOR
    PORT MAP (
        A => S7166,
        B => S7352,
        Y => S7353
    );
NOT_527: ENTITY WORK.NOT
    PORT MAP (
        A => S7353,
        Y => S7354
    );
NAND_4276: ENTITY WORK.NAND
    PORT MAP (
        A => S7166,
        B => S7352,
        Y => S7355
    );
NAND_4277: ENTITY WORK.NAND
    PORT MAP (
        A => S7354,
        B => S7355,
        Y => S7356
    );
NOT_528: ENTITY WORK.NOT
    PORT MAP (
        A => S7356,
        Y => S7357
    );
NOR_2675: ENTITY WORK.NOR
    PORT MAP (
        A => S7313,
        B => S7319,
        Y => S7358
    );
NAND_4278: ENTITY WORK.NAND
    PORT MAP (
        A => S7314,
        B => S7320,
        Y => S7359
    );
NOR_2676: ENTITY WORK.NOR
    PORT MAP (
        A => S7189,
        B => S7197,
        Y => S7360
    );
NAND_4279: ENTITY WORK.NAND
    PORT MAP (
        A => S7190,
        B => S7198,
        Y => S7361
    );
NAND_4280: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_0,
        B => S3036,
        Y => S7362
    );
NOT_529: ENTITY WORK.NOT
    PORT MAP (
        A => S7362,
        Y => S7363
    );
NOR_2677: ENTITY WORK.NOR
    PORT MAP (
        A => S1116,
        B => S2817,
        Y => S7364
    );
NOR_2678: ENTITY WORK.NOR
    PORT MAP (
        A => S7163,
        B => S7364,
        Y => S7365
    );
NOT_530: ENTITY WORK.NOT
    PORT MAP (
        A => S7365,
        Y => S7366
    );
NOR_2679: ENTITY WORK.NOR
    PORT MAP (
        A => S1116,
        B => S2920,
        Y => S7367
    );
NAND_4281: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_2,
        B => S2919,
        Y => S7368
    );
NOR_2680: ENTITY WORK.NOR
    PORT MAP (
        A => S7160,
        B => S7368,
        Y => S7369
    );
NAND_4282: ENTITY WORK.NAND
    PORT MAP (
        A => S7159,
        B => S7367,
        Y => S7370
    );
NOR_2681: ENTITY WORK.NOR
    PORT MAP (
        A => S7365,
        B => S7369,
        Y => S7371
    );
NAND_4283: ENTITY WORK.NAND
    PORT MAP (
        A => S7366,
        B => S7370,
        Y => S7372
    );
NOR_2682: ENTITY WORK.NOR
    PORT MAP (
        A => S7362,
        B => S7372,
        Y => S7373
    );
NAND_4284: ENTITY WORK.NAND
    PORT MAP (
        A => S7363,
        B => S7371,
        Y => S7374
    );
NOR_2683: ENTITY WORK.NOR
    PORT MAP (
        A => S7363,
        B => S7371,
        Y => S7375
    );
NAND_4285: ENTITY WORK.NAND
    PORT MAP (
        A => S7362,
        B => S7372,
        Y => S7376
    );
NOR_2684: ENTITY WORK.NOR
    PORT MAP (
        A => S7373,
        B => S7375,
        Y => S7377
    );
NAND_4286: ENTITY WORK.NAND
    PORT MAP (
        A => S7374,
        B => S7376,
        Y => S7378
    );
NOR_2685: ENTITY WORK.NOR
    PORT MAP (
        A => S7179,
        B => S7183,
        Y => S7379
    );
NAND_4287: ENTITY WORK.NAND
    PORT MAP (
        A => S7180,
        B => S7184,
        Y => S7380
    );
NOR_2686: ENTITY WORK.NOR
    PORT MAP (
        A => S1065,
        B => S2718,
        Y => S7381
    );
NAND_4288: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_3,
        B => S2717,
        Y => S7382
    );
NOR_2687: ENTITY WORK.NOR
    PORT MAP (
        A => S963,
        B => S2518,
        Y => S7383
    );
NAND_4289: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_5,
        B => S2517,
        Y => S7384
    );
NOR_2688: ENTITY WORK.NOR
    PORT MAP (
        A => S7177,
        B => S7383,
        Y => S7385
    );
NAND_4290: ENTITY WORK.NAND
    PORT MAP (
        A => S7178,
        B => S7384,
        Y => S7386
    );
NOR_2689: ENTITY WORK.NOR
    PORT MAP (
        A => S963,
        B => S2618,
        Y => S7387
    );
NAND_4291: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_5,
        B => S2617,
        Y => S7388
    );
NOR_2690: ENTITY WORK.NOR
    PORT MAP (
        A => S7174,
        B => S7388,
        Y => S7389
    );
NAND_4292: ENTITY WORK.NAND
    PORT MAP (
        A => S7173,
        B => S7387,
        Y => S7390
    );
NOR_2691: ENTITY WORK.NOR
    PORT MAP (
        A => S7385,
        B => S7389,
        Y => S7391
    );
NAND_4293: ENTITY WORK.NAND
    PORT MAP (
        A => S7386,
        B => S7390,
        Y => S7392
    );
NOR_2692: ENTITY WORK.NOR
    PORT MAP (
        A => S7382,
        B => S7392,
        Y => S7393
    );
NAND_4294: ENTITY WORK.NAND
    PORT MAP (
        A => S7381,
        B => S7391,
        Y => S7394
    );
NOR_2693: ENTITY WORK.NOR
    PORT MAP (
        A => S7381,
        B => S7391,
        Y => S7395
    );
NAND_4295: ENTITY WORK.NAND
    PORT MAP (
        A => S7382,
        B => S7392,
        Y => S7396
    );
NOR_2694: ENTITY WORK.NOR
    PORT MAP (
        A => S7393,
        B => S7395,
        Y => S7397
    );
NAND_4296: ENTITY WORK.NAND
    PORT MAP (
        A => S7394,
        B => S7396,
        Y => S7398
    );
NOR_2695: ENTITY WORK.NOR
    PORT MAP (
        A => S7379,
        B => S7398,
        Y => S7399
    );
NAND_4297: ENTITY WORK.NAND
    PORT MAP (
        A => S7380,
        B => S7397,
        Y => S7400
    );
NOR_2696: ENTITY WORK.NOR
    PORT MAP (
        A => S7380,
        B => S7397,
        Y => S7401
    );
NAND_4298: ENTITY WORK.NAND
    PORT MAP (
        A => S7379,
        B => S7398,
        Y => S7402
    );
NOR_2697: ENTITY WORK.NOR
    PORT MAP (
        A => S7399,
        B => S7401,
        Y => S7403
    );
NAND_4299: ENTITY WORK.NAND
    PORT MAP (
        A => S7400,
        B => S7402,
        Y => S7404
    );
NOR_2698: ENTITY WORK.NOR
    PORT MAP (
        A => S7377,
        B => S7403,
        Y => S7405
    );
NAND_4300: ENTITY WORK.NAND
    PORT MAP (
        A => S7378,
        B => S7404,
        Y => S7406
    );
NOR_2699: ENTITY WORK.NOR
    PORT MAP (
        A => S7378,
        B => S7404,
        Y => S7407
    );
NAND_4301: ENTITY WORK.NAND
    PORT MAP (
        A => S7377,
        B => S7403,
        Y => S7408
    );
NOR_2700: ENTITY WORK.NOR
    PORT MAP (
        A => S7405,
        B => S7407,
        Y => S7409
    );
NAND_4302: ENTITY WORK.NAND
    PORT MAP (
        A => S7406,
        B => S7408,
        Y => S7410
    );
NOR_2701: ENTITY WORK.NOR
    PORT MAP (
        A => S7239,
        B => S7247,
        Y => S7411
    );
NAND_4303: ENTITY WORK.NAND
    PORT MAP (
        A => S7240,
        B => S7248,
        Y => S7412
    );
NOR_2702: ENTITY WORK.NOR
    PORT MAP (
        A => S7410,
        B => S7411,
        Y => S7413
    );
NAND_4304: ENTITY WORK.NAND
    PORT MAP (
        A => S7409,
        B => S7412,
        Y => S7414
    );
NOR_2703: ENTITY WORK.NOR
    PORT MAP (
        A => S7409,
        B => S7412,
        Y => S7415
    );
NAND_4305: ENTITY WORK.NAND
    PORT MAP (
        A => S7410,
        B => S7411,
        Y => S7416
    );
NOR_2704: ENTITY WORK.NOR
    PORT MAP (
        A => S7413,
        B => S7415,
        Y => S7417
    );
NAND_4306: ENTITY WORK.NAND
    PORT MAP (
        A => S7414,
        B => S7416,
        Y => S7418
    );
NOR_2705: ENTITY WORK.NOR
    PORT MAP (
        A => S7361,
        B => S7417,
        Y => S7419
    );
NAND_4307: ENTITY WORK.NAND
    PORT MAP (
        A => S7360,
        B => S7418,
        Y => S7420
    );
NOR_2706: ENTITY WORK.NOR
    PORT MAP (
        A => S7360,
        B => S7418,
        Y => S7421
    );
NAND_4308: ENTITY WORK.NAND
    PORT MAP (
        A => S7361,
        B => S7417,
        Y => S7422
    );
NOR_2707: ENTITY WORK.NOR
    PORT MAP (
        A => S7419,
        B => S7421,
        Y => S7423
    );
NAND_4309: ENTITY WORK.NAND
    PORT MAP (
        A => S7420,
        B => S7422,
        Y => S7424
    );
NOR_2708: ENTITY WORK.NOR
    PORT MAP (
        A => S7301,
        B => S7307,
        Y => S7425
    );
NAND_4310: ENTITY WORK.NAND
    PORT MAP (
        A => S7302,
        B => S7308,
        Y => S7426
    );
NOR_2709: ENTITY WORK.NOR
    PORT MAP (
        A => S7227,
        B => S7231,
        Y => S7427
    );
NAND_4311: ENTITY WORK.NAND
    PORT MAP (
        A => S7228,
        B => S7232,
        Y => S7428
    );
NOR_2710: ENTITY WORK.NOR
    PORT MAP (
        A => S910,
        B => S2418,
        Y => S7429
    );
NAND_4312: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_6,
        B => S2417,
        Y => S7430
    );
NOR_2711: ENTITY WORK.NOR
    PORT MAP (
        A => S805,
        B => S2206,
        Y => S7431
    );
NAND_4313: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_8,
        B => S2205,
        Y => S7432
    );
NOR_2712: ENTITY WORK.NOR
    PORT MAP (
        A => S7225,
        B => S7431,
        Y => S7433
    );
NAND_4314: ENTITY WORK.NAND
    PORT MAP (
        A => S7226,
        B => S7432,
        Y => S7434
    );
NOR_2713: ENTITY WORK.NOR
    PORT MAP (
        A => S805,
        B => S2312,
        Y => S7435
    );
NAND_4315: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_8,
        B => S2311,
        Y => S7436
    );
NOR_2714: ENTITY WORK.NOR
    PORT MAP (
        A => S7222,
        B => S7436,
        Y => S7437
    );
NAND_4316: ENTITY WORK.NAND
    PORT MAP (
        A => S7221,
        B => S7435,
        Y => S7438
    );
NOR_2715: ENTITY WORK.NOR
    PORT MAP (
        A => S7433,
        B => S7437,
        Y => S7439
    );
NAND_4317: ENTITY WORK.NAND
    PORT MAP (
        A => S7434,
        B => S7438,
        Y => S7440
    );
NOR_2716: ENTITY WORK.NOR
    PORT MAP (
        A => S7430,
        B => S7440,
        Y => S7441
    );
NAND_4318: ENTITY WORK.NAND
    PORT MAP (
        A => S7429,
        B => S7439,
        Y => S7442
    );
NOR_2717: ENTITY WORK.NOR
    PORT MAP (
        A => S7429,
        B => S7439,
        Y => S7443
    );
NAND_4319: ENTITY WORK.NAND
    PORT MAP (
        A => S7430,
        B => S7440,
        Y => S7444
    );
NOR_2718: ENTITY WORK.NOR
    PORT MAP (
        A => S7441,
        B => S7443,
        Y => S7445
    );
NAND_4320: ENTITY WORK.NAND
    PORT MAP (
        A => S7442,
        B => S7444,
        Y => S7446
    );
NOR_2719: ENTITY WORK.NOR
    PORT MAP (
        A => S7260,
        B => S7264,
        Y => S7447
    );
NAND_4321: ENTITY WORK.NAND
    PORT MAP (
        A => S7261,
        B => S7265,
        Y => S7448
    );
NOR_2720: ENTITY WORK.NOR
    PORT MAP (
        A => S7446,
        B => S7447,
        Y => S7449
    );
NAND_4322: ENTITY WORK.NAND
    PORT MAP (
        A => S7445,
        B => S7448,
        Y => S7450
    );
NOR_2721: ENTITY WORK.NOR
    PORT MAP (
        A => S7445,
        B => S7448,
        Y => S7451
    );
NAND_4323: ENTITY WORK.NAND
    PORT MAP (
        A => S7446,
        B => S7447,
        Y => S7452
    );
NOR_2722: ENTITY WORK.NOR
    PORT MAP (
        A => S7449,
        B => S7451,
        Y => S7453
    );
NAND_4324: ENTITY WORK.NAND
    PORT MAP (
        A => S7450,
        B => S7452,
        Y => S7454
    );
NOR_2723: ENTITY WORK.NOR
    PORT MAP (
        A => S7428,
        B => S7453,
        Y => S7455
    );
NAND_4325: ENTITY WORK.NAND
    PORT MAP (
        A => S7427,
        B => S7454,
        Y => S7456
    );
NOR_2724: ENTITY WORK.NOR
    PORT MAP (
        A => S7427,
        B => S7454,
        Y => S7457
    );
NAND_4326: ENTITY WORK.NAND
    PORT MAP (
        A => S7428,
        B => S7453,
        Y => S7458
    );
NOR_2725: ENTITY WORK.NOR
    PORT MAP (
        A => S7455,
        B => S7457,
        Y => S7459
    );
NAND_4327: ENTITY WORK.NAND
    PORT MAP (
        A => S7456,
        B => S7458,
        Y => S7460
    );
NOR_2726: ENTITY WORK.NOR
    PORT MAP (
        A => S7289,
        B => S7295,
        Y => S7461
    );
NAND_4328: ENTITY WORK.NAND
    PORT MAP (
        A => S7290,
        B => S7296,
        Y => S7462
    );
NOR_2727: ENTITY WORK.NOR
    PORT MAP (
        A => S754,
        B => S2107,
        Y => S7463
    );
NAND_4329: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_9,
        B => S2106,
        Y => S7464
    );
NAND_4330: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_11,
        B => S1952,
        Y => S7465
    );
NAND_4331: ENTITY WORK.NAND
    PORT MAP (
        A => S7259,
        B => S7465,
        Y => S7466
    );
NOT_531: ENTITY WORK.NOT
    PORT MAP (
        A => S7466,
        Y => S7467
    );
NOR_2728: ENTITY WORK.NOR
    PORT MAP (
        A => S651,
        B => S1598,
        Y => S7468
    );
NAND_4332: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_11,
        B => S1597,
        Y => S7469
    );
NOR_2729: ENTITY WORK.NOR
    PORT MAP (
        A => S7256,
        B => S7469,
        Y => S7470
    );
NAND_4333: ENTITY WORK.NAND
    PORT MAP (
        A => S7255,
        B => S7468,
        Y => S7471
    );
NOR_2730: ENTITY WORK.NOR
    PORT MAP (
        A => S7467,
        B => S7470,
        Y => S7472
    );
NAND_4334: ENTITY WORK.NAND
    PORT MAP (
        A => S7466,
        B => S7471,
        Y => S7473
    );
NOR_2731: ENTITY WORK.NOR
    PORT MAP (
        A => S7464,
        B => S7473,
        Y => S7474
    );
NAND_4335: ENTITY WORK.NAND
    PORT MAP (
        A => S7463,
        B => S7472,
        Y => S7475
    );
NOR_2732: ENTITY WORK.NOR
    PORT MAP (
        A => S7463,
        B => S7472,
        Y => S7477
    );
NAND_4336: ENTITY WORK.NAND
    PORT MAP (
        A => S7464,
        B => S7473,
        Y => S7478
    );
NOR_2733: ENTITY WORK.NOR
    PORT MAP (
        A => S7474,
        B => S7477,
        Y => S7479
    );
NAND_4337: ENTITY WORK.NAND
    PORT MAP (
        A => S7475,
        B => S7478,
        Y => S7480
    );
NOR_2734: ENTITY WORK.NOR
    PORT MAP (
        A => S7279,
        B => S7283,
        Y => S7481
    );
NAND_4338: ENTITY WORK.NAND
    PORT MAP (
        A => S7280,
        B => S7284,
        Y => S7482
    );
NOR_2735: ENTITY WORK.NOR
    PORT MAP (
        A => S599,
        B => S1849,
        Y => S7483
    );
NAND_4339: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_12,
        B => S1848,
        Y => S7484
    );
NAND_4340: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_14,
        B => S1515,
        Y => S7485
    );
NAND_4341: ENTITY WORK.NAND
    PORT MAP (
        A => S7278,
        B => S7485,
        Y => S7486
    );
NOT_532: ENTITY WORK.NOT
    PORT MAP (
        A => S7486,
        Y => S7488
    );
NOR_2736: ENTITY WORK.NOR
    PORT MAP (
        A => S492,
        B => S1746,
        Y => S7489
    );
NAND_4342: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_14,
        B => S1745,
        Y => S7490
    );
NOR_2737: ENTITY WORK.NOR
    PORT MAP (
        A => S7275,
        B => S7490,
        Y => S7491
    );
NAND_4343: ENTITY WORK.NAND
    PORT MAP (
        A => S7274,
        B => S7489,
        Y => S7492
    );
NOR_2738: ENTITY WORK.NOR
    PORT MAP (
        A => S7488,
        B => S7491,
        Y => S7493
    );
NAND_4344: ENTITY WORK.NAND
    PORT MAP (
        A => S7486,
        B => S7492,
        Y => S7494
    );
NOR_2739: ENTITY WORK.NOR
    PORT MAP (
        A => S7484,
        B => S7494,
        Y => S7495
    );
NAND_4345: ENTITY WORK.NAND
    PORT MAP (
        A => S7483,
        B => S7493,
        Y => S7496
    );
NOR_2740: ENTITY WORK.NOR
    PORT MAP (
        A => S7483,
        B => S7493,
        Y => S7497
    );
NAND_4346: ENTITY WORK.NAND
    PORT MAP (
        A => S7484,
        B => S7494,
        Y => S7499
    );
NOR_2741: ENTITY WORK.NOR
    PORT MAP (
        A => S7495,
        B => S7497,
        Y => S7500
    );
NAND_4347: ENTITY WORK.NAND
    PORT MAP (
        A => S7496,
        B => S7499,
        Y => S7501
    );
NOR_2742: ENTITY WORK.NOR
    PORT MAP (
        A => S7481,
        B => S7501,
        Y => S7502
    );
NAND_4348: ENTITY WORK.NAND
    PORT MAP (
        A => S7482,
        B => S7500,
        Y => S7503
    );
NOR_2743: ENTITY WORK.NOR
    PORT MAP (
        A => S7482,
        B => S7500,
        Y => S7504
    );
NAND_4349: ENTITY WORK.NAND
    PORT MAP (
        A => S7481,
        B => S7501,
        Y => S7505
    );
NOR_2744: ENTITY WORK.NOR
    PORT MAP (
        A => S7502,
        B => S7504,
        Y => S7506
    );
NAND_4350: ENTITY WORK.NAND
    PORT MAP (
        A => S7503,
        B => S7505,
        Y => S7507
    );
NOR_2745: ENTITY WORK.NOR
    PORT MAP (
        A => S7480,
        B => S7507,
        Y => S7508
    );
NAND_4351: ENTITY WORK.NAND
    PORT MAP (
        A => S7479,
        B => S7506,
        Y => S7510
    );
NOR_2746: ENTITY WORK.NOR
    PORT MAP (
        A => S7479,
        B => S7506,
        Y => S7511
    );
NAND_4352: ENTITY WORK.NAND
    PORT MAP (
        A => S7480,
        B => S7507,
        Y => S7512
    );
NOR_2747: ENTITY WORK.NOR
    PORT MAP (
        A => S7508,
        B => S7511,
        Y => S7513
    );
NAND_4353: ENTITY WORK.NAND
    PORT MAP (
        A => S7510,
        B => S7512,
        Y => S7514
    );
NOR_2748: ENTITY WORK.NOR
    PORT MAP (
        A => S7461,
        B => S7514,
        Y => S7515
    );
NAND_4354: ENTITY WORK.NAND
    PORT MAP (
        A => S7462,
        B => S7513,
        Y => S7516
    );
NOR_2749: ENTITY WORK.NOR
    PORT MAP (
        A => S7462,
        B => S7513,
        Y => S7517
    );
NAND_4355: ENTITY WORK.NAND
    PORT MAP (
        A => S7461,
        B => S7514,
        Y => S7518
    );
NOR_2750: ENTITY WORK.NOR
    PORT MAP (
        A => S7515,
        B => S7517,
        Y => S7519
    );
NAND_4356: ENTITY WORK.NAND
    PORT MAP (
        A => S7516,
        B => S7518,
        Y => S7521
    );
NOR_2751: ENTITY WORK.NOR
    PORT MAP (
        A => S7460,
        B => S7521,
        Y => S7522
    );
NAND_4357: ENTITY WORK.NAND
    PORT MAP (
        A => S7459,
        B => S7519,
        Y => S7523
    );
NOR_2752: ENTITY WORK.NOR
    PORT MAP (
        A => S7459,
        B => S7519,
        Y => S7524
    );
NAND_4358: ENTITY WORK.NAND
    PORT MAP (
        A => S7460,
        B => S7521,
        Y => S7525
    );
NOR_2753: ENTITY WORK.NOR
    PORT MAP (
        A => S7522,
        B => S7524,
        Y => S7526
    );
NAND_4359: ENTITY WORK.NAND
    PORT MAP (
        A => S7523,
        B => S7525,
        Y => S7527
    );
NOR_2754: ENTITY WORK.NOR
    PORT MAP (
        A => S7425,
        B => S7527,
        Y => S7528
    );
NAND_4360: ENTITY WORK.NAND
    PORT MAP (
        A => S7426,
        B => S7526,
        Y => S7529
    );
NOR_2755: ENTITY WORK.NOR
    PORT MAP (
        A => S7426,
        B => S7526,
        Y => S7530
    );
NAND_4361: ENTITY WORK.NAND
    PORT MAP (
        A => S7425,
        B => S7527,
        Y => S7532
    );
NOR_2756: ENTITY WORK.NOR
    PORT MAP (
        A => S7528,
        B => S7530,
        Y => S7533
    );
NAND_4362: ENTITY WORK.NAND
    PORT MAP (
        A => S7529,
        B => S7532,
        Y => S7534
    );
NOR_2757: ENTITY WORK.NOR
    PORT MAP (
        A => S7424,
        B => S7534,
        Y => S7535
    );
NAND_4363: ENTITY WORK.NAND
    PORT MAP (
        A => S7423,
        B => S7533,
        Y => S7536
    );
NOR_2758: ENTITY WORK.NOR
    PORT MAP (
        A => S7423,
        B => S7533,
        Y => S7537
    );
NAND_4364: ENTITY WORK.NAND
    PORT MAP (
        A => S7424,
        B => S7534,
        Y => S7538
    );
NOR_2759: ENTITY WORK.NOR
    PORT MAP (
        A => S7535,
        B => S7537,
        Y => S7539
    );
NAND_4365: ENTITY WORK.NAND
    PORT MAP (
        A => S7536,
        B => S7538,
        Y => S7540
    );
NOR_2760: ENTITY WORK.NOR
    PORT MAP (
        A => S7358,
        B => S7540,
        Y => S7541
    );
NAND_4366: ENTITY WORK.NAND
    PORT MAP (
        A => S7359,
        B => S7539,
        Y => S7543
    );
NAND_4367: ENTITY WORK.NAND
    PORT MAP (
        A => S7358,
        B => S7540,
        Y => S7544
    );
NAND_4368: ENTITY WORK.NAND
    PORT MAP (
        A => S7543,
        B => S7544,
        Y => S7545
    );
NOT_533: ENTITY WORK.NOT
    PORT MAP (
        A => S7545,
        Y => S7546
    );
NAND_4369: ENTITY WORK.NAND
    PORT MAP (
        A => S7357,
        B => S7546,
        Y => S7547
    );
NOT_534: ENTITY WORK.NOT
    PORT MAP (
        A => S7547,
        Y => S7548
    );
NAND_4370: ENTITY WORK.NAND
    PORT MAP (
        A => S7356,
        B => S7545,
        Y => S7549
    );
NAND_4371: ENTITY WORK.NAND
    PORT MAP (
        A => S7547,
        B => S7549,
        Y => S7550
    );
NOT_535: ENTITY WORK.NOT
    PORT MAP (
        A => S7550,
        Y => S7551
    );
NAND_4372: ENTITY WORK.NAND
    PORT MAP (
        A => S7350,
        B => S7550,
        Y => S7552
    );
NAND_4373: ENTITY WORK.NAND
    PORT MAP (
        A => S7351,
        B => S7551,
        Y => S7554
    );
NAND_4374: ENTITY WORK.NAND
    PORT MAP (
        A => S7552,
        B => S7554,
        Y => S7555
    );
NOR_2761: ENTITY WORK.NOR
    PORT MAP (
        A => S7336,
        B => S7555,
        Y => S7556
    );
NOT_536: ENTITY WORK.NOT
    PORT MAP (
        A => S7556,
        Y => S7557
    );
NAND_4375: ENTITY WORK.NAND
    PORT MAP (
        A => S7336,
        B => S7555,
        Y => S7558
    );
NAND_4376: ENTITY WORK.NAND
    PORT MAP (
        A => S7557,
        B => S7558,
        Y => S7559
    );
NOR_2762: ENTITY WORK.NOR
    PORT MAP (
        A => S7338,
        B => S7342,
        Y => S7560
    );
NAND_4377: ENTITY WORK.NAND
    PORT MAP (
        A => S7559,
        B => S7560,
        Y => S7561
    );
NOR_2763: ENTITY WORK.NOR
    PORT MAP (
        A => S7559,
        B => S7560,
        Y => S7562
    );
NOR_2764: ENTITY WORK.NOR
    PORT MAP (
        A => S5949,
        B => S7562,
        Y => S7563
    );
NAND_4378: ENTITY WORK.NAND
    PORT MAP (
        A => S7561,
        B => S7563,
        Y => S7565
    );
NAND_4379: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu1_14,
        B => S5950,
        Y => S7566
    );
NOT_537: ENTITY WORK.NOT
    PORT MAP (
        A => S7566,
        Y => S7567
    );
NOR_2765: ENTITY WORK.NOR
    PORT MAP (
        A => S3899,
        B => S3945,
        Y => S7568
    );
NOR_2766: ENTITY WORK.NOR
    PORT MAP (
        A => S7567,
        B => S7568,
        Y => S7569
    );
NAND_4380: ENTITY WORK.NAND
    PORT MAP (
        A => S7565,
        B => S7569,
        Y => S296
    );
NOR_2767: ENTITY WORK.NOR
    PORT MAP (
        A => S7556,
        B => S7562,
        Y => S7570
    );
NOR_2768: ENTITY WORK.NOR
    PORT MAP (
        A => S7541,
        B => S7548,
        Y => S7571
    );
NAND_4381: ENTITY WORK.NAND
    PORT MAP (
        A => S7543,
        B => S7547,
        Y => S7572
    );
NOR_2769: ENTITY WORK.NOR
    PORT MAP (
        A => S7449,
        B => S7457,
        Y => S7573
    );
NAND_4382: ENTITY WORK.NAND
    PORT MAP (
        A => S7450,
        B => S7458,
        Y => S7575
    );
NOR_2770: ENTITY WORK.NOR
    PORT MAP (
        A => S548,
        B => S1849,
        Y => S7576
    );
NAND_4383: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_13,
        B => S1848,
        Y => S7577
    );
NOR_2771: ENTITY WORK.NOR
    PORT MAP (
        A => S1304,
        B => S1516,
        Y => S7578
    );
NAND_4384: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_15,
        B => S1515,
        Y => S7579
    );
NOR_2772: ENTITY WORK.NOR
    PORT MAP (
        A => S7490,
        B => S7578,
        Y => S7580
    );
NAND_4385: ENTITY WORK.NAND
    PORT MAP (
        A => S7489,
        B => S7579,
        Y => S7581
    );
NOR_2773: ENTITY WORK.NOR
    PORT MAP (
        A => S7489,
        B => S7579,
        Y => S7582
    );
NAND_4386: ENTITY WORK.NAND
    PORT MAP (
        A => S7490,
        B => S7578,
        Y => S7583
    );
NOR_2774: ENTITY WORK.NOR
    PORT MAP (
        A => S7580,
        B => S7582,
        Y => S7584
    );
NAND_4387: ENTITY WORK.NAND
    PORT MAP (
        A => S7581,
        B => S7583,
        Y => S7586
    );
NOR_2775: ENTITY WORK.NOR
    PORT MAP (
        A => S599,
        B => S1953,
        Y => S7587
    );
NAND_4388: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_12,
        B => S1952,
        Y => S7588
    );
NOR_2776: ENTITY WORK.NOR
    PORT MAP (
        A => S7469,
        B => S7587,
        Y => S7589
    );
NAND_4389: ENTITY WORK.NAND
    PORT MAP (
        A => S7468,
        B => S7588,
        Y => S7590
    );
NOR_2777: ENTITY WORK.NOR
    PORT MAP (
        A => S7468,
        B => S7588,
        Y => S7591
    );
NAND_4390: ENTITY WORK.NAND
    PORT MAP (
        A => S7469,
        B => S7587,
        Y => S7592
    );
NOR_2778: ENTITY WORK.NOR
    PORT MAP (
        A => S7589,
        B => S7591,
        Y => S7593
    );
NAND_4391: ENTITY WORK.NAND
    PORT MAP (
        A => S7590,
        B => S7592,
        Y => S7594
    );
NOR_2779: ENTITY WORK.NOR
    PORT MAP (
        A => S7584,
        B => S7593,
        Y => S7595
    );
NAND_4392: ENTITY WORK.NAND
    PORT MAP (
        A => S7586,
        B => S7594,
        Y => S7597
    );
NOR_2780: ENTITY WORK.NOR
    PORT MAP (
        A => S7586,
        B => S7594,
        Y => S7598
    );
NAND_4393: ENTITY WORK.NAND
    PORT MAP (
        A => S7584,
        B => S7593,
        Y => S7599
    );
NOR_2781: ENTITY WORK.NOR
    PORT MAP (
        A => S7595,
        B => S7598,
        Y => S7600
    );
NAND_4394: ENTITY WORK.NAND
    PORT MAP (
        A => S7597,
        B => S7599,
        Y => S7601
    );
NOR_2782: ENTITY WORK.NOR
    PORT MAP (
        A => S7576,
        B => S7601,
        Y => S7602
    );
NAND_4395: ENTITY WORK.NAND
    PORT MAP (
        A => S7577,
        B => S7600,
        Y => S7603
    );
NOR_2783: ENTITY WORK.NOR
    PORT MAP (
        A => S7577,
        B => S7600,
        Y => S7604
    );
NAND_4396: ENTITY WORK.NAND
    PORT MAP (
        A => S7576,
        B => S7601,
        Y => S7605
    );
NOR_2784: ENTITY WORK.NOR
    PORT MAP (
        A => S7602,
        B => S7604,
        Y => S7606
    );
NAND_4397: ENTITY WORK.NAND
    PORT MAP (
        A => S7603,
        B => S7605,
        Y => S7608
    );
NOR_2785: ENTITY WORK.NOR
    PORT MAP (
        A => S702,
        B => S2107,
        Y => S7609
    );
NAND_4398: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_10,
        B => S2106,
        Y => S7610
    );
NOR_2786: ENTITY WORK.NOR
    PORT MAP (
        A => S7491,
        B => S7495,
        Y => S7611
    );
NAND_4399: ENTITY WORK.NAND
    PORT MAP (
        A => S7492,
        B => S7496,
        Y => S7612
    );
NOR_2787: ENTITY WORK.NOR
    PORT MAP (
        A => S7609,
        B => S7611,
        Y => S7613
    );
NAND_4400: ENTITY WORK.NAND
    PORT MAP (
        A => S7610,
        B => S7612,
        Y => S7614
    );
NOR_2788: ENTITY WORK.NOR
    PORT MAP (
        A => S7610,
        B => S7612,
        Y => S7615
    );
NAND_4401: ENTITY WORK.NAND
    PORT MAP (
        A => S7609,
        B => S7611,
        Y => S7616
    );
NOR_2789: ENTITY WORK.NOR
    PORT MAP (
        A => S7613,
        B => S7615,
        Y => S7617
    );
NAND_4402: ENTITY WORK.NAND
    PORT MAP (
        A => S7614,
        B => S7616,
        Y => S7619
    );
NOR_2790: ENTITY WORK.NOR
    PORT MAP (
        A => S7470,
        B => S7474,
        Y => S7620
    );
NAND_4403: ENTITY WORK.NAND
    PORT MAP (
        A => S7471,
        B => S7475,
        Y => S7621
    );
NOR_2791: ENTITY WORK.NOR
    PORT MAP (
        A => S858,
        B => S2418,
        Y => S7622
    );
NAND_4404: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_7,
        B => S2417,
        Y => S7623
    );
NOR_2792: ENTITY WORK.NOR
    PORT MAP (
        A => S754,
        B => S2206,
        Y => S7624
    );
NAND_4405: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_9,
        B => S2205,
        Y => S7625
    );
NOR_2793: ENTITY WORK.NOR
    PORT MAP (
        A => S7435,
        B => S7625,
        Y => S7626
    );
NAND_4406: ENTITY WORK.NAND
    PORT MAP (
        A => S7436,
        B => S7624,
        Y => S7627
    );
NOR_2794: ENTITY WORK.NOR
    PORT MAP (
        A => S7436,
        B => S7624,
        Y => S7628
    );
NAND_4407: ENTITY WORK.NAND
    PORT MAP (
        A => S7435,
        B => S7625,
        Y => S7630
    );
NOR_2795: ENTITY WORK.NOR
    PORT MAP (
        A => S7626,
        B => S7628,
        Y => S7631
    );
NAND_4408: ENTITY WORK.NAND
    PORT MAP (
        A => S7627,
        B => S7630,
        Y => S7632
    );
NOR_2796: ENTITY WORK.NOR
    PORT MAP (
        A => S7623,
        B => S7632,
        Y => S7633
    );
NAND_4409: ENTITY WORK.NAND
    PORT MAP (
        A => S7622,
        B => S7631,
        Y => S7634
    );
NOR_2797: ENTITY WORK.NOR
    PORT MAP (
        A => S7622,
        B => S7631,
        Y => S7635
    );
NAND_4410: ENTITY WORK.NAND
    PORT MAP (
        A => S7623,
        B => S7632,
        Y => S7636
    );
NOR_2798: ENTITY WORK.NOR
    PORT MAP (
        A => S7633,
        B => S7635,
        Y => S7637
    );
NAND_4411: ENTITY WORK.NAND
    PORT MAP (
        A => S7634,
        B => S7636,
        Y => S7638
    );
NOR_2799: ENTITY WORK.NOR
    PORT MAP (
        A => S7620,
        B => S7637,
        Y => S7639
    );
NAND_4412: ENTITY WORK.NAND
    PORT MAP (
        A => S7621,
        B => S7638,
        Y => S7641
    );
NOR_2800: ENTITY WORK.NOR
    PORT MAP (
        A => S7621,
        B => S7638,
        Y => S7642
    );
NAND_4413: ENTITY WORK.NAND
    PORT MAP (
        A => S7620,
        B => S7637,
        Y => S7643
    );
NOR_2801: ENTITY WORK.NOR
    PORT MAP (
        A => S7639,
        B => S7642,
        Y => S7644
    );
NAND_4414: ENTITY WORK.NAND
    PORT MAP (
        A => S7641,
        B => S7643,
        Y => S7645
    );
NOR_2802: ENTITY WORK.NOR
    PORT MAP (
        A => S7617,
        B => S7645,
        Y => S7646
    );
NAND_4415: ENTITY WORK.NAND
    PORT MAP (
        A => S7619,
        B => S7644,
        Y => S7647
    );
NOR_2803: ENTITY WORK.NOR
    PORT MAP (
        A => S7619,
        B => S7644,
        Y => S7648
    );
NAND_4416: ENTITY WORK.NAND
    PORT MAP (
        A => S7617,
        B => S7645,
        Y => S7649
    );
NOR_2804: ENTITY WORK.NOR
    PORT MAP (
        A => S7646,
        B => S7648,
        Y => S7650
    );
NAND_4417: ENTITY WORK.NAND
    PORT MAP (
        A => S7647,
        B => S7649,
        Y => S7652
    );
NOR_2805: ENTITY WORK.NOR
    PORT MAP (
        A => S7606,
        B => S7650,
        Y => S7653
    );
NAND_4418: ENTITY WORK.NAND
    PORT MAP (
        A => S7608,
        B => S7652,
        Y => S7654
    );
NOR_2806: ENTITY WORK.NOR
    PORT MAP (
        A => S7608,
        B => S7652,
        Y => S7655
    );
NAND_4419: ENTITY WORK.NAND
    PORT MAP (
        A => S7606,
        B => S7650,
        Y => S7656
    );
NOR_2807: ENTITY WORK.NOR
    PORT MAP (
        A => S7653,
        B => S7655,
        Y => S7657
    );
NAND_4420: ENTITY WORK.NAND
    PORT MAP (
        A => S7654,
        B => S7656,
        Y => S7658
    );
NOR_2808: ENTITY WORK.NOR
    PORT MAP (
        A => S7573,
        B => S7657,
        Y => S7659
    );
NAND_4421: ENTITY WORK.NAND
    PORT MAP (
        A => S7575,
        B => S7658,
        Y => S7660
    );
NOR_2809: ENTITY WORK.NOR
    PORT MAP (
        A => S7575,
        B => S7658,
        Y => S7661
    );
NAND_4422: ENTITY WORK.NAND
    PORT MAP (
        A => S7573,
        B => S7657,
        Y => S7663
    );
NOR_2810: ENTITY WORK.NOR
    PORT MAP (
        A => S7659,
        B => S7661,
        Y => S7664
    );
NAND_4423: ENTITY WORK.NAND
    PORT MAP (
        A => S7660,
        B => S7663,
        Y => S7665
    );
NOR_2811: ENTITY WORK.NOR
    PORT MAP (
        A => S1065,
        B => S2817,
        Y => S7666
    );
NAND_4424: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_3,
        B => S2816,
        Y => S7667
    );
NOR_2812: ENTITY WORK.NOR
    PORT MAP (
        A => S7367,
        B => S7667,
        Y => S7668
    );
NAND_4425: ENTITY WORK.NAND
    PORT MAP (
        A => S7368,
        B => S7666,
        Y => S7669
    );
NOR_2813: ENTITY WORK.NOR
    PORT MAP (
        A => S7368,
        B => S7666,
        Y => S7670
    );
NAND_4426: ENTITY WORK.NAND
    PORT MAP (
        A => S7367,
        B => S7667,
        Y => S7671
    );
NOR_2814: ENTITY WORK.NOR
    PORT MAP (
        A => S7668,
        B => S7670,
        Y => S7672
    );
NAND_4427: ENTITY WORK.NAND
    PORT MAP (
        A => S7669,
        B => S7671,
        Y => S7674
    );
NOR_2815: ENTITY WORK.NOR
    PORT MAP (
        A => S910,
        B => S2518,
        Y => S7675
    );
NAND_4428: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_6,
        B => S2517,
        Y => S7676
    );
NOR_2816: ENTITY WORK.NOR
    PORT MAP (
        A => S7387,
        B => S7675,
        Y => S7677
    );
NAND_4429: ENTITY WORK.NAND
    PORT MAP (
        A => S7388,
        B => S7676,
        Y => S7678
    );
NOR_2817: ENTITY WORK.NOR
    PORT MAP (
        A => S7388,
        B => S7676,
        Y => S7679
    );
NAND_4430: ENTITY WORK.NAND
    PORT MAP (
        A => S7387,
        B => S7675,
        Y => S7680
    );
NOR_2818: ENTITY WORK.NOR
    PORT MAP (
        A => S7677,
        B => S7679,
        Y => S7681
    );
NAND_4431: ENTITY WORK.NAND
    PORT MAP (
        A => S7678,
        B => S7680,
        Y => S7682
    );
NOR_2819: ENTITY WORK.NOR
    PORT MAP (
        A => S1013,
        B => S2718,
        Y => S7683
    );
NAND_4432: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_4,
        B => S2717,
        Y => S7685
    );
NOR_2820: ENTITY WORK.NOR
    PORT MAP (
        A => S7672,
        B => S7685,
        Y => S7686
    );
NAND_4433: ENTITY WORK.NAND
    PORT MAP (
        A => S7674,
        B => S7683,
        Y => S7687
    );
NOR_2821: ENTITY WORK.NOR
    PORT MAP (
        A => S7674,
        B => S7683,
        Y => S7688
    );
NAND_4434: ENTITY WORK.NAND
    PORT MAP (
        A => S7672,
        B => S7685,
        Y => S7689
    );
NOR_2822: ENTITY WORK.NOR
    PORT MAP (
        A => S7686,
        B => S7688,
        Y => S7690
    );
NAND_4435: ENTITY WORK.NAND
    PORT MAP (
        A => S7687,
        B => S7689,
        Y => S7691
    );
NOR_2823: ENTITY WORK.NOR
    PORT MAP (
        A => S7682,
        B => S7691,
        Y => S7692
    );
NAND_4436: ENTITY WORK.NAND
    PORT MAP (
        A => S7681,
        B => S7690,
        Y => S7693
    );
NOR_2824: ENTITY WORK.NOR
    PORT MAP (
        A => S7681,
        B => S7690,
        Y => S7694
    );
NAND_4437: ENTITY WORK.NAND
    PORT MAP (
        A => S7682,
        B => S7691,
        Y => S7696
    );
NAND_4438: ENTITY WORK.NAND
    PORT MAP (
        A => S7693,
        B => S7696,
        Y => S7697
    );
NOR_2825: ENTITY WORK.NOR
    PORT MAP (
        A => S7692,
        B => S7694,
        Y => S7698
    );
NAND_4439: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_1,
        B => S3036,
        Y => S7699
    );
NOT_538: ENTITY WORK.NOT
    PORT MAP (
        A => S7699,
        Y => S7700
    );
NOR_2826: ENTITY WORK.NOR
    PORT MAP (
        A => S7389,
        B => S7393,
        Y => S7701
    );
NAND_4440: ENTITY WORK.NAND
    PORT MAP (
        A => S7390,
        B => S7394,
        Y => S7702
    );
NOR_2827: ENTITY WORK.NOR
    PORT MAP (
        A => S7699,
        B => S7702,
        Y => S7703
    );
NAND_4441: ENTITY WORK.NAND
    PORT MAP (
        A => S7700,
        B => S7701,
        Y => S7704
    );
NOR_2828: ENTITY WORK.NOR
    PORT MAP (
        A => S7700,
        B => S7701,
        Y => S7705
    );
NAND_4442: ENTITY WORK.NAND
    PORT MAP (
        A => S7699,
        B => S7702,
        Y => S7707
    );
NOR_2829: ENTITY WORK.NOR
    PORT MAP (
        A => S7703,
        B => S7705,
        Y => S7708
    );
NAND_4443: ENTITY WORK.NAND
    PORT MAP (
        A => S7704,
        B => S7707,
        Y => S7709
    );
NOR_2830: ENTITY WORK.NOR
    PORT MAP (
        A => S7697,
        B => S7709,
        Y => S7710
    );
NAND_4444: ENTITY WORK.NAND
    PORT MAP (
        A => S7698,
        B => S7708,
        Y => S7711
    );
NOR_2831: ENTITY WORK.NOR
    PORT MAP (
        A => S7698,
        B => S7708,
        Y => S7712
    );
NAND_4445: ENTITY WORK.NAND
    PORT MAP (
        A => S7697,
        B => S7709,
        Y => S7713
    );
NOR_2832: ENTITY WORK.NOR
    PORT MAP (
        A => S7710,
        B => S7712,
        Y => S7714
    );
NAND_4446: ENTITY WORK.NAND
    PORT MAP (
        A => S7711,
        B => S7713,
        Y => S7715
    );
NOR_2833: ENTITY WORK.NOR
    PORT MAP (
        A => S7437,
        B => S7441,
        Y => S7716
    );
NAND_4447: ENTITY WORK.NAND
    PORT MAP (
        A => S7438,
        B => S7442,
        Y => S7718
    );
NOR_2834: ENTITY WORK.NOR
    PORT MAP (
        A => S7502,
        B => S7508,
        Y => S7719
    );
NAND_4448: ENTITY WORK.NAND
    PORT MAP (
        A => S7503,
        B => S7510,
        Y => S7720
    );
NOR_2835: ENTITY WORK.NOR
    PORT MAP (
        A => S7718,
        B => S7720,
        Y => S7721
    );
NAND_4449: ENTITY WORK.NAND
    PORT MAP (
        A => S7716,
        B => S7719,
        Y => S7722
    );
NOR_2836: ENTITY WORK.NOR
    PORT MAP (
        A => S7716,
        B => S7719,
        Y => S7723
    );
NAND_4450: ENTITY WORK.NAND
    PORT MAP (
        A => S7718,
        B => S7720,
        Y => S7724
    );
NOR_2837: ENTITY WORK.NOR
    PORT MAP (
        A => S7721,
        B => S7723,
        Y => S7725
    );
NAND_4451: ENTITY WORK.NAND
    PORT MAP (
        A => S7722,
        B => S7724,
        Y => S7726
    );
NOR_2838: ENTITY WORK.NOR
    PORT MAP (
        A => S7714,
        B => S7726,
        Y => S7727
    );
NAND_4452: ENTITY WORK.NAND
    PORT MAP (
        A => S7715,
        B => S7725,
        Y => S7729
    );
NOR_2839: ENTITY WORK.NOR
    PORT MAP (
        A => S7715,
        B => S7725,
        Y => S7730
    );
NAND_4453: ENTITY WORK.NAND
    PORT MAP (
        A => S7714,
        B => S7726,
        Y => S7731
    );
NOR_2840: ENTITY WORK.NOR
    PORT MAP (
        A => S7727,
        B => S7730,
        Y => S7732
    );
NAND_4454: ENTITY WORK.NAND
    PORT MAP (
        A => S7729,
        B => S7731,
        Y => S7733
    );
NOR_2841: ENTITY WORK.NOR
    PORT MAP (
        A => S7664,
        B => S7733,
        Y => S7734
    );
NAND_4455: ENTITY WORK.NAND
    PORT MAP (
        A => S7665,
        B => S7732,
        Y => S7735
    );
NOR_2842: ENTITY WORK.NOR
    PORT MAP (
        A => S7665,
        B => S7732,
        Y => S7736
    );
NAND_4456: ENTITY WORK.NAND
    PORT MAP (
        A => S7664,
        B => S7733,
        Y => S7737
    );
NOR_2843: ENTITY WORK.NOR
    PORT MAP (
        A => S7734,
        B => S7736,
        Y => S7738
    );
NAND_4457: ENTITY WORK.NAND
    PORT MAP (
        A => S7735,
        B => S7737,
        Y => S7740
    );
NOR_2844: ENTITY WORK.NOR
    PORT MAP (
        A => S7528,
        B => S7535,
        Y => S7741
    );
NAND_4458: ENTITY WORK.NAND
    PORT MAP (
        A => S7529,
        B => S7536,
        Y => S7742
    );
NOR_2845: ENTITY WORK.NOR
    PORT MAP (
        A => S7515,
        B => S7522,
        Y => S7743
    );
NAND_4459: ENTITY WORK.NAND
    PORT MAP (
        A => S7516,
        B => S7523,
        Y => S7744
    );
NOR_2846: ENTITY WORK.NOR
    PORT MAP (
        A => S1220,
        B => S3142,
        Y => S7745
    );
NAND_4460: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_0,
        B => S3141,
        Y => S7746
    );
NOR_2847: ENTITY WORK.NOR
    PORT MAP (
        A => S7369,
        B => S7373,
        Y => S7747
    );
NAND_4461: ENTITY WORK.NAND
    PORT MAP (
        A => S7370,
        B => S7374,
        Y => S7748
    );
NOR_2848: ENTITY WORK.NOR
    PORT MAP (
        A => S7745,
        B => S7748,
        Y => S7749
    );
NAND_4462: ENTITY WORK.NAND
    PORT MAP (
        A => S7746,
        B => S7747,
        Y => S7751
    );
NOR_2849: ENTITY WORK.NOR
    PORT MAP (
        A => S7746,
        B => S7747,
        Y => S7752
    );
NAND_4463: ENTITY WORK.NAND
    PORT MAP (
        A => S7745,
        B => S7748,
        Y => S7753
    );
NOR_2850: ENTITY WORK.NOR
    PORT MAP (
        A => S7749,
        B => S7752,
        Y => S7754
    );
NAND_4464: ENTITY WORK.NAND
    PORT MAP (
        A => S7751,
        B => S7753,
        Y => S7755
    );
NOR_2851: ENTITY WORK.NOR
    PORT MAP (
        A => S7399,
        B => S7407,
        Y => S7756
    );
NAND_4465: ENTITY WORK.NAND
    PORT MAP (
        A => S7400,
        B => S7408,
        Y => S7757
    );
NOR_2852: ENTITY WORK.NOR
    PORT MAP (
        A => S7755,
        B => S7757,
        Y => S7758
    );
NAND_4466: ENTITY WORK.NAND
    PORT MAP (
        A => S7754,
        B => S7756,
        Y => S7759
    );
NOR_2853: ENTITY WORK.NOR
    PORT MAP (
        A => S7754,
        B => S7756,
        Y => S7760
    );
NAND_4467: ENTITY WORK.NAND
    PORT MAP (
        A => S7755,
        B => S7757,
        Y => S7762
    );
NOR_2854: ENTITY WORK.NOR
    PORT MAP (
        A => S7758,
        B => S7760,
        Y => S7763
    );
NAND_4468: ENTITY WORK.NAND
    PORT MAP (
        A => S7759,
        B => S7762,
        Y => S7764
    );
NOR_2855: ENTITY WORK.NOR
    PORT MAP (
        A => S7743,
        B => S7764,
        Y => S7765
    );
NAND_4469: ENTITY WORK.NAND
    PORT MAP (
        A => S7744,
        B => S7763,
        Y => S7766
    );
NOR_2856: ENTITY WORK.NOR
    PORT MAP (
        A => S7744,
        B => S7763,
        Y => S7767
    );
NAND_4470: ENTITY WORK.NAND
    PORT MAP (
        A => S7743,
        B => S7764,
        Y => S7768
    );
NOR_2857: ENTITY WORK.NOR
    PORT MAP (
        A => S7765,
        B => S7767,
        Y => S7769
    );
NAND_4471: ENTITY WORK.NAND
    PORT MAP (
        A => S7766,
        B => S7768,
        Y => S7770
    );
NOR_2858: ENTITY WORK.NOR
    PORT MAP (
        A => S7413,
        B => S7421,
        Y => S7771
    );
NAND_4472: ENTITY WORK.NAND
    PORT MAP (
        A => S7414,
        B => S7422,
        Y => S7773
    );
NOR_2859: ENTITY WORK.NOR
    PORT MAP (
        A => S7770,
        B => S7773,
        Y => S7774
    );
NAND_4473: ENTITY WORK.NAND
    PORT MAP (
        A => S7769,
        B => S7771,
        Y => S7775
    );
NOR_2860: ENTITY WORK.NOR
    PORT MAP (
        A => S7769,
        B => S7771,
        Y => S7776
    );
NAND_4474: ENTITY WORK.NAND
    PORT MAP (
        A => S7770,
        B => S7773,
        Y => S7777
    );
NOR_2861: ENTITY WORK.NOR
    PORT MAP (
        A => S7774,
        B => S7776,
        Y => S7778
    );
NAND_4475: ENTITY WORK.NAND
    PORT MAP (
        A => S7775,
        B => S7777,
        Y => S7779
    );
NOR_2862: ENTITY WORK.NOR
    PORT MAP (
        A => S7741,
        B => S7778,
        Y => S7780
    );
NAND_4476: ENTITY WORK.NAND
    PORT MAP (
        A => S7742,
        B => S7779,
        Y => S7781
    );
NOR_2863: ENTITY WORK.NOR
    PORT MAP (
        A => S7742,
        B => S7779,
        Y => S7782
    );
NAND_4477: ENTITY WORK.NAND
    PORT MAP (
        A => S7741,
        B => S7778,
        Y => S7784
    );
NOR_2864: ENTITY WORK.NOR
    PORT MAP (
        A => S7780,
        B => S7782,
        Y => S7785
    );
NAND_4478: ENTITY WORK.NAND
    PORT MAP (
        A => S7781,
        B => S7784,
        Y => S7786
    );
NOR_2865: ENTITY WORK.NOR
    PORT MAP (
        A => S7738,
        B => S7785,
        Y => S7787
    );
NAND_4479: ENTITY WORK.NAND
    PORT MAP (
        A => S7740,
        B => S7786,
        Y => S7788
    );
NOR_2866: ENTITY WORK.NOR
    PORT MAP (
        A => S7740,
        B => S7786,
        Y => S7789
    );
NAND_4480: ENTITY WORK.NAND
    PORT MAP (
        A => S7738,
        B => S7785,
        Y => S7790
    );
NOR_2867: ENTITY WORK.NOR
    PORT MAP (
        A => S7787,
        B => S7789,
        Y => S7791
    );
NAND_4481: ENTITY WORK.NAND
    PORT MAP (
        A => S7788,
        B => S7790,
        Y => S7792
    );
NOR_2868: ENTITY WORK.NOR
    PORT MAP (
        A => S7571,
        B => S7792,
        Y => S7793
    );
NAND_4482: ENTITY WORK.NAND
    PORT MAP (
        A => S7572,
        B => S7791,
        Y => S7795
    );
NOR_2869: ENTITY WORK.NOR
    PORT MAP (
        A => S7572,
        B => S7791,
        Y => S7796
    );
NAND_4483: ENTITY WORK.NAND
    PORT MAP (
        A => S7571,
        B => S7792,
        Y => S7797
    );
NOR_2870: ENTITY WORK.NOR
    PORT MAP (
        A => S7793,
        B => S7796,
        Y => S7798
    );
NAND_4484: ENTITY WORK.NAND
    PORT MAP (
        A => S7795,
        B => S7797,
        Y => S7799
    );
NAND_4485: ENTITY WORK.NAND
    PORT MAP (
        A => S7353,
        B => S7554,
        Y => S7800
    );
NOT_539: ENTITY WORK.NOT
    PORT MAP (
        A => S7800,
        Y => S7801
    );
NOR_2871: ENTITY WORK.NOR
    PORT MAP (
        A => S7353,
        B => S7554,
        Y => S7802
    );
NOT_540: ENTITY WORK.NOT
    PORT MAP (
        A => S7802,
        Y => S7803
    );
NOR_2872: ENTITY WORK.NOR
    PORT MAP (
        A => S7801,
        B => S7802,
        Y => S7804
    );
NAND_4486: ENTITY WORK.NAND
    PORT MAP (
        A => S7800,
        B => S7803,
        Y => S7806
    );
NAND_4487: ENTITY WORK.NAND
    PORT MAP (
        A => S7798,
        B => S7806,
        Y => S7807
    );
NAND_4488: ENTITY WORK.NAND
    PORT MAP (
        A => S7799,
        B => S7804,
        Y => S7808
    );
NAND_4489: ENTITY WORK.NAND
    PORT MAP (
        A => S7807,
        B => S7808,
        Y => S7809
    );
NOR_2873: ENTITY WORK.NOR
    PORT MAP (
        A => S7570,
        B => S7809,
        Y => S7810
    );
NAND_4490: ENTITY WORK.NAND
    PORT MAP (
        A => S7570,
        B => S7809,
        Y => S7811
    );
NOR_2874: ENTITY WORK.NOR
    PORT MAP (
        A => S5949,
        B => S7810,
        Y => S7812
    );
NAND_4491: ENTITY WORK.NAND
    PORT MAP (
        A => S7811,
        B => S7812,
        Y => S7813
    );
NAND_4492: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_multdivunit_outmdu1_15,
        B => S5950,
        Y => S7814
    );
NOT_541: ENTITY WORK.NOT
    PORT MAP (
        A => S7814,
        Y => S7815
    );
NOR_2875: ENTITY WORK.NOR
    PORT MAP (
        A => datapath_addsubunit_in1_15,
        B => S1516,
        Y => S7817
    );
NOR_2876: ENTITY WORK.NOR
    PORT MAP (
        A => S3899,
        B => S7817,
        Y => S7818
    );
NOT_542: ENTITY WORK.NOT
    PORT MAP (
        A => S7818,
        Y => S7819
    );
NOR_2877: ENTITY WORK.NOR
    PORT MAP (
        A => S3927,
        B => S7819,
        Y => S7820
    );
NOR_2878: ENTITY WORK.NOR
    PORT MAP (
        A => S7815,
        B => S7820,
        Y => S7821
    );
NAND_4493: ENTITY WORK.NAND
    PORT MAP (
        A => S7813,
        B => S7821,
        Y => S297
    );
NOR_2879: ENTITY WORK.NOR
    PORT MAP (
        A => S8033,
        B => S1377,
        Y => S298
    );
NOR_2880: ENTITY WORK.NOR
    PORT MAP (
        A => S8044,
        B => S1377,
        Y => S299
    );
NOR_2881: ENTITY WORK.NOR
    PORT MAP (
        A => S8054,
        B => S1377,
        Y => S300
    );
NOR_2882: ENTITY WORK.NOR
    PORT MAP (
        A => S8065,
        B => S1377,
        Y => S301
    );
NOR_2883: ENTITY WORK.NOR
    PORT MAP (
        A => S8076,
        B => S1377,
        Y => S302
    );
NOR_2884: ENTITY WORK.NOR
    PORT MAP (
        A => S8087,
        B => S1377,
        Y => S303
    );
NOR_2885: ENTITY WORK.NOR
    PORT MAP (
        A => S8097,
        B => S1377,
        Y => S304
    );
NOR_2886: ENTITY WORK.NOR
    PORT MAP (
        A => S8108,
        B => S1377,
        Y => S305
    );
NOR_2887: ENTITY WORK.NOR
    PORT MAP (
        A => S8119,
        B => S1377,
        Y => S306
    );
NOR_2888: ENTITY WORK.NOR
    PORT MAP (
        A => S8129,
        B => S1377,
        Y => S307
    );
NOR_2889: ENTITY WORK.NOR
    PORT MAP (
        A => S8140,
        B => S1377,
        Y => S308
    );
NOR_2890: ENTITY WORK.NOR
    PORT MAP (
        A => S8151,
        B => S1377,
        Y => S309
    );
NOR_2891: ENTITY WORK.NOR
    PORT MAP (
        A => S8161,
        B => S1377,
        Y => S310
    );
NOR_2892: ENTITY WORK.NOR
    PORT MAP (
        A => S8172,
        B => S1377,
        Y => S311
    );
NOR_2893: ENTITY WORK.NOR
    PORT MAP (
        A => S8183,
        B => S1377,
        Y => S312
    );
NAND_4494: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_databusin_0,
        B => controller_1115_S_0,
        Y => S7824
    );
NAND_4495: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_instruction_0,
        B => S1379,
        Y => S7825
    );
NAND_4496: ENTITY WORK.NAND
    PORT MAP (
        A => S7824,
        B => S7825,
        Y => S313
    );
NAND_4497: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_databusin_1,
        B => controller_1115_S_0,
        Y => S7826
    );
NAND_4498: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_instruction_1,
        B => S1379,
        Y => S7827
    );
NAND_4499: ENTITY WORK.NAND
    PORT MAP (
        A => S7826,
        B => S7827,
        Y => S314
    );
NAND_4500: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_databusin_2,
        B => controller_1115_S_0,
        Y => S7828
    );
NAND_4501: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_instruction_2,
        B => S1379,
        Y => S7829
    );
NAND_4502: ENTITY WORK.NAND
    PORT MAP (
        A => S7828,
        B => S7829,
        Y => S315
    );
NAND_4503: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_databusin_3,
        B => controller_1115_S_0,
        Y => S7831
    );
NAND_4504: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_instruction_3,
        B => S1379,
        Y => S7832
    );
NAND_4505: ENTITY WORK.NAND
    PORT MAP (
        A => S7831,
        B => S7832,
        Y => S316
    );
NAND_4506: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_databusin_4,
        B => controller_1115_S_0,
        Y => S7833
    );
NAND_4507: ENTITY WORK.NAND
    PORT MAP (
        A => controller_fib_0,
        B => S1379,
        Y => S7834
    );
NAND_4508: ENTITY WORK.NAND
    PORT MAP (
        A => S7833,
        B => S7834,
        Y => S317
    );
NAND_4509: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_databusin_5,
        B => controller_1115_S_0,
        Y => S7835
    );
NAND_4510: ENTITY WORK.NAND
    PORT MAP (
        A => controller_fib_1,
        B => S1379,
        Y => S7836
    );
NAND_4511: ENTITY WORK.NAND
    PORT MAP (
        A => S7835,
        B => S7836,
        Y => S318
    );
NAND_4512: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_databusin_6,
        B => controller_1115_S_0,
        Y => S7837
    );
NAND_4513: ENTITY WORK.NAND
    PORT MAP (
        A => controller_fib_2,
        B => S1379,
        Y => S7839
    );
NAND_4514: ENTITY WORK.NAND
    PORT MAP (
        A => S7837,
        B => S7839,
        Y => S319
    );
NAND_4515: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_databusin_7,
        B => controller_1115_S_0,
        Y => S7840
    );
NAND_4516: ENTITY WORK.NAND
    PORT MAP (
        A => controller_fib_3,
        B => S1379,
        Y => S7841
    );
NAND_4517: ENTITY WORK.NAND
    PORT MAP (
        A => S7840,
        B => S7841,
        Y => S320
    );
NAND_4518: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_databusin_8,
        B => controller_1115_S_0,
        Y => S7842
    );
NAND_4519: ENTITY WORK.NAND
    PORT MAP (
        A => controller_fib_4,
        B => S1379,
        Y => S7843
    );
NAND_4520: ENTITY WORK.NAND
    PORT MAP (
        A => S7842,
        B => S7843,
        Y => S321
    );
NAND_4521: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_databusin_9,
        B => controller_1115_S_0,
        Y => S7844
    );
NAND_4522: ENTITY WORK.NAND
    PORT MAP (
        A => controller_216_B_0,
        B => S1379,
        Y => S7845
    );
NAND_4523: ENTITY WORK.NAND
    PORT MAP (
        A => S7844,
        B => S7845,
        Y => S322
    );
NAND_4524: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_databusin_10,
        B => controller_1115_S_0,
        Y => S7847
    );
NAND_4525: ENTITY WORK.NAND
    PORT MAP (
        A => controller_opcode_2,
        B => S1379,
        Y => S7848
    );
NAND_4526: ENTITY WORK.NAND
    PORT MAP (
        A => S7847,
        B => S7848,
        Y => S323
    );
NAND_4527: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_databusin_11,
        B => controller_1115_S_0,
        Y => S7849
    );
NAND_4528: ENTITY WORK.NAND
    PORT MAP (
        A => controller_opcode_3,
        B => S1379,
        Y => S7850
    );
NAND_4529: ENTITY WORK.NAND
    PORT MAP (
        A => S7849,
        B => S7850,
        Y => S324
    );
NAND_4530: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_databusin_12,
        B => controller_1115_S_0,
        Y => S7851
    );
NAND_4531: ENTITY WORK.NAND
    PORT MAP (
        A => controller_opcode_4,
        B => S1379,
        Y => S7852
    );
NAND_4532: ENTITY WORK.NAND
    PORT MAP (
        A => S7851,
        B => S7852,
        Y => S325
    );
NAND_4533: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_databusin_13,
        B => controller_1115_S_0,
        Y => S7854
    );
NAND_4534: ENTITY WORK.NAND
    PORT MAP (
        A => controller_opcode_5,
        B => S1379,
        Y => S7855
    );
NAND_4535: ENTITY WORK.NAND
    PORT MAP (
        A => S7854,
        B => S7855,
        Y => S326
    );
NAND_4536: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_databusin_14,
        B => controller_1115_S_0,
        Y => S7856
    );
NAND_4537: ENTITY WORK.NAND
    PORT MAP (
        A => controller_opcode_6,
        B => S1379,
        Y => S7857
    );
NAND_4538: ENTITY WORK.NAND
    PORT MAP (
        A => S7856,
        B => S7857,
        Y => S327
    );
NAND_4539: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_adr_outreg_0,
        B => S1383,
        Y => S7858
    );
NAND_4540: ENTITY WORK.NAND
    PORT MAP (
        A => S1222,
        B => S1382,
        Y => S7859
    );
NAND_4541: ENTITY WORK.NAND
    PORT MAP (
        A => S7858,
        B => S7859,
        Y => S328
    );
NAND_4542: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_adr_outreg_1,
        B => S1383,
        Y => S7860
    );
NAND_4543: ENTITY WORK.NAND
    PORT MAP (
        A => S1170,
        B => S1382,
        Y => S7862
    );
NAND_4544: ENTITY WORK.NAND
    PORT MAP (
        A => S7860,
        B => S7862,
        Y => S329
    );
NAND_4545: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_adr_outreg_2,
        B => S1383,
        Y => S7863
    );
NAND_4546: ENTITY WORK.NAND
    PORT MAP (
        A => S1118,
        B => S1382,
        Y => S7864
    );
NAND_4547: ENTITY WORK.NAND
    PORT MAP (
        A => S7863,
        B => S7864,
        Y => S330
    );
NAND_4548: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_adr_outreg_3,
        B => S1383,
        Y => S7865
    );
NAND_4549: ENTITY WORK.NAND
    PORT MAP (
        A => S1067,
        B => S1382,
        Y => S7866
    );
NAND_4550: ENTITY WORK.NAND
    PORT MAP (
        A => S7865,
        B => S7866,
        Y => S331
    );
NAND_4551: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_adr_outreg_4,
        B => S1383,
        Y => S7867
    );
NAND_4552: ENTITY WORK.NAND
    PORT MAP (
        A => S1015,
        B => S1382,
        Y => S7868
    );
NAND_4553: ENTITY WORK.NAND
    PORT MAP (
        A => S7867,
        B => S7868,
        Y => S332
    );
NAND_4554: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_adr_outreg_5,
        B => S1383,
        Y => S7870
    );
NAND_4555: ENTITY WORK.NAND
    PORT MAP (
        A => S965,
        B => S1382,
        Y => S7871
    );
NAND_4556: ENTITY WORK.NAND
    PORT MAP (
        A => S7870,
        B => S7871,
        Y => S333
    );
NAND_4557: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_adr_outreg_6,
        B => S1383,
        Y => S7872
    );
NAND_4558: ENTITY WORK.NAND
    PORT MAP (
        A => S912,
        B => S1382,
        Y => S7873
    );
NAND_4559: ENTITY WORK.NAND
    PORT MAP (
        A => S7872,
        B => S7873,
        Y => S334
    );
NAND_4560: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_adr_outreg_7,
        B => S1383,
        Y => S7874
    );
NAND_4561: ENTITY WORK.NAND
    PORT MAP (
        A => S860,
        B => S1382,
        Y => S7875
    );
NAND_4562: ENTITY WORK.NAND
    PORT MAP (
        A => S7874,
        B => S7875,
        Y => S335
    );
NAND_4563: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_adr_outreg_8,
        B => S1383,
        Y => S7877
    );
NAND_4564: ENTITY WORK.NAND
    PORT MAP (
        A => S807,
        B => S1382,
        Y => S7878
    );
NAND_4565: ENTITY WORK.NAND
    PORT MAP (
        A => S7877,
        B => S7878,
        Y => S336
    );
NAND_4566: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_adr_outreg_9,
        B => S1383,
        Y => S7879
    );
NAND_4567: ENTITY WORK.NAND
    PORT MAP (
        A => S756,
        B => S1382,
        Y => S7880
    );
NAND_4568: ENTITY WORK.NAND
    PORT MAP (
        A => S7879,
        B => S7880,
        Y => S337
    );
NAND_4569: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_adr_outreg_10,
        B => S1383,
        Y => S7881
    );
NAND_4570: ENTITY WORK.NAND
    PORT MAP (
        A => S704,
        B => S1382,
        Y => S7882
    );
NAND_4571: ENTITY WORK.NAND
    PORT MAP (
        A => S7881,
        B => S7882,
        Y => S338
    );
NAND_4572: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_adr_outreg_11,
        B => S1383,
        Y => S7883
    );
NAND_4573: ENTITY WORK.NAND
    PORT MAP (
        A => S653,
        B => S1382,
        Y => S7885
    );
NAND_4574: ENTITY WORK.NAND
    PORT MAP (
        A => S7883,
        B => S7885,
        Y => S339
    );
NAND_4575: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_adr_outreg_12,
        B => S1383,
        Y => S7886
    );
NAND_4576: ENTITY WORK.NAND
    PORT MAP (
        A => S601,
        B => S1382,
        Y => S7887
    );
NAND_4577: ENTITY WORK.NAND
    PORT MAP (
        A => S7886,
        B => S7887,
        Y => S340
    );
NAND_4578: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_adr_outreg_13,
        B => S1383,
        Y => S7888
    );
NAND_4579: ENTITY WORK.NAND
    PORT MAP (
        A => S550,
        B => S1382,
        Y => S7889
    );
NAND_4580: ENTITY WORK.NAND
    PORT MAP (
        A => S7888,
        B => S7889,
        Y => S341
    );
NAND_4581: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_adr_outreg_14,
        B => S1383,
        Y => S7890
    );
NAND_4582: ENTITY WORK.NAND
    PORT MAP (
        A => S498,
        B => S1382,
        Y => S7891
    );
NAND_4583: ENTITY WORK.NAND
    PORT MAP (
        A => S7890,
        B => S7891,
        Y => S342
    );
NOR_2894: ENTITY WORK.NOR
    PORT MAP (
        A => controller_216_B_0,
        B => S1628,
        Y => controller_readmem
    );
NOR_2895: ENTITY WORK.NOR
    PORT MAP (
        A => controller_216_B_0,
        B => S403,
        Y => controller_writemem
    );
NAND_4584: ENTITY WORK.NAND
    PORT MAP (
        A => controller_216_B_0,
        B => S1627,
        Y => S7893
    );
NOT_543: ENTITY WORK.NOT
    PORT MAP (
        A => S7893,
        Y => controller_readio
    );
NOR_2896: ENTITY WORK.NOR
    PORT MAP (
        A => S8278,
        B => S403,
        Y => controller_writeio
    );
NOR_2897: ENTITY WORK.NOR
    PORT MAP (
        A => S1377,
        B => controller_1115_S_0,
        Y => S7894
    );
NOT_544: ENTITY WORK.NOT
    PORT MAP (
        A => S7894,
        Y => controller_1405_Y_0
    );
NAND_4585: ENTITY WORK.NAND
    PORT MAP (
        A => S8572,
        B => S8576,
        Y => S7895
    );
NOT_545: ENTITY WORK.NOT
    PORT MAP (
        A => S7895,
        Y => S7896
    );
NAND_4586: ENTITY WORK.NAND
    PORT MAP (
        A => S1383,
        B => S5950,
        Y => S7898
    );
NOR_2898: ENTITY WORK.NOR
    PORT MAP (
        A => S7896,
        B => S7898,
        Y => S7899
    );
NAND_4587: ENTITY WORK.NAND
    PORT MAP (
        A => S1378,
        B => S7899,
        Y => controller_1405_Y_1
    );
NAND_4588: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_0,
        B => controller_1115_S_0,
        Y => S7900
    );
NAND_4589: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_adr_outreg_0,
        B => S8576,
        Y => S7901
    );
NAND_4590: ENTITY WORK.NAND
    PORT MAP (
        A => S7900,
        B => S7901,
        Y => datapath_addrbus_0
    );
NAND_4591: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_1,
        B => controller_1115_S_0,
        Y => S7902
    );
NAND_4592: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_adr_outreg_1,
        B => S8576,
        Y => S7903
    );
NAND_4593: ENTITY WORK.NAND
    PORT MAP (
        A => S7902,
        B => S7903,
        Y => datapath_addrbus_1
    );
NAND_4594: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_2,
        B => controller_1115_S_0,
        Y => S7904
    );
NAND_4595: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_adr_outreg_2,
        B => S8576,
        Y => S7906
    );
NAND_4596: ENTITY WORK.NAND
    PORT MAP (
        A => S7904,
        B => S7906,
        Y => datapath_addrbus_2
    );
NAND_4597: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_3,
        B => controller_1115_S_0,
        Y => S7907
    );
NAND_4598: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_adr_outreg_3,
        B => S8576,
        Y => S7908
    );
NAND_4599: ENTITY WORK.NAND
    PORT MAP (
        A => S7907,
        B => S7908,
        Y => datapath_addrbus_3
    );
NAND_4600: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_4,
        B => controller_1115_S_0,
        Y => S7909
    );
NAND_4601: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_adr_outreg_4,
        B => S8576,
        Y => S7910
    );
NAND_4602: ENTITY WORK.NAND
    PORT MAP (
        A => S7909,
        B => S7910,
        Y => datapath_addrbus_4
    );
NAND_4603: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_5,
        B => controller_1115_S_0,
        Y => S7911
    );
NAND_4604: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_adr_outreg_5,
        B => S8576,
        Y => S7912
    );
NAND_4605: ENTITY WORK.NAND
    PORT MAP (
        A => S7911,
        B => S7912,
        Y => datapath_addrbus_5
    );
NAND_4606: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_6,
        B => controller_1115_S_0,
        Y => S7914
    );
NAND_4607: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_adr_outreg_6,
        B => S8576,
        Y => S7915
    );
NAND_4608: ENTITY WORK.NAND
    PORT MAP (
        A => S7914,
        B => S7915,
        Y => datapath_addrbus_6
    );
NAND_4609: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_7,
        B => controller_1115_S_0,
        Y => S7916
    );
NAND_4610: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_adr_outreg_7,
        B => S8576,
        Y => S7917
    );
NAND_4611: ENTITY WORK.NAND
    PORT MAP (
        A => S7916,
        B => S7917,
        Y => datapath_addrbus_7
    );
NAND_4612: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_8,
        B => controller_1115_S_0,
        Y => S7918
    );
NAND_4613: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_adr_outreg_8,
        B => S8576,
        Y => S7919
    );
NAND_4614: ENTITY WORK.NAND
    PORT MAP (
        A => S7918,
        B => S7919,
        Y => datapath_addrbus_8
    );
NAND_4615: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_9,
        B => controller_1115_S_0,
        Y => S7921
    );
NAND_4616: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_adr_outreg_9,
        B => S8576,
        Y => S7922
    );
NAND_4617: ENTITY WORK.NAND
    PORT MAP (
        A => S7921,
        B => S7922,
        Y => datapath_addrbus_9
    );
NAND_4618: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_10,
        B => controller_1115_S_0,
        Y => S7923
    );
NAND_4619: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_adr_outreg_10,
        B => S8576,
        Y => S7924
    );
NAND_4620: ENTITY WORK.NAND
    PORT MAP (
        A => S7923,
        B => S7924,
        Y => datapath_addrbus_10
    );
NAND_4621: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_11,
        B => controller_1115_S_0,
        Y => S7925
    );
NAND_4622: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_adr_outreg_11,
        B => S8576,
        Y => S7926
    );
NAND_4623: ENTITY WORK.NAND
    PORT MAP (
        A => S7925,
        B => S7926,
        Y => datapath_addrbus_11
    );
NAND_4624: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_12,
        B => controller_1115_S_0,
        Y => S7927
    );
NAND_4625: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_adr_outreg_12,
        B => S8576,
        Y => S7929
    );
NAND_4626: ENTITY WORK.NAND
    PORT MAP (
        A => S7927,
        B => S7929,
        Y => datapath_addrbus_12
    );
NAND_4627: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_13,
        B => controller_1115_S_0,
        Y => S7930
    );
NAND_4628: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_adr_outreg_13,
        B => S8576,
        Y => S7931
    );
NAND_4629: ENTITY WORK.NAND
    PORT MAP (
        A => S7930,
        B => S7931,
        Y => datapath_addrbus_13
    );
NAND_4630: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_14,
        B => controller_1115_S_0,
        Y => S7932
    );
NAND_4631: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_adr_outreg_14,
        B => S8576,
        Y => S7933
    );
NAND_4632: ENTITY WORK.NAND
    PORT MAP (
        A => S7932,
        B => S7933,
        Y => datapath_addrbus_14
    );
NAND_4633: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_muxmem_in2_15,
        B => controller_1115_S_0,
        Y => S7934
    );
NAND_4634: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_adr_outreg_15,
        B => S8576,
        Y => S7935
    );
NAND_4635: ENTITY WORK.NAND
    PORT MAP (
        A => S7934,
        B => S7935,
        Y => datapath_addrbus_15
    );
NOR_2899: ENTITY WORK.NOR
    PORT MAP (
        A => S1604,
        B => S1746,
        Y => S7937
    );
NAND_4636: ENTITY WORK.NAND
    PORT MAP (
        A => S1605,
        B => S1745,
        Y => S7938
    );
NAND_4637: ENTITY WORK.NAND
    PORT MAP (
        A => controller_fib_1,
        B => S1607,
        Y => S7939
    );
NOT_546: ENTITY WORK.NOT
    PORT MAP (
        A => S7939,
        Y => S7940
    );
NOR_2900: ENTITY WORK.NOR
    PORT MAP (
        A => S7937,
        B => S7940,
        Y => S7941
    );
NAND_4638: ENTITY WORK.NAND
    PORT MAP (
        A => S7938,
        B => S7939,
        Y => S7942
    );
NOR_2901: ENTITY WORK.NOR
    PORT MAP (
        A => S1516,
        B => S1604,
        Y => S7943
    );
NAND_4639: ENTITY WORK.NAND
    PORT MAP (
        A => S1515,
        B => S1605,
        Y => S7944
    );
NAND_4640: ENTITY WORK.NAND
    PORT MAP (
        A => controller_fib_0,
        B => S1607,
        Y => S7945
    );
NOT_547: ENTITY WORK.NOT
    PORT MAP (
        A => S7945,
        Y => S7947
    );
NOR_2902: ENTITY WORK.NOR
    PORT MAP (
        A => S7943,
        B => S7947,
        Y => S7948
    );
NAND_4641: ENTITY WORK.NAND
    PORT MAP (
        A => S7944,
        B => S7945,
        Y => S7949
    );
NOR_2903: ENTITY WORK.NOR
    PORT MAP (
        A => S7942,
        B => S7949,
        Y => S7950
    );
NAND_4642: ENTITY WORK.NAND
    PORT MAP (
        A => S7941,
        B => S7948,
        Y => S7951
    );
NOR_2904: ENTITY WORK.NOR
    PORT MAP (
        A => S1604,
        B => S1953,
        Y => S7952
    );
NAND_4643: ENTITY WORK.NAND
    PORT MAP (
        A => S1605,
        B => S1952,
        Y => S7953
    );
NAND_4644: ENTITY WORK.NAND
    PORT MAP (
        A => controller_fib_3,
        B => S1607,
        Y => S7954
    );
NOT_548: ENTITY WORK.NOT
    PORT MAP (
        A => S7954,
        Y => S7955
    );
NOR_2905: ENTITY WORK.NOR
    PORT MAP (
        A => S7952,
        B => S7955,
        Y => S7956
    );
NAND_4645: ENTITY WORK.NAND
    PORT MAP (
        A => S7953,
        B => S7954,
        Y => S7958
    );
NOR_2906: ENTITY WORK.NOR
    PORT MAP (
        A => S1604,
        B => S1849,
        Y => S7959
    );
NAND_4646: ENTITY WORK.NAND
    PORT MAP (
        A => S1605,
        B => S1848,
        Y => S7960
    );
NAND_4647: ENTITY WORK.NAND
    PORT MAP (
        A => controller_fib_2,
        B => S1607,
        Y => S7961
    );
NOT_549: ENTITY WORK.NOT
    PORT MAP (
        A => S7961,
        Y => S7962
    );
NOR_2907: ENTITY WORK.NOR
    PORT MAP (
        A => S7959,
        B => S7962,
        Y => S7963
    );
NAND_4648: ENTITY WORK.NAND
    PORT MAP (
        A => S7960,
        B => S7961,
        Y => S7964
    );
NOR_2908: ENTITY WORK.NOR
    PORT MAP (
        A => S7958,
        B => S7964,
        Y => S7965
    );
NAND_4649: ENTITY WORK.NAND
    PORT MAP (
        A => S7956,
        B => S7963,
        Y => S7966
    );
NOR_2909: ENTITY WORK.NOR
    PORT MAP (
        A => S7951,
        B => S7966,
        Y => S7967
    );
NAND_4650: ENTITY WORK.NAND
    PORT MAP (
        A => S7950,
        B => S7965,
        Y => S7969
    );
NAND_4651: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_0,
        B => S7967,
        Y => S7970
    );
NOT_550: ENTITY WORK.NOT
    PORT MAP (
        A => S7970,
        Y => datapath_shiftunit_2439_A
    );
NOR_2910: ENTITY WORK.NOR
    PORT MAP (
        A => S7941,
        B => S7948,
        Y => S7971
    );
NAND_4652: ENTITY WORK.NAND
    PORT MAP (
        A => S7942,
        B => S7949,
        Y => S7972
    );
NOR_2911: ENTITY WORK.NOR
    PORT MAP (
        A => S7966,
        B => S7972,
        Y => S7973
    );
NAND_4653: ENTITY WORK.NAND
    PORT MAP (
        A => S7965,
        B => S7971,
        Y => S7974
    );
NAND_4654: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_3,
        B => S7973,
        Y => S7975
    );
NOR_2912: ENTITY WORK.NOR
    PORT MAP (
        A => S7956,
        B => S7964,
        Y => S7976
    );
NAND_4655: ENTITY WORK.NAND
    PORT MAP (
        A => S7958,
        B => S7963,
        Y => S7977
    );
NOR_2913: ENTITY WORK.NOR
    PORT MAP (
        A => S7941,
        B => S7949,
        Y => S7979
    );
NAND_4656: ENTITY WORK.NAND
    PORT MAP (
        A => S7942,
        B => S7948,
        Y => S7980
    );
NAND_4657: ENTITY WORK.NAND
    PORT MAP (
        A => S7976,
        B => S7979,
        Y => S7981
    );
NOT_551: ENTITY WORK.NOT
    PORT MAP (
        A => S7981,
        Y => S7982
    );
NAND_4658: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_10,
        B => S7982,
        Y => S7983
    );
NOR_2914: ENTITY WORK.NOR
    PORT MAP (
        A => S7951,
        B => S7977,
        Y => S7984
    );
NAND_4659: ENTITY WORK.NAND
    PORT MAP (
        A => S7950,
        B => S7976,
        Y => S7985
    );
NAND_4660: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_8,
        B => S7984,
        Y => S7986
    );
NOR_2915: ENTITY WORK.NOR
    PORT MAP (
        A => S7942,
        B => S7948,
        Y => S7987
    );
NAND_4661: ENTITY WORK.NAND
    PORT MAP (
        A => S7941,
        B => S7949,
        Y => S7988
    );
NOR_2916: ENTITY WORK.NOR
    PORT MAP (
        A => S7956,
        B => S7963,
        Y => S7990
    );
NAND_4662: ENTITY WORK.NAND
    PORT MAP (
        A => S7958,
        B => S7964,
        Y => S7991
    );
NAND_4663: ENTITY WORK.NAND
    PORT MAP (
        A => S7987,
        B => S7990,
        Y => S7992
    );
NOT_552: ENTITY WORK.NOT
    PORT MAP (
        A => S7992,
        Y => S7993
    );
NAND_4664: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_13,
        B => S7993,
        Y => S7994
    );
NOR_2917: ENTITY WORK.NOR
    PORT MAP (
        A => S7951,
        B => S7991,
        Y => S7995
    );
NAND_4665: ENTITY WORK.NAND
    PORT MAP (
        A => S7950,
        B => S7990,
        Y => S7996
    );
NAND_4666: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_12,
        B => S7995,
        Y => S7997
    );
NAND_4667: ENTITY WORK.NAND
    PORT MAP (
        A => S7994,
        B => S7997,
        Y => S7998
    );
NOR_2918: ENTITY WORK.NOR
    PORT MAP (
        A => S7958,
        B => S7963,
        Y => S7999
    );
NAND_4668: ENTITY WORK.NAND
    PORT MAP (
        A => S7956,
        B => S7964,
        Y => S8001
    );
NOR_2919: ENTITY WORK.NOR
    PORT MAP (
        A => S7951,
        B => S8001,
        Y => S8002
    );
NAND_4669: ENTITY WORK.NAND
    PORT MAP (
        A => S7950,
        B => S7999,
        Y => S8003
    );
NOR_2920: ENTITY WORK.NOR
    PORT MAP (
        A => S1013,
        B => S8003,
        Y => S8004
    );
NAND_4670: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_4,
        B => S8002,
        Y => S8005
    );
NOR_2921: ENTITY WORK.NOR
    PORT MAP (
        A => S7972,
        B => S7977,
        Y => S8006
    );
NAND_4671: ENTITY WORK.NAND
    PORT MAP (
        A => S7971,
        B => S7976,
        Y => S8007
    );
NAND_4672: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_11,
        B => S8006,
        Y => S8008
    );
NOR_2922: ENTITY WORK.NOR
    PORT MAP (
        A => S7966,
        B => S7988,
        Y => S8009
    );
NAND_4673: ENTITY WORK.NAND
    PORT MAP (
        A => S7965,
        B => S7987,
        Y => S8010
    );
NOR_2923: ENTITY WORK.NOR
    PORT MAP (
        A => S1168,
        B => S8010,
        Y => S8012
    );
NAND_4674: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_1,
        B => S8009,
        Y => S8013
    );
NOR_2924: ENTITY WORK.NOR
    PORT MAP (
        A => S7966,
        B => S7980,
        Y => S8014
    );
NAND_4675: ENTITY WORK.NAND
    PORT MAP (
        A => S7965,
        B => S7979,
        Y => S8015
    );
NAND_4676: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_2,
        B => S8014,
        Y => S8016
    );
NOR_2925: ENTITY WORK.NOR
    PORT MAP (
        A => S7980,
        B => S8001,
        Y => S8017
    );
NAND_4677: ENTITY WORK.NAND
    PORT MAP (
        A => S7979,
        B => S7999,
        Y => S8018
    );
NOR_2926: ENTITY WORK.NOR
    PORT MAP (
        A => S910,
        B => S8018,
        Y => S8019
    );
NOR_2927: ENTITY WORK.NOR
    PORT MAP (
        A => S7977,
        B => S7988,
        Y => S8020
    );
NAND_4678: ENTITY WORK.NAND
    PORT MAP (
        A => S7976,
        B => S7987,
        Y => S8021
    );
NAND_4679: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_9,
        B => S8020,
        Y => S8023
    );
NOR_2928: ENTITY WORK.NOR
    PORT MAP (
        A => S7988,
        B => S8001,
        Y => S8024
    );
NAND_4680: ENTITY WORK.NAND
    PORT MAP (
        A => S7987,
        B => S7999,
        Y => S8025
    );
NOR_2929: ENTITY WORK.NOR
    PORT MAP (
        A => S963,
        B => S8025,
        Y => S8026
    );
NOR_2930: ENTITY WORK.NOR
    PORT MAP (
        A => S7980,
        B => S7991,
        Y => S8027
    );
NAND_4681: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_14,
        B => S8027,
        Y => S8028
    );
NAND_4682: ENTITY WORK.NAND
    PORT MAP (
        A => S7964,
        B => S7971,
        Y => S8029
    );
NOR_2931: ENTITY WORK.NOR
    PORT MAP (
        A => S7972,
        B => S8001,
        Y => S8030
    );
NAND_4683: ENTITY WORK.NAND
    PORT MAP (
        A => S7971,
        B => S7999,
        Y => S8031
    );
NOR_2932: ENTITY WORK.NOR
    PORT MAP (
        A => S858,
        B => S8031,
        Y => S8032
    );
NAND_4684: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_7,
        B => S8030,
        Y => S8034
    );
NOR_2933: ENTITY WORK.NOR
    PORT MAP (
        A => S7956,
        B => S8029,
        Y => S8035
    );
NAND_4685: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_15,
        B => S8035,
        Y => S8036
    );
NOR_2934: ENTITY WORK.NOR
    PORT MAP (
        A => S8004,
        B => S8032,
        Y => S8037
    );
NAND_4686: ENTITY WORK.NAND
    PORT MAP (
        A => S7971,
        B => S7990,
        Y => S8038
    );
NAND_4687: ENTITY WORK.NAND
    PORT MAP (
        A => S7986,
        B => S8023,
        Y => S8039
    );
NAND_4688: ENTITY WORK.NAND
    PORT MAP (
        A => S7970,
        B => S8013,
        Y => S8040
    );
NAND_4689: ENTITY WORK.NAND
    PORT MAP (
        A => S7975,
        B => S8016,
        Y => S8041
    );
NOR_2935: ENTITY WORK.NOR
    PORT MAP (
        A => S8040,
        B => S8041,
        Y => S8042
    );
NAND_4690: ENTITY WORK.NAND
    PORT MAP (
        A => S7983,
        B => S8042,
        Y => S8043
    );
NOR_2936: ENTITY WORK.NOR
    PORT MAP (
        A => S7998,
        B => S8043,
        Y => S8045
    );
NOR_2937: ENTITY WORK.NOR
    PORT MAP (
        A => S8019,
        B => S8026,
        Y => S8046
    );
NAND_4691: ENTITY WORK.NAND
    PORT MAP (
        A => S8037,
        B => S8046,
        Y => S8047
    );
NAND_4692: ENTITY WORK.NAND
    PORT MAP (
        A => S8008,
        B => S8028,
        Y => S8048
    );
NOR_2938: ENTITY WORK.NOR
    PORT MAP (
        A => S8039,
        B => S8048,
        Y => S8049
    );
NAND_4693: ENTITY WORK.NAND
    PORT MAP (
        A => S8036,
        B => S8049,
        Y => S8050
    );
NOR_2939: ENTITY WORK.NOR
    PORT MAP (
        A => S8047,
        B => S8050,
        Y => S8051
    );
NAND_4694: ENTITY WORK.NAND
    PORT MAP (
        A => S8045,
        B => S8051,
        Y => datapath_shiftunit_2135_A
    );
NOR_2940: ENTITY WORK.NOR
    PORT MAP (
        A => S910,
        B => S8025,
        Y => S8052
    );
NAND_4695: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_6,
        B => S8024,
        Y => S8053
    );
NOR_2941: ENTITY WORK.NOR
    PORT MAP (
        A => S1116,
        B => S8010,
        Y => S8055
    );
NAND_4696: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_2,
        B => S8009,
        Y => S8056
    );
NOR_2942: ENTITY WORK.NOR
    PORT MAP (
        A => S548,
        B => S7996,
        Y => S8057
    );
NAND_4697: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_5,
        B => S8002,
        Y => S8058
    );
NAND_4698: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_9,
        B => S7984,
        Y => S8059
    );
NAND_4699: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_3,
        B => S8014,
        Y => S8060
    );
NOR_2943: ENTITY WORK.NOR
    PORT MAP (
        A => S858,
        B => S8018,
        Y => S8061
    );
NAND_4700: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_10,
        B => S8020,
        Y => S8062
    );
NOR_2944: ENTITY WORK.NOR
    PORT MAP (
        A => S1013,
        B => S7974,
        Y => S8063
    );
NAND_4701: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_4,
        B => S7973,
        Y => S8064
    );
NAND_4702: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_11,
        B => S7982,
        Y => S8066
    );
NAND_4703: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_1,
        B => S7967,
        Y => S8067
    );
NAND_4704: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_12,
        B => S8006,
        Y => S8068
    );
NAND_4705: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_14,
        B => S7993,
        Y => S8069
    );
NAND_4706: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_8,
        B => S8030,
        Y => S8070
    );
NAND_4707: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_15,
        B => S8027,
        Y => S8071
    );
NAND_4708: ENTITY WORK.NAND
    PORT MAP (
        A => S8062,
        B => S8070,
        Y => S8072
    );
NAND_4709: ENTITY WORK.NAND
    PORT MAP (
        A => S8056,
        B => S8069,
        Y => S8073
    );
NOR_2945: ENTITY WORK.NOR
    PORT MAP (
        A => S8072,
        B => S8073,
        Y => S8074
    );
NOR_2946: ENTITY WORK.NOR
    PORT MAP (
        A => S8052,
        B => S8057,
        Y => S8075
    );
NAND_4710: ENTITY WORK.NAND
    PORT MAP (
        A => S8058,
        B => S8059,
        Y => S8077
    );
NOR_2947: ENTITY WORK.NOR
    PORT MAP (
        A => S1304,
        B => S1612,
        Y => S8078
    );
NAND_4711: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_15,
        B => S1611,
        Y => S8079
    );
NOR_2948: ENTITY WORK.NOR
    PORT MAP (
        A => S8038,
        B => S8079,
        Y => S8080
    );
NOR_2949: ENTITY WORK.NOR
    PORT MAP (
        A => S8077,
        B => S8080,
        Y => S8081
    );
NAND_4712: ENTITY WORK.NAND
    PORT MAP (
        A => S8075,
        B => S8081,
        Y => S8082
    );
NAND_4713: ENTITY WORK.NAND
    PORT MAP (
        A => S8068,
        B => S8071,
        Y => S8083
    );
NOR_2950: ENTITY WORK.NOR
    PORT MAP (
        A => S8061,
        B => S8083,
        Y => S8084
    );
NAND_4714: ENTITY WORK.NAND
    PORT MAP (
        A => S8060,
        B => S8067,
        Y => S8085
    );
NAND_4715: ENTITY WORK.NAND
    PORT MAP (
        A => S8064,
        B => S8066,
        Y => S8086
    );
NOR_2951: ENTITY WORK.NOR
    PORT MAP (
        A => S8085,
        B => S8086,
        Y => S8088
    );
NAND_4716: ENTITY WORK.NAND
    PORT MAP (
        A => S8084,
        B => S8088,
        Y => S8089
    );
NOR_2952: ENTITY WORK.NOR
    PORT MAP (
        A => S8082,
        B => S8089,
        Y => S8090
    );
NAND_4717: ENTITY WORK.NAND
    PORT MAP (
        A => S8074,
        B => S8090,
        Y => datapath_shiftunit_2153_A
    );
NAND_4718: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_4,
        B => S8014,
        Y => S8091
    );
NAND_4719: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_5,
        B => S7973,
        Y => S8092
    );
NAND_4720: ENTITY WORK.NAND
    PORT MAP (
        A => S8091,
        B => S8092,
        Y => S8093
    );
NOR_2953: ENTITY WORK.NOR
    PORT MAP (
        A => S599,
        B => S7981,
        Y => S8094
    );
NOR_2954: ENTITY WORK.NOR
    PORT MAP (
        A => S1304,
        B => S7992,
        Y => S8095
    );
NOR_2955: ENTITY WORK.NOR
    PORT MAP (
        A => S8094,
        B => S8095,
        Y => S8096
    );
NOR_2956: ENTITY WORK.NOR
    PORT MAP (
        A => S858,
        B => S8025,
        Y => S8098
    );
NOR_2957: ENTITY WORK.NOR
    PORT MAP (
        A => S548,
        B => S8007,
        Y => S8099
    );
NOR_2958: ENTITY WORK.NOR
    PORT MAP (
        A => S8098,
        B => S8099,
        Y => S8100
    );
NAND_4721: ENTITY WORK.NAND
    PORT MAP (
        A => S8096,
        B => S8100,
        Y => S8101
    );
NOR_2959: ENTITY WORK.NOR
    PORT MAP (
        A => S8093,
        B => S8101,
        Y => S8102
    );
NOR_2960: ENTITY WORK.NOR
    PORT MAP (
        A => S7941,
        B => S8079,
        Y => S8103
    );
NAND_4722: ENTITY WORK.NAND
    PORT MAP (
        A => S7942,
        B => S8078,
        Y => S8104
    );
NOR_2961: ENTITY WORK.NOR
    PORT MAP (
        A => S7991,
        B => S8104,
        Y => S8105
    );
NOR_2962: ENTITY WORK.NOR
    PORT MAP (
        A => S805,
        B => S8018,
        Y => S8106
    );
NAND_4723: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_8,
        B => S8017,
        Y => S8107
    );
NOR_2963: ENTITY WORK.NOR
    PORT MAP (
        A => S910,
        B => S8003,
        Y => S8109
    );
NAND_4724: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_6,
        B => S8002,
        Y => S8110
    );
NAND_4725: ENTITY WORK.NAND
    PORT MAP (
        A => S8107,
        B => S8110,
        Y => S8111
    );
NAND_4726: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_2,
        B => S7967,
        Y => S8112
    );
NAND_4727: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_14,
        B => S7995,
        Y => S8113
    );
NAND_4728: ENTITY WORK.NAND
    PORT MAP (
        A => S8112,
        B => S8113,
        Y => S8114
    );
NOR_2964: ENTITY WORK.NOR
    PORT MAP (
        A => S8111,
        B => S8114,
        Y => S8115
    );
NAND_4729: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_10,
        B => S7984,
        Y => S8116
    );
NAND_4730: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_11,
        B => S8020,
        Y => S8117
    );
NAND_4731: ENTITY WORK.NAND
    PORT MAP (
        A => S8116,
        B => S8117,
        Y => S8118
    );
NAND_4732: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_3,
        B => S8009,
        Y => S8120
    );
NAND_4733: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_9,
        B => S8030,
        Y => S8121
    );
NAND_4734: ENTITY WORK.NAND
    PORT MAP (
        A => S8120,
        B => S8121,
        Y => S8122
    );
NOR_2965: ENTITY WORK.NOR
    PORT MAP (
        A => S8118,
        B => S8122,
        Y => S8123
    );
NAND_4735: ENTITY WORK.NAND
    PORT MAP (
        A => S8115,
        B => S8123,
        Y => S8124
    );
NOR_2966: ENTITY WORK.NOR
    PORT MAP (
        A => S8105,
        B => S8124,
        Y => S8125
    );
NAND_4736: ENTITY WORK.NAND
    PORT MAP (
        A => S7958,
        B => S8078,
        Y => S8126
    );
NOR_2967: ENTITY WORK.NOR
    PORT MAP (
        A => S7991,
        B => S8079,
        Y => S8127
    );
NAND_4737: ENTITY WORK.NAND
    PORT MAP (
        A => S8102,
        B => S8125,
        Y => datapath_shiftunit_2171_A
    );
NAND_4738: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_7,
        B => S8002,
        Y => S8128
    );
NAND_4739: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_10,
        B => S8030,
        Y => S8130
    );
NAND_4740: ENTITY WORK.NAND
    PORT MAP (
        A => S8128,
        B => S8130,
        Y => S8131
    );
NOR_2968: ENTITY WORK.NOR
    PORT MAP (
        A => S1065,
        B => S7969,
        Y => S8132
    );
NAND_4741: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_3,
        B => S7967,
        Y => S8133
    );
NAND_4742: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_11,
        B => S7984,
        Y => S8134
    );
NAND_4743: ENTITY WORK.NAND
    PORT MAP (
        A => S8133,
        B => S8134,
        Y => S8135
    );
NAND_4744: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_14,
        B => S8006,
        Y => S8136
    );
NOR_2969: ENTITY WORK.NOR
    PORT MAP (
        A => S1611,
        B => S7950,
        Y => S8137
    );
NOR_2970: ENTITY WORK.NOR
    PORT MAP (
        A => S7991,
        B => S8137,
        Y => S8138
    );
NAND_4745: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_15,
        B => S8138,
        Y => S8139
    );
NAND_4746: ENTITY WORK.NAND
    PORT MAP (
        A => S8136,
        B => S8139,
        Y => S8141
    );
NOR_2971: ENTITY WORK.NOR
    PORT MAP (
        A => S8135,
        B => S8141,
        Y => S8142
    );
NOT_553: ENTITY WORK.NOT
    PORT MAP (
        A => S8142,
        Y => S8143
    );
NOR_2972: ENTITY WORK.NOR
    PORT MAP (
        A => S8131,
        B => S8143,
        Y => S8144
    );
NAND_4747: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_4,
        B => S8009,
        Y => S8145
    );
NOR_2973: ENTITY WORK.NOR
    PORT MAP (
        A => S599,
        B => S8021,
        Y => S8146
    );
NOR_2974: ENTITY WORK.NOR
    PORT MAP (
        A => S910,
        B => S7974,
        Y => S8147
    );
NAND_4748: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_6,
        B => S7973,
        Y => S8148
    );
NOR_2975: ENTITY WORK.NOR
    PORT MAP (
        A => S8146,
        B => S8147,
        Y => S8149
    );
NAND_4749: ENTITY WORK.NAND
    PORT MAP (
        A => S8145,
        B => S8149,
        Y => S8150
    );
NOR_2976: ENTITY WORK.NOR
    PORT MAP (
        A => S805,
        B => S8025,
        Y => S8152
    );
NOR_2977: ENTITY WORK.NOR
    PORT MAP (
        A => S963,
        B => S8015,
        Y => S8153
    );
NOR_2978: ENTITY WORK.NOR
    PORT MAP (
        A => S8152,
        B => S8153,
        Y => S8154
    );
NOR_2979: ENTITY WORK.NOR
    PORT MAP (
        A => S548,
        B => S7981,
        Y => S8155
    );
NOR_2980: ENTITY WORK.NOR
    PORT MAP (
        A => S754,
        B => S8018,
        Y => S8156
    );
NAND_4750: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_9,
        B => S8017,
        Y => S8157
    );
NOR_2981: ENTITY WORK.NOR
    PORT MAP (
        A => S8155,
        B => S8156,
        Y => S8158
    );
NAND_4751: ENTITY WORK.NAND
    PORT MAP (
        A => S8154,
        B => S8158,
        Y => S8159
    );
NOR_2982: ENTITY WORK.NOR
    PORT MAP (
        A => S8150,
        B => S8159,
        Y => S8160
    );
NAND_4752: ENTITY WORK.NAND
    PORT MAP (
        A => S8144,
        B => S8160,
        Y => datapath_shiftunit_2189_A
    );
NOR_2983: ENTITY WORK.NOR
    PORT MAP (
        A => S805,
        B => S8003,
        Y => S8162
    );
NOR_2984: ENTITY WORK.NOR
    PORT MAP (
        A => S1304,
        B => S8007,
        Y => S8163
    );
NOR_2985: ENTITY WORK.NOR
    PORT MAP (
        A => S8162,
        B => S8163,
        Y => S8164
    );
NOR_2986: ENTITY WORK.NOR
    PORT MAP (
        A => S754,
        B => S8025,
        Y => S8165
    );
NAND_4753: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_9,
        B => S8024,
        Y => S8166
    );
NOR_2987: ENTITY WORK.NOR
    PORT MAP (
        A => S651,
        B => S8031,
        Y => S8167
    );
NOR_2988: ENTITY WORK.NOR
    PORT MAP (
        A => S8165,
        B => S8167,
        Y => S8168
    );
NAND_4754: ENTITY WORK.NAND
    PORT MAP (
        A => S8164,
        B => S8168,
        Y => S8169
    );
NOR_2989: ENTITY WORK.NOR
    PORT MAP (
        A => S8127,
        B => S8169,
        Y => S8170
    );
NOR_2990: ENTITY WORK.NOR
    PORT MAP (
        A => S858,
        B => S7974,
        Y => S8171
    );
NOR_2991: ENTITY WORK.NOR
    PORT MAP (
        A => S910,
        B => S8015,
        Y => S8173
    );
NOR_2992: ENTITY WORK.NOR
    PORT MAP (
        A => S8171,
        B => S8173,
        Y => S8174
    );
NOR_2993: ENTITY WORK.NOR
    PORT MAP (
        A => S963,
        B => S8010,
        Y => S8175
    );
NAND_4755: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_5,
        B => S8009,
        Y => S8176
    );
NOR_2994: ENTITY WORK.NOR
    PORT MAP (
        A => S1013,
        B => S7969,
        Y => S8177
    );
NAND_4756: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_4,
        B => S7967,
        Y => S8178
    );
NOR_2995: ENTITY WORK.NOR
    PORT MAP (
        A => S8175,
        B => S8177,
        Y => S8179
    );
NAND_4757: ENTITY WORK.NAND
    PORT MAP (
        A => S8174,
        B => S8179,
        Y => S8180
    );
NOR_2996: ENTITY WORK.NOR
    PORT MAP (
        A => S548,
        B => S8021,
        Y => S8181
    );
NOR_2997: ENTITY WORK.NOR
    PORT MAP (
        A => S702,
        B => S8018,
        Y => S8182
    );
NOR_2998: ENTITY WORK.NOR
    PORT MAP (
        A => S8181,
        B => S8182,
        Y => S8184
    );
NOR_2999: ENTITY WORK.NOR
    PORT MAP (
        A => S492,
        B => S7981,
        Y => S8185
    );
NOR_3000: ENTITY WORK.NOR
    PORT MAP (
        A => S599,
        B => S7985,
        Y => S8186
    );
NOR_3001: ENTITY WORK.NOR
    PORT MAP (
        A => S8185,
        B => S8186,
        Y => S8187
    );
NAND_4758: ENTITY WORK.NAND
    PORT MAP (
        A => S8184,
        B => S8187,
        Y => S8188
    );
NOR_3002: ENTITY WORK.NOR
    PORT MAP (
        A => S8180,
        B => S8188,
        Y => S8189
    );
NAND_4759: ENTITY WORK.NAND
    PORT MAP (
        A => S8170,
        B => S8189,
        Y => datapath_shiftunit_2207_A
    );
NOR_3003: ENTITY WORK.NOR
    PORT MAP (
        A => S7990,
        B => S8006,
        Y => S8190
    );
NOR_3004: ENTITY WORK.NOR
    PORT MAP (
        A => S8079,
        B => S8190,
        Y => S8191
    );
NOR_3005: ENTITY WORK.NOR
    PORT MAP (
        A => S492,
        B => S8021,
        Y => S8192
    );
NOR_3006: ENTITY WORK.NOR
    PORT MAP (
        A => S910,
        B => S8010,
        Y => S8194
    );
NOR_3007: ENTITY WORK.NOR
    PORT MAP (
        A => S8192,
        B => S8194,
        Y => S8195
    );
NOR_3008: ENTITY WORK.NOR
    PORT MAP (
        A => S651,
        B => S8018,
        Y => S8196
    );
NOR_3009: ENTITY WORK.NOR
    PORT MAP (
        A => S805,
        B => S7974,
        Y => S8197
    );
NOR_3010: ENTITY WORK.NOR
    PORT MAP (
        A => S8196,
        B => S8197,
        Y => S8198
    );
NAND_4760: ENTITY WORK.NAND
    PORT MAP (
        A => S8195,
        B => S8198,
        Y => S8199
    );
NOR_3011: ENTITY WORK.NOR
    PORT MAP (
        A => S8191,
        B => S8199,
        Y => S8200
    );
NAND_4761: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_10,
        B => S8024,
        Y => S8201
    );
NOR_3012: ENTITY WORK.NOR
    PORT MAP (
        A => S858,
        B => S8015,
        Y => S8202
    );
NOR_3013: ENTITY WORK.NOR
    PORT MAP (
        A => S754,
        B => S8003,
        Y => S8203
    );
NOR_3014: ENTITY WORK.NOR
    PORT MAP (
        A => S8202,
        B => S8203,
        Y => S8205
    );
NAND_4762: ENTITY WORK.NAND
    PORT MAP (
        A => S8201,
        B => S8205,
        Y => S8206
    );
NOR_3015: ENTITY WORK.NOR
    PORT MAP (
        A => S1304,
        B => S7981,
        Y => S8207
    );
NOR_3016: ENTITY WORK.NOR
    PORT MAP (
        A => S599,
        B => S8031,
        Y => S8208
    );
NOR_3017: ENTITY WORK.NOR
    PORT MAP (
        A => S8207,
        B => S8208,
        Y => S8209
    );
NOR_3018: ENTITY WORK.NOR
    PORT MAP (
        A => S963,
        B => S7969,
        Y => S8210
    );
NOR_3019: ENTITY WORK.NOR
    PORT MAP (
        A => S548,
        B => S7985,
        Y => S8211
    );
NOR_3020: ENTITY WORK.NOR
    PORT MAP (
        A => S8210,
        B => S8211,
        Y => S8212
    );
NAND_4763: ENTITY WORK.NAND
    PORT MAP (
        A => S8209,
        B => S8212,
        Y => S8213
    );
NOR_3021: ENTITY WORK.NOR
    PORT MAP (
        A => S8206,
        B => S8213,
        Y => S8214
    );
NAND_4764: ENTITY WORK.NAND
    PORT MAP (
        A => S8200,
        B => S8214,
        Y => datapath_shiftunit_2225_A
    );
NOR_3022: ENTITY WORK.NOR
    PORT MAP (
        A => S548,
        B => S8031,
        Y => S8216
    );
NOR_3023: ENTITY WORK.NOR
    PORT MAP (
        A => S651,
        B => S8025,
        Y => S8217
    );
NOR_3024: ENTITY WORK.NOR
    PORT MAP (
        A => S805,
        B => S8015,
        Y => S8218
    );
NAND_4765: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_15,
        B => S8020,
        Y => S8219
    );
NOR_3025: ENTITY WORK.NOR
    PORT MAP (
        A => S858,
        B => S8010,
        Y => S8220
    );
NAND_4766: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_7,
        B => S8009,
        Y => S8221
    );
NAND_4767: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_9,
        B => S7973,
        Y => S8222
    );
NAND_4768: ENTITY WORK.NAND
    PORT MAP (
        A => S7981,
        B => S8190,
        Y => S8223
    );
NAND_4769: ENTITY WORK.NAND
    PORT MAP (
        A => S8078,
        B => S8223,
        Y => S8224
    );
NOR_3026: ENTITY WORK.NOR
    PORT MAP (
        A => S492,
        B => S7985,
        Y => S8226
    );
NOR_3027: ENTITY WORK.NOR
    PORT MAP (
        A => S599,
        B => S8018,
        Y => S8227
    );
NAND_4770: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_10,
        B => S8002,
        Y => S8228
    );
NOR_3028: ENTITY WORK.NOR
    PORT MAP (
        A => S910,
        B => S7969,
        Y => S8229
    );
NAND_4771: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_6,
        B => S7967,
        Y => S8230
    );
NOR_3029: ENTITY WORK.NOR
    PORT MAP (
        A => S8217,
        B => S8218,
        Y => S8231
    );
NOR_3030: ENTITY WORK.NOR
    PORT MAP (
        A => S8216,
        B => S8226,
        Y => S8232
    );
NAND_4772: ENTITY WORK.NAND
    PORT MAP (
        A => S8221,
        B => S8232,
        Y => S8233
    );
NAND_4773: ENTITY WORK.NAND
    PORT MAP (
        A => S8224,
        B => S8231,
        Y => S8234
    );
NOR_3031: ENTITY WORK.NOR
    PORT MAP (
        A => S8233,
        B => S8234,
        Y => S8235
    );
NAND_4774: ENTITY WORK.NAND
    PORT MAP (
        A => S8219,
        B => S8228,
        Y => S8237
    );
NOR_3032: ENTITY WORK.NOR
    PORT MAP (
        A => S8227,
        B => S8229,
        Y => S8238
    );
NAND_4775: ENTITY WORK.NAND
    PORT MAP (
        A => S8222,
        B => S8238,
        Y => S8239
    );
NOR_3033: ENTITY WORK.NOR
    PORT MAP (
        A => S8237,
        B => S8239,
        Y => S8240
    );
NAND_4776: ENTITY WORK.NAND
    PORT MAP (
        A => S8235,
        B => S8240,
        Y => datapath_shiftunit_2243_A
    );
NOR_3034: ENTITY WORK.NOR
    PORT MAP (
        A => S702,
        B => S7974,
        Y => S8241
    );
NAND_4777: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_10,
        B => S7973,
        Y => S8242
    );
NOR_3035: ENTITY WORK.NOR
    PORT MAP (
        A => S548,
        B => S8018,
        Y => S8243
    );
NOR_3036: ENTITY WORK.NOR
    PORT MAP (
        A => S754,
        B => S8015,
        Y => S8244
    );
NAND_4778: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_11,
        B => S8002,
        Y => S8245
    );
NOR_3037: ENTITY WORK.NOR
    PORT MAP (
        A => S858,
        B => S7969,
        Y => S8247
    );
NOR_3038: ENTITY WORK.NOR
    PORT MAP (
        A => S1304,
        B => S7985,
        Y => S8248
    );
NOR_3039: ENTITY WORK.NOR
    PORT MAP (
        A => S599,
        B => S8025,
        Y => S8249
    );
NOR_3040: ENTITY WORK.NOR
    PORT MAP (
        A => S492,
        B => S8031,
        Y => S8250
    );
NOR_3041: ENTITY WORK.NOR
    PORT MAP (
        A => S805,
        B => S8010,
        Y => S8251
    );
NOR_3042: ENTITY WORK.NOR
    PORT MAP (
        A => S8247,
        B => S8249,
        Y => S8252
    );
NOR_3043: ENTITY WORK.NOR
    PORT MAP (
        A => S8241,
        B => S8251,
        Y => S8253
    );
NAND_4779: ENTITY WORK.NAND
    PORT MAP (
        A => S8252,
        B => S8253,
        Y => S8254
    );
NOR_3044: ENTITY WORK.NOR
    PORT MAP (
        A => S8021,
        B => S8079,
        Y => S8255
    );
NOR_3045: ENTITY WORK.NOR
    PORT MAP (
        A => S8254,
        B => S8255,
        Y => S8256
    );
NOR_3046: ENTITY WORK.NOR
    PORT MAP (
        A => S8243,
        B => S8248,
        Y => S8258
    );
NAND_4780: ENTITY WORK.NAND
    PORT MAP (
        A => S8245,
        B => S8258,
        Y => S8259
    );
NOR_3047: ENTITY WORK.NOR
    PORT MAP (
        A => S8244,
        B => S8250,
        Y => S8260
    );
NAND_4781: ENTITY WORK.NAND
    PORT MAP (
        A => S8224,
        B => S8260,
        Y => S8261
    );
NOR_3048: ENTITY WORK.NOR
    PORT MAP (
        A => S8259,
        B => S8261,
        Y => S8262
    );
NAND_4782: ENTITY WORK.NAND
    PORT MAP (
        A => S8256,
        B => S8262,
        Y => datapath_shiftunit_2261_A
    );
NOR_3049: ENTITY WORK.NOR
    PORT MAP (
        A => S1304,
        B => S8031,
        Y => S8263
    );
NOR_3050: ENTITY WORK.NOR
    PORT MAP (
        A => S548,
        B => S8025,
        Y => S8264
    );
NOR_3051: ENTITY WORK.NOR
    PORT MAP (
        A => S754,
        B => S8010,
        Y => S8265
    );
NOR_3052: ENTITY WORK.NOR
    PORT MAP (
        A => S599,
        B => S8003,
        Y => S8266
    );
NOR_3053: ENTITY WORK.NOR
    PORT MAP (
        A => S492,
        B => S8018,
        Y => S8268
    );
NOR_3054: ENTITY WORK.NOR
    PORT MAP (
        A => S651,
        B => S7974,
        Y => S8269
    );
NOR_3055: ENTITY WORK.NOR
    PORT MAP (
        A => S805,
        B => S7969,
        Y => S8270
    );
NOR_3056: ENTITY WORK.NOR
    PORT MAP (
        A => S702,
        B => S8015,
        Y => S8271
    );
NAND_4783: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_10,
        B => S8014,
        Y => S8272
    );
NOR_3057: ENTITY WORK.NOR
    PORT MAP (
        A => S8265,
        B => S8268,
        Y => S8273
    );
NOR_3058: ENTITY WORK.NOR
    PORT MAP (
        A => S8266,
        B => S8270,
        Y => S8274
    );
NAND_4784: ENTITY WORK.NAND
    PORT MAP (
        A => S8126,
        B => S8274,
        Y => S8275
    );
NOR_3059: ENTITY WORK.NOR
    PORT MAP (
        A => S8263,
        B => S8269,
        Y => S8276
    );
NOR_3060: ENTITY WORK.NOR
    PORT MAP (
        A => S8264,
        B => S8271,
        Y => S8277
    );
NAND_4785: ENTITY WORK.NAND
    PORT MAP (
        A => S8276,
        B => S8277,
        Y => S8279
    );
NOR_3061: ENTITY WORK.NOR
    PORT MAP (
        A => S8275,
        B => S8279,
        Y => S8280
    );
NAND_4786: ENTITY WORK.NAND
    PORT MAP (
        A => S8273,
        B => S8280,
        Y => datapath_shiftunit_2279_A
    );
NAND_4787: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_12,
        B => S7973,
        Y => S8281
    );
NAND_4788: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_13,
        B => S8002,
        Y => S8282
    );
NAND_4789: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_14,
        B => S8024,
        Y => S8283
    );
NOR_3062: ENTITY WORK.NOR
    PORT MAP (
        A => S7941,
        B => S7963,
        Y => S8284
    );
NOR_3063: ENTITY WORK.NOR
    PORT MAP (
        A => S7958,
        B => S8284,
        Y => S8285
    );
NAND_4790: ENTITY WORK.NAND
    PORT MAP (
        A => S1612,
        B => S8018,
        Y => S8286
    );
NAND_4791: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_15,
        B => S8286,
        Y => S8287
    );
NOR_3064: ENTITY WORK.NOR
    PORT MAP (
        A => S8285,
        B => S8287,
        Y => S8289
    );
NAND_4792: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_10,
        B => S8009,
        Y => S8290
    );
NAND_4793: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_11,
        B => S8014,
        Y => S8291
    );
NOR_3065: ENTITY WORK.NOR
    PORT MAP (
        A => S754,
        B => S7969,
        Y => S8292
    );
NAND_4794: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_9,
        B => S7967,
        Y => S8293
    );
NAND_4795: ENTITY WORK.NAND
    PORT MAP (
        A => S8283,
        B => S8293,
        Y => S8294
    );
NAND_4796: ENTITY WORK.NAND
    PORT MAP (
        A => S8281,
        B => S8290,
        Y => S8295
    );
NOR_3066: ENTITY WORK.NOR
    PORT MAP (
        A => S8294,
        B => S8295,
        Y => S8296
    );
NAND_4797: ENTITY WORK.NAND
    PORT MAP (
        A => S8282,
        B => S8291,
        Y => S8297
    );
NOR_3067: ENTITY WORK.NOR
    PORT MAP (
        A => S8289,
        B => S8297,
        Y => S8298
    );
NAND_4798: ENTITY WORK.NAND
    PORT MAP (
        A => S8296,
        B => S8298,
        Y => datapath_shiftunit_2297_A
    );
NOR_3068: ENTITY WORK.NOR
    PORT MAP (
        A => S651,
        B => S8010,
        Y => S8300
    );
NAND_4799: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_11,
        B => S8009,
        Y => S8301
    );
NOR_3069: ENTITY WORK.NOR
    PORT MAP (
        A => S702,
        B => S7969,
        Y => S8302
    );
NAND_4800: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_10,
        B => S7967,
        Y => S8303
    );
NAND_4801: ENTITY WORK.NAND
    PORT MAP (
        A => S8301,
        B => S8303,
        Y => S8304
    );
NAND_4802: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_13,
        B => S7973,
        Y => S8305
    );
NAND_4803: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_15,
        B => S8024,
        Y => S8306
    );
NAND_4804: ENTITY WORK.NAND
    PORT MAP (
        A => S8305,
        B => S8306,
        Y => S8307
    );
NOR_3070: ENTITY WORK.NOR
    PORT MAP (
        A => S8304,
        B => S8307,
        Y => S8308
    );
NAND_4805: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_12,
        B => S8014,
        Y => S8310
    );
NAND_4806: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_14,
        B => S8002,
        Y => S8311
    );
NAND_4807: ENTITY WORK.NAND
    PORT MAP (
        A => S8310,
        B => S8311,
        Y => S8312
    );
NOR_3071: ENTITY WORK.NOR
    PORT MAP (
        A => S8079,
        B => S8285,
        Y => S8313
    );
NOR_3072: ENTITY WORK.NOR
    PORT MAP (
        A => S8312,
        B => S8313,
        Y => S8314
    );
NAND_4808: ENTITY WORK.NAND
    PORT MAP (
        A => S8308,
        B => S8314,
        Y => datapath_shiftunit_2315_A
    );
NAND_4809: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_15,
        B => S8002,
        Y => S8315
    );
NAND_4810: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_13,
        B => S8014,
        Y => S8316
    );
NOR_3073: ENTITY WORK.NOR
    PORT MAP (
        A => S492,
        B => S7974,
        Y => S8317
    );
NOR_3074: ENTITY WORK.NOR
    PORT MAP (
        A => S8025,
        B => S8079,
        Y => S8318
    );
NAND_4811: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_11,
        B => S7967,
        Y => S8320
    );
NOR_3075: ENTITY WORK.NOR
    PORT MAP (
        A => S599,
        B => S8010,
        Y => S8321
    );
NAND_4812: ENTITY WORK.NAND
    PORT MAP (
        A => S8315,
        B => S8316,
        Y => S8322
    );
NOR_3076: ENTITY WORK.NOR
    PORT MAP (
        A => S8313,
        B => S8322,
        Y => S8323
    );
NOR_3077: ENTITY WORK.NOR
    PORT MAP (
        A => S8317,
        B => S8321,
        Y => S8324
    );
NAND_4813: ENTITY WORK.NAND
    PORT MAP (
        A => S8320,
        B => S8324,
        Y => S8325
    );
NOR_3078: ENTITY WORK.NOR
    PORT MAP (
        A => S8318,
        B => S8325,
        Y => S8326
    );
NAND_4814: ENTITY WORK.NAND
    PORT MAP (
        A => S8323,
        B => S8326,
        Y => datapath_shiftunit_2333_A
    );
NAND_4815: ENTITY WORK.NAND
    PORT MAP (
        A => S7966,
        B => S8078,
        Y => S8327
    );
NOR_3079: ENTITY WORK.NOR
    PORT MAP (
        A => S599,
        B => S7969,
        Y => S8328
    );
NAND_4816: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_12,
        B => S7967,
        Y => S8330
    );
NAND_4817: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_15,
        B => S7973,
        Y => S8331
    );
NAND_4818: ENTITY WORK.NAND
    PORT MAP (
        A => S8330,
        B => S8331,
        Y => S8332
    );
NAND_4819: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_13,
        B => S8009,
        Y => S8333
    );
NAND_4820: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_14,
        B => S8014,
        Y => S8334
    );
NAND_4821: ENTITY WORK.NAND
    PORT MAP (
        A => S8333,
        B => S8334,
        Y => S8335
    );
NOR_3080: ENTITY WORK.NOR
    PORT MAP (
        A => S8332,
        B => S8335,
        Y => S8336
    );
NAND_4822: ENTITY WORK.NAND
    PORT MAP (
        A => S8327,
        B => S8336,
        Y => datapath_shiftunit_2351_A
    );
NOR_3081: ENTITY WORK.NOR
    PORT MAP (
        A => S7966,
        B => S7971,
        Y => S8337
    );
NOR_3082: ENTITY WORK.NOR
    PORT MAP (
        A => S8079,
        B => S8337,
        Y => S8338
    );
NAND_4823: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_14,
        B => S8009,
        Y => S8340
    );
NOR_3083: ENTITY WORK.NOR
    PORT MAP (
        A => S548,
        B => S7969,
        Y => S8341
    );
NAND_4824: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_13,
        B => S7967,
        Y => S8342
    );
NAND_4825: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_15,
        B => S8014,
        Y => S8343
    );
NAND_4826: ENTITY WORK.NAND
    PORT MAP (
        A => S8340,
        B => S8342,
        Y => S8344
    );
NOR_3084: ENTITY WORK.NOR
    PORT MAP (
        A => S8338,
        B => S8344,
        Y => S8345
    );
NAND_4827: ENTITY WORK.NAND
    PORT MAP (
        A => S8343,
        B => S8345,
        Y => datapath_shiftunit_2369_A
    );
NAND_4828: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_15,
        B => S8009,
        Y => S8346
    );
NAND_4829: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_14,
        B => S7967,
        Y => S8347
    );
NAND_4830: ENTITY WORK.NAND
    PORT MAP (
        A => S8346,
        B => S8347,
        Y => S8348
    );
NOR_3085: ENTITY WORK.NOR
    PORT MAP (
        A => S8103,
        B => S8348,
        Y => S8350
    );
NAND_4831: ENTITY WORK.NAND
    PORT MAP (
        A => S8327,
        B => S8350,
        Y => datapath_shiftunit_2387_A
    );
NAND_4832: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_15,
        B => S7967,
        Y => S8351
    );
NAND_4833: ENTITY WORK.NAND
    PORT MAP (
        A => S8079,
        B => S8351,
        Y => datapath_shiftunit_2405_A
    );
NAND_4834: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_0,
        B => S8009,
        Y => S8352
    );
NAND_4835: ENTITY WORK.NAND
    PORT MAP (
        A => S8067,
        B => S8352,
        Y => datapath_shiftunit_2457_A
    );
NOR_3086: ENTITY WORK.NOR
    PORT MAP (
        A => S1220,
        B => S8015,
        Y => S8353
    );
NOR_3087: ENTITY WORK.NOR
    PORT MAP (
        A => S8012,
        B => S8353,
        Y => S8354
    );
NAND_4836: ENTITY WORK.NAND
    PORT MAP (
        A => S8112,
        B => S8354,
        Y => datapath_shiftunit_2475_A
    );
NOR_3088: ENTITY WORK.NOR
    PORT MAP (
        A => S8055,
        B => S8132,
        Y => S8355
    );
NOR_3089: ENTITY WORK.NOR
    PORT MAP (
        A => S1220,
        B => S7974,
        Y => S8357
    );
NOR_3090: ENTITY WORK.NOR
    PORT MAP (
        A => S1168,
        B => S8015,
        Y => S8358
    );
NOR_3091: ENTITY WORK.NOR
    PORT MAP (
        A => S8357,
        B => S8358,
        Y => S8359
    );
NAND_4837: ENTITY WORK.NAND
    PORT MAP (
        A => S8355,
        B => S8359,
        Y => datapath_shiftunit_2493_A
    );
NAND_4838: ENTITY WORK.NAND
    PORT MAP (
        A => S8016,
        B => S8120,
        Y => S8360
    );
NAND_4839: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_1,
        B => S7973,
        Y => S8361
    );
NAND_4840: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_0,
        B => S8002,
        Y => S8362
    );
NAND_4841: ENTITY WORK.NAND
    PORT MAP (
        A => S8178,
        B => S8362,
        Y => S8363
    );
NOR_3092: ENTITY WORK.NOR
    PORT MAP (
        A => S8360,
        B => S8363,
        Y => S8364
    );
NAND_4842: ENTITY WORK.NAND
    PORT MAP (
        A => S8361,
        B => S8364,
        Y => datapath_shiftunit_2511_A
    );
NAND_4843: ENTITY WORK.NAND
    PORT MAP (
        A => S8060,
        B => S8145,
        Y => S8366
    );
NAND_4844: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_0,
        B => S8024,
        Y => S8367
    );
NAND_4845: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_2,
        B => S7973,
        Y => S8368
    );
NOR_3093: ENTITY WORK.NOR
    PORT MAP (
        A => S1168,
        B => S8003,
        Y => S8369
    );
NOR_3094: ENTITY WORK.NOR
    PORT MAP (
        A => S8210,
        B => S8369,
        Y => S8370
    );
NAND_4846: ENTITY WORK.NAND
    PORT MAP (
        A => S8367,
        B => S8368,
        Y => S8371
    );
NOR_3095: ENTITY WORK.NOR
    PORT MAP (
        A => S8366,
        B => S8371,
        Y => S8372
    );
NAND_4847: ENTITY WORK.NAND
    PORT MAP (
        A => S8370,
        B => S8372,
        Y => datapath_shiftunit_2529_A
    );
NOR_3096: ENTITY WORK.NOR
    PORT MAP (
        A => S1116,
        B => S8003,
        Y => S8373
    );
NAND_4848: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_1,
        B => S8024,
        Y => S8374
    );
NAND_4849: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_0,
        B => S8017,
        Y => S8376
    );
NAND_4850: ENTITY WORK.NAND
    PORT MAP (
        A => S8374,
        B => S8376,
        Y => S8377
    );
NOR_3097: ENTITY WORK.NOR
    PORT MAP (
        A => S8373,
        B => S8377,
        Y => S8378
    );
NAND_4851: ENTITY WORK.NAND
    PORT MAP (
        A => S7975,
        B => S8091,
        Y => S8379
    );
NAND_4852: ENTITY WORK.NAND
    PORT MAP (
        A => S8176,
        B => S8230,
        Y => S8380
    );
NOR_3098: ENTITY WORK.NOR
    PORT MAP (
        A => S8379,
        B => S8380,
        Y => S8381
    );
NAND_4853: ENTITY WORK.NAND
    PORT MAP (
        A => S8378,
        B => S8381,
        Y => datapath_shiftunit_2547_A
    );
NOR_3099: ENTITY WORK.NOR
    PORT MAP (
        A => S8153,
        B => S8194,
        Y => S8382
    );
NOR_3100: ENTITY WORK.NOR
    PORT MAP (
        A => S8063,
        B => S8247,
        Y => S8383
    );
NAND_4854: ENTITY WORK.NAND
    PORT MAP (
        A => S8382,
        B => S8383,
        Y => S8384
    );
NAND_4855: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_1,
        B => S8017,
        Y => S8386
    );
NOR_3101: ENTITY WORK.NOR
    PORT MAP (
        A => S1220,
        B => S8031,
        Y => S8387
    );
NAND_4856: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_2,
        B => S8024,
        Y => S8388
    );
NOR_3102: ENTITY WORK.NOR
    PORT MAP (
        A => S1065,
        B => S8003,
        Y => S8389
    );
NAND_4857: ENTITY WORK.NAND
    PORT MAP (
        A => S8386,
        B => S8388,
        Y => S8390
    );
NOR_3103: ENTITY WORK.NOR
    PORT MAP (
        A => S8389,
        B => S8390,
        Y => S8391
    );
NOR_3104: ENTITY WORK.NOR
    PORT MAP (
        A => S8384,
        B => S8387,
        Y => S8392
    );
NAND_4858: ENTITY WORK.NAND
    PORT MAP (
        A => S8391,
        B => S8392,
        Y => datapath_shiftunit_2565_A
    );
NOR_3105: ENTITY WORK.NOR
    PORT MAP (
        A => S1220,
        B => S7985,
        Y => S8393
    );
NAND_4859: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_2,
        B => S8017,
        Y => S8394
    );
NAND_4860: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_3,
        B => S8024,
        Y => S8396
    );
NAND_4861: ENTITY WORK.NAND
    PORT MAP (
        A => S8394,
        B => S8396,
        Y => S8397
    );
NOR_3106: ENTITY WORK.NOR
    PORT MAP (
        A => S8393,
        B => S8397,
        Y => S8398
    );
NAND_4862: ENTITY WORK.NAND
    PORT MAP (
        A => S8005,
        B => S8092,
        Y => S8399
    );
NOR_3107: ENTITY WORK.NOR
    PORT MAP (
        A => S8173,
        B => S8220,
        Y => S8400
    );
NOR_3108: ENTITY WORK.NOR
    PORT MAP (
        A => S1168,
        B => S8031,
        Y => S8401
    );
NOR_3109: ENTITY WORK.NOR
    PORT MAP (
        A => S8270,
        B => S8401,
        Y => S8402
    );
NAND_4863: ENTITY WORK.NAND
    PORT MAP (
        A => S8400,
        B => S8402,
        Y => S8403
    );
NOR_3110: ENTITY WORK.NOR
    PORT MAP (
        A => S8399,
        B => S8403,
        Y => S8404
    );
NAND_4864: ENTITY WORK.NAND
    PORT MAP (
        A => S8398,
        B => S8404,
        Y => datapath_shiftunit_2583_A
    );
NAND_4865: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_1,
        B => S7984,
        Y => S8406
    );
NAND_4866: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_0,
        B => S8020,
        Y => S8407
    );
NAND_4867: ENTITY WORK.NAND
    PORT MAP (
        A => S8406,
        B => S8407,
        Y => S8408
    );
NAND_4868: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_3,
        B => S8017,
        Y => S8409
    );
NAND_4869: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_4,
        B => S8024,
        Y => S8410
    );
NAND_4870: ENTITY WORK.NAND
    PORT MAP (
        A => S8409,
        B => S8410,
        Y => S8411
    );
NOR_3111: ENTITY WORK.NOR
    PORT MAP (
        A => S8408,
        B => S8411,
        Y => S8412
    );
NAND_4871: ENTITY WORK.NAND
    PORT MAP (
        A => S8058,
        B => S8148,
        Y => S8413
    );
NOR_3112: ENTITY WORK.NOR
    PORT MAP (
        A => S8202,
        B => S8251,
        Y => S8414
    );
NOR_3113: ENTITY WORK.NOR
    PORT MAP (
        A => S1116,
        B => S8031,
        Y => S8415
    );
NOR_3114: ENTITY WORK.NOR
    PORT MAP (
        A => S8292,
        B => S8415,
        Y => S8417
    );
NAND_4872: ENTITY WORK.NAND
    PORT MAP (
        A => S8414,
        B => S8417,
        Y => S8418
    );
NOR_3115: ENTITY WORK.NOR
    PORT MAP (
        A => S8413,
        B => S8418,
        Y => S8419
    );
NAND_4873: ENTITY WORK.NAND
    PORT MAP (
        A => S8412,
        B => S8419,
        Y => datapath_shiftunit_2601_A
    );
NOR_3116: ENTITY WORK.NOR
    PORT MAP (
        A => S1220,
        B => S7981,
        Y => S8420
    );
NAND_4874: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_2,
        B => S7984,
        Y => S8421
    );
NAND_4875: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_1,
        B => S8020,
        Y => S8422
    );
NAND_4876: ENTITY WORK.NAND
    PORT MAP (
        A => S8421,
        B => S8422,
        Y => S8423
    );
NOR_3117: ENTITY WORK.NOR
    PORT MAP (
        A => S8420,
        B => S8423,
        Y => S8424
    );
NOR_3118: ENTITY WORK.NOR
    PORT MAP (
        A => S8265,
        B => S8302,
        Y => S8425
    );
NOR_3119: ENTITY WORK.NOR
    PORT MAP (
        A => S1065,
        B => S8031,
        Y => S8427
    );
NOR_3120: ENTITY WORK.NOR
    PORT MAP (
        A => S1013,
        B => S8018,
        Y => S8428
    );
NOR_3121: ENTITY WORK.NOR
    PORT MAP (
        A => S8427,
        B => S8428,
        Y => S8429
    );
NAND_4877: ENTITY WORK.NAND
    PORT MAP (
        A => S8425,
        B => S8429,
        Y => S8430
    );
NOR_3122: ENTITY WORK.NOR
    PORT MAP (
        A => S8026,
        B => S8109,
        Y => S8431
    );
NOR_3123: ENTITY WORK.NOR
    PORT MAP (
        A => S8171,
        B => S8218,
        Y => S8432
    );
NAND_4878: ENTITY WORK.NAND
    PORT MAP (
        A => S8431,
        B => S8432,
        Y => S8433
    );
NOR_3124: ENTITY WORK.NOR
    PORT MAP (
        A => S8430,
        B => S8433,
        Y => S8434
    );
NAND_4879: ENTITY WORK.NAND
    PORT MAP (
        A => S8424,
        B => S8434,
        Y => datapath_shiftunit_2619_A
    );
NOR_3125: ENTITY WORK.NOR
    PORT MAP (
        A => S1065,
        B => S7985,
        Y => S8435
    );
NOR_3126: ENTITY WORK.NOR
    PORT MAP (
        A => S1116,
        B => S8021,
        Y => S8437
    );
NOR_3127: ENTITY WORK.NOR
    PORT MAP (
        A => S1220,
        B => S8007,
        Y => S8438
    );
NOR_3128: ENTITY WORK.NOR
    PORT MAP (
        A => S963,
        B => S8018,
        Y => S8439
    );
NOR_3129: ENTITY WORK.NOR
    PORT MAP (
        A => S1168,
        B => S7981,
        Y => S8440
    );
NOR_3130: ENTITY WORK.NOR
    PORT MAP (
        A => S1013,
        B => S8031,
        Y => S8441
    );
NOR_3131: ENTITY WORK.NOR
    PORT MAP (
        A => S8197,
        B => S8438,
        Y => S8442
    );
NOR_3132: ENTITY WORK.NOR
    PORT MAP (
        A => S8439,
        B => S8440,
        Y => S8443
    );
NAND_4880: ENTITY WORK.NAND
    PORT MAP (
        A => S8442,
        B => S8443,
        Y => S8444
    );
NAND_4881: ENTITY WORK.NAND
    PORT MAP (
        A => S8053,
        B => S8290,
        Y => S8445
    );
NOR_3133: ENTITY WORK.NOR
    PORT MAP (
        A => S8444,
        B => S8445,
        Y => S8446
    );
NAND_4882: ENTITY WORK.NAND
    PORT MAP (
        A => S8128,
        B => S8320,
        Y => S8448
    );
NOR_3134: ENTITY WORK.NOR
    PORT MAP (
        A => S8244,
        B => S8435,
        Y => S8449
    );
NOR_3135: ENTITY WORK.NOR
    PORT MAP (
        A => S8437,
        B => S8441,
        Y => S8450
    );
NAND_4883: ENTITY WORK.NAND
    PORT MAP (
        A => S8449,
        B => S8450,
        Y => S8451
    );
NOR_3136: ENTITY WORK.NOR
    PORT MAP (
        A => S8448,
        B => S8451,
        Y => S8452
    );
NAND_4884: ENTITY WORK.NAND
    PORT MAP (
        A => S8446,
        B => S8452,
        Y => datapath_shiftunit_2637_A
    );
NOR_3137: ENTITY WORK.NOR
    PORT MAP (
        A => S8019,
        B => S8098,
        Y => S8453
    );
NOR_3138: ENTITY WORK.NOR
    PORT MAP (
        A => S963,
        B => S8031,
        Y => S8454
    );
NOR_3139: ENTITY WORK.NOR
    PORT MAP (
        A => S1065,
        B => S8021,
        Y => S8455
    );
NOR_3140: ENTITY WORK.NOR
    PORT MAP (
        A => S1013,
        B => S7985,
        Y => S8456
    );
NAND_4885: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_0,
        B => S7995,
        Y => S8458
    );
NOR_3141: ENTITY WORK.NOR
    PORT MAP (
        A => S1168,
        B => S8007,
        Y => S8459
    );
NOR_3142: ENTITY WORK.NOR
    PORT MAP (
        A => S1116,
        B => S7981,
        Y => S8460
    );
NOR_3143: ENTITY WORK.NOR
    PORT MAP (
        A => S8162,
        B => S8300,
        Y => S8461
    );
NAND_4886: ENTITY WORK.NAND
    PORT MAP (
        A => S8453,
        B => S8461,
        Y => S8462
    );
NOR_3144: ENTITY WORK.NOR
    PORT MAP (
        A => S8455,
        B => S8459,
        Y => S8463
    );
NAND_4887: ENTITY WORK.NAND
    PORT MAP (
        A => S8458,
        B => S8463,
        Y => S8464
    );
NOR_3145: ENTITY WORK.NOR
    PORT MAP (
        A => S8462,
        B => S8464,
        Y => S8465
    );
NAND_4888: ENTITY WORK.NAND
    PORT MAP (
        A => S8222,
        B => S8272,
        Y => S8466
    );
NOR_3146: ENTITY WORK.NOR
    PORT MAP (
        A => S8456,
        B => S8460,
        Y => S8467
    );
NOR_3147: ENTITY WORK.NOR
    PORT MAP (
        A => S8328,
        B => S8454,
        Y => S8469
    );
NAND_4889: ENTITY WORK.NAND
    PORT MAP (
        A => S8467,
        B => S8469,
        Y => S8470
    );
NOR_3148: ENTITY WORK.NOR
    PORT MAP (
        A => S8466,
        B => S8470,
        Y => S8471
    );
NAND_4890: ENTITY WORK.NAND
    PORT MAP (
        A => S8465,
        B => S8471,
        Y => datapath_shiftunit_2655_A
    );
NOR_3149: ENTITY WORK.NOR
    PORT MAP (
        A => S8061,
        B => S8152,
        Y => S8472
    );
NOR_3150: ENTITY WORK.NOR
    PORT MAP (
        A => S1168,
        B => S7996,
        Y => S8473
    );
NOR_3151: ENTITY WORK.NOR
    PORT MAP (
        A => S1013,
        B => S8021,
        Y => S8474
    );
NOR_3152: ENTITY WORK.NOR
    PORT MAP (
        A => S8473,
        B => S8474,
        Y => S8475
    );
NOR_3153: ENTITY WORK.NOR
    PORT MAP (
        A => S1116,
        B => S8007,
        Y => S8476
    );
NOR_3154: ENTITY WORK.NOR
    PORT MAP (
        A => S1065,
        B => S7981,
        Y => S8477
    );
NOR_3155: ENTITY WORK.NOR
    PORT MAP (
        A => S910,
        B => S8031,
        Y => S8479
    );
NOR_3156: ENTITY WORK.NOR
    PORT MAP (
        A => S963,
        B => S7985,
        Y => S8480
    );
NOR_3157: ENTITY WORK.NOR
    PORT MAP (
        A => S1220,
        B => S7992,
        Y => S8481
    );
NOR_3158: ENTITY WORK.NOR
    PORT MAP (
        A => S8203,
        B => S8321,
        Y => S8482
    );
NAND_4891: ENTITY WORK.NAND
    PORT MAP (
        A => S8472,
        B => S8482,
        Y => S8483
    );
NOR_3159: ENTITY WORK.NOR
    PORT MAP (
        A => S8479,
        B => S8480,
        Y => S8484
    );
NOR_3160: ENTITY WORK.NOR
    PORT MAP (
        A => S8477,
        B => S8481,
        Y => S8485
    );
NAND_4892: ENTITY WORK.NAND
    PORT MAP (
        A => S8484,
        B => S8485,
        Y => S8486
    );
NOR_3161: ENTITY WORK.NOR
    PORT MAP (
        A => S8483,
        B => S8486,
        Y => S8487
    );
NOR_3162: ENTITY WORK.NOR
    PORT MAP (
        A => S8341,
        B => S8476,
        Y => S8488
    );
NAND_4893: ENTITY WORK.NAND
    PORT MAP (
        A => S8475,
        B => S8488,
        Y => S8490
    );
NAND_4894: ENTITY WORK.NAND
    PORT MAP (
        A => S8242,
        B => S8291,
        Y => S8491
    );
NOR_3163: ENTITY WORK.NOR
    PORT MAP (
        A => S8490,
        B => S8491,
        Y => S8492
    );
NAND_4895: ENTITY WORK.NAND
    PORT MAP (
        A => S8487,
        B => S8492,
        Y => datapath_shiftunit_2673_A
    );
NOR_3164: ENTITY WORK.NOR
    PORT MAP (
        A => S963,
        B => S8021,
        Y => S8493
    );
NAND_4896: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_6,
        B => S7984,
        Y => S8494
    );
NAND_4897: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_3,
        B => S8006,
        Y => S8495
    );
NAND_4898: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_0,
        B => S8027,
        Y => S8496
    );
NOR_3165: ENTITY WORK.NOR
    PORT MAP (
        A => S1013,
        B => S7981,
        Y => S8497
    );
NAND_4899: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_2,
        B => S7995,
        Y => S8498
    );
NOR_3166: ENTITY WORK.NOR
    PORT MAP (
        A => S1168,
        B => S7992,
        Y => S8500
    );
NOR_3167: ENTITY WORK.NOR
    PORT MAP (
        A => S8106,
        B => S8269,
        Y => S8501
    );
NAND_4900: ENTITY WORK.NAND
    PORT MAP (
        A => S8496,
        B => S8498,
        Y => S8502
    );
NOR_3168: ENTITY WORK.NOR
    PORT MAP (
        A => S8493,
        B => S8502,
        Y => S8503
    );
NAND_4901: ENTITY WORK.NAND
    PORT MAP (
        A => S8034,
        B => S8166,
        Y => S8504
    );
NAND_4902: ENTITY WORK.NAND
    PORT MAP (
        A => S8333,
        B => S8494,
        Y => S8505
    );
NOR_3169: ENTITY WORK.NOR
    PORT MAP (
        A => S8504,
        B => S8505,
        Y => S8506
    );
NAND_4903: ENTITY WORK.NAND
    PORT MAP (
        A => S8503,
        B => S8506,
        Y => S8507
    );
NAND_4904: ENTITY WORK.NAND
    PORT MAP (
        A => S8228,
        B => S8495,
        Y => S8508
    );
NOR_3170: ENTITY WORK.NOR
    PORT MAP (
        A => S8497,
        B => S8508,
        Y => S8509
    );
NAND_4905: ENTITY WORK.NAND
    PORT MAP (
        A => S8310,
        B => S8347,
        Y => S8511
    );
NOR_3171: ENTITY WORK.NOR
    PORT MAP (
        A => S8500,
        B => S8511,
        Y => S8512
    );
NAND_4906: ENTITY WORK.NAND
    PORT MAP (
        A => S8509,
        B => S8512,
        Y => S8513
    );
NOR_3172: ENTITY WORK.NOR
    PORT MAP (
        A => S8507,
        B => S8513,
        Y => S8514
    );
NAND_4907: ENTITY WORK.NAND
    PORT MAP (
        A => S8501,
        B => S8514,
        Y => datapath_shiftunit_2691_A
    );
NAND_4908: ENTITY WORK.NAND
    PORT MAP (
        A => S8281,
        B => S8316,
        Y => S8515
    );
NAND_4909: ENTITY WORK.NAND
    PORT MAP (
        A => S8340,
        B => S8351,
        Y => S8516
    );
NOR_3173: ENTITY WORK.NOR
    PORT MAP (
        A => S8515,
        B => S8516,
        Y => S8517
    );
NAND_4910: ENTITY WORK.NAND
    PORT MAP (
        A => S8070,
        B => S8157,
        Y => S8518
    );
NAND_4911: ENTITY WORK.NAND
    PORT MAP (
        A => S8201,
        B => S8245,
        Y => S8519
    );
NOR_3174: ENTITY WORK.NOR
    PORT MAP (
        A => S8518,
        B => S8519,
        Y => S8521
    );
NAND_4912: ENTITY WORK.NAND
    PORT MAP (
        A => S8517,
        B => S8521,
        Y => S8522
    );
NAND_4913: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_2,
        B => S7993,
        Y => S8523
    );
NAND_4914: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_7,
        B => S7984,
        Y => S8524
    );
NAND_4915: ENTITY WORK.NAND
    PORT MAP (
        A => S8523,
        B => S8524,
        Y => S8525
    );
NAND_4916: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_3,
        B => S7995,
        Y => S8526
    );
NAND_4917: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_1,
        B => S8027,
        Y => S8527
    );
NAND_4918: ENTITY WORK.NAND
    PORT MAP (
        A => S8526,
        B => S8527,
        Y => S8528
    );
NOR_3175: ENTITY WORK.NOR
    PORT MAP (
        A => S8525,
        B => S8528,
        Y => S8529
    );
NAND_4919: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_6,
        B => S8020,
        Y => S8530
    );
NAND_4920: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_4,
        B => S8006,
        Y => S8532
    );
NAND_4921: ENTITY WORK.NAND
    PORT MAP (
        A => S8530,
        B => S8532,
        Y => S8533
    );
NOR_3176: ENTITY WORK.NOR
    PORT MAP (
        A => S963,
        B => S7981,
        Y => S8534
    );
NOT_554: ENTITY WORK.NOT
    PORT MAP (
        A => S8534,
        Y => S8535
    );
NAND_4922: ENTITY WORK.NAND
    PORT MAP (
        A => datapath_addsubunit_in1_0,
        B => S8035,
        Y => S8536
    );
NAND_4923: ENTITY WORK.NAND
    PORT MAP (
        A => S8535,
        B => S8536,
        Y => S8537
    );
NOR_3177: ENTITY WORK.NOR
    PORT MAP (
        A => S8533,
        B => S8537,
        Y => S8538
    );
NAND_4924: ENTITY WORK.NAND
    PORT MAP (
        A => S8529,
        B => S8538,
        Y => S8539
    );
NOR_3178: ENTITY WORK.NOR
    PORT MAP (
        A => S8522,
        B => S8539,
        Y => S8540
    );
NOT_555: ENTITY WORK.NOT
    PORT MAP (
        A => S8540,
        Y => datapath_shiftunit_2708_A
    );
BUF_1: ENTITY WORK.BUF
    PORT MAP (
        A => datapath_theregisterfile_memtrf_240,
        Y => S244
    );
BUF_2: ENTITY WORK.BUF
    PORT MAP (
        A => datapath_theregisterfile_memtrf_241,
        Y => S245
    );
BUF_3: ENTITY WORK.BUF
    PORT MAP (
        A => datapath_theregisterfile_memtrf_242,
        Y => S246
    );
BUF_4: ENTITY WORK.BUF
    PORT MAP (
        A => datapath_theregisterfile_memtrf_243,
        Y => S247
    );
BUF_5: ENTITY WORK.BUF
    PORT MAP (
        A => datapath_theregisterfile_memtrf_244,
        Y => S248
    );
BUF_6: ENTITY WORK.BUF
    PORT MAP (
        A => datapath_theregisterfile_memtrf_245,
        Y => S249
    );
BUF_7: ENTITY WORK.BUF
    PORT MAP (
        A => datapath_theregisterfile_memtrf_246,
        Y => S250
    );
BUF_8: ENTITY WORK.BUF
    PORT MAP (
        A => datapath_theregisterfile_memtrf_247,
        Y => S251
    );
BUF_9: ENTITY WORK.BUF
    PORT MAP (
        A => datapath_theregisterfile_memtrf_248,
        Y => S252
    );
BUF_10: ENTITY WORK.BUF
    PORT MAP (
        A => datapath_theregisterfile_memtrf_249,
        Y => S253
    );
BUF_11: ENTITY WORK.BUF
    PORT MAP (
        A => datapath_theregisterfile_memtrf_250,
        Y => S254
    );
BUF_12: ENTITY WORK.BUF
    PORT MAP (
        A => datapath_theregisterfile_memtrf_251,
        Y => S255
    );
BUF_13: ENTITY WORK.BUF
    PORT MAP (
        A => datapath_theregisterfile_memtrf_252,
        Y => S256
    );
BUF_14: ENTITY WORK.BUF
    PORT MAP (
        A => datapath_theregisterfile_memtrf_253,
        Y => S257
    );
BUF_15: ENTITY WORK.BUF
    PORT MAP (
        A => datapath_theregisterfile_memtrf_254,
        Y => S258
    );
BUF_16: ENTITY WORK.BUF
    PORT MAP (
        A => datapath_theregisterfile_memtrf_255,
        Y => S259
    );
BUF_17: ENTITY WORK.BUF
    PORT MAP (
        A => controller_outflag_0,
        Y => S260
    );
BUF_18: ENTITY WORK.BUF
    PORT MAP (
        A => controller_outflag_1,
        Y => S261
    );
BUF_19: ENTITY WORK.BUF
    PORT MAP (
        A => controller_outflag_2,
        Y => S262
    );
BUF_20: ENTITY WORK.BUF
    PORT MAP (
        A => controller_outflag_3,
        Y => S263
    );
BUF_21: ENTITY WORK.BUF
    PORT MAP (
        A => controller_outflag_6,
        Y => S266
    );
BUF_22: ENTITY WORK.BUF
    PORT MAP (
        A => controller_outflag_7,
        Y => S343
    );
DFF_PP0_1: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => controller_1405_Y_0,
        Q => controller_pstate_0,
        R => controller_rst
    );
DFF_PP0_2: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => controller_1405_Y_1,
        Q => controller_pstate_1,
        R => controller_rst
    );
DFF_PP0_3: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S328,
        Q => datapath_adr_outreg_0,
        R => controller_rst
    );
DFF_PP0_4: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S329,
        Q => datapath_adr_outreg_1,
        R => controller_rst
    );
DFF_PP0_5: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S330,
        Q => datapath_adr_outreg_2,
        R => controller_rst
    );
DFF_PP0_6: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S331,
        Q => datapath_adr_outreg_3,
        R => controller_rst
    );
DFF_PP0_7: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S332,
        Q => datapath_adr_outreg_4,
        R => controller_rst
    );
DFF_PP0_8: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S333,
        Q => datapath_adr_outreg_5,
        R => controller_rst
    );
DFF_PP0_9: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S334,
        Q => datapath_adr_outreg_6,
        R => controller_rst
    );
DFF_PP0_10: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S335,
        Q => datapath_adr_outreg_7,
        R => controller_rst
    );
DFF_PP0_11: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S336,
        Q => datapath_adr_outreg_8,
        R => controller_rst
    );
DFF_PP0_12: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S337,
        Q => datapath_adr_outreg_9,
        R => controller_rst
    );
DFF_PP0_13: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S338,
        Q => datapath_adr_outreg_10,
        R => controller_rst
    );
DFF_PP0_14: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S339,
        Q => datapath_adr_outreg_11,
        R => controller_rst
    );
DFF_PP0_15: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S340,
        Q => datapath_adr_outreg_12,
        R => controller_rst
    );
DFF_PP0_16: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S341,
        Q => datapath_adr_outreg_13,
        R => controller_rst
    );
DFF_PP0_17: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S342,
        Q => datapath_adr_outreg_14,
        R => controller_rst
    );
DFF_PP0_18: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S3,
        Q => datapath_adr_outreg_15,
        R => controller_rst
    );
DFF_PP0_19: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S313,
        Q => datapath_instruction_0,
        R => controller_rst
    );
DFF_PP0_20: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S314,
        Q => datapath_instruction_1,
        R => controller_rst
    );
DFF_PP0_21: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S315,
        Q => datapath_instruction_2,
        R => controller_rst
    );
DFF_PP0_22: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S316,
        Q => datapath_instruction_3,
        R => controller_rst
    );
DFF_PP0_23: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S317,
        Q => controller_fib_0,
        R => controller_rst
    );
DFF_PP0_24: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S318,
        Q => controller_fib_1,
        R => controller_rst
    );
DFF_PP0_25: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S319,
        Q => controller_fib_2,
        R => controller_rst
    );
DFF_PP0_26: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S320,
        Q => controller_fib_3,
        R => controller_rst
    );
DFF_PP0_27: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S321,
        Q => controller_fib_4,
        R => controller_rst
    );
DFF_PP0_28: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S322,
        Q => controller_216_B_0,
        R => controller_rst
    );
DFF_PP0_29: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S323,
        Q => controller_opcode_2,
        R => controller_rst
    );
DFF_PP0_30: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S324,
        Q => controller_opcode_3,
        R => controller_rst
    );
DFF_PP0_31: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S325,
        Q => controller_opcode_4,
        R => controller_rst
    );
DFF_PP0_32: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S326,
        Q => controller_opcode_5,
        R => controller_rst
    );
DFF_PP0_33: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S327,
        Q => controller_opcode_6,
        R => controller_rst
    );
DFF_PP0_34: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S2,
        Q => controller_opcode_7,
        R => controller_rst
    );
DFF_PP0_35: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S282,
        Q => datapath_multdivunit_outmdu1_0,
        R => controller_rst
    );
DFF_PP0_36: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S283,
        Q => datapath_multdivunit_outmdu1_1,
        R => controller_rst
    );
DFF_PP0_37: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S284,
        Q => datapath_multdivunit_outmdu1_2,
        R => controller_rst
    );
DFF_PP0_38: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S285,
        Q => datapath_multdivunit_outmdu1_3,
        R => controller_rst
    );
DFF_PP0_39: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S286,
        Q => datapath_multdivunit_outmdu1_4,
        R => controller_rst
    );
DFF_PP0_40: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S287,
        Q => datapath_multdivunit_outmdu1_5,
        R => controller_rst
    );
DFF_PP0_41: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S288,
        Q => datapath_multdivunit_outmdu1_6,
        R => controller_rst
    );
DFF_PP0_42: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S289,
        Q => datapath_multdivunit_outmdu1_7,
        R => controller_rst
    );
DFF_PP0_43: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S290,
        Q => datapath_multdivunit_outmdu1_8,
        R => controller_rst
    );
DFF_PP0_44: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S291,
        Q => datapath_multdivunit_outmdu1_9,
        R => controller_rst
    );
DFF_PP0_45: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S292,
        Q => datapath_multdivunit_outmdu1_10,
        R => controller_rst
    );
DFF_PP0_46: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S293,
        Q => datapath_multdivunit_outmdu1_11,
        R => controller_rst
    );
DFF_PP0_47: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S294,
        Q => datapath_multdivunit_outmdu1_12,
        R => controller_rst
    );
DFF_PP0_48: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S295,
        Q => datapath_multdivunit_outmdu1_13,
        R => controller_rst
    );
DFF_PP0_49: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S296,
        Q => datapath_multdivunit_outmdu1_14,
        R => controller_rst
    );
DFF_PP0_50: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S297,
        Q => datapath_multdivunit_outmdu1_15,
        R => controller_rst
    );
DFF_PP0_51: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S298,
        Q => datapath_multdivunit_outmdu2_0,
        R => controller_rst
    );
DFF_PP0_52: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S299,
        Q => datapath_multdivunit_outmdu2_1,
        R => controller_rst
    );
DFF_PP0_53: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S300,
        Q => datapath_multdivunit_outmdu2_2,
        R => controller_rst
    );
DFF_PP0_54: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S301,
        Q => datapath_multdivunit_outmdu2_3,
        R => controller_rst
    );
DFF_PP0_55: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S302,
        Q => datapath_multdivunit_outmdu2_4,
        R => controller_rst
    );
DFF_PP0_56: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S303,
        Q => datapath_multdivunit_outmdu2_5,
        R => controller_rst
    );
DFF_PP0_57: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S304,
        Q => datapath_multdivunit_outmdu2_6,
        R => controller_rst
    );
DFF_PP0_58: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S305,
        Q => datapath_multdivunit_outmdu2_7,
        R => controller_rst
    );
DFF_PP0_59: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S306,
        Q => datapath_multdivunit_outmdu2_8,
        R => controller_rst
    );
DFF_PP0_60: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S307,
        Q => datapath_multdivunit_outmdu2_9,
        R => controller_rst
    );
DFF_PP0_61: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S308,
        Q => datapath_multdivunit_outmdu2_10,
        R => controller_rst
    );
DFF_PP0_62: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S309,
        Q => datapath_multdivunit_outmdu2_11,
        R => controller_rst
    );
DFF_PP0_63: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S310,
        Q => datapath_multdivunit_outmdu2_12,
        R => controller_rst
    );
DFF_PP0_64: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S311,
        Q => datapath_multdivunit_outmdu2_13,
        R => controller_rst
    );
DFF_PP0_65: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S312,
        Q => datapath_multdivunit_outmdu2_14,
        R => controller_rst
    );
DFF_PP0_66: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S1,
        Q => datapath_multdivunit_outmdu2_15,
        R => controller_rst
    );
DFF_PP0_67: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S267,
        Q => datapath_muxmem_in2_0,
        R => controller_rst
    );
DFF_PP0_68: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S268,
        Q => datapath_muxmem_in2_1,
        R => controller_rst
    );
DFF_PP0_69: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S269,
        Q => datapath_muxmem_in2_2,
        R => controller_rst
    );
DFF_PP0_70: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S270,
        Q => datapath_muxmem_in2_3,
        R => controller_rst
    );
DFF_PP0_71: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S271,
        Q => datapath_muxmem_in2_4,
        R => controller_rst
    );
DFF_PP0_72: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S272,
        Q => datapath_muxmem_in2_5,
        R => controller_rst
    );
DFF_PP0_73: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S273,
        Q => datapath_muxmem_in2_6,
        R => controller_rst
    );
DFF_PP0_74: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S274,
        Q => datapath_muxmem_in2_7,
        R => controller_rst
    );
DFF_PP0_75: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S275,
        Q => datapath_muxmem_in2_8,
        R => controller_rst
    );
DFF_PP0_76: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S276,
        Q => datapath_muxmem_in2_9,
        R => controller_rst
    );
DFF_PP0_77: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S277,
        Q => datapath_muxmem_in2_10,
        R => controller_rst
    );
DFF_PP0_78: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S278,
        Q => datapath_muxmem_in2_11,
        R => controller_rst
    );
DFF_PP0_79: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S279,
        Q => datapath_muxmem_in2_12,
        R => controller_rst
    );
DFF_PP0_80: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S280,
        Q => datapath_muxmem_in2_13,
        R => controller_rst
    );
DFF_PP0_81: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S281,
        Q => datapath_muxmem_in2_14,
        R => controller_rst
    );
DFF_PP0_82: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S0,
        Q => datapath_muxmem_in2_15,
        R => controller_rst
    );
DFF_NP1_1: ENTITY WORK.DFF_NP1
    PORT MAP (
        C => controller_clk,
        D => S4,
        Q => datapath_theregisterfile_memtrf_64,
        R => controller_rst
    );
DFF_NP1_2: ENTITY WORK.DFF_NP1
    PORT MAP (
        C => controller_clk,
        D => S5,
        Q => datapath_theregisterfile_memtrf_65,
        R => controller_rst
    );
DFF_NP0_1: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S6,
        Q => datapath_theregisterfile_memtrf_66,
        R => controller_rst
    );
DFF_NP1_3: ENTITY WORK.DFF_NP1
    PORT MAP (
        C => controller_clk,
        D => S7,
        Q => datapath_theregisterfile_memtrf_67,
        R => controller_rst
    );
DFF_NP0_2: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S8,
        Q => datapath_theregisterfile_memtrf_68,
        R => controller_rst
    );
DFF_NP0_3: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S9,
        Q => datapath_theregisterfile_memtrf_69,
        R => controller_rst
    );
DFF_NP0_4: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S10,
        Q => datapath_theregisterfile_memtrf_70,
        R => controller_rst
    );
DFF_NP0_5: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S11,
        Q => datapath_theregisterfile_memtrf_71,
        R => controller_rst
    );
DFF_NP0_6: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S12,
        Q => datapath_theregisterfile_memtrf_72,
        R => controller_rst
    );
DFF_NP0_7: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S13,
        Q => datapath_theregisterfile_memtrf_73,
        R => controller_rst
    );
DFF_NP0_8: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S14,
        Q => datapath_theregisterfile_memtrf_74,
        R => controller_rst
    );
DFF_NP0_9: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S15,
        Q => datapath_theregisterfile_memtrf_75,
        R => controller_rst
    );
DFF_NP0_10: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S16,
        Q => datapath_theregisterfile_memtrf_76,
        R => controller_rst
    );
DFF_NP0_11: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S17,
        Q => datapath_theregisterfile_memtrf_77,
        R => controller_rst
    );
DFF_NP0_12: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S18,
        Q => datapath_theregisterfile_memtrf_78,
        R => controller_rst
    );
DFF_NP0_13: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S19,
        Q => datapath_theregisterfile_memtrf_79,
        R => controller_rst
    );
DFF_NP1_4: ENTITY WORK.DFF_NP1
    PORT MAP (
        C => controller_clk,
        D => S20,
        Q => datapath_theregisterfile_memtrf_32,
        R => controller_rst
    );
DFF_NP0_14: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S21,
        Q => datapath_theregisterfile_memtrf_33,
        R => controller_rst
    );
DFF_NP1_5: ENTITY WORK.DFF_NP1
    PORT MAP (
        C => controller_clk,
        D => S22,
        Q => datapath_theregisterfile_memtrf_34,
        R => controller_rst
    );
DFF_NP1_6: ENTITY WORK.DFF_NP1
    PORT MAP (
        C => controller_clk,
        D => S23,
        Q => datapath_theregisterfile_memtrf_35,
        R => controller_rst
    );
DFF_NP0_15: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S24,
        Q => datapath_theregisterfile_memtrf_36,
        R => controller_rst
    );
DFF_NP0_16: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S25,
        Q => datapath_theregisterfile_memtrf_37,
        R => controller_rst
    );
DFF_NP0_17: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S26,
        Q => datapath_theregisterfile_memtrf_38,
        R => controller_rst
    );
DFF_NP0_18: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S27,
        Q => datapath_theregisterfile_memtrf_39,
        R => controller_rst
    );
DFF_NP0_19: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S28,
        Q => datapath_theregisterfile_memtrf_40,
        R => controller_rst
    );
DFF_NP0_20: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S29,
        Q => datapath_theregisterfile_memtrf_41,
        R => controller_rst
    );
DFF_NP0_21: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S30,
        Q => datapath_theregisterfile_memtrf_42,
        R => controller_rst
    );
DFF_NP0_22: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S31,
        Q => datapath_theregisterfile_memtrf_43,
        R => controller_rst
    );
DFF_NP0_23: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S32,
        Q => datapath_theregisterfile_memtrf_44,
        R => controller_rst
    );
DFF_NP0_24: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S33,
        Q => datapath_theregisterfile_memtrf_45,
        R => controller_rst
    );
DFF_NP0_25: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S34,
        Q => datapath_theregisterfile_memtrf_46,
        R => controller_rst
    );
DFF_NP0_26: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S35,
        Q => datapath_theregisterfile_memtrf_47,
        R => controller_rst
    );
DFF_NP0_27: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S36,
        Q => datapath_theregisterfile_memtrf_48,
        R => controller_rst
    );
DFF_NP0_28: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S37,
        Q => datapath_theregisterfile_memtrf_49,
        R => controller_rst
    );
DFF_NP1_7: ENTITY WORK.DFF_NP1
    PORT MAP (
        C => controller_clk,
        D => S38,
        Q => datapath_theregisterfile_memtrf_50,
        R => controller_rst
    );
DFF_NP1_8: ENTITY WORK.DFF_NP1
    PORT MAP (
        C => controller_clk,
        D => S39,
        Q => datapath_theregisterfile_memtrf_51,
        R => controller_rst
    );
DFF_NP0_29: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S40,
        Q => datapath_theregisterfile_memtrf_52,
        R => controller_rst
    );
DFF_NP0_30: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S41,
        Q => datapath_theregisterfile_memtrf_53,
        R => controller_rst
    );
DFF_NP0_31: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S42,
        Q => datapath_theregisterfile_memtrf_54,
        R => controller_rst
    );
DFF_NP0_32: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S43,
        Q => datapath_theregisterfile_memtrf_55,
        R => controller_rst
    );
DFF_NP0_33: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S44,
        Q => datapath_theregisterfile_memtrf_56,
        R => controller_rst
    );
DFF_NP0_34: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S45,
        Q => datapath_theregisterfile_memtrf_57,
        R => controller_rst
    );
DFF_NP0_35: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S46,
        Q => datapath_theregisterfile_memtrf_58,
        R => controller_rst
    );
DFF_NP0_36: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S47,
        Q => datapath_theregisterfile_memtrf_59,
        R => controller_rst
    );
DFF_NP0_37: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S48,
        Q => datapath_theregisterfile_memtrf_60,
        R => controller_rst
    );
DFF_NP0_38: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S49,
        Q => datapath_theregisterfile_memtrf_61,
        R => controller_rst
    );
DFF_NP0_39: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S50,
        Q => datapath_theregisterfile_memtrf_62,
        R => controller_rst
    );
DFF_NP0_40: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S51,
        Q => datapath_theregisterfile_memtrf_63,
        R => controller_rst
    );
DFF_NP1_9: ENTITY WORK.DFF_NP1
    PORT MAP (
        C => controller_clk,
        D => S52,
        Q => datapath_theregisterfile_memtrf_128,
        R => controller_rst
    );
DFF_NP1_10: ENTITY WORK.DFF_NP1
    PORT MAP (
        C => controller_clk,
        D => S53,
        Q => datapath_theregisterfile_memtrf_129,
        R => controller_rst
    );
DFF_NP1_11: ENTITY WORK.DFF_NP1
    PORT MAP (
        C => controller_clk,
        D => S54,
        Q => datapath_theregisterfile_memtrf_130,
        R => controller_rst
    );
DFF_NP0_41: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S55,
        Q => datapath_theregisterfile_memtrf_131,
        R => controller_rst
    );
DFF_NP0_42: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S56,
        Q => datapath_theregisterfile_memtrf_132,
        R => controller_rst
    );
DFF_NP0_43: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S57,
        Q => datapath_theregisterfile_memtrf_133,
        R => controller_rst
    );
DFF_NP0_44: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S58,
        Q => datapath_theregisterfile_memtrf_134,
        R => controller_rst
    );
DFF_NP0_45: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S59,
        Q => datapath_theregisterfile_memtrf_135,
        R => controller_rst
    );
DFF_NP0_46: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S60,
        Q => datapath_theregisterfile_memtrf_136,
        R => controller_rst
    );
DFF_NP0_47: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S61,
        Q => datapath_theregisterfile_memtrf_137,
        R => controller_rst
    );
DFF_NP0_48: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S62,
        Q => datapath_theregisterfile_memtrf_138,
        R => controller_rst
    );
DFF_NP0_49: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S63,
        Q => datapath_theregisterfile_memtrf_139,
        R => controller_rst
    );
DFF_NP0_50: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S64,
        Q => datapath_theregisterfile_memtrf_140,
        R => controller_rst
    );
DFF_NP0_51: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S65,
        Q => datapath_theregisterfile_memtrf_141,
        R => controller_rst
    );
DFF_NP0_52: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S66,
        Q => datapath_theregisterfile_memtrf_142,
        R => controller_rst
    );
DFF_NP0_53: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S67,
        Q => datapath_theregisterfile_memtrf_143,
        R => controller_rst
    );
DFF_NP0_54: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S68,
        Q => datapath_theregisterfile_memtrf_16,
        R => controller_rst
    );
DFF_NP1_12: ENTITY WORK.DFF_NP1
    PORT MAP (
        C => controller_clk,
        D => S69,
        Q => datapath_theregisterfile_memtrf_17,
        R => controller_rst
    );
DFF_NP1_13: ENTITY WORK.DFF_NP1
    PORT MAP (
        C => controller_clk,
        D => S70,
        Q => datapath_theregisterfile_memtrf_18,
        R => controller_rst
    );
DFF_NP1_14: ENTITY WORK.DFF_NP1
    PORT MAP (
        C => controller_clk,
        D => S71,
        Q => datapath_theregisterfile_memtrf_19,
        R => controller_rst
    );
DFF_NP0_55: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S72,
        Q => datapath_theregisterfile_memtrf_20,
        R => controller_rst
    );
DFF_NP0_56: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S73,
        Q => datapath_theregisterfile_memtrf_21,
        R => controller_rst
    );
DFF_NP0_57: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S74,
        Q => datapath_theregisterfile_memtrf_22,
        R => controller_rst
    );
DFF_NP0_58: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S75,
        Q => datapath_theregisterfile_memtrf_23,
        R => controller_rst
    );
DFF_NP0_59: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S76,
        Q => datapath_theregisterfile_memtrf_24,
        R => controller_rst
    );
DFF_NP0_60: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S77,
        Q => datapath_theregisterfile_memtrf_25,
        R => controller_rst
    );
DFF_NP0_61: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S78,
        Q => datapath_theregisterfile_memtrf_26,
        R => controller_rst
    );
DFF_NP0_62: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S79,
        Q => datapath_theregisterfile_memtrf_27,
        R => controller_rst
    );
DFF_NP0_63: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S80,
        Q => datapath_theregisterfile_memtrf_28,
        R => controller_rst
    );
DFF_NP0_64: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S81,
        Q => datapath_theregisterfile_memtrf_29,
        R => controller_rst
    );
DFF_NP0_65: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S82,
        Q => datapath_theregisterfile_memtrf_30,
        R => controller_rst
    );
DFF_NP0_66: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S83,
        Q => datapath_theregisterfile_memtrf_31,
        R => controller_rst
    );
DFF_NP0_67: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S84,
        Q => datapath_theregisterfile_memtrf_80,
        R => controller_rst
    );
DFF_NP1_15: ENTITY WORK.DFF_NP1
    PORT MAP (
        C => controller_clk,
        D => S85,
        Q => datapath_theregisterfile_memtrf_81,
        R => controller_rst
    );
DFF_NP0_68: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S86,
        Q => datapath_theregisterfile_memtrf_82,
        R => controller_rst
    );
DFF_NP1_16: ENTITY WORK.DFF_NP1
    PORT MAP (
        C => controller_clk,
        D => S87,
        Q => datapath_theregisterfile_memtrf_83,
        R => controller_rst
    );
DFF_NP0_69: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S88,
        Q => datapath_theregisterfile_memtrf_84,
        R => controller_rst
    );
DFF_NP0_70: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S89,
        Q => datapath_theregisterfile_memtrf_85,
        R => controller_rst
    );
DFF_NP0_71: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S90,
        Q => datapath_theregisterfile_memtrf_86,
        R => controller_rst
    );
DFF_NP0_72: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S91,
        Q => datapath_theregisterfile_memtrf_87,
        R => controller_rst
    );
DFF_NP0_73: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S92,
        Q => datapath_theregisterfile_memtrf_88,
        R => controller_rst
    );
DFF_NP0_74: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S93,
        Q => datapath_theregisterfile_memtrf_89,
        R => controller_rst
    );
DFF_NP0_75: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S94,
        Q => datapath_theregisterfile_memtrf_90,
        R => controller_rst
    );
DFF_NP0_76: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S95,
        Q => datapath_theregisterfile_memtrf_91,
        R => controller_rst
    );
DFF_NP0_77: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S96,
        Q => datapath_theregisterfile_memtrf_92,
        R => controller_rst
    );
DFF_NP0_78: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S97,
        Q => datapath_theregisterfile_memtrf_93,
        R => controller_rst
    );
DFF_NP0_79: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S98,
        Q => datapath_theregisterfile_memtrf_94,
        R => controller_rst
    );
DFF_NP0_80: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S99,
        Q => datapath_theregisterfile_memtrf_95,
        R => controller_rst
    );
DFF_NP1_17: ENTITY WORK.DFF_NP1
    PORT MAP (
        C => controller_clk,
        D => S100,
        Q => datapath_theregisterfile_memtrf_96,
        R => controller_rst
    );
DFF_NP0_81: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S101,
        Q => datapath_theregisterfile_memtrf_97,
        R => controller_rst
    );
DFF_NP0_82: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S102,
        Q => datapath_theregisterfile_memtrf_98,
        R => controller_rst
    );
DFF_NP1_18: ENTITY WORK.DFF_NP1
    PORT MAP (
        C => controller_clk,
        D => S103,
        Q => datapath_theregisterfile_memtrf_99,
        R => controller_rst
    );
DFF_NP0_83: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S104,
        Q => datapath_theregisterfile_memtrf_100,
        R => controller_rst
    );
DFF_NP0_84: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S105,
        Q => datapath_theregisterfile_memtrf_101,
        R => controller_rst
    );
DFF_NP0_85: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S106,
        Q => datapath_theregisterfile_memtrf_102,
        R => controller_rst
    );
DFF_NP0_86: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S107,
        Q => datapath_theregisterfile_memtrf_103,
        R => controller_rst
    );
DFF_NP0_87: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S108,
        Q => datapath_theregisterfile_memtrf_104,
        R => controller_rst
    );
DFF_NP0_88: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S109,
        Q => datapath_theregisterfile_memtrf_105,
        R => controller_rst
    );
DFF_NP0_89: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S110,
        Q => datapath_theregisterfile_memtrf_106,
        R => controller_rst
    );
DFF_NP0_90: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S111,
        Q => datapath_theregisterfile_memtrf_107,
        R => controller_rst
    );
DFF_NP0_91: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S112,
        Q => datapath_theregisterfile_memtrf_108,
        R => controller_rst
    );
DFF_NP0_92: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S113,
        Q => datapath_theregisterfile_memtrf_109,
        R => controller_rst
    );
DFF_NP0_93: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S114,
        Q => datapath_theregisterfile_memtrf_110,
        R => controller_rst
    );
DFF_NP0_94: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S115,
        Q => datapath_theregisterfile_memtrf_111,
        R => controller_rst
    );
DFF_NP0_95: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S116,
        Q => datapath_theregisterfile_memtrf_112,
        R => controller_rst
    );
DFF_NP0_96: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S117,
        Q => datapath_theregisterfile_memtrf_113,
        R => controller_rst
    );
DFF_NP0_97: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S118,
        Q => datapath_theregisterfile_memtrf_114,
        R => controller_rst
    );
DFF_NP1_19: ENTITY WORK.DFF_NP1
    PORT MAP (
        C => controller_clk,
        D => S119,
        Q => datapath_theregisterfile_memtrf_115,
        R => controller_rst
    );
DFF_NP0_98: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S120,
        Q => datapath_theregisterfile_memtrf_116,
        R => controller_rst
    );
DFF_NP0_99: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S121,
        Q => datapath_theregisterfile_memtrf_117,
        R => controller_rst
    );
DFF_NP0_100: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S122,
        Q => datapath_theregisterfile_memtrf_118,
        R => controller_rst
    );
DFF_NP0_101: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S123,
        Q => datapath_theregisterfile_memtrf_119,
        R => controller_rst
    );
DFF_NP0_102: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S124,
        Q => datapath_theregisterfile_memtrf_120,
        R => controller_rst
    );
DFF_NP0_103: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S125,
        Q => datapath_theregisterfile_memtrf_121,
        R => controller_rst
    );
DFF_NP0_104: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S126,
        Q => datapath_theregisterfile_memtrf_122,
        R => controller_rst
    );
DFF_NP0_105: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S127,
        Q => datapath_theregisterfile_memtrf_123,
        R => controller_rst
    );
DFF_NP0_106: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S128,
        Q => datapath_theregisterfile_memtrf_124,
        R => controller_rst
    );
DFF_NP0_107: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S129,
        Q => datapath_theregisterfile_memtrf_125,
        R => controller_rst
    );
DFF_NP0_108: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S130,
        Q => datapath_theregisterfile_memtrf_126,
        R => controller_rst
    );
DFF_NP0_109: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S131,
        Q => datapath_theregisterfile_memtrf_127,
        R => controller_rst
    );
DFF_NP1_20: ENTITY WORK.DFF_NP1
    PORT MAP (
        C => controller_clk,
        D => S132,
        Q => datapath_theregisterfile_memtrf_0,
        R => controller_rst
    );
DFF_NP1_21: ENTITY WORK.DFF_NP1
    PORT MAP (
        C => controller_clk,
        D => S133,
        Q => datapath_theregisterfile_memtrf_1,
        R => controller_rst
    );
DFF_NP1_22: ENTITY WORK.DFF_NP1
    PORT MAP (
        C => controller_clk,
        D => S134,
        Q => datapath_theregisterfile_memtrf_2,
        R => controller_rst
    );
DFF_NP1_23: ENTITY WORK.DFF_NP1
    PORT MAP (
        C => controller_clk,
        D => S135,
        Q => datapath_theregisterfile_memtrf_3,
        R => controller_rst
    );
DFF_NP0_110: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S136,
        Q => datapath_theregisterfile_memtrf_4,
        R => controller_rst
    );
DFF_NP0_111: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S137,
        Q => datapath_theregisterfile_memtrf_5,
        R => controller_rst
    );
DFF_NP0_112: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S138,
        Q => datapath_theregisterfile_memtrf_6,
        R => controller_rst
    );
DFF_NP0_113: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S139,
        Q => datapath_theregisterfile_memtrf_7,
        R => controller_rst
    );
DFF_NP0_114: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S140,
        Q => datapath_theregisterfile_memtrf_8,
        R => controller_rst
    );
DFF_NP0_115: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S141,
        Q => datapath_theregisterfile_memtrf_9,
        R => controller_rst
    );
DFF_NP0_116: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S142,
        Q => datapath_theregisterfile_memtrf_10,
        R => controller_rst
    );
DFF_NP0_117: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S143,
        Q => datapath_theregisterfile_memtrf_11,
        R => controller_rst
    );
DFF_NP0_118: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S144,
        Q => datapath_theregisterfile_memtrf_12,
        R => controller_rst
    );
DFF_NP0_119: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S145,
        Q => datapath_theregisterfile_memtrf_13,
        R => controller_rst
    );
DFF_NP0_120: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S146,
        Q => datapath_theregisterfile_memtrf_14,
        R => controller_rst
    );
DFF_NP0_121: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S147,
        Q => datapath_theregisterfile_memtrf_15,
        R => controller_rst
    );
DFF_NP0_122: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S148,
        Q => datapath_theregisterfile_memtrf_144,
        R => controller_rst
    );
DFF_NP1_24: ENTITY WORK.DFF_NP1
    PORT MAP (
        C => controller_clk,
        D => S149,
        Q => datapath_theregisterfile_memtrf_145,
        R => controller_rst
    );
DFF_NP1_25: ENTITY WORK.DFF_NP1
    PORT MAP (
        C => controller_clk,
        D => S150,
        Q => datapath_theregisterfile_memtrf_146,
        R => controller_rst
    );
DFF_NP0_123: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S151,
        Q => datapath_theregisterfile_memtrf_147,
        R => controller_rst
    );
DFF_NP0_124: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S152,
        Q => datapath_theregisterfile_memtrf_148,
        R => controller_rst
    );
DFF_NP0_125: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S153,
        Q => datapath_theregisterfile_memtrf_149,
        R => controller_rst
    );
DFF_NP0_126: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S154,
        Q => datapath_theregisterfile_memtrf_150,
        R => controller_rst
    );
DFF_NP0_127: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S155,
        Q => datapath_theregisterfile_memtrf_151,
        R => controller_rst
    );
DFF_NP0_128: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S156,
        Q => datapath_theregisterfile_memtrf_152,
        R => controller_rst
    );
DFF_NP0_129: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S157,
        Q => datapath_theregisterfile_memtrf_153,
        R => controller_rst
    );
DFF_NP0_130: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S158,
        Q => datapath_theregisterfile_memtrf_154,
        R => controller_rst
    );
DFF_NP0_131: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S159,
        Q => datapath_theregisterfile_memtrf_155,
        R => controller_rst
    );
DFF_NP0_132: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S160,
        Q => datapath_theregisterfile_memtrf_156,
        R => controller_rst
    );
DFF_NP0_133: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S161,
        Q => datapath_theregisterfile_memtrf_157,
        R => controller_rst
    );
DFF_NP0_134: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S162,
        Q => datapath_theregisterfile_memtrf_158,
        R => controller_rst
    );
DFF_NP0_135: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S163,
        Q => datapath_theregisterfile_memtrf_159,
        R => controller_rst
    );
DFF_NP1_26: ENTITY WORK.DFF_NP1
    PORT MAP (
        C => controller_clk,
        D => S164,
        Q => datapath_theregisterfile_memtrf_160,
        R => controller_rst
    );
DFF_NP0_136: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S165,
        Q => datapath_theregisterfile_memtrf_161,
        R => controller_rst
    );
DFF_NP1_27: ENTITY WORK.DFF_NP1
    PORT MAP (
        C => controller_clk,
        D => S166,
        Q => datapath_theregisterfile_memtrf_162,
        R => controller_rst
    );
DFF_NP0_137: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S167,
        Q => datapath_theregisterfile_memtrf_163,
        R => controller_rst
    );
DFF_NP0_138: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S168,
        Q => datapath_theregisterfile_memtrf_164,
        R => controller_rst
    );
DFF_NP0_139: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S169,
        Q => datapath_theregisterfile_memtrf_165,
        R => controller_rst
    );
DFF_NP0_140: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S170,
        Q => datapath_theregisterfile_memtrf_166,
        R => controller_rst
    );
DFF_NP0_141: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S171,
        Q => datapath_theregisterfile_memtrf_167,
        R => controller_rst
    );
DFF_NP0_142: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S172,
        Q => datapath_theregisterfile_memtrf_168,
        R => controller_rst
    );
DFF_NP0_143: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S173,
        Q => datapath_theregisterfile_memtrf_169,
        R => controller_rst
    );
DFF_NP0_144: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S174,
        Q => datapath_theregisterfile_memtrf_170,
        R => controller_rst
    );
DFF_NP0_145: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S175,
        Q => datapath_theregisterfile_memtrf_171,
        R => controller_rst
    );
DFF_NP0_146: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S176,
        Q => datapath_theregisterfile_memtrf_172,
        R => controller_rst
    );
DFF_NP0_147: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S177,
        Q => datapath_theregisterfile_memtrf_173,
        R => controller_rst
    );
DFF_NP0_148: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S178,
        Q => datapath_theregisterfile_memtrf_174,
        R => controller_rst
    );
DFF_NP0_149: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S179,
        Q => datapath_theregisterfile_memtrf_175,
        R => controller_rst
    );
DFF_NP0_150: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S180,
        Q => datapath_theregisterfile_memtrf_176,
        R => controller_rst
    );
DFF_NP0_151: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S181,
        Q => datapath_theregisterfile_memtrf_177,
        R => controller_rst
    );
DFF_NP1_28: ENTITY WORK.DFF_NP1
    PORT MAP (
        C => controller_clk,
        D => S182,
        Q => datapath_theregisterfile_memtrf_178,
        R => controller_rst
    );
DFF_NP0_152: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S183,
        Q => datapath_theregisterfile_memtrf_179,
        R => controller_rst
    );
DFF_NP0_153: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S184,
        Q => datapath_theregisterfile_memtrf_180,
        R => controller_rst
    );
DFF_NP0_154: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S185,
        Q => datapath_theregisterfile_memtrf_181,
        R => controller_rst
    );
DFF_NP0_155: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S186,
        Q => datapath_theregisterfile_memtrf_182,
        R => controller_rst
    );
DFF_NP0_156: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S187,
        Q => datapath_theregisterfile_memtrf_183,
        R => controller_rst
    );
DFF_NP0_157: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S188,
        Q => datapath_theregisterfile_memtrf_184,
        R => controller_rst
    );
DFF_NP0_158: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S189,
        Q => datapath_theregisterfile_memtrf_185,
        R => controller_rst
    );
DFF_NP0_159: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S190,
        Q => datapath_theregisterfile_memtrf_186,
        R => controller_rst
    );
DFF_NP0_160: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S191,
        Q => datapath_theregisterfile_memtrf_187,
        R => controller_rst
    );
DFF_NP0_161: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S192,
        Q => datapath_theregisterfile_memtrf_188,
        R => controller_rst
    );
DFF_NP0_162: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S193,
        Q => datapath_theregisterfile_memtrf_189,
        R => controller_rst
    );
DFF_NP0_163: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S194,
        Q => datapath_theregisterfile_memtrf_190,
        R => controller_rst
    );
DFF_NP0_164: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S195,
        Q => datapath_theregisterfile_memtrf_191,
        R => controller_rst
    );
DFF_NP1_29: ENTITY WORK.DFF_NP1
    PORT MAP (
        C => controller_clk,
        D => S196,
        Q => datapath_theregisterfile_memtrf_192,
        R => controller_rst
    );
DFF_NP1_30: ENTITY WORK.DFF_NP1
    PORT MAP (
        C => controller_clk,
        D => S197,
        Q => datapath_theregisterfile_memtrf_193,
        R => controller_rst
    );
DFF_NP0_165: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S198,
        Q => datapath_theregisterfile_memtrf_194,
        R => controller_rst
    );
DFF_NP0_166: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S199,
        Q => datapath_theregisterfile_memtrf_195,
        R => controller_rst
    );
DFF_NP0_167: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S200,
        Q => datapath_theregisterfile_memtrf_196,
        R => controller_rst
    );
DFF_NP0_168: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S201,
        Q => datapath_theregisterfile_memtrf_197,
        R => controller_rst
    );
DFF_NP0_169: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S202,
        Q => datapath_theregisterfile_memtrf_198,
        R => controller_rst
    );
DFF_NP0_170: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S203,
        Q => datapath_theregisterfile_memtrf_199,
        R => controller_rst
    );
DFF_NP0_171: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S204,
        Q => datapath_theregisterfile_memtrf_200,
        R => controller_rst
    );
DFF_NP0_172: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S205,
        Q => datapath_theregisterfile_memtrf_201,
        R => controller_rst
    );
DFF_NP0_173: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S206,
        Q => datapath_theregisterfile_memtrf_202,
        R => controller_rst
    );
DFF_NP0_174: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S207,
        Q => datapath_theregisterfile_memtrf_203,
        R => controller_rst
    );
DFF_NP0_175: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S208,
        Q => datapath_theregisterfile_memtrf_204,
        R => controller_rst
    );
DFF_NP0_176: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S209,
        Q => datapath_theregisterfile_memtrf_205,
        R => controller_rst
    );
DFF_NP0_177: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S210,
        Q => datapath_theregisterfile_memtrf_206,
        R => controller_rst
    );
DFF_NP0_178: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S211,
        Q => datapath_theregisterfile_memtrf_207,
        R => controller_rst
    );
DFF_NP0_179: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S212,
        Q => datapath_theregisterfile_memtrf_208,
        R => controller_rst
    );
DFF_NP1_31: ENTITY WORK.DFF_NP1
    PORT MAP (
        C => controller_clk,
        D => S213,
        Q => datapath_theregisterfile_memtrf_209,
        R => controller_rst
    );
DFF_NP0_180: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S214,
        Q => datapath_theregisterfile_memtrf_210,
        R => controller_rst
    );
DFF_NP0_181: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S215,
        Q => datapath_theregisterfile_memtrf_211,
        R => controller_rst
    );
DFF_NP0_182: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S216,
        Q => datapath_theregisterfile_memtrf_212,
        R => controller_rst
    );
DFF_NP0_183: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S217,
        Q => datapath_theregisterfile_memtrf_213,
        R => controller_rst
    );
DFF_NP0_184: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S218,
        Q => datapath_theregisterfile_memtrf_214,
        R => controller_rst
    );
DFF_NP0_185: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S219,
        Q => datapath_theregisterfile_memtrf_215,
        R => controller_rst
    );
DFF_NP0_186: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S220,
        Q => datapath_theregisterfile_memtrf_216,
        R => controller_rst
    );
DFF_NP0_187: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S221,
        Q => datapath_theregisterfile_memtrf_217,
        R => controller_rst
    );
DFF_NP0_188: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S222,
        Q => datapath_theregisterfile_memtrf_218,
        R => controller_rst
    );
DFF_NP0_189: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S223,
        Q => datapath_theregisterfile_memtrf_219,
        R => controller_rst
    );
DFF_NP0_190: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S224,
        Q => datapath_theregisterfile_memtrf_220,
        R => controller_rst
    );
DFF_NP0_191: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S225,
        Q => datapath_theregisterfile_memtrf_221,
        R => controller_rst
    );
DFF_NP0_192: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S226,
        Q => datapath_theregisterfile_memtrf_222,
        R => controller_rst
    );
DFF_NP0_193: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S227,
        Q => datapath_theregisterfile_memtrf_223,
        R => controller_rst
    );
DFF_NP1_32: ENTITY WORK.DFF_NP1
    PORT MAP (
        C => controller_clk,
        D => S228,
        Q => datapath_theregisterfile_memtrf_224,
        R => controller_rst
    );
DFF_NP0_194: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S229,
        Q => datapath_theregisterfile_memtrf_225,
        R => controller_rst
    );
DFF_NP0_195: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S230,
        Q => datapath_theregisterfile_memtrf_226,
        R => controller_rst
    );
DFF_NP0_196: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S231,
        Q => datapath_theregisterfile_memtrf_227,
        R => controller_rst
    );
DFF_NP0_197: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S232,
        Q => datapath_theregisterfile_memtrf_228,
        R => controller_rst
    );
DFF_NP0_198: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S233,
        Q => datapath_theregisterfile_memtrf_229,
        R => controller_rst
    );
DFF_NP0_199: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S234,
        Q => datapath_theregisterfile_memtrf_230,
        R => controller_rst
    );
DFF_NP0_200: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S235,
        Q => datapath_theregisterfile_memtrf_231,
        R => controller_rst
    );
DFF_NP0_201: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S236,
        Q => datapath_theregisterfile_memtrf_232,
        R => controller_rst
    );
DFF_NP0_202: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S237,
        Q => datapath_theregisterfile_memtrf_233,
        R => controller_rst
    );
DFF_NP0_203: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S238,
        Q => datapath_theregisterfile_memtrf_234,
        R => controller_rst
    );
DFF_NP0_204: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S239,
        Q => datapath_theregisterfile_memtrf_235,
        R => controller_rst
    );
DFF_NP0_205: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S240,
        Q => datapath_theregisterfile_memtrf_236,
        R => controller_rst
    );
DFF_NP0_206: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S241,
        Q => datapath_theregisterfile_memtrf_237,
        R => controller_rst
    );
DFF_NP0_207: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S242,
        Q => datapath_theregisterfile_memtrf_238,
        R => controller_rst
    );
DFF_NP0_208: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S243,
        Q => datapath_theregisterfile_memtrf_239,
        R => controller_rst
    );
DFF_NP0_209: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S244,
        Q => datapath_theregisterfile_memtrf_240,
        R => controller_rst
    );
DFF_NP0_210: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S245,
        Q => datapath_theregisterfile_memtrf_241,
        R => controller_rst
    );
DFF_NP0_211: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S246,
        Q => datapath_theregisterfile_memtrf_242,
        R => controller_rst
    );
DFF_NP0_212: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S247,
        Q => datapath_theregisterfile_memtrf_243,
        R => controller_rst
    );
DFF_NP0_213: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S248,
        Q => datapath_theregisterfile_memtrf_244,
        R => controller_rst
    );
DFF_NP0_214: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S249,
        Q => datapath_theregisterfile_memtrf_245,
        R => controller_rst
    );
DFF_NP0_215: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S250,
        Q => datapath_theregisterfile_memtrf_246,
        R => controller_rst
    );
DFF_NP0_216: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S251,
        Q => datapath_theregisterfile_memtrf_247,
        R => controller_rst
    );
DFF_NP0_217: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S252,
        Q => datapath_theregisterfile_memtrf_248,
        R => controller_rst
    );
DFF_NP0_218: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S253,
        Q => datapath_theregisterfile_memtrf_249,
        R => controller_rst
    );
DFF_NP0_219: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S254,
        Q => datapath_theregisterfile_memtrf_250,
        R => controller_rst
    );
DFF_NP0_220: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S255,
        Q => datapath_theregisterfile_memtrf_251,
        R => controller_rst
    );
DFF_NP0_221: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S256,
        Q => datapath_theregisterfile_memtrf_252,
        R => controller_rst
    );
DFF_NP0_222: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S257,
        Q => datapath_theregisterfile_memtrf_253,
        R => controller_rst
    );
DFF_NP0_223: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S258,
        Q => datapath_theregisterfile_memtrf_254,
        R => controller_rst
    );
DFF_NP0_224: ENTITY WORK.DFF_NP0
    PORT MAP (
        C => controller_clk,
        D => S259,
        Q => datapath_theregisterfile_memtrf_255,
        R => controller_rst
    );
DFF_PP0_83: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S260,
        Q => controller_outflag_0,
        R => controller_rst
    );
DFF_PP0_84: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S261,
        Q => controller_outflag_1,
        R => controller_rst
    );
DFF_PP0_85: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S262,
        Q => controller_outflag_2,
        R => controller_rst
    );
DFF_PP0_86: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S263,
        Q => controller_outflag_3,
        R => controller_rst
    );
DFF_PP0_87: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S264,
        Q => controller_389_B_0,
        R => controller_rst
    );
DFF_PP0_88: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S265,
        Q => controller_389_B_2,
        R => controller_rst
    );
DFF_PP0_89: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S266,
        Q => controller_outflag_6,
        R => controller_rst
    );
DFF_PP0_90: ENTITY WORK.DFF_PP0
    PORT MAP (
        C => controller_clk,
        D => S343,
        Q => controller_outflag_7,
        R => controller_rst
    );
OBUF_1: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_muxmem_in2_0,
        O => PCout(0)
    );
OBUF_2: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_muxmem_in2_1,
        O => PCout(1)
    );
OBUF_3: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_muxmem_in2_10,
        O => PCout(10)
    );
OBUF_4: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_muxmem_in2_11,
        O => PCout(11)
    );
OBUF_5: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_muxmem_in2_12,
        O => PCout(12)
    );
OBUF_6: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_muxmem_in2_13,
        O => PCout(13)
    );
OBUF_7: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_muxmem_in2_14,
        O => PCout(14)
    );
OBUF_8: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_muxmem_in2_15,
        O => PCout(15)
    );
OBUF_9: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_muxmem_in2_2,
        O => PCout(2)
    );
OBUF_10: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_muxmem_in2_3,
        O => PCout(3)
    );
OBUF_11: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_muxmem_in2_4,
        O => PCout(4)
    );
OBUF_12: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_muxmem_in2_5,
        O => PCout(5)
    );
OBUF_13: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_muxmem_in2_6,
        O => PCout(6)
    );
OBUF_14: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_muxmem_in2_7,
        O => PCout(7)
    );
OBUF_15: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_muxmem_in2_8,
        O => PCout(8)
    );
OBUF_16: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_muxmem_in2_9,
        O => PCout(9)
    );
OBUF_17: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_addrbus_0,
        O => addrBus(0)
    );
OBUF_18: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_addrbus_1,
        O => addrBus(1)
    );
OBUF_19: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_addrbus_10,
        O => addrBus(10)
    );
OBUF_20: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_addrbus_11,
        O => addrBus(11)
    );
OBUF_21: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_addrbus_12,
        O => addrBus(12)
    );
OBUF_22: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_addrbus_13,
        O => addrBus(13)
    );
OBUF_23: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_addrbus_14,
        O => addrBus(14)
    );
OBUF_24: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_addrbus_15,
        O => addrBus(15)
    );
OBUF_25: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_addrbus_2,
        O => addrBus(2)
    );
OBUF_26: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_addrbus_3,
        O => addrBus(3)
    );
OBUF_27: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_addrbus_4,
        O => addrBus(4)
    );
OBUF_28: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_addrbus_5,
        O => addrBus(5)
    );
OBUF_29: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_addrbus_6,
        O => addrBus(6)
    );
OBUF_30: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_addrbus_7,
        O => addrBus(7)
    );
OBUF_31: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_addrbus_8,
        O => addrBus(8)
    );
OBUF_32: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_addrbus_9,
        O => addrBus(9)
    );
IBUF_1: ENTITY WORK.IBUF
    PORT MAP (
        I => clk,
        O => controller_clk
    );
IBUF_2: ENTITY WORK.IBUF
    PORT MAP (
        I => dataBusIn(0),
        O => datapath_databusin_0
    );
IBUF_3: ENTITY WORK.IBUF
    PORT MAP (
        I => dataBusIn(1),
        O => datapath_databusin_1
    );
IBUF_4: ENTITY WORK.IBUF
    PORT MAP (
        I => dataBusIn(10),
        O => datapath_databusin_10
    );
IBUF_5: ENTITY WORK.IBUF
    PORT MAP (
        I => dataBusIn(11),
        O => datapath_databusin_11
    );
IBUF_6: ENTITY WORK.IBUF
    PORT MAP (
        I => dataBusIn(12),
        O => datapath_databusin_12
    );
IBUF_7: ENTITY WORK.IBUF
    PORT MAP (
        I => dataBusIn(13),
        O => datapath_databusin_13
    );
IBUF_8: ENTITY WORK.IBUF
    PORT MAP (
        I => dataBusIn(14),
        O => datapath_databusin_14
    );
IBUF_9: ENTITY WORK.IBUF
    PORT MAP (
        I => dataBusIn(15),
        O => datapath_databusin_15
    );
IBUF_10: ENTITY WORK.IBUF
    PORT MAP (
        I => dataBusIn(2),
        O => datapath_databusin_2
    );
IBUF_11: ENTITY WORK.IBUF
    PORT MAP (
        I => dataBusIn(3),
        O => datapath_databusin_3
    );
IBUF_12: ENTITY WORK.IBUF
    PORT MAP (
        I => dataBusIn(4),
        O => datapath_databusin_4
    );
IBUF_13: ENTITY WORK.IBUF
    PORT MAP (
        I => dataBusIn(5),
        O => datapath_databusin_5
    );
IBUF_14: ENTITY WORK.IBUF
    PORT MAP (
        I => dataBusIn(6),
        O => datapath_databusin_6
    );
IBUF_15: ENTITY WORK.IBUF
    PORT MAP (
        I => dataBusIn(7),
        O => datapath_databusin_7
    );
IBUF_16: ENTITY WORK.IBUF
    PORT MAP (
        I => dataBusIn(8),
        O => datapath_databusin_8
    );
IBUF_17: ENTITY WORK.IBUF
    PORT MAP (
        I => dataBusIn(9),
        O => datapath_databusin_9
    );
OBUF_33: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_addsubunit_in1_0,
        O => dataBusOut(0)
    );
OBUF_34: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_addsubunit_in1_1,
        O => dataBusOut(1)
    );
OBUF_35: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_addsubunit_in1_10,
        O => dataBusOut(10)
    );
OBUF_36: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_addsubunit_in1_11,
        O => dataBusOut(11)
    );
OBUF_37: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_addsubunit_in1_12,
        O => dataBusOut(12)
    );
OBUF_38: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_addsubunit_in1_13,
        O => dataBusOut(13)
    );
OBUF_39: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_addsubunit_in1_14,
        O => dataBusOut(14)
    );
OBUF_40: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_addsubunit_in1_15,
        O => dataBusOut(15)
    );
OBUF_41: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_addsubunit_in1_2,
        O => dataBusOut(2)
    );
OBUF_42: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_addsubunit_in1_3,
        O => dataBusOut(3)
    );
OBUF_43: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_addsubunit_in1_4,
        O => dataBusOut(4)
    );
OBUF_44: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_addsubunit_in1_5,
        O => dataBusOut(5)
    );
OBUF_45: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_addsubunit_in1_6,
        O => dataBusOut(6)
    );
OBUF_46: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_addsubunit_in1_7,
        O => dataBusOut(7)
    );
OBUF_47: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_addsubunit_in1_8,
        O => dataBusOut(8)
    );
OBUF_48: ENTITY WORK.OBUF
    PORT MAP (
        I => datapath_addsubunit_in1_9,
        O => dataBusOut(9)
    );
OBUF_49: ENTITY WORK.OBUF
    PORT MAP (
        I => controller_readio,
        O => readIO
    );
OBUF_50: ENTITY WORK.OBUF
    PORT MAP (
        I => controller_1115_S_0,
        O => readInst
    );
OBUF_51: ENTITY WORK.OBUF
    PORT MAP (
        I => controller_readmem,
        O => readMEM
    );
IBUF_18: ENTITY WORK.IBUF
    PORT MAP (
        I => readyMEM,
        O => controller_readymem
    );
IBUF_19: ENTITY WORK.IBUF
    PORT MAP (
        I => rst,
        O => controller_rst
    );
OBUF_52: ENTITY WORK.OBUF
    PORT MAP (
        I => controller_writeio,
        O => writeIO
    );
OBUF_53: ENTITY WORK.OBUF
    PORT MAP (
        I => controller_writemem,
        O => writeMEM
    );

END ARCHITECTURE arch;
