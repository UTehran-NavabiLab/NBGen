module counter(clk, rst, en, clkEn, count, co);

wire _0_;
wire _10_;
wire _11_;
wire _12_;
wire _13_;
wire _14_;
wire _15_;
wire _16_;
wire _17_;
wire _18_;
wire _19_;
wire _1_;
wire _20_;
wire _21_;
wire _22_;
wire _23_;
wire _24_;
wire _25_;
wire _2_;
wire _3_;
wire _4_;
wire _5_;
wire _6_;
wire _7_;
wire _8_;
wire _9_;
input clk;
input rst;
input en;
input clkEn;
output [3:0] count;output co;

INV_X1 #() 
INV_X1_1_ (
  .A({ _20_[2] }),
  .ZN({ _4_ })
);
AND4_X1 #() 
AND4_X1_1_ (
  .A1({ _4_ }),
  .A2({ _20_[3] }),
  .A3({ _20_[1] }),
  .A4({ _20_[0] }),
  .ZN({ _24_ })
);
INV_X1 #() 
INV_X1_2_ (
  .A({ _25_[0] }),
  .ZN({ _5_ })
);
NAND2_X1 #() 
NAND2_X1_1_ (
  .A1({ clkEn }),
  .A2({ en }),
  .ZN({ _6_ })
);
INV_X1 #() 
INV_X1_3_ (
  .A({ rst }),
  .ZN({ _7_ })
);
OAI21_X1 #() 
OAI21_X1_1_ (
  .A({ _7_ }),
  .B1({ _6_ }),
  .B2({ _20_[0] }),
  .ZN({ _8_ })
);
AOI21_X1 #() 
AOI21_X1_1_ (
  .A({ _8_ }),
  .B1({ _6_ }),
  .B2({ _5_ }),
  .ZN({ _0_ })
);
INV_X1 #() 
INV_X1_4_ (
  .A({ _20_[1] }),
  .ZN({ _9_ })
);
NAND3_X1 #() 
NAND3_X1_1_ (
  .A1({ clkEn }),
  .A2({ en }),
  .A3({ _25_[0] }),
  .ZN({ _10_ })
);
NAND4_X1 #() 
NAND4_X1_1_ (
  .A1({ _20_[1] }),
  .A2({ _25_[0] }),
  .A3({ clkEn }),
  .A4({ en }),
  .ZN({ _11_ })
);
NAND2_X1 #() 
NAND2_X1_2_ (
  .A1({ _11_ }),
  .A2({ _7_ }),
  .ZN({ _12_ })
);
AOI21_X1 #() 
AOI21_X1_2_ (
  .A({ _12_ }),
  .B1({ _10_ }),
  .B2({ _9_ }),
  .ZN({ _1_ })
);
NAND2_X1 #() 
NAND2_X1_3_ (
  .A1({ _20_[2] }),
  .A2({ _20_[1] }),
  .ZN({ _13_ })
);
OAI21_X1 #() 
OAI21_X1_2_ (
  .A({ _7_ }),
  .B1({ _10_ }),
  .B2({ _13_ }),
  .ZN({ _14_ })
);
AOI21_X1 #() 
AOI21_X1_3_ (
  .A({ _14_ }),
  .B1({ _11_ }),
  .B2({ _4_ }),
  .ZN({ _2_ })
);
OAI21_X1 #() 
OAI21_X1_3_ (
  .A({ _20_[3] }),
  .B1({ _10_ }),
  .B2({ _13_ }),
  .ZN({ _15_ })
);
INV_X1 #() 
INV_X1_5_ (
  .A({ _20_[3] }),
  .ZN({ _16_ })
);
AND3_X1 #() 
AND3_X1_1_ (
  .A1({ _25_[0] }),
  .A2({ en }),
  .A3({ clkEn }),
  .ZN({ _17_ })
);
AND2_X1 #() 
AND2_X1_1_ (
  .A1({ _20_[1] }),
  .A2({ _20_[2] }),
  .ZN({ _18_ })
);
NAND3_X1 #() 
NAND3_X1_2_ (
  .A1({ _17_ }),
  .A2({ _16_ }),
  .A3({ _18_ }),
  .ZN({ _19_ })
);
AOI21_X1 #() 
AOI21_X1_4_ (
  .A({ rst }),
  .B1({ _19_ }),
  .B2({ _15_ }),
  .ZN({ _3_ })
);
DFF_X1 #() 
DFF_X1_1_ (
  .CK({ clk }),
  .D({ _0_ }),
  .Q({ _25_[0] }),
  .QN({ _20_[0] })
);
DFF_X1 #() 
DFF_X1_2_ (
  .CK({ clk }),
  .D({ _1_ }),
  .Q({ _20_[1] }),
  .QN({ _21_ })
);
DFF_X1 #() 
DFF_X1_3_ (
  .CK({ clk }),
  .D({ _2_ }),
  .Q({ _20_[2] }),
  .QN({ _22_ })
);
DFF_X1 #() 
DFF_X1_4_ (
  .CK({ clk }),
  .D({ _3_ }),
  .Q({ _20_[3] }),
  .QN({ _23_ })
);
BUF_X1 #() 
BUF_X1_1_ (
  .A({ _24_ }),
  .Z({ co })
);
BUF_X1 #() 
BUF_X1_2_ (
  .A({ _25_[0] }),
  .Z({ count[0] })
);
BUF_X1 #() 
BUF_X1_3_ (
  .A({ _20_[1] }),
  .Z({ count[1] })
);
BUF_X1 #() 
BUF_X1_4_ (
  .A({ _20_[2] }),
  .Z({ count[2] })
);
BUF_X1 #() 
BUF_X1_5_ (
  .A({ _20_[3] }),
  .Z({ count[3] })
);

endmodule