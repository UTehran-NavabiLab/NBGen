module sequence(clk, rst, x, out);

wire S0;
wire S1;
wire S2;
wire S3;
wire S4;
wire S5;
wire S6;
wire S7;
wire S8;
wire S9;
wire S10;
wire S11;
wire ns_0;
wire ns_1;
wire ps_0;
wire ps_1;
input clk;
input rst;
input x;
output out;

notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_1_ (
  .A({ ps_1 }),
  .Y({ S3 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_2_ (
  .A({ S9 }),
  .Y({ S4 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_1_ (
  .A({ ps_0, ps_1 }),
  .Y({ S5 })
);
notg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
notg_3_ (
  .A({ S5 }),
  .Y({ S7 })
);
nor_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nor_n_1_ (
  .A({ ps_0, S3 }),
  .Y({ S0 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_2_ (
  .A({ S0, S9 }),
  .Y({ S1 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_3_ (
  .A({ S4, ps_0 }),
  .Y({ S2 })
);
nand_n #( 
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
nand_n_4_ (
  .A({ S2, S1 }),
  .Y({ ns_1 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_1_ (
  .A({ S9 }),
  .Y({ ns_0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_1_ (
  .C({ S6 }),
  .CE({ 1'b1 }),
  .D({ ns_0 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ ps_0 }),
  .R({ S8 }),
  .Si({ S10 }),
  .global_reset({ 1'b0 })
);
dff #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
dff_2_ (
  .C({ S6 }),
  .CE({ 1'b1 }),
  .D({ ns_1 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ ps_1 }),
  .R({ S8 }),
  .Si({ S11 }),
  .global_reset({ 1'b0 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_2_ (
  .A({ clk }),
  .Y({ S6 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_3_ (
  .A({ S7 }),
  .Y({ out })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_4_ (
  .A({ rst }),
  .Y({ S8 })
);
bufg #( 
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)) 
bufg_5_ (
  .A({ x }),
  .Y({ S9 })
);

endmodule