LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

ENTITY MAPn IS
    PORT (
        clk : IN STD_LOGIC;
        rst : IN STD_LOGIC;
        run : IN STD_LOGIC;
        pause : IN STD_LOGIC;
        din : IN STD_LOGIC_VECTOR (383 DOWNTO 0);
        w : IN STD_LOGIC_VECTOR (383 DOWNTO 0);
        reg_out : OUT STD_LOGIC;
        dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0));
END ENTITY MAPn;

ARCHITECTURE arch OF MAPn IS
    SIGNAL S0 : STD_LOGIC;
    SIGNAL S1 : STD_LOGIC;
    SIGNAL S2 : STD_LOGIC;
    SIGNAL S3 : STD_LOGIC;
    SIGNAL S4 : STD_LOGIC;
    SIGNAL S5 : STD_LOGIC;
    SIGNAL S6 : STD_LOGIC;
    SIGNAL S7 : STD_LOGIC;
    SIGNAL data_out_map_0 : STD_LOGIC;
    SIGNAL data_out_map_100 : STD_LOGIC;
    SIGNAL data_out_map_101 : STD_LOGIC;
    SIGNAL data_out_map_102 : STD_LOGIC;
    SIGNAL data_out_map_103 : STD_LOGIC;
    SIGNAL data_out_map_104 : STD_LOGIC;
    SIGNAL data_out_map_105 : STD_LOGIC;
    SIGNAL data_out_map_106 : STD_LOGIC;
    SIGNAL data_out_map_107 : STD_LOGIC;
    SIGNAL data_out_map_108 : STD_LOGIC;
    SIGNAL data_out_map_109 : STD_LOGIC;
    SIGNAL data_out_map_10 : STD_LOGIC;
    SIGNAL data_out_map_110 : STD_LOGIC;
    SIGNAL data_out_map_111 : STD_LOGIC;
    SIGNAL data_out_map_112 : STD_LOGIC;
    SIGNAL data_out_map_113 : STD_LOGIC;
    SIGNAL data_out_map_114 : STD_LOGIC;
    SIGNAL data_out_map_115 : STD_LOGIC;
    SIGNAL data_out_map_116 : STD_LOGIC;
    SIGNAL data_out_map_117 : STD_LOGIC;
    SIGNAL data_out_map_118 : STD_LOGIC;
    SIGNAL data_out_map_119 : STD_LOGIC;
    SIGNAL data_out_map_11 : STD_LOGIC;
    SIGNAL data_out_map_120 : STD_LOGIC;
    SIGNAL data_out_map_121 : STD_LOGIC;
    SIGNAL data_out_map_122 : STD_LOGIC;
    SIGNAL data_out_map_123 : STD_LOGIC;
    SIGNAL data_out_map_124 : STD_LOGIC;
    SIGNAL data_out_map_125 : STD_LOGIC;
    SIGNAL data_out_map_126 : STD_LOGIC;
    SIGNAL data_out_map_127 : STD_LOGIC;
    SIGNAL data_out_map_12 : STD_LOGIC;
    SIGNAL data_out_map_13 : STD_LOGIC;
    SIGNAL data_out_map_14 : STD_LOGIC;
    SIGNAL data_out_map_15 : STD_LOGIC;
    SIGNAL data_out_map_16 : STD_LOGIC;
    SIGNAL data_out_map_17 : STD_LOGIC;
    SIGNAL data_out_map_18 : STD_LOGIC;
    SIGNAL data_out_map_19 : STD_LOGIC;
    SIGNAL data_out_map_1 : STD_LOGIC;
    SIGNAL data_out_map_20 : STD_LOGIC;
    SIGNAL data_out_map_21 : STD_LOGIC;
    SIGNAL data_out_map_22 : STD_LOGIC;
    SIGNAL data_out_map_23 : STD_LOGIC;
    SIGNAL data_out_map_24 : STD_LOGIC;
    SIGNAL data_out_map_25 : STD_LOGIC;
    SIGNAL data_out_map_26 : STD_LOGIC;
    SIGNAL data_out_map_27 : STD_LOGIC;
    SIGNAL data_out_map_28 : STD_LOGIC;
    SIGNAL data_out_map_29 : STD_LOGIC;
    SIGNAL data_out_map_2 : STD_LOGIC;
    SIGNAL data_out_map_30 : STD_LOGIC;
    SIGNAL data_out_map_31 : STD_LOGIC;
    SIGNAL data_out_map_32 : STD_LOGIC;
    SIGNAL data_out_map_33 : STD_LOGIC;
    SIGNAL data_out_map_34 : STD_LOGIC;
    SIGNAL data_out_map_35 : STD_LOGIC;
    SIGNAL data_out_map_36 : STD_LOGIC;
    SIGNAL data_out_map_37 : STD_LOGIC;
    SIGNAL data_out_map_38 : STD_LOGIC;
    SIGNAL data_out_map_39 : STD_LOGIC;
    SIGNAL data_out_map_3 : STD_LOGIC;
    SIGNAL data_out_map_40 : STD_LOGIC;
    SIGNAL data_out_map_41 : STD_LOGIC;
    SIGNAL data_out_map_42 : STD_LOGIC;
    SIGNAL data_out_map_43 : STD_LOGIC;
    SIGNAL data_out_map_44 : STD_LOGIC;
    SIGNAL data_out_map_45 : STD_LOGIC;
    SIGNAL data_out_map_46 : STD_LOGIC;
    SIGNAL data_out_map_47 : STD_LOGIC;
    SIGNAL data_out_map_48 : STD_LOGIC;
    SIGNAL data_out_map_49 : STD_LOGIC;
    SIGNAL data_out_map_4 : STD_LOGIC;
    SIGNAL data_out_map_50 : STD_LOGIC;
    SIGNAL data_out_map_51 : STD_LOGIC;
    SIGNAL data_out_map_52 : STD_LOGIC;
    SIGNAL data_out_map_53 : STD_LOGIC;
    SIGNAL data_out_map_54 : STD_LOGIC;
    SIGNAL data_out_map_55 : STD_LOGIC;
    SIGNAL data_out_map_56 : STD_LOGIC;
    SIGNAL data_out_map_57 : STD_LOGIC;
    SIGNAL data_out_map_58 : STD_LOGIC;
    SIGNAL data_out_map_59 : STD_LOGIC;
    SIGNAL data_out_map_5 : STD_LOGIC;
    SIGNAL data_out_map_60 : STD_LOGIC;
    SIGNAL data_out_map_61 : STD_LOGIC;
    SIGNAL data_out_map_62 : STD_LOGIC;
    SIGNAL data_out_map_63 : STD_LOGIC;
    SIGNAL data_out_map_64 : STD_LOGIC;
    SIGNAL data_out_map_65 : STD_LOGIC;
    SIGNAL data_out_map_66 : STD_LOGIC;
    SIGNAL data_out_map_67 : STD_LOGIC;
    SIGNAL data_out_map_68 : STD_LOGIC;
    SIGNAL data_out_map_69 : STD_LOGIC;
    SIGNAL data_out_map_6 : STD_LOGIC;
    SIGNAL data_out_map_70 : STD_LOGIC;
    SIGNAL data_out_map_71 : STD_LOGIC;
    SIGNAL data_out_map_72 : STD_LOGIC;
    SIGNAL data_out_map_73 : STD_LOGIC;
    SIGNAL data_out_map_74 : STD_LOGIC;
    SIGNAL data_out_map_75 : STD_LOGIC;
    SIGNAL data_out_map_76 : STD_LOGIC;
    SIGNAL data_out_map_77 : STD_LOGIC;
    SIGNAL data_out_map_78 : STD_LOGIC;
    SIGNAL data_out_map_79 : STD_LOGIC;
    SIGNAL data_out_map_7 : STD_LOGIC;
    SIGNAL data_out_map_80 : STD_LOGIC;
    SIGNAL data_out_map_81 : STD_LOGIC;
    SIGNAL data_out_map_82 : STD_LOGIC;
    SIGNAL data_out_map_83 : STD_LOGIC;
    SIGNAL data_out_map_84 : STD_LOGIC;
    SIGNAL data_out_map_85 : STD_LOGIC;
    SIGNAL data_out_map_86 : STD_LOGIC;
    SIGNAL data_out_map_87 : STD_LOGIC;
    SIGNAL data_out_map_88 : STD_LOGIC;
    SIGNAL data_out_map_89 : STD_LOGIC;
    SIGNAL data_out_map_8 : STD_LOGIC;
    SIGNAL data_out_map_90 : STD_LOGIC;
    SIGNAL data_out_map_91 : STD_LOGIC;
    SIGNAL data_out_map_92 : STD_LOGIC;
    SIGNAL data_out_map_93 : STD_LOGIC;
    SIGNAL data_out_map_94 : STD_LOGIC;
    SIGNAL data_out_map_95 : STD_LOGIC;
    SIGNAL data_out_map_96 : STD_LOGIC;
    SIGNAL data_out_map_97 : STD_LOGIC;
    SIGNAL data_out_map_98 : STD_LOGIC;
    SIGNAL data_out_map_99 : STD_LOGIC;
    SIGNAL data_out_map_9 : STD_LOGIC;
    SIGNAL hb0_map_ns_for:1_map_ns:4 : STD_LOGIC;
    SIGNAL hb0_map_ns_for:2_map_ns:13 : STD_LOGIC;
    SIGNAL hb0_map_ns_for:3_map_ns:22 : STD_LOGIC;
    SIGNAL hb0_map_ns_for:4_map_ns:31 : STD_LOGIC;

BEGIN
BUF_X1_1: ENTITY WORK.BUF_X1
    PORT MAP (
        A => clk,
        Z => S0
    );
BUF_X1_2: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(0),
        Z => S1(0)
    );
BUF_X1_3: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(1),
        Z => S1(1)
    );
BUF_X1_4: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(10),
        Z => S1(10)
    );
BUF_X1_5: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(100),
        Z => S1(100)
    );
BUF_X1_6: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(101),
        Z => S1(101)
    );
BUF_X1_7: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(102),
        Z => S1(102)
    );
BUF_X1_8: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(103),
        Z => S1(103)
    );
BUF_X1_9: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(104),
        Z => S1(104)
    );
BUF_X1_10: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(105),
        Z => S1(105)
    );
BUF_X1_11: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(106),
        Z => S1(106)
    );
BUF_X1_12: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(107),
        Z => S1(107)
    );
BUF_X1_13: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(108),
        Z => S1(108)
    );
BUF_X1_14: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(109),
        Z => S1(109)
    );
BUF_X1_15: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(11),
        Z => S1(11)
    );
BUF_X1_16: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(110),
        Z => S1(110)
    );
BUF_X1_17: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(111),
        Z => S1(111)
    );
BUF_X1_18: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(112),
        Z => S1(112)
    );
BUF_X1_19: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(113),
        Z => S1(113)
    );
BUF_X1_20: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(114),
        Z => S1(114)
    );
BUF_X1_21: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(115),
        Z => S1(115)
    );
BUF_X1_22: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(116),
        Z => S1(116)
    );
BUF_X1_23: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(117),
        Z => S1(117)
    );
BUF_X1_24: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(118),
        Z => S1(118)
    );
BUF_X1_25: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(119),
        Z => S1(119)
    );
BUF_X1_26: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(12),
        Z => S1(12)
    );
BUF_X1_27: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(120),
        Z => S1(120)
    );
BUF_X1_28: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(121),
        Z => S1(121)
    );
BUF_X1_29: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(122),
        Z => S1(122)
    );
BUF_X1_30: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(123),
        Z => S1(123)
    );
BUF_X1_31: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(124),
        Z => S1(124)
    );
BUF_X1_32: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(125),
        Z => S1(125)
    );
BUF_X1_33: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(126),
        Z => S1(126)
    );
BUF_X1_34: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(127),
        Z => S1(127)
    );
BUF_X1_35: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(128),
        Z => S1(128)
    );
BUF_X1_36: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(129),
        Z => S1(129)
    );
BUF_X1_37: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(13),
        Z => S1(13)
    );
BUF_X1_38: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(130),
        Z => S1(130)
    );
BUF_X1_39: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(131),
        Z => S1(131)
    );
BUF_X1_40: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(132),
        Z => S1(132)
    );
BUF_X1_41: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(133),
        Z => S1(133)
    );
BUF_X1_42: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(134),
        Z => S1(134)
    );
BUF_X1_43: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(135),
        Z => S1(135)
    );
BUF_X1_44: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(136),
        Z => S1(136)
    );
BUF_X1_45: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(137),
        Z => S1(137)
    );
BUF_X1_46: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(138),
        Z => S1(138)
    );
BUF_X1_47: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(139),
        Z => S1(139)
    );
BUF_X1_48: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(14),
        Z => S1(14)
    );
BUF_X1_49: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(140),
        Z => S1(140)
    );
BUF_X1_50: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(141),
        Z => S1(141)
    );
BUF_X1_51: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(142),
        Z => S1(142)
    );
BUF_X1_52: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(143),
        Z => S1(143)
    );
BUF_X1_53: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(144),
        Z => S1(144)
    );
BUF_X1_54: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(145),
        Z => S1(145)
    );
BUF_X1_55: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(146),
        Z => S1(146)
    );
BUF_X1_56: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(147),
        Z => S1(147)
    );
BUF_X1_57: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(148),
        Z => S1(148)
    );
BUF_X1_58: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(149),
        Z => S1(149)
    );
BUF_X1_59: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(15),
        Z => S1(15)
    );
BUF_X1_60: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(150),
        Z => S1(150)
    );
BUF_X1_61: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(151),
        Z => S1(151)
    );
BUF_X1_62: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(152),
        Z => S1(152)
    );
BUF_X1_63: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(153),
        Z => S1(153)
    );
BUF_X1_64: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(154),
        Z => S1(154)
    );
BUF_X1_65: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(155),
        Z => S1(155)
    );
BUF_X1_66: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(156),
        Z => S1(156)
    );
BUF_X1_67: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(157),
        Z => S1(157)
    );
BUF_X1_68: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(158),
        Z => S1(158)
    );
BUF_X1_69: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(159),
        Z => S1(159)
    );
BUF_X1_70: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(16),
        Z => S1(16)
    );
BUF_X1_71: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(160),
        Z => S1(160)
    );
BUF_X1_72: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(161),
        Z => S1(161)
    );
BUF_X1_73: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(162),
        Z => S1(162)
    );
BUF_X1_74: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(163),
        Z => S1(163)
    );
BUF_X1_75: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(164),
        Z => S1(164)
    );
BUF_X1_76: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(165),
        Z => S1(165)
    );
BUF_X1_77: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(166),
        Z => S1(166)
    );
BUF_X1_78: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(167),
        Z => S1(167)
    );
BUF_X1_79: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(168),
        Z => S1(168)
    );
BUF_X1_80: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(169),
        Z => S1(169)
    );
BUF_X1_81: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(17),
        Z => S1(17)
    );
BUF_X1_82: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(170),
        Z => S1(170)
    );
BUF_X1_83: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(171),
        Z => S1(171)
    );
BUF_X1_84: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(172),
        Z => S1(172)
    );
BUF_X1_85: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(173),
        Z => S1(173)
    );
BUF_X1_86: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(174),
        Z => S1(174)
    );
BUF_X1_87: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(175),
        Z => S1(175)
    );
BUF_X1_88: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(176),
        Z => S1(176)
    );
BUF_X1_89: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(177),
        Z => S1(177)
    );
BUF_X1_90: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(178),
        Z => S1(178)
    );
BUF_X1_91: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(179),
        Z => S1(179)
    );
BUF_X1_92: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(18),
        Z => S1(18)
    );
BUF_X1_93: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(180),
        Z => S1(180)
    );
BUF_X1_94: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(181),
        Z => S1(181)
    );
BUF_X1_95: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(182),
        Z => S1(182)
    );
BUF_X1_96: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(183),
        Z => S1(183)
    );
BUF_X1_97: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(184),
        Z => S1(184)
    );
BUF_X1_98: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(185),
        Z => S1(185)
    );
BUF_X1_99: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(186),
        Z => S1(186)
    );
BUF_X1_100: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(187),
        Z => S1(187)
    );
BUF_X1_101: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(188),
        Z => S1(188)
    );
BUF_X1_102: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(189),
        Z => S1(189)
    );
BUF_X1_103: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(19),
        Z => S1(19)
    );
BUF_X1_104: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(190),
        Z => S1(190)
    );
BUF_X1_105: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(191),
        Z => S1(191)
    );
BUF_X1_106: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(192),
        Z => S1(192)
    );
BUF_X1_107: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(193),
        Z => S1(193)
    );
BUF_X1_108: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(194),
        Z => S1(194)
    );
BUF_X1_109: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(195),
        Z => S1(195)
    );
BUF_X1_110: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(196),
        Z => S1(196)
    );
BUF_X1_111: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(197),
        Z => S1(197)
    );
BUF_X1_112: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(198),
        Z => S1(198)
    );
BUF_X1_113: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(199),
        Z => S1(199)
    );
BUF_X1_114: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(2),
        Z => S1(2)
    );
BUF_X1_115: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(20),
        Z => S1(20)
    );
BUF_X1_116: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(200),
        Z => S1(200)
    );
BUF_X1_117: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(201),
        Z => S1(201)
    );
BUF_X1_118: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(202),
        Z => S1(202)
    );
BUF_X1_119: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(203),
        Z => S1(203)
    );
BUF_X1_120: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(204),
        Z => S1(204)
    );
BUF_X1_121: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(205),
        Z => S1(205)
    );
BUF_X1_122: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(206),
        Z => S1(206)
    );
BUF_X1_123: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(207),
        Z => S1(207)
    );
BUF_X1_124: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(208),
        Z => S1(208)
    );
BUF_X1_125: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(209),
        Z => S1(209)
    );
BUF_X1_126: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(21),
        Z => S1(21)
    );
BUF_X1_127: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(210),
        Z => S1(210)
    );
BUF_X1_128: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(211),
        Z => S1(211)
    );
BUF_X1_129: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(212),
        Z => S1(212)
    );
BUF_X1_130: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(213),
        Z => S1(213)
    );
BUF_X1_131: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(214),
        Z => S1(214)
    );
BUF_X1_132: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(215),
        Z => S1(215)
    );
BUF_X1_133: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(216),
        Z => S1(216)
    );
BUF_X1_134: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(217),
        Z => S1(217)
    );
BUF_X1_135: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(218),
        Z => S1(218)
    );
BUF_X1_136: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(219),
        Z => S1(219)
    );
BUF_X1_137: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(22),
        Z => S1(22)
    );
BUF_X1_138: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(220),
        Z => S1(220)
    );
BUF_X1_139: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(221),
        Z => S1(221)
    );
BUF_X1_140: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(222),
        Z => S1(222)
    );
BUF_X1_141: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(223),
        Z => S1(223)
    );
BUF_X1_142: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(224),
        Z => S1(224)
    );
BUF_X1_143: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(225),
        Z => S1(225)
    );
BUF_X1_144: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(226),
        Z => S1(226)
    );
BUF_X1_145: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(227),
        Z => S1(227)
    );
BUF_X1_146: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(228),
        Z => S1(228)
    );
BUF_X1_147: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(229),
        Z => S1(229)
    );
BUF_X1_148: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(23),
        Z => S1(23)
    );
BUF_X1_149: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(230),
        Z => S1(230)
    );
BUF_X1_150: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(231),
        Z => S1(231)
    );
BUF_X1_151: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(232),
        Z => S1(232)
    );
BUF_X1_152: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(233),
        Z => S1(233)
    );
BUF_X1_153: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(234),
        Z => S1(234)
    );
BUF_X1_154: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(235),
        Z => S1(235)
    );
BUF_X1_155: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(236),
        Z => S1(236)
    );
BUF_X1_156: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(237),
        Z => S1(237)
    );
BUF_X1_157: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(238),
        Z => S1(238)
    );
BUF_X1_158: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(239),
        Z => S1(239)
    );
BUF_X1_159: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(24),
        Z => S1(24)
    );
BUF_X1_160: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(240),
        Z => S1(240)
    );
BUF_X1_161: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(241),
        Z => S1(241)
    );
BUF_X1_162: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(242),
        Z => S1(242)
    );
BUF_X1_163: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(243),
        Z => S1(243)
    );
BUF_X1_164: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(244),
        Z => S1(244)
    );
BUF_X1_165: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(245),
        Z => S1(245)
    );
BUF_X1_166: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(246),
        Z => S1(246)
    );
BUF_X1_167: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(247),
        Z => S1(247)
    );
BUF_X1_168: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(248),
        Z => S1(248)
    );
BUF_X1_169: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(249),
        Z => S1(249)
    );
BUF_X1_170: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(25),
        Z => S1(25)
    );
BUF_X1_171: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(250),
        Z => S1(250)
    );
BUF_X1_172: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(251),
        Z => S1(251)
    );
BUF_X1_173: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(252),
        Z => S1(252)
    );
BUF_X1_174: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(253),
        Z => S1(253)
    );
BUF_X1_175: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(254),
        Z => S1(254)
    );
BUF_X1_176: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(255),
        Z => S1(255)
    );
BUF_X1_177: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(256),
        Z => S1(256)
    );
BUF_X1_178: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(257),
        Z => S1(257)
    );
BUF_X1_179: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(258),
        Z => S1(258)
    );
BUF_X1_180: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(259),
        Z => S1(259)
    );
BUF_X1_181: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(26),
        Z => S1(26)
    );
BUF_X1_182: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(260),
        Z => S1(260)
    );
BUF_X1_183: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(261),
        Z => S1(261)
    );
BUF_X1_184: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(262),
        Z => S1(262)
    );
BUF_X1_185: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(263),
        Z => S1(263)
    );
BUF_X1_186: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(264),
        Z => S1(264)
    );
BUF_X1_187: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(265),
        Z => S1(265)
    );
BUF_X1_188: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(266),
        Z => S1(266)
    );
BUF_X1_189: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(267),
        Z => S1(267)
    );
BUF_X1_190: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(268),
        Z => S1(268)
    );
BUF_X1_191: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(269),
        Z => S1(269)
    );
BUF_X1_192: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(27),
        Z => S1(27)
    );
BUF_X1_193: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(270),
        Z => S1(270)
    );
BUF_X1_194: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(271),
        Z => S1(271)
    );
BUF_X1_195: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(272),
        Z => S1(272)
    );
BUF_X1_196: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(273),
        Z => S1(273)
    );
BUF_X1_197: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(274),
        Z => S1(274)
    );
BUF_X1_198: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(275),
        Z => S1(275)
    );
BUF_X1_199: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(276),
        Z => S1(276)
    );
BUF_X1_200: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(277),
        Z => S1(277)
    );
BUF_X1_201: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(278),
        Z => S1(278)
    );
BUF_X1_202: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(279),
        Z => S1(279)
    );
BUF_X1_203: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(28),
        Z => S1(28)
    );
BUF_X1_204: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(280),
        Z => S1(280)
    );
BUF_X1_205: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(281),
        Z => S1(281)
    );
BUF_X1_206: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(282),
        Z => S1(282)
    );
BUF_X1_207: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(283),
        Z => S1(283)
    );
BUF_X1_208: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(284),
        Z => S1(284)
    );
BUF_X1_209: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(285),
        Z => S1(285)
    );
BUF_X1_210: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(286),
        Z => S1(286)
    );
BUF_X1_211: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(287),
        Z => S1(287)
    );
BUF_X1_212: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(288),
        Z => S1(288)
    );
BUF_X1_213: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(289),
        Z => S1(289)
    );
BUF_X1_214: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(29),
        Z => S1(29)
    );
BUF_X1_215: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(290),
        Z => S1(290)
    );
BUF_X1_216: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(291),
        Z => S1(291)
    );
BUF_X1_217: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(292),
        Z => S1(292)
    );
BUF_X1_218: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(293),
        Z => S1(293)
    );
BUF_X1_219: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(294),
        Z => S1(294)
    );
BUF_X1_220: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(295),
        Z => S1(295)
    );
BUF_X1_221: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(296),
        Z => S1(296)
    );
BUF_X1_222: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(297),
        Z => S1(297)
    );
BUF_X1_223: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(298),
        Z => S1(298)
    );
BUF_X1_224: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(299),
        Z => S1(299)
    );
BUF_X1_225: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(3),
        Z => S1(3)
    );
BUF_X1_226: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(30),
        Z => S1(30)
    );
BUF_X1_227: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(300),
        Z => S1(300)
    );
BUF_X1_228: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(301),
        Z => S1(301)
    );
BUF_X1_229: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(302),
        Z => S1(302)
    );
BUF_X1_230: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(303),
        Z => S1(303)
    );
BUF_X1_231: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(304),
        Z => S1(304)
    );
BUF_X1_232: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(305),
        Z => S1(305)
    );
BUF_X1_233: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(306),
        Z => S1(306)
    );
BUF_X1_234: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(307),
        Z => S1(307)
    );
BUF_X1_235: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(308),
        Z => S1(308)
    );
BUF_X1_236: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(309),
        Z => S1(309)
    );
BUF_X1_237: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(31),
        Z => S1(31)
    );
BUF_X1_238: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(310),
        Z => S1(310)
    );
BUF_X1_239: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(311),
        Z => S1(311)
    );
BUF_X1_240: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(312),
        Z => S1(312)
    );
BUF_X1_241: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(313),
        Z => S1(313)
    );
BUF_X1_242: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(314),
        Z => S1(314)
    );
BUF_X1_243: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(315),
        Z => S1(315)
    );
BUF_X1_244: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(316),
        Z => S1(316)
    );
BUF_X1_245: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(317),
        Z => S1(317)
    );
BUF_X1_246: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(318),
        Z => S1(318)
    );
BUF_X1_247: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(319),
        Z => S1(319)
    );
BUF_X1_248: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(32),
        Z => S1(32)
    );
BUF_X1_249: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(320),
        Z => S1(320)
    );
BUF_X1_250: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(321),
        Z => S1(321)
    );
BUF_X1_251: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(322),
        Z => S1(322)
    );
BUF_X1_252: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(323),
        Z => S1(323)
    );
BUF_X1_253: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(324),
        Z => S1(324)
    );
BUF_X1_254: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(325),
        Z => S1(325)
    );
BUF_X1_255: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(326),
        Z => S1(326)
    );
BUF_X1_256: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(327),
        Z => S1(327)
    );
BUF_X1_257: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(328),
        Z => S1(328)
    );
BUF_X1_258: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(329),
        Z => S1(329)
    );
BUF_X1_259: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(33),
        Z => S1(33)
    );
BUF_X1_260: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(330),
        Z => S1(330)
    );
BUF_X1_261: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(331),
        Z => S1(331)
    );
BUF_X1_262: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(332),
        Z => S1(332)
    );
BUF_X1_263: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(333),
        Z => S1(333)
    );
BUF_X1_264: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(334),
        Z => S1(334)
    );
BUF_X1_265: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(335),
        Z => S1(335)
    );
BUF_X1_266: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(336),
        Z => S1(336)
    );
BUF_X1_267: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(337),
        Z => S1(337)
    );
BUF_X1_268: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(338),
        Z => S1(338)
    );
BUF_X1_269: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(339),
        Z => S1(339)
    );
BUF_X1_270: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(34),
        Z => S1(34)
    );
BUF_X1_271: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(340),
        Z => S1(340)
    );
BUF_X1_272: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(341),
        Z => S1(341)
    );
BUF_X1_273: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(342),
        Z => S1(342)
    );
BUF_X1_274: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(343),
        Z => S1(343)
    );
BUF_X1_275: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(344),
        Z => S1(344)
    );
BUF_X1_276: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(345),
        Z => S1(345)
    );
BUF_X1_277: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(346),
        Z => S1(346)
    );
BUF_X1_278: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(347),
        Z => S1(347)
    );
BUF_X1_279: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(348),
        Z => S1(348)
    );
BUF_X1_280: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(349),
        Z => S1(349)
    );
BUF_X1_281: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(35),
        Z => S1(35)
    );
BUF_X1_282: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(350),
        Z => S1(350)
    );
BUF_X1_283: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(351),
        Z => S1(351)
    );
BUF_X1_284: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(352),
        Z => S1(352)
    );
BUF_X1_285: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(353),
        Z => S1(353)
    );
BUF_X1_286: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(354),
        Z => S1(354)
    );
BUF_X1_287: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(355),
        Z => S1(355)
    );
BUF_X1_288: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(356),
        Z => S1(356)
    );
BUF_X1_289: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(357),
        Z => S1(357)
    );
BUF_X1_290: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(358),
        Z => S1(358)
    );
BUF_X1_291: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(359),
        Z => S1(359)
    );
BUF_X1_292: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(36),
        Z => S1(36)
    );
BUF_X1_293: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(360),
        Z => S1(360)
    );
BUF_X1_294: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(361),
        Z => S1(361)
    );
BUF_X1_295: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(362),
        Z => S1(362)
    );
BUF_X1_296: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(363),
        Z => S1(363)
    );
BUF_X1_297: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(364),
        Z => S1(364)
    );
BUF_X1_298: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(365),
        Z => S1(365)
    );
BUF_X1_299: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(366),
        Z => S1(366)
    );
BUF_X1_300: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(367),
        Z => S1(367)
    );
BUF_X1_301: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(368),
        Z => S1(368)
    );
BUF_X1_302: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(369),
        Z => S1(369)
    );
BUF_X1_303: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(37),
        Z => S1(37)
    );
BUF_X1_304: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(370),
        Z => S1(370)
    );
BUF_X1_305: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(371),
        Z => S1(371)
    );
BUF_X1_306: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(372),
        Z => S1(372)
    );
BUF_X1_307: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(373),
        Z => S1(373)
    );
BUF_X1_308: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(374),
        Z => S1(374)
    );
BUF_X1_309: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(375),
        Z => S1(375)
    );
BUF_X1_310: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(376),
        Z => S1(376)
    );
BUF_X1_311: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(377),
        Z => S1(377)
    );
BUF_X1_312: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(378),
        Z => S1(378)
    );
BUF_X1_313: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(379),
        Z => S1(379)
    );
BUF_X1_314: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(38),
        Z => S1(38)
    );
BUF_X1_315: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(380),
        Z => S1(380)
    );
BUF_X1_316: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(381),
        Z => S1(381)
    );
BUF_X1_317: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(382),
        Z => S1(382)
    );
BUF_X1_318: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(383),
        Z => S1(383)
    );
BUF_X1_319: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(39),
        Z => S1(39)
    );
BUF_X1_320: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(4),
        Z => S1(4)
    );
BUF_X1_321: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(40),
        Z => S1(40)
    );
BUF_X1_322: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(41),
        Z => S1(41)
    );
BUF_X1_323: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(42),
        Z => S1(42)
    );
BUF_X1_324: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(43),
        Z => S1(43)
    );
BUF_X1_325: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(44),
        Z => S1(44)
    );
BUF_X1_326: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(45),
        Z => S1(45)
    );
BUF_X1_327: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(46),
        Z => S1(46)
    );
BUF_X1_328: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(47),
        Z => S1(47)
    );
BUF_X1_329: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(48),
        Z => S1(48)
    );
BUF_X1_330: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(49),
        Z => S1(49)
    );
BUF_X1_331: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(5),
        Z => S1(5)
    );
BUF_X1_332: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(50),
        Z => S1(50)
    );
BUF_X1_333: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(51),
        Z => S1(51)
    );
BUF_X1_334: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(52),
        Z => S1(52)
    );
BUF_X1_335: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(53),
        Z => S1(53)
    );
BUF_X1_336: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(54),
        Z => S1(54)
    );
BUF_X1_337: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(55),
        Z => S1(55)
    );
BUF_X1_338: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(56),
        Z => S1(56)
    );
BUF_X1_339: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(57),
        Z => S1(57)
    );
BUF_X1_340: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(58),
        Z => S1(58)
    );
BUF_X1_341: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(59),
        Z => S1(59)
    );
BUF_X1_342: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(6),
        Z => S1(6)
    );
BUF_X1_343: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(60),
        Z => S1(60)
    );
BUF_X1_344: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(61),
        Z => S1(61)
    );
BUF_X1_345: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(62),
        Z => S1(62)
    );
BUF_X1_346: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(63),
        Z => S1(63)
    );
BUF_X1_347: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(64),
        Z => S1(64)
    );
BUF_X1_348: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(65),
        Z => S1(65)
    );
BUF_X1_349: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(66),
        Z => S1(66)
    );
BUF_X1_350: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(67),
        Z => S1(67)
    );
BUF_X1_351: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(68),
        Z => S1(68)
    );
BUF_X1_352: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(69),
        Z => S1(69)
    );
BUF_X1_353: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(7),
        Z => S1(7)
    );
BUF_X1_354: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(70),
        Z => S1(70)
    );
BUF_X1_355: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(71),
        Z => S1(71)
    );
BUF_X1_356: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(72),
        Z => S1(72)
    );
BUF_X1_357: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(73),
        Z => S1(73)
    );
BUF_X1_358: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(74),
        Z => S1(74)
    );
BUF_X1_359: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(75),
        Z => S1(75)
    );
BUF_X1_360: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(76),
        Z => S1(76)
    );
BUF_X1_361: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(77),
        Z => S1(77)
    );
BUF_X1_362: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(78),
        Z => S1(78)
    );
BUF_X1_363: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(79),
        Z => S1(79)
    );
BUF_X1_364: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(8),
        Z => S1(8)
    );
BUF_X1_365: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(80),
        Z => S1(80)
    );
BUF_X1_366: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(81),
        Z => S1(81)
    );
BUF_X1_367: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(82),
        Z => S1(82)
    );
BUF_X1_368: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(83),
        Z => S1(83)
    );
BUF_X1_369: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(84),
        Z => S1(84)
    );
BUF_X1_370: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(85),
        Z => S1(85)
    );
BUF_X1_371: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(86),
        Z => S1(86)
    );
BUF_X1_372: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(87),
        Z => S1(87)
    );
BUF_X1_373: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(88),
        Z => S1(88)
    );
BUF_X1_374: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(89),
        Z => S1(89)
    );
BUF_X1_375: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(9),
        Z => S1(9)
    );
BUF_X1_376: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(90),
        Z => S1(90)
    );
BUF_X1_377: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(91),
        Z => S1(91)
    );
BUF_X1_378: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(92),
        Z => S1(92)
    );
BUF_X1_379: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(93),
        Z => S1(93)
    );
BUF_X1_380: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(94),
        Z => S1(94)
    );
BUF_X1_381: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(95),
        Z => S1(95)
    );
BUF_X1_382: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(96),
        Z => S1(96)
    );
BUF_X1_383: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(97),
        Z => S1(97)
    );
BUF_X1_384: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(98),
        Z => S1(98)
    );
BUF_X1_385: ENTITY WORK.BUF_X1
    PORT MAP (
        A => din(99),
        Z => S1(99)
    );
BUF_X1_386: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S2(0),
        Z => dout(0)
    );
BUF_X1_387: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S2(1),
        Z => dout(1)
    );
BUF_X1_388: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S2(10),
        Z => dout(10)
    );
BUF_X1_389: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S2(11),
        Z => dout(11)
    );
BUF_X1_390: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S2(12),
        Z => dout(12)
    );
BUF_X1_391: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S2(13),
        Z => dout(13)
    );
BUF_X1_392: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S2(14),
        Z => dout(14)
    );
BUF_X1_393: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S2(15),
        Z => dout(15)
    );
BUF_X1_394: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S2(16),
        Z => dout(16)
    );
BUF_X1_395: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S2(17),
        Z => dout(17)
    );
BUF_X1_396: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S2(18),
        Z => dout(18)
    );
BUF_X1_397: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S2(19),
        Z => dout(19)
    );
BUF_X1_398: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S2(2),
        Z => dout(2)
    );
BUF_X1_399: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S2(20),
        Z => dout(20)
    );
BUF_X1_400: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S2(21),
        Z => dout(21)
    );
BUF_X1_401: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S2(22),
        Z => dout(22)
    );
BUF_X1_402: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S2(23),
        Z => dout(23)
    );
BUF_X1_403: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S2(24),
        Z => dout(24)
    );
BUF_X1_404: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S2(25),
        Z => dout(25)
    );
BUF_X1_405: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S2(26),
        Z => dout(26)
    );
BUF_X1_406: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S2(27),
        Z => dout(27)
    );
BUF_X1_407: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S2(28),
        Z => dout(28)
    );
BUF_X1_408: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S2(29),
        Z => dout(29)
    );
BUF_X1_409: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S2(3),
        Z => dout(3)
    );
BUF_X1_410: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S2(30),
        Z => dout(30)
    );
BUF_X1_411: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S2(31),
        Z => dout(31)
    );
BUF_X1_412: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S2(4),
        Z => dout(4)
    );
BUF_X1_413: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S2(5),
        Z => dout(5)
    );
BUF_X1_414: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S2(6),
        Z => dout(6)
    );
BUF_X1_415: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S2(7),
        Z => dout(7)
    );
BUF_X1_416: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S2(8),
        Z => dout(8)
    );
BUF_X1_417: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S2(9),
        Z => dout(9)
    );
BUF_X1_418: ENTITY WORK.BUF_X1
    PORT MAP (
        A => pause,
        Z => S3
    );
BUF_X1_419: ENTITY WORK.BUF_X1
    PORT MAP (
        A => S4,
        Z => reg_out
    );
BUF_X1_420: ENTITY WORK.BUF_X1
    PORT MAP (
        A => rst,
        Z => S5
    );
BUF_X1_421: ENTITY WORK.BUF_X1
    PORT MAP (
        A => run,
        Z => S6
    );
BUF_X1_422: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(0),
        Z => S7(0)
    );
BUF_X1_423: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(1),
        Z => S7(1)
    );
BUF_X1_424: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(10),
        Z => S7(10)
    );
BUF_X1_425: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(100),
        Z => S7(100)
    );
BUF_X1_426: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(101),
        Z => S7(101)
    );
BUF_X1_427: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(102),
        Z => S7(102)
    );
BUF_X1_428: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(103),
        Z => S7(103)
    );
BUF_X1_429: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(104),
        Z => S7(104)
    );
BUF_X1_430: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(105),
        Z => S7(105)
    );
BUF_X1_431: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(106),
        Z => S7(106)
    );
BUF_X1_432: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(107),
        Z => S7(107)
    );
BUF_X1_433: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(108),
        Z => S7(108)
    );
BUF_X1_434: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(109),
        Z => S7(109)
    );
BUF_X1_435: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(11),
        Z => S7(11)
    );
BUF_X1_436: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(110),
        Z => S7(110)
    );
BUF_X1_437: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(111),
        Z => S7(111)
    );
BUF_X1_438: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(112),
        Z => S7(112)
    );
BUF_X1_439: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(113),
        Z => S7(113)
    );
BUF_X1_440: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(114),
        Z => S7(114)
    );
BUF_X1_441: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(115),
        Z => S7(115)
    );
BUF_X1_442: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(116),
        Z => S7(116)
    );
BUF_X1_443: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(117),
        Z => S7(117)
    );
BUF_X1_444: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(118),
        Z => S7(118)
    );
BUF_X1_445: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(119),
        Z => S7(119)
    );
BUF_X1_446: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(12),
        Z => S7(12)
    );
BUF_X1_447: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(120),
        Z => S7(120)
    );
BUF_X1_448: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(121),
        Z => S7(121)
    );
BUF_X1_449: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(122),
        Z => S7(122)
    );
BUF_X1_450: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(123),
        Z => S7(123)
    );
BUF_X1_451: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(124),
        Z => S7(124)
    );
BUF_X1_452: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(125),
        Z => S7(125)
    );
BUF_X1_453: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(126),
        Z => S7(126)
    );
BUF_X1_454: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(127),
        Z => S7(127)
    );
BUF_X1_455: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(128),
        Z => S7(128)
    );
BUF_X1_456: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(129),
        Z => S7(129)
    );
BUF_X1_457: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(13),
        Z => S7(13)
    );
BUF_X1_458: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(130),
        Z => S7(130)
    );
BUF_X1_459: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(131),
        Z => S7(131)
    );
BUF_X1_460: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(132),
        Z => S7(132)
    );
BUF_X1_461: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(133),
        Z => S7(133)
    );
BUF_X1_462: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(134),
        Z => S7(134)
    );
BUF_X1_463: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(135),
        Z => S7(135)
    );
BUF_X1_464: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(136),
        Z => S7(136)
    );
BUF_X1_465: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(137),
        Z => S7(137)
    );
BUF_X1_466: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(138),
        Z => S7(138)
    );
BUF_X1_467: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(139),
        Z => S7(139)
    );
BUF_X1_468: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(14),
        Z => S7(14)
    );
BUF_X1_469: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(140),
        Z => S7(140)
    );
BUF_X1_470: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(141),
        Z => S7(141)
    );
BUF_X1_471: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(142),
        Z => S7(142)
    );
BUF_X1_472: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(143),
        Z => S7(143)
    );
BUF_X1_473: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(144),
        Z => S7(144)
    );
BUF_X1_474: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(145),
        Z => S7(145)
    );
BUF_X1_475: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(146),
        Z => S7(146)
    );
BUF_X1_476: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(147),
        Z => S7(147)
    );
BUF_X1_477: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(148),
        Z => S7(148)
    );
BUF_X1_478: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(149),
        Z => S7(149)
    );
BUF_X1_479: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(15),
        Z => S7(15)
    );
BUF_X1_480: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(150),
        Z => S7(150)
    );
BUF_X1_481: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(151),
        Z => S7(151)
    );
BUF_X1_482: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(152),
        Z => S7(152)
    );
BUF_X1_483: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(153),
        Z => S7(153)
    );
BUF_X1_484: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(154),
        Z => S7(154)
    );
BUF_X1_485: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(155),
        Z => S7(155)
    );
BUF_X1_486: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(156),
        Z => S7(156)
    );
BUF_X1_487: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(157),
        Z => S7(157)
    );
BUF_X1_488: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(158),
        Z => S7(158)
    );
BUF_X1_489: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(159),
        Z => S7(159)
    );
BUF_X1_490: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(16),
        Z => S7(16)
    );
BUF_X1_491: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(160),
        Z => S7(160)
    );
BUF_X1_492: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(161),
        Z => S7(161)
    );
BUF_X1_493: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(162),
        Z => S7(162)
    );
BUF_X1_494: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(163),
        Z => S7(163)
    );
BUF_X1_495: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(164),
        Z => S7(164)
    );
BUF_X1_496: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(165),
        Z => S7(165)
    );
BUF_X1_497: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(166),
        Z => S7(166)
    );
BUF_X1_498: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(167),
        Z => S7(167)
    );
BUF_X1_499: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(168),
        Z => S7(168)
    );
BUF_X1_500: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(169),
        Z => S7(169)
    );
BUF_X1_501: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(17),
        Z => S7(17)
    );
BUF_X1_502: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(170),
        Z => S7(170)
    );
BUF_X1_503: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(171),
        Z => S7(171)
    );
BUF_X1_504: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(172),
        Z => S7(172)
    );
BUF_X1_505: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(173),
        Z => S7(173)
    );
BUF_X1_506: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(174),
        Z => S7(174)
    );
BUF_X1_507: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(175),
        Z => S7(175)
    );
BUF_X1_508: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(176),
        Z => S7(176)
    );
BUF_X1_509: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(177),
        Z => S7(177)
    );
BUF_X1_510: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(178),
        Z => S7(178)
    );
BUF_X1_511: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(179),
        Z => S7(179)
    );
BUF_X1_512: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(18),
        Z => S7(18)
    );
BUF_X1_513: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(180),
        Z => S7(180)
    );
BUF_X1_514: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(181),
        Z => S7(181)
    );
BUF_X1_515: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(182),
        Z => S7(182)
    );
BUF_X1_516: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(183),
        Z => S7(183)
    );
BUF_X1_517: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(184),
        Z => S7(184)
    );
BUF_X1_518: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(185),
        Z => S7(185)
    );
BUF_X1_519: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(186),
        Z => S7(186)
    );
BUF_X1_520: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(187),
        Z => S7(187)
    );
BUF_X1_521: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(188),
        Z => S7(188)
    );
BUF_X1_522: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(189),
        Z => S7(189)
    );
BUF_X1_523: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(19),
        Z => S7(19)
    );
BUF_X1_524: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(190),
        Z => S7(190)
    );
BUF_X1_525: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(191),
        Z => S7(191)
    );
BUF_X1_526: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(192),
        Z => S7(192)
    );
BUF_X1_527: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(193),
        Z => S7(193)
    );
BUF_X1_528: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(194),
        Z => S7(194)
    );
BUF_X1_529: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(195),
        Z => S7(195)
    );
BUF_X1_530: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(196),
        Z => S7(196)
    );
BUF_X1_531: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(197),
        Z => S7(197)
    );
BUF_X1_532: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(198),
        Z => S7(198)
    );
BUF_X1_533: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(199),
        Z => S7(199)
    );
BUF_X1_534: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(2),
        Z => S7(2)
    );
BUF_X1_535: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(20),
        Z => S7(20)
    );
BUF_X1_536: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(200),
        Z => S7(200)
    );
BUF_X1_537: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(201),
        Z => S7(201)
    );
BUF_X1_538: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(202),
        Z => S7(202)
    );
BUF_X1_539: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(203),
        Z => S7(203)
    );
BUF_X1_540: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(204),
        Z => S7(204)
    );
BUF_X1_541: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(205),
        Z => S7(205)
    );
BUF_X1_542: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(206),
        Z => S7(206)
    );
BUF_X1_543: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(207),
        Z => S7(207)
    );
BUF_X1_544: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(208),
        Z => S7(208)
    );
BUF_X1_545: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(209),
        Z => S7(209)
    );
BUF_X1_546: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(21),
        Z => S7(21)
    );
BUF_X1_547: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(210),
        Z => S7(210)
    );
BUF_X1_548: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(211),
        Z => S7(211)
    );
BUF_X1_549: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(212),
        Z => S7(212)
    );
BUF_X1_550: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(213),
        Z => S7(213)
    );
BUF_X1_551: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(214),
        Z => S7(214)
    );
BUF_X1_552: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(215),
        Z => S7(215)
    );
BUF_X1_553: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(216),
        Z => S7(216)
    );
BUF_X1_554: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(217),
        Z => S7(217)
    );
BUF_X1_555: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(218),
        Z => S7(218)
    );
BUF_X1_556: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(219),
        Z => S7(219)
    );
BUF_X1_557: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(22),
        Z => S7(22)
    );
BUF_X1_558: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(220),
        Z => S7(220)
    );
BUF_X1_559: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(221),
        Z => S7(221)
    );
BUF_X1_560: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(222),
        Z => S7(222)
    );
BUF_X1_561: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(223),
        Z => S7(223)
    );
BUF_X1_562: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(224),
        Z => S7(224)
    );
BUF_X1_563: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(225),
        Z => S7(225)
    );
BUF_X1_564: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(226),
        Z => S7(226)
    );
BUF_X1_565: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(227),
        Z => S7(227)
    );
BUF_X1_566: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(228),
        Z => S7(228)
    );
BUF_X1_567: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(229),
        Z => S7(229)
    );
BUF_X1_568: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(23),
        Z => S7(23)
    );
BUF_X1_569: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(230),
        Z => S7(230)
    );
BUF_X1_570: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(231),
        Z => S7(231)
    );
BUF_X1_571: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(232),
        Z => S7(232)
    );
BUF_X1_572: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(233),
        Z => S7(233)
    );
BUF_X1_573: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(234),
        Z => S7(234)
    );
BUF_X1_574: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(235),
        Z => S7(235)
    );
BUF_X1_575: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(236),
        Z => S7(236)
    );
BUF_X1_576: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(237),
        Z => S7(237)
    );
BUF_X1_577: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(238),
        Z => S7(238)
    );
BUF_X1_578: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(239),
        Z => S7(239)
    );
BUF_X1_579: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(24),
        Z => S7(24)
    );
BUF_X1_580: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(240),
        Z => S7(240)
    );
BUF_X1_581: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(241),
        Z => S7(241)
    );
BUF_X1_582: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(242),
        Z => S7(242)
    );
BUF_X1_583: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(243),
        Z => S7(243)
    );
BUF_X1_584: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(244),
        Z => S7(244)
    );
BUF_X1_585: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(245),
        Z => S7(245)
    );
BUF_X1_586: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(246),
        Z => S7(246)
    );
BUF_X1_587: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(247),
        Z => S7(247)
    );
BUF_X1_588: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(248),
        Z => S7(248)
    );
BUF_X1_589: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(249),
        Z => S7(249)
    );
BUF_X1_590: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(25),
        Z => S7(25)
    );
BUF_X1_591: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(250),
        Z => S7(250)
    );
BUF_X1_592: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(251),
        Z => S7(251)
    );
BUF_X1_593: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(252),
        Z => S7(252)
    );
BUF_X1_594: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(253),
        Z => S7(253)
    );
BUF_X1_595: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(254),
        Z => S7(254)
    );
BUF_X1_596: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(255),
        Z => S7(255)
    );
BUF_X1_597: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(256),
        Z => S7(256)
    );
BUF_X1_598: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(257),
        Z => S7(257)
    );
BUF_X1_599: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(258),
        Z => S7(258)
    );
BUF_X1_600: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(259),
        Z => S7(259)
    );
BUF_X1_601: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(26),
        Z => S7(26)
    );
BUF_X1_602: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(260),
        Z => S7(260)
    );
BUF_X1_603: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(261),
        Z => S7(261)
    );
BUF_X1_604: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(262),
        Z => S7(262)
    );
BUF_X1_605: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(263),
        Z => S7(263)
    );
BUF_X1_606: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(264),
        Z => S7(264)
    );
BUF_X1_607: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(265),
        Z => S7(265)
    );
BUF_X1_608: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(266),
        Z => S7(266)
    );
BUF_X1_609: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(267),
        Z => S7(267)
    );
BUF_X1_610: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(268),
        Z => S7(268)
    );
BUF_X1_611: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(269),
        Z => S7(269)
    );
BUF_X1_612: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(27),
        Z => S7(27)
    );
BUF_X1_613: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(270),
        Z => S7(270)
    );
BUF_X1_614: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(271),
        Z => S7(271)
    );
BUF_X1_615: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(272),
        Z => S7(272)
    );
BUF_X1_616: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(273),
        Z => S7(273)
    );
BUF_X1_617: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(274),
        Z => S7(274)
    );
BUF_X1_618: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(275),
        Z => S7(275)
    );
BUF_X1_619: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(276),
        Z => S7(276)
    );
BUF_X1_620: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(277),
        Z => S7(277)
    );
BUF_X1_621: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(278),
        Z => S7(278)
    );
BUF_X1_622: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(279),
        Z => S7(279)
    );
BUF_X1_623: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(28),
        Z => S7(28)
    );
BUF_X1_624: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(280),
        Z => S7(280)
    );
BUF_X1_625: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(281),
        Z => S7(281)
    );
BUF_X1_626: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(282),
        Z => S7(282)
    );
BUF_X1_627: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(283),
        Z => S7(283)
    );
BUF_X1_628: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(284),
        Z => S7(284)
    );
BUF_X1_629: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(285),
        Z => S7(285)
    );
BUF_X1_630: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(286),
        Z => S7(286)
    );
BUF_X1_631: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(287),
        Z => S7(287)
    );
BUF_X1_632: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(288),
        Z => S7(288)
    );
BUF_X1_633: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(289),
        Z => S7(289)
    );
BUF_X1_634: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(29),
        Z => S7(29)
    );
BUF_X1_635: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(290),
        Z => S7(290)
    );
BUF_X1_636: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(291),
        Z => S7(291)
    );
BUF_X1_637: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(292),
        Z => S7(292)
    );
BUF_X1_638: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(293),
        Z => S7(293)
    );
BUF_X1_639: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(294),
        Z => S7(294)
    );
BUF_X1_640: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(295),
        Z => S7(295)
    );
BUF_X1_641: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(296),
        Z => S7(296)
    );
BUF_X1_642: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(297),
        Z => S7(297)
    );
BUF_X1_643: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(298),
        Z => S7(298)
    );
BUF_X1_644: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(299),
        Z => S7(299)
    );
BUF_X1_645: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(3),
        Z => S7(3)
    );
BUF_X1_646: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(30),
        Z => S7(30)
    );
BUF_X1_647: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(300),
        Z => S7(300)
    );
BUF_X1_648: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(301),
        Z => S7(301)
    );
BUF_X1_649: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(302),
        Z => S7(302)
    );
BUF_X1_650: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(303),
        Z => S7(303)
    );
BUF_X1_651: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(304),
        Z => S7(304)
    );
BUF_X1_652: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(305),
        Z => S7(305)
    );
BUF_X1_653: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(306),
        Z => S7(306)
    );
BUF_X1_654: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(307),
        Z => S7(307)
    );
BUF_X1_655: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(308),
        Z => S7(308)
    );
BUF_X1_656: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(309),
        Z => S7(309)
    );
BUF_X1_657: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(31),
        Z => S7(31)
    );
BUF_X1_658: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(310),
        Z => S7(310)
    );
BUF_X1_659: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(311),
        Z => S7(311)
    );
BUF_X1_660: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(312),
        Z => S7(312)
    );
BUF_X1_661: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(313),
        Z => S7(313)
    );
BUF_X1_662: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(314),
        Z => S7(314)
    );
BUF_X1_663: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(315),
        Z => S7(315)
    );
BUF_X1_664: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(316),
        Z => S7(316)
    );
BUF_X1_665: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(317),
        Z => S7(317)
    );
BUF_X1_666: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(318),
        Z => S7(318)
    );
BUF_X1_667: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(319),
        Z => S7(319)
    );
BUF_X1_668: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(32),
        Z => S7(32)
    );
BUF_X1_669: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(320),
        Z => S7(320)
    );
BUF_X1_670: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(321),
        Z => S7(321)
    );
BUF_X1_671: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(322),
        Z => S7(322)
    );
BUF_X1_672: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(323),
        Z => S7(323)
    );
BUF_X1_673: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(324),
        Z => S7(324)
    );
BUF_X1_674: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(325),
        Z => S7(325)
    );
BUF_X1_675: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(326),
        Z => S7(326)
    );
BUF_X1_676: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(327),
        Z => S7(327)
    );
BUF_X1_677: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(328),
        Z => S7(328)
    );
BUF_X1_678: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(329),
        Z => S7(329)
    );
BUF_X1_679: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(33),
        Z => S7(33)
    );
BUF_X1_680: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(330),
        Z => S7(330)
    );
BUF_X1_681: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(331),
        Z => S7(331)
    );
BUF_X1_682: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(332),
        Z => S7(332)
    );
BUF_X1_683: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(333),
        Z => S7(333)
    );
BUF_X1_684: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(334),
        Z => S7(334)
    );
BUF_X1_685: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(335),
        Z => S7(335)
    );
BUF_X1_686: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(336),
        Z => S7(336)
    );
BUF_X1_687: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(337),
        Z => S7(337)
    );
BUF_X1_688: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(338),
        Z => S7(338)
    );
BUF_X1_689: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(339),
        Z => S7(339)
    );
BUF_X1_690: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(34),
        Z => S7(34)
    );
BUF_X1_691: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(340),
        Z => S7(340)
    );
BUF_X1_692: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(341),
        Z => S7(341)
    );
BUF_X1_693: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(342),
        Z => S7(342)
    );
BUF_X1_694: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(343),
        Z => S7(343)
    );
BUF_X1_695: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(344),
        Z => S7(344)
    );
BUF_X1_696: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(345),
        Z => S7(345)
    );
BUF_X1_697: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(346),
        Z => S7(346)
    );
BUF_X1_698: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(347),
        Z => S7(347)
    );
BUF_X1_699: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(348),
        Z => S7(348)
    );
BUF_X1_700: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(349),
        Z => S7(349)
    );
BUF_X1_701: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(35),
        Z => S7(35)
    );
BUF_X1_702: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(350),
        Z => S7(350)
    );
BUF_X1_703: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(351),
        Z => S7(351)
    );
BUF_X1_704: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(352),
        Z => S7(352)
    );
BUF_X1_705: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(353),
        Z => S7(353)
    );
BUF_X1_706: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(354),
        Z => S7(354)
    );
BUF_X1_707: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(355),
        Z => S7(355)
    );
BUF_X1_708: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(356),
        Z => S7(356)
    );
BUF_X1_709: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(357),
        Z => S7(357)
    );
BUF_X1_710: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(358),
        Z => S7(358)
    );
BUF_X1_711: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(359),
        Z => S7(359)
    );
BUF_X1_712: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(36),
        Z => S7(36)
    );
BUF_X1_713: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(360),
        Z => S7(360)
    );
BUF_X1_714: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(361),
        Z => S7(361)
    );
BUF_X1_715: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(362),
        Z => S7(362)
    );
BUF_X1_716: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(363),
        Z => S7(363)
    );
BUF_X1_717: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(364),
        Z => S7(364)
    );
BUF_X1_718: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(365),
        Z => S7(365)
    );
BUF_X1_719: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(366),
        Z => S7(366)
    );
BUF_X1_720: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(367),
        Z => S7(367)
    );
BUF_X1_721: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(368),
        Z => S7(368)
    );
BUF_X1_722: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(369),
        Z => S7(369)
    );
BUF_X1_723: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(37),
        Z => S7(37)
    );
BUF_X1_724: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(370),
        Z => S7(370)
    );
BUF_X1_725: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(371),
        Z => S7(371)
    );
BUF_X1_726: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(372),
        Z => S7(372)
    );
BUF_X1_727: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(373),
        Z => S7(373)
    );
BUF_X1_728: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(374),
        Z => S7(374)
    );
BUF_X1_729: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(375),
        Z => S7(375)
    );
BUF_X1_730: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(376),
        Z => S7(376)
    );
BUF_X1_731: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(377),
        Z => S7(377)
    );
BUF_X1_732: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(378),
        Z => S7(378)
    );
BUF_X1_733: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(379),
        Z => S7(379)
    );
BUF_X1_734: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(38),
        Z => S7(38)
    );
BUF_X1_735: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(380),
        Z => S7(380)
    );
BUF_X1_736: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(381),
        Z => S7(381)
    );
BUF_X1_737: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(382),
        Z => S7(382)
    );
BUF_X1_738: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(383),
        Z => S7(383)
    );
BUF_X1_739: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(39),
        Z => S7(39)
    );
BUF_X1_740: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(4),
        Z => S7(4)
    );
BUF_X1_741: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(40),
        Z => S7(40)
    );
BUF_X1_742: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(41),
        Z => S7(41)
    );
BUF_X1_743: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(42),
        Z => S7(42)
    );
BUF_X1_744: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(43),
        Z => S7(43)
    );
BUF_X1_745: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(44),
        Z => S7(44)
    );
BUF_X1_746: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(45),
        Z => S7(45)
    );
BUF_X1_747: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(46),
        Z => S7(46)
    );
BUF_X1_748: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(47),
        Z => S7(47)
    );
BUF_X1_749: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(48),
        Z => S7(48)
    );
BUF_X1_750: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(49),
        Z => S7(49)
    );
BUF_X1_751: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(5),
        Z => S7(5)
    );
BUF_X1_752: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(50),
        Z => S7(50)
    );
BUF_X1_753: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(51),
        Z => S7(51)
    );
BUF_X1_754: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(52),
        Z => S7(52)
    );
BUF_X1_755: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(53),
        Z => S7(53)
    );
BUF_X1_756: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(54),
        Z => S7(54)
    );
BUF_X1_757: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(55),
        Z => S7(55)
    );
BUF_X1_758: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(56),
        Z => S7(56)
    );
BUF_X1_759: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(57),
        Z => S7(57)
    );
BUF_X1_760: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(58),
        Z => S7(58)
    );
BUF_X1_761: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(59),
        Z => S7(59)
    );
BUF_X1_762: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(6),
        Z => S7(6)
    );
BUF_X1_763: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(60),
        Z => S7(60)
    );
BUF_X1_764: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(61),
        Z => S7(61)
    );
BUF_X1_765: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(62),
        Z => S7(62)
    );
BUF_X1_766: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(63),
        Z => S7(63)
    );
BUF_X1_767: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(64),
        Z => S7(64)
    );
BUF_X1_768: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(65),
        Z => S7(65)
    );
BUF_X1_769: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(66),
        Z => S7(66)
    );
BUF_X1_770: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(67),
        Z => S7(67)
    );
BUF_X1_771: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(68),
        Z => S7(68)
    );
BUF_X1_772: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(69),
        Z => S7(69)
    );
BUF_X1_773: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(7),
        Z => S7(7)
    );
BUF_X1_774: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(70),
        Z => S7(70)
    );
BUF_X1_775: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(71),
        Z => S7(71)
    );
BUF_X1_776: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(72),
        Z => S7(72)
    );
BUF_X1_777: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(73),
        Z => S7(73)
    );
BUF_X1_778: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(74),
        Z => S7(74)
    );
BUF_X1_779: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(75),
        Z => S7(75)
    );
BUF_X1_780: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(76),
        Z => S7(76)
    );
BUF_X1_781: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(77),
        Z => S7(77)
    );
BUF_X1_782: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(78),
        Z => S7(78)
    );
BUF_X1_783: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(79),
        Z => S7(79)
    );
BUF_X1_784: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(8),
        Z => S7(8)
    );
BUF_X1_785: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(80),
        Z => S7(80)
    );
BUF_X1_786: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(81),
        Z => S7(81)
    );
BUF_X1_787: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(82),
        Z => S7(82)
    );
BUF_X1_788: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(83),
        Z => S7(83)
    );
BUF_X1_789: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(84),
        Z => S7(84)
    );
BUF_X1_790: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(85),
        Z => S7(85)
    );
BUF_X1_791: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(86),
        Z => S7(86)
    );
BUF_X1_792: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(87),
        Z => S7(87)
    );
BUF_X1_793: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(88),
        Z => S7(88)
    );
BUF_X1_794: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(89),
        Z => S7(89)
    );
BUF_X1_795: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(9),
        Z => S7(9)
    );
BUF_X1_796: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(90),
        Z => S7(90)
    );
BUF_X1_797: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(91),
        Z => S7(91)
    );
BUF_X1_798: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(92),
        Z => S7(92)
    );
BUF_X1_799: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(93),
        Z => S7(93)
    );
BUF_X1_800: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(94),
        Z => S7(94)
    );
BUF_X1_801: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(95),
        Z => S7(95)
    );
BUF_X1_802: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(96),
        Z => S7(96)
    );
BUF_X1_803: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(97),
        Z => S7(97)
    );
BUF_X1_804: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(98),
        Z => S7(98)
    );
BUF_X1_805: ENTITY WORK.BUF_X1
    PORT MAP (
        A => w(99),
        Z => S7(99)
    );
convergence_accumulator_plate_4_1: ENTITY WORK.convergence_accumulator_plate_4
    PORT MAP (
        clk => S0,
        din(0) => data_out_map_0,
        din(1) => data_out_map_1,
        din(2) => data_out_map_2,
        din(3) => data_out_map_3,
        din(4) => data_out_map_4,
        din(5) => data_out_map_5,
        din(6) => data_out_map_6,
        din(7) => data_out_map_7,
        din(8) => data_out_map_8,
        din(9) => data_out_map_9,
        din(10) => data_out_map_10,
        din(11) => data_out_map_11,
        din(12) => data_out_map_12,
        din(13) => data_out_map_13,
        din(14) => data_out_map_14,
        din(15) => data_out_map_15,
        din(16) => data_out_map_16,
        din(17) => data_out_map_17,
        din(18) => data_out_map_18,
        din(19) => data_out_map_19,
        din(20) => data_out_map_20,
        din(21) => data_out_map_21,
        din(22) => data_out_map_22,
        din(23) => data_out_map_23,
        din(24) => data_out_map_24,
        din(25) => data_out_map_25,
        din(26) => data_out_map_26,
        din(27) => data_out_map_27,
        din(28) => data_out_map_28,
        din(29) => data_out_map_29,
        din(30) => data_out_map_30,
        din(31) => data_out_map_31,
        din(32) => data_out_map_32,
        din(33) => data_out_map_33,
        din(34) => data_out_map_34,
        din(35) => data_out_map_35,
        din(36) => data_out_map_36,
        din(37) => data_out_map_37,
        din(38) => data_out_map_38,
        din(39) => data_out_map_39,
        din(40) => data_out_map_40,
        din(41) => data_out_map_41,
        din(42) => data_out_map_42,
        din(43) => data_out_map_43,
        din(44) => data_out_map_44,
        din(45) => data_out_map_45,
        din(46) => data_out_map_46,
        din(47) => data_out_map_47,
        din(48) => data_out_map_48,
        din(49) => data_out_map_49,
        din(50) => data_out_map_50,
        din(51) => data_out_map_51,
        din(52) => data_out_map_52,
        din(53) => data_out_map_53,
        din(54) => data_out_map_54,
        din(55) => data_out_map_55,
        din(56) => data_out_map_56,
        din(57) => data_out_map_57,
        din(58) => data_out_map_58,
        din(59) => data_out_map_59,
        din(60) => data_out_map_60,
        din(61) => data_out_map_61,
        din(62) => data_out_map_62,
        din(63) => data_out_map_63,
        din(64) => data_out_map_64,
        din(65) => data_out_map_65,
        din(66) => data_out_map_66,
        din(67) => data_out_map_67,
        din(68) => data_out_map_68,
        din(69) => data_out_map_69,
        din(70) => data_out_map_70,
        din(71) => data_out_map_71,
        din(72) => data_out_map_72,
        din(73) => data_out_map_73,
        din(74) => data_out_map_74,
        din(75) => data_out_map_75,
        din(76) => data_out_map_76,
        din(77) => data_out_map_77,
        din(78) => data_out_map_78,
        din(79) => data_out_map_79,
        din(80) => data_out_map_80,
        din(81) => data_out_map_81,
        din(82) => data_out_map_82,
        din(83) => data_out_map_83,
        din(84) => data_out_map_84,
        din(85) => data_out_map_85,
        din(86) => data_out_map_86,
        din(87) => data_out_map_87,
        din(88) => data_out_map_88,
        din(89) => data_out_map_89,
        din(90) => data_out_map_90,
        din(91) => data_out_map_91,
        din(92) => data_out_map_92,
        din(93) => data_out_map_93,
        din(94) => data_out_map_94,
        din(95) => data_out_map_95,
        din(96) => data_out_map_96,
        din(97) => data_out_map_97,
        din(98) => data_out_map_98,
        din(99) => data_out_map_99,
        din(100) => data_out_map_100,
        din(101) => data_out_map_101,
        din(102) => data_out_map_102,
        din(103) => data_out_map_103,
        din(104) => data_out_map_104,
        din(105) => data_out_map_105,
        din(106) => data_out_map_106,
        din(107) => data_out_map_107,
        din(108) => data_out_map_108,
        din(109) => data_out_map_109,
        din(110) => data_out_map_110,
        din(111) => data_out_map_111,
        din(112) => data_out_map_112,
        din(113) => data_out_map_113,
        din(114) => data_out_map_114,
        din(115) => data_out_map_115,
        din(116) => data_out_map_116,
        din(117) => data_out_map_117,
        din(118) => data_out_map_118,
        din(119) => data_out_map_119,
        din(120) => data_out_map_120,
        din(121) => data_out_map_121,
        din(122) => data_out_map_122,
        din(123) => data_out_map_123,
        din(124) => data_out_map_124,
        din(125) => data_out_map_125,
        din(126) => data_out_map_126,
        din(127) => data_out_map_127,
        dout(0) => S2(0),
        dout(1) => S2(1),
        dout(2) => S2(2),
        dout(3) => S2(3),
        dout(4) => S2(4),
        dout(5) => S2(5),
        dout(6) => S2(6),
        dout(7) => S2(7),
        dout(8) => S2(8),
        dout(9) => S2(9),
        dout(10) => S2(10),
        dout(11) => S2(11),
        dout(12) => S2(12),
        dout(13) => S2(13),
        dout(14) => S2(14),
        dout(15) => S2(15),
        dout(16) => S2(16),
        dout(17) => S2(17),
        dout(18) => S2(18),
        dout(19) => S2(19),
        dout(20) => S2(20),
        dout(21) => S2(21),
        dout(22) => S2(22),
        dout(23) => S2(23),
        dout(24) => S2(24),
        dout(25) => S2(25),
        dout(26) => S2(26),
        dout(27) => S2(27),
        dout(28) => S2(28),
        dout(29) => S2(29),
        dout(30) => S2(30),
        dout(31) => S2(31),
        reg_out => S4,
        rst => S5,
        run => hb0_map_ns_for:1_map_ns:4
    );
mapn_1_6_1_1_1_1_1_12_1: ENTITY WORK.mapn_1_6_1_1_1_1_1_12
    PORT MAP (
        clk => S0,
        din(0) => S1(0),
        din(1) => S1(1),
        din(2) => S1(2),
        din(3) => S1(3),
        din(4) => S1(4),
        din(5) => S1(5),
        din(6) => S1(6),
        din(7) => S1(7),
        din(8) => S1(8),
        din(9) => S1(9),
        din(10) => S1(10),
        din(11) => S1(11),
        din(12) => S1(12),
        din(13) => S1(13),
        din(14) => S1(14),
        din(15) => S1(15),
        din(16) => S1(16),
        din(17) => S1(17),
        din(18) => S1(18),
        din(19) => S1(19),
        din(20) => S1(20),
        din(21) => S1(21),
        din(22) => S1(22),
        din(23) => S1(23),
        din(24) => S1(24),
        din(25) => S1(25),
        din(26) => S1(26),
        din(27) => S1(27),
        din(28) => S1(28),
        din(29) => S1(29),
        din(30) => S1(30),
        din(31) => S1(31),
        din(32) => S1(32),
        din(33) => S1(33),
        din(34) => S1(34),
        din(35) => S1(35),
        din(36) => S1(36),
        din(37) => S1(37),
        din(38) => S1(38),
        din(39) => S1(39),
        din(40) => S1(40),
        din(41) => S1(41),
        din(42) => S1(42),
        din(43) => S1(43),
        din(44) => S1(44),
        din(45) => S1(45),
        din(46) => S1(46),
        din(47) => S1(47),
        din(48) => S1(48),
        din(49) => S1(49),
        din(50) => S1(50),
        din(51) => S1(51),
        din(52) => S1(52),
        din(53) => S1(53),
        din(54) => S1(54),
        din(55) => S1(55),
        din(56) => S1(56),
        din(57) => S1(57),
        din(58) => S1(58),
        din(59) => S1(59),
        din(60) => S1(60),
        din(61) => S1(61),
        din(62) => S1(62),
        din(63) => S1(63),
        din(64) => S1(64),
        din(65) => S1(65),
        din(66) => S1(66),
        din(67) => S1(67),
        din(68) => S1(68),
        din(69) => S1(69),
        din(70) => S1(70),
        din(71) => S1(71),
        din(72) => S1(72),
        din(73) => S1(73),
        din(74) => S1(74),
        din(75) => S1(75),
        din(76) => S1(76),
        din(77) => S1(77),
        din(78) => S1(78),
        din(79) => S1(79),
        din(80) => S1(80),
        din(81) => S1(81),
        din(82) => S1(82),
        din(83) => S1(83),
        din(84) => S1(84),
        din(85) => S1(85),
        din(86) => S1(86),
        din(87) => S1(87),
        din(88) => S1(88),
        din(89) => S1(89),
        din(90) => S1(90),
        din(91) => S1(91),
        din(92) => S1(92),
        din(93) => S1(93),
        din(94) => S1(94),
        din(95) => S1(95),
        dout(0) => data_out_map_0,
        dout(1) => data_out_map_1,
        dout(2) => data_out_map_2,
        dout(3) => data_out_map_3,
        dout(4) => data_out_map_4,
        dout(5) => data_out_map_5,
        dout(6) => data_out_map_6,
        dout(7) => data_out_map_7,
        dout(8) => data_out_map_8,
        dout(9) => data_out_map_9,
        dout(10) => data_out_map_10,
        dout(11) => data_out_map_11,
        dout(12) => data_out_map_12,
        dout(13) => data_out_map_13,
        dout(14) => data_out_map_14,
        dout(15) => data_out_map_15,
        dout(16) => data_out_map_16,
        dout(17) => data_out_map_17,
        dout(18) => data_out_map_18,
        dout(19) => data_out_map_19,
        dout(20) => data_out_map_20,
        dout(21) => data_out_map_21,
        dout(22) => data_out_map_22,
        dout(23) => data_out_map_23,
        dout(24) => data_out_map_24,
        dout(25) => data_out_map_25,
        dout(26) => data_out_map_26,
        dout(27) => data_out_map_27,
        dout(28) => data_out_map_28,
        dout(29) => data_out_map_29,
        dout(30) => data_out_map_30,
        dout(31) => data_out_map_31,
        pause => S3,
        reg_out => hb0_map_ns_for:1_map_ns:4,
        rst => S5,
        run => S6,
        w(0) => S7(0),
        w(1) => S7(1),
        w(2) => S7(2),
        w(3) => S7(3),
        w(4) => S7(4),
        w(5) => S7(5),
        w(6) => S7(6),
        w(7) => S7(7),
        w(8) => S7(8),
        w(9) => S7(9),
        w(10) => S7(10),
        w(11) => S7(11),
        w(12) => S7(12),
        w(13) => S7(13),
        w(14) => S7(14),
        w(15) => S7(15),
        w(16) => S7(16),
        w(17) => S7(17),
        w(18) => S7(18),
        w(19) => S7(19),
        w(20) => S7(20),
        w(21) => S7(21),
        w(22) => S7(22),
        w(23) => S7(23),
        w(24) => S7(24),
        w(25) => S7(25),
        w(26) => S7(26),
        w(27) => S7(27),
        w(28) => S7(28),
        w(29) => S7(29),
        w(30) => S7(30),
        w(31) => S7(31),
        w(32) => S7(32),
        w(33) => S7(33),
        w(34) => S7(34),
        w(35) => S7(35),
        w(36) => S7(36),
        w(37) => S7(37),
        w(38) => S7(38),
        w(39) => S7(39),
        w(40) => S7(40),
        w(41) => S7(41),
        w(42) => S7(42),
        w(43) => S7(43),
        w(44) => S7(44),
        w(45) => S7(45),
        w(46) => S7(46),
        w(47) => S7(47),
        w(48) => S7(48),
        w(49) => S7(49),
        w(50) => S7(50),
        w(51) => S7(51),
        w(52) => S7(52),
        w(53) => S7(53),
        w(54) => S7(54),
        w(55) => S7(55),
        w(56) => S7(56),
        w(57) => S7(57),
        w(58) => S7(58),
        w(59) => S7(59),
        w(60) => S7(60),
        w(61) => S7(61),
        w(62) => S7(62),
        w(63) => S7(63),
        w(64) => S7(64),
        w(65) => S7(65),
        w(66) => S7(66),
        w(67) => S7(67),
        w(68) => S7(68),
        w(69) => S7(69),
        w(70) => S7(70),
        w(71) => S7(71),
        w(72) => S7(72),
        w(73) => S7(73),
        w(74) => S7(74),
        w(75) => S7(75),
        w(76) => S7(76),
        w(77) => S7(77),
        w(78) => S7(78),
        w(79) => S7(79),
        w(80) => S7(80),
        w(81) => S7(81),
        w(82) => S7(82),
        w(83) => S7(83),
        w(84) => S7(84),
        w(85) => S7(85),
        w(86) => S7(86),
        w(87) => S7(87),
        w(88) => S7(88),
        w(89) => S7(89),
        w(90) => S7(90),
        w(91) => S7(91),
        w(92) => S7(92),
        w(93) => S7(93),
        w(94) => S7(94),
        w(95) => S7(95)
    );
mapn_1_6_1_1_1_1_1_12_2: ENTITY WORK.mapn_1_6_1_1_1_1_1_12
    PORT MAP (
        clk => S0,
        din(0) => S1(96),
        din(1) => S1(97),
        din(2) => S1(98),
        din(3) => S1(99),
        din(4) => S1(100),
        din(5) => S1(101),
        din(6) => S1(102),
        din(7) => S1(103),
        din(8) => S1(104),
        din(9) => S1(105),
        din(10) => S1(106),
        din(11) => S1(107),
        din(12) => S1(108),
        din(13) => S1(109),
        din(14) => S1(110),
        din(15) => S1(111),
        din(16) => S1(112),
        din(17) => S1(113),
        din(18) => S1(114),
        din(19) => S1(115),
        din(20) => S1(116),
        din(21) => S1(117),
        din(22) => S1(118),
        din(23) => S1(119),
        din(24) => S1(120),
        din(25) => S1(121),
        din(26) => S1(122),
        din(27) => S1(123),
        din(28) => S1(124),
        din(29) => S1(125),
        din(30) => S1(126),
        din(31) => S1(127),
        din(32) => S1(128),
        din(33) => S1(129),
        din(34) => S1(130),
        din(35) => S1(131),
        din(36) => S1(132),
        din(37) => S1(133),
        din(38) => S1(134),
        din(39) => S1(135),
        din(40) => S1(136),
        din(41) => S1(137),
        din(42) => S1(138),
        din(43) => S1(139),
        din(44) => S1(140),
        din(45) => S1(141),
        din(46) => S1(142),
        din(47) => S1(143),
        din(48) => S1(144),
        din(49) => S1(145),
        din(50) => S1(146),
        din(51) => S1(147),
        din(52) => S1(148),
        din(53) => S1(149),
        din(54) => S1(150),
        din(55) => S1(151),
        din(56) => S1(152),
        din(57) => S1(153),
        din(58) => S1(154),
        din(59) => S1(155),
        din(60) => S1(156),
        din(61) => S1(157),
        din(62) => S1(158),
        din(63) => S1(159),
        din(64) => S1(160),
        din(65) => S1(161),
        din(66) => S1(162),
        din(67) => S1(163),
        din(68) => S1(164),
        din(69) => S1(165),
        din(70) => S1(166),
        din(71) => S1(167),
        din(72) => S1(168),
        din(73) => S1(169),
        din(74) => S1(170),
        din(75) => S1(171),
        din(76) => S1(172),
        din(77) => S1(173),
        din(78) => S1(174),
        din(79) => S1(175),
        din(80) => S1(176),
        din(81) => S1(177),
        din(82) => S1(178),
        din(83) => S1(179),
        din(84) => S1(180),
        din(85) => S1(181),
        din(86) => S1(182),
        din(87) => S1(183),
        din(88) => S1(184),
        din(89) => S1(185),
        din(90) => S1(186),
        din(91) => S1(187),
        din(92) => S1(188),
        din(93) => S1(189),
        din(94) => S1(190),
        din(95) => S1(191),
        dout(0) => data_out_map_32,
        dout(1) => data_out_map_33,
        dout(2) => data_out_map_34,
        dout(3) => data_out_map_35,
        dout(4) => data_out_map_36,
        dout(5) => data_out_map_37,
        dout(6) => data_out_map_38,
        dout(7) => data_out_map_39,
        dout(8) => data_out_map_40,
        dout(9) => data_out_map_41,
        dout(10) => data_out_map_42,
        dout(11) => data_out_map_43,
        dout(12) => data_out_map_44,
        dout(13) => data_out_map_45,
        dout(14) => data_out_map_46,
        dout(15) => data_out_map_47,
        dout(16) => data_out_map_48,
        dout(17) => data_out_map_49,
        dout(18) => data_out_map_50,
        dout(19) => data_out_map_51,
        dout(20) => data_out_map_52,
        dout(21) => data_out_map_53,
        dout(22) => data_out_map_54,
        dout(23) => data_out_map_55,
        dout(24) => data_out_map_56,
        dout(25) => data_out_map_57,
        dout(26) => data_out_map_58,
        dout(27) => data_out_map_59,
        dout(28) => data_out_map_60,
        dout(29) => data_out_map_61,
        dout(30) => data_out_map_62,
        dout(31) => data_out_map_63,
        pause => S3,
        reg_out => hb0_map_ns_for:2_map_ns:13,
        rst => S5,
        run => S6,
        w(0) => S7(96),
        w(1) => S7(97),
        w(2) => S7(98),
        w(3) => S7(99),
        w(4) => S7(100),
        w(5) => S7(101),
        w(6) => S7(102),
        w(7) => S7(103),
        w(8) => S7(104),
        w(9) => S7(105),
        w(10) => S7(106),
        w(11) => S7(107),
        w(12) => S7(108),
        w(13) => S7(109),
        w(14) => S7(110),
        w(15) => S7(111),
        w(16) => S7(112),
        w(17) => S7(113),
        w(18) => S7(114),
        w(19) => S7(115),
        w(20) => S7(116),
        w(21) => S7(117),
        w(22) => S7(118),
        w(23) => S7(119),
        w(24) => S7(120),
        w(25) => S7(121),
        w(26) => S7(122),
        w(27) => S7(123),
        w(28) => S7(124),
        w(29) => S7(125),
        w(30) => S7(126),
        w(31) => S7(127),
        w(32) => S7(128),
        w(33) => S7(129),
        w(34) => S7(130),
        w(35) => S7(131),
        w(36) => S7(132),
        w(37) => S7(133),
        w(38) => S7(134),
        w(39) => S7(135),
        w(40) => S7(136),
        w(41) => S7(137),
        w(42) => S7(138),
        w(43) => S7(139),
        w(44) => S7(140),
        w(45) => S7(141),
        w(46) => S7(142),
        w(47) => S7(143),
        w(48) => S7(144),
        w(49) => S7(145),
        w(50) => S7(146),
        w(51) => S7(147),
        w(52) => S7(148),
        w(53) => S7(149),
        w(54) => S7(150),
        w(55) => S7(151),
        w(56) => S7(152),
        w(57) => S7(153),
        w(58) => S7(154),
        w(59) => S7(155),
        w(60) => S7(156),
        w(61) => S7(157),
        w(62) => S7(158),
        w(63) => S7(159),
        w(64) => S7(160),
        w(65) => S7(161),
        w(66) => S7(162),
        w(67) => S7(163),
        w(68) => S7(164),
        w(69) => S7(165),
        w(70) => S7(166),
        w(71) => S7(167),
        w(72) => S7(168),
        w(73) => S7(169),
        w(74) => S7(170),
        w(75) => S7(171),
        w(76) => S7(172),
        w(77) => S7(173),
        w(78) => S7(174),
        w(79) => S7(175),
        w(80) => S7(176),
        w(81) => S7(177),
        w(82) => S7(178),
        w(83) => S7(179),
        w(84) => S7(180),
        w(85) => S7(181),
        w(86) => S7(182),
        w(87) => S7(183),
        w(88) => S7(184),
        w(89) => S7(185),
        w(90) => S7(186),
        w(91) => S7(187),
        w(92) => S7(188),
        w(93) => S7(189),
        w(94) => S7(190),
        w(95) => S7(191)
    );
mapn_1_6_1_1_1_1_1_12_3: ENTITY WORK.mapn_1_6_1_1_1_1_1_12
    PORT MAP (
        clk => S0,
        din(0) => S1(192),
        din(1) => S1(193),
        din(2) => S1(194),
        din(3) => S1(195),
        din(4) => S1(196),
        din(5) => S1(197),
        din(6) => S1(198),
        din(7) => S1(199),
        din(8) => S1(200),
        din(9) => S1(201),
        din(10) => S1(202),
        din(11) => S1(203),
        din(12) => S1(204),
        din(13) => S1(205),
        din(14) => S1(206),
        din(15) => S1(207),
        din(16) => S1(208),
        din(17) => S1(209),
        din(18) => S1(210),
        din(19) => S1(211),
        din(20) => S1(212),
        din(21) => S1(213),
        din(22) => S1(214),
        din(23) => S1(215),
        din(24) => S1(216),
        din(25) => S1(217),
        din(26) => S1(218),
        din(27) => S1(219),
        din(28) => S1(220),
        din(29) => S1(221),
        din(30) => S1(222),
        din(31) => S1(223),
        din(32) => S1(224),
        din(33) => S1(225),
        din(34) => S1(226),
        din(35) => S1(227),
        din(36) => S1(228),
        din(37) => S1(229),
        din(38) => S1(230),
        din(39) => S1(231),
        din(40) => S1(232),
        din(41) => S1(233),
        din(42) => S1(234),
        din(43) => S1(235),
        din(44) => S1(236),
        din(45) => S1(237),
        din(46) => S1(238),
        din(47) => S1(239),
        din(48) => S1(240),
        din(49) => S1(241),
        din(50) => S1(242),
        din(51) => S1(243),
        din(52) => S1(244),
        din(53) => S1(245),
        din(54) => S1(246),
        din(55) => S1(247),
        din(56) => S1(248),
        din(57) => S1(249),
        din(58) => S1(250),
        din(59) => S1(251),
        din(60) => S1(252),
        din(61) => S1(253),
        din(62) => S1(254),
        din(63) => S1(255),
        din(64) => S1(256),
        din(65) => S1(257),
        din(66) => S1(258),
        din(67) => S1(259),
        din(68) => S1(260),
        din(69) => S1(261),
        din(70) => S1(262),
        din(71) => S1(263),
        din(72) => S1(264),
        din(73) => S1(265),
        din(74) => S1(266),
        din(75) => S1(267),
        din(76) => S1(268),
        din(77) => S1(269),
        din(78) => S1(270),
        din(79) => S1(271),
        din(80) => S1(272),
        din(81) => S1(273),
        din(82) => S1(274),
        din(83) => S1(275),
        din(84) => S1(276),
        din(85) => S1(277),
        din(86) => S1(278),
        din(87) => S1(279),
        din(88) => S1(280),
        din(89) => S1(281),
        din(90) => S1(282),
        din(91) => S1(283),
        din(92) => S1(284),
        din(93) => S1(285),
        din(94) => S1(286),
        din(95) => S1(287),
        dout(0) => data_out_map_64,
        dout(1) => data_out_map_65,
        dout(2) => data_out_map_66,
        dout(3) => data_out_map_67,
        dout(4) => data_out_map_68,
        dout(5) => data_out_map_69,
        dout(6) => data_out_map_70,
        dout(7) => data_out_map_71,
        dout(8) => data_out_map_72,
        dout(9) => data_out_map_73,
        dout(10) => data_out_map_74,
        dout(11) => data_out_map_75,
        dout(12) => data_out_map_76,
        dout(13) => data_out_map_77,
        dout(14) => data_out_map_78,
        dout(15) => data_out_map_79,
        dout(16) => data_out_map_80,
        dout(17) => data_out_map_81,
        dout(18) => data_out_map_82,
        dout(19) => data_out_map_83,
        dout(20) => data_out_map_84,
        dout(21) => data_out_map_85,
        dout(22) => data_out_map_86,
        dout(23) => data_out_map_87,
        dout(24) => data_out_map_88,
        dout(25) => data_out_map_89,
        dout(26) => data_out_map_90,
        dout(27) => data_out_map_91,
        dout(28) => data_out_map_92,
        dout(29) => data_out_map_93,
        dout(30) => data_out_map_94,
        dout(31) => data_out_map_95,
        pause => S3,
        reg_out => hb0_map_ns_for:3_map_ns:22,
        rst => S5,
        run => S6,
        w(0) => S7(192),
        w(1) => S7(193),
        w(2) => S7(194),
        w(3) => S7(195),
        w(4) => S7(196),
        w(5) => S7(197),
        w(6) => S7(198),
        w(7) => S7(199),
        w(8) => S7(200),
        w(9) => S7(201),
        w(10) => S7(202),
        w(11) => S7(203),
        w(12) => S7(204),
        w(13) => S7(205),
        w(14) => S7(206),
        w(15) => S7(207),
        w(16) => S7(208),
        w(17) => S7(209),
        w(18) => S7(210),
        w(19) => S7(211),
        w(20) => S7(212),
        w(21) => S7(213),
        w(22) => S7(214),
        w(23) => S7(215),
        w(24) => S7(216),
        w(25) => S7(217),
        w(26) => S7(218),
        w(27) => S7(219),
        w(28) => S7(220),
        w(29) => S7(221),
        w(30) => S7(222),
        w(31) => S7(223),
        w(32) => S7(224),
        w(33) => S7(225),
        w(34) => S7(226),
        w(35) => S7(227),
        w(36) => S7(228),
        w(37) => S7(229),
        w(38) => S7(230),
        w(39) => S7(231),
        w(40) => S7(232),
        w(41) => S7(233),
        w(42) => S7(234),
        w(43) => S7(235),
        w(44) => S7(236),
        w(45) => S7(237),
        w(46) => S7(238),
        w(47) => S7(239),
        w(48) => S7(240),
        w(49) => S7(241),
        w(50) => S7(242),
        w(51) => S7(243),
        w(52) => S7(244),
        w(53) => S7(245),
        w(54) => S7(246),
        w(55) => S7(247),
        w(56) => S7(248),
        w(57) => S7(249),
        w(58) => S7(250),
        w(59) => S7(251),
        w(60) => S7(252),
        w(61) => S7(253),
        w(62) => S7(254),
        w(63) => S7(255),
        w(64) => S7(256),
        w(65) => S7(257),
        w(66) => S7(258),
        w(67) => S7(259),
        w(68) => S7(260),
        w(69) => S7(261),
        w(70) => S7(262),
        w(71) => S7(263),
        w(72) => S7(264),
        w(73) => S7(265),
        w(74) => S7(266),
        w(75) => S7(267),
        w(76) => S7(268),
        w(77) => S7(269),
        w(78) => S7(270),
        w(79) => S7(271),
        w(80) => S7(272),
        w(81) => S7(273),
        w(82) => S7(274),
        w(83) => S7(275),
        w(84) => S7(276),
        w(85) => S7(277),
        w(86) => S7(278),
        w(87) => S7(279),
        w(88) => S7(280),
        w(89) => S7(281),
        w(90) => S7(282),
        w(91) => S7(283),
        w(92) => S7(284),
        w(93) => S7(285),
        w(94) => S7(286),
        w(95) => S7(287)
    );
mapn_1_6_1_1_1_1_1_12_4: ENTITY WORK.mapn_1_6_1_1_1_1_1_12
    PORT MAP (
        clk => S0,
        din(0) => S1(288),
        din(1) => S1(289),
        din(2) => S1(290),
        din(3) => S1(291),
        din(4) => S1(292),
        din(5) => S1(293),
        din(6) => S1(294),
        din(7) => S1(295),
        din(8) => S1(296),
        din(9) => S1(297),
        din(10) => S1(298),
        din(11) => S1(299),
        din(12) => S1(300),
        din(13) => S1(301),
        din(14) => S1(302),
        din(15) => S1(303),
        din(16) => S1(304),
        din(17) => S1(305),
        din(18) => S1(306),
        din(19) => S1(307),
        din(20) => S1(308),
        din(21) => S1(309),
        din(22) => S1(310),
        din(23) => S1(311),
        din(24) => S1(312),
        din(25) => S1(313),
        din(26) => S1(314),
        din(27) => S1(315),
        din(28) => S1(316),
        din(29) => S1(317),
        din(30) => S1(318),
        din(31) => S1(319),
        din(32) => S1(320),
        din(33) => S1(321),
        din(34) => S1(322),
        din(35) => S1(323),
        din(36) => S1(324),
        din(37) => S1(325),
        din(38) => S1(326),
        din(39) => S1(327),
        din(40) => S1(328),
        din(41) => S1(329),
        din(42) => S1(330),
        din(43) => S1(331),
        din(44) => S1(332),
        din(45) => S1(333),
        din(46) => S1(334),
        din(47) => S1(335),
        din(48) => S1(336),
        din(49) => S1(337),
        din(50) => S1(338),
        din(51) => S1(339),
        din(52) => S1(340),
        din(53) => S1(341),
        din(54) => S1(342),
        din(55) => S1(343),
        din(56) => S1(344),
        din(57) => S1(345),
        din(58) => S1(346),
        din(59) => S1(347),
        din(60) => S1(348),
        din(61) => S1(349),
        din(62) => S1(350),
        din(63) => S1(351),
        din(64) => S1(352),
        din(65) => S1(353),
        din(66) => S1(354),
        din(67) => S1(355),
        din(68) => S1(356),
        din(69) => S1(357),
        din(70) => S1(358),
        din(71) => S1(359),
        din(72) => S1(360),
        din(73) => S1(361),
        din(74) => S1(362),
        din(75) => S1(363),
        din(76) => S1(364),
        din(77) => S1(365),
        din(78) => S1(366),
        din(79) => S1(367),
        din(80) => S1(368),
        din(81) => S1(369),
        din(82) => S1(370),
        din(83) => S1(371),
        din(84) => S1(372),
        din(85) => S1(373),
        din(86) => S1(374),
        din(87) => S1(375),
        din(88) => S1(376),
        din(89) => S1(377),
        din(90) => S1(378),
        din(91) => S1(379),
        din(92) => S1(380),
        din(93) => S1(381),
        din(94) => S1(382),
        din(95) => S1(383),
        dout(0) => data_out_map_96,
        dout(1) => data_out_map_97,
        dout(2) => data_out_map_98,
        dout(3) => data_out_map_99,
        dout(4) => data_out_map_100,
        dout(5) => data_out_map_101,
        dout(6) => data_out_map_102,
        dout(7) => data_out_map_103,
        dout(8) => data_out_map_104,
        dout(9) => data_out_map_105,
        dout(10) => data_out_map_106,
        dout(11) => data_out_map_107,
        dout(12) => data_out_map_108,
        dout(13) => data_out_map_109,
        dout(14) => data_out_map_110,
        dout(15) => data_out_map_111,
        dout(16) => data_out_map_112,
        dout(17) => data_out_map_113,
        dout(18) => data_out_map_114,
        dout(19) => data_out_map_115,
        dout(20) => data_out_map_116,
        dout(21) => data_out_map_117,
        dout(22) => data_out_map_118,
        dout(23) => data_out_map_119,
        dout(24) => data_out_map_120,
        dout(25) => data_out_map_121,
        dout(26) => data_out_map_122,
        dout(27) => data_out_map_123,
        dout(28) => data_out_map_124,
        dout(29) => data_out_map_125,
        dout(30) => data_out_map_126,
        dout(31) => data_out_map_127,
        pause => S3,
        reg_out => hb0_map_ns_for:4_map_ns:31,
        rst => S5,
        run => S6,
        w(0) => S7(288),
        w(1) => S7(289),
        w(2) => S7(290),
        w(3) => S7(291),
        w(4) => S7(292),
        w(5) => S7(293),
        w(6) => S7(294),
        w(7) => S7(295),
        w(8) => S7(296),
        w(9) => S7(297),
        w(10) => S7(298),
        w(11) => S7(299),
        w(12) => S7(300),
        w(13) => S7(301),
        w(14) => S7(302),
        w(15) => S7(303),
        w(16) => S7(304),
        w(17) => S7(305),
        w(18) => S7(306),
        w(19) => S7(307),
        w(20) => S7(308),
        w(21) => S7(309),
        w(22) => S7(310),
        w(23) => S7(311),
        w(24) => S7(312),
        w(25) => S7(313),
        w(26) => S7(314),
        w(27) => S7(315),
        w(28) => S7(316),
        w(29) => S7(317),
        w(30) => S7(318),
        w(31) => S7(319),
        w(32) => S7(320),
        w(33) => S7(321),
        w(34) => S7(322),
        w(35) => S7(323),
        w(36) => S7(324),
        w(37) => S7(325),
        w(38) => S7(326),
        w(39) => S7(327),
        w(40) => S7(328),
        w(41) => S7(329),
        w(42) => S7(330),
        w(43) => S7(331),
        w(44) => S7(332),
        w(45) => S7(333),
        w(46) => S7(334),
        w(47) => S7(335),
        w(48) => S7(336),
        w(49) => S7(337),
        w(50) => S7(338),
        w(51) => S7(339),
        w(52) => S7(340),
        w(53) => S7(341),
        w(54) => S7(342),
        w(55) => S7(343),
        w(56) => S7(344),
        w(57) => S7(345),
        w(58) => S7(346),
        w(59) => S7(347),
        w(60) => S7(348),
        w(61) => S7(349),
        w(62) => S7(350),
        w(63) => S7(351),
        w(64) => S7(352),
        w(65) => S7(353),
        w(66) => S7(354),
        w(67) => S7(355),
        w(68) => S7(356),
        w(69) => S7(357),
        w(70) => S7(358),
        w(71) => S7(359),
        w(72) => S7(360),
        w(73) => S7(361),
        w(74) => S7(362),
        w(75) => S7(363),
        w(76) => S7(364),
        w(77) => S7(365),
        w(78) => S7(366),
        w(79) => S7(367),
        w(80) => S7(368),
        w(81) => S7(369),
        w(82) => S7(370),
        w(83) => S7(371),
        w(84) => S7(372),
        w(85) => S7(373),
        w(86) => S7(374),
        w(87) => S7(375),
        w(88) => S7(376),
        w(89) => S7(377),
        w(90) => S7(378),
        w(91) => S7(379),
        w(92) => S7(380),
        w(93) => S7(381),
        w(94) => S7(382),
        w(95) => S7(383)
    );

END ARCHITECTURE arch;
